MACRO r2r_dac
  CLASS BLOCK ;
  FOREIGN r2r_dac ;
  ORIGIN -5.000 27.290 ;
  SIZE 13.860 BY 26.330 ;
  PIN out
    PORT
      LAYER met1 ;
        RECT 5.200 -20.400 6.200 -19.400 ;
    END
  END out
  PIN vdd
    ANTENNADIFFAREA 29.199598 ;
    PORT
      LAYER met1 ;
        RECT 7.930 -1.960 8.930 -0.960 ;
    END
  END vdd
  PIN b0
    ANTENNAGATEAREA 1.200000 ;
    PORT
      LAYER met1 ;
        RECT 16.870 -10.170 17.870 -9.170 ;
    END
  END b0
  PIN b1
    ANTENNAGATEAREA 1.200000 ;
    PORT
      LAYER met1 ;
        RECT 15.210 -10.120 16.210 -9.120 ;
    END
  END b1
  PIN b2
    ANTENNAGATEAREA 1.200000 ;
    PORT
      LAYER met1 ;
        RECT 13.640 -10.120 14.640 -9.120 ;
    END
  END b2
  PIN b3
    ANTENNAGATEAREA 1.200000 ;
    PORT
      LAYER met1 ;
        RECT 12.020 -10.090 13.020 -9.090 ;
    END
  END b3
  PIN b4
    ANTENNAGATEAREA 1.200000 ;
    PORT
      LAYER met1 ;
        RECT 10.470 -10.120 11.470 -9.120 ;
    END
  END b4
  PIN b5
    ANTENNAGATEAREA 1.200000 ;
    PORT
      LAYER met1 ;
        RECT 8.860 -10.090 9.860 -9.090 ;
    END
  END b5
  PIN b6
    ANTENNAGATEAREA 1.200000 ;
    PORT
      LAYER met1 ;
        RECT 7.350 -10.120 8.350 -9.120 ;
    END
  END b6
  PIN b7
    ANTENNAGATEAREA 1.200000 ;
    PORT
      LAYER met1 ;
        RECT 5.850 -10.100 6.850 -9.100 ;
    END
  END b7
  PIN vss
    ANTENNADIFFAREA 39.098999 ;
    PORT
      LAYER met1 ;
        RECT 5.200 -14.400 6.200 -13.400 ;
    END
  END vss
  OBS
      LAYER nwell ;
        RECT 5.000 -9.310 18.170 -1.470 ;
      LAYER pwell ;
        RECT 5.010 -13.810 18.180 -10.020 ;
        RECT 5.010 -21.300 18.860 -14.080 ;
        RECT 5.010 -27.290 15.900 -21.300 ;
      LAYER li1 ;
        RECT 5.230 -1.650 17.940 -1.040 ;
        RECT 5.180 -1.850 17.990 -1.650 ;
        RECT 5.180 -8.960 5.350 -1.850 ;
        RECT 5.750 -8.230 5.920 -2.190 ;
        RECT 6.190 -8.230 6.360 -2.190 ;
        RECT 5.890 -8.615 6.220 -8.445 ;
        RECT 6.760 -8.960 6.930 -1.850 ;
        RECT 7.330 -8.230 7.500 -2.190 ;
        RECT 7.770 -8.230 7.940 -2.190 ;
        RECT 7.470 -8.615 7.800 -8.445 ;
        RECT 8.340 -8.960 8.510 -1.850 ;
        RECT 8.910 -8.230 9.080 -2.190 ;
        RECT 9.350 -8.230 9.520 -2.190 ;
        RECT 9.050 -8.615 9.380 -8.445 ;
        RECT 9.920 -8.960 10.090 -1.850 ;
        RECT 10.490 -8.230 10.660 -2.190 ;
        RECT 10.930 -8.230 11.100 -2.190 ;
        RECT 10.630 -8.615 10.960 -8.445 ;
        RECT 11.500 -8.960 11.670 -1.850 ;
        RECT 12.070 -8.230 12.240 -2.190 ;
        RECT 12.510 -8.230 12.680 -2.190 ;
        RECT 12.210 -8.615 12.540 -8.445 ;
        RECT 13.080 -8.960 13.250 -1.850 ;
        RECT 13.650 -8.230 13.820 -2.190 ;
        RECT 14.090 -8.230 14.260 -2.190 ;
        RECT 13.790 -8.615 14.120 -8.445 ;
        RECT 14.660 -8.960 14.830 -1.850 ;
        RECT 15.230 -8.230 15.400 -2.190 ;
        RECT 15.670 -8.230 15.840 -2.190 ;
        RECT 15.370 -8.615 15.700 -8.445 ;
        RECT 16.240 -8.960 16.410 -1.850 ;
        RECT 16.810 -8.230 16.980 -2.190 ;
        RECT 17.250 -8.230 17.420 -2.190 ;
        RECT 16.950 -8.615 17.280 -8.445 ;
        RECT 17.820 -8.960 17.990 -1.850 ;
        RECT 5.180 -9.130 17.990 -8.960 ;
        RECT 5.190 -10.370 18.000 -10.200 ;
        RECT 5.190 -13.440 5.360 -10.370 ;
        RECT 5.900 -10.880 6.230 -10.710 ;
        RECT 5.760 -13.090 5.930 -11.050 ;
        RECT 6.200 -13.090 6.370 -11.050 ;
        RECT 6.770 -13.440 6.940 -10.370 ;
        RECT 7.480 -10.880 7.810 -10.710 ;
        RECT 7.340 -13.090 7.510 -11.050 ;
        RECT 7.780 -13.090 7.950 -11.050 ;
        RECT 8.350 -13.440 8.520 -10.370 ;
        RECT 9.060 -10.880 9.390 -10.710 ;
        RECT 8.920 -13.090 9.090 -11.050 ;
        RECT 9.360 -13.090 9.530 -11.050 ;
        RECT 9.930 -13.440 10.100 -10.370 ;
        RECT 10.640 -10.880 10.970 -10.710 ;
        RECT 10.500 -13.090 10.670 -11.050 ;
        RECT 10.940 -13.090 11.110 -11.050 ;
        RECT 11.510 -13.440 11.680 -10.370 ;
        RECT 12.220 -10.880 12.550 -10.710 ;
        RECT 12.080 -13.090 12.250 -11.050 ;
        RECT 12.520 -13.090 12.690 -11.050 ;
        RECT 13.090 -13.440 13.260 -10.370 ;
        RECT 13.800 -10.880 14.130 -10.710 ;
        RECT 13.660 -13.090 13.830 -11.050 ;
        RECT 14.100 -13.090 14.270 -11.050 ;
        RECT 14.670 -13.440 14.840 -10.370 ;
        RECT 15.380 -10.880 15.710 -10.710 ;
        RECT 15.240 -13.090 15.410 -11.050 ;
        RECT 15.680 -13.090 15.850 -11.050 ;
        RECT 16.250 -13.440 16.420 -10.370 ;
        RECT 16.960 -10.880 17.290 -10.710 ;
        RECT 16.820 -13.090 16.990 -11.050 ;
        RECT 17.260 -13.090 17.430 -11.050 ;
        RECT 17.830 -13.440 18.000 -10.370 ;
        RECT 5.190 -13.630 18.000 -13.440 ;
        RECT 5.270 -14.260 17.960 -13.630 ;
        RECT 5.190 -14.430 18.680 -14.260 ;
        RECT 5.190 -20.950 5.360 -14.430 ;
        RECT 5.840 -17.070 6.190 -14.910 ;
        RECT 5.840 -20.470 6.190 -18.310 ;
        RECT 6.670 -20.950 6.840 -14.430 ;
        RECT 7.320 -17.070 7.670 -14.910 ;
        RECT 7.320 -20.470 7.670 -18.310 ;
        RECT 8.150 -20.950 8.320 -14.430 ;
        RECT 8.800 -17.070 9.150 -14.910 ;
        RECT 8.800 -20.470 9.150 -18.310 ;
        RECT 9.630 -20.950 9.800 -14.430 ;
        RECT 10.280 -17.070 10.630 -14.910 ;
        RECT 10.280 -20.470 10.630 -18.310 ;
        RECT 11.110 -20.950 11.280 -14.430 ;
        RECT 11.760 -17.070 12.110 -14.910 ;
        RECT 11.760 -20.470 12.110 -18.310 ;
        RECT 12.590 -20.950 12.760 -14.430 ;
        RECT 13.240 -17.070 13.590 -14.910 ;
        RECT 13.240 -20.470 13.590 -18.310 ;
        RECT 14.070 -20.950 14.240 -14.430 ;
        RECT 14.720 -17.070 15.070 -14.910 ;
        RECT 14.720 -20.470 15.070 -18.310 ;
        RECT 15.550 -20.950 15.720 -14.430 ;
        RECT 16.200 -17.070 16.550 -14.910 ;
        RECT 16.200 -20.470 16.550 -18.310 ;
        RECT 17.030 -20.950 17.200 -14.430 ;
        RECT 17.680 -17.070 18.030 -14.910 ;
        RECT 17.680 -20.470 18.030 -18.310 ;
        RECT 18.510 -20.950 18.680 -14.430 ;
        RECT 5.190 -21.120 18.680 -20.950 ;
        RECT 5.190 -26.940 5.360 -21.120 ;
        RECT 5.840 -23.760 6.190 -21.600 ;
        RECT 5.840 -26.460 6.190 -24.300 ;
        RECT 6.670 -26.940 6.840 -21.120 ;
        RECT 7.320 -23.760 7.670 -21.600 ;
        RECT 7.320 -26.460 7.670 -24.300 ;
        RECT 8.150 -26.940 8.320 -21.120 ;
        RECT 8.800 -23.760 9.150 -21.600 ;
        RECT 8.800 -26.460 9.150 -24.300 ;
        RECT 9.630 -26.940 9.800 -21.120 ;
        RECT 10.280 -23.760 10.630 -21.600 ;
        RECT 10.280 -26.460 10.630 -24.300 ;
        RECT 11.110 -26.940 11.280 -21.120 ;
        RECT 11.760 -23.760 12.110 -21.600 ;
        RECT 11.760 -26.460 12.110 -24.300 ;
        RECT 12.590 -26.940 12.760 -21.120 ;
        RECT 13.240 -23.760 13.590 -21.600 ;
        RECT 13.240 -26.460 13.590 -24.300 ;
        RECT 14.070 -26.940 14.240 -21.120 ;
        RECT 14.720 -23.760 15.070 -21.600 ;
        RECT 14.720 -26.460 15.070 -24.300 ;
        RECT 15.550 -26.940 15.720 -21.120 ;
        RECT 5.190 -27.110 15.720 -26.940 ;
      LAYER met1 ;
        RECT 5.190 -0.980 7.930 -0.960 ;
        RECT 5.170 -1.790 7.930 -0.980 ;
        RECT 5.190 -1.850 7.930 -1.790 ;
        RECT 8.930 -0.980 18.000 -0.960 ;
        RECT 8.930 -1.790 18.010 -0.980 ;
        RECT 8.930 -1.850 18.000 -1.790 ;
        RECT 6.190 -2.210 6.630 -1.850 ;
        RECT 7.770 -1.960 7.930 -1.850 ;
        RECT 7.770 -2.210 8.210 -1.960 ;
        RECT 9.360 -2.210 9.800 -1.850 ;
        RECT 10.950 -2.210 11.390 -1.850 ;
        RECT 5.330 -2.260 5.560 -2.230 ;
        RECT 5.720 -2.260 5.950 -2.210 ;
        RECT 5.330 -8.150 5.950 -2.260 ;
        RECT 5.330 -8.430 5.570 -8.150 ;
        RECT 5.720 -8.210 5.950 -8.150 ;
        RECT 6.160 -8.150 6.630 -2.210 ;
        RECT 7.300 -2.280 7.530 -2.210 ;
        RECT 7.000 -8.130 7.530 -2.280 ;
        RECT 7.000 -8.150 7.160 -8.130 ;
        RECT 6.160 -8.210 6.390 -8.150 ;
        RECT 7.010 -8.390 7.160 -8.150 ;
        RECT 7.300 -8.210 7.530 -8.130 ;
        RECT 7.740 -8.130 8.210 -2.210 ;
        RECT 8.880 -2.280 9.110 -2.210 ;
        RECT 8.510 -6.870 9.120 -2.280 ;
        RECT 7.740 -8.210 7.970 -8.130 ;
        RECT 8.490 -8.160 9.120 -6.870 ;
        RECT 9.320 -8.120 9.800 -2.210 ;
        RECT 10.460 -2.260 10.690 -2.210 ;
        RECT 5.330 -10.860 5.710 -8.430 ;
        RECT 5.910 -8.440 6.200 -8.415 ;
        RECT 5.900 -9.100 6.220 -8.440 ;
        RECT 5.850 -10.170 6.850 -10.100 ;
        RECT 5.900 -10.860 6.220 -10.170 ;
        RECT 5.330 -11.170 5.570 -10.860 ;
        RECT 5.920 -10.900 6.220 -10.860 ;
        RECT 5.920 -10.910 6.210 -10.900 ;
        RECT 7.010 -10.920 7.210 -8.390 ;
        RECT 7.490 -8.420 7.780 -8.415 ;
        RECT 7.480 -9.120 7.820 -8.420 ;
        RECT 7.480 -10.890 7.820 -10.120 ;
        RECT 7.500 -10.910 7.790 -10.890 ;
        RECT 5.730 -11.170 5.960 -11.070 ;
        RECT 5.330 -11.180 5.960 -11.170 ;
        RECT 5.300 -12.980 5.960 -11.180 ;
        RECT 5.330 -13.000 5.560 -12.980 ;
        RECT 5.730 -13.070 5.960 -12.980 ;
        RECT 6.170 -11.140 6.400 -11.070 ;
        RECT 6.170 -12.950 6.730 -11.140 ;
        RECT 7.010 -11.180 7.160 -10.920 ;
        RECT 7.310 -11.180 7.540 -11.070 ;
        RECT 7.010 -11.190 7.540 -11.180 ;
        RECT 6.170 -13.070 6.400 -12.950 ;
        RECT 6.560 -13.270 6.730 -12.950 ;
        RECT 6.970 -12.990 7.540 -11.190 ;
        RECT 7.020 -13.000 7.540 -12.990 ;
        RECT 7.310 -13.070 7.540 -13.000 ;
        RECT 7.750 -11.120 7.980 -11.070 ;
        RECT 7.750 -11.150 8.260 -11.120 ;
        RECT 7.750 -12.960 8.290 -11.150 ;
        RECT 8.490 -11.170 8.680 -8.160 ;
        RECT 8.880 -8.210 9.110 -8.160 ;
        RECT 9.320 -8.210 9.550 -8.120 ;
        RECT 10.070 -8.160 10.690 -2.260 ;
        RECT 9.040 -9.090 9.400 -8.410 ;
        RECT 8.860 -10.120 9.860 -10.090 ;
        RECT 9.040 -10.910 9.400 -10.120 ;
        RECT 8.890 -11.170 9.120 -11.070 ;
        RECT 8.490 -11.840 9.120 -11.170 ;
        RECT 7.750 -13.070 7.980 -12.960 ;
        RECT 8.120 -13.190 8.290 -12.960 ;
        RECT 8.510 -13.040 9.120 -11.840 ;
        RECT 8.890 -13.070 9.120 -13.040 ;
        RECT 9.330 -11.120 9.560 -11.070 ;
        RECT 9.330 -13.000 9.870 -11.120 ;
        RECT 10.090 -11.140 10.260 -8.160 ;
        RECT 10.460 -8.210 10.690 -8.160 ;
        RECT 10.900 -8.130 11.390 -2.210 ;
        RECT 12.040 -2.290 12.270 -2.210 ;
        RECT 10.900 -8.210 11.130 -8.130 ;
        RECT 11.630 -8.170 12.270 -2.290 ;
        RECT 10.650 -8.420 10.940 -8.415 ;
        RECT 10.640 -9.090 10.980 -8.420 ;
        RECT 10.470 -9.120 11.470 -9.090 ;
        RECT 10.640 -10.900 10.980 -10.120 ;
        RECT 10.660 -10.910 10.950 -10.900 ;
        RECT 10.470 -11.140 10.700 -11.070 ;
        RECT 10.090 -11.180 10.700 -11.140 ;
        RECT 10.070 -12.980 10.700 -11.180 ;
        RECT 10.100 -13.000 10.700 -12.980 ;
        RECT 9.330 -13.070 9.560 -13.000 ;
        RECT 6.480 -13.410 6.730 -13.270 ;
        RECT 8.110 -13.410 8.290 -13.190 ;
        RECT 9.700 -13.240 9.870 -13.000 ;
        RECT 10.470 -13.070 10.700 -13.000 ;
        RECT 10.910 -11.140 11.140 -11.070 ;
        RECT 10.910 -13.020 11.450 -11.140 ;
        RECT 11.640 -11.150 11.830 -8.170 ;
        RECT 12.040 -8.210 12.270 -8.170 ;
        RECT 12.470 -8.180 12.910 -1.850 ;
        RECT 14.090 -2.210 14.530 -1.850 ;
        RECT 15.680 -2.210 16.120 -1.850 ;
        RECT 17.260 -2.210 17.700 -1.850 ;
        RECT 13.620 -2.230 13.850 -2.210 ;
        RECT 13.170 -8.160 13.850 -2.230 ;
        RECT 12.480 -8.210 12.710 -8.180 ;
        RECT 12.230 -8.420 12.520 -8.415 ;
        RECT 12.210 -9.090 12.570 -8.420 ;
        RECT 12.020 -10.120 13.020 -10.090 ;
        RECT 12.210 -10.910 12.570 -10.120 ;
        RECT 12.050 -11.150 12.280 -11.070 ;
        RECT 11.640 -13.000 12.280 -11.150 ;
        RECT 10.910 -13.070 11.140 -13.020 ;
        RECT 9.690 -13.410 9.870 -13.240 ;
        RECT 11.280 -13.410 11.450 -13.020 ;
        RECT 12.050 -13.070 12.280 -13.000 ;
        RECT 12.490 -11.120 12.720 -11.070 ;
        RECT 13.180 -11.110 13.440 -8.160 ;
        RECT 13.620 -8.210 13.850 -8.160 ;
        RECT 14.060 -8.150 14.530 -2.210 ;
        RECT 15.200 -2.250 15.430 -2.210 ;
        RECT 14.060 -8.210 14.290 -8.150 ;
        RECT 14.750 -8.160 15.430 -2.250 ;
        RECT 13.810 -8.420 14.100 -8.415 ;
        RECT 13.780 -9.090 14.120 -8.420 ;
        RECT 13.640 -9.120 14.640 -9.090 ;
        RECT 13.780 -10.910 14.120 -10.120 ;
        RECT 13.630 -11.110 13.860 -11.070 ;
        RECT 12.490 -13.000 13.030 -11.120 ;
        RECT 12.490 -13.070 12.720 -13.000 ;
        RECT 12.860 -13.410 13.030 -13.000 ;
        RECT 13.180 -13.030 13.860 -11.110 ;
        RECT 13.630 -13.070 13.860 -13.030 ;
        RECT 14.070 -11.130 14.300 -11.070 ;
        RECT 14.070 -13.010 14.620 -11.130 ;
        RECT 14.800 -11.150 15.060 -8.160 ;
        RECT 15.200 -8.210 15.430 -8.160 ;
        RECT 15.640 -8.170 16.120 -2.210 ;
        RECT 16.780 -2.250 17.010 -2.210 ;
        RECT 16.350 -8.140 17.010 -2.250 ;
        RECT 16.350 -8.160 16.610 -8.140 ;
        RECT 15.640 -8.210 15.870 -8.170 ;
        RECT 16.360 -8.370 16.610 -8.160 ;
        RECT 16.780 -8.210 17.010 -8.140 ;
        RECT 17.220 -8.120 17.700 -2.210 ;
        RECT 17.220 -8.210 17.450 -8.120 ;
        RECT 15.390 -8.420 15.680 -8.415 ;
        RECT 15.380 -9.120 15.710 -8.420 ;
        RECT 15.380 -10.910 15.710 -10.120 ;
        RECT 16.360 -10.470 16.660 -8.370 ;
        RECT 16.970 -8.420 17.260 -8.415 ;
        RECT 16.950 -9.100 17.310 -8.420 ;
        RECT 16.870 -9.170 17.870 -9.100 ;
        RECT 16.440 -10.920 16.660 -10.470 ;
        RECT 16.950 -10.910 17.310 -10.170 ;
        RECT 15.210 -11.150 15.440 -11.070 ;
        RECT 14.780 -13.000 15.440 -11.150 ;
        RECT 14.070 -13.070 14.300 -13.010 ;
        RECT 14.460 -13.410 14.620 -13.010 ;
        RECT 15.210 -13.070 15.440 -13.000 ;
        RECT 15.650 -11.130 15.880 -11.070 ;
        RECT 15.650 -13.020 16.200 -11.130 ;
        RECT 16.440 -11.160 16.620 -10.920 ;
        RECT 16.790 -11.160 17.020 -11.070 ;
        RECT 16.440 -11.310 17.020 -11.160 ;
        RECT 16.410 -12.980 17.020 -11.310 ;
        RECT 16.420 -13.010 17.020 -12.980 ;
        RECT 15.650 -13.070 15.880 -13.020 ;
        RECT 16.030 -13.410 16.200 -13.020 ;
        RECT 16.790 -13.070 17.020 -13.010 ;
        RECT 17.230 -11.130 17.460 -11.070 ;
        RECT 17.230 -12.980 17.920 -11.130 ;
        RECT 17.230 -13.070 17.460 -12.980 ;
        RECT 17.610 -13.230 17.920 -12.980 ;
        RECT 17.590 -13.270 17.920 -13.230 ;
        RECT 17.590 -13.410 18.080 -13.270 ;
        RECT 5.180 -14.400 5.200 -13.440 ;
        RECT 6.200 -14.400 18.080 -13.410 ;
        RECT 5.180 -14.430 18.080 -14.400 ;
        RECT 5.200 -14.470 18.080 -14.430 ;
        RECT 5.740 -17.150 6.350 -14.810 ;
        RECT 7.180 -15.000 7.840 -14.680 ;
        RECT 7.230 -17.120 7.840 -15.000 ;
        RECT 7.680 -17.150 7.840 -17.120 ;
        RECT 8.700 -17.160 9.250 -14.810 ;
        RECT 10.210 -17.180 10.760 -14.830 ;
        RECT 11.670 -17.150 12.220 -14.800 ;
        RECT 13.150 -17.120 13.700 -14.770 ;
        RECT 14.600 -17.130 15.150 -14.780 ;
        RECT 16.100 -17.120 16.650 -14.770 ;
        RECT 17.520 -14.910 18.080 -14.470 ;
        RECT 17.520 -17.070 18.090 -14.910 ;
        RECT 17.520 -17.080 18.080 -17.070 ;
        RECT 5.180 -18.330 5.570 -18.320 ;
        RECT 5.180 -19.400 6.200 -18.330 ;
        RECT 5.180 -20.400 5.200 -19.400 ;
        RECT 5.180 -20.490 6.200 -20.400 ;
        RECT 5.180 -24.310 5.570 -20.490 ;
        RECT 6.660 -20.730 7.660 -18.330 ;
        RECT 8.150 -20.460 9.150 -18.310 ;
        RECT 6.410 -20.960 7.660 -20.730 ;
        RECT 5.850 -21.120 7.660 -20.960 ;
        RECT 7.920 -21.100 9.150 -20.460 ;
        RECT 9.630 -20.470 10.630 -18.320 ;
        RECT 11.090 -20.470 12.090 -18.330 ;
        RECT 5.850 -21.420 7.130 -21.120 ;
        RECT 5.850 -23.300 6.850 -21.420 ;
        RECT 7.920 -21.570 8.600 -21.100 ;
        RECT 9.410 -21.110 10.630 -20.470 ;
        RECT 9.410 -21.570 10.090 -21.110 ;
        RECT 10.900 -21.120 12.090 -20.470 ;
        RECT 12.590 -20.500 13.590 -18.310 ;
        RECT 15.530 -18.330 17.840 -18.320 ;
        RECT 12.350 -21.100 13.590 -20.500 ;
        RECT 14.100 -20.510 15.100 -18.330 ;
        RECT 15.530 -20.500 18.010 -18.330 ;
        RECT 10.900 -21.570 11.580 -21.120 ;
        RECT 12.350 -21.570 13.030 -21.100 ;
        RECT 7.300 -22.040 8.600 -21.570 ;
        RECT 7.300 -23.210 8.340 -22.040 ;
        RECT 8.810 -22.050 10.090 -21.570 ;
        RECT 10.280 -22.050 11.580 -21.570 ;
        RECT 8.810 -23.210 9.850 -22.050 ;
        RECT 10.280 -23.210 11.320 -22.050 ;
        RECT 11.770 -22.080 13.030 -21.570 ;
        RECT 13.850 -21.120 15.100 -20.510 ;
        RECT 15.360 -21.110 18.010 -20.500 ;
        RECT 13.850 -21.580 14.530 -21.120 ;
        RECT 15.360 -21.570 16.040 -21.110 ;
        RECT 17.010 -21.120 18.010 -21.110 ;
        RECT 5.850 -23.750 7.080 -23.300 ;
        RECT 7.300 -23.750 8.630 -23.210 ;
        RECT 8.810 -23.750 10.120 -23.210 ;
        RECT 10.280 -23.750 11.610 -23.210 ;
        RECT 11.770 -23.220 12.810 -22.080 ;
        RECT 13.250 -22.090 14.530 -21.580 ;
        RECT 14.730 -22.080 16.040 -21.570 ;
        RECT 13.250 -23.220 14.290 -22.090 ;
        RECT 11.770 -23.750 13.040 -23.220 ;
        RECT 6.400 -24.310 7.080 -23.750 ;
        RECT 7.950 -24.300 8.630 -23.750 ;
        RECT 9.440 -24.290 10.120 -23.750 ;
        RECT 10.930 -24.290 11.610 -23.750 ;
        RECT 12.360 -24.290 13.040 -23.750 ;
        RECT 13.250 -23.760 14.550 -23.220 ;
        RECT 14.730 -23.750 15.770 -22.080 ;
        RECT 13.870 -24.290 14.550 -23.760 ;
        RECT 5.180 -26.460 6.200 -24.310 ;
        RECT 6.400 -24.880 7.710 -24.310 ;
        RECT 7.950 -24.790 9.160 -24.300 ;
        RECT 9.440 -24.790 10.670 -24.290 ;
        RECT 10.930 -24.790 12.140 -24.290 ;
        RECT 6.670 -26.470 7.710 -24.880 ;
        RECT 8.120 -26.480 9.160 -24.790 ;
        RECT 9.630 -26.470 10.670 -24.790 ;
        RECT 11.100 -26.470 12.140 -24.790 ;
        RECT 12.360 -24.800 13.630 -24.290 ;
        RECT 13.870 -24.800 15.100 -24.290 ;
        RECT 12.590 -26.470 13.630 -24.800 ;
        RECT 14.060 -26.470 15.100 -24.800 ;
      LAYER met2 ;
        RECT 5.350 -12.000 5.670 -11.130 ;
        RECT 5.340 -13.030 5.670 -12.000 ;
        RECT 7.020 -12.020 7.340 -11.140 ;
        RECT 5.340 -14.790 5.650 -13.030 ;
        RECT 7.000 -13.040 7.340 -12.020 ;
        RECT 8.580 -13.040 8.900 -11.140 ;
        RECT 10.120 -12.030 10.440 -11.130 ;
        RECT 10.100 -13.030 10.440 -12.030 ;
        RECT 11.710 -12.220 12.030 -11.110 ;
        RECT 7.000 -14.680 7.310 -13.040 ;
        RECT 5.340 -14.950 5.560 -14.790 ;
        RECT 5.810 -14.950 6.350 -14.810 ;
        RECT 5.340 -17.040 6.350 -14.950 ;
        RECT 5.380 -17.060 6.350 -17.040 ;
        RECT 7.000 -15.000 7.810 -14.680 ;
        RECT 8.580 -14.810 8.890 -13.040 ;
        RECT 7.000 -17.060 7.730 -15.000 ;
        RECT 5.740 -17.150 6.350 -17.060 ;
        RECT 7.280 -17.090 7.730 -17.060 ;
        RECT 7.310 -17.120 7.680 -17.090 ;
        RECT 8.580 -17.100 9.250 -14.810 ;
        RECT 10.100 -14.830 10.410 -13.030 ;
        RECT 11.670 -14.800 12.040 -12.220 ;
        RECT 13.270 -12.230 13.590 -11.140 ;
        RECT 14.860 -12.190 15.180 -11.120 ;
        RECT 16.460 -11.880 16.740 -11.130 ;
        RECT 13.250 -14.770 13.620 -12.230 ;
        RECT 10.100 -17.070 10.760 -14.830 ;
        RECT 8.700 -17.160 9.250 -17.100 ;
        RECT 10.210 -17.180 10.760 -17.070 ;
        RECT 11.670 -17.150 12.220 -14.800 ;
        RECT 13.150 -17.120 13.700 -14.770 ;
        RECT 14.860 -14.780 15.210 -12.190 ;
        RECT 16.440 -14.770 16.740 -11.880 ;
        RECT 14.600 -17.030 15.210 -14.780 ;
        RECT 14.600 -17.130 15.150 -17.030 ;
        RECT 16.100 -17.060 16.740 -14.770 ;
        RECT 16.100 -17.120 16.650 -17.060 ;
  END
END r2r_dac
END LIBRARY

