VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_tim2305_adc_dac
  CLASS BLOCK ;
  FOREIGN tt_um_tim2305_adc_dac ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 13.475 211.915 13.645 212.105 ;
        RECT 14.855 211.915 15.025 212.105 ;
        RECT 20.375 211.915 20.545 212.105 ;
        RECT 25.890 211.965 26.010 212.075 ;
        RECT 26.815 211.915 26.985 212.105 ;
        RECT 32.335 211.915 32.505 212.105 ;
        RECT 37.855 211.915 38.025 212.105 ;
        RECT 39.695 211.915 39.865 212.105 ;
        RECT 45.215 211.915 45.385 212.105 ;
        RECT 50.735 211.915 50.905 212.105 ;
        RECT 52.575 211.915 52.745 212.105 ;
        RECT 58.095 211.915 58.265 212.105 ;
        RECT 63.615 211.915 63.785 212.105 ;
        RECT 65.455 211.915 65.625 212.105 ;
        RECT 70.975 211.915 71.145 212.105 ;
        RECT 74.195 211.915 74.365 212.105 ;
        RECT 74.655 211.915 74.825 212.105 ;
        RECT 77.410 211.965 77.530 212.075 ;
        RECT 78.335 211.915 78.505 212.105 ;
        RECT 83.855 211.915 84.025 212.105 ;
        RECT 89.375 211.915 89.545 212.105 ;
        RECT 91.215 211.915 91.385 212.105 ;
        RECT 96.735 211.915 96.905 212.105 ;
        RECT 102.255 211.915 102.425 212.105 ;
        RECT 104.095 211.915 104.265 212.105 ;
        RECT 109.615 211.915 109.785 212.105 ;
        RECT 115.135 211.915 115.305 212.105 ;
        RECT 116.975 211.915 117.145 212.105 ;
        RECT 122.495 211.915 122.665 212.105 ;
        RECT 128.015 211.915 128.185 212.105 ;
        RECT 129.855 211.915 130.025 212.105 ;
        RECT 135.375 211.915 135.545 212.105 ;
        RECT 137.210 211.965 137.330 212.075 ;
        RECT 138.595 211.915 138.765 212.105 ;
        RECT 13.335 211.105 14.705 211.915 ;
        RECT 14.715 211.105 20.225 211.915 ;
        RECT 20.235 211.105 25.745 211.915 ;
        RECT 26.225 211.045 26.655 211.830 ;
        RECT 26.675 211.105 32.185 211.915 ;
        RECT 32.195 211.105 37.705 211.915 ;
        RECT 37.715 211.105 39.085 211.915 ;
        RECT 39.105 211.045 39.535 211.830 ;
        RECT 39.555 211.105 45.065 211.915 ;
        RECT 45.075 211.105 50.585 211.915 ;
        RECT 50.595 211.105 51.965 211.915 ;
        RECT 51.985 211.045 52.415 211.830 ;
        RECT 52.435 211.105 57.945 211.915 ;
        RECT 57.955 211.105 63.465 211.915 ;
        RECT 63.475 211.105 64.845 211.915 ;
        RECT 64.865 211.045 65.295 211.830 ;
        RECT 65.315 211.105 70.825 211.915 ;
        RECT 70.835 211.105 72.665 211.915 ;
        RECT 72.675 211.235 74.505 211.915 ;
        RECT 72.675 211.005 74.020 211.235 ;
        RECT 74.515 211.105 77.265 211.915 ;
        RECT 77.745 211.045 78.175 211.830 ;
        RECT 78.195 211.105 83.705 211.915 ;
        RECT 83.715 211.105 89.225 211.915 ;
        RECT 89.235 211.105 90.605 211.915 ;
        RECT 90.625 211.045 91.055 211.830 ;
        RECT 91.075 211.105 96.585 211.915 ;
        RECT 96.595 211.105 102.105 211.915 ;
        RECT 102.115 211.105 103.485 211.915 ;
        RECT 103.505 211.045 103.935 211.830 ;
        RECT 103.955 211.105 109.465 211.915 ;
        RECT 109.475 211.105 114.985 211.915 ;
        RECT 114.995 211.105 116.365 211.915 ;
        RECT 116.385 211.045 116.815 211.830 ;
        RECT 116.835 211.105 122.345 211.915 ;
        RECT 122.355 211.105 127.865 211.915 ;
        RECT 127.875 211.105 129.245 211.915 ;
        RECT 129.265 211.045 129.695 211.830 ;
        RECT 129.715 211.105 135.225 211.915 ;
        RECT 135.235 211.105 137.065 211.915 ;
        RECT 137.535 211.105 138.905 211.915 ;
      LAYER nwell ;
        RECT 13.140 207.885 139.100 210.715 ;
      LAYER pwell ;
        RECT 13.335 206.685 14.705 207.495 ;
        RECT 14.715 206.685 20.225 207.495 ;
        RECT 20.235 206.685 25.745 207.495 ;
        RECT 26.225 206.770 26.655 207.555 ;
        RECT 26.675 206.685 32.185 207.495 ;
        RECT 32.195 206.685 37.705 207.495 ;
        RECT 37.715 206.685 43.225 207.495 ;
        RECT 43.235 206.685 48.745 207.495 ;
        RECT 48.755 206.685 51.505 207.495 ;
        RECT 51.985 206.770 52.415 207.555 ;
        RECT 52.435 206.685 57.945 207.495 ;
        RECT 57.955 206.685 63.465 207.495 ;
        RECT 63.475 206.685 68.985 207.495 ;
        RECT 68.995 206.685 74.505 207.495 ;
        RECT 74.515 206.685 77.265 207.495 ;
        RECT 77.745 206.770 78.175 207.555 ;
        RECT 78.195 206.685 83.705 207.495 ;
        RECT 83.715 206.685 89.225 207.495 ;
        RECT 89.235 206.685 94.745 207.495 ;
        RECT 94.755 206.685 100.265 207.495 ;
        RECT 100.275 206.685 103.025 207.495 ;
        RECT 103.505 206.770 103.935 207.555 ;
        RECT 103.955 206.685 109.465 207.495 ;
        RECT 109.475 206.685 114.985 207.495 ;
        RECT 114.995 206.685 120.505 207.495 ;
        RECT 120.515 206.685 126.025 207.495 ;
        RECT 126.035 206.685 128.785 207.495 ;
        RECT 129.265 206.770 129.695 207.555 ;
        RECT 129.715 206.685 135.225 207.495 ;
        RECT 135.235 206.685 137.065 207.495 ;
        RECT 137.535 206.685 138.905 207.495 ;
        RECT 13.475 206.475 13.645 206.685 ;
        RECT 14.855 206.475 15.025 206.685 ;
        RECT 20.375 206.475 20.545 206.685 ;
        RECT 25.895 206.635 26.065 206.665 ;
        RECT 25.890 206.525 26.065 206.635 ;
        RECT 25.895 206.475 26.065 206.525 ;
        RECT 26.815 206.495 26.985 206.685 ;
        RECT 31.415 206.475 31.585 206.665 ;
        RECT 32.335 206.495 32.505 206.685 ;
        RECT 36.935 206.475 37.105 206.665 ;
        RECT 37.855 206.495 38.025 206.685 ;
        RECT 38.770 206.525 38.890 206.635 ;
        RECT 39.695 206.475 39.865 206.665 ;
        RECT 43.375 206.495 43.545 206.685 ;
        RECT 45.215 206.475 45.385 206.665 ;
        RECT 48.895 206.495 49.065 206.685 ;
        RECT 50.735 206.475 50.905 206.665 ;
        RECT 51.650 206.525 51.770 206.635 ;
        RECT 52.575 206.495 52.745 206.685 ;
        RECT 56.255 206.475 56.425 206.665 ;
        RECT 58.095 206.495 58.265 206.685 ;
        RECT 61.775 206.475 61.945 206.665 ;
        RECT 63.615 206.495 63.785 206.685 ;
        RECT 64.530 206.525 64.650 206.635 ;
        RECT 65.455 206.475 65.625 206.665 ;
        RECT 69.135 206.495 69.305 206.685 ;
        RECT 70.975 206.475 71.145 206.665 ;
        RECT 74.655 206.495 74.825 206.685 ;
        RECT 76.495 206.475 76.665 206.665 ;
        RECT 77.410 206.525 77.530 206.635 ;
        RECT 78.335 206.495 78.505 206.685 ;
        RECT 82.015 206.475 82.185 206.665 ;
        RECT 83.855 206.495 84.025 206.685 ;
        RECT 87.535 206.475 87.705 206.665 ;
        RECT 89.375 206.495 89.545 206.685 ;
        RECT 90.290 206.525 90.410 206.635 ;
        RECT 91.215 206.475 91.385 206.665 ;
        RECT 94.895 206.495 95.065 206.685 ;
        RECT 96.735 206.475 96.905 206.665 ;
        RECT 100.415 206.495 100.585 206.685 ;
        RECT 102.255 206.475 102.425 206.665 ;
        RECT 103.170 206.525 103.290 206.635 ;
        RECT 104.095 206.495 104.265 206.685 ;
        RECT 107.775 206.475 107.945 206.665 ;
        RECT 109.615 206.495 109.785 206.685 ;
        RECT 113.295 206.475 113.465 206.665 ;
        RECT 115.135 206.495 115.305 206.685 ;
        RECT 116.050 206.525 116.170 206.635 ;
        RECT 116.975 206.475 117.145 206.665 ;
        RECT 120.655 206.495 120.825 206.685 ;
        RECT 122.495 206.475 122.665 206.665 ;
        RECT 126.175 206.495 126.345 206.685 ;
        RECT 128.015 206.475 128.185 206.665 ;
        RECT 128.930 206.525 129.050 206.635 ;
        RECT 129.855 206.495 130.025 206.685 ;
        RECT 133.535 206.475 133.705 206.665 ;
        RECT 135.375 206.495 135.545 206.685 ;
        RECT 137.210 206.525 137.330 206.635 ;
        RECT 138.595 206.475 138.765 206.685 ;
        RECT 13.335 205.665 14.705 206.475 ;
        RECT 14.715 205.665 20.225 206.475 ;
        RECT 20.235 205.665 25.745 206.475 ;
        RECT 25.755 205.665 31.265 206.475 ;
        RECT 31.275 205.665 36.785 206.475 ;
        RECT 36.795 205.665 38.625 206.475 ;
        RECT 39.105 205.605 39.535 206.390 ;
        RECT 39.555 205.665 45.065 206.475 ;
        RECT 45.075 205.665 50.585 206.475 ;
        RECT 50.595 205.665 56.105 206.475 ;
        RECT 56.115 205.665 61.625 206.475 ;
        RECT 61.635 205.665 64.385 206.475 ;
        RECT 64.865 205.605 65.295 206.390 ;
        RECT 65.315 205.665 70.825 206.475 ;
        RECT 70.835 205.665 76.345 206.475 ;
        RECT 76.355 205.665 81.865 206.475 ;
        RECT 81.875 205.665 87.385 206.475 ;
        RECT 87.395 205.665 90.145 206.475 ;
        RECT 90.625 205.605 91.055 206.390 ;
        RECT 91.075 205.665 96.585 206.475 ;
        RECT 96.595 205.665 102.105 206.475 ;
        RECT 102.115 205.665 107.625 206.475 ;
        RECT 107.635 205.665 113.145 206.475 ;
        RECT 113.155 205.665 115.905 206.475 ;
        RECT 116.385 205.605 116.815 206.390 ;
        RECT 116.835 205.665 122.345 206.475 ;
        RECT 122.355 205.665 127.865 206.475 ;
        RECT 127.875 205.665 133.385 206.475 ;
        RECT 133.395 205.665 137.065 206.475 ;
        RECT 137.535 205.665 138.905 206.475 ;
      LAYER nwell ;
        RECT 13.140 202.445 139.100 205.275 ;
      LAYER pwell ;
        RECT 13.335 201.245 14.705 202.055 ;
        RECT 14.715 201.245 20.225 202.055 ;
        RECT 20.235 201.245 25.745 202.055 ;
        RECT 26.225 201.330 26.655 202.115 ;
        RECT 26.675 201.245 32.185 202.055 ;
        RECT 32.195 201.245 37.705 202.055 ;
        RECT 37.715 201.245 43.225 202.055 ;
        RECT 43.235 201.245 48.745 202.055 ;
        RECT 48.755 201.245 51.505 202.055 ;
        RECT 51.985 201.330 52.415 202.115 ;
        RECT 52.435 201.245 57.945 202.055 ;
        RECT 57.955 201.245 63.465 202.055 ;
        RECT 63.475 201.245 68.985 202.055 ;
        RECT 68.995 201.245 74.505 202.055 ;
        RECT 74.515 201.245 77.265 202.055 ;
        RECT 77.745 201.330 78.175 202.115 ;
        RECT 78.195 201.245 83.705 202.055 ;
        RECT 83.715 201.245 89.225 202.055 ;
        RECT 89.235 201.245 94.745 202.055 ;
        RECT 94.755 201.245 100.265 202.055 ;
        RECT 100.275 201.245 103.025 202.055 ;
        RECT 103.505 201.330 103.935 202.115 ;
        RECT 103.955 201.245 109.465 202.055 ;
        RECT 109.475 201.245 114.985 202.055 ;
        RECT 114.995 201.245 120.505 202.055 ;
        RECT 120.515 201.245 126.025 202.055 ;
        RECT 126.035 201.245 128.785 202.055 ;
        RECT 129.265 201.330 129.695 202.115 ;
        RECT 129.715 201.245 135.225 202.055 ;
        RECT 135.235 201.245 137.065 202.055 ;
        RECT 137.535 201.245 138.905 202.055 ;
        RECT 13.475 201.035 13.645 201.245 ;
        RECT 14.855 201.035 15.025 201.245 ;
        RECT 20.375 201.035 20.545 201.245 ;
        RECT 25.895 201.195 26.065 201.225 ;
        RECT 25.890 201.085 26.065 201.195 ;
        RECT 25.895 201.035 26.065 201.085 ;
        RECT 26.815 201.055 26.985 201.245 ;
        RECT 31.415 201.035 31.585 201.225 ;
        RECT 32.335 201.055 32.505 201.245 ;
        RECT 36.935 201.035 37.105 201.225 ;
        RECT 37.855 201.055 38.025 201.245 ;
        RECT 38.770 201.085 38.890 201.195 ;
        RECT 39.695 201.035 39.865 201.225 ;
        RECT 43.375 201.055 43.545 201.245 ;
        RECT 45.215 201.035 45.385 201.225 ;
        RECT 48.895 201.055 49.065 201.245 ;
        RECT 50.735 201.035 50.905 201.225 ;
        RECT 51.650 201.085 51.770 201.195 ;
        RECT 52.575 201.055 52.745 201.245 ;
        RECT 56.255 201.035 56.425 201.225 ;
        RECT 58.095 201.055 58.265 201.245 ;
        RECT 61.775 201.035 61.945 201.225 ;
        RECT 63.615 201.055 63.785 201.245 ;
        RECT 64.075 201.035 64.245 201.225 ;
        RECT 64.530 201.085 64.650 201.195 ;
        RECT 66.375 201.035 66.545 201.225 ;
        RECT 66.835 201.035 67.005 201.225 ;
        RECT 69.135 201.055 69.305 201.245 ;
        RECT 74.655 201.055 74.825 201.245 ;
        RECT 77.415 201.195 77.585 201.225 ;
        RECT 77.410 201.085 77.585 201.195 ;
        RECT 77.415 201.035 77.585 201.085 ;
        RECT 78.335 201.055 78.505 201.245 ;
        RECT 80.175 201.035 80.345 201.225 ;
        RECT 80.635 201.035 80.805 201.225 ;
        RECT 83.855 201.055 84.025 201.245 ;
        RECT 86.155 201.035 86.325 201.225 ;
        RECT 89.375 201.055 89.545 201.245 ;
        RECT 89.845 201.080 90.005 201.190 ;
        RECT 91.215 201.035 91.385 201.225 ;
        RECT 94.895 201.055 95.065 201.245 ;
        RECT 96.735 201.035 96.905 201.225 ;
        RECT 100.415 201.055 100.585 201.245 ;
        RECT 102.255 201.035 102.425 201.225 ;
        RECT 103.170 201.085 103.290 201.195 ;
        RECT 104.095 201.055 104.265 201.245 ;
        RECT 107.775 201.035 107.945 201.225 ;
        RECT 109.615 201.055 109.785 201.245 ;
        RECT 114.675 201.035 114.845 201.225 ;
        RECT 115.135 201.035 115.305 201.245 ;
        RECT 116.975 201.035 117.145 201.225 ;
        RECT 120.655 201.055 120.825 201.245 ;
        RECT 122.495 201.035 122.665 201.225 ;
        RECT 126.175 201.055 126.345 201.245 ;
        RECT 128.015 201.035 128.185 201.225 ;
        RECT 128.930 201.085 129.050 201.195 ;
        RECT 129.855 201.055 130.025 201.245 ;
        RECT 133.535 201.035 133.705 201.225 ;
        RECT 135.375 201.055 135.545 201.245 ;
        RECT 137.210 201.085 137.330 201.195 ;
        RECT 138.595 201.035 138.765 201.245 ;
        RECT 13.335 200.225 14.705 201.035 ;
        RECT 14.715 200.225 20.225 201.035 ;
        RECT 20.235 200.225 25.745 201.035 ;
        RECT 25.755 200.225 31.265 201.035 ;
        RECT 31.275 200.225 36.785 201.035 ;
        RECT 36.795 200.225 38.625 201.035 ;
        RECT 39.105 200.165 39.535 200.950 ;
        RECT 39.555 200.225 45.065 201.035 ;
        RECT 45.075 200.225 50.585 201.035 ;
        RECT 50.595 200.225 56.105 201.035 ;
        RECT 56.115 200.225 61.625 201.035 ;
        RECT 61.635 200.225 63.005 201.035 ;
        RECT 63.015 200.255 64.385 201.035 ;
        RECT 64.865 200.165 65.295 200.950 ;
        RECT 65.325 200.125 66.675 201.035 ;
        RECT 66.695 200.355 74.005 201.035 ;
        RECT 70.210 200.135 71.120 200.355 ;
        RECT 72.655 200.125 74.005 200.355 ;
        RECT 74.150 200.355 77.615 201.035 ;
        RECT 77.745 200.355 80.485 201.035 ;
        RECT 74.150 200.125 75.070 200.355 ;
        RECT 80.495 200.225 86.005 201.035 ;
        RECT 86.015 200.225 89.685 201.035 ;
        RECT 90.625 200.165 91.055 200.950 ;
        RECT 91.075 200.225 96.585 201.035 ;
        RECT 96.595 200.225 102.105 201.035 ;
        RECT 102.115 200.225 107.625 201.035 ;
        RECT 107.635 200.225 113.145 201.035 ;
        RECT 113.155 200.355 114.985 201.035 ;
        RECT 113.155 200.125 114.500 200.355 ;
        RECT 114.995 200.225 116.365 201.035 ;
        RECT 116.385 200.165 116.815 200.950 ;
        RECT 116.835 200.225 122.345 201.035 ;
        RECT 122.355 200.225 127.865 201.035 ;
        RECT 127.875 200.225 133.385 201.035 ;
        RECT 133.395 200.225 137.065 201.035 ;
        RECT 137.535 200.225 138.905 201.035 ;
      LAYER nwell ;
        RECT 13.140 197.005 139.100 199.835 ;
      LAYER pwell ;
        RECT 13.335 195.805 14.705 196.615 ;
        RECT 14.715 195.805 20.225 196.615 ;
        RECT 20.235 195.805 25.745 196.615 ;
        RECT 26.225 195.890 26.655 196.675 ;
        RECT 26.675 195.805 32.185 196.615 ;
        RECT 32.195 195.805 37.705 196.615 ;
        RECT 37.715 195.805 43.225 196.615 ;
        RECT 43.235 195.805 48.745 196.615 ;
        RECT 48.755 195.805 51.505 196.615 ;
        RECT 51.985 195.890 52.415 196.675 ;
        RECT 52.435 195.805 57.945 196.615 ;
        RECT 57.955 195.805 60.705 196.615 ;
        RECT 61.270 196.485 62.190 196.715 ;
        RECT 61.270 195.805 64.735 196.485 ;
        RECT 65.795 195.805 67.145 196.715 ;
        RECT 67.255 195.805 70.365 196.715 ;
        RECT 73.890 196.485 74.800 196.705 ;
        RECT 76.335 196.485 77.685 196.715 ;
        RECT 70.375 195.805 77.685 196.485 ;
        RECT 77.745 195.890 78.175 196.675 ;
        RECT 79.245 196.485 80.175 196.715 ;
        RECT 78.340 195.805 80.175 196.485 ;
        RECT 80.495 195.805 86.005 196.615 ;
        RECT 86.015 195.805 88.765 196.615 ;
        RECT 89.255 195.805 90.605 196.715 ;
        RECT 91.575 196.485 92.925 196.715 ;
        RECT 94.460 196.485 95.370 196.705 ;
        RECT 91.575 195.805 98.885 196.485 ;
        RECT 98.895 195.805 101.185 196.715 ;
        RECT 101.195 195.805 103.025 196.715 ;
        RECT 103.505 195.890 103.935 196.675 ;
        RECT 103.955 195.805 107.625 196.615 ;
        RECT 108.595 196.485 109.945 196.715 ;
        RECT 111.480 196.485 112.390 196.705 ;
        RECT 115.955 196.485 117.305 196.715 ;
        RECT 118.840 196.485 119.750 196.705 ;
        RECT 108.595 195.805 115.905 196.485 ;
        RECT 115.955 195.805 123.265 196.485 ;
        RECT 123.275 195.805 128.785 196.615 ;
        RECT 129.265 195.890 129.695 196.675 ;
        RECT 129.715 195.805 135.225 196.615 ;
        RECT 135.235 195.805 137.065 196.615 ;
        RECT 137.535 195.805 138.905 196.615 ;
        RECT 13.475 195.595 13.645 195.805 ;
        RECT 14.855 195.595 15.025 195.805 ;
        RECT 20.375 195.595 20.545 195.805 ;
        RECT 25.895 195.755 26.065 195.785 ;
        RECT 25.890 195.645 26.065 195.755 ;
        RECT 25.895 195.595 26.065 195.645 ;
        RECT 26.815 195.615 26.985 195.805 ;
        RECT 31.425 195.640 31.585 195.750 ;
        RECT 32.335 195.595 32.505 195.805 ;
        RECT 36.015 195.595 36.185 195.785 ;
        RECT 37.855 195.615 38.025 195.805 ;
        RECT 38.770 195.645 38.890 195.755 ;
        RECT 39.695 195.595 39.865 195.785 ;
        RECT 43.375 195.615 43.545 195.805 ;
        RECT 45.215 195.595 45.385 195.785 ;
        RECT 48.895 195.615 49.065 195.805 ;
        RECT 51.650 195.645 51.770 195.755 ;
        RECT 52.115 195.595 52.285 195.785 ;
        RECT 52.575 195.595 52.745 195.805 ;
        RECT 54.410 195.645 54.530 195.755 ;
        RECT 58.095 195.615 58.265 195.805 ;
        RECT 60.850 195.645 60.970 195.755 ;
        RECT 61.775 195.595 61.945 195.785 ;
        RECT 62.235 195.595 62.405 195.785 ;
        RECT 64.535 195.615 64.705 195.805 ;
        RECT 65.005 195.650 65.165 195.760 ;
        RECT 65.455 195.595 65.625 195.785 ;
        RECT 66.830 195.615 67.000 195.805 ;
        RECT 67.295 195.615 67.465 195.805 ;
        RECT 70.515 195.615 70.685 195.805 ;
        RECT 78.340 195.785 78.505 195.805 ;
        RECT 72.820 195.595 72.990 195.785 ;
        RECT 78.335 195.615 78.505 195.785 ;
        RECT 79.715 195.595 79.885 195.785 ;
        RECT 80.170 195.645 80.290 195.755 ;
        RECT 80.635 195.615 80.805 195.805 ;
        RECT 81.550 195.595 81.720 195.785 ;
        RECT 82.015 195.595 82.185 195.785 ;
        RECT 85.690 195.645 85.810 195.755 ;
        RECT 86.155 195.615 86.325 195.805 ;
        RECT 88.910 195.645 89.030 195.755 ;
        RECT 89.375 195.595 89.545 195.785 ;
        RECT 89.845 195.640 90.005 195.750 ;
        RECT 90.290 195.615 90.460 195.805 ;
        RECT 90.765 195.650 90.925 195.760 ;
        RECT 98.115 195.595 98.285 195.785 ;
        RECT 98.575 195.595 98.745 195.805 ;
        RECT 99.035 195.615 99.205 195.805 ;
        RECT 101.340 195.615 101.510 195.805 ;
        RECT 103.175 195.755 103.345 195.785 ;
        RECT 102.265 195.640 102.425 195.750 ;
        RECT 103.170 195.645 103.345 195.755 ;
        RECT 103.175 195.595 103.345 195.645 ;
        RECT 104.095 195.615 104.265 195.805 ;
        RECT 107.785 195.650 107.945 195.760 ;
        RECT 110.530 195.645 110.650 195.755 ;
        RECT 114.400 195.595 114.570 195.785 ;
        RECT 115.135 195.595 115.305 195.785 ;
        RECT 115.595 195.615 115.765 195.805 ;
        RECT 116.975 195.595 117.145 195.785 ;
        RECT 122.495 195.595 122.665 195.785 ;
        RECT 122.955 195.615 123.125 195.805 ;
        RECT 123.415 195.615 123.585 195.805 ;
        RECT 128.015 195.595 128.185 195.785 ;
        RECT 128.930 195.645 129.050 195.755 ;
        RECT 129.855 195.615 130.025 195.805 ;
        RECT 133.535 195.595 133.705 195.785 ;
        RECT 135.375 195.615 135.545 195.805 ;
        RECT 137.210 195.645 137.330 195.755 ;
        RECT 138.595 195.595 138.765 195.805 ;
        RECT 13.335 194.785 14.705 195.595 ;
        RECT 14.715 194.785 20.225 195.595 ;
        RECT 20.235 194.785 25.745 195.595 ;
        RECT 25.755 194.785 31.265 195.595 ;
        RECT 32.195 194.915 35.865 195.595 ;
        RECT 34.935 194.685 35.865 194.915 ;
        RECT 35.875 194.785 38.625 195.595 ;
        RECT 39.105 194.725 39.535 195.510 ;
        RECT 39.555 194.785 45.065 195.595 ;
        RECT 45.075 194.785 50.585 195.595 ;
        RECT 50.595 194.915 52.425 195.595 ;
        RECT 52.435 194.785 54.265 195.595 ;
        RECT 54.775 194.915 62.085 195.595 ;
        RECT 54.775 194.685 56.125 194.915 ;
        RECT 57.660 194.695 58.570 194.915 ;
        RECT 62.095 194.685 64.815 195.595 ;
        RECT 64.865 194.725 65.295 195.510 ;
        RECT 65.315 194.915 72.625 195.595 ;
        RECT 68.830 194.695 69.740 194.915 ;
        RECT 71.275 194.685 72.625 194.915 ;
        RECT 72.675 194.915 76.260 195.595 ;
        RECT 76.450 194.915 79.915 195.595 ;
        RECT 72.675 194.685 73.595 194.915 ;
        RECT 76.450 194.685 77.370 194.915 ;
        RECT 80.515 194.685 81.865 195.595 ;
        RECT 81.875 194.785 85.545 195.595 ;
        RECT 86.110 194.915 89.575 195.595 ;
        RECT 86.110 194.685 87.030 194.915 ;
        RECT 90.625 194.725 91.055 195.510 ;
        RECT 91.115 194.915 98.425 195.595 ;
        RECT 98.545 194.915 102.010 195.595 ;
        RECT 103.035 194.915 110.345 195.595 ;
        RECT 111.085 194.915 114.985 195.595 ;
        RECT 91.115 194.685 92.465 194.915 ;
        RECT 94.000 194.695 94.910 194.915 ;
        RECT 101.090 194.685 102.010 194.915 ;
        RECT 106.550 194.695 107.460 194.915 ;
        RECT 108.995 194.685 110.345 194.915 ;
        RECT 114.055 194.685 114.985 194.915 ;
        RECT 114.995 194.785 116.365 195.595 ;
        RECT 116.385 194.725 116.815 195.510 ;
        RECT 116.835 194.785 122.345 195.595 ;
        RECT 122.355 194.785 127.865 195.595 ;
        RECT 127.875 194.785 133.385 195.595 ;
        RECT 133.395 194.785 137.065 195.595 ;
        RECT 137.535 194.785 138.905 195.595 ;
      LAYER nwell ;
        RECT 13.140 191.565 139.100 194.395 ;
      LAYER pwell ;
        RECT 13.335 190.365 14.705 191.175 ;
        RECT 14.715 190.365 18.385 191.175 ;
        RECT 22.370 191.045 23.280 191.265 ;
        RECT 24.815 191.045 26.165 191.275 ;
        RECT 18.855 190.365 26.165 191.045 ;
        RECT 26.225 190.450 26.655 191.235 ;
        RECT 26.675 190.365 28.505 191.175 ;
        RECT 31.715 191.045 32.645 191.275 ;
        RECT 36.170 191.045 37.080 191.265 ;
        RECT 38.615 191.045 39.965 191.275 ;
        RECT 28.975 190.365 32.645 191.045 ;
        RECT 32.655 190.365 39.965 191.045 ;
        RECT 40.015 190.365 43.685 191.175 ;
        RECT 47.210 191.045 48.120 191.265 ;
        RECT 49.655 191.045 51.005 191.275 ;
        RECT 43.695 190.365 51.005 191.045 ;
        RECT 51.985 190.450 52.415 191.235 ;
        RECT 55.950 191.045 56.860 191.265 ;
        RECT 58.395 191.045 59.745 191.275 ;
        RECT 52.435 190.365 59.745 191.045 ;
        RECT 60.255 191.045 61.175 191.275 ;
        RECT 60.255 190.365 63.840 191.045 ;
        RECT 63.955 190.365 65.305 191.275 ;
        RECT 67.970 191.045 68.890 191.275 ;
        RECT 65.425 190.365 68.890 191.045 ;
        RECT 69.005 190.365 72.665 191.275 ;
        RECT 72.675 190.365 74.045 191.175 ;
        RECT 75.390 191.075 76.345 191.275 ;
        RECT 74.065 190.395 76.345 191.075 ;
        RECT 13.475 190.155 13.645 190.365 ;
        RECT 14.855 190.155 15.025 190.365 ;
        RECT 18.530 190.205 18.650 190.315 ;
        RECT 18.995 190.175 19.165 190.365 ;
        RECT 23.595 190.155 23.765 190.345 ;
        RECT 26.815 190.155 26.985 190.365 ;
        RECT 27.275 190.155 27.445 190.345 ;
        RECT 28.655 190.315 28.825 190.345 ;
        RECT 28.650 190.205 28.825 190.315 ;
        RECT 28.655 190.155 28.825 190.205 ;
        RECT 29.115 190.175 29.285 190.365 ;
        RECT 30.955 190.155 31.125 190.345 ;
        RECT 32.795 190.175 32.965 190.365 ;
        RECT 38.325 190.200 38.485 190.310 ;
        RECT 39.695 190.155 39.865 190.345 ;
        RECT 40.155 190.175 40.325 190.365 ;
        RECT 43.835 190.175 44.005 190.365 ;
        RECT 46.135 190.155 46.305 190.345 ;
        RECT 46.595 190.155 46.765 190.345 ;
        RECT 51.205 190.210 51.365 190.320 ;
        RECT 51.655 190.155 51.825 190.345 ;
        RECT 52.115 190.155 52.285 190.345 ;
        RECT 52.575 190.175 52.745 190.365 ;
        RECT 57.635 190.155 57.805 190.345 ;
        RECT 59.930 190.205 60.050 190.315 ;
        RECT 60.400 190.175 60.570 190.365 ;
        RECT 63.150 190.205 63.270 190.315 ;
        RECT 64.070 190.175 64.240 190.365 ;
        RECT 64.535 190.155 64.705 190.345 ;
        RECT 65.455 190.175 65.625 190.365 ;
        RECT 13.335 189.345 14.705 190.155 ;
        RECT 14.715 189.345 20.225 190.155 ;
        RECT 20.235 189.475 23.905 190.155 ;
        RECT 20.235 189.245 21.165 189.475 ;
        RECT 23.915 189.245 27.085 190.155 ;
        RECT 27.135 189.345 28.505 190.155 ;
        RECT 28.515 189.475 30.805 190.155 ;
        RECT 30.815 189.475 38.125 190.155 ;
        RECT 29.885 189.245 30.805 189.475 ;
        RECT 34.330 189.255 35.240 189.475 ;
        RECT 36.775 189.245 38.125 189.475 ;
        RECT 39.105 189.285 39.535 190.070 ;
        RECT 39.595 189.245 42.765 190.155 ;
        RECT 42.775 189.475 46.445 190.155 ;
        RECT 42.775 189.245 43.705 189.475 ;
        RECT 46.455 189.345 50.125 190.155 ;
        RECT 50.135 189.245 51.950 190.155 ;
        RECT 51.975 189.345 57.485 190.155 ;
        RECT 57.495 189.345 63.005 190.155 ;
        RECT 63.485 189.245 64.835 190.155 ;
        RECT 65.315 190.125 66.270 190.155 ;
        RECT 67.300 190.125 67.470 190.345 ;
        RECT 67.755 190.175 67.925 190.345 ;
        RECT 69.130 190.175 69.300 190.365 ;
        RECT 67.760 190.155 67.925 190.175 ;
        RECT 70.055 190.155 70.225 190.345 ;
        RECT 72.815 190.175 72.985 190.365 ;
        RECT 74.190 190.175 74.360 190.395 ;
        RECT 75.390 190.365 76.345 190.395 ;
        RECT 76.355 190.365 77.705 191.275 ;
        RECT 77.745 190.450 78.175 191.235 ;
        RECT 79.155 191.045 80.505 191.275 ;
        RECT 82.040 191.045 82.950 191.265 ;
        RECT 89.130 191.045 90.050 191.275 ;
        RECT 93.670 191.045 94.580 191.265 ;
        RECT 96.115 191.045 97.465 191.275 ;
        RECT 79.155 190.365 86.465 191.045 ;
        RECT 86.585 190.365 90.050 191.045 ;
        RECT 90.155 190.365 97.465 191.045 ;
        RECT 97.610 191.045 98.530 191.275 ;
        RECT 102.530 191.075 103.485 191.275 ;
        RECT 97.610 190.365 101.075 191.045 ;
        RECT 101.205 190.395 103.485 191.075 ;
        RECT 103.505 190.450 103.935 191.235 ;
        RECT 75.575 190.155 75.745 190.345 ;
        RECT 77.420 190.175 77.590 190.365 ;
        RECT 78.345 190.210 78.505 190.320 ;
        RECT 82.935 190.155 83.105 190.345 ;
        RECT 86.155 190.175 86.325 190.365 ;
        RECT 86.615 190.345 86.785 190.365 ;
        RECT 86.615 190.175 86.790 190.345 ;
        RECT 90.295 190.315 90.465 190.365 ;
        RECT 90.290 190.205 90.465 190.315 ;
        RECT 91.210 190.205 91.330 190.315 ;
        RECT 90.295 190.175 90.465 190.205 ;
        RECT 86.620 190.155 86.790 190.175 ;
        RECT 91.675 190.155 91.845 190.345 ;
        RECT 64.865 189.285 65.295 190.070 ;
        RECT 65.315 189.445 67.595 190.125 ;
        RECT 67.760 189.475 69.595 190.155 ;
        RECT 65.315 189.245 66.270 189.445 ;
        RECT 68.665 189.245 69.595 189.475 ;
        RECT 69.915 189.345 75.425 190.155 ;
        RECT 75.435 189.475 82.745 190.155 ;
        RECT 78.950 189.255 79.860 189.475 ;
        RECT 81.395 189.245 82.745 189.475 ;
        RECT 82.795 189.345 86.465 190.155 ;
        RECT 86.475 189.245 89.950 190.155 ;
        RECT 90.625 189.285 91.055 190.070 ;
        RECT 91.535 189.475 95.205 190.155 ;
        RECT 95.360 190.125 95.530 190.345 ;
        RECT 100.875 190.175 101.045 190.365 ;
        RECT 101.330 190.345 101.500 190.395 ;
        RECT 102.530 190.365 103.485 190.395 ;
        RECT 103.955 190.365 107.165 191.275 ;
        RECT 107.175 190.365 109.365 191.275 ;
        RECT 109.935 190.365 113.605 191.275 ;
        RECT 113.925 191.045 114.855 191.275 ;
        RECT 113.925 190.365 115.760 191.045 ;
        RECT 115.915 190.365 117.265 191.275 ;
        RECT 117.295 190.365 118.645 191.275 ;
        RECT 118.675 190.365 124.185 191.175 ;
        RECT 124.195 190.365 127.865 191.175 ;
        RECT 127.875 190.365 129.245 191.175 ;
        RECT 129.265 190.450 129.695 191.235 ;
        RECT 129.715 190.365 133.385 191.175 ;
        RECT 133.855 190.365 135.225 191.145 ;
        RECT 136.155 190.365 137.525 191.145 ;
        RECT 137.535 190.365 138.905 191.175 ;
        RECT 101.330 190.175 101.505 190.345 ;
        RECT 101.335 190.155 101.505 190.175 ;
        RECT 101.795 190.155 101.965 190.345 ;
        RECT 104.085 190.175 104.255 190.365 ;
        RECT 104.560 190.155 104.730 190.345 ;
        RECT 107.320 190.175 107.490 190.365 ;
        RECT 108.695 190.155 108.865 190.345 ;
        RECT 109.165 190.200 109.325 190.310 ;
        RECT 109.610 190.205 109.730 190.315 ;
        RECT 110.075 190.155 110.245 190.345 ;
        RECT 97.490 190.125 98.425 190.155 ;
        RECT 95.360 189.925 98.425 190.125 ;
        RECT 94.275 189.245 95.205 189.475 ;
        RECT 95.215 189.445 98.425 189.925 ;
        RECT 95.215 189.245 96.145 189.445 ;
        RECT 97.475 189.245 98.425 189.445 ;
        RECT 98.435 189.245 101.645 190.155 ;
        RECT 101.655 189.245 104.405 190.155 ;
        RECT 104.415 189.245 106.605 190.155 ;
        RECT 106.715 189.475 109.005 190.155 ;
        RECT 109.935 189.475 112.225 190.155 ;
        RECT 112.380 190.125 112.550 190.345 ;
        RECT 113.290 190.175 113.460 190.365 ;
        RECT 115.595 190.345 115.760 190.365 ;
        RECT 115.595 190.175 115.765 190.345 ;
        RECT 116.060 190.175 116.230 190.365 ;
        RECT 116.975 190.155 117.145 190.345 ;
        RECT 118.360 190.175 118.530 190.365 ;
        RECT 118.815 190.175 118.985 190.365 ;
        RECT 122.495 190.155 122.665 190.345 ;
        RECT 124.335 190.315 124.505 190.365 ;
        RECT 124.330 190.205 124.505 190.315 ;
        RECT 124.335 190.175 124.505 190.205 ;
        RECT 124.795 190.155 124.965 190.345 ;
        RECT 128.015 190.175 128.185 190.365 ;
        RECT 129.855 190.175 130.025 190.365 ;
        RECT 133.530 190.205 133.650 190.315 ;
        RECT 133.995 190.175 134.165 190.365 ;
        RECT 135.375 190.155 135.545 190.345 ;
        RECT 135.835 190.155 136.005 190.345 ;
        RECT 137.205 190.175 137.375 190.365 ;
        RECT 138.595 190.155 138.765 190.365 ;
        RECT 114.510 190.125 115.445 190.155 ;
        RECT 112.380 189.925 115.445 190.125 ;
        RECT 106.715 189.245 107.635 189.475 ;
        RECT 111.305 189.245 112.225 189.475 ;
        RECT 112.235 189.445 115.445 189.925 ;
        RECT 112.235 189.245 113.165 189.445 ;
        RECT 114.495 189.245 115.445 189.445 ;
        RECT 116.385 189.285 116.815 190.070 ;
        RECT 116.835 189.345 122.345 190.155 ;
        RECT 122.355 189.345 124.185 190.155 ;
        RECT 124.655 189.475 131.965 190.155 ;
        RECT 128.170 189.255 129.080 189.475 ;
        RECT 130.615 189.245 131.965 189.475 ;
        RECT 132.110 189.475 135.575 190.155 ;
        RECT 135.695 189.475 137.525 190.155 ;
        RECT 132.110 189.245 133.030 189.475 ;
        RECT 136.180 189.245 137.525 189.475 ;
        RECT 137.535 189.345 138.905 190.155 ;
      LAYER nwell ;
        RECT 13.140 186.125 139.100 188.955 ;
      LAYER pwell ;
        RECT 13.335 184.925 14.705 185.735 ;
        RECT 14.715 184.925 18.385 185.735 ;
        RECT 18.395 185.605 19.325 185.835 ;
        RECT 18.395 184.925 22.065 185.605 ;
        RECT 22.075 184.925 25.745 185.735 ;
        RECT 26.225 185.010 26.655 185.795 ;
        RECT 26.675 184.925 30.345 185.735 ;
        RECT 30.835 184.925 32.185 185.835 ;
        RECT 32.210 184.925 34.025 185.835 ;
        RECT 36.110 185.605 37.245 185.835 ;
        RECT 34.035 184.925 37.245 185.605 ;
        RECT 37.275 184.925 38.625 185.835 ;
        RECT 38.635 184.925 39.985 185.835 ;
        RECT 40.015 184.925 45.525 185.735 ;
        RECT 48.275 185.605 49.205 185.835 ;
        RECT 45.535 184.925 49.205 185.605 ;
        RECT 49.215 184.925 50.565 185.835 ;
        RECT 50.595 184.925 51.965 185.735 ;
        RECT 51.985 185.010 52.415 185.795 ;
        RECT 52.435 184.925 57.945 185.735 ;
        RECT 58.875 184.925 61.795 185.835 ;
        RECT 62.190 185.605 63.110 185.835 ;
        RECT 65.870 185.605 66.790 185.835 ;
        RECT 62.190 184.925 65.655 185.605 ;
        RECT 65.870 184.925 69.335 185.605 ;
        RECT 69.475 184.925 70.825 185.835 ;
        RECT 70.835 184.925 72.185 185.835 ;
        RECT 72.215 184.925 77.725 185.735 ;
        RECT 77.745 185.010 78.175 185.795 ;
        RECT 80.850 185.605 81.770 185.835 ;
        RECT 78.305 184.925 81.770 185.605 ;
        RECT 81.875 184.925 87.385 185.735 ;
        RECT 87.855 184.925 89.205 185.835 ;
        RECT 89.255 184.925 90.605 185.835 ;
        RECT 90.615 184.925 92.445 185.735 ;
        RECT 94.275 185.605 95.205 185.835 ;
        RECT 92.455 184.925 95.205 185.605 ;
        RECT 95.225 184.925 96.575 185.835 ;
        RECT 97.065 184.925 98.415 185.835 ;
        RECT 98.435 184.925 99.805 185.735 ;
        RECT 100.270 185.155 102.105 185.835 ;
        RECT 100.270 184.925 101.960 185.155 ;
        RECT 102.115 184.925 103.485 185.735 ;
        RECT 103.505 185.010 103.935 185.795 ;
        RECT 103.955 184.925 106.705 185.735 ;
        RECT 107.175 185.605 108.095 185.835 ;
        RECT 111.295 185.605 112.225 185.835 ;
        RECT 107.175 184.925 109.465 185.605 ;
        RECT 109.475 184.925 112.225 185.605 ;
        RECT 112.235 185.605 113.165 185.835 ;
        RECT 116.330 185.635 117.285 185.835 ;
        RECT 112.235 184.925 114.985 185.605 ;
        RECT 115.005 184.955 117.285 185.635 ;
        RECT 13.475 184.715 13.645 184.925 ;
        RECT 14.855 184.715 15.025 184.925 ;
        RECT 16.235 184.715 16.405 184.905 ;
        RECT 18.075 184.715 18.245 184.905 ;
        RECT 21.755 184.735 21.925 184.925 ;
        RECT 22.215 184.735 22.385 184.925 ;
        RECT 25.440 184.715 25.610 184.905 ;
        RECT 25.890 184.765 26.010 184.875 ;
        RECT 26.815 184.715 26.985 184.925 ;
        RECT 30.490 184.765 30.610 184.875 ;
        RECT 31.870 184.735 32.040 184.925 ;
        RECT 32.335 184.715 32.505 184.925 ;
        RECT 34.175 184.735 34.345 184.925 ;
        RECT 37.855 184.715 38.025 184.905 ;
        RECT 38.310 184.735 38.480 184.925 ;
        RECT 38.780 184.735 38.950 184.925 ;
        RECT 39.695 184.715 39.865 184.905 ;
        RECT 40.155 184.735 40.325 184.925 ;
        RECT 41.530 184.765 41.650 184.875 ;
        RECT 43.375 184.715 43.545 184.905 ;
        RECT 43.835 184.715 44.005 184.905 ;
        RECT 45.675 184.735 45.845 184.925 ;
        RECT 46.135 184.715 46.305 184.905 ;
        RECT 49.360 184.735 49.530 184.925 ;
        RECT 50.735 184.735 50.905 184.925 ;
        RECT 52.575 184.735 52.745 184.925 ;
        RECT 53.495 184.715 53.665 184.905 ;
        RECT 57.170 184.765 57.290 184.875 ;
        RECT 57.635 184.715 57.805 184.905 ;
        RECT 58.105 184.770 58.265 184.880 ;
        RECT 59.020 184.735 59.190 184.925 ;
        RECT 65.455 184.715 65.625 184.925 ;
        RECT 68.215 184.715 68.385 184.905 ;
        RECT 69.135 184.735 69.305 184.925 ;
        RECT 69.590 184.735 69.760 184.925 ;
        RECT 71.900 184.735 72.070 184.925 ;
        RECT 72.355 184.735 72.525 184.925 ;
        RECT 78.335 184.735 78.505 184.925 ;
        RECT 82.015 184.735 82.185 184.925 ;
        RECT 82.475 184.715 82.645 184.905 ;
        RECT 86.155 184.715 86.325 184.905 ;
        RECT 86.615 184.715 86.785 184.905 ;
        RECT 87.530 184.765 87.650 184.875 ;
        RECT 88.920 184.735 89.090 184.925 ;
        RECT 90.290 184.735 90.460 184.925 ;
        RECT 90.755 184.735 90.925 184.925 ;
        RECT 91.215 184.715 91.385 184.905 ;
        RECT 92.595 184.735 92.765 184.925 ;
        RECT 96.275 184.735 96.445 184.925 ;
        RECT 96.735 184.875 96.905 184.905 ;
        RECT 96.730 184.765 96.905 184.875 ;
        RECT 96.735 184.715 96.905 184.765 ;
        RECT 97.195 184.735 97.365 184.925 ;
        RECT 98.575 184.735 98.745 184.925 ;
        RECT 101.790 184.735 101.960 184.925 ;
        RECT 102.255 184.715 102.425 184.925 ;
        RECT 104.095 184.735 104.265 184.925 ;
        RECT 105.930 184.765 106.050 184.875 ;
        RECT 106.850 184.765 106.970 184.875 ;
        RECT 109.155 184.715 109.325 184.925 ;
        RECT 109.615 184.905 109.785 184.925 ;
        RECT 109.615 184.735 109.790 184.905 ;
        RECT 109.620 184.715 109.790 184.735 ;
        RECT 111.920 184.715 112.090 184.905 ;
        RECT 114.675 184.735 114.845 184.925 ;
        RECT 115.130 184.735 115.300 184.955 ;
        RECT 116.330 184.925 117.285 184.955 ;
        RECT 117.295 184.925 119.125 185.835 ;
        RECT 119.620 185.605 120.965 185.835 ;
        RECT 119.135 184.925 120.965 185.605 ;
        RECT 120.975 184.925 126.485 185.735 ;
        RECT 126.495 184.925 129.245 185.735 ;
        RECT 129.265 185.010 129.695 185.795 ;
        RECT 129.715 185.605 130.645 185.835 ;
        RECT 134.340 185.605 135.685 185.835 ;
        RECT 136.180 185.605 137.525 185.835 ;
        RECT 129.715 184.925 133.615 185.605 ;
        RECT 133.855 184.925 135.685 185.605 ;
        RECT 135.695 184.925 137.525 185.605 ;
        RECT 137.535 184.925 138.905 185.735 ;
        RECT 115.590 184.715 115.760 184.905 ;
        RECT 116.050 184.765 116.170 184.875 ;
        RECT 117.440 184.735 117.610 184.925 ;
        RECT 119.275 184.735 119.445 184.925 ;
        RECT 120.190 184.715 120.360 184.905 ;
        RECT 120.660 184.715 120.830 184.905 ;
        RECT 121.115 184.735 121.285 184.925 ;
        RECT 122.955 184.715 123.125 184.905 ;
        RECT 124.790 184.765 124.910 184.875 ;
        RECT 125.255 184.715 125.425 184.905 ;
        RECT 126.635 184.715 126.805 184.925 ;
        RECT 130.130 184.735 130.300 184.925 ;
        RECT 133.995 184.735 134.165 184.925 ;
        RECT 135.835 184.735 136.005 184.925 ;
        RECT 137.215 184.715 137.385 184.905 ;
        RECT 138.595 184.715 138.765 184.925 ;
        RECT 13.335 183.905 14.705 184.715 ;
        RECT 14.715 183.935 16.085 184.715 ;
        RECT 16.095 183.905 17.925 184.715 ;
        RECT 17.935 184.035 25.245 184.715 ;
        RECT 21.450 183.815 22.360 184.035 ;
        RECT 23.895 183.805 25.245 184.035 ;
        RECT 25.295 183.805 26.645 184.715 ;
        RECT 26.675 183.905 32.185 184.715 ;
        RECT 32.195 183.905 37.705 184.715 ;
        RECT 37.715 183.905 39.085 184.715 ;
        RECT 39.105 183.845 39.535 184.630 ;
        RECT 39.555 183.905 41.385 184.715 ;
        RECT 41.855 183.805 43.670 184.715 ;
        RECT 43.695 184.035 45.985 184.715 ;
        RECT 45.995 184.035 53.305 184.715 ;
        RECT 45.065 183.805 45.985 184.035 ;
        RECT 49.510 183.815 50.420 184.035 ;
        RECT 51.955 183.805 53.305 184.035 ;
        RECT 53.355 183.905 57.025 184.715 ;
        RECT 57.495 184.035 64.805 184.715 ;
        RECT 61.010 183.815 61.920 184.035 ;
        RECT 63.455 183.805 64.805 184.035 ;
        RECT 64.865 183.845 65.295 184.630 ;
        RECT 65.325 183.805 68.055 184.715 ;
        RECT 68.075 184.035 75.385 184.715 ;
        RECT 71.590 183.815 72.500 184.035 ;
        RECT 74.035 183.805 75.385 184.035 ;
        RECT 75.475 184.035 82.785 184.715 ;
        RECT 82.890 184.035 86.355 184.715 ;
        RECT 75.475 183.805 76.825 184.035 ;
        RECT 78.360 183.815 79.270 184.035 ;
        RECT 82.890 183.805 83.810 184.035 ;
        RECT 86.475 183.905 90.145 184.715 ;
        RECT 90.625 183.845 91.055 184.630 ;
        RECT 91.075 183.905 96.585 184.715 ;
        RECT 96.595 183.905 102.105 184.715 ;
        RECT 102.115 183.905 105.785 184.715 ;
        RECT 106.385 183.805 109.385 184.715 ;
        RECT 109.475 184.035 111.750 184.715 ;
        RECT 110.380 183.805 111.750 184.035 ;
        RECT 111.775 183.805 113.605 184.715 ;
        RECT 113.630 184.035 115.905 184.715 ;
        RECT 113.630 183.805 115.000 184.035 ;
        RECT 116.385 183.845 116.815 184.630 ;
        RECT 117.030 183.805 120.505 184.715 ;
        RECT 120.515 183.805 122.725 184.715 ;
        RECT 122.815 183.905 124.645 184.715 ;
        RECT 125.115 183.935 126.485 184.715 ;
        RECT 126.495 184.035 133.805 184.715 ;
        RECT 130.010 183.815 130.920 184.035 ;
        RECT 132.455 183.805 133.805 184.035 ;
        RECT 133.950 184.035 137.415 184.715 ;
        RECT 133.950 183.805 134.870 184.035 ;
        RECT 137.535 183.905 138.905 184.715 ;
      LAYER nwell ;
        RECT 13.140 180.685 139.100 183.515 ;
      LAYER pwell ;
        RECT 13.335 179.485 14.705 180.295 ;
        RECT 14.715 179.485 16.545 180.295 ;
        RECT 20.530 180.165 21.440 180.385 ;
        RECT 22.975 180.165 24.325 180.395 ;
        RECT 17.015 179.485 24.325 180.165 ;
        RECT 24.375 179.485 25.725 180.395 ;
        RECT 26.225 179.570 26.655 180.355 ;
        RECT 26.675 179.485 28.505 180.295 ;
        RECT 29.460 180.165 30.805 180.395 ;
        RECT 28.975 179.485 30.805 180.165 ;
        RECT 31.270 179.715 33.105 180.395 ;
        RECT 31.270 179.485 32.960 179.715 ;
        RECT 33.115 179.485 35.865 180.395 ;
        RECT 35.875 179.485 39.085 180.395 ;
        RECT 42.055 180.305 43.005 180.395 ;
        RECT 39.105 179.485 41.845 180.165 ;
        RECT 42.055 179.485 43.985 180.305 ;
        RECT 44.655 180.165 46.005 180.395 ;
        RECT 47.540 180.165 48.450 180.385 ;
        RECT 44.655 179.485 51.965 180.165 ;
        RECT 51.985 179.570 52.415 180.355 ;
        RECT 52.435 180.165 53.570 180.395 ;
        RECT 52.435 179.485 55.645 180.165 ;
        RECT 55.655 179.485 57.025 180.295 ;
        RECT 60.550 180.165 61.460 180.385 ;
        RECT 62.995 180.165 64.345 180.395 ;
        RECT 57.035 179.485 64.345 180.165 ;
        RECT 64.415 179.485 65.765 180.395 ;
        RECT 65.775 179.485 67.145 180.295 ;
        RECT 67.250 180.165 68.170 180.395 ;
        RECT 67.250 179.485 70.715 180.165 ;
        RECT 71.005 179.485 74.505 180.395 ;
        RECT 74.515 180.195 75.460 180.395 ;
        RECT 76.795 180.195 77.725 180.395 ;
        RECT 74.515 179.715 77.725 180.195 ;
        RECT 74.515 179.515 77.585 179.715 ;
        RECT 77.745 179.570 78.175 180.355 ;
        RECT 81.855 180.165 82.785 180.395 ;
        RECT 74.515 179.485 75.460 179.515 ;
        RECT 13.475 179.275 13.645 179.485 ;
        RECT 14.855 179.275 15.025 179.485 ;
        RECT 16.690 179.325 16.810 179.435 ;
        RECT 17.155 179.295 17.325 179.485 ;
        RECT 17.610 179.275 17.780 179.465 ;
        RECT 21.295 179.275 21.465 179.465 ;
        RECT 23.595 179.275 23.765 179.465 ;
        RECT 24.055 179.275 24.225 179.465 ;
        RECT 24.520 179.295 24.690 179.485 ;
        RECT 25.890 179.325 26.010 179.435 ;
        RECT 26.815 179.295 26.985 179.485 ;
        RECT 27.275 179.275 27.445 179.465 ;
        RECT 28.650 179.325 28.770 179.435 ;
        RECT 29.115 179.295 29.285 179.485 ;
        RECT 32.790 179.295 32.960 179.485 ;
        RECT 33.250 179.275 33.420 179.465 ;
        RECT 33.710 179.325 33.830 179.435 ;
        RECT 35.555 179.295 35.725 179.485 ;
        RECT 36.015 179.295 36.185 179.485 ;
        RECT 38.775 179.275 38.945 179.465 ;
        RECT 39.700 179.275 39.870 179.465 ;
        RECT 41.535 179.295 41.705 179.485 ;
        RECT 43.835 179.465 43.985 179.485 ;
        RECT 43.835 179.295 44.005 179.465 ;
        RECT 44.290 179.325 44.410 179.435 ;
        RECT 51.655 179.295 51.825 179.485 ;
        RECT 55.335 179.275 55.505 179.485 ;
        RECT 55.795 179.465 55.965 179.485 ;
        RECT 55.795 179.295 55.970 179.465 ;
        RECT 55.800 179.275 55.970 179.295 ;
        RECT 57.175 179.275 57.345 179.485 ;
        RECT 62.695 179.275 62.865 179.465 ;
        RECT 64.530 179.295 64.700 179.485 ;
        RECT 65.915 179.295 66.085 179.485 ;
        RECT 70.515 179.295 70.685 179.485 ;
        RECT 71.005 179.465 71.140 179.485 ;
        RECT 70.970 179.295 71.140 179.465 ;
        RECT 72.355 179.275 72.525 179.465 ;
        RECT 72.815 179.275 72.985 179.465 ;
        RECT 77.415 179.295 77.585 179.515 ;
        RECT 78.885 179.485 82.785 180.165 ;
        RECT 82.795 179.485 84.145 180.395 ;
        RECT 84.175 179.485 89.685 180.295 ;
        RECT 89.695 179.485 91.065 180.295 ;
        RECT 91.075 180.165 92.005 180.395 ;
        RECT 95.310 180.165 96.230 180.395 ;
        RECT 101.550 180.165 102.470 180.395 ;
        RECT 91.075 179.485 94.975 180.165 ;
        RECT 95.310 179.485 98.775 180.165 ;
        RECT 99.005 179.485 102.470 180.165 ;
        RECT 103.505 179.570 103.935 180.355 ;
        RECT 104.035 179.485 106.245 180.395 ;
        RECT 106.255 179.485 107.605 180.395 ;
        RECT 107.635 179.485 108.985 180.395 ;
        RECT 110.810 180.195 111.765 180.395 ;
        RECT 109.485 179.515 111.765 180.195 ;
        RECT 78.330 179.325 78.450 179.435 ;
        RECT 79.715 179.295 79.885 179.465 ;
        RECT 77.415 179.275 77.580 179.295 ;
        RECT 79.715 179.275 79.865 179.295 ;
        RECT 80.175 179.275 80.345 179.465 ;
        RECT 82.200 179.295 82.370 179.485 ;
        RECT 82.940 179.295 83.110 179.485 ;
        RECT 84.130 179.275 84.300 179.465 ;
        RECT 84.315 179.295 84.485 179.485 ;
        RECT 87.995 179.275 88.165 179.465 ;
        RECT 89.835 179.295 90.005 179.485 ;
        RECT 91.490 179.295 91.660 179.485 ;
        RECT 98.115 179.275 98.285 179.465 ;
        RECT 98.575 179.295 98.745 179.485 ;
        RECT 99.035 179.295 99.205 179.485 ;
        RECT 101.335 179.275 101.505 179.465 ;
        RECT 101.785 179.275 101.955 179.465 ;
        RECT 102.725 179.330 102.885 179.440 ;
        RECT 105.015 179.275 105.185 179.465 ;
        RECT 105.930 179.295 106.100 179.485 ;
        RECT 106.400 179.295 106.570 179.485 ;
        RECT 108.700 179.295 108.870 179.485 ;
        RECT 109.610 179.465 109.780 179.515 ;
        RECT 110.810 179.485 111.765 179.515 ;
        RECT 111.925 179.485 115.580 180.395 ;
        RECT 117.250 180.195 118.205 180.395 ;
        RECT 115.925 179.515 118.205 180.195 ;
        RECT 119.265 180.165 120.195 180.395 ;
        RECT 111.925 179.465 112.085 179.485 ;
        RECT 109.150 179.325 109.270 179.435 ;
        RECT 109.610 179.295 109.785 179.465 ;
        RECT 111.915 179.295 112.085 179.465 ;
        RECT 109.615 179.275 109.785 179.295 ;
        RECT 112.835 179.275 113.005 179.465 ;
        RECT 115.605 179.320 115.765 179.430 ;
        RECT 116.050 179.295 116.220 179.515 ;
        RECT 117.250 179.485 118.205 179.515 ;
        RECT 118.360 179.485 120.195 180.165 ;
        RECT 120.515 179.485 121.885 180.295 ;
        RECT 121.895 179.485 125.105 180.395 ;
        RECT 128.315 180.165 129.245 180.395 ;
        RECT 125.345 179.485 129.245 180.165 ;
        RECT 129.265 179.570 129.695 180.355 ;
        RECT 133.230 180.165 134.140 180.385 ;
        RECT 135.675 180.165 137.025 180.395 ;
        RECT 129.715 179.485 137.025 180.165 ;
        RECT 137.535 179.485 138.905 180.295 ;
        RECT 118.360 179.465 118.525 179.485 ;
        RECT 116.975 179.295 117.145 179.465 ;
        RECT 118.355 179.295 118.525 179.465 ;
        RECT 120.655 179.295 120.825 179.485 ;
        RECT 116.985 179.275 117.145 179.295 ;
        RECT 121.115 179.275 121.285 179.465 ;
        RECT 122.035 179.295 122.205 179.485 ;
        RECT 124.335 179.275 124.505 179.465 ;
        RECT 128.660 179.295 128.830 179.485 ;
        RECT 129.855 179.295 130.025 179.485 ;
        RECT 130.960 179.275 131.130 179.465 ;
        RECT 131.695 179.275 131.865 179.465 ;
        RECT 136.295 179.275 136.465 179.465 ;
        RECT 136.765 179.320 136.925 179.430 ;
        RECT 137.210 179.325 137.330 179.435 ;
        RECT 138.595 179.275 138.765 179.485 ;
        RECT 13.335 178.465 14.705 179.275 ;
        RECT 14.715 178.465 16.545 179.275 ;
        RECT 16.575 178.365 17.925 179.275 ;
        RECT 17.935 178.595 21.605 179.275 ;
        RECT 21.615 178.595 23.905 179.275 ;
        RECT 23.915 178.595 27.125 179.275 ;
        RECT 17.935 178.365 18.865 178.595 ;
        RECT 21.615 178.365 22.535 178.595 ;
        RECT 25.990 178.365 27.125 178.595 ;
        RECT 27.135 178.465 29.885 179.275 ;
        RECT 30.090 178.365 33.565 179.275 ;
        RECT 34.270 178.595 39.085 179.275 ;
        RECT 39.105 178.405 39.535 179.190 ;
        RECT 39.555 178.365 50.565 179.275 ;
        RECT 50.830 178.595 55.645 179.275 ;
        RECT 55.655 178.365 57.005 179.275 ;
        RECT 57.035 178.465 62.545 179.275 ;
        RECT 62.555 178.465 64.385 179.275 ;
        RECT 64.865 178.405 65.295 179.190 ;
        RECT 65.355 178.595 72.665 179.275 ;
        RECT 65.355 178.365 66.705 178.595 ;
        RECT 68.240 178.375 69.150 178.595 ;
        RECT 72.685 178.365 75.415 179.275 ;
        RECT 75.745 178.595 77.580 179.275 ;
        RECT 75.745 178.365 76.675 178.595 ;
        RECT 77.935 178.455 79.865 179.275 ;
        RECT 80.145 178.595 83.610 179.275 ;
        RECT 77.935 178.365 78.885 178.455 ;
        RECT 82.690 178.365 83.610 178.595 ;
        RECT 83.715 178.595 87.615 179.275 ;
        RECT 83.715 178.365 84.645 178.595 ;
        RECT 87.855 178.465 90.605 179.275 ;
        RECT 90.625 178.405 91.055 179.190 ;
        RECT 91.115 178.595 98.425 179.275 ;
        RECT 91.115 178.365 92.465 178.595 ;
        RECT 94.000 178.375 94.910 178.595 ;
        RECT 98.435 178.365 101.645 179.275 ;
        RECT 101.655 178.365 104.865 179.275 ;
        RECT 104.875 178.465 108.545 179.275 ;
        RECT 109.475 178.365 112.685 179.275 ;
        RECT 112.705 178.365 115.435 179.275 ;
        RECT 116.385 178.405 116.815 179.190 ;
        RECT 116.985 178.365 120.640 179.275 ;
        RECT 120.975 178.365 124.185 179.275 ;
        RECT 124.195 178.365 127.405 179.275 ;
        RECT 127.645 178.595 131.545 179.275 ;
        RECT 130.615 178.365 131.545 178.595 ;
        RECT 131.555 178.495 132.925 179.275 ;
        RECT 133.030 178.595 136.495 179.275 ;
        RECT 133.030 178.365 133.950 178.595 ;
        RECT 137.535 178.465 138.905 179.275 ;
      LAYER nwell ;
        RECT 13.140 175.245 139.100 178.075 ;
      LAYER pwell ;
        RECT 13.335 174.045 14.705 174.855 ;
        RECT 14.715 174.045 20.225 174.855 ;
        RECT 21.155 174.045 22.970 174.955 ;
        RECT 22.995 174.045 25.745 174.855 ;
        RECT 26.225 174.130 26.655 174.915 ;
        RECT 26.675 174.045 28.505 174.855 ;
        RECT 30.310 174.755 31.265 174.955 ;
        RECT 28.985 174.075 31.265 174.755 ;
        RECT 13.475 173.835 13.645 174.045 ;
        RECT 14.855 173.835 15.025 174.045 ;
        RECT 17.610 173.885 17.730 173.995 ;
        RECT 18.075 173.835 18.245 174.025 ;
        RECT 20.385 173.890 20.545 174.000 ;
        RECT 22.675 173.835 22.845 174.045 ;
        RECT 23.135 173.835 23.305 174.045 ;
        RECT 25.895 173.995 26.065 174.025 ;
        RECT 25.890 173.885 26.065 173.995 ;
        RECT 25.895 173.835 26.065 173.885 ;
        RECT 26.815 173.855 26.985 174.045 ;
        RECT 29.110 174.025 29.280 174.075 ;
        RECT 30.310 174.045 31.265 174.075 ;
        RECT 32.215 174.045 33.565 174.955 ;
        RECT 33.770 174.045 37.245 174.955 ;
        RECT 37.255 174.755 38.200 174.955 ;
        RECT 39.535 174.755 40.465 174.955 ;
        RECT 37.255 174.275 40.465 174.755 ;
        RECT 41.525 174.725 42.455 174.955 ;
        RECT 37.255 174.075 40.325 174.275 ;
        RECT 37.255 174.045 38.200 174.075 ;
        RECT 32.330 174.025 32.500 174.045 ;
        RECT 28.650 173.885 28.770 173.995 ;
        RECT 29.110 173.855 29.285 174.025 ;
        RECT 31.425 173.890 31.585 174.000 ;
        RECT 32.330 173.855 32.505 174.025 ;
        RECT 35.090 173.885 35.210 173.995 ;
        RECT 29.115 173.835 29.285 173.855 ;
        RECT 32.335 173.835 32.505 173.855 ;
        RECT 13.335 173.025 14.705 173.835 ;
        RECT 14.715 173.025 17.465 173.835 ;
        RECT 17.975 172.925 21.145 173.835 ;
        RECT 21.155 173.155 22.985 173.835 ;
        RECT 22.995 173.025 25.745 173.835 ;
        RECT 25.855 172.925 28.965 173.835 ;
        RECT 29.075 172.925 32.185 173.835 ;
        RECT 32.195 173.025 34.945 173.835 ;
        RECT 35.550 173.805 35.720 174.025 ;
        RECT 36.930 173.855 37.100 174.045 ;
        RECT 37.855 173.835 38.025 174.025 ;
        RECT 39.700 173.835 39.870 174.025 ;
        RECT 40.155 173.855 40.325 174.075 ;
        RECT 40.620 174.045 42.455 174.725 ;
        RECT 42.775 174.045 46.445 174.855 ;
        RECT 49.195 174.725 50.125 174.955 ;
        RECT 46.455 174.045 50.125 174.725 ;
        RECT 50.155 174.045 51.505 174.955 ;
        RECT 51.985 174.130 52.415 174.915 ;
        RECT 52.815 174.045 55.240 174.725 ;
        RECT 55.655 174.045 59.325 174.855 ;
        RECT 60.255 174.045 65.070 174.725 ;
        RECT 65.315 174.045 76.325 174.955 ;
        RECT 76.355 174.045 77.705 174.955 ;
        RECT 77.745 174.130 78.175 174.915 ;
        RECT 78.695 174.725 80.045 174.955 ;
        RECT 81.580 174.725 82.490 174.945 ;
        RECT 89.530 174.725 90.440 174.945 ;
        RECT 91.975 174.725 93.325 174.955 ;
        RECT 78.695 174.045 86.005 174.725 ;
        RECT 86.015 174.045 93.325 174.725 ;
        RECT 93.375 174.045 95.205 174.855 ;
        RECT 95.255 174.725 96.605 174.955 ;
        RECT 98.140 174.725 99.050 174.945 ;
        RECT 95.255 174.045 102.565 174.725 ;
        RECT 103.505 174.130 103.935 174.915 ;
        RECT 106.610 174.725 107.530 174.955 ;
        RECT 104.065 174.045 107.530 174.725 ;
        RECT 107.715 174.045 110.715 174.955 ;
        RECT 110.855 174.045 113.775 174.955 ;
        RECT 114.075 174.045 115.905 174.855 ;
        RECT 115.925 174.045 118.655 174.955 ;
        RECT 118.985 174.725 119.915 174.955 ;
        RECT 118.985 174.045 120.820 174.725 ;
        RECT 120.975 174.045 126.485 174.855 ;
        RECT 127.900 174.725 129.245 174.955 ;
        RECT 127.415 174.045 129.245 174.725 ;
        RECT 129.265 174.130 129.695 174.915 ;
        RECT 129.715 174.725 130.645 174.955 ;
        RECT 133.950 174.725 134.870 174.955 ;
        RECT 129.715 174.045 133.615 174.725 ;
        RECT 133.950 174.045 137.415 174.725 ;
        RECT 137.535 174.045 138.905 174.855 ;
        RECT 40.620 174.025 40.785 174.045 ;
        RECT 40.615 173.855 40.785 174.025 ;
        RECT 42.915 173.855 43.085 174.045 ;
        RECT 43.375 173.835 43.545 174.025 ;
        RECT 46.595 173.855 46.765 174.045 ;
        RECT 48.895 173.835 49.065 174.025 ;
        RECT 51.190 173.855 51.360 174.045 ;
        RECT 51.650 173.885 51.770 173.995 ;
        RECT 53.495 173.835 53.665 174.025 ;
        RECT 53.955 173.835 54.125 174.025 ;
        RECT 55.335 173.855 55.505 174.025 ;
        RECT 55.795 173.855 55.965 174.045 ;
        RECT 59.475 173.835 59.645 174.025 ;
        RECT 60.395 173.855 60.565 174.045 ;
        RECT 65.460 174.025 65.630 174.045 ;
        RECT 61.320 173.835 61.490 174.025 ;
        RECT 63.155 173.835 63.325 174.025 ;
        RECT 65.455 173.855 65.630 174.025 ;
        RECT 65.455 173.835 65.625 173.855 ;
        RECT 72.815 173.835 72.985 174.025 ;
        RECT 74.195 173.835 74.365 174.025 ;
        RECT 77.420 173.855 77.590 174.045 ;
        RECT 78.150 173.835 78.320 174.025 ;
        RECT 78.330 173.885 78.450 173.995 ;
        RECT 82.290 173.835 82.460 174.025 ;
        RECT 85.695 173.855 85.865 174.045 ;
        RECT 86.155 173.835 86.325 174.045 ;
        RECT 89.845 173.880 90.005 173.990 ;
        RECT 91.215 173.835 91.385 174.025 ;
        RECT 93.515 173.855 93.685 174.045 ;
        RECT 102.255 174.025 102.425 174.045 ;
        RECT 93.975 173.835 94.145 174.025 ;
        RECT 99.035 173.835 99.205 174.025 ;
        RECT 101.790 173.885 101.910 173.995 ;
        RECT 102.250 173.855 102.425 174.025 ;
        RECT 102.725 173.890 102.885 174.000 ;
        RECT 102.250 173.835 102.420 173.855 ;
        RECT 103.635 173.835 103.805 174.025 ;
        RECT 104.095 173.855 104.265 174.045 ;
        RECT 107.775 173.855 107.945 174.045 ;
        RECT 109.155 173.835 109.325 174.025 ;
        RECT 111.000 173.855 111.170 174.045 ;
        RECT 112.830 173.885 112.950 173.995 ;
        RECT 114.215 173.855 114.385 174.045 ;
        RECT 115.135 173.835 115.305 174.025 ;
        RECT 115.605 173.880 115.765 173.990 ;
        RECT 118.355 173.855 118.525 174.045 ;
        RECT 120.655 174.025 120.820 174.045 ;
        RECT 120.190 173.835 120.360 174.025 ;
        RECT 120.655 173.835 120.825 174.025 ;
        RECT 121.115 173.855 121.285 174.045 ;
        RECT 124.335 173.835 124.505 174.025 ;
        RECT 125.715 173.835 125.885 174.025 ;
        RECT 126.645 173.890 126.805 174.000 ;
        RECT 127.095 173.835 127.265 174.025 ;
        RECT 127.555 173.855 127.725 174.045 ;
        RECT 130.130 173.855 130.300 174.045 ;
        RECT 135.375 173.835 135.545 174.025 ;
        RECT 135.835 173.835 136.005 174.025 ;
        RECT 137.215 173.855 137.385 174.045 ;
        RECT 138.595 173.835 138.765 174.045 ;
        RECT 36.750 173.805 37.705 173.835 ;
        RECT 35.425 173.125 37.705 173.805 ;
        RECT 36.750 172.925 37.705 173.125 ;
        RECT 37.715 173.025 39.085 173.835 ;
        RECT 39.105 172.965 39.535 173.750 ;
        RECT 39.555 172.925 43.210 173.835 ;
        RECT 43.235 173.025 48.745 173.835 ;
        RECT 48.795 172.925 51.965 173.835 ;
        RECT 51.975 173.155 53.805 173.835 ;
        RECT 53.815 173.025 59.325 173.835 ;
        RECT 59.335 173.025 61.165 173.835 ;
        RECT 61.175 172.925 63.005 173.835 ;
        RECT 63.015 173.025 64.845 173.835 ;
        RECT 64.865 172.965 65.295 173.750 ;
        RECT 65.315 173.155 72.625 173.835 ;
        RECT 68.830 172.935 69.740 173.155 ;
        RECT 71.275 172.925 72.625 173.155 ;
        RECT 72.675 173.025 74.045 173.835 ;
        RECT 74.165 173.155 77.630 173.835 ;
        RECT 76.710 172.925 77.630 173.155 ;
        RECT 77.735 173.155 81.635 173.835 ;
        RECT 81.875 173.155 85.775 173.835 ;
        RECT 77.735 172.925 78.665 173.155 ;
        RECT 81.875 172.925 82.805 173.155 ;
        RECT 86.015 173.025 89.685 173.835 ;
        RECT 90.625 172.965 91.055 173.750 ;
        RECT 91.075 173.025 93.825 173.835 ;
        RECT 93.835 173.155 98.650 173.835 ;
        RECT 98.895 173.025 101.645 173.835 ;
        RECT 102.135 172.925 103.485 173.835 ;
        RECT 103.495 173.025 109.005 173.835 ;
        RECT 109.015 173.025 112.685 173.835 ;
        RECT 113.155 173.155 115.445 173.835 ;
        RECT 113.155 172.925 114.075 173.155 ;
        RECT 116.385 172.965 116.815 173.750 ;
        RECT 117.030 172.925 120.505 173.835 ;
        RECT 120.515 173.025 124.185 173.835 ;
        RECT 124.195 173.025 125.565 173.835 ;
        RECT 125.575 173.055 126.945 173.835 ;
        RECT 126.955 173.155 134.265 173.835 ;
        RECT 130.470 172.935 131.380 173.155 ;
        RECT 132.915 172.925 134.265 173.155 ;
        RECT 134.315 173.055 135.685 173.835 ;
        RECT 135.695 173.155 137.525 173.835 ;
        RECT 136.180 172.925 137.525 173.155 ;
        RECT 137.535 173.025 138.905 173.835 ;
      LAYER nwell ;
        RECT 13.140 169.805 139.100 172.635 ;
      LAYER pwell ;
        RECT 13.335 168.605 14.705 169.415 ;
        RECT 14.715 168.605 16.085 169.385 ;
        RECT 16.095 168.605 17.465 169.415 ;
        RECT 17.485 169.285 20.485 169.515 ;
        RECT 22.075 169.285 23.005 169.515 ;
        RECT 17.485 169.195 22.065 169.285 ;
        RECT 17.475 168.835 22.065 169.195 ;
        RECT 17.475 168.645 18.405 168.835 ;
        RECT 17.485 168.605 18.405 168.645 ;
        RECT 20.495 168.605 22.065 168.835 ;
        RECT 22.075 168.605 25.745 169.285 ;
        RECT 26.225 168.690 26.655 169.475 ;
        RECT 27.155 168.605 28.505 169.515 ;
        RECT 28.515 168.605 31.265 169.415 ;
        RECT 31.275 168.605 34.485 169.515 ;
        RECT 37.215 169.315 38.165 169.515 ;
        RECT 34.495 168.635 38.165 169.315 ;
        RECT 13.475 168.395 13.645 168.605 ;
        RECT 14.865 168.585 15.035 168.605 ;
        RECT 14.855 168.415 15.035 168.585 ;
        RECT 16.235 168.415 16.405 168.605 ;
        RECT 16.690 168.445 16.810 168.555 ;
        RECT 21.755 168.415 21.925 168.605 ;
        RECT 14.855 168.395 15.025 168.415 ;
        RECT 24.055 168.395 24.225 168.585 ;
        RECT 24.515 168.395 24.685 168.585 ;
        RECT 25.435 168.415 25.605 168.605 ;
        RECT 25.890 168.445 26.010 168.555 ;
        RECT 26.810 168.445 26.930 168.555 ;
        RECT 27.270 168.445 27.390 168.555 ;
        RECT 27.740 168.395 27.910 168.585 ;
        RECT 28.190 168.415 28.360 168.605 ;
        RECT 28.655 168.415 28.825 168.605 ;
        RECT 30.035 168.395 30.205 168.585 ;
        RECT 33.255 168.395 33.425 168.585 ;
        RECT 34.185 168.415 34.355 168.605 ;
        RECT 34.640 168.395 34.810 168.635 ;
        RECT 37.215 168.605 38.165 168.635 ;
        RECT 39.405 169.285 40.335 169.515 ;
        RECT 39.405 168.605 41.240 169.285 ;
        RECT 41.395 168.605 45.065 169.415 ;
        RECT 45.545 168.605 48.275 169.515 ;
        RECT 49.045 168.605 51.965 169.515 ;
        RECT 51.985 168.690 52.415 169.475 ;
        RECT 52.475 169.285 53.825 169.515 ;
        RECT 55.360 169.285 56.270 169.505 ;
        RECT 52.475 168.605 59.785 169.285 ;
        RECT 59.795 168.605 65.305 169.415 ;
        RECT 66.685 169.285 67.605 169.515 ;
        RECT 69.445 169.285 70.365 169.515 ;
        RECT 65.315 168.605 67.605 169.285 ;
        RECT 68.075 168.605 70.365 169.285 ;
        RECT 70.375 168.605 73.850 169.515 ;
        RECT 74.055 169.315 75.005 169.515 ;
        RECT 74.055 168.635 77.725 169.315 ;
        RECT 77.745 168.690 78.175 169.475 ;
        RECT 81.770 169.285 82.690 169.515 ;
        RECT 85.995 169.285 86.925 169.515 ;
        RECT 89.590 169.285 90.510 169.515 ;
        RECT 74.055 168.605 75.005 168.635 ;
        RECT 41.075 168.585 41.240 168.605 ;
        RECT 38.325 168.440 38.485 168.560 ;
        RECT 39.695 168.395 39.865 168.585 ;
        RECT 41.075 168.415 41.245 168.585 ;
        RECT 41.535 168.395 41.705 168.605 ;
        RECT 45.210 168.445 45.330 168.555 ;
        RECT 45.675 168.415 45.845 168.605 ;
        RECT 47.060 168.395 47.230 168.585 ;
        RECT 47.515 168.395 47.685 168.585 ;
        RECT 48.430 168.445 48.550 168.555 ;
        RECT 51.650 168.415 51.820 168.605 ;
        RECT 58.095 168.395 58.265 168.585 ;
        RECT 59.475 168.415 59.645 168.605 ;
        RECT 59.935 168.415 60.105 168.605 ;
        RECT 61.775 168.395 61.945 168.585 ;
        RECT 62.235 168.395 62.405 168.585 ;
        RECT 65.455 168.395 65.625 168.605 ;
        RECT 67.295 168.395 67.465 168.585 ;
        RECT 67.750 168.445 67.870 168.555 ;
        RECT 68.215 168.415 68.385 168.605 ;
        RECT 13.335 167.585 14.705 168.395 ;
        RECT 14.715 167.585 16.545 168.395 ;
        RECT 17.055 167.715 24.365 168.395 ;
        RECT 17.055 167.485 18.405 167.715 ;
        RECT 19.940 167.495 20.850 167.715 ;
        RECT 24.375 167.585 27.125 168.395 ;
        RECT 27.740 168.165 29.430 168.395 ;
        RECT 27.595 167.485 29.430 168.165 ;
        RECT 29.895 167.485 33.105 168.395 ;
        RECT 33.115 167.585 34.485 168.395 ;
        RECT 34.495 167.715 38.165 168.395 ;
        RECT 34.495 167.485 35.420 167.715 ;
        RECT 39.105 167.525 39.535 168.310 ;
        RECT 39.555 167.585 41.385 168.395 ;
        RECT 41.395 167.485 45.945 168.395 ;
        RECT 45.995 167.485 47.345 168.395 ;
        RECT 47.375 167.715 51.045 168.395 ;
        RECT 50.115 167.485 51.045 167.715 ;
        RECT 51.095 167.715 58.405 168.395 ;
        RECT 58.415 167.715 62.085 168.395 ;
        RECT 51.095 167.485 52.445 167.715 ;
        RECT 53.980 167.495 54.890 167.715 ;
        RECT 58.415 167.485 59.345 167.715 ;
        RECT 62.095 167.585 64.845 168.395 ;
        RECT 64.865 167.525 65.295 168.310 ;
        RECT 65.315 167.585 67.145 168.395 ;
        RECT 67.155 167.715 69.905 168.395 ;
        RECT 70.060 168.365 70.230 168.585 ;
        RECT 70.520 168.415 70.690 168.605 ;
        RECT 75.585 168.395 75.755 168.585 ;
        RECT 76.045 168.440 76.205 168.550 ;
        RECT 77.410 168.415 77.580 168.635 ;
        RECT 79.225 168.605 82.690 169.285 ;
        RECT 83.025 168.605 86.925 169.285 ;
        RECT 87.045 168.605 90.510 169.285 ;
        RECT 91.075 169.285 92.005 169.515 ;
        RECT 91.075 168.605 94.975 169.285 ;
        RECT 95.215 168.605 96.585 169.415 ;
        RECT 99.250 169.285 100.170 169.515 ;
        RECT 96.705 168.605 100.170 169.285 ;
        RECT 100.275 168.605 103.025 169.415 ;
        RECT 103.505 168.690 103.935 169.475 ;
        RECT 114.755 169.425 115.705 169.515 ;
        RECT 103.955 168.605 109.465 169.415 ;
        RECT 109.475 168.605 113.145 169.415 ;
        RECT 113.775 168.605 115.705 169.425 ;
        RECT 115.915 169.285 116.835 169.515 ;
        RECT 115.915 168.605 119.500 169.285 ;
        RECT 119.790 168.605 123.265 169.515 ;
        RECT 123.275 168.605 126.485 169.515 ;
        RECT 126.495 168.605 129.245 169.415 ;
        RECT 129.265 168.690 129.695 169.475 ;
        RECT 129.715 169.285 130.645 169.515 ;
        RECT 133.950 169.285 134.870 169.515 ;
        RECT 129.715 168.605 133.615 169.285 ;
        RECT 133.950 168.605 137.415 169.285 ;
        RECT 137.535 168.605 138.905 169.415 ;
        RECT 78.345 168.450 78.505 168.560 ;
        RECT 79.255 168.415 79.425 168.605 ;
        RECT 71.720 168.365 72.665 168.395 ;
        RECT 68.975 167.485 69.905 167.715 ;
        RECT 69.915 167.685 72.665 168.365 ;
        RECT 71.720 167.485 72.665 167.685 ;
        RECT 72.675 167.485 75.885 168.395 ;
        RECT 76.815 168.365 77.750 168.395 ;
        RECT 79.710 168.365 79.880 168.585 ;
        RECT 86.340 168.415 86.510 168.605 ;
        RECT 87.075 168.395 87.245 168.605 ;
        RECT 87.535 168.395 87.705 168.585 ;
        RECT 90.290 168.445 90.410 168.555 ;
        RECT 90.750 168.445 90.870 168.555 ;
        RECT 91.225 168.440 91.385 168.550 ;
        RECT 91.490 168.415 91.660 168.605 ;
        RECT 95.355 168.415 95.525 168.605 ;
        RECT 96.735 168.415 96.905 168.605 ;
        RECT 99.035 168.395 99.205 168.585 ;
        RECT 99.495 168.395 99.665 168.585 ;
        RECT 100.415 168.415 100.585 168.605 ;
        RECT 102.715 168.395 102.885 168.585 ;
        RECT 103.170 168.445 103.290 168.555 ;
        RECT 104.095 168.415 104.265 168.605 ;
        RECT 109.615 168.585 109.785 168.605 ;
        RECT 113.775 168.585 113.925 168.605 ;
        RECT 104.550 168.445 104.670 168.555 ;
        RECT 105.015 168.415 105.185 168.585 ;
        RECT 105.035 168.395 105.185 168.415 ;
        RECT 108.235 168.395 108.405 168.585 ;
        RECT 109.615 168.415 109.790 168.585 ;
        RECT 109.620 168.395 109.790 168.415 ;
        RECT 110.990 168.395 111.160 168.585 ;
        RECT 112.380 168.395 112.550 168.585 ;
        RECT 112.845 168.440 113.005 168.550 ;
        RECT 113.290 168.445 113.410 168.555 ;
        RECT 113.755 168.415 113.925 168.585 ;
        RECT 116.060 168.415 116.230 168.605 ;
        RECT 113.905 168.395 113.925 168.415 ;
        RECT 76.815 168.165 79.880 168.365 ;
        RECT 76.815 167.685 80.025 168.165 ;
        RECT 76.815 167.485 77.765 167.685 ;
        RECT 79.095 167.485 80.025 167.685 ;
        RECT 80.075 167.715 87.385 168.395 ;
        RECT 80.075 167.485 81.425 167.715 ;
        RECT 82.960 167.495 83.870 167.715 ;
        RECT 87.395 167.585 90.145 168.395 ;
        RECT 90.625 167.525 91.055 168.310 ;
        RECT 92.035 167.715 99.345 168.395 ;
        RECT 92.035 167.485 93.385 167.715 ;
        RECT 94.920 167.495 95.830 167.715 ;
        RECT 99.355 167.485 102.565 168.395 ;
        RECT 102.575 167.585 104.405 168.395 ;
        RECT 105.035 167.575 106.965 168.395 ;
        RECT 106.015 167.485 106.965 167.575 ;
        RECT 107.185 167.485 108.535 168.395 ;
        RECT 108.555 167.485 109.905 168.395 ;
        RECT 109.955 167.485 111.305 168.395 ;
        RECT 111.315 167.485 112.665 168.395 ;
        RECT 113.905 167.715 116.355 168.395 ;
        RECT 116.970 168.365 117.140 168.585 ;
        RECT 119.275 168.395 119.445 168.585 ;
        RECT 122.950 168.415 123.120 168.605 ;
        RECT 123.415 168.415 123.585 168.605 ;
        RECT 125.260 168.395 125.430 168.585 ;
        RECT 125.725 168.440 125.885 168.550 ;
        RECT 126.635 168.395 126.805 168.605 ;
        RECT 130.130 168.415 130.300 168.605 ;
        RECT 133.995 168.395 134.165 168.585 ;
        RECT 135.835 168.395 136.005 168.585 ;
        RECT 137.215 168.415 137.385 168.605 ;
        RECT 138.595 168.395 138.765 168.605 ;
        RECT 118.170 168.365 119.125 168.395 ;
        RECT 114.395 167.485 116.355 167.715 ;
        RECT 116.385 167.525 116.815 168.310 ;
        RECT 116.845 167.685 119.125 168.365 ;
        RECT 119.135 167.715 123.950 168.395 ;
        RECT 118.170 167.485 119.125 167.685 ;
        RECT 124.195 167.485 125.545 168.395 ;
        RECT 126.495 167.715 133.805 168.395 ;
        RECT 133.855 167.715 135.685 168.395 ;
        RECT 135.695 167.715 137.525 168.395 ;
        RECT 130.010 167.495 130.920 167.715 ;
        RECT 132.455 167.485 133.805 167.715 ;
        RECT 134.340 167.485 135.685 167.715 ;
        RECT 136.180 167.485 137.525 167.715 ;
        RECT 137.535 167.585 138.905 168.395 ;
      LAYER nwell ;
        RECT 13.140 164.365 139.100 167.195 ;
      LAYER pwell ;
        RECT 13.335 163.165 14.705 163.975 ;
        RECT 19.150 163.845 20.060 164.065 ;
        RECT 21.595 163.845 22.945 164.075 ;
        RECT 15.635 163.165 22.945 163.845 ;
        RECT 22.995 163.165 25.745 163.975 ;
        RECT 26.225 163.250 26.655 164.035 ;
        RECT 26.685 163.165 29.425 163.845 ;
        RECT 29.435 163.165 34.945 163.975 ;
        RECT 34.955 163.165 37.705 164.075 ;
        RECT 37.715 163.165 39.545 163.975 ;
        RECT 39.555 163.875 40.500 164.075 ;
        RECT 39.555 163.195 42.305 163.875 ;
        RECT 39.555 163.165 40.500 163.195 ;
        RECT 13.475 162.955 13.645 163.165 ;
        RECT 14.855 162.955 15.025 163.145 ;
        RECT 15.775 162.975 15.945 163.165 ;
        RECT 20.375 162.955 20.545 163.145 ;
        RECT 22.210 163.005 22.330 163.115 ;
        RECT 22.675 162.955 22.845 163.145 ;
        RECT 23.135 162.975 23.305 163.165 ;
        RECT 29.115 163.145 29.285 163.165 ;
        RECT 25.895 163.115 26.065 163.145 ;
        RECT 25.890 163.005 26.065 163.115 ;
        RECT 28.650 163.005 28.770 163.115 ;
        RECT 25.895 162.955 26.065 163.005 ;
        RECT 29.115 162.975 29.290 163.145 ;
        RECT 29.575 162.975 29.745 163.165 ;
        RECT 29.120 162.955 29.290 162.975 ;
        RECT 31.415 162.955 31.585 163.145 ;
        RECT 35.095 162.975 35.265 163.165 ;
        RECT 36.935 162.955 37.105 163.145 ;
        RECT 37.855 162.975 38.025 163.165 ;
        RECT 38.770 163.005 38.890 163.115 ;
        RECT 39.695 162.955 39.865 163.145 ;
        RECT 41.070 163.005 41.190 163.115 ;
        RECT 41.535 162.955 41.705 163.145 ;
        RECT 41.990 162.975 42.160 163.195 ;
        RECT 42.445 163.165 45.445 164.075 ;
        RECT 45.535 163.165 46.885 164.075 ;
        RECT 50.575 163.845 51.505 164.075 ;
        RECT 47.835 163.165 51.505 163.845 ;
        RECT 51.985 163.250 52.415 164.035 ;
        RECT 52.475 163.845 53.825 164.075 ;
        RECT 55.360 163.845 56.270 164.065 ;
        RECT 68.075 163.875 69.005 164.075 ;
        RECT 70.335 163.875 71.285 164.075 ;
        RECT 52.475 163.165 59.785 163.845 ;
        RECT 60.255 163.165 62.995 163.845 ;
        RECT 63.015 163.165 67.830 163.845 ;
        RECT 68.075 163.395 71.285 163.875 ;
        RECT 73.115 163.845 74.045 164.075 ;
        RECT 76.710 163.845 77.630 164.075 ;
        RECT 68.220 163.195 71.285 163.395 ;
        RECT 13.335 162.145 14.705 162.955 ;
        RECT 14.715 162.145 20.225 162.955 ;
        RECT 20.235 162.145 22.065 162.955 ;
        RECT 22.575 162.045 25.745 162.955 ;
        RECT 25.755 162.145 28.505 162.955 ;
        RECT 29.120 162.725 30.810 162.955 ;
        RECT 28.975 162.045 30.810 162.725 ;
        RECT 31.275 162.145 36.785 162.955 ;
        RECT 36.795 162.145 38.625 162.955 ;
        RECT 39.105 162.085 39.535 162.870 ;
        RECT 39.565 162.045 40.915 162.955 ;
        RECT 41.495 162.045 44.605 162.955 ;
        RECT 44.760 162.925 44.930 163.145 ;
        RECT 45.215 162.975 45.385 163.165 ;
        RECT 45.680 162.975 45.850 163.165 ;
        RECT 47.065 163.010 47.225 163.120 ;
        RECT 47.515 162.955 47.685 163.145 ;
        RECT 47.975 162.975 48.145 163.165 ;
        RECT 51.650 163.005 51.770 163.115 ;
        RECT 52.115 162.955 52.285 163.145 ;
        RECT 52.575 162.955 52.745 163.145 ;
        RECT 58.095 162.955 58.265 163.145 ;
        RECT 59.475 162.975 59.645 163.165 ;
        RECT 59.930 163.005 60.050 163.115 ;
        RECT 60.395 162.975 60.565 163.165 ;
        RECT 63.155 162.975 63.325 163.165 ;
        RECT 63.615 162.955 63.785 163.145 ;
        RECT 65.455 162.955 65.625 163.145 ;
        RECT 68.220 162.975 68.390 163.195 ;
        RECT 70.350 163.165 71.285 163.195 ;
        RECT 71.295 163.165 74.045 163.845 ;
        RECT 74.165 163.165 77.630 163.845 ;
        RECT 77.745 163.250 78.175 164.035 ;
        RECT 78.235 163.845 79.585 164.075 ;
        RECT 81.120 163.845 82.030 164.065 ;
        RECT 85.555 163.845 86.485 164.075 ;
        RECT 78.235 163.165 85.545 163.845 ;
        RECT 85.555 163.165 89.455 163.845 ;
        RECT 89.695 163.165 91.525 163.975 ;
        RECT 97.055 163.845 97.985 164.075 ;
        RECT 91.995 163.165 96.810 163.845 ;
        RECT 97.055 163.165 100.955 163.845 ;
        RECT 101.195 163.165 103.025 163.975 ;
        RECT 103.505 163.250 103.935 164.035 ;
        RECT 103.955 163.165 105.785 164.075 ;
        RECT 106.265 163.165 107.615 164.075 ;
        RECT 107.635 163.165 111.305 163.975 ;
        RECT 111.925 163.165 115.580 164.075 ;
        RECT 115.915 163.165 117.745 164.075 ;
        RECT 118.215 163.165 129.225 164.075 ;
        RECT 129.265 163.250 129.695 164.035 ;
        RECT 129.715 163.845 130.645 164.075 ;
        RECT 133.950 163.845 134.870 164.075 ;
        RECT 129.715 163.165 133.615 163.845 ;
        RECT 133.950 163.165 137.415 163.845 ;
        RECT 137.535 163.165 138.905 163.975 ;
        RECT 71.435 162.975 71.605 163.165 ;
        RECT 74.195 162.975 74.365 163.165 ;
        RECT 76.035 162.955 76.205 163.145 ;
        RECT 76.495 162.955 76.665 163.145 ;
        RECT 85.235 162.955 85.405 163.165 ;
        RECT 85.970 162.955 86.140 163.165 ;
        RECT 89.835 162.975 90.005 163.165 ;
        RECT 91.225 163.000 91.385 163.110 ;
        RECT 91.670 163.005 91.790 163.115 ;
        RECT 92.135 162.955 92.305 163.165 ;
        RECT 97.470 162.955 97.640 163.165 ;
        RECT 101.335 162.975 101.505 163.165 ;
        RECT 101.610 162.955 101.780 163.145 ;
        RECT 103.170 163.005 103.290 163.115 ;
        RECT 104.100 162.975 104.270 163.165 ;
        RECT 105.930 163.005 106.050 163.115 ;
        RECT 106.395 162.975 106.565 163.165 ;
        RECT 107.775 162.975 107.945 163.165 ;
        RECT 111.925 163.145 112.085 163.165 ;
        RECT 108.695 162.955 108.865 163.145 ;
        RECT 109.155 162.955 109.325 163.145 ;
        RECT 111.450 163.005 111.570 163.115 ;
        RECT 111.915 162.975 112.085 163.145 ;
        RECT 112.380 162.955 112.550 163.145 ;
        RECT 115.605 163.000 115.765 163.110 ;
        RECT 116.060 162.975 116.230 163.165 ;
        RECT 46.420 162.925 47.365 162.955 ;
        RECT 44.615 162.245 47.365 162.925 ;
        RECT 46.420 162.045 47.365 162.245 ;
        RECT 47.375 162.145 49.205 162.955 ;
        RECT 49.215 162.045 52.325 162.955 ;
        RECT 52.435 162.145 57.945 162.955 ;
        RECT 57.955 162.145 63.465 162.955 ;
        RECT 63.475 162.145 64.845 162.955 ;
        RECT 64.865 162.085 65.295 162.870 ;
        RECT 65.315 162.275 72.625 162.955 ;
        RECT 68.830 162.055 69.740 162.275 ;
        RECT 71.275 162.045 72.625 162.275 ;
        RECT 72.770 162.275 76.235 162.955 ;
        RECT 72.770 162.045 73.690 162.275 ;
        RECT 76.355 162.145 78.185 162.955 ;
        RECT 78.235 162.275 85.545 162.955 ;
        RECT 85.555 162.275 89.455 162.955 ;
        RECT 78.235 162.045 79.585 162.275 ;
        RECT 81.120 162.055 82.030 162.275 ;
        RECT 85.555 162.045 86.485 162.275 ;
        RECT 90.625 162.085 91.055 162.870 ;
        RECT 91.995 162.275 96.810 162.955 ;
        RECT 97.055 162.275 100.955 162.955 ;
        RECT 101.195 162.275 105.095 162.955 ;
        RECT 105.430 162.275 108.895 162.955 ;
        RECT 97.055 162.045 97.985 162.275 ;
        RECT 101.195 162.045 102.125 162.275 ;
        RECT 105.430 162.045 106.350 162.275 ;
        RECT 109.015 162.045 112.225 162.955 ;
        RECT 112.235 162.045 115.155 162.955 ;
        RECT 116.970 162.925 117.140 163.145 ;
        RECT 117.890 163.005 118.010 163.115 ;
        RECT 118.360 162.975 118.530 163.165 ;
        RECT 119.275 162.955 119.445 163.145 ;
        RECT 124.335 162.975 124.505 163.145 ;
        RECT 124.340 162.955 124.505 162.975 ;
        RECT 126.635 162.955 126.805 163.145 ;
        RECT 130.130 162.975 130.300 163.165 ;
        RECT 133.995 162.955 134.165 163.145 ;
        RECT 135.370 163.005 135.490 163.115 ;
        RECT 135.835 162.955 136.005 163.145 ;
        RECT 137.215 162.975 137.385 163.165 ;
        RECT 138.595 162.955 138.765 163.165 ;
        RECT 118.170 162.925 119.125 162.955 ;
        RECT 116.385 162.085 116.815 162.870 ;
        RECT 116.845 162.245 119.125 162.925 ;
        RECT 119.135 162.275 123.950 162.955 ;
        RECT 124.340 162.275 126.175 162.955 ;
        RECT 126.495 162.275 133.805 162.955 ;
        RECT 118.170 162.045 119.125 162.245 ;
        RECT 125.245 162.045 126.175 162.275 ;
        RECT 130.010 162.055 130.920 162.275 ;
        RECT 132.455 162.045 133.805 162.275 ;
        RECT 133.855 162.175 135.225 162.955 ;
        RECT 135.695 162.275 137.525 162.955 ;
        RECT 136.180 162.045 137.525 162.275 ;
        RECT 137.535 162.145 138.905 162.955 ;
      LAYER nwell ;
        RECT 13.140 158.925 139.100 161.755 ;
      LAYER pwell ;
        RECT 13.335 157.725 14.705 158.535 ;
        RECT 14.715 157.725 20.225 158.535 ;
        RECT 20.235 157.725 25.745 158.535 ;
        RECT 26.225 157.810 26.655 158.595 ;
        RECT 26.675 157.725 32.185 158.535 ;
        RECT 32.195 157.725 34.025 158.535 ;
        RECT 34.090 157.725 44.110 158.635 ;
        RECT 44.155 157.725 49.665 158.535 ;
        RECT 49.675 157.725 51.505 158.535 ;
        RECT 51.985 157.810 52.415 158.595 ;
        RECT 52.435 157.725 57.945 158.535 ;
        RECT 57.955 157.725 63.465 158.535 ;
        RECT 63.475 157.725 66.225 158.535 ;
        RECT 66.695 158.405 67.625 158.635 ;
        RECT 66.695 157.725 70.595 158.405 ;
        RECT 70.835 157.725 72.205 158.535 ;
        RECT 72.310 158.405 73.230 158.635 ;
        RECT 72.310 157.725 75.775 158.405 ;
        RECT 75.895 157.725 77.725 158.535 ;
        RECT 77.745 157.810 78.175 158.595 ;
        RECT 78.195 157.725 83.705 158.535 ;
        RECT 83.715 157.725 85.085 158.535 ;
        RECT 88.295 158.405 89.225 158.635 ;
        RECT 85.325 157.725 89.225 158.405 ;
        RECT 89.235 157.725 91.985 158.535 ;
        RECT 95.970 158.405 96.880 158.625 ;
        RECT 98.415 158.405 99.765 158.635 ;
        RECT 92.455 157.725 99.765 158.405 ;
        RECT 99.815 157.725 103.485 158.535 ;
        RECT 103.505 157.810 103.935 158.595 ;
        RECT 106.610 158.405 107.530 158.635 ;
        RECT 104.065 157.725 107.530 158.405 ;
        RECT 107.635 157.725 109.465 158.635 ;
        RECT 109.495 157.725 110.845 158.635 ;
        RECT 114.430 158.405 115.350 158.635 ;
        RECT 111.885 157.725 115.350 158.405 ;
        RECT 115.455 157.725 118.665 158.635 ;
        RECT 128.315 158.405 129.245 158.635 ;
        RECT 119.135 157.725 123.950 158.405 ;
        RECT 125.345 157.725 129.245 158.405 ;
        RECT 129.265 157.810 129.695 158.595 ;
        RECT 133.230 158.405 134.140 158.625 ;
        RECT 135.675 158.405 137.025 158.635 ;
        RECT 129.715 157.725 137.025 158.405 ;
        RECT 137.535 157.725 138.905 158.535 ;
        RECT 13.475 157.515 13.645 157.725 ;
        RECT 14.855 157.515 15.025 157.725 ;
        RECT 16.695 157.515 16.865 157.705 ;
        RECT 19.455 157.515 19.625 157.705 ;
        RECT 20.375 157.535 20.545 157.725 ;
        RECT 25.890 157.565 26.010 157.675 ;
        RECT 26.815 157.535 26.985 157.725 ;
        RECT 30.950 157.515 31.120 157.705 ;
        RECT 31.415 157.515 31.585 157.705 ;
        RECT 32.335 157.535 32.505 157.725 ;
        RECT 34.175 157.535 34.345 157.725 ;
        RECT 35.105 157.560 35.265 157.670 ;
        RECT 36.015 157.515 36.185 157.705 ;
        RECT 38.770 157.565 38.890 157.675 ;
        RECT 39.695 157.535 39.865 157.705 ;
        RECT 39.700 157.515 39.865 157.535 ;
        RECT 41.995 157.515 42.165 157.705 ;
        RECT 44.295 157.535 44.465 157.725 ;
        RECT 47.515 157.515 47.685 157.705 ;
        RECT 49.815 157.535 49.985 157.725 ;
        RECT 51.650 157.565 51.770 157.675 ;
        RECT 52.575 157.535 52.745 157.725 ;
        RECT 53.035 157.515 53.205 157.705 ;
        RECT 58.095 157.535 58.265 157.725 ;
        RECT 58.555 157.515 58.725 157.705 ;
        RECT 63.615 157.535 63.785 157.725 ;
        RECT 64.085 157.560 64.245 157.670 ;
        RECT 65.455 157.515 65.625 157.705 ;
        RECT 66.370 157.565 66.490 157.675 ;
        RECT 67.110 157.535 67.280 157.725 ;
        RECT 70.975 157.535 71.145 157.725 ;
        RECT 73.090 157.515 73.260 157.705 ;
        RECT 75.575 157.535 75.745 157.725 ;
        RECT 76.035 157.535 76.205 157.725 ;
        RECT 78.335 157.535 78.505 157.725 ;
        RECT 80.175 157.515 80.345 157.705 ;
        RECT 80.635 157.515 80.805 157.705 ;
        RECT 83.855 157.535 84.025 157.725 ;
        RECT 86.155 157.515 86.325 157.705 ;
        RECT 88.640 157.535 88.810 157.725 ;
        RECT 89.375 157.535 89.545 157.725 ;
        RECT 89.845 157.560 90.005 157.670 ;
        RECT 91.215 157.515 91.385 157.705 ;
        RECT 92.130 157.565 92.250 157.675 ;
        RECT 92.595 157.515 92.765 157.725 ;
        RECT 99.955 157.535 100.125 157.725 ;
        RECT 104.095 157.535 104.265 157.725 ;
        RECT 107.780 157.705 107.950 157.725 ;
        RECT 107.775 157.535 107.950 157.705 ;
        RECT 108.245 157.560 108.405 157.670 ;
        RECT 109.610 157.535 109.780 157.725 ;
        RECT 111.005 157.570 111.165 157.680 ;
        RECT 111.915 157.535 112.085 157.725 ;
        RECT 107.775 157.515 107.945 157.535 ;
        RECT 116.055 157.515 116.225 157.705 ;
        RECT 116.970 157.515 117.140 157.705 ;
        RECT 118.355 157.535 118.525 157.725 ;
        RECT 118.810 157.565 118.930 157.675 ;
        RECT 119.275 157.515 119.445 157.725 ;
        RECT 122.495 157.515 122.665 157.705 ;
        RECT 124.345 157.570 124.505 157.680 ;
        RECT 125.715 157.515 125.885 157.705 ;
        RECT 128.660 157.535 128.830 157.725 ;
        RECT 128.935 157.515 129.105 157.705 ;
        RECT 129.855 157.535 130.025 157.725 ;
        RECT 130.775 157.515 130.945 157.705 ;
        RECT 135.375 157.515 135.545 157.705 ;
        RECT 135.835 157.515 136.005 157.705 ;
        RECT 137.210 157.565 137.330 157.675 ;
        RECT 138.595 157.515 138.765 157.725 ;
        RECT 13.335 156.705 14.705 157.515 ;
        RECT 14.715 156.835 16.545 157.515 ;
        RECT 15.200 156.605 16.545 156.835 ;
        RECT 16.555 156.705 19.305 157.515 ;
        RECT 19.315 156.835 26.625 157.515 ;
        RECT 27.595 156.835 31.265 157.515 ;
        RECT 22.830 156.615 23.740 156.835 ;
        RECT 25.275 156.605 26.625 156.835 ;
        RECT 30.340 156.605 31.265 156.835 ;
        RECT 31.275 156.705 34.945 157.515 ;
        RECT 35.875 156.835 38.625 157.515 ;
        RECT 37.695 156.605 38.625 156.835 ;
        RECT 39.105 156.645 39.535 157.430 ;
        RECT 39.700 156.835 41.535 157.515 ;
        RECT 40.605 156.605 41.535 156.835 ;
        RECT 41.855 156.705 47.365 157.515 ;
        RECT 47.375 156.705 52.885 157.515 ;
        RECT 52.895 156.705 58.405 157.515 ;
        RECT 58.415 156.705 63.925 157.515 ;
        RECT 64.865 156.645 65.295 157.430 ;
        RECT 65.315 156.835 72.625 157.515 ;
        RECT 68.830 156.615 69.740 156.835 ;
        RECT 71.275 156.605 72.625 156.835 ;
        RECT 72.675 156.835 76.575 157.515 ;
        RECT 76.910 156.835 80.375 157.515 ;
        RECT 72.675 156.605 73.605 156.835 ;
        RECT 76.910 156.605 77.830 156.835 ;
        RECT 80.495 156.705 86.005 157.515 ;
        RECT 86.015 156.705 89.685 157.515 ;
        RECT 90.625 156.645 91.055 157.430 ;
        RECT 91.075 156.705 92.445 157.515 ;
        RECT 92.455 156.835 99.765 157.515 ;
        RECT 95.970 156.615 96.880 156.835 ;
        RECT 98.415 156.605 99.765 156.835 ;
        RECT 100.775 156.835 108.085 157.515 ;
        RECT 109.055 156.835 116.365 157.515 ;
        RECT 100.775 156.605 102.125 156.835 ;
        RECT 103.660 156.615 104.570 156.835 ;
        RECT 109.055 156.605 110.405 156.835 ;
        RECT 111.940 156.615 112.850 156.835 ;
        RECT 116.385 156.645 116.815 157.430 ;
        RECT 116.855 156.605 118.205 157.515 ;
        RECT 119.135 156.605 122.345 157.515 ;
        RECT 122.355 156.605 125.565 157.515 ;
        RECT 125.575 156.605 128.785 157.515 ;
        RECT 128.795 156.705 130.625 157.515 ;
        RECT 130.635 156.735 132.005 157.515 ;
        RECT 132.110 156.835 135.575 157.515 ;
        RECT 135.695 156.835 137.525 157.515 ;
        RECT 132.110 156.605 133.030 156.835 ;
        RECT 136.180 156.605 137.525 156.835 ;
        RECT 137.535 156.705 138.905 157.515 ;
      LAYER nwell ;
        RECT 13.140 153.485 139.100 156.315 ;
      LAYER pwell ;
        RECT 13.335 152.285 14.705 153.095 ;
        RECT 14.715 152.285 16.545 152.965 ;
        RECT 16.555 152.285 18.385 153.095 ;
        RECT 18.415 152.285 19.765 153.195 ;
        RECT 19.775 152.965 20.695 153.195 ;
        RECT 19.775 152.285 22.065 152.965 ;
        RECT 22.075 152.285 23.425 153.195 ;
        RECT 23.765 152.965 24.695 153.195 ;
        RECT 23.765 152.285 25.600 152.965 ;
        RECT 26.225 152.370 26.655 153.155 ;
        RECT 26.675 152.965 27.810 153.195 ;
        RECT 26.675 152.285 29.885 152.965 ;
        RECT 29.895 152.285 33.565 153.095 ;
        RECT 34.950 152.515 36.785 153.195 ;
        RECT 34.950 152.285 36.640 152.515 ;
        RECT 36.795 152.285 39.545 153.095 ;
        RECT 41.880 152.965 43.225 153.195 ;
        RECT 39.555 152.285 41.385 152.965 ;
        RECT 41.395 152.285 43.225 152.965 ;
        RECT 43.235 152.285 48.745 153.095 ;
        RECT 48.755 152.285 51.505 153.095 ;
        RECT 51.985 152.370 52.415 153.155 ;
        RECT 52.435 152.285 54.265 153.095 ;
        RECT 54.275 152.285 56.105 152.965 ;
        RECT 56.115 152.285 57.945 152.965 ;
        RECT 57.975 152.285 59.325 153.195 ;
        RECT 59.335 152.285 62.085 153.095 ;
        RECT 62.595 152.965 63.945 153.195 ;
        RECT 65.480 152.965 66.390 153.185 ;
        RECT 69.915 152.965 70.845 153.195 ;
        RECT 62.595 152.285 69.905 152.965 ;
        RECT 69.915 152.285 73.815 152.965 ;
        RECT 74.065 152.285 76.805 152.965 ;
        RECT 77.745 152.370 78.175 153.155 ;
        RECT 78.195 152.285 80.025 153.095 ;
        RECT 80.035 152.965 80.965 153.195 ;
        RECT 86.830 152.965 87.750 153.195 ;
        RECT 80.035 152.285 83.935 152.965 ;
        RECT 84.285 152.285 87.750 152.965 ;
        RECT 87.855 152.285 93.365 153.095 ;
        RECT 93.375 152.285 94.745 153.095 ;
        RECT 94.755 152.965 95.685 153.195 ;
        RECT 98.895 152.965 99.825 153.195 ;
        RECT 94.755 152.285 98.655 152.965 ;
        RECT 98.895 152.285 102.795 152.965 ;
        RECT 103.505 152.370 103.935 153.155 ;
        RECT 107.070 152.965 107.990 153.195 ;
        RECT 104.525 152.285 107.990 152.965 ;
        RECT 108.105 152.285 109.455 153.195 ;
        RECT 110.395 152.285 111.745 153.195 ;
        RECT 111.775 152.285 115.445 153.095 ;
        RECT 118.655 152.965 119.585 153.195 ;
        RECT 115.685 152.285 119.585 152.965 ;
        RECT 119.595 152.965 120.940 153.195 ;
        RECT 125.410 152.965 126.320 153.185 ;
        RECT 127.855 152.965 129.205 153.195 ;
        RECT 119.595 152.285 121.425 152.965 ;
        RECT 121.895 152.285 129.205 152.965 ;
        RECT 129.265 152.370 129.695 153.155 ;
        RECT 129.810 152.965 130.730 153.195 ;
        RECT 134.340 152.965 135.685 153.195 ;
        RECT 136.180 152.965 137.525 153.195 ;
        RECT 129.810 152.285 133.275 152.965 ;
        RECT 133.855 152.285 135.685 152.965 ;
        RECT 135.695 152.285 137.525 152.965 ;
        RECT 137.535 152.285 138.905 153.095 ;
        RECT 13.475 152.075 13.645 152.285 ;
        RECT 14.855 152.075 15.025 152.285 ;
        RECT 16.695 152.095 16.865 152.285 ;
        RECT 13.335 151.265 14.705 152.075 ;
        RECT 14.715 151.265 16.545 152.075 ;
        RECT 16.555 152.045 17.490 152.075 ;
        RECT 19.450 152.045 19.620 152.285 ;
        RECT 19.915 152.075 20.085 152.265 ;
        RECT 21.755 152.095 21.925 152.285 ;
        RECT 22.220 152.095 22.390 152.285 ;
        RECT 25.435 152.265 25.600 152.285 ;
        RECT 23.135 152.075 23.305 152.265 ;
        RECT 25.435 152.095 25.605 152.265 ;
        RECT 25.890 152.125 26.010 152.235 ;
        RECT 29.575 152.095 29.745 152.285 ;
        RECT 30.035 152.095 30.205 152.285 ;
        RECT 30.495 152.075 30.665 152.265 ;
        RECT 33.710 152.240 33.880 152.265 ;
        RECT 31.885 152.120 32.045 152.230 ;
        RECT 33.710 152.130 33.885 152.240 ;
        RECT 33.710 152.075 33.880 152.130 ;
        RECT 34.175 152.075 34.345 152.265 ;
        RECT 36.470 152.095 36.640 152.285 ;
        RECT 36.935 152.095 37.105 152.285 ;
        RECT 37.395 152.075 37.565 152.265 ;
        RECT 39.695 152.075 39.865 152.265 ;
        RECT 41.075 152.095 41.245 152.285 ;
        RECT 41.535 152.095 41.705 152.285 ;
        RECT 41.995 152.075 42.165 152.265 ;
        RECT 43.375 152.095 43.545 152.285 ;
        RECT 47.515 152.075 47.685 152.265 ;
        RECT 48.895 152.095 49.065 152.285 ;
        RECT 51.650 152.125 51.770 152.235 ;
        RECT 52.575 152.095 52.745 152.285 ;
        RECT 55.795 152.095 55.965 152.285 ;
        RECT 57.175 152.075 57.345 152.265 ;
        RECT 57.635 152.075 57.805 152.285 ;
        RECT 58.090 152.095 58.260 152.285 ;
        RECT 59.475 152.095 59.645 152.285 ;
        RECT 62.230 152.125 62.350 152.235 ;
        RECT 65.450 152.125 65.570 152.235 ;
        RECT 65.920 152.075 66.090 152.265 ;
        RECT 69.595 152.095 69.765 152.285 ;
        RECT 70.330 152.095 70.500 152.285 ;
        RECT 76.035 152.075 76.205 152.265 ;
        RECT 76.495 152.075 76.665 152.285 ;
        RECT 76.965 152.130 77.125 152.240 ;
        RECT 78.335 152.095 78.505 152.285 ;
        RECT 80.450 152.095 80.620 152.285 ;
        RECT 84.130 152.075 84.300 152.265 ;
        RECT 84.315 152.095 84.485 152.285 ;
        RECT 87.995 152.075 88.165 152.285 ;
        RECT 91.490 152.075 91.660 152.265 ;
        RECT 93.515 152.095 93.685 152.285 ;
        RECT 95.170 152.095 95.340 152.285 ;
        RECT 98.575 152.075 98.745 152.265 ;
        RECT 99.035 152.075 99.205 152.265 ;
        RECT 99.310 152.095 99.480 152.285 ;
        RECT 103.170 152.125 103.290 152.235 ;
        RECT 104.090 152.125 104.210 152.235 ;
        RECT 104.555 152.075 104.725 152.285 ;
        RECT 108.235 152.095 108.405 152.285 ;
        RECT 109.625 152.130 109.785 152.240 ;
        RECT 110.075 152.075 110.245 152.265 ;
        RECT 111.460 152.095 111.630 152.285 ;
        RECT 111.915 152.095 112.085 152.285 ;
        RECT 115.605 152.120 115.765 152.230 ;
        RECT 116.985 152.120 117.145 152.230 ;
        RECT 117.890 152.075 118.060 152.265 ;
        RECT 119.000 152.095 119.170 152.285 ;
        RECT 119.275 152.075 119.445 152.265 ;
        RECT 121.115 152.095 121.285 152.285 ;
        RECT 121.570 152.125 121.690 152.235 ;
        RECT 122.035 152.095 122.205 152.285 ;
        RECT 122.955 152.075 123.125 152.265 ;
        RECT 124.610 152.075 124.780 152.265 ;
        RECT 128.475 152.075 128.645 152.265 ;
        RECT 132.150 152.125 132.270 152.235 ;
        RECT 132.615 152.075 132.785 152.265 ;
        RECT 133.075 152.095 133.245 152.285 ;
        RECT 133.530 152.125 133.650 152.235 ;
        RECT 133.995 152.075 134.165 152.285 ;
        RECT 135.835 152.095 136.005 152.285 ;
        RECT 138.595 152.075 138.765 152.285 ;
        RECT 16.555 151.845 19.620 152.045 ;
        RECT 16.555 151.365 19.765 151.845 ;
        RECT 19.775 151.395 22.985 152.075 ;
        RECT 22.995 151.395 30.305 152.075 ;
        RECT 16.555 151.165 17.505 151.365 ;
        RECT 18.835 151.165 19.765 151.365 ;
        RECT 21.850 151.165 22.985 151.395 ;
        RECT 26.510 151.175 27.420 151.395 ;
        RECT 28.955 151.165 30.305 151.395 ;
        RECT 30.365 151.165 31.715 152.075 ;
        RECT 32.675 151.165 34.025 152.075 ;
        RECT 34.035 151.165 37.245 152.075 ;
        RECT 37.255 151.265 39.085 152.075 ;
        RECT 39.105 151.205 39.535 151.990 ;
        RECT 39.555 151.165 41.845 152.075 ;
        RECT 41.855 151.265 47.365 152.075 ;
        RECT 47.375 151.265 50.125 152.075 ;
        RECT 50.175 151.395 57.485 152.075 ;
        RECT 57.495 151.395 64.805 152.075 ;
        RECT 50.175 151.165 51.525 151.395 ;
        RECT 53.060 151.175 53.970 151.395 ;
        RECT 61.010 151.175 61.920 151.395 ;
        RECT 63.455 151.165 64.805 151.395 ;
        RECT 64.865 151.205 65.295 151.990 ;
        RECT 65.775 151.165 68.890 152.075 ;
        RECT 69.035 151.395 76.345 152.075 ;
        RECT 76.355 151.395 83.665 152.075 ;
        RECT 69.035 151.165 70.385 151.395 ;
        RECT 71.920 151.175 72.830 151.395 ;
        RECT 79.870 151.175 80.780 151.395 ;
        RECT 82.315 151.165 83.665 151.395 ;
        RECT 83.715 151.395 87.615 152.075 ;
        RECT 83.715 151.165 84.645 151.395 ;
        RECT 87.855 151.265 90.605 152.075 ;
        RECT 90.625 151.205 91.055 151.990 ;
        RECT 91.075 151.395 94.975 152.075 ;
        RECT 95.310 151.395 98.775 152.075 ;
        RECT 91.075 151.165 92.005 151.395 ;
        RECT 95.310 151.165 96.230 151.395 ;
        RECT 98.895 151.265 104.405 152.075 ;
        RECT 104.415 151.265 109.925 152.075 ;
        RECT 109.935 151.265 115.445 152.075 ;
        RECT 116.385 151.205 116.815 151.990 ;
        RECT 117.775 151.165 119.125 152.075 ;
        RECT 119.135 151.265 122.805 152.075 ;
        RECT 122.815 151.265 124.185 152.075 ;
        RECT 124.195 151.395 128.095 152.075 ;
        RECT 124.195 151.165 125.125 151.395 ;
        RECT 128.335 151.265 132.005 152.075 ;
        RECT 132.475 151.295 133.845 152.075 ;
        RECT 133.855 151.265 137.525 152.075 ;
        RECT 137.535 151.265 138.905 152.075 ;
      LAYER nwell ;
        RECT 13.140 148.045 139.100 150.875 ;
      LAYER pwell ;
        RECT 13.335 146.845 14.705 147.655 ;
        RECT 14.715 146.845 16.545 147.655 ;
        RECT 20.070 147.525 20.980 147.745 ;
        RECT 22.515 147.525 23.865 147.755 ;
        RECT 16.555 146.845 23.865 147.525 ;
        RECT 24.115 147.665 25.065 147.755 ;
        RECT 24.115 146.845 26.045 147.665 ;
        RECT 26.225 146.930 26.655 147.715 ;
        RECT 26.675 146.845 28.025 147.755 ;
        RECT 28.055 147.555 28.985 147.755 ;
        RECT 30.320 147.555 31.265 147.755 ;
        RECT 28.055 147.075 31.265 147.555 ;
        RECT 28.195 146.875 31.265 147.075 ;
        RECT 13.475 146.635 13.645 146.845 ;
        RECT 14.855 146.655 15.025 146.845 ;
        RECT 15.775 146.635 15.945 146.825 ;
        RECT 16.695 146.655 16.865 146.845 ;
        RECT 25.895 146.825 26.045 146.845 ;
        RECT 23.140 146.635 23.310 146.825 ;
        RECT 24.520 146.635 24.690 146.825 ;
        RECT 25.895 146.635 26.065 146.825 ;
        RECT 27.740 146.655 27.910 146.845 ;
        RECT 28.195 146.655 28.365 146.875 ;
        RECT 30.320 146.845 31.265 146.875 ;
        RECT 31.470 146.845 34.945 147.755 ;
        RECT 34.955 147.555 35.905 147.755 ;
        RECT 37.235 147.555 38.165 147.755 ;
        RECT 34.955 147.075 38.165 147.555 ;
        RECT 34.955 146.875 38.020 147.075 ;
        RECT 34.955 146.845 35.890 146.875 ;
        RECT 34.630 146.825 34.800 146.845 ;
        RECT 31.425 146.680 31.585 146.790 ;
        RECT 32.335 146.635 32.505 146.825 ;
        RECT 34.630 146.655 34.810 146.825 ;
        RECT 37.850 146.655 38.020 146.875 ;
        RECT 38.235 146.845 40.005 147.755 ;
        RECT 40.015 146.845 42.765 147.655 ;
        RECT 43.245 146.845 45.975 147.755 ;
        RECT 45.995 146.845 49.665 147.655 ;
        RECT 51.045 147.525 51.965 147.755 ;
        RECT 49.675 146.845 51.965 147.525 ;
        RECT 51.985 146.930 52.415 147.715 ;
        RECT 55.950 147.525 56.860 147.745 ;
        RECT 58.395 147.525 59.745 147.755 ;
        RECT 52.435 146.845 59.745 147.525 ;
        RECT 59.795 146.845 63.465 147.655 ;
        RECT 65.765 147.525 66.685 147.755 ;
        RECT 64.395 146.845 66.685 147.525 ;
        RECT 66.695 146.845 73.805 147.755 ;
        RECT 74.150 147.525 75.070 147.755 ;
        RECT 74.150 146.845 77.615 147.525 ;
        RECT 77.745 146.930 78.175 147.715 ;
        RECT 79.155 147.525 80.505 147.755 ;
        RECT 82.040 147.525 82.950 147.745 ;
        RECT 89.990 147.525 90.900 147.745 ;
        RECT 92.435 147.525 93.785 147.755 ;
        RECT 98.270 147.525 99.180 147.745 ;
        RECT 100.715 147.525 102.065 147.755 ;
        RECT 79.155 146.845 86.465 147.525 ;
        RECT 86.475 146.845 93.785 147.525 ;
        RECT 94.755 146.845 102.065 147.525 ;
        RECT 102.115 146.845 103.485 147.655 ;
        RECT 103.505 146.930 103.935 147.715 ;
        RECT 104.050 147.525 104.970 147.755 ;
        RECT 107.730 147.525 108.650 147.755 ;
        RECT 104.050 146.845 107.515 147.525 ;
        RECT 107.730 146.845 111.195 147.525 ;
        RECT 111.510 146.845 114.985 147.755 ;
        RECT 115.305 147.525 116.235 147.755 ;
        RECT 115.305 146.845 117.140 147.525 ;
        RECT 117.295 146.845 122.805 147.655 ;
        RECT 122.815 146.845 128.325 147.655 ;
        RECT 129.265 146.930 129.695 147.715 ;
        RECT 133.230 147.525 134.140 147.745 ;
        RECT 135.675 147.525 137.025 147.755 ;
        RECT 129.715 146.845 137.025 147.525 ;
        RECT 137.535 146.845 138.905 147.655 ;
        RECT 39.690 146.825 39.860 146.845 ;
        RECT 34.640 146.635 34.810 146.655 ;
        RECT 38.315 146.635 38.485 146.825 ;
        RECT 38.770 146.685 38.890 146.795 ;
        RECT 39.690 146.655 39.865 146.825 ;
        RECT 40.155 146.655 40.325 146.845 ;
        RECT 39.695 146.635 39.865 146.655 ;
        RECT 41.995 146.635 42.165 146.825 ;
        RECT 42.910 146.685 43.030 146.795 ;
        RECT 43.380 146.635 43.550 146.825 ;
        RECT 45.675 146.655 45.845 146.845 ;
        RECT 46.135 146.655 46.305 146.845 ;
        RECT 49.350 146.635 49.520 146.825 ;
        RECT 49.815 146.655 49.985 146.845 ;
        RECT 50.740 146.635 50.910 146.825 ;
        RECT 52.575 146.655 52.745 146.845 ;
        RECT 54.410 146.635 54.580 146.825 ;
        RECT 54.875 146.635 55.045 146.825 ;
        RECT 57.180 146.635 57.350 146.825 ;
        RECT 58.555 146.635 58.725 146.825 ;
        RECT 59.935 146.655 60.105 146.845 ;
        RECT 63.625 146.690 63.785 146.800 ;
        RECT 64.085 146.680 64.245 146.790 ;
        RECT 64.535 146.655 64.705 146.845 ;
        RECT 65.455 146.635 65.625 146.825 ;
        RECT 13.335 145.825 14.705 146.635 ;
        RECT 15.635 145.955 22.945 146.635 ;
        RECT 19.150 145.735 20.060 145.955 ;
        RECT 21.595 145.725 22.945 145.955 ;
        RECT 22.995 145.725 24.345 146.635 ;
        RECT 24.375 145.725 25.725 146.635 ;
        RECT 25.755 145.825 31.265 146.635 ;
        RECT 32.205 145.725 33.555 146.635 ;
        RECT 33.575 145.725 34.925 146.635 ;
        RECT 34.955 145.725 38.625 146.635 ;
        RECT 39.105 145.765 39.535 146.550 ;
        RECT 39.555 145.955 41.845 146.635 ;
        RECT 40.925 145.725 41.845 145.955 ;
        RECT 41.855 145.825 43.225 146.635 ;
        RECT 43.235 145.725 47.625 146.635 ;
        RECT 47.835 145.725 49.665 146.635 ;
        RECT 49.675 145.725 51.025 146.635 ;
        RECT 51.250 145.725 54.725 146.635 ;
        RECT 54.735 145.955 57.025 146.635 ;
        RECT 56.105 145.725 57.025 145.955 ;
        RECT 57.035 145.725 58.385 146.635 ;
        RECT 58.415 145.825 63.925 146.635 ;
        RECT 64.865 145.765 65.295 146.550 ;
        RECT 65.315 145.825 66.685 146.635 ;
        RECT 66.840 146.605 67.010 146.845 ;
        RECT 70.055 146.635 70.225 146.825 ;
        RECT 73.275 146.635 73.445 146.825 ;
        RECT 73.730 146.685 73.850 146.795 ;
        RECT 74.195 146.635 74.365 146.825 ;
        RECT 77.415 146.655 77.585 146.845 ;
        RECT 78.345 146.690 78.505 146.800 ;
        RECT 83.395 146.635 83.565 146.825 ;
        RECT 86.155 146.655 86.325 146.845 ;
        RECT 86.615 146.655 86.785 146.845 ;
        RECT 91.215 146.635 91.385 146.825 ;
        RECT 93.050 146.685 93.170 146.795 ;
        RECT 93.515 146.635 93.685 146.825 ;
        RECT 93.985 146.690 94.145 146.800 ;
        RECT 94.895 146.655 95.065 146.845 ;
        RECT 101.150 146.635 101.320 146.825 ;
        RECT 102.255 146.655 102.425 146.845 ;
        RECT 105.290 146.635 105.460 146.825 ;
        RECT 107.315 146.655 107.485 146.845 ;
        RECT 109.155 146.635 109.325 146.825 ;
        RECT 110.995 146.655 111.165 146.845 ;
        RECT 114.670 146.655 114.840 146.845 ;
        RECT 116.975 146.825 117.140 146.845 ;
        RECT 116.975 146.635 117.145 146.825 ;
        RECT 117.435 146.655 117.605 146.845 ;
        RECT 122.955 146.655 123.125 146.845 ;
        RECT 124.335 146.635 124.505 146.825 ;
        RECT 128.485 146.690 128.645 146.800 ;
        RECT 129.390 146.635 129.560 146.825 ;
        RECT 129.855 146.655 130.025 146.845 ;
        RECT 129.860 146.635 130.025 146.655 ;
        RECT 132.155 146.635 132.325 146.825 ;
        RECT 133.995 146.635 134.165 146.825 ;
        RECT 135.835 146.635 136.005 146.825 ;
        RECT 137.210 146.685 137.330 146.795 ;
        RECT 138.595 146.635 138.765 146.845 ;
        RECT 68.970 146.605 69.905 146.635 ;
        RECT 66.840 146.405 69.905 146.605 ;
        RECT 66.695 145.925 69.905 146.405 ;
        RECT 69.915 145.955 72.205 146.635 ;
        RECT 66.695 145.725 67.625 145.925 ;
        RECT 68.955 145.725 69.905 145.925 ;
        RECT 71.285 145.725 72.205 145.955 ;
        RECT 72.225 145.725 73.575 146.635 ;
        RECT 74.055 145.955 83.160 146.635 ;
        RECT 83.255 145.955 90.565 146.635 ;
        RECT 86.770 145.735 87.680 145.955 ;
        RECT 89.215 145.725 90.565 145.955 ;
        RECT 90.625 145.765 91.055 146.550 ;
        RECT 91.075 145.825 92.905 146.635 ;
        RECT 93.375 145.955 100.685 146.635 ;
        RECT 96.890 145.735 97.800 145.955 ;
        RECT 99.335 145.725 100.685 145.955 ;
        RECT 100.735 145.955 104.635 146.635 ;
        RECT 104.875 145.955 108.775 146.635 ;
        RECT 109.015 145.955 116.325 146.635 ;
        RECT 100.735 145.725 101.665 145.955 ;
        RECT 104.875 145.725 105.805 145.955 ;
        RECT 112.530 145.735 113.440 145.955 ;
        RECT 114.975 145.725 116.325 145.955 ;
        RECT 116.385 145.765 116.815 146.550 ;
        RECT 116.835 145.955 124.145 146.635 ;
        RECT 120.350 145.735 121.260 145.955 ;
        RECT 122.795 145.725 124.145 145.955 ;
        RECT 124.195 145.825 126.025 146.635 ;
        RECT 126.230 145.725 129.705 146.635 ;
        RECT 129.860 145.955 131.695 146.635 ;
        RECT 130.765 145.725 131.695 145.955 ;
        RECT 132.015 145.825 133.845 146.635 ;
        RECT 133.855 145.955 135.685 146.635 ;
        RECT 135.695 145.955 137.525 146.635 ;
        RECT 134.340 145.725 135.685 145.955 ;
        RECT 136.180 145.725 137.525 145.955 ;
        RECT 137.535 145.825 138.905 146.635 ;
      LAYER nwell ;
        RECT 13.140 142.605 139.100 145.435 ;
      LAYER pwell ;
        RECT 13.335 141.405 14.705 142.215 ;
        RECT 14.715 141.405 18.385 142.215 ;
        RECT 18.395 142.085 19.315 142.315 ;
        RECT 18.395 141.405 20.685 142.085 ;
        RECT 20.695 141.405 26.205 142.215 ;
        RECT 26.225 141.490 26.655 142.275 ;
        RECT 26.675 141.405 32.185 142.215 ;
        RECT 32.195 141.405 33.565 142.215 ;
        RECT 33.585 141.405 37.245 142.315 ;
        RECT 38.395 142.225 39.345 142.315 ;
        RECT 37.415 141.405 39.345 142.225 ;
        RECT 39.555 141.405 42.305 142.215 ;
        RECT 42.315 142.115 43.260 142.315 ;
        RECT 42.315 141.435 45.065 142.115 ;
        RECT 45.075 142.085 46.005 142.315 ;
        RECT 42.315 141.405 43.260 141.435 ;
        RECT 13.475 141.195 13.645 141.405 ;
        RECT 14.855 141.195 15.025 141.405 ;
        RECT 20.375 141.195 20.545 141.405 ;
        RECT 20.835 141.215 21.005 141.405 ;
        RECT 23.130 141.195 23.300 141.385 ;
        RECT 23.595 141.195 23.765 141.385 ;
        RECT 26.815 141.215 26.985 141.405 ;
        RECT 29.115 141.195 29.285 141.385 ;
        RECT 32.335 141.215 32.505 141.405 ;
        RECT 32.790 141.245 32.910 141.355 ;
        RECT 33.710 141.215 33.880 141.405 ;
        RECT 37.415 141.385 37.565 141.405 ;
        RECT 34.630 141.195 34.800 141.385 ;
        RECT 36.475 141.195 36.645 141.385 ;
        RECT 36.935 141.195 37.105 141.385 ;
        RECT 37.395 141.215 37.565 141.385 ;
        RECT 38.770 141.245 38.890 141.355 ;
        RECT 39.695 141.195 39.865 141.405 ;
        RECT 44.750 141.215 44.920 141.435 ;
        RECT 45.075 141.405 48.745 142.085 ;
        RECT 48.755 141.405 51.965 142.315 ;
        RECT 51.985 141.490 52.415 142.275 ;
        RECT 52.435 141.405 54.250 142.315 ;
        RECT 68.275 142.225 69.225 142.315 ;
        RECT 54.275 141.405 59.785 142.215 ;
        RECT 59.795 141.405 65.305 142.215 ;
        RECT 65.315 141.405 68.065 142.215 ;
        RECT 68.275 141.405 70.205 142.225 ;
        RECT 70.375 141.405 73.125 142.215 ;
        RECT 76.795 142.085 77.725 142.315 ;
        RECT 73.825 141.405 77.725 142.085 ;
        RECT 77.745 141.490 78.175 142.275 ;
        RECT 78.195 141.405 81.865 142.215 ;
        RECT 85.075 142.085 86.005 142.315 ;
        RECT 82.105 141.405 86.005 142.085 ;
        RECT 86.110 142.085 87.030 142.315 ;
        RECT 86.110 141.405 89.575 142.085 ;
        RECT 89.695 141.405 93.365 142.215 ;
        RECT 96.890 142.085 97.800 142.305 ;
        RECT 99.335 142.085 100.685 142.315 ;
        RECT 93.375 141.405 100.685 142.085 ;
        RECT 100.735 141.405 103.485 142.215 ;
        RECT 103.505 141.490 103.935 142.275 ;
        RECT 104.050 142.085 104.970 142.315 ;
        RECT 104.050 141.405 107.515 142.085 ;
        RECT 108.555 141.405 112.030 142.315 ;
        RECT 115.750 142.085 116.660 142.305 ;
        RECT 118.195 142.085 119.545 142.315 ;
        RECT 120.645 142.085 121.575 142.315 ;
        RECT 112.235 141.405 119.545 142.085 ;
        RECT 119.740 141.405 121.575 142.085 ;
        RECT 121.895 141.405 123.265 142.215 ;
        RECT 124.325 142.085 125.255 142.315 ;
        RECT 123.420 141.405 125.255 142.085 ;
        RECT 125.770 141.405 129.245 142.315 ;
        RECT 129.265 141.490 129.695 142.275 ;
        RECT 133.230 142.085 134.140 142.305 ;
        RECT 135.675 142.085 137.025 142.315 ;
        RECT 129.715 141.405 137.025 142.085 ;
        RECT 137.535 141.405 138.905 142.215 ;
        RECT 45.225 141.240 45.385 141.350 ;
        RECT 46.135 141.215 46.305 141.385 ;
        RECT 48.435 141.215 48.605 141.405 ;
        RECT 48.895 141.215 49.065 141.405 ;
        RECT 50.275 141.215 50.445 141.385 ;
        RECT 50.745 141.240 50.905 141.350 ;
        RECT 46.140 141.195 46.305 141.215 ;
        RECT 50.275 141.195 50.440 141.215 ;
        RECT 51.655 141.195 51.825 141.385 ;
        RECT 53.955 141.215 54.125 141.405 ;
        RECT 54.415 141.215 54.585 141.405 ;
        RECT 59.935 141.215 60.105 141.405 ;
        RECT 60.855 141.195 61.025 141.385 ;
        RECT 61.315 141.195 61.485 141.385 ;
        RECT 65.455 141.215 65.625 141.405 ;
        RECT 70.055 141.385 70.205 141.405 ;
        RECT 66.375 141.195 66.545 141.385 ;
        RECT 70.055 141.215 70.225 141.385 ;
        RECT 70.515 141.215 70.685 141.405 ;
        RECT 73.270 141.245 73.390 141.355 ;
        RECT 73.735 141.195 73.905 141.385 ;
        RECT 77.140 141.215 77.310 141.405 ;
        RECT 78.335 141.215 78.505 141.405 ;
        RECT 79.255 141.195 79.425 141.385 ;
        RECT 84.775 141.195 84.945 141.385 ;
        RECT 85.420 141.215 85.590 141.405 ;
        RECT 89.375 141.215 89.545 141.405 ;
        RECT 89.835 141.215 90.005 141.405 ;
        RECT 90.290 141.245 90.410 141.355 ;
        RECT 91.215 141.195 91.385 141.385 ;
        RECT 93.515 141.215 93.685 141.405 ;
        RECT 96.730 141.245 96.850 141.355 ;
        RECT 97.470 141.195 97.640 141.385 ;
        RECT 100.875 141.215 101.045 141.405 ;
        RECT 101.335 141.195 101.505 141.385 ;
        RECT 105.010 141.245 105.130 141.355 ;
        RECT 105.465 141.195 105.635 141.385 ;
        RECT 107.315 141.215 107.485 141.405 ;
        RECT 108.700 141.385 108.870 141.405 ;
        RECT 107.785 141.250 107.945 141.360 ;
        RECT 108.695 141.215 108.870 141.385 ;
        RECT 112.375 141.215 112.545 141.405 ;
        RECT 119.740 141.385 119.905 141.405 ;
        RECT 108.695 141.195 108.865 141.215 ;
        RECT 113.750 141.195 113.920 141.385 ;
        RECT 116.055 141.215 116.225 141.385 ;
        RECT 116.055 141.195 116.220 141.215 ;
        RECT 116.975 141.195 117.145 141.385 ;
        RECT 119.735 141.215 119.905 141.385 ;
        RECT 122.035 141.215 122.205 141.405 ;
        RECT 123.420 141.385 123.585 141.405 ;
        RECT 122.495 141.195 122.665 141.385 ;
        RECT 123.415 141.215 123.585 141.385 ;
        RECT 124.330 141.245 124.450 141.355 ;
        RECT 127.555 141.195 127.725 141.385 ;
        RECT 128.015 141.195 128.185 141.385 ;
        RECT 128.930 141.215 129.100 141.405 ;
        RECT 129.855 141.215 130.025 141.405 ;
        RECT 135.370 141.245 135.490 141.355 ;
        RECT 135.835 141.195 136.005 141.385 ;
        RECT 137.210 141.245 137.330 141.355 ;
        RECT 138.595 141.195 138.765 141.405 ;
        RECT 13.335 140.385 14.705 141.195 ;
        RECT 14.715 140.385 20.225 141.195 ;
        RECT 20.235 140.385 22.065 141.195 ;
        RECT 22.095 140.285 23.445 141.195 ;
        RECT 23.455 140.385 28.965 141.195 ;
        RECT 28.975 140.385 32.645 141.195 ;
        RECT 33.115 140.285 34.945 141.195 ;
        RECT 34.955 140.285 36.770 141.195 ;
        RECT 36.795 140.385 38.625 141.195 ;
        RECT 39.105 140.325 39.535 141.110 ;
        RECT 39.555 140.385 45.065 141.195 ;
        RECT 46.140 140.515 47.975 141.195 ;
        RECT 47.045 140.285 47.975 140.515 ;
        RECT 48.605 140.515 50.440 141.195 ;
        RECT 51.515 140.515 53.805 141.195 ;
        RECT 48.605 140.285 49.535 140.515 ;
        RECT 52.885 140.285 53.805 140.515 ;
        RECT 53.855 140.515 61.165 141.195 ;
        RECT 53.855 140.285 55.205 140.515 ;
        RECT 56.740 140.295 57.650 140.515 ;
        RECT 61.175 140.385 64.845 141.195 ;
        RECT 64.865 140.325 65.295 141.110 ;
        RECT 66.235 140.515 73.545 141.195 ;
        RECT 69.750 140.295 70.660 140.515 ;
        RECT 72.195 140.285 73.545 140.515 ;
        RECT 73.595 140.385 79.105 141.195 ;
        RECT 79.115 140.385 84.625 141.195 ;
        RECT 84.635 140.385 90.145 141.195 ;
        RECT 90.625 140.325 91.055 141.110 ;
        RECT 91.075 140.385 96.585 141.195 ;
        RECT 97.055 140.515 100.955 141.195 ;
        RECT 97.055 140.285 97.985 140.515 ;
        RECT 101.195 140.385 104.865 141.195 ;
        RECT 105.335 140.285 108.545 141.195 ;
        RECT 108.555 140.385 110.385 141.195 ;
        RECT 110.590 140.285 114.065 141.195 ;
        RECT 114.385 140.515 116.220 141.195 ;
        RECT 114.385 140.285 115.315 140.515 ;
        RECT 116.385 140.325 116.815 141.110 ;
        RECT 116.835 140.385 122.345 141.195 ;
        RECT 122.355 140.385 124.185 141.195 ;
        RECT 124.655 140.285 127.865 141.195 ;
        RECT 127.875 140.515 135.185 141.195 ;
        RECT 135.695 140.515 137.525 141.195 ;
        RECT 131.390 140.295 132.300 140.515 ;
        RECT 133.835 140.285 135.185 140.515 ;
        RECT 136.180 140.285 137.525 140.515 ;
        RECT 137.535 140.385 138.905 141.195 ;
      LAYER nwell ;
        RECT 13.140 137.165 139.100 139.995 ;
      LAYER pwell ;
        RECT 13.335 135.965 14.705 136.775 ;
        RECT 14.715 135.965 18.385 136.775 ;
        RECT 18.395 136.645 19.530 136.875 ;
        RECT 21.925 136.645 22.855 136.875 ;
        RECT 23.915 136.645 24.835 136.875 ;
        RECT 18.395 135.965 21.605 136.645 ;
        RECT 21.925 135.965 23.760 136.645 ;
        RECT 23.915 135.965 26.205 136.645 ;
        RECT 26.225 136.050 26.655 136.835 ;
        RECT 26.675 135.965 28.025 136.875 ;
        RECT 28.055 135.965 33.565 136.775 ;
        RECT 33.590 135.965 35.405 136.875 ;
        RECT 35.415 135.965 40.925 136.775 ;
        RECT 40.935 135.965 46.445 136.775 ;
        RECT 46.455 135.965 49.205 136.775 ;
        RECT 49.215 135.965 50.565 136.875 ;
        RECT 50.595 135.965 51.945 136.875 ;
        RECT 51.985 136.050 52.415 136.835 ;
        RECT 52.435 135.965 55.605 136.875 ;
        RECT 55.655 135.965 61.165 136.775 ;
        RECT 61.175 135.965 63.925 136.775 ;
        RECT 67.910 136.645 68.820 136.865 ;
        RECT 70.355 136.645 72.125 136.875 ;
        RECT 64.395 135.965 72.125 136.645 ;
        RECT 72.215 136.645 73.145 136.875 ;
        RECT 72.215 135.965 76.115 136.645 ;
        RECT 76.355 135.965 77.725 136.775 ;
        RECT 77.745 136.050 78.175 136.835 ;
        RECT 81.710 136.645 82.620 136.865 ;
        RECT 84.155 136.645 85.925 136.875 ;
        RECT 78.195 135.965 85.925 136.645 ;
        RECT 86.015 136.645 86.945 136.875 ;
        RECT 86.015 135.965 89.915 136.645 ;
        RECT 90.155 135.965 93.825 136.775 ;
        RECT 94.295 136.645 95.225 136.875 ;
        RECT 98.530 136.645 99.450 136.875 ;
        RECT 94.295 135.965 98.195 136.645 ;
        RECT 98.530 135.965 101.995 136.645 ;
        RECT 102.115 135.965 103.485 136.775 ;
        RECT 103.505 136.050 103.935 136.835 ;
        RECT 103.955 135.965 106.705 136.775 ;
        RECT 107.175 135.965 110.385 136.875 ;
        RECT 110.395 135.965 113.605 136.875 ;
        RECT 113.925 136.645 114.855 136.875 ;
        RECT 113.925 135.965 115.760 136.645 ;
        RECT 115.915 135.965 117.745 136.775 ;
        RECT 117.755 135.965 120.965 136.875 ;
        RECT 120.975 135.965 126.485 136.775 ;
        RECT 128.005 136.645 128.935 136.875 ;
        RECT 127.100 135.965 128.935 136.645 ;
        RECT 129.265 136.050 129.695 136.835 ;
        RECT 129.910 135.965 133.385 136.875 ;
        RECT 133.395 135.965 136.605 136.875 ;
        RECT 137.535 135.965 138.905 136.775 ;
        RECT 13.475 135.755 13.645 135.965 ;
        RECT 14.855 135.945 15.025 135.965 ;
        RECT 14.850 135.775 15.025 135.945 ;
        RECT 14.850 135.755 15.020 135.775 ;
        RECT 16.235 135.755 16.405 135.945 ;
        RECT 21.295 135.775 21.465 135.965 ;
        RECT 23.595 135.945 23.760 135.965 ;
        RECT 23.595 135.775 23.765 135.945 ;
        RECT 25.435 135.755 25.605 135.945 ;
        RECT 25.895 135.755 26.065 135.965 ;
        RECT 26.820 135.775 26.990 135.965 ;
        RECT 28.195 135.775 28.365 135.965 ;
        RECT 30.495 135.755 30.665 135.945 ;
        RECT 33.255 135.755 33.425 135.945 ;
        RECT 33.715 135.775 33.885 135.965 ;
        RECT 35.555 135.775 35.725 135.965 ;
        RECT 36.475 135.755 36.645 135.945 ;
        RECT 36.935 135.755 37.105 135.945 ;
        RECT 38.770 135.805 38.890 135.915 ;
        RECT 39.695 135.755 39.865 135.945 ;
        RECT 41.075 135.775 41.245 135.965 ;
        RECT 45.225 135.800 45.385 135.910 ;
        RECT 46.135 135.755 46.305 135.945 ;
        RECT 46.595 135.775 46.765 135.965 ;
        RECT 49.360 135.775 49.530 135.965 ;
        RECT 50.740 135.775 50.910 135.965 ;
        RECT 55.335 135.775 55.505 135.965 ;
        RECT 55.795 135.775 55.965 135.965 ;
        RECT 56.255 135.755 56.425 135.945 ;
        RECT 56.715 135.755 56.885 135.945 ;
        RECT 61.315 135.775 61.485 135.965 ;
        RECT 62.235 135.755 62.405 135.945 ;
        RECT 64.070 135.805 64.190 135.915 ;
        RECT 64.535 135.775 64.705 135.965 ;
        RECT 65.455 135.755 65.625 135.945 ;
        RECT 72.630 135.775 72.800 135.965 ;
        RECT 72.820 135.755 72.990 135.945 ;
        RECT 13.335 134.945 14.705 135.755 ;
        RECT 14.735 134.845 16.085 135.755 ;
        RECT 16.095 135.075 23.405 135.755 ;
        RECT 19.610 134.855 20.520 135.075 ;
        RECT 22.055 134.845 23.405 135.075 ;
        RECT 23.455 135.075 25.745 135.755 ;
        RECT 25.755 135.075 28.965 135.755 ;
        RECT 23.455 134.845 24.375 135.075 ;
        RECT 27.830 134.845 28.965 135.075 ;
        RECT 28.975 134.845 30.790 135.755 ;
        RECT 30.815 134.845 33.565 135.755 ;
        RECT 33.575 134.845 36.785 135.755 ;
        RECT 36.795 134.945 38.625 135.755 ;
        RECT 39.105 134.885 39.535 135.670 ;
        RECT 39.555 134.945 45.065 135.755 ;
        RECT 45.995 135.075 49.205 135.755 ;
        RECT 48.070 134.845 49.205 135.075 ;
        RECT 49.255 135.075 56.565 135.755 ;
        RECT 49.255 134.845 50.605 135.075 ;
        RECT 52.140 134.855 53.050 135.075 ;
        RECT 56.575 134.945 62.085 135.755 ;
        RECT 62.095 134.945 64.845 135.755 ;
        RECT 64.865 134.885 65.295 135.670 ;
        RECT 65.315 135.075 72.625 135.755 ;
        RECT 68.830 134.855 69.740 135.075 ;
        RECT 71.275 134.845 72.625 135.075 ;
        RECT 72.675 134.845 74.025 135.755 ;
        RECT 74.200 135.725 74.370 135.945 ;
        RECT 76.495 135.775 76.665 135.965 ;
        RECT 78.335 135.775 78.505 135.965 ;
        RECT 80.820 135.755 80.990 135.945 ;
        RECT 81.555 135.755 81.725 135.945 ;
        RECT 86.430 135.775 86.600 135.965 ;
        RECT 89.375 135.755 89.545 135.945 ;
        RECT 90.295 135.775 90.465 135.965 ;
        RECT 91.215 135.755 91.385 135.945 ;
        RECT 93.055 135.755 93.225 135.945 ;
        RECT 93.970 135.805 94.090 135.915 ;
        RECT 94.710 135.775 94.880 135.965 ;
        RECT 100.690 135.755 100.860 135.945 ;
        RECT 101.795 135.775 101.965 135.965 ;
        RECT 102.255 135.775 102.425 135.965 ;
        RECT 104.095 135.775 104.265 135.965 ;
        RECT 104.555 135.755 104.725 135.945 ;
        RECT 105.935 135.755 106.105 135.945 ;
        RECT 106.850 135.805 106.970 135.915 ;
        RECT 107.305 135.775 107.475 135.965 ;
        RECT 110.525 135.775 110.695 135.965 ;
        RECT 115.595 135.945 115.760 135.965 ;
        RECT 113.295 135.755 113.465 135.945 ;
        RECT 115.595 135.775 115.765 135.945 ;
        RECT 116.055 135.915 116.225 135.965 ;
        RECT 116.050 135.805 116.225 135.915 ;
        RECT 116.055 135.775 116.225 135.805 ;
        RECT 116.975 135.755 117.145 135.945 ;
        RECT 120.655 135.775 120.825 135.965 ;
        RECT 121.115 135.775 121.285 135.965 ;
        RECT 127.100 135.945 127.265 135.965 ;
        RECT 124.335 135.755 124.505 135.945 ;
        RECT 126.630 135.805 126.750 135.915 ;
        RECT 127.095 135.755 127.265 135.945 ;
        RECT 133.070 135.775 133.240 135.965 ;
        RECT 134.455 135.755 134.625 135.945 ;
        RECT 135.835 135.755 136.005 135.945 ;
        RECT 136.295 135.775 136.465 135.965 ;
        RECT 136.765 135.810 136.925 135.920 ;
        RECT 138.595 135.755 138.765 135.965 ;
        RECT 76.330 135.725 77.265 135.755 ;
        RECT 74.200 135.525 77.265 135.725 ;
        RECT 74.055 135.045 77.265 135.525 ;
        RECT 77.505 135.075 81.405 135.755 ;
        RECT 81.415 135.075 89.145 135.755 ;
        RECT 74.055 134.845 74.985 135.045 ;
        RECT 76.315 134.845 77.265 135.045 ;
        RECT 80.475 134.845 81.405 135.075 ;
        RECT 84.930 134.855 85.840 135.075 ;
        RECT 87.375 134.845 89.145 135.075 ;
        RECT 89.235 134.945 90.605 135.755 ;
        RECT 90.625 134.885 91.055 135.670 ;
        RECT 91.075 134.945 92.905 135.755 ;
        RECT 92.915 135.075 100.225 135.755 ;
        RECT 96.430 134.855 97.340 135.075 ;
        RECT 98.875 134.845 100.225 135.075 ;
        RECT 100.275 135.075 104.175 135.755 ;
        RECT 100.275 134.845 101.205 135.075 ;
        RECT 104.415 134.945 105.785 135.755 ;
        RECT 105.795 135.075 113.105 135.755 ;
        RECT 113.155 135.075 115.895 135.755 ;
        RECT 109.310 134.855 110.220 135.075 ;
        RECT 111.755 134.845 113.105 135.075 ;
        RECT 116.385 134.885 116.815 135.670 ;
        RECT 116.835 135.075 124.145 135.755 ;
        RECT 120.350 134.855 121.260 135.075 ;
        RECT 122.795 134.845 124.145 135.075 ;
        RECT 124.195 134.945 126.945 135.755 ;
        RECT 126.955 135.075 134.265 135.755 ;
        RECT 130.470 134.855 131.380 135.075 ;
        RECT 132.915 134.845 134.265 135.075 ;
        RECT 134.315 134.945 135.685 135.755 ;
        RECT 135.695 135.075 137.525 135.755 ;
        RECT 136.180 134.845 137.525 135.075 ;
        RECT 137.535 134.945 138.905 135.755 ;
      LAYER nwell ;
        RECT 13.140 131.725 139.100 134.555 ;
      LAYER pwell ;
        RECT 13.335 130.525 14.705 131.335 ;
        RECT 14.715 130.525 17.465 131.335 ;
        RECT 21.450 131.205 22.360 131.425 ;
        RECT 23.895 131.205 25.245 131.435 ;
        RECT 17.935 130.525 25.245 131.205 ;
        RECT 26.225 130.610 26.655 131.395 ;
        RECT 28.045 131.205 28.965 131.435 ;
        RECT 26.675 130.525 28.965 131.205 ;
        RECT 28.975 130.525 30.325 131.435 ;
        RECT 31.315 130.525 34.485 131.435 ;
        RECT 38.010 131.205 38.920 131.425 ;
        RECT 40.455 131.205 41.805 131.435 ;
        RECT 34.495 130.525 41.805 131.205 ;
        RECT 41.855 130.525 43.670 131.435 ;
        RECT 45.065 131.205 45.985 131.435 ;
        RECT 47.365 131.205 48.285 131.435 ;
        RECT 43.695 130.525 45.985 131.205 ;
        RECT 45.995 130.525 48.285 131.205 ;
        RECT 48.295 130.525 49.645 131.435 ;
        RECT 51.045 131.205 51.965 131.435 ;
        RECT 49.675 130.525 51.965 131.205 ;
        RECT 51.985 130.610 52.415 131.395 ;
        RECT 52.435 130.525 57.945 131.335 ;
        RECT 57.955 130.525 63.465 131.335 ;
        RECT 63.475 130.525 67.145 131.335 ;
        RECT 67.925 131.205 68.855 131.435 ;
        RECT 70.965 131.205 71.895 131.435 ;
        RECT 67.925 130.525 69.760 131.205 ;
        RECT 13.475 130.315 13.645 130.525 ;
        RECT 14.855 130.315 15.025 130.525 ;
        RECT 17.610 130.365 17.730 130.475 ;
        RECT 18.075 130.335 18.245 130.525 ;
        RECT 20.375 130.315 20.545 130.505 ;
        RECT 25.445 130.370 25.605 130.480 ;
        RECT 26.815 130.335 26.985 130.525 ;
        RECT 29.120 130.505 29.290 130.525 ;
        RECT 29.115 130.335 29.290 130.505 ;
        RECT 29.115 130.315 29.285 130.335 ;
        RECT 29.575 130.315 29.745 130.505 ;
        RECT 30.505 130.370 30.665 130.480 ;
        RECT 31.415 130.335 31.585 130.525 ;
        RECT 34.635 130.335 34.805 130.525 ;
        RECT 36.935 130.315 37.105 130.505 ;
        RECT 37.395 130.315 37.565 130.505 ;
        RECT 39.695 130.315 39.865 130.505 ;
        RECT 41.075 130.315 41.245 130.505 ;
        RECT 43.375 130.335 43.545 130.525 ;
        RECT 43.835 130.335 44.005 130.525 ;
        RECT 44.295 130.315 44.465 130.505 ;
        RECT 46.135 130.335 46.305 130.525 ;
        RECT 48.440 130.335 48.610 130.525 ;
        RECT 49.815 130.335 49.985 130.525 ;
        RECT 52.575 130.315 52.745 130.525 ;
        RECT 53.035 130.315 53.205 130.505 ;
        RECT 58.095 130.335 58.265 130.525 ;
        RECT 58.550 130.365 58.670 130.475 ;
        RECT 59.015 130.315 59.185 130.505 ;
        RECT 63.615 130.335 63.785 130.525 ;
        RECT 69.595 130.505 69.760 130.525 ;
        RECT 70.060 130.525 71.895 131.205 ;
        RECT 72.415 131.345 73.365 131.435 ;
        RECT 72.415 130.525 74.345 131.345 ;
        RECT 74.515 130.525 77.265 131.335 ;
        RECT 77.745 130.610 78.175 131.395 ;
        RECT 78.655 131.235 79.585 131.435 ;
        RECT 80.920 131.235 81.865 131.435 ;
        RECT 78.655 130.755 81.865 131.235 ;
        RECT 83.245 131.205 84.165 131.435 ;
        RECT 87.690 131.205 88.600 131.425 ;
        RECT 90.135 131.205 91.905 131.435 ;
        RECT 78.795 130.555 81.865 130.755 ;
        RECT 70.060 130.505 70.225 130.525 ;
        RECT 74.195 130.505 74.345 130.525 ;
        RECT 64.085 130.360 64.245 130.470 ;
        RECT 66.370 130.315 66.540 130.505 ;
        RECT 66.835 130.315 67.005 130.505 ;
        RECT 67.290 130.365 67.410 130.475 ;
        RECT 69.140 130.315 69.310 130.505 ;
        RECT 69.595 130.475 69.765 130.505 ;
        RECT 69.590 130.365 69.765 130.475 ;
        RECT 69.595 130.335 69.765 130.365 ;
        RECT 70.050 130.335 70.225 130.505 ;
        RECT 70.050 130.315 70.220 130.335 ;
        RECT 71.435 130.315 71.605 130.505 ;
        RECT 74.195 130.335 74.365 130.505 ;
        RECT 74.655 130.335 74.825 130.525 ;
        RECT 76.955 130.315 77.125 130.505 ;
        RECT 78.795 130.475 78.965 130.555 ;
        RECT 80.920 130.525 81.865 130.555 ;
        RECT 81.875 130.525 84.165 131.205 ;
        RECT 84.175 130.525 91.905 131.205 ;
        RECT 91.995 130.525 93.825 131.335 ;
        RECT 97.810 131.205 98.720 131.425 ;
        RECT 100.255 131.205 101.605 131.435 ;
        RECT 94.295 130.525 101.605 131.205 ;
        RECT 101.655 130.525 103.485 131.335 ;
        RECT 103.505 130.610 103.935 131.395 ;
        RECT 104.050 131.205 104.970 131.435 ;
        RECT 104.050 130.525 107.515 131.205 ;
        RECT 107.635 130.525 111.110 131.435 ;
        RECT 111.315 130.525 114.525 131.435 ;
        RECT 114.535 130.525 116.365 131.335 ;
        RECT 116.375 130.525 119.850 131.435 ;
        RECT 120.365 131.205 121.295 131.435 ;
        RECT 120.365 130.525 122.200 131.205 ;
        RECT 122.355 130.525 125.105 131.335 ;
        RECT 125.770 130.525 129.245 131.435 ;
        RECT 129.265 130.610 129.695 131.395 ;
        RECT 130.025 131.205 130.955 131.435 ;
        RECT 132.325 131.205 133.255 131.435 ;
        RECT 130.025 130.525 131.860 131.205 ;
        RECT 132.325 130.525 134.160 131.205 ;
        RECT 134.315 130.525 135.685 131.335 ;
        RECT 136.180 131.205 137.525 131.435 ;
        RECT 135.695 130.525 137.525 131.205 ;
        RECT 137.535 130.525 138.905 131.335 ;
        RECT 77.410 130.365 77.530 130.475 ;
        RECT 78.330 130.365 78.450 130.475 ;
        RECT 78.790 130.365 78.965 130.475 ;
        RECT 78.795 130.335 78.965 130.365 ;
        RECT 79.255 130.315 79.425 130.505 ;
        RECT 13.335 129.505 14.705 130.315 ;
        RECT 14.715 129.505 20.225 130.315 ;
        RECT 20.235 129.505 22.065 130.315 ;
        RECT 22.115 129.635 29.425 130.315 ;
        RECT 22.115 129.405 23.465 129.635 ;
        RECT 25.000 129.415 25.910 129.635 ;
        RECT 29.435 129.505 34.945 130.315 ;
        RECT 34.955 129.635 37.245 130.315 ;
        RECT 34.955 129.405 35.875 129.635 ;
        RECT 37.255 129.505 39.085 130.315 ;
        RECT 39.105 129.445 39.535 130.230 ;
        RECT 39.555 129.505 40.925 130.315 ;
        RECT 41.035 129.405 44.145 130.315 ;
        RECT 44.155 129.505 45.525 130.315 ;
        RECT 45.575 129.635 52.885 130.315 ;
        RECT 45.575 129.405 46.925 129.635 ;
        RECT 48.460 129.415 49.370 129.635 ;
        RECT 52.895 129.505 58.405 130.315 ;
        RECT 58.875 129.635 63.690 130.315 ;
        RECT 64.865 129.445 65.295 130.230 ;
        RECT 65.335 129.405 66.685 130.315 ;
        RECT 66.695 129.505 68.065 130.315 ;
        RECT 68.075 129.405 69.425 130.315 ;
        RECT 69.935 129.405 71.285 130.315 ;
        RECT 71.295 129.505 76.805 130.315 ;
        RECT 76.815 129.505 78.645 130.315 ;
        RECT 79.125 129.405 80.475 130.315 ;
        RECT 80.635 130.285 80.805 130.505 ;
        RECT 82.015 130.335 82.185 130.525 ;
        RECT 83.865 130.360 84.025 130.470 ;
        RECT 84.315 130.335 84.485 130.525 ;
        RECT 85.050 130.315 85.220 130.505 ;
        RECT 88.915 130.315 89.085 130.505 ;
        RECT 91.215 130.315 91.385 130.505 ;
        RECT 92.135 130.335 92.305 130.525 ;
        RECT 93.970 130.365 94.090 130.475 ;
        RECT 94.435 130.335 94.605 130.525 ;
        RECT 96.745 130.360 96.905 130.470 ;
        RECT 97.930 130.315 98.100 130.505 ;
        RECT 101.795 130.315 101.965 130.525 ;
        RECT 107.315 130.315 107.485 130.525 ;
        RECT 107.780 130.335 107.950 130.525 ;
        RECT 111.445 130.335 111.615 130.525 ;
        RECT 112.840 130.315 113.010 130.505 ;
        RECT 114.675 130.335 114.845 130.525 ;
        RECT 116.520 130.335 116.690 130.525 ;
        RECT 122.035 130.505 122.200 130.525 ;
        RECT 118.815 130.335 118.985 130.505 ;
        RECT 118.815 130.315 118.980 130.335 ;
        RECT 119.275 130.315 119.445 130.505 ;
        RECT 122.035 130.335 122.205 130.505 ;
        RECT 122.495 130.335 122.665 130.525 ;
        RECT 125.250 130.365 125.370 130.475 ;
        RECT 128.010 130.315 128.180 130.505 ;
        RECT 128.475 130.315 128.645 130.505 ;
        RECT 128.930 130.335 129.100 130.525 ;
        RECT 131.695 130.505 131.860 130.525 ;
        RECT 133.995 130.505 134.160 130.525 ;
        RECT 131.695 130.335 131.865 130.505 ;
        RECT 133.995 130.335 134.165 130.505 ;
        RECT 134.455 130.335 134.625 130.525 ;
        RECT 135.835 130.315 136.005 130.525 ;
        RECT 138.595 130.315 138.765 130.525 ;
        RECT 82.760 130.285 83.705 130.315 ;
        RECT 80.635 130.085 83.705 130.285 ;
        RECT 80.495 129.605 83.705 130.085 ;
        RECT 80.495 129.405 81.425 129.605 ;
        RECT 82.760 129.405 83.705 129.605 ;
        RECT 84.635 129.635 88.535 130.315 ;
        RECT 84.635 129.405 85.565 129.635 ;
        RECT 88.775 129.505 90.605 130.315 ;
        RECT 90.625 129.445 91.055 130.230 ;
        RECT 91.075 129.505 96.585 130.315 ;
        RECT 97.515 129.635 101.415 130.315 ;
        RECT 97.515 129.405 98.445 129.635 ;
        RECT 101.655 129.505 107.165 130.315 ;
        RECT 107.175 129.505 112.685 130.315 ;
        RECT 112.695 129.405 116.170 130.315 ;
        RECT 116.385 129.445 116.815 130.230 ;
        RECT 117.145 129.635 118.980 130.315 ;
        RECT 117.145 129.405 118.075 129.635 ;
        RECT 119.135 129.505 124.645 130.315 ;
        RECT 124.850 129.405 128.325 130.315 ;
        RECT 128.335 129.635 135.645 130.315 ;
        RECT 135.695 129.635 137.525 130.315 ;
        RECT 131.850 129.415 132.760 129.635 ;
        RECT 134.295 129.405 135.645 129.635 ;
        RECT 136.180 129.405 137.525 129.635 ;
        RECT 137.535 129.505 138.905 130.315 ;
      LAYER nwell ;
        RECT 13.140 126.285 139.100 129.115 ;
      LAYER pwell ;
        RECT 13.335 125.085 14.705 125.895 ;
        RECT 14.715 125.085 20.225 125.895 ;
        RECT 20.235 125.085 22.985 125.895 ;
        RECT 24.115 125.085 26.205 125.895 ;
        RECT 26.225 125.170 26.655 125.955 ;
        RECT 26.910 125.085 31.725 125.765 ;
        RECT 31.735 125.085 37.245 125.895 ;
        RECT 37.255 125.085 42.765 125.895 ;
        RECT 42.775 125.085 48.285 125.895 ;
        RECT 48.295 125.085 51.965 125.895 ;
        RECT 51.985 125.170 52.415 125.955 ;
        RECT 52.435 125.085 56.105 125.895 ;
        RECT 56.115 125.085 57.465 125.995 ;
        RECT 57.495 125.085 58.865 125.895 ;
        RECT 58.875 125.085 69.885 125.995 ;
        RECT 69.915 125.085 71.285 125.895 ;
        RECT 71.390 125.765 72.310 125.995 ;
        RECT 74.975 125.765 75.895 125.995 ;
        RECT 71.390 125.085 74.855 125.765 ;
        RECT 74.975 125.085 77.265 125.765 ;
        RECT 77.745 125.170 78.175 125.955 ;
        RECT 79.530 125.795 80.485 125.995 ;
        RECT 78.205 125.115 80.485 125.795 ;
        RECT 80.955 125.795 81.885 125.995 ;
        RECT 83.220 125.795 84.165 125.995 ;
        RECT 80.955 125.315 84.165 125.795 ;
        RECT 13.475 124.875 13.645 125.085 ;
        RECT 14.855 124.875 15.025 125.085 ;
        RECT 20.375 124.875 20.545 125.085 ;
        RECT 23.130 124.925 23.250 125.035 ;
        RECT 25.435 124.875 25.605 125.065 ;
        RECT 25.895 124.875 26.065 125.085 ;
        RECT 27.730 124.925 27.850 125.035 ;
        RECT 28.200 124.875 28.370 125.065 ;
        RECT 31.415 124.895 31.585 125.085 ;
        RECT 31.875 124.895 32.045 125.085 ;
        RECT 37.395 124.895 37.565 125.085 ;
        RECT 39.695 124.875 39.865 125.065 ;
        RECT 42.915 124.895 43.085 125.085 ;
        RECT 45.215 124.875 45.385 125.065 ;
        RECT 48.435 124.895 48.605 125.085 ;
        RECT 50.735 124.875 50.905 125.065 ;
        RECT 52.575 124.895 52.745 125.085 ;
        RECT 53.490 124.925 53.610 125.035 ;
        RECT 53.955 124.875 54.125 125.065 ;
        RECT 56.260 124.895 56.430 125.085 ;
        RECT 57.635 124.875 57.805 125.085 ;
        RECT 59.020 124.895 59.190 125.085 ;
        RECT 65.455 124.875 65.625 125.065 ;
        RECT 70.055 124.895 70.225 125.085 ;
        RECT 72.815 124.875 72.985 125.065 ;
        RECT 74.655 124.895 74.825 125.085 ;
        RECT 76.495 124.875 76.665 125.065 ;
        RECT 76.955 124.895 77.125 125.085 ;
        RECT 77.410 124.925 77.530 125.035 ;
        RECT 78.330 124.895 78.500 125.115 ;
        RECT 79.530 125.085 80.485 125.115 ;
        RECT 81.095 125.115 84.165 125.315 ;
        RECT 78.610 124.875 78.780 125.065 ;
        RECT 80.630 124.925 80.750 125.035 ;
        RECT 81.095 124.895 81.265 125.115 ;
        RECT 83.220 125.085 84.165 125.115 ;
        RECT 84.635 125.765 85.565 125.995 ;
        RECT 84.635 125.085 88.535 125.765 ;
        RECT 88.775 125.085 94.285 125.895 ;
        RECT 94.295 125.085 95.665 125.895 ;
        RECT 99.190 125.765 100.100 125.985 ;
        RECT 101.635 125.765 102.985 125.995 ;
        RECT 95.675 125.085 102.985 125.765 ;
        RECT 103.505 125.170 103.935 125.955 ;
        RECT 103.955 125.765 104.885 125.995 ;
        RECT 108.190 125.765 109.110 125.995 ;
        RECT 115.750 125.765 116.660 125.985 ;
        RECT 118.195 125.765 119.545 125.995 ;
        RECT 103.955 125.085 107.855 125.765 ;
        RECT 108.190 125.085 111.655 125.765 ;
        RECT 112.235 125.085 119.545 125.765 ;
        RECT 119.595 125.085 125.105 125.895 ;
        RECT 125.115 125.085 128.785 125.895 ;
        RECT 129.265 125.170 129.695 125.955 ;
        RECT 129.715 125.085 132.925 125.995 ;
        RECT 134.340 125.765 135.685 125.995 ;
        RECT 136.180 125.765 137.525 125.995 ;
        RECT 133.855 125.085 135.685 125.765 ;
        RECT 135.695 125.085 137.525 125.765 ;
        RECT 137.535 125.085 138.905 125.895 ;
        RECT 82.470 124.925 82.590 125.035 ;
        RECT 82.935 124.875 83.105 125.065 ;
        RECT 84.310 124.925 84.430 125.035 ;
        RECT 85.050 124.895 85.220 125.085 ;
        RECT 88.915 124.895 89.085 125.085 ;
        RECT 91.490 124.875 91.660 125.065 ;
        RECT 94.435 124.895 94.605 125.085 ;
        RECT 95.350 124.925 95.470 125.035 ;
        RECT 95.815 124.875 95.985 125.085 ;
        RECT 103.170 124.925 103.290 125.035 ;
        RECT 104.370 124.895 104.540 125.085 ;
        RECT 106.390 124.875 106.560 125.065 ;
        RECT 106.855 124.875 107.025 125.065 ;
        RECT 111.455 124.895 111.625 125.085 ;
        RECT 111.910 124.925 112.030 125.035 ;
        RECT 112.375 124.875 112.545 125.085 ;
        RECT 116.050 124.925 116.170 125.035 ;
        RECT 116.970 124.925 117.090 125.035 ;
        RECT 117.435 124.875 117.605 125.065 ;
        RECT 119.275 124.875 119.445 125.065 ;
        RECT 119.735 124.895 119.905 125.085 ;
        RECT 122.950 124.925 123.070 125.035 ;
        RECT 125.255 124.895 125.425 125.085 ;
        RECT 126.630 124.875 126.800 125.065 ;
        RECT 127.095 124.875 127.265 125.065 ;
        RECT 128.930 124.925 129.050 125.035 ;
        RECT 132.615 124.895 132.785 125.085 ;
        RECT 133.085 124.930 133.245 125.040 ;
        RECT 133.995 124.895 134.165 125.085 ;
        RECT 134.455 124.875 134.625 125.065 ;
        RECT 135.835 124.895 136.005 125.085 ;
        RECT 137.210 124.925 137.330 125.035 ;
        RECT 138.595 124.875 138.765 125.085 ;
        RECT 13.335 124.065 14.705 124.875 ;
        RECT 14.715 124.065 20.225 124.875 ;
        RECT 20.235 124.065 22.985 124.875 ;
        RECT 23.455 124.195 25.745 124.875 ;
        RECT 23.455 123.965 24.375 124.195 ;
        RECT 25.755 124.065 27.585 124.875 ;
        RECT 28.055 123.965 39.065 124.875 ;
        RECT 39.105 124.005 39.535 124.790 ;
        RECT 39.555 124.065 45.065 124.875 ;
        RECT 45.075 124.065 50.585 124.875 ;
        RECT 50.595 124.065 53.345 124.875 ;
        RECT 53.925 124.195 57.390 124.875 ;
        RECT 57.495 124.195 64.805 124.875 ;
        RECT 56.470 123.965 57.390 124.195 ;
        RECT 61.010 123.975 61.920 124.195 ;
        RECT 63.455 123.965 64.805 124.195 ;
        RECT 64.865 124.005 65.295 124.790 ;
        RECT 65.315 124.195 72.625 124.875 ;
        RECT 72.785 124.195 76.250 124.875 ;
        RECT 68.830 123.975 69.740 124.195 ;
        RECT 71.275 123.965 72.625 124.195 ;
        RECT 75.330 123.965 76.250 124.195 ;
        RECT 76.355 124.065 78.185 124.875 ;
        RECT 78.195 124.195 82.095 124.875 ;
        RECT 82.795 124.195 90.525 124.875 ;
        RECT 78.195 123.965 79.125 124.195 ;
        RECT 86.310 123.975 87.220 124.195 ;
        RECT 88.755 123.965 90.525 124.195 ;
        RECT 90.625 124.005 91.055 124.790 ;
        RECT 91.075 124.195 94.975 124.875 ;
        RECT 95.675 124.195 102.985 124.875 ;
        RECT 91.075 123.965 92.005 124.195 ;
        RECT 99.190 123.975 100.100 124.195 ;
        RECT 101.635 123.965 102.985 124.195 ;
        RECT 103.115 123.965 106.700 124.875 ;
        RECT 106.715 124.065 112.225 124.875 ;
        RECT 112.235 124.065 115.905 124.875 ;
        RECT 116.385 124.005 116.815 124.790 ;
        RECT 117.295 124.195 119.125 124.875 ;
        RECT 117.780 123.965 119.125 124.195 ;
        RECT 119.135 124.065 122.805 124.875 ;
        RECT 123.470 123.965 126.945 124.875 ;
        RECT 126.955 124.195 134.265 124.875 ;
        RECT 130.470 123.975 131.380 124.195 ;
        RECT 132.915 123.965 134.265 124.195 ;
        RECT 134.315 124.065 137.065 124.875 ;
        RECT 137.535 124.065 138.905 124.875 ;
      LAYER nwell ;
        RECT 13.140 120.845 139.100 123.675 ;
      LAYER pwell ;
        RECT 13.335 119.645 14.705 120.455 ;
        RECT 14.715 119.645 16.085 120.455 ;
        RECT 16.135 120.325 17.485 120.555 ;
        RECT 19.020 120.325 19.930 120.545 ;
        RECT 16.135 119.645 23.445 120.325 ;
        RECT 23.465 119.645 26.195 120.555 ;
        RECT 26.225 119.730 26.655 120.515 ;
        RECT 26.675 119.645 28.045 120.455 ;
        RECT 33.115 120.325 34.250 120.555 ;
        RECT 38.155 120.325 39.085 120.555 ;
        RECT 28.055 119.645 32.870 120.325 ;
        RECT 33.115 119.645 36.325 120.325 ;
        RECT 36.335 119.645 39.085 120.325 ;
        RECT 39.095 119.645 41.845 120.555 ;
        RECT 41.855 119.875 43.690 120.555 ;
        RECT 42.000 119.645 43.690 119.875 ;
        RECT 44.155 119.645 49.665 120.455 ;
        RECT 49.675 119.645 51.505 120.455 ;
        RECT 51.985 119.730 52.415 120.515 ;
        RECT 52.435 119.645 54.250 120.555 ;
        RECT 57.790 120.325 58.700 120.545 ;
        RECT 60.235 120.325 61.585 120.555 ;
        RECT 69.435 120.325 70.365 120.555 ;
        RECT 54.275 119.645 61.585 120.325 ;
        RECT 61.635 119.645 66.450 120.325 ;
        RECT 66.695 119.645 70.365 120.325 ;
        RECT 70.470 120.325 71.390 120.555 ;
        RECT 75.395 120.355 76.775 120.555 ;
        RECT 70.470 119.645 73.935 120.325 ;
        RECT 74.070 119.675 76.775 120.355 ;
        RECT 77.745 119.730 78.175 120.515 ;
        RECT 13.475 119.435 13.645 119.645 ;
        RECT 14.855 119.435 15.025 119.645 ;
        RECT 18.535 119.455 18.705 119.625 ;
        RECT 18.535 119.435 18.700 119.455 ;
        RECT 13.335 118.625 14.705 119.435 ;
        RECT 14.715 118.625 16.545 119.435 ;
        RECT 16.865 118.755 18.700 119.435 ;
        RECT 19.000 119.405 19.170 119.625 ;
        RECT 22.215 119.435 22.385 119.625 ;
        RECT 23.135 119.455 23.305 119.645 ;
        RECT 25.895 119.455 26.065 119.645 ;
        RECT 26.815 119.455 26.985 119.645 ;
        RECT 28.195 119.455 28.365 119.645 ;
        RECT 29.575 119.455 29.745 119.625 ;
        RECT 29.580 119.435 29.745 119.455 ;
        RECT 31.875 119.435 32.045 119.625 ;
        RECT 36.015 119.455 36.185 119.645 ;
        RECT 36.475 119.455 36.645 119.645 ;
        RECT 39.235 119.455 39.405 119.645 ;
        RECT 39.695 119.435 39.865 119.625 ;
        RECT 42.000 119.455 42.170 119.645 ;
        RECT 42.455 119.455 42.625 119.625 ;
        RECT 44.295 119.455 44.465 119.645 ;
        RECT 42.475 119.435 42.625 119.455 ;
        RECT 44.755 119.435 44.925 119.625 ;
        RECT 46.590 119.485 46.710 119.595 ;
        RECT 48.435 119.435 48.605 119.625 ;
        RECT 48.895 119.435 49.065 119.625 ;
        RECT 49.815 119.455 49.985 119.645 ;
        RECT 51.650 119.485 51.770 119.595 ;
        RECT 53.955 119.455 54.125 119.645 ;
        RECT 54.415 119.455 54.585 119.645 ;
        RECT 56.255 119.435 56.425 119.625 ;
        RECT 61.315 119.435 61.485 119.625 ;
        RECT 61.775 119.455 61.945 119.645 ;
        RECT 65.455 119.435 65.625 119.625 ;
        RECT 66.835 119.455 67.005 119.645 ;
        RECT 73.735 119.455 73.905 119.645 ;
        RECT 74.195 119.455 74.365 119.675 ;
        RECT 75.395 119.645 76.775 119.675 ;
        RECT 78.195 119.645 79.545 120.555 ;
        RECT 79.575 119.645 83.245 120.455 ;
        RECT 87.230 120.325 88.140 120.545 ;
        RECT 89.675 120.325 91.445 120.555 ;
        RECT 83.715 119.645 91.445 120.325 ;
        RECT 91.535 119.645 97.045 120.455 ;
        RECT 97.055 119.645 100.725 120.455 ;
        RECT 101.665 119.645 103.015 120.555 ;
        RECT 103.505 119.730 103.935 120.515 ;
        RECT 105.295 120.355 106.705 120.555 ;
        RECT 103.970 119.675 106.705 120.355 ;
        RECT 74.655 119.455 74.825 119.625 ;
        RECT 74.655 119.435 74.820 119.455 ;
        RECT 75.120 119.435 75.290 119.625 ;
        RECT 76.955 119.435 77.125 119.625 ;
        RECT 79.260 119.455 79.430 119.645 ;
        RECT 79.715 119.455 79.885 119.645 ;
        RECT 83.390 119.485 83.510 119.595 ;
        RECT 83.855 119.455 84.025 119.645 ;
        RECT 84.775 119.435 84.945 119.625 ;
        RECT 87.535 119.435 87.705 119.625 ;
        RECT 90.290 119.485 90.410 119.595 ;
        RECT 91.215 119.435 91.385 119.625 ;
        RECT 91.675 119.455 91.845 119.645 ;
        RECT 96.275 119.435 96.445 119.625 ;
        RECT 97.195 119.455 97.365 119.645 ;
        RECT 97.655 119.435 97.825 119.625 ;
        RECT 100.885 119.490 101.045 119.600 ;
        RECT 21.130 119.405 22.065 119.435 ;
        RECT 19.000 119.205 22.065 119.405 ;
        RECT 16.865 118.525 17.795 118.755 ;
        RECT 18.855 118.725 22.065 119.205 ;
        RECT 22.075 118.755 29.385 119.435 ;
        RECT 29.580 118.755 31.415 119.435 ;
        RECT 31.735 118.755 39.045 119.435 ;
        RECT 18.855 118.525 19.785 118.725 ;
        RECT 21.115 118.525 22.065 118.725 ;
        RECT 25.590 118.535 26.500 118.755 ;
        RECT 28.035 118.525 29.385 118.755 ;
        RECT 30.485 118.525 31.415 118.755 ;
        RECT 35.250 118.535 36.160 118.755 ;
        RECT 37.695 118.525 39.045 118.755 ;
        RECT 39.105 118.565 39.535 119.350 ;
        RECT 39.555 118.525 42.305 119.435 ;
        RECT 42.475 118.615 44.405 119.435 ;
        RECT 44.615 118.625 46.445 119.435 ;
        RECT 43.455 118.525 44.405 118.615 ;
        RECT 46.915 118.525 48.730 119.435 ;
        RECT 48.755 118.755 56.065 119.435 ;
        RECT 56.115 118.755 60.930 119.435 ;
        RECT 61.285 118.755 64.750 119.435 ;
        RECT 52.270 118.535 53.180 118.755 ;
        RECT 54.715 118.525 56.065 118.755 ;
        RECT 63.830 118.525 64.750 118.755 ;
        RECT 64.865 118.565 65.295 119.350 ;
        RECT 65.315 118.755 72.625 119.435 ;
        RECT 68.830 118.535 69.740 118.755 ;
        RECT 71.275 118.525 72.625 118.755 ;
        RECT 72.985 118.755 74.820 119.435 ;
        RECT 72.985 118.525 73.915 118.755 ;
        RECT 74.975 118.525 76.805 119.435 ;
        RECT 76.815 118.755 84.545 119.435 ;
        RECT 80.330 118.535 81.240 118.755 ;
        RECT 82.775 118.525 84.545 118.755 ;
        RECT 84.635 118.625 87.385 119.435 ;
        RECT 87.395 118.755 90.135 119.435 ;
        RECT 90.625 118.565 91.055 119.350 ;
        RECT 91.075 118.755 95.890 119.435 ;
        RECT 96.145 118.525 97.495 119.435 ;
        RECT 97.515 118.625 98.885 119.435 ;
        RECT 98.895 119.405 100.290 119.435 ;
        RECT 101.335 119.405 101.505 119.625 ;
        RECT 102.715 119.455 102.885 119.645 ;
        RECT 103.170 119.485 103.290 119.595 ;
        RECT 104.095 119.455 104.265 119.675 ;
        RECT 105.310 119.645 106.705 119.675 ;
        RECT 106.715 119.645 109.465 120.455 ;
        RECT 109.475 119.645 112.950 120.555 ;
        RECT 116.670 120.325 117.580 120.545 ;
        RECT 119.115 120.325 120.465 120.555 ;
        RECT 113.155 119.645 120.465 120.325 ;
        RECT 120.825 120.325 121.755 120.555 ;
        RECT 120.825 119.645 122.660 120.325 ;
        RECT 122.815 119.645 128.325 120.455 ;
        RECT 129.265 119.730 129.695 120.515 ;
        RECT 130.765 120.325 131.695 120.555 ;
        RECT 129.860 119.645 131.695 120.325 ;
        RECT 132.325 120.325 133.255 120.555 ;
        RECT 132.325 119.645 134.160 120.325 ;
        RECT 134.315 119.645 135.685 120.455 ;
        RECT 136.180 120.325 137.525 120.555 ;
        RECT 135.695 119.645 137.525 120.325 ;
        RECT 137.535 119.645 138.905 120.455 ;
        RECT 106.855 119.455 107.025 119.645 ;
        RECT 109.620 119.625 109.790 119.645 ;
        RECT 107.310 119.435 107.480 119.625 ;
        RECT 107.775 119.435 107.945 119.625 ;
        RECT 109.615 119.455 109.790 119.625 ;
        RECT 113.295 119.455 113.465 119.645 ;
        RECT 122.495 119.625 122.660 119.645 ;
        RECT 109.615 119.435 109.785 119.455 ;
        RECT 116.050 119.435 116.220 119.625 ;
        RECT 119.735 119.435 119.905 119.625 ;
        RECT 120.195 119.435 120.365 119.625 ;
        RECT 122.495 119.455 122.665 119.625 ;
        RECT 122.955 119.595 123.125 119.645 ;
        RECT 129.860 119.625 130.025 119.645 ;
        RECT 122.950 119.485 123.125 119.595 ;
        RECT 122.955 119.455 123.125 119.485 ;
        RECT 126.630 119.435 126.800 119.625 ;
        RECT 127.095 119.435 127.265 119.625 ;
        RECT 128.485 119.490 128.645 119.600 ;
        RECT 129.855 119.455 130.025 119.625 ;
        RECT 133.995 119.625 134.160 119.645 ;
        RECT 133.995 119.455 134.165 119.625 ;
        RECT 134.455 119.455 134.625 119.645 ;
        RECT 135.835 119.455 136.005 119.645 ;
        RECT 136.765 119.480 136.925 119.590 ;
        RECT 134.460 119.435 134.625 119.455 ;
        RECT 138.595 119.435 138.765 119.645 ;
        RECT 98.895 118.725 101.630 119.405 ;
        RECT 98.895 118.525 100.305 118.725 ;
        RECT 102.055 118.525 107.625 119.435 ;
        RECT 107.635 118.755 109.465 119.435 ;
        RECT 109.475 118.625 113.145 119.435 ;
        RECT 114.175 118.525 116.365 119.435 ;
        RECT 116.385 118.565 116.815 119.350 ;
        RECT 116.835 118.525 120.045 119.435 ;
        RECT 120.055 118.755 122.795 119.435 ;
        RECT 123.470 118.525 126.945 119.435 ;
        RECT 126.955 118.755 134.265 119.435 ;
        RECT 134.460 118.755 136.295 119.435 ;
        RECT 130.470 118.535 131.380 118.755 ;
        RECT 132.915 118.525 134.265 118.755 ;
        RECT 135.365 118.525 136.295 118.755 ;
        RECT 137.535 118.625 138.905 119.435 ;
      LAYER nwell ;
        RECT 13.140 115.405 139.100 118.235 ;
      LAYER pwell ;
        RECT 13.335 114.205 14.705 115.015 ;
        RECT 14.715 114.205 18.385 115.015 ;
        RECT 18.855 114.915 19.805 115.115 ;
        RECT 21.135 114.915 22.065 115.115 ;
        RECT 18.855 114.435 22.065 114.915 ;
        RECT 18.855 114.235 21.920 114.435 ;
        RECT 18.855 114.205 19.790 114.235 ;
        RECT 13.475 113.995 13.645 114.205 ;
        RECT 14.855 113.995 15.025 114.205 ;
        RECT 17.610 114.045 17.730 114.155 ;
        RECT 18.075 113.995 18.245 114.185 ;
        RECT 18.530 114.045 18.650 114.155 ;
        RECT 21.750 114.015 21.920 114.235 ;
        RECT 22.095 114.205 23.445 115.115 ;
        RECT 23.465 114.205 26.195 115.115 ;
        RECT 26.225 114.290 26.655 115.075 ;
        RECT 26.805 114.205 29.805 115.115 ;
        RECT 29.895 114.205 31.725 115.015 ;
        RECT 31.885 114.205 35.540 115.115 ;
        RECT 35.875 114.915 36.825 115.115 ;
        RECT 38.155 114.915 39.085 115.115 ;
        RECT 35.875 114.435 39.085 114.915 ;
        RECT 35.875 114.235 38.940 114.435 ;
        RECT 35.875 114.205 36.810 114.235 ;
        RECT 22.210 114.015 22.380 114.205 ;
        RECT 23.595 114.015 23.765 114.205 ;
        RECT 25.435 113.995 25.605 114.185 ;
        RECT 29.115 113.995 29.285 114.185 ;
        RECT 29.575 114.015 29.745 114.205 ;
        RECT 30.035 114.015 30.205 114.205 ;
        RECT 31.885 114.185 32.045 114.205 ;
        RECT 31.415 114.015 31.585 114.185 ;
        RECT 31.415 113.995 31.565 114.015 ;
        RECT 31.875 113.995 32.045 114.185 ;
        RECT 37.395 113.995 37.565 114.185 ;
        RECT 38.770 114.015 38.940 114.235 ;
        RECT 39.095 114.205 40.465 115.015 ;
        RECT 40.475 114.205 44.130 115.115 ;
        RECT 45.075 114.915 46.025 115.115 ;
        RECT 47.355 114.915 48.285 115.115 ;
        RECT 45.075 114.435 48.285 114.915 ;
        RECT 50.950 114.885 51.870 115.115 ;
        RECT 45.075 114.235 48.140 114.435 ;
        RECT 45.075 114.205 46.010 114.235 ;
        RECT 39.235 114.015 39.405 114.205 ;
        RECT 39.695 113.995 39.865 114.185 ;
        RECT 40.620 114.015 40.790 114.205 ;
        RECT 41.530 114.045 41.650 114.155 ;
        RECT 44.305 114.050 44.465 114.160 ;
        RECT 44.750 113.995 44.920 114.185 ;
        RECT 45.215 113.995 45.385 114.185 ;
        RECT 47.970 114.015 48.140 114.235 ;
        RECT 48.405 114.205 51.870 114.885 ;
        RECT 51.985 114.290 52.415 115.075 ;
        RECT 52.475 114.885 53.825 115.115 ;
        RECT 55.360 114.885 56.270 115.105 ;
        RECT 52.475 114.205 59.785 114.885 ;
        RECT 59.795 114.205 61.165 115.015 ;
        RECT 61.175 114.205 63.925 115.115 ;
        RECT 63.935 114.205 65.305 115.015 ;
        RECT 65.315 114.915 66.270 115.115 ;
        RECT 65.315 114.235 67.595 114.915 ;
        RECT 67.615 114.885 68.535 115.115 ;
        RECT 70.010 114.885 70.930 115.115 ;
        RECT 76.795 114.885 77.725 115.115 ;
        RECT 65.315 114.205 66.270 114.235 ;
        RECT 48.435 114.015 48.605 114.205 ;
        RECT 13.335 113.185 14.705 113.995 ;
        RECT 14.715 113.185 17.465 113.995 ;
        RECT 17.935 113.315 25.245 113.995 ;
        RECT 21.450 113.095 22.360 113.315 ;
        RECT 23.895 113.085 25.245 113.315 ;
        RECT 25.295 113.185 27.125 113.995 ;
        RECT 27.135 113.315 29.425 113.995 ;
        RECT 27.135 113.085 28.055 113.315 ;
        RECT 29.635 113.175 31.565 113.995 ;
        RECT 31.735 113.185 37.245 113.995 ;
        RECT 37.255 113.185 39.085 113.995 ;
        RECT 29.635 113.085 30.585 113.175 ;
        RECT 39.105 113.125 39.535 113.910 ;
        RECT 39.555 113.185 41.385 113.995 ;
        RECT 42.000 113.085 45.065 113.995 ;
        RECT 45.085 113.085 47.815 113.995 ;
        RECT 47.835 113.965 48.785 113.995 ;
        RECT 51.190 113.965 51.360 114.185 ;
        RECT 51.655 114.015 51.825 114.185 ;
        RECT 51.660 113.995 51.825 114.015 ;
        RECT 53.955 113.995 54.125 114.185 ;
        RECT 59.475 114.155 59.645 114.205 ;
        RECT 59.470 114.045 59.645 114.155 ;
        RECT 59.475 114.015 59.645 114.045 ;
        RECT 59.935 114.185 60.105 114.205 ;
        RECT 59.935 114.015 60.110 114.185 ;
        RECT 61.315 114.015 61.485 114.205 ;
        RECT 59.940 113.995 60.110 114.015 ;
        RECT 61.775 113.995 61.945 114.185 ;
        RECT 64.075 114.015 64.245 114.205 ;
        RECT 66.380 113.995 66.550 114.185 ;
        RECT 67.300 114.015 67.470 114.235 ;
        RECT 67.615 114.205 69.905 114.885 ;
        RECT 70.010 114.205 73.475 114.885 ;
        RECT 73.825 114.205 77.725 114.885 ;
        RECT 77.745 114.290 78.175 115.075 ;
        RECT 81.710 114.885 82.620 115.105 ;
        RECT 84.155 114.885 85.925 115.115 ;
        RECT 78.195 114.205 85.925 114.885 ;
        RECT 86.485 114.205 89.225 114.885 ;
        RECT 89.235 114.205 92.905 115.015 ;
        RECT 92.915 114.205 94.285 115.015 ;
        RECT 94.310 114.885 95.680 115.115 ;
        RECT 94.310 114.205 96.585 114.885 ;
        RECT 96.595 114.205 98.805 115.115 ;
        RECT 98.905 114.205 100.255 115.115 ;
        RECT 102.335 115.025 103.285 115.115 ;
        RECT 101.355 114.205 103.285 115.025 ;
        RECT 103.505 114.290 103.935 115.075 ;
        RECT 103.955 114.205 106.145 115.115 ;
        RECT 106.255 114.205 109.925 115.015 ;
        RECT 109.935 114.205 111.305 115.015 ;
        RECT 114.830 114.885 115.740 115.105 ;
        RECT 117.275 114.885 118.625 115.115 ;
        RECT 111.315 114.205 118.625 114.885 ;
        RECT 118.675 114.205 123.490 114.885 ;
        RECT 123.930 114.205 127.405 115.115 ;
        RECT 127.415 114.205 129.245 115.015 ;
        RECT 129.265 114.290 129.695 115.075 ;
        RECT 133.230 114.885 134.140 115.105 ;
        RECT 135.675 114.885 137.025 115.115 ;
        RECT 129.715 114.205 137.025 114.885 ;
        RECT 137.535 114.205 138.905 115.015 ;
        RECT 69.595 113.995 69.765 114.205 ;
        RECT 71.430 113.995 71.600 114.185 ;
        RECT 71.895 113.995 72.065 114.185 ;
        RECT 73.275 114.015 73.445 114.205 ;
        RECT 77.140 114.015 77.310 114.205 ;
        RECT 77.415 113.995 77.585 114.185 ;
        RECT 78.335 114.015 78.505 114.205 ;
        RECT 82.930 114.045 83.050 114.155 ;
        RECT 83.395 113.995 83.565 114.185 ;
        RECT 86.150 114.045 86.270 114.155 ;
        RECT 88.915 114.015 89.085 114.205 ;
        RECT 89.375 114.015 89.545 114.205 ;
        RECT 91.205 113.995 91.375 114.185 ;
        RECT 93.055 114.015 93.225 114.205 ;
        RECT 94.435 113.995 94.605 114.185 ;
        RECT 96.270 114.015 96.440 114.205 ;
        RECT 96.740 114.015 96.910 114.205 ;
        RECT 99.035 114.015 99.205 114.205 ;
        RECT 101.355 114.185 101.505 114.205 ;
        RECT 99.955 113.995 100.125 114.185 ;
        RECT 100.425 114.050 100.585 114.160 ;
        RECT 101.335 114.015 101.505 114.185 ;
        RECT 101.790 114.045 101.910 114.155 ;
        RECT 102.260 113.995 102.430 114.185 ;
        RECT 104.100 114.015 104.270 114.205 ;
        RECT 106.395 114.015 106.565 114.205 ;
        RECT 107.775 114.015 107.945 114.185 ;
        RECT 107.775 113.995 107.940 114.015 ;
        RECT 108.235 113.995 108.405 114.185 ;
        RECT 109.615 114.015 109.785 114.185 ;
        RECT 110.075 114.015 110.245 114.205 ;
        RECT 111.455 114.015 111.625 114.205 ;
        RECT 109.620 113.995 109.785 114.015 ;
        RECT 111.920 113.995 112.090 114.185 ;
        RECT 115.605 114.040 115.765 114.150 ;
        RECT 116.975 113.995 117.145 114.185 ;
        RECT 118.815 114.015 118.985 114.205 ;
        RECT 122.035 113.995 122.205 114.185 ;
        RECT 127.090 113.995 127.260 114.205 ;
        RECT 127.555 113.995 127.725 114.205 ;
        RECT 129.855 114.015 130.025 114.205 ;
        RECT 134.925 114.040 135.085 114.150 ;
        RECT 135.835 113.995 136.005 114.185 ;
        RECT 137.210 114.045 137.330 114.155 ;
        RECT 138.595 113.995 138.765 114.205 ;
        RECT 47.835 113.285 51.505 113.965 ;
        RECT 51.660 113.315 53.495 113.995 ;
        RECT 47.835 113.085 48.785 113.285 ;
        RECT 52.565 113.085 53.495 113.315 ;
        RECT 53.815 113.185 59.325 113.995 ;
        RECT 59.795 113.085 61.625 113.995 ;
        RECT 61.735 113.085 64.845 113.995 ;
        RECT 64.865 113.125 65.295 113.910 ;
        RECT 65.315 113.085 66.665 113.995 ;
        RECT 68.065 113.965 69.905 113.995 ;
        RECT 66.740 113.315 69.905 113.965 ;
        RECT 66.740 113.285 69.420 113.315 ;
        RECT 68.065 113.085 69.420 113.285 ;
        RECT 69.915 113.085 71.745 113.995 ;
        RECT 71.755 113.185 77.265 113.995 ;
        RECT 77.275 113.185 82.785 113.995 ;
        RECT 83.255 113.315 90.565 113.995 ;
        RECT 86.770 113.095 87.680 113.315 ;
        RECT 89.215 113.085 90.565 113.315 ;
        RECT 90.625 113.125 91.055 113.910 ;
        RECT 91.075 113.085 94.285 113.995 ;
        RECT 94.295 113.185 99.805 113.995 ;
        RECT 99.815 113.185 101.645 113.995 ;
        RECT 102.115 113.085 105.590 113.995 ;
        RECT 106.105 113.315 107.940 113.995 ;
        RECT 106.105 113.085 107.035 113.315 ;
        RECT 108.095 113.185 109.465 113.995 ;
        RECT 109.620 113.315 111.455 113.995 ;
        RECT 110.525 113.085 111.455 113.315 ;
        RECT 111.775 113.085 115.250 113.995 ;
        RECT 116.385 113.125 116.815 113.910 ;
        RECT 116.835 113.315 121.650 113.995 ;
        RECT 121.895 113.185 123.725 113.995 ;
        RECT 123.930 113.085 127.405 113.995 ;
        RECT 127.415 113.315 134.725 113.995 ;
        RECT 135.695 113.315 137.525 113.995 ;
        RECT 130.930 113.095 131.840 113.315 ;
        RECT 133.375 113.085 134.725 113.315 ;
        RECT 136.180 113.085 137.525 113.315 ;
        RECT 137.535 113.185 138.905 113.995 ;
      LAYER nwell ;
        RECT 13.140 109.965 139.100 112.795 ;
      LAYER pwell ;
        RECT 13.335 108.765 14.705 109.575 ;
        RECT 14.715 108.765 17.465 109.575 ;
        RECT 20.990 109.445 21.900 109.665 ;
        RECT 23.435 109.445 24.785 109.675 ;
        RECT 17.475 108.765 24.785 109.445 ;
        RECT 24.835 108.765 26.205 109.575 ;
        RECT 26.225 108.850 26.655 109.635 ;
        RECT 28.750 109.445 29.885 109.675 ;
        RECT 26.675 108.765 29.885 109.445 ;
        RECT 29.895 108.765 35.405 109.575 ;
        RECT 35.415 108.765 40.925 109.575 ;
        RECT 40.935 108.765 42.765 109.575 ;
        RECT 44.655 109.445 46.005 109.675 ;
        RECT 47.540 109.445 48.450 109.665 ;
        RECT 42.775 108.765 44.605 109.445 ;
        RECT 44.655 108.765 51.965 109.445 ;
        RECT 51.985 108.850 52.415 109.635 ;
        RECT 55.090 109.445 56.010 109.675 ;
        RECT 52.545 108.765 56.010 109.445 ;
        RECT 56.125 108.765 57.475 109.675 ;
        RECT 57.495 108.765 61.165 109.575 ;
        RECT 61.175 108.765 63.005 109.675 ;
        RECT 66.530 109.445 67.440 109.665 ;
        RECT 68.975 109.445 70.325 109.675 ;
        RECT 63.015 108.765 70.325 109.445 ;
        RECT 70.375 108.765 75.885 109.575 ;
        RECT 75.895 108.765 77.725 109.575 ;
        RECT 77.745 108.850 78.175 109.635 ;
        RECT 79.245 109.445 80.175 109.675 ;
        RECT 78.340 108.765 80.175 109.445 ;
        RECT 80.495 108.765 82.325 109.575 ;
        RECT 82.335 108.765 85.545 109.675 ;
        RECT 91.845 109.445 92.775 109.675 ;
        RECT 86.710 108.765 91.525 109.445 ;
        RECT 91.845 108.765 93.680 109.445 ;
        RECT 93.835 108.765 97.505 109.575 ;
        RECT 97.825 109.445 98.755 109.675 ;
        RECT 97.825 108.765 99.660 109.445 ;
        RECT 100.010 108.765 103.485 109.675 ;
        RECT 103.505 108.850 103.935 109.635 ;
        RECT 107.470 109.445 108.380 109.665 ;
        RECT 109.915 109.445 111.265 109.675 ;
        RECT 103.955 108.765 111.265 109.445 ;
        RECT 111.510 108.765 114.985 109.675 ;
        RECT 119.815 109.585 120.765 109.675 ;
        RECT 114.995 108.765 118.665 109.575 ;
        RECT 118.835 108.765 120.765 109.585 ;
        RECT 121.285 109.445 122.215 109.675 ;
        RECT 121.285 108.765 123.120 109.445 ;
        RECT 123.275 108.765 125.105 109.575 ;
        RECT 125.425 109.445 126.355 109.675 ;
        RECT 125.425 108.765 127.260 109.445 ;
        RECT 127.415 108.765 129.245 109.575 ;
        RECT 129.265 108.850 129.695 109.635 ;
        RECT 129.715 108.765 132.925 109.675 ;
        RECT 134.340 109.445 135.685 109.675 ;
        RECT 136.180 109.445 137.525 109.675 ;
        RECT 133.855 108.765 135.685 109.445 ;
        RECT 135.695 108.765 137.525 109.445 ;
        RECT 137.535 108.765 138.905 109.575 ;
        RECT 13.475 108.555 13.645 108.765 ;
        RECT 14.855 108.555 15.025 108.765 ;
        RECT 17.615 108.745 17.785 108.765 ;
        RECT 17.615 108.575 17.790 108.745 ;
        RECT 17.620 108.555 17.790 108.575 ;
        RECT 21.295 108.555 21.465 108.745 ;
        RECT 21.760 108.555 21.930 108.745 ;
        RECT 24.975 108.575 25.145 108.765 ;
        RECT 26.815 108.575 26.985 108.765 ;
        RECT 27.275 108.555 27.445 108.745 ;
        RECT 27.735 108.555 27.905 108.745 ;
        RECT 30.035 108.575 30.205 108.765 ;
        RECT 33.250 108.605 33.370 108.715 ;
        RECT 33.715 108.555 33.885 108.745 ;
        RECT 35.555 108.575 35.725 108.765 ;
        RECT 36.015 108.555 36.185 108.745 ;
        RECT 38.770 108.605 38.890 108.715 ;
        RECT 40.620 108.555 40.790 108.745 ;
        RECT 41.075 108.555 41.245 108.765 ;
        RECT 42.915 108.575 43.085 108.765 ;
        RECT 43.830 108.605 43.950 108.715 ;
        RECT 44.295 108.575 44.465 108.745 ;
        RECT 46.595 108.575 46.765 108.745 ;
        RECT 44.315 108.555 44.465 108.575 ;
        RECT 46.745 108.555 46.765 108.575 ;
        RECT 49.355 108.555 49.525 108.745 ;
        RECT 51.655 108.575 51.825 108.765 ;
        RECT 52.575 108.575 52.745 108.765 ;
        RECT 53.035 108.575 53.205 108.745 ;
        RECT 56.255 108.575 56.425 108.765 ;
        RECT 53.040 108.555 53.205 108.575 ;
        RECT 57.175 108.555 57.345 108.745 ;
        RECT 57.635 108.555 57.805 108.765 ;
        RECT 61.320 108.555 61.490 108.765 ;
        RECT 63.155 108.575 63.325 108.765 ;
        RECT 65.455 108.555 65.625 108.745 ;
        RECT 70.055 108.555 70.225 108.745 ;
        RECT 70.515 108.555 70.685 108.765 ;
        RECT 74.195 108.555 74.365 108.745 ;
        RECT 76.035 108.575 76.205 108.765 ;
        RECT 78.340 108.745 78.505 108.765 ;
        RECT 78.335 108.575 78.505 108.745 ;
        RECT 80.635 108.575 80.805 108.765 ;
        RECT 81.555 108.555 81.725 108.745 ;
        RECT 82.465 108.575 82.635 108.765 ;
        RECT 85.230 108.605 85.350 108.715 ;
        RECT 85.700 108.555 85.870 108.745 ;
        RECT 89.375 108.555 89.545 108.745 ;
        RECT 91.215 108.575 91.385 108.765 ;
        RECT 93.515 108.745 93.680 108.765 ;
        RECT 93.515 108.575 93.685 108.745 ;
        RECT 93.975 108.555 94.145 108.765 ;
        RECT 99.495 108.745 99.660 108.765 ;
        RECT 103.170 108.745 103.340 108.765 ;
        RECT 94.435 108.555 94.605 108.745 ;
        RECT 99.495 108.575 99.665 108.745 ;
        RECT 99.955 108.555 100.125 108.745 ;
        RECT 102.710 108.605 102.830 108.715 ;
        RECT 103.170 108.575 103.345 108.745 ;
        RECT 104.095 108.575 104.265 108.765 ;
        RECT 103.175 108.555 103.345 108.575 ;
        RECT 110.535 108.555 110.705 108.745 ;
        RECT 113.290 108.605 113.410 108.715 ;
        RECT 113.755 108.575 113.925 108.745 ;
        RECT 114.670 108.575 114.840 108.765 ;
        RECT 115.135 108.575 115.305 108.765 ;
        RECT 118.835 108.745 118.985 108.765 ;
        RECT 116.050 108.605 116.170 108.715 ;
        RECT 113.775 108.555 113.925 108.575 ;
        RECT 116.975 108.555 117.145 108.745 ;
        RECT 118.815 108.575 118.985 108.745 ;
        RECT 122.955 108.745 123.120 108.765 ;
        RECT 122.955 108.575 123.125 108.745 ;
        RECT 123.415 108.575 123.585 108.765 ;
        RECT 127.095 108.745 127.260 108.765 ;
        RECT 125.710 108.555 125.880 108.745 ;
        RECT 126.175 108.555 126.345 108.745 ;
        RECT 127.095 108.575 127.265 108.745 ;
        RECT 127.555 108.575 127.725 108.765 ;
        RECT 132.615 108.575 132.785 108.765 ;
        RECT 133.085 108.610 133.245 108.720 ;
        RECT 133.995 108.575 134.165 108.765 ;
        RECT 135.835 108.575 136.005 108.765 ;
        RECT 136.295 108.555 136.465 108.745 ;
        RECT 136.765 108.600 136.925 108.710 ;
        RECT 138.595 108.555 138.765 108.765 ;
        RECT 13.335 107.745 14.705 108.555 ;
        RECT 14.715 107.745 17.465 108.555 ;
        RECT 17.475 107.645 19.305 108.555 ;
        RECT 19.315 107.875 21.605 108.555 ;
        RECT 19.315 107.645 20.235 107.875 ;
        RECT 21.615 107.645 24.535 108.555 ;
        RECT 24.845 107.645 27.575 108.555 ;
        RECT 27.595 107.745 33.105 108.555 ;
        RECT 33.575 107.875 35.865 108.555 ;
        RECT 34.945 107.645 35.865 107.875 ;
        RECT 35.885 107.645 38.615 108.555 ;
        RECT 39.105 107.685 39.535 108.470 ;
        RECT 39.555 107.645 40.905 108.555 ;
        RECT 40.935 107.745 43.685 108.555 ;
        RECT 44.315 107.735 46.245 108.555 ;
        RECT 46.745 107.875 49.195 108.555 ;
        RECT 49.325 107.875 52.790 108.555 ;
        RECT 53.040 107.875 54.875 108.555 ;
        RECT 45.295 107.645 46.245 107.735 ;
        RECT 47.235 107.645 49.195 107.875 ;
        RECT 51.870 107.645 52.790 107.875 ;
        RECT 53.945 107.645 54.875 107.875 ;
        RECT 55.195 107.875 57.485 108.555 ;
        RECT 55.195 107.645 56.115 107.875 ;
        RECT 57.495 107.745 61.165 108.555 ;
        RECT 61.175 107.645 64.845 108.555 ;
        RECT 64.865 107.685 65.295 108.470 ;
        RECT 65.315 107.745 66.685 108.555 ;
        RECT 66.790 107.875 70.255 108.555 ;
        RECT 66.790 107.645 67.710 107.875 ;
        RECT 70.375 107.745 74.045 108.555 ;
        RECT 74.055 107.875 81.365 108.555 ;
        RECT 77.570 107.655 78.480 107.875 ;
        RECT 80.015 107.645 81.365 107.875 ;
        RECT 81.415 107.745 85.085 108.555 ;
        RECT 85.555 107.645 89.030 108.555 ;
        RECT 89.235 107.745 90.605 108.555 ;
        RECT 90.625 107.685 91.055 108.470 ;
        RECT 91.075 107.645 94.285 108.555 ;
        RECT 94.295 107.745 99.805 108.555 ;
        RECT 99.815 107.745 102.565 108.555 ;
        RECT 103.035 107.875 110.345 108.555 ;
        RECT 106.550 107.655 107.460 107.875 ;
        RECT 108.995 107.645 110.345 107.875 ;
        RECT 110.395 107.745 113.145 108.555 ;
        RECT 113.775 107.735 115.705 108.555 ;
        RECT 114.755 107.645 115.705 107.735 ;
        RECT 116.385 107.685 116.815 108.470 ;
        RECT 116.835 107.745 122.345 108.555 ;
        RECT 122.550 107.645 126.025 108.555 ;
        RECT 126.035 107.875 133.345 108.555 ;
        RECT 129.550 107.655 130.460 107.875 ;
        RECT 131.995 107.645 133.345 107.875 ;
        RECT 133.395 107.645 136.605 108.555 ;
        RECT 137.535 107.745 138.905 108.555 ;
      LAYER nwell ;
        RECT 13.140 104.525 139.100 107.355 ;
      LAYER pwell ;
        RECT 13.335 103.325 14.705 104.135 ;
        RECT 14.715 103.325 20.225 104.135 ;
        RECT 20.235 103.325 22.065 104.135 ;
        RECT 23.125 104.005 24.055 104.235 ;
        RECT 22.220 103.325 24.055 104.005 ;
        RECT 24.375 103.325 26.205 104.135 ;
        RECT 26.225 103.410 26.655 104.195 ;
        RECT 26.675 103.325 30.345 104.135 ;
        RECT 30.355 103.325 31.725 104.135 ;
        RECT 32.045 104.005 32.975 104.235 ;
        RECT 37.550 104.005 38.460 104.225 ;
        RECT 39.995 104.005 41.345 104.235 ;
        RECT 32.045 103.325 33.880 104.005 ;
        RECT 34.035 103.325 41.345 104.005 ;
        RECT 41.435 104.005 42.785 104.235 ;
        RECT 44.320 104.005 45.230 104.225 ;
        RECT 48.755 104.035 49.685 104.235 ;
        RECT 51.015 104.035 51.965 104.235 ;
        RECT 41.435 103.325 48.745 104.005 ;
        RECT 48.755 103.555 51.965 104.035 ;
        RECT 48.900 103.355 51.965 103.555 ;
        RECT 51.985 103.410 52.415 104.195 ;
        RECT 52.475 104.005 53.825 104.235 ;
        RECT 55.360 104.005 56.270 104.225 ;
        RECT 63.770 104.005 64.680 104.225 ;
        RECT 66.215 104.005 67.565 104.235 ;
        RECT 13.475 103.115 13.645 103.325 ;
        RECT 14.855 103.115 15.025 103.325 ;
        RECT 17.610 103.115 17.780 103.305 ;
        RECT 20.375 103.135 20.545 103.325 ;
        RECT 22.220 103.305 22.385 103.325 ;
        RECT 21.295 103.115 21.465 103.305 ;
        RECT 22.215 103.135 22.385 103.305 ;
        RECT 24.515 103.135 24.685 103.325 ;
        RECT 26.815 103.135 26.985 103.325 ;
        RECT 28.655 103.115 28.825 103.305 ;
        RECT 30.495 103.135 30.665 103.325 ;
        RECT 33.715 103.305 33.880 103.325 ;
        RECT 30.955 103.115 31.125 103.305 ;
        RECT 31.415 103.115 31.585 103.305 ;
        RECT 33.715 103.135 33.885 103.305 ;
        RECT 34.175 103.135 34.345 103.325 ;
        RECT 35.090 103.165 35.210 103.275 ;
        RECT 13.335 102.305 14.705 103.115 ;
        RECT 14.715 102.305 17.465 103.115 ;
        RECT 17.495 102.205 18.845 103.115 ;
        RECT 18.855 102.435 21.605 103.115 ;
        RECT 21.655 102.435 28.965 103.115 ;
        RECT 28.975 102.435 31.265 103.115 ;
        RECT 18.855 102.205 19.785 102.435 ;
        RECT 21.655 102.205 23.005 102.435 ;
        RECT 24.540 102.215 25.450 102.435 ;
        RECT 28.975 102.205 29.895 102.435 ;
        RECT 31.275 102.305 34.945 103.115 ;
        RECT 35.415 103.085 36.350 103.115 ;
        RECT 38.310 103.085 38.480 103.305 ;
        RECT 38.770 103.165 38.890 103.275 ;
        RECT 39.695 103.115 39.865 103.305 ;
        RECT 41.995 103.115 42.165 103.305 ;
        RECT 44.750 103.165 44.870 103.275 ;
        RECT 45.215 103.135 45.385 103.305 ;
        RECT 48.435 103.135 48.605 103.325 ;
        RECT 48.900 103.135 49.070 103.355 ;
        RECT 51.030 103.325 51.965 103.355 ;
        RECT 52.475 103.325 59.785 104.005 ;
        RECT 60.255 103.325 67.565 104.005 ;
        RECT 67.615 103.325 73.125 104.135 ;
        RECT 73.135 103.325 74.965 104.135 ;
        RECT 75.745 104.005 76.675 104.235 ;
        RECT 75.745 103.325 77.580 104.005 ;
        RECT 77.745 103.410 78.175 104.195 ;
        RECT 78.195 103.325 81.670 104.235 ;
        RECT 82.335 103.325 85.545 104.235 ;
        RECT 89.070 104.005 89.980 104.225 ;
        RECT 91.515 104.005 92.865 104.235 ;
        RECT 85.555 103.325 92.865 104.005 ;
        RECT 93.225 104.005 94.155 104.235 ;
        RECT 93.225 103.325 95.060 104.005 ;
        RECT 95.675 103.325 97.865 104.235 ;
        RECT 98.175 104.145 99.125 104.235 ;
        RECT 98.175 103.325 100.105 104.145 ;
        RECT 100.275 103.325 103.025 104.135 ;
        RECT 103.505 103.410 103.935 104.195 ;
        RECT 103.955 103.325 107.625 104.135 ;
        RECT 107.635 103.325 109.005 104.135 ;
        RECT 109.015 103.325 111.205 104.235 ;
        RECT 114.830 104.005 115.740 104.225 ;
        RECT 117.275 104.005 118.625 104.235 ;
        RECT 111.315 103.325 118.625 104.005 ;
        RECT 118.675 103.325 124.185 104.135 ;
        RECT 124.965 104.005 125.895 104.235 ;
        RECT 127.265 104.005 128.195 104.235 ;
        RECT 124.965 103.325 126.800 104.005 ;
        RECT 127.265 103.325 129.100 104.005 ;
        RECT 129.265 103.410 129.695 104.195 ;
        RECT 129.715 103.325 132.925 104.235 ;
        RECT 133.985 104.005 134.915 104.235 ;
        RECT 136.180 104.005 137.525 104.235 ;
        RECT 133.080 103.325 134.915 104.005 ;
        RECT 135.695 103.325 137.525 104.005 ;
        RECT 137.535 103.325 138.905 104.135 ;
        RECT 45.220 103.115 45.385 103.135 ;
        RECT 54.415 103.115 54.585 103.305 ;
        RECT 54.875 103.115 55.045 103.305 ;
        RECT 59.475 103.135 59.645 103.325 ;
        RECT 59.930 103.165 60.050 103.275 ;
        RECT 60.395 103.115 60.565 103.325 ;
        RECT 64.085 103.160 64.245 103.270 ;
        RECT 65.455 103.115 65.625 103.305 ;
        RECT 67.755 103.135 67.925 103.325 ;
        RECT 70.975 103.115 71.145 103.305 ;
        RECT 73.275 103.135 73.445 103.325 ;
        RECT 77.415 103.305 77.580 103.325 ;
        RECT 73.730 103.165 73.850 103.275 ;
        RECT 74.200 103.115 74.370 103.305 ;
        RECT 75.110 103.165 75.230 103.275 ;
        RECT 77.415 103.135 77.585 103.305 ;
        RECT 78.340 103.135 78.510 103.325 ;
        RECT 79.715 103.135 79.885 103.305 ;
        RECT 79.715 103.115 79.880 103.135 ;
        RECT 80.175 103.115 80.345 103.305 ;
        RECT 82.010 103.165 82.130 103.275 ;
        RECT 82.465 103.135 82.635 103.325 ;
        RECT 82.925 103.115 83.095 103.305 ;
        RECT 85.695 103.135 85.865 103.325 ;
        RECT 94.895 103.305 95.060 103.325 ;
        RECT 86.150 103.165 86.270 103.275 ;
        RECT 86.620 103.115 86.790 103.305 ;
        RECT 90.290 103.165 90.410 103.275 ;
        RECT 91.215 103.115 91.385 103.305 ;
        RECT 94.895 103.135 95.065 103.305 ;
        RECT 95.350 103.165 95.470 103.275 ;
        RECT 95.820 103.135 95.990 103.325 ;
        RECT 99.955 103.305 100.105 103.325 ;
        RECT 96.735 103.115 96.905 103.305 ;
        RECT 98.575 103.115 98.745 103.305 ;
        RECT 99.955 103.135 100.125 103.305 ;
        RECT 100.415 103.135 100.585 103.325 ;
        RECT 103.170 103.165 103.290 103.275 ;
        RECT 104.095 103.135 104.265 103.325 ;
        RECT 105.935 103.115 106.105 103.305 ;
        RECT 107.775 103.135 107.945 103.325 ;
        RECT 109.160 103.135 109.330 103.325 ;
        RECT 110.535 103.115 110.705 103.305 ;
        RECT 110.995 103.115 111.165 103.305 ;
        RECT 111.455 103.135 111.625 103.325 ;
        RECT 112.840 103.115 113.010 103.305 ;
        RECT 116.975 103.115 117.145 103.305 ;
        RECT 118.815 103.135 118.985 103.325 ;
        RECT 126.635 103.305 126.800 103.325 ;
        RECT 128.935 103.305 129.100 103.325 ;
        RECT 124.330 103.165 124.450 103.275 ;
        RECT 126.635 103.135 126.805 103.305 ;
        RECT 128.010 103.115 128.180 103.305 ;
        RECT 128.475 103.115 128.645 103.305 ;
        RECT 128.935 103.135 129.105 103.305 ;
        RECT 132.615 103.135 132.785 103.325 ;
        RECT 133.080 103.305 133.245 103.325 ;
        RECT 133.075 103.135 133.245 103.305 ;
        RECT 135.370 103.165 135.490 103.275 ;
        RECT 135.835 103.115 136.005 103.325 ;
        RECT 138.595 103.115 138.765 103.325 ;
        RECT 35.415 102.885 38.480 103.085 ;
        RECT 35.415 102.405 38.625 102.885 ;
        RECT 35.415 102.205 36.365 102.405 ;
        RECT 37.695 102.205 38.625 102.405 ;
        RECT 39.105 102.245 39.535 103.030 ;
        RECT 39.555 102.435 41.845 103.115 ;
        RECT 40.925 102.205 41.845 102.435 ;
        RECT 41.855 102.305 44.605 103.115 ;
        RECT 45.220 102.435 47.055 103.115 ;
        RECT 46.125 102.205 47.055 102.435 ;
        RECT 47.415 102.435 54.725 103.115 ;
        RECT 47.415 102.205 48.765 102.435 ;
        RECT 50.300 102.215 51.210 102.435 ;
        RECT 54.735 102.305 60.245 103.115 ;
        RECT 60.255 102.305 63.925 103.115 ;
        RECT 64.865 102.245 65.295 103.030 ;
        RECT 65.315 102.305 70.825 103.115 ;
        RECT 70.835 102.305 73.585 103.115 ;
        RECT 74.055 102.205 77.530 103.115 ;
        RECT 78.045 102.435 79.880 103.115 ;
        RECT 78.045 102.205 78.975 102.435 ;
        RECT 80.035 102.305 82.785 103.115 ;
        RECT 82.795 102.205 86.005 103.115 ;
        RECT 86.475 102.205 89.950 103.115 ;
        RECT 90.625 102.245 91.055 103.030 ;
        RECT 91.075 102.305 96.585 103.115 ;
        RECT 96.595 102.305 98.425 103.115 ;
        RECT 98.435 102.435 105.745 103.115 ;
        RECT 101.950 102.215 102.860 102.435 ;
        RECT 104.395 102.205 105.745 102.435 ;
        RECT 105.795 102.305 107.625 103.115 ;
        RECT 107.635 102.205 110.845 103.115 ;
        RECT 110.855 102.305 112.685 103.115 ;
        RECT 112.695 102.205 116.170 103.115 ;
        RECT 116.385 102.245 116.815 103.030 ;
        RECT 116.835 102.435 124.145 103.115 ;
        RECT 120.350 102.215 121.260 102.435 ;
        RECT 122.795 102.205 124.145 102.435 ;
        RECT 124.850 102.205 128.325 103.115 ;
        RECT 128.335 102.435 135.645 103.115 ;
        RECT 135.695 102.435 137.525 103.115 ;
        RECT 131.850 102.215 132.760 102.435 ;
        RECT 134.295 102.205 135.645 102.435 ;
        RECT 136.180 102.205 137.525 102.435 ;
        RECT 137.535 102.305 138.905 103.115 ;
      LAYER nwell ;
        RECT 13.140 99.085 139.100 101.915 ;
      LAYER pwell ;
        RECT 13.335 97.885 14.705 98.695 ;
        RECT 14.715 97.885 18.385 98.695 ;
        RECT 21.910 98.565 22.820 98.785 ;
        RECT 24.355 98.565 25.705 98.795 ;
        RECT 18.395 97.885 25.705 98.565 ;
        RECT 26.225 97.970 26.655 98.755 ;
        RECT 26.675 97.885 32.185 98.695 ;
        RECT 32.195 97.885 37.705 98.695 ;
        RECT 37.715 97.885 43.225 98.695 ;
        RECT 43.235 97.885 48.745 98.695 ;
        RECT 48.755 97.885 50.105 98.795 ;
        RECT 50.135 97.885 51.965 98.695 ;
        RECT 51.985 97.970 52.415 98.755 ;
        RECT 52.435 97.885 57.945 98.695 ;
        RECT 57.955 97.885 63.465 98.695 ;
        RECT 63.475 97.885 68.985 98.695 ;
        RECT 68.995 97.885 70.365 98.695 ;
        RECT 73.890 98.565 74.800 98.785 ;
        RECT 76.335 98.565 77.685 98.795 ;
        RECT 70.375 97.885 77.685 98.565 ;
        RECT 77.745 97.970 78.175 98.755 ;
        RECT 78.195 97.885 81.670 98.795 ;
        RECT 82.820 98.565 84.165 98.795 ;
        RECT 82.335 97.885 84.165 98.565 ;
        RECT 84.175 97.885 86.925 98.695 ;
        RECT 86.935 97.885 90.145 98.795 ;
        RECT 90.155 97.885 95.665 98.695 ;
        RECT 95.675 97.885 97.505 98.695 ;
        RECT 97.975 97.885 101.450 98.795 ;
        RECT 101.655 98.565 103.000 98.795 ;
        RECT 101.655 97.885 103.485 98.565 ;
        RECT 103.505 97.970 103.935 98.755 ;
        RECT 104.265 98.565 105.195 98.795 ;
        RECT 104.265 97.885 106.100 98.565 ;
        RECT 106.255 97.885 111.765 98.695 ;
        RECT 111.775 97.885 113.605 98.695 ;
        RECT 115.125 98.565 116.055 98.795 ;
        RECT 116.860 98.565 118.205 98.795 ;
        RECT 114.220 97.885 116.055 98.565 ;
        RECT 116.375 97.885 118.205 98.565 ;
        RECT 118.215 97.885 123.725 98.695 ;
        RECT 123.735 97.885 125.565 98.695 ;
        RECT 125.770 97.885 129.245 98.795 ;
        RECT 129.265 97.970 129.695 98.755 ;
        RECT 133.230 98.565 134.140 98.785 ;
        RECT 135.675 98.565 137.025 98.795 ;
        RECT 129.715 97.885 137.025 98.565 ;
        RECT 137.535 97.885 138.905 98.695 ;
        RECT 13.475 97.675 13.645 97.885 ;
        RECT 14.855 97.675 15.025 97.885 ;
        RECT 18.535 97.695 18.705 97.885 ;
        RECT 20.375 97.675 20.545 97.865 ;
        RECT 25.895 97.835 26.065 97.865 ;
        RECT 25.890 97.725 26.065 97.835 ;
        RECT 25.895 97.675 26.065 97.725 ;
        RECT 26.815 97.695 26.985 97.885 ;
        RECT 31.415 97.675 31.585 97.865 ;
        RECT 32.335 97.695 32.505 97.885 ;
        RECT 36.935 97.675 37.105 97.865 ;
        RECT 37.855 97.695 38.025 97.885 ;
        RECT 38.770 97.725 38.890 97.835 ;
        RECT 39.695 97.675 39.865 97.865 ;
        RECT 43.375 97.695 43.545 97.885 ;
        RECT 45.215 97.675 45.385 97.865 ;
        RECT 49.820 97.695 49.990 97.885 ;
        RECT 50.275 97.695 50.445 97.885 ;
        RECT 50.735 97.675 50.905 97.865 ;
        RECT 52.575 97.695 52.745 97.885 ;
        RECT 56.255 97.675 56.425 97.865 ;
        RECT 58.095 97.695 58.265 97.885 ;
        RECT 61.775 97.675 61.945 97.865 ;
        RECT 63.615 97.695 63.785 97.885 ;
        RECT 64.530 97.725 64.650 97.835 ;
        RECT 65.455 97.675 65.625 97.865 ;
        RECT 69.135 97.695 69.305 97.885 ;
        RECT 70.515 97.695 70.685 97.885 ;
        RECT 78.340 97.865 78.510 97.885 ;
        RECT 70.975 97.675 71.145 97.865 ;
        RECT 78.335 97.695 78.510 97.865 ;
        RECT 78.335 97.675 78.505 97.695 ;
        RECT 79.720 97.675 79.890 97.865 ;
        RECT 82.010 97.725 82.130 97.835 ;
        RECT 82.475 97.695 82.645 97.885 ;
        RECT 83.400 97.675 83.570 97.865 ;
        RECT 84.315 97.695 84.485 97.885 ;
        RECT 89.835 97.675 90.005 97.885 ;
        RECT 90.295 97.835 90.465 97.885 ;
        RECT 90.290 97.725 90.465 97.835 ;
        RECT 90.295 97.695 90.465 97.725 ;
        RECT 91.215 97.695 91.385 97.865 ;
        RECT 95.815 97.695 95.985 97.885 ;
        RECT 91.220 97.675 91.385 97.695 ;
        RECT 96.730 97.675 96.900 97.865 ;
        RECT 97.195 97.675 97.365 97.865 ;
        RECT 97.650 97.725 97.770 97.835 ;
        RECT 98.120 97.695 98.290 97.885 ;
        RECT 98.575 97.675 98.745 97.865 ;
        RECT 103.175 97.695 103.345 97.885 ;
        RECT 105.935 97.865 106.100 97.885 ;
        RECT 105.935 97.695 106.110 97.865 ;
        RECT 106.395 97.695 106.565 97.885 ;
        RECT 105.940 97.675 106.110 97.695 ;
        RECT 109.615 97.675 109.785 97.865 ;
        RECT 111.915 97.695 112.085 97.885 ;
        RECT 114.220 97.865 114.385 97.885 ;
        RECT 112.835 97.675 113.005 97.865 ;
        RECT 113.750 97.725 113.870 97.835 ;
        RECT 114.215 97.695 114.385 97.865 ;
        RECT 116.515 97.695 116.685 97.885 ;
        RECT 118.355 97.695 118.525 97.885 ;
        RECT 114.220 97.675 114.385 97.695 ;
        RECT 120.190 97.675 120.360 97.865 ;
        RECT 120.650 97.725 120.770 97.835 ;
        RECT 121.120 97.675 121.290 97.865 ;
        RECT 123.875 97.695 124.045 97.885 ;
        RECT 124.790 97.725 124.910 97.835 ;
        RECT 128.930 97.695 129.100 97.885 ;
        RECT 129.855 97.695 130.025 97.885 ;
        RECT 132.155 97.675 132.325 97.865 ;
        RECT 132.615 97.675 132.785 97.865 ;
        RECT 133.995 97.675 134.165 97.865 ;
        RECT 135.835 97.675 136.005 97.865 ;
        RECT 137.210 97.725 137.330 97.835 ;
        RECT 138.595 97.675 138.765 97.885 ;
        RECT 13.335 96.865 14.705 97.675 ;
        RECT 14.715 96.865 20.225 97.675 ;
        RECT 20.235 96.865 25.745 97.675 ;
        RECT 25.755 96.865 31.265 97.675 ;
        RECT 31.275 96.865 36.785 97.675 ;
        RECT 36.795 96.865 38.625 97.675 ;
        RECT 39.105 96.805 39.535 97.590 ;
        RECT 39.555 96.865 45.065 97.675 ;
        RECT 45.075 96.865 50.585 97.675 ;
        RECT 50.595 96.865 56.105 97.675 ;
        RECT 56.115 96.865 61.625 97.675 ;
        RECT 61.635 96.865 64.385 97.675 ;
        RECT 64.865 96.805 65.295 97.590 ;
        RECT 65.315 96.865 70.825 97.675 ;
        RECT 70.835 96.995 78.145 97.675 ;
        RECT 74.350 96.775 75.260 96.995 ;
        RECT 76.795 96.765 78.145 96.995 ;
        RECT 78.195 96.865 79.565 97.675 ;
        RECT 79.575 96.765 83.050 97.675 ;
        RECT 83.255 96.765 86.730 97.675 ;
        RECT 86.935 96.765 90.145 97.675 ;
        RECT 90.625 96.805 91.055 97.590 ;
        RECT 91.220 96.995 93.055 97.675 ;
        RECT 92.125 96.765 93.055 96.995 ;
        RECT 93.570 96.765 97.045 97.675 ;
        RECT 97.055 96.865 98.425 97.675 ;
        RECT 98.435 96.995 105.745 97.675 ;
        RECT 101.950 96.775 102.860 96.995 ;
        RECT 104.395 96.765 105.745 96.995 ;
        RECT 105.795 96.765 109.270 97.675 ;
        RECT 109.475 96.765 112.685 97.675 ;
        RECT 112.695 96.865 114.065 97.675 ;
        RECT 114.220 96.995 116.055 97.675 ;
        RECT 115.125 96.765 116.055 96.995 ;
        RECT 116.385 96.805 116.815 97.590 ;
        RECT 117.030 96.765 120.505 97.675 ;
        RECT 120.975 96.765 124.450 97.675 ;
        RECT 125.155 96.995 132.465 97.675 ;
        RECT 125.155 96.765 126.505 96.995 ;
        RECT 128.040 96.775 128.950 96.995 ;
        RECT 132.475 96.865 133.845 97.675 ;
        RECT 133.855 96.995 135.685 97.675 ;
        RECT 135.695 96.995 137.525 97.675 ;
        RECT 134.340 96.765 135.685 96.995 ;
        RECT 136.180 96.765 137.525 96.995 ;
        RECT 137.535 96.865 138.905 97.675 ;
      LAYER nwell ;
        RECT 13.140 93.645 139.100 96.475 ;
      LAYER pwell ;
        RECT 13.335 92.445 14.705 93.255 ;
        RECT 14.715 92.445 20.225 93.255 ;
        RECT 20.235 92.445 25.745 93.255 ;
        RECT 26.225 92.530 26.655 93.315 ;
        RECT 26.675 92.445 32.185 93.255 ;
        RECT 32.195 92.445 37.705 93.255 ;
        RECT 37.715 92.445 43.225 93.255 ;
        RECT 43.235 92.445 48.745 93.255 ;
        RECT 48.755 92.445 51.505 93.255 ;
        RECT 51.985 92.530 52.415 93.315 ;
        RECT 52.435 92.445 57.945 93.255 ;
        RECT 57.955 92.445 63.465 93.255 ;
        RECT 63.475 92.445 68.985 93.255 ;
        RECT 68.995 92.445 74.505 93.255 ;
        RECT 74.515 92.445 77.265 93.255 ;
        RECT 77.745 92.530 78.175 93.315 ;
        RECT 81.710 93.125 82.620 93.345 ;
        RECT 84.155 93.125 85.505 93.355 ;
        RECT 78.195 92.445 85.505 93.125 ;
        RECT 85.555 92.445 86.925 93.255 ;
        RECT 90.450 93.125 91.360 93.345 ;
        RECT 92.895 93.125 94.245 93.355 ;
        RECT 97.810 93.125 98.720 93.345 ;
        RECT 100.255 93.125 101.605 93.355 ;
        RECT 86.935 92.445 94.245 93.125 ;
        RECT 94.295 92.445 101.605 93.125 ;
        RECT 101.655 92.445 103.485 93.125 ;
        RECT 103.505 92.530 103.935 93.315 ;
        RECT 103.955 92.445 107.430 93.355 ;
        RECT 107.635 92.445 110.845 93.355 ;
        RECT 111.355 93.125 112.705 93.355 ;
        RECT 114.240 93.125 115.150 93.345 ;
        RECT 122.190 93.125 123.100 93.345 ;
        RECT 124.635 93.125 125.985 93.355 ;
        RECT 111.355 92.445 118.665 93.125 ;
        RECT 118.675 92.445 125.985 93.125 ;
        RECT 126.345 93.125 127.275 93.355 ;
        RECT 126.345 92.445 128.180 93.125 ;
        RECT 129.265 92.530 129.695 93.315 ;
        RECT 129.910 92.445 133.385 93.355 ;
        RECT 133.395 92.445 135.225 93.255 ;
        RECT 136.180 93.125 137.525 93.355 ;
        RECT 135.695 92.445 137.525 93.125 ;
        RECT 137.535 92.445 138.905 93.255 ;
        RECT 13.475 92.235 13.645 92.445 ;
        RECT 14.855 92.235 15.025 92.445 ;
        RECT 20.375 92.235 20.545 92.445 ;
        RECT 25.895 92.395 26.065 92.425 ;
        RECT 25.890 92.285 26.065 92.395 ;
        RECT 25.895 92.235 26.065 92.285 ;
        RECT 26.815 92.255 26.985 92.445 ;
        RECT 31.415 92.235 31.585 92.425 ;
        RECT 32.335 92.255 32.505 92.445 ;
        RECT 36.935 92.235 37.105 92.425 ;
        RECT 37.855 92.255 38.025 92.445 ;
        RECT 38.770 92.285 38.890 92.395 ;
        RECT 39.695 92.235 39.865 92.425 ;
        RECT 43.375 92.255 43.545 92.445 ;
        RECT 45.215 92.235 45.385 92.425 ;
        RECT 48.895 92.255 49.065 92.445 ;
        RECT 50.735 92.235 50.905 92.425 ;
        RECT 51.650 92.285 51.770 92.395 ;
        RECT 52.575 92.255 52.745 92.445 ;
        RECT 56.255 92.235 56.425 92.425 ;
        RECT 58.095 92.255 58.265 92.445 ;
        RECT 61.775 92.235 61.945 92.425 ;
        RECT 63.615 92.255 63.785 92.445 ;
        RECT 64.530 92.285 64.650 92.395 ;
        RECT 65.455 92.235 65.625 92.425 ;
        RECT 69.135 92.255 69.305 92.445 ;
        RECT 70.975 92.235 71.145 92.425 ;
        RECT 74.655 92.255 74.825 92.445 ;
        RECT 76.495 92.235 76.665 92.425 ;
        RECT 77.410 92.285 77.530 92.395 ;
        RECT 78.335 92.255 78.505 92.445 ;
        RECT 85.695 92.255 85.865 92.445 ;
        RECT 87.075 92.255 87.245 92.445 ;
        RECT 87.995 92.255 88.165 92.425 ;
        RECT 85.695 92.235 85.860 92.255 ;
        RECT 87.995 92.235 88.160 92.255 ;
        RECT 88.455 92.235 88.625 92.425 ;
        RECT 90.290 92.285 90.410 92.395 ;
        RECT 91.220 92.235 91.390 92.425 ;
        RECT 94.435 92.255 94.605 92.445 ;
        RECT 94.890 92.285 95.010 92.395 ;
        RECT 97.195 92.255 97.365 92.425 ;
        RECT 101.795 92.255 101.965 92.445 ;
        RECT 104.100 92.255 104.270 92.445 ;
        RECT 97.195 92.235 97.360 92.255 ;
        RECT 104.555 92.235 104.725 92.425 ;
        RECT 105.015 92.255 105.185 92.425 ;
        RECT 105.020 92.235 105.185 92.255 ;
        RECT 107.315 92.235 107.485 92.425 ;
        RECT 107.775 92.255 107.945 92.445 ;
        RECT 110.990 92.285 111.110 92.395 ;
        RECT 111.915 92.235 112.085 92.425 ;
        RECT 112.375 92.235 112.545 92.425 ;
        RECT 115.605 92.280 115.765 92.390 ;
        RECT 116.980 92.235 117.150 92.425 ;
        RECT 118.355 92.255 118.525 92.445 ;
        RECT 118.815 92.255 118.985 92.445 ;
        RECT 128.015 92.425 128.180 92.445 ;
        RECT 120.650 92.285 120.770 92.395 ;
        RECT 121.115 92.235 121.285 92.425 ;
        RECT 128.015 92.255 128.185 92.425 ;
        RECT 128.475 92.255 128.645 92.425 ;
        RECT 128.480 92.235 128.645 92.255 ;
        RECT 130.775 92.235 130.945 92.425 ;
        RECT 133.070 92.255 133.240 92.445 ;
        RECT 133.535 92.255 133.705 92.445 ;
        RECT 134.455 92.235 134.625 92.425 ;
        RECT 135.370 92.285 135.490 92.395 ;
        RECT 135.835 92.235 136.005 92.445 ;
        RECT 138.595 92.235 138.765 92.445 ;
        RECT 13.335 91.425 14.705 92.235 ;
        RECT 14.715 91.425 20.225 92.235 ;
        RECT 20.235 91.425 25.745 92.235 ;
        RECT 25.755 91.425 31.265 92.235 ;
        RECT 31.275 91.425 36.785 92.235 ;
        RECT 36.795 91.425 38.625 92.235 ;
        RECT 39.105 91.365 39.535 92.150 ;
        RECT 39.555 91.425 45.065 92.235 ;
        RECT 45.075 91.425 50.585 92.235 ;
        RECT 50.595 91.425 56.105 92.235 ;
        RECT 56.115 91.425 61.625 92.235 ;
        RECT 61.635 91.425 64.385 92.235 ;
        RECT 64.865 91.365 65.295 92.150 ;
        RECT 65.315 91.425 70.825 92.235 ;
        RECT 70.835 91.425 76.345 92.235 ;
        RECT 76.355 91.555 83.665 92.235 ;
        RECT 79.870 91.335 80.780 91.555 ;
        RECT 82.315 91.325 83.665 91.555 ;
        RECT 84.025 91.555 85.860 92.235 ;
        RECT 86.325 91.555 88.160 92.235 ;
        RECT 84.025 91.325 84.955 91.555 ;
        RECT 86.325 91.325 87.255 91.555 ;
        RECT 88.315 91.425 90.145 92.235 ;
        RECT 90.625 91.365 91.055 92.150 ;
        RECT 91.075 91.325 94.550 92.235 ;
        RECT 95.525 91.555 97.360 92.235 ;
        RECT 97.555 91.555 104.865 92.235 ;
        RECT 105.020 91.555 106.855 92.235 ;
        RECT 95.525 91.325 96.455 91.555 ;
        RECT 97.555 91.325 98.905 91.555 ;
        RECT 100.440 91.335 101.350 91.555 ;
        RECT 105.925 91.325 106.855 91.555 ;
        RECT 107.175 91.425 109.005 92.235 ;
        RECT 109.015 91.325 112.225 92.235 ;
        RECT 112.235 91.325 115.445 92.235 ;
        RECT 116.385 91.365 116.815 92.150 ;
        RECT 116.835 91.325 120.310 92.235 ;
        RECT 120.975 91.555 128.285 92.235 ;
        RECT 128.480 91.555 130.315 92.235 ;
        RECT 124.490 91.335 125.400 91.555 ;
        RECT 126.935 91.325 128.285 91.555 ;
        RECT 129.385 91.325 130.315 91.555 ;
        RECT 130.635 91.425 134.305 92.235 ;
        RECT 134.315 91.425 135.685 92.235 ;
        RECT 135.695 91.555 137.525 92.235 ;
        RECT 136.180 91.325 137.525 91.555 ;
        RECT 137.535 91.425 138.905 92.235 ;
      LAYER nwell ;
        RECT 13.140 88.205 139.100 91.035 ;
      LAYER pwell ;
        RECT 13.335 87.005 14.705 87.815 ;
        RECT 14.715 87.005 20.225 87.815 ;
        RECT 20.235 87.005 25.745 87.815 ;
        RECT 26.225 87.090 26.655 87.875 ;
        RECT 26.675 87.005 32.185 87.815 ;
        RECT 32.195 87.005 37.705 87.815 ;
        RECT 37.715 87.005 39.085 87.815 ;
        RECT 39.105 87.090 39.535 87.875 ;
        RECT 39.555 87.005 45.065 87.815 ;
        RECT 45.075 87.005 50.585 87.815 ;
        RECT 50.595 87.005 51.965 87.815 ;
        RECT 51.985 87.090 52.415 87.875 ;
        RECT 52.435 87.005 57.945 87.815 ;
        RECT 57.955 87.005 59.785 87.815 ;
        RECT 60.280 87.685 61.625 87.915 ;
        RECT 59.795 87.005 61.625 87.685 ;
        RECT 61.635 87.005 64.385 87.815 ;
        RECT 64.865 87.090 65.295 87.875 ;
        RECT 66.235 87.685 67.580 87.915 ;
        RECT 66.235 87.005 68.065 87.685 ;
        RECT 68.075 87.005 69.445 87.815 ;
        RECT 70.115 87.685 74.045 87.915 ;
        RECT 69.630 87.005 74.045 87.685 ;
        RECT 74.055 87.685 75.400 87.915 ;
        RECT 75.895 87.685 77.240 87.915 ;
        RECT 74.055 87.005 75.885 87.685 ;
        RECT 75.895 87.005 77.725 87.685 ;
        RECT 77.745 87.090 78.175 87.875 ;
        RECT 79.115 87.685 80.460 87.915 ;
        RECT 79.115 87.005 80.945 87.685 ;
        RECT 80.955 87.005 82.325 87.815 ;
        RECT 82.335 87.685 83.680 87.915 ;
        RECT 82.335 87.005 84.165 87.685 ;
        RECT 84.175 87.005 85.545 87.815 ;
        RECT 85.555 87.685 86.900 87.915 ;
        RECT 85.555 87.005 87.385 87.685 ;
        RECT 87.395 87.005 88.765 87.815 ;
        RECT 88.775 87.685 90.120 87.915 ;
        RECT 88.775 87.005 90.605 87.685 ;
        RECT 90.625 87.090 91.055 87.875 ;
        RECT 91.995 87.685 93.340 87.915 ;
        RECT 91.995 87.005 93.825 87.685 ;
        RECT 93.835 87.005 95.205 87.815 ;
        RECT 95.215 87.685 96.560 87.915 ;
        RECT 97.975 87.685 99.320 87.915 ;
        RECT 100.865 87.685 101.795 87.915 ;
        RECT 95.215 87.005 97.045 87.685 ;
        RECT 97.975 87.005 99.805 87.685 ;
        RECT 99.960 87.005 101.795 87.685 ;
        RECT 102.115 87.005 103.485 87.815 ;
        RECT 103.505 87.090 103.935 87.875 ;
        RECT 103.955 87.685 105.300 87.915 ;
        RECT 105.795 87.685 107.140 87.915 ;
        RECT 108.095 87.685 109.440 87.915 ;
        RECT 103.955 87.005 105.785 87.685 ;
        RECT 105.795 87.005 107.625 87.685 ;
        RECT 108.095 87.005 109.925 87.685 ;
        RECT 109.935 87.005 111.305 87.815 ;
        RECT 111.800 87.685 113.145 87.915 ;
        RECT 114.665 87.685 115.595 87.915 ;
        RECT 111.315 87.005 113.145 87.685 ;
        RECT 113.760 87.005 115.595 87.685 ;
        RECT 116.385 87.090 116.815 87.875 ;
        RECT 117.320 87.685 118.665 87.915 ;
        RECT 119.160 87.685 120.505 87.915 ;
        RECT 116.835 87.005 118.665 87.685 ;
        RECT 118.675 87.005 120.505 87.685 ;
        RECT 120.975 87.685 122.320 87.915 ;
        RECT 120.975 87.005 122.805 87.685 ;
        RECT 122.815 87.005 124.185 87.815 ;
        RECT 124.680 87.685 126.025 87.915 ;
        RECT 124.195 87.005 126.025 87.685 ;
        RECT 126.035 87.005 127.405 87.815 ;
        RECT 127.900 87.685 129.245 87.915 ;
        RECT 127.415 87.005 129.245 87.685 ;
        RECT 129.265 87.090 129.695 87.875 ;
        RECT 130.635 87.685 131.980 87.915 ;
        RECT 130.635 87.005 132.465 87.685 ;
        RECT 132.475 87.005 136.145 87.815 ;
        RECT 136.155 87.005 137.525 87.815 ;
        RECT 137.535 87.005 138.905 87.815 ;
        RECT 13.475 86.815 13.645 87.005 ;
        RECT 14.855 86.815 15.025 87.005 ;
        RECT 20.375 86.815 20.545 87.005 ;
        RECT 25.890 86.845 26.010 86.955 ;
        RECT 26.815 86.815 26.985 87.005 ;
        RECT 32.335 86.815 32.505 87.005 ;
        RECT 37.855 86.815 38.025 87.005 ;
        RECT 39.695 86.815 39.865 87.005 ;
        RECT 45.215 86.815 45.385 87.005 ;
        RECT 50.735 86.815 50.905 87.005 ;
        RECT 52.575 86.815 52.745 87.005 ;
        RECT 58.095 86.815 58.265 87.005 ;
        RECT 59.935 86.815 60.105 87.005 ;
        RECT 61.775 86.815 61.945 87.005 ;
        RECT 64.530 86.845 64.650 86.955 ;
        RECT 65.465 86.850 65.625 86.960 ;
        RECT 67.755 86.815 67.925 87.005 ;
        RECT 68.215 86.815 68.385 87.005 ;
        RECT 69.630 86.985 69.740 87.005 ;
        RECT 69.570 86.815 69.740 86.985 ;
        RECT 75.575 86.815 75.745 87.005 ;
        RECT 77.415 86.815 77.585 87.005 ;
        RECT 78.345 86.850 78.505 86.960 ;
        RECT 80.635 86.815 80.805 87.005 ;
        RECT 81.095 86.815 81.265 87.005 ;
        RECT 83.855 86.815 84.025 87.005 ;
        RECT 84.315 86.815 84.485 87.005 ;
        RECT 87.075 86.815 87.245 87.005 ;
        RECT 87.535 86.815 87.705 87.005 ;
        RECT 90.295 86.815 90.465 87.005 ;
        RECT 91.225 86.850 91.385 86.960 ;
        RECT 93.515 86.815 93.685 87.005 ;
        RECT 93.975 86.815 94.145 87.005 ;
        RECT 96.735 86.815 96.905 87.005 ;
        RECT 97.205 86.850 97.365 86.960 ;
        RECT 99.495 86.815 99.665 87.005 ;
        RECT 99.960 86.985 100.125 87.005 ;
        RECT 99.955 86.815 100.125 86.985 ;
        RECT 102.255 86.815 102.425 87.005 ;
        RECT 105.475 86.815 105.645 87.005 ;
        RECT 107.315 86.815 107.485 87.005 ;
        RECT 107.770 86.845 107.890 86.955 ;
        RECT 109.615 86.815 109.785 87.005 ;
        RECT 110.075 86.815 110.245 87.005 ;
        RECT 111.455 86.815 111.625 87.005 ;
        RECT 113.760 86.985 113.925 87.005 ;
        RECT 113.290 86.845 113.410 86.955 ;
        RECT 113.755 86.815 113.925 86.985 ;
        RECT 116.050 86.845 116.170 86.955 ;
        RECT 116.975 86.815 117.145 87.005 ;
        RECT 118.815 86.815 118.985 87.005 ;
        RECT 120.650 86.845 120.770 86.955 ;
        RECT 122.495 86.815 122.665 87.005 ;
        RECT 122.955 86.815 123.125 87.005 ;
        RECT 124.335 86.815 124.505 87.005 ;
        RECT 126.175 86.815 126.345 87.005 ;
        RECT 127.555 86.815 127.725 87.005 ;
        RECT 129.865 86.850 130.025 86.960 ;
        RECT 132.155 86.815 132.325 87.005 ;
        RECT 132.615 86.815 132.785 87.005 ;
        RECT 136.295 86.815 136.465 87.005 ;
        RECT 138.595 86.815 138.765 87.005 ;
      LAYER nwell ;
        RECT 12.730 50.225 48.990 51.830 ;
      LAYER pwell ;
        RECT 12.925 49.025 14.295 49.835 ;
        RECT 14.305 49.025 19.815 49.835 ;
        RECT 21.230 49.705 22.575 49.935 ;
        RECT 20.745 49.025 22.575 49.705 ;
        RECT 22.715 49.025 25.715 49.935 ;
        RECT 25.815 49.110 26.245 49.895 ;
        RECT 29.840 49.705 30.760 49.935 ;
        RECT 27.295 49.025 30.760 49.705 ;
        RECT 31.785 49.705 33.130 49.935 ;
        RECT 36.280 49.705 37.200 49.935 ;
        RECT 31.785 49.025 33.615 49.705 ;
        RECT 33.735 49.025 37.200 49.705 ;
        RECT 37.305 49.025 38.675 49.805 ;
        RECT 38.695 49.110 39.125 49.895 ;
        RECT 40.065 49.705 41.410 49.935 ;
        RECT 40.065 49.025 41.895 49.705 ;
        RECT 41.905 49.025 43.275 49.835 ;
        RECT 43.285 49.025 44.655 49.805 ;
        RECT 44.665 49.025 46.035 49.805 ;
        RECT 46.045 49.025 47.415 49.805 ;
        RECT 47.425 49.025 48.795 49.835 ;
        RECT 13.065 48.815 13.235 49.025 ;
        RECT 14.445 48.815 14.615 49.025 ;
        RECT 18.120 48.865 18.240 48.975 ;
        RECT 19.975 48.870 20.135 48.980 ;
        RECT 20.885 48.835 21.055 49.025 ;
        RECT 25.485 48.815 25.655 49.025 ;
        RECT 25.945 48.815 26.115 49.005 ;
        RECT 26.415 48.870 26.575 48.980 ;
        RECT 27.325 48.835 27.495 49.025 ;
        RECT 31.015 48.870 31.175 48.980 ;
        RECT 33.305 48.835 33.475 49.025 ;
        RECT 33.765 48.835 33.935 49.025 ;
        RECT 37.455 49.005 37.625 49.025 ;
        RECT 35.145 48.835 35.315 49.005 ;
        RECT 35.145 48.815 35.310 48.835 ;
        RECT 35.605 48.815 35.775 49.005 ;
        RECT 37.445 48.835 37.625 49.005 ;
        RECT 37.445 48.815 37.615 48.835 ;
        RECT 39.285 48.815 39.455 49.005 ;
        RECT 41.585 48.835 41.755 49.025 ;
        RECT 42.045 48.835 42.215 49.025 ;
        RECT 42.505 48.815 42.675 49.005 ;
        RECT 44.345 48.835 44.515 49.025 ;
        RECT 45.725 48.835 45.895 49.025 ;
        RECT 47.095 48.815 47.265 49.025 ;
        RECT 48.485 48.815 48.655 49.025 ;
        RECT 12.925 48.005 14.295 48.815 ;
        RECT 14.305 48.005 17.975 48.815 ;
        RECT 18.485 48.135 25.795 48.815 ;
        RECT 25.805 48.135 33.115 48.815 ;
        RECT 18.485 47.905 19.835 48.135 ;
        RECT 21.370 47.915 22.280 48.135 ;
        RECT 29.320 47.915 30.230 48.135 ;
        RECT 31.765 47.905 33.115 48.135 ;
        RECT 33.475 48.135 35.310 48.815 ;
        RECT 35.465 48.135 37.295 48.815 ;
        RECT 33.475 47.905 34.405 48.135 ;
        RECT 35.950 47.905 37.295 48.135 ;
        RECT 37.315 47.905 38.665 48.815 ;
        RECT 38.695 47.945 39.125 48.730 ;
        RECT 39.225 47.905 42.225 48.815 ;
        RECT 42.475 48.135 45.940 48.815 ;
        RECT 45.020 47.905 45.940 48.135 ;
        RECT 46.045 48.035 47.415 48.815 ;
        RECT 47.425 48.005 48.795 48.815 ;
      LAYER nwell ;
        RECT 12.730 44.785 48.990 47.615 ;
      LAYER pwell ;
        RECT 12.925 43.585 14.295 44.395 ;
        RECT 17.820 44.265 18.730 44.485 ;
        RECT 20.265 44.265 21.615 44.495 ;
        RECT 14.305 43.585 21.615 44.265 ;
        RECT 21.760 44.265 22.680 44.495 ;
        RECT 21.760 43.585 25.225 44.265 ;
        RECT 25.815 43.670 26.245 44.455 ;
        RECT 26.265 44.265 27.195 44.495 ;
        RECT 31.915 44.265 32.845 44.495 ;
        RECT 26.265 43.585 30.165 44.265 ;
        RECT 31.010 43.585 32.845 44.265 ;
        RECT 33.175 43.585 34.525 44.495 ;
        RECT 38.060 44.265 38.970 44.485 ;
        RECT 40.505 44.265 41.855 44.495 ;
        RECT 43.415 44.265 44.345 44.495 ;
        RECT 34.545 43.585 41.855 44.265 ;
        RECT 42.510 43.585 44.345 44.265 ;
        RECT 44.665 43.585 46.035 44.365 ;
        RECT 46.045 43.585 47.415 44.365 ;
        RECT 47.425 43.585 48.795 44.395 ;
        RECT 13.065 43.375 13.235 43.585 ;
        RECT 14.445 43.395 14.615 43.585 ;
        RECT 15.825 43.375 15.995 43.565 ;
        RECT 16.560 43.375 16.730 43.565 ;
        RECT 20.425 43.375 20.595 43.565 ;
        RECT 25.025 43.395 25.195 43.585 ;
        RECT 25.480 43.425 25.600 43.535 ;
        RECT 26.680 43.395 26.850 43.585 ;
        RECT 31.010 43.565 31.175 43.585 ;
        RECT 30.545 43.535 30.715 43.565 ;
        RECT 30.540 43.425 30.715 43.535 ;
        RECT 30.545 43.375 30.715 43.425 ;
        RECT 31.005 43.395 31.175 43.565 ;
        RECT 34.225 43.375 34.395 43.585 ;
        RECT 34.685 43.375 34.855 43.585 ;
        RECT 42.510 43.565 42.675 43.585 ;
        RECT 12.925 42.565 14.295 43.375 ;
        RECT 14.305 42.695 16.135 43.375 ;
        RECT 16.145 42.695 20.045 43.375 ;
        RECT 14.305 42.465 15.650 42.695 ;
        RECT 16.145 42.465 17.075 42.695 ;
        RECT 20.285 42.565 21.655 43.375 ;
        RECT 21.750 42.695 30.855 43.375 ;
        RECT 30.960 42.695 34.425 43.375 ;
        RECT 30.960 42.465 31.880 42.695 ;
        RECT 34.545 42.565 35.915 43.375 ;
        RECT 36.070 43.345 36.240 43.565 ;
        RECT 39.285 43.375 39.455 43.565 ;
        RECT 42.040 43.425 42.160 43.535 ;
        RECT 42.505 43.395 42.675 43.565 ;
        RECT 42.965 43.375 43.135 43.565 ;
        RECT 44.805 43.395 44.975 43.585 ;
        RECT 46.655 43.420 46.815 43.530 ;
        RECT 47.095 43.395 47.265 43.585 ;
        RECT 48.485 43.375 48.655 43.585 ;
        RECT 37.730 43.345 38.675 43.375 ;
        RECT 35.925 42.665 38.675 43.345 ;
        RECT 37.730 42.465 38.675 42.665 ;
        RECT 38.695 42.505 39.125 43.290 ;
        RECT 39.225 42.465 42.675 43.375 ;
        RECT 42.905 42.465 46.355 43.375 ;
        RECT 47.425 42.565 48.795 43.375 ;
      LAYER nwell ;
        RECT 12.730 39.345 48.990 42.175 ;
      LAYER pwell ;
        RECT 12.925 38.145 14.295 38.955 ;
        RECT 14.305 38.825 15.235 39.055 ;
        RECT 21.960 38.825 22.870 39.045 ;
        RECT 24.405 38.825 25.755 39.055 ;
        RECT 14.305 38.145 18.205 38.825 ;
        RECT 18.445 38.145 25.755 38.825 ;
        RECT 25.815 38.230 26.245 39.015 ;
        RECT 29.780 38.825 30.690 39.045 ;
        RECT 32.225 38.825 33.575 39.055 ;
        RECT 26.265 38.145 33.575 38.825 ;
        RECT 34.085 38.825 35.450 39.055 ;
        RECT 34.085 38.145 37.295 38.825 ;
        RECT 38.305 38.145 41.305 39.055 ;
        RECT 41.445 38.145 42.795 39.055 ;
        RECT 43.365 38.145 46.815 39.055 ;
        RECT 47.425 38.145 48.795 38.955 ;
        RECT 13.065 37.935 13.235 38.145 ;
        RECT 14.720 37.955 14.890 38.145 ;
        RECT 18.585 37.955 18.755 38.145 ;
        RECT 21.345 37.935 21.515 38.125 ;
        RECT 21.805 37.935 21.975 38.125 ;
        RECT 24.560 37.985 24.680 38.095 ;
        RECT 25.025 37.935 25.195 38.125 ;
        RECT 26.405 37.955 26.575 38.145 ;
        RECT 33.760 37.985 33.880 38.095 ;
        RECT 36.980 37.955 37.150 38.145 ;
        RECT 37.445 37.935 37.615 38.125 ;
        RECT 37.915 37.980 38.075 38.090 ;
        RECT 38.365 37.955 38.535 38.145 ;
        RECT 41.590 38.125 41.760 38.145 ;
        RECT 12.925 37.125 14.295 37.935 ;
        RECT 14.345 37.255 21.655 37.935 ;
        RECT 14.345 37.025 15.695 37.255 ;
        RECT 17.230 37.035 18.140 37.255 ;
        RECT 21.665 37.125 24.415 37.935 ;
        RECT 24.885 37.255 33.990 37.935 ;
        RECT 34.180 37.255 37.645 37.935 ;
        RECT 39.280 37.905 39.450 38.125 ;
        RECT 41.585 37.955 41.760 38.125 ;
        RECT 42.960 37.985 43.080 38.095 ;
        RECT 43.425 37.955 43.595 38.145 ;
        RECT 44.340 37.985 44.460 38.095 ;
        RECT 41.585 37.935 41.755 37.955 ;
        RECT 45.720 37.935 45.890 38.125 ;
        RECT 47.105 38.095 47.275 38.125 ;
        RECT 47.100 37.985 47.275 38.095 ;
        RECT 47.105 37.935 47.275 37.985 ;
        RECT 48.485 37.935 48.655 38.145 ;
        RECT 40.480 37.905 41.435 37.935 ;
        RECT 34.180 37.025 35.100 37.255 ;
        RECT 38.695 37.065 39.125 37.850 ;
        RECT 39.155 37.225 41.435 37.905 ;
        RECT 40.480 37.025 41.435 37.225 ;
        RECT 41.445 37.125 44.195 37.935 ;
        RECT 44.685 37.025 46.035 37.935 ;
        RECT 46.045 37.155 47.415 37.935 ;
        RECT 47.425 37.125 48.795 37.935 ;
      LAYER nwell ;
        RECT 12.730 33.905 48.990 36.735 ;
      LAYER pwell ;
        RECT 12.925 32.705 14.295 33.515 ;
        RECT 14.305 32.705 15.675 33.515 ;
        RECT 18.340 33.385 19.260 33.615 ;
        RECT 15.795 32.705 19.260 33.385 ;
        RECT 19.460 33.385 20.380 33.615 ;
        RECT 19.460 32.705 22.925 33.385 ;
        RECT 23.045 32.705 25.795 33.515 ;
        RECT 25.815 32.790 26.245 33.575 ;
        RECT 26.285 32.705 27.635 33.615 ;
        RECT 27.715 32.705 31.775 33.615 ;
        RECT 31.880 33.385 32.800 33.615 ;
        RECT 31.880 32.705 35.345 33.385 ;
        RECT 35.465 32.705 36.835 33.515 ;
        RECT 36.845 33.415 37.795 33.615 ;
        RECT 36.845 32.735 40.515 33.415 ;
        RECT 36.845 32.705 37.795 32.735 ;
        RECT 13.065 32.495 13.235 32.705 ;
        RECT 14.445 32.515 14.615 32.705 ;
        RECT 15.825 32.495 15.995 32.705 ;
        RECT 16.280 32.545 16.400 32.655 ;
        RECT 17.020 32.495 17.190 32.685 ;
        RECT 20.885 32.495 21.055 32.685 ;
        RECT 22.725 32.515 22.895 32.705 ;
        RECT 23.185 32.515 23.355 32.705 ;
        RECT 27.320 32.515 27.490 32.705 ;
        RECT 28.520 32.495 28.690 32.685 ;
        RECT 31.465 32.515 31.635 32.705 ;
        RECT 35.145 32.515 35.315 32.705 ;
        RECT 35.605 32.495 35.775 32.705 ;
        RECT 36.065 32.495 36.235 32.685 ;
        RECT 40.200 32.515 40.370 32.735 ;
        RECT 40.525 32.705 41.875 33.615 ;
        RECT 41.905 32.705 43.275 33.485 ;
        RECT 43.425 32.705 46.875 33.615 ;
        RECT 47.425 32.705 48.795 33.515 ;
        RECT 40.670 32.515 40.840 32.705 ;
        RECT 42.055 32.685 42.225 32.705 ;
        RECT 42.040 32.515 42.225 32.685 ;
        RECT 42.515 32.540 42.675 32.650 ;
        RECT 42.040 32.495 42.210 32.515 ;
        RECT 46.645 32.495 46.815 32.705 ;
        RECT 47.100 32.545 47.220 32.655 ;
        RECT 48.485 32.495 48.655 32.705 ;
        RECT 12.925 31.685 14.295 32.495 ;
        RECT 14.305 31.815 16.135 32.495 ;
        RECT 16.605 31.815 20.505 32.495 ;
        RECT 20.745 31.815 28.055 32.495 ;
        RECT 14.305 31.585 15.650 31.815 ;
        RECT 16.605 31.585 17.535 31.815 ;
        RECT 24.260 31.595 25.170 31.815 ;
        RECT 26.705 31.585 28.055 31.815 ;
        RECT 28.105 31.815 32.005 32.495 ;
        RECT 32.340 31.815 35.805 32.495 ;
        RECT 28.105 31.585 29.035 31.815 ;
        RECT 32.340 31.585 33.260 31.815 ;
        RECT 35.925 31.685 38.675 32.495 ;
        RECT 38.695 31.625 39.125 32.410 ;
        RECT 39.435 31.585 42.355 32.495 ;
        RECT 43.425 31.585 46.875 32.495 ;
        RECT 47.425 31.685 48.795 32.495 ;
      LAYER nwell ;
        RECT 12.730 28.465 48.990 31.295 ;
      LAYER pwell ;
        RECT 12.925 27.265 14.295 28.075 ;
        RECT 17.820 27.945 18.730 28.165 ;
        RECT 20.265 27.945 21.615 28.175 ;
        RECT 14.305 27.265 21.615 27.945 ;
        RECT 21.665 27.265 25.335 28.075 ;
        RECT 25.815 27.350 26.245 28.135 ;
        RECT 29.780 27.945 30.690 28.165 ;
        RECT 32.225 27.945 33.575 28.175 ;
        RECT 35.470 27.945 36.835 28.175 ;
        RECT 26.265 27.265 33.575 27.945 ;
        RECT 33.625 27.265 36.835 27.945 ;
        RECT 36.845 27.265 39.595 28.075 ;
        RECT 42.720 27.945 43.640 28.175 ;
        RECT 40.175 27.265 43.640 27.945 ;
        RECT 43.825 27.265 46.825 28.175 ;
        RECT 47.425 27.265 48.795 28.075 ;
        RECT 13.065 27.055 13.235 27.265 ;
        RECT 14.445 27.075 14.615 27.265 ;
        RECT 15.825 27.055 15.995 27.245 ;
        RECT 16.295 27.100 16.455 27.210 ;
        RECT 17.205 27.055 17.375 27.245 ;
        RECT 20.895 27.100 21.055 27.210 ;
        RECT 21.805 27.055 21.975 27.265 ;
        RECT 25.480 27.105 25.600 27.215 ;
        RECT 26.405 27.075 26.575 27.265 ;
        RECT 28.890 27.055 29.060 27.245 ;
        RECT 29.625 27.055 29.795 27.245 ;
        RECT 31.465 27.055 31.635 27.245 ;
        RECT 33.770 27.075 33.940 27.265 ;
        RECT 36.985 27.075 37.155 27.265 ;
        RECT 39.560 27.055 39.730 27.245 ;
        RECT 39.740 27.105 39.860 27.215 ;
        RECT 40.205 27.075 40.375 27.265 ;
        RECT 43.425 27.055 43.595 27.245 ;
        RECT 43.885 27.075 44.055 27.265 ;
        RECT 12.925 26.245 14.295 27.055 ;
        RECT 14.305 26.375 16.135 27.055 ;
        RECT 17.175 26.375 20.640 27.055 ;
        RECT 21.775 26.375 25.240 27.055 ;
        RECT 25.575 26.375 29.475 27.055 ;
        RECT 14.305 26.145 15.650 26.375 ;
        RECT 19.720 26.145 20.640 26.375 ;
        RECT 24.320 26.145 25.240 26.375 ;
        RECT 28.545 26.145 29.475 26.375 ;
        RECT 29.485 26.245 31.315 27.055 ;
        RECT 31.325 26.375 38.635 27.055 ;
        RECT 34.840 26.155 35.750 26.375 ;
        RECT 37.285 26.145 38.635 26.375 ;
        RECT 38.695 26.185 39.125 26.970 ;
        RECT 39.145 26.375 43.045 27.055 ;
        RECT 39.145 26.145 40.075 26.375 ;
        RECT 43.285 26.275 44.655 27.055 ;
        RECT 44.665 27.025 45.610 27.055 ;
        RECT 47.100 27.025 47.270 27.245 ;
        RECT 48.485 27.055 48.655 27.265 ;
        RECT 44.665 26.345 47.415 27.025 ;
        RECT 44.665 26.145 45.610 26.345 ;
        RECT 47.425 26.245 48.795 27.055 ;
      LAYER nwell ;
        RECT 12.730 23.025 48.990 25.855 ;
      LAYER pwell ;
        RECT 12.925 21.825 14.295 22.635 ;
        RECT 14.345 22.505 15.695 22.735 ;
        RECT 17.230 22.505 18.140 22.725 ;
        RECT 14.345 21.825 21.655 22.505 ;
        RECT 21.665 21.825 25.335 22.635 ;
        RECT 25.815 21.910 26.245 22.695 ;
        RECT 26.265 21.825 35.370 22.505 ;
        RECT 35.465 21.825 36.835 22.635 ;
        RECT 36.845 21.825 38.215 22.605 ;
        RECT 38.225 21.825 39.595 22.605 ;
        RECT 39.605 21.825 40.975 22.605 ;
        RECT 40.985 21.825 42.355 22.605 ;
        RECT 42.385 21.825 43.735 22.735 ;
        RECT 43.825 21.825 47.275 22.735 ;
        RECT 47.425 21.825 48.795 22.635 ;
        RECT 13.065 21.615 13.235 21.825 ;
        RECT 15.825 21.615 15.995 21.805 ;
        RECT 16.295 21.660 16.455 21.770 ;
        RECT 17.480 21.615 17.650 21.805 ;
        RECT 21.345 21.615 21.515 21.825 ;
        RECT 21.805 21.635 21.975 21.825 ;
        RECT 25.025 21.615 25.195 21.805 ;
        RECT 25.480 21.665 25.600 21.775 ;
        RECT 26.405 21.635 26.575 21.825 ;
        RECT 33.305 21.615 33.475 21.805 ;
        RECT 34.040 21.615 34.210 21.805 ;
        RECT 35.605 21.635 35.775 21.825 ;
        RECT 36.985 21.635 37.155 21.825 ;
        RECT 37.915 21.660 38.075 21.770 ;
        RECT 38.365 21.635 38.535 21.825 ;
        RECT 39.745 21.635 39.915 21.825 ;
        RECT 41.125 21.635 41.295 21.825 ;
        RECT 42.505 21.615 42.675 21.805 ;
        RECT 42.975 21.660 43.135 21.770 ;
        RECT 43.420 21.635 43.590 21.825 ;
        RECT 43.885 21.635 44.055 21.825 ;
        RECT 46.185 21.615 46.355 21.805 ;
        RECT 46.655 21.660 46.815 21.770 ;
        RECT 48.485 21.615 48.655 21.825 ;
        RECT 12.925 20.805 14.295 21.615 ;
        RECT 14.305 20.935 16.135 21.615 ;
        RECT 17.065 20.935 20.965 21.615 ;
        RECT 14.305 20.705 15.650 20.935 ;
        RECT 17.065 20.705 17.995 20.935 ;
        RECT 21.205 20.805 24.875 21.615 ;
        RECT 24.885 20.805 26.255 21.615 ;
        RECT 26.305 20.935 33.615 21.615 ;
        RECT 33.625 20.935 37.525 21.615 ;
        RECT 26.305 20.705 27.655 20.935 ;
        RECT 29.190 20.715 30.100 20.935 ;
        RECT 33.625 20.705 34.555 20.935 ;
        RECT 38.695 20.745 39.125 21.530 ;
        RECT 39.240 20.935 42.705 21.615 ;
        RECT 39.240 20.705 40.160 20.935 ;
        RECT 43.745 20.705 46.495 21.615 ;
        RECT 47.425 20.805 48.795 21.615 ;
      LAYER nwell ;
        RECT 12.730 17.585 48.990 20.415 ;
      LAYER pwell ;
        RECT 12.925 16.385 14.295 17.195 ;
        RECT 14.305 16.385 19.815 17.195 ;
        RECT 19.825 16.385 23.495 17.195 ;
        RECT 24.450 17.065 25.795 17.295 ;
        RECT 23.965 16.385 25.795 17.065 ;
        RECT 25.815 16.470 26.245 17.255 ;
        RECT 26.725 17.065 28.070 17.295 ;
        RECT 32.080 17.065 32.990 17.285 ;
        RECT 34.525 17.065 35.875 17.295 ;
        RECT 26.725 16.385 28.555 17.065 ;
        RECT 28.565 16.385 35.875 17.065 ;
        RECT 35.925 17.065 37.270 17.295 ;
        RECT 35.925 16.385 37.755 17.065 ;
        RECT 38.695 16.470 39.125 17.255 ;
        RECT 40.550 17.065 41.895 17.295 ;
        RECT 40.065 16.385 41.895 17.065 ;
        RECT 41.905 16.385 43.275 17.165 ;
        RECT 46.025 17.065 46.955 17.295 ;
        RECT 44.205 16.385 46.955 17.065 ;
        RECT 47.425 16.385 48.795 17.195 ;
        RECT 13.065 16.195 13.235 16.385 ;
        RECT 14.445 16.195 14.615 16.385 ;
        RECT 19.965 16.195 20.135 16.385 ;
        RECT 23.640 16.225 23.760 16.335 ;
        RECT 24.105 16.195 24.275 16.385 ;
        RECT 26.400 16.225 26.520 16.335 ;
        RECT 28.245 16.195 28.415 16.385 ;
        RECT 28.705 16.195 28.875 16.385 ;
        RECT 37.445 16.195 37.615 16.385 ;
        RECT 37.915 16.230 38.075 16.340 ;
        RECT 39.295 16.230 39.455 16.340 ;
        RECT 40.205 16.195 40.375 16.385 ;
        RECT 42.955 16.195 43.125 16.385 ;
        RECT 43.435 16.230 43.595 16.340 ;
        RECT 44.345 16.195 44.515 16.385 ;
        RECT 47.100 16.225 47.220 16.335 ;
        RECT 48.485 16.195 48.655 16.385 ;
      LAYER li1 ;
        RECT 13.330 211.935 138.910 212.105 ;
        RECT 13.415 211.185 14.625 211.935 ;
        RECT 14.795 211.390 20.140 211.935 ;
        RECT 20.315 211.390 25.660 211.935 ;
        RECT 13.415 210.645 13.935 211.185 ;
        RECT 14.105 210.475 14.625 211.015 ;
        RECT 16.380 210.560 16.720 211.390 ;
        RECT 13.415 209.385 14.625 210.475 ;
        RECT 18.200 209.820 18.550 211.070 ;
        RECT 21.900 210.560 22.240 211.390 ;
        RECT 26.295 211.210 26.585 211.935 ;
        RECT 26.755 211.390 32.100 211.935 ;
        RECT 32.275 211.390 37.620 211.935 ;
        RECT 23.720 209.820 24.070 211.070 ;
        RECT 28.340 210.560 28.680 211.390 ;
        RECT 14.795 209.385 20.140 209.820 ;
        RECT 20.315 209.385 25.660 209.820 ;
        RECT 26.295 209.385 26.585 210.550 ;
        RECT 30.160 209.820 30.510 211.070 ;
        RECT 33.860 210.560 34.200 211.390 ;
        RECT 37.795 211.185 39.005 211.935 ;
        RECT 39.175 211.210 39.465 211.935 ;
        RECT 39.635 211.390 44.980 211.935 ;
        RECT 45.155 211.390 50.500 211.935 ;
        RECT 35.680 209.820 36.030 211.070 ;
        RECT 37.795 210.645 38.315 211.185 ;
        RECT 38.485 210.475 39.005 211.015 ;
        RECT 41.220 210.560 41.560 211.390 ;
        RECT 26.755 209.385 32.100 209.820 ;
        RECT 32.275 209.385 37.620 209.820 ;
        RECT 37.795 209.385 39.005 210.475 ;
        RECT 39.175 209.385 39.465 210.550 ;
        RECT 43.040 209.820 43.390 211.070 ;
        RECT 46.740 210.560 47.080 211.390 ;
        RECT 50.675 211.185 51.885 211.935 ;
        RECT 52.055 211.210 52.345 211.935 ;
        RECT 52.515 211.390 57.860 211.935 ;
        RECT 58.035 211.390 63.380 211.935 ;
        RECT 48.560 209.820 48.910 211.070 ;
        RECT 50.675 210.645 51.195 211.185 ;
        RECT 51.365 210.475 51.885 211.015 ;
        RECT 54.100 210.560 54.440 211.390 ;
        RECT 39.635 209.385 44.980 209.820 ;
        RECT 45.155 209.385 50.500 209.820 ;
        RECT 50.675 209.385 51.885 210.475 ;
        RECT 52.055 209.385 52.345 210.550 ;
        RECT 55.920 209.820 56.270 211.070 ;
        RECT 59.620 210.560 59.960 211.390 ;
        RECT 63.555 211.185 64.765 211.935 ;
        RECT 64.935 211.210 65.225 211.935 ;
        RECT 65.395 211.390 70.740 211.935 ;
        RECT 61.440 209.820 61.790 211.070 ;
        RECT 63.555 210.645 64.075 211.185 ;
        RECT 64.245 210.475 64.765 211.015 ;
        RECT 66.980 210.560 67.320 211.390 ;
        RECT 70.915 211.165 72.585 211.935 ;
        RECT 52.515 209.385 57.860 209.820 ;
        RECT 58.035 209.385 63.380 209.820 ;
        RECT 63.555 209.385 64.765 210.475 ;
        RECT 64.935 209.385 65.225 210.550 ;
        RECT 68.800 209.820 69.150 211.070 ;
        RECT 70.915 210.645 71.665 211.165 ;
        RECT 72.760 211.095 73.020 211.935 ;
        RECT 73.195 211.190 73.450 211.765 ;
        RECT 73.620 211.555 73.950 211.935 ;
        RECT 74.165 211.385 74.335 211.765 ;
        RECT 73.620 211.215 74.335 211.385 ;
        RECT 71.835 210.475 72.585 210.995 ;
        RECT 65.395 209.385 70.740 209.820 ;
        RECT 70.915 209.385 72.585 210.475 ;
        RECT 72.760 209.385 73.020 210.535 ;
        RECT 73.195 210.460 73.365 211.190 ;
        RECT 73.620 211.025 73.790 211.215 ;
        RECT 74.595 211.165 77.185 211.935 ;
        RECT 77.815 211.210 78.105 211.935 ;
        RECT 78.275 211.390 83.620 211.935 ;
        RECT 83.795 211.390 89.140 211.935 ;
        RECT 73.535 210.695 73.790 211.025 ;
        RECT 73.620 210.485 73.790 210.695 ;
        RECT 74.070 210.665 74.425 211.035 ;
        RECT 74.595 210.645 75.805 211.165 ;
        RECT 73.195 209.555 73.450 210.460 ;
        RECT 73.620 210.315 74.335 210.485 ;
        RECT 75.975 210.475 77.185 210.995 ;
        RECT 79.860 210.560 80.200 211.390 ;
        RECT 73.620 209.385 73.950 210.145 ;
        RECT 74.165 209.555 74.335 210.315 ;
        RECT 74.595 209.385 77.185 210.475 ;
        RECT 77.815 209.385 78.105 210.550 ;
        RECT 81.680 209.820 82.030 211.070 ;
        RECT 85.380 210.560 85.720 211.390 ;
        RECT 89.315 211.185 90.525 211.935 ;
        RECT 90.695 211.210 90.985 211.935 ;
        RECT 91.155 211.390 96.500 211.935 ;
        RECT 96.675 211.390 102.020 211.935 ;
        RECT 87.200 209.820 87.550 211.070 ;
        RECT 89.315 210.645 89.835 211.185 ;
        RECT 90.005 210.475 90.525 211.015 ;
        RECT 92.740 210.560 93.080 211.390 ;
        RECT 78.275 209.385 83.620 209.820 ;
        RECT 83.795 209.385 89.140 209.820 ;
        RECT 89.315 209.385 90.525 210.475 ;
        RECT 90.695 209.385 90.985 210.550 ;
        RECT 94.560 209.820 94.910 211.070 ;
        RECT 98.260 210.560 98.600 211.390 ;
        RECT 102.195 211.185 103.405 211.935 ;
        RECT 103.575 211.210 103.865 211.935 ;
        RECT 104.035 211.390 109.380 211.935 ;
        RECT 109.555 211.390 114.900 211.935 ;
        RECT 100.080 209.820 100.430 211.070 ;
        RECT 102.195 210.645 102.715 211.185 ;
        RECT 102.885 210.475 103.405 211.015 ;
        RECT 105.620 210.560 105.960 211.390 ;
        RECT 91.155 209.385 96.500 209.820 ;
        RECT 96.675 209.385 102.020 209.820 ;
        RECT 102.195 209.385 103.405 210.475 ;
        RECT 103.575 209.385 103.865 210.550 ;
        RECT 107.440 209.820 107.790 211.070 ;
        RECT 111.140 210.560 111.480 211.390 ;
        RECT 115.075 211.185 116.285 211.935 ;
        RECT 116.455 211.210 116.745 211.935 ;
        RECT 116.915 211.390 122.260 211.935 ;
        RECT 122.435 211.390 127.780 211.935 ;
        RECT 112.960 209.820 113.310 211.070 ;
        RECT 115.075 210.645 115.595 211.185 ;
        RECT 115.765 210.475 116.285 211.015 ;
        RECT 118.500 210.560 118.840 211.390 ;
        RECT 104.035 209.385 109.380 209.820 ;
        RECT 109.555 209.385 114.900 209.820 ;
        RECT 115.075 209.385 116.285 210.475 ;
        RECT 116.455 209.385 116.745 210.550 ;
        RECT 120.320 209.820 120.670 211.070 ;
        RECT 124.020 210.560 124.360 211.390 ;
        RECT 127.955 211.185 129.165 211.935 ;
        RECT 129.335 211.210 129.625 211.935 ;
        RECT 129.795 211.390 135.140 211.935 ;
        RECT 125.840 209.820 126.190 211.070 ;
        RECT 127.955 210.645 128.475 211.185 ;
        RECT 128.645 210.475 129.165 211.015 ;
        RECT 131.380 210.560 131.720 211.390 ;
        RECT 135.315 211.165 136.985 211.935 ;
        RECT 137.615 211.185 138.825 211.935 ;
        RECT 116.915 209.385 122.260 209.820 ;
        RECT 122.435 209.385 127.780 209.820 ;
        RECT 127.955 209.385 129.165 210.475 ;
        RECT 129.335 209.385 129.625 210.550 ;
        RECT 133.200 209.820 133.550 211.070 ;
        RECT 135.315 210.645 136.065 211.165 ;
        RECT 136.235 210.475 136.985 210.995 ;
        RECT 129.795 209.385 135.140 209.820 ;
        RECT 135.315 209.385 136.985 210.475 ;
        RECT 137.615 210.475 138.135 211.015 ;
        RECT 138.305 210.645 138.825 211.185 ;
        RECT 137.615 209.385 138.825 210.475 ;
        RECT 13.330 209.215 138.910 209.385 ;
        RECT 13.415 208.125 14.625 209.215 ;
        RECT 14.795 208.780 20.140 209.215 ;
        RECT 20.315 208.780 25.660 209.215 ;
        RECT 13.415 207.415 13.935 207.955 ;
        RECT 14.105 207.585 14.625 208.125 ;
        RECT 13.415 206.665 14.625 207.415 ;
        RECT 16.380 207.210 16.720 208.040 ;
        RECT 18.200 207.530 18.550 208.780 ;
        RECT 21.900 207.210 22.240 208.040 ;
        RECT 23.720 207.530 24.070 208.780 ;
        RECT 26.295 208.050 26.585 209.215 ;
        RECT 26.755 208.780 32.100 209.215 ;
        RECT 32.275 208.780 37.620 209.215 ;
        RECT 37.795 208.780 43.140 209.215 ;
        RECT 43.315 208.780 48.660 209.215 ;
        RECT 14.795 206.665 20.140 207.210 ;
        RECT 20.315 206.665 25.660 207.210 ;
        RECT 26.295 206.665 26.585 207.390 ;
        RECT 28.340 207.210 28.680 208.040 ;
        RECT 30.160 207.530 30.510 208.780 ;
        RECT 33.860 207.210 34.200 208.040 ;
        RECT 35.680 207.530 36.030 208.780 ;
        RECT 39.380 207.210 39.720 208.040 ;
        RECT 41.200 207.530 41.550 208.780 ;
        RECT 44.900 207.210 45.240 208.040 ;
        RECT 46.720 207.530 47.070 208.780 ;
        RECT 48.835 208.125 51.425 209.215 ;
        RECT 48.835 207.435 50.045 207.955 ;
        RECT 50.215 207.605 51.425 208.125 ;
        RECT 52.055 208.050 52.345 209.215 ;
        RECT 52.515 208.780 57.860 209.215 ;
        RECT 58.035 208.780 63.380 209.215 ;
        RECT 63.555 208.780 68.900 209.215 ;
        RECT 69.075 208.780 74.420 209.215 ;
        RECT 26.755 206.665 32.100 207.210 ;
        RECT 32.275 206.665 37.620 207.210 ;
        RECT 37.795 206.665 43.140 207.210 ;
        RECT 43.315 206.665 48.660 207.210 ;
        RECT 48.835 206.665 51.425 207.435 ;
        RECT 52.055 206.665 52.345 207.390 ;
        RECT 54.100 207.210 54.440 208.040 ;
        RECT 55.920 207.530 56.270 208.780 ;
        RECT 59.620 207.210 59.960 208.040 ;
        RECT 61.440 207.530 61.790 208.780 ;
        RECT 65.140 207.210 65.480 208.040 ;
        RECT 66.960 207.530 67.310 208.780 ;
        RECT 70.660 207.210 71.000 208.040 ;
        RECT 72.480 207.530 72.830 208.780 ;
        RECT 74.595 208.125 77.185 209.215 ;
        RECT 74.595 207.435 75.805 207.955 ;
        RECT 75.975 207.605 77.185 208.125 ;
        RECT 77.815 208.050 78.105 209.215 ;
        RECT 78.275 208.780 83.620 209.215 ;
        RECT 83.795 208.780 89.140 209.215 ;
        RECT 89.315 208.780 94.660 209.215 ;
        RECT 94.835 208.780 100.180 209.215 ;
        RECT 52.515 206.665 57.860 207.210 ;
        RECT 58.035 206.665 63.380 207.210 ;
        RECT 63.555 206.665 68.900 207.210 ;
        RECT 69.075 206.665 74.420 207.210 ;
        RECT 74.595 206.665 77.185 207.435 ;
        RECT 77.815 206.665 78.105 207.390 ;
        RECT 79.860 207.210 80.200 208.040 ;
        RECT 81.680 207.530 82.030 208.780 ;
        RECT 85.380 207.210 85.720 208.040 ;
        RECT 87.200 207.530 87.550 208.780 ;
        RECT 90.900 207.210 91.240 208.040 ;
        RECT 92.720 207.530 93.070 208.780 ;
        RECT 96.420 207.210 96.760 208.040 ;
        RECT 98.240 207.530 98.590 208.780 ;
        RECT 100.355 208.125 102.945 209.215 ;
        RECT 100.355 207.435 101.565 207.955 ;
        RECT 101.735 207.605 102.945 208.125 ;
        RECT 103.575 208.050 103.865 209.215 ;
        RECT 104.035 208.780 109.380 209.215 ;
        RECT 109.555 208.780 114.900 209.215 ;
        RECT 115.075 208.780 120.420 209.215 ;
        RECT 120.595 208.780 125.940 209.215 ;
        RECT 78.275 206.665 83.620 207.210 ;
        RECT 83.795 206.665 89.140 207.210 ;
        RECT 89.315 206.665 94.660 207.210 ;
        RECT 94.835 206.665 100.180 207.210 ;
        RECT 100.355 206.665 102.945 207.435 ;
        RECT 103.575 206.665 103.865 207.390 ;
        RECT 105.620 207.210 105.960 208.040 ;
        RECT 107.440 207.530 107.790 208.780 ;
        RECT 111.140 207.210 111.480 208.040 ;
        RECT 112.960 207.530 113.310 208.780 ;
        RECT 116.660 207.210 117.000 208.040 ;
        RECT 118.480 207.530 118.830 208.780 ;
        RECT 122.180 207.210 122.520 208.040 ;
        RECT 124.000 207.530 124.350 208.780 ;
        RECT 126.115 208.125 128.705 209.215 ;
        RECT 126.115 207.435 127.325 207.955 ;
        RECT 127.495 207.605 128.705 208.125 ;
        RECT 129.335 208.050 129.625 209.215 ;
        RECT 129.795 208.780 135.140 209.215 ;
        RECT 104.035 206.665 109.380 207.210 ;
        RECT 109.555 206.665 114.900 207.210 ;
        RECT 115.075 206.665 120.420 207.210 ;
        RECT 120.595 206.665 125.940 207.210 ;
        RECT 126.115 206.665 128.705 207.435 ;
        RECT 129.335 206.665 129.625 207.390 ;
        RECT 131.380 207.210 131.720 208.040 ;
        RECT 133.200 207.530 133.550 208.780 ;
        RECT 135.315 208.125 136.985 209.215 ;
        RECT 135.315 207.435 136.065 207.955 ;
        RECT 136.235 207.605 136.985 208.125 ;
        RECT 137.615 208.125 138.825 209.215 ;
        RECT 137.615 207.585 138.135 208.125 ;
        RECT 129.795 206.665 135.140 207.210 ;
        RECT 135.315 206.665 136.985 207.435 ;
        RECT 138.305 207.415 138.825 207.955 ;
        RECT 137.615 206.665 138.825 207.415 ;
        RECT 13.330 206.495 138.910 206.665 ;
        RECT 13.415 205.745 14.625 206.495 ;
        RECT 14.795 205.950 20.140 206.495 ;
        RECT 20.315 205.950 25.660 206.495 ;
        RECT 25.835 205.950 31.180 206.495 ;
        RECT 31.355 205.950 36.700 206.495 ;
        RECT 13.415 205.205 13.935 205.745 ;
        RECT 14.105 205.035 14.625 205.575 ;
        RECT 16.380 205.120 16.720 205.950 ;
        RECT 13.415 203.945 14.625 205.035 ;
        RECT 18.200 204.380 18.550 205.630 ;
        RECT 21.900 205.120 22.240 205.950 ;
        RECT 23.720 204.380 24.070 205.630 ;
        RECT 27.420 205.120 27.760 205.950 ;
        RECT 29.240 204.380 29.590 205.630 ;
        RECT 32.940 205.120 33.280 205.950 ;
        RECT 36.875 205.725 38.545 206.495 ;
        RECT 39.175 205.770 39.465 206.495 ;
        RECT 39.635 205.950 44.980 206.495 ;
        RECT 45.155 205.950 50.500 206.495 ;
        RECT 50.675 205.950 56.020 206.495 ;
        RECT 56.195 205.950 61.540 206.495 ;
        RECT 34.760 204.380 35.110 205.630 ;
        RECT 36.875 205.205 37.625 205.725 ;
        RECT 37.795 205.035 38.545 205.555 ;
        RECT 41.220 205.120 41.560 205.950 ;
        RECT 14.795 203.945 20.140 204.380 ;
        RECT 20.315 203.945 25.660 204.380 ;
        RECT 25.835 203.945 31.180 204.380 ;
        RECT 31.355 203.945 36.700 204.380 ;
        RECT 36.875 203.945 38.545 205.035 ;
        RECT 39.175 203.945 39.465 205.110 ;
        RECT 43.040 204.380 43.390 205.630 ;
        RECT 46.740 205.120 47.080 205.950 ;
        RECT 48.560 204.380 48.910 205.630 ;
        RECT 52.260 205.120 52.600 205.950 ;
        RECT 54.080 204.380 54.430 205.630 ;
        RECT 57.780 205.120 58.120 205.950 ;
        RECT 61.715 205.725 64.305 206.495 ;
        RECT 64.935 205.770 65.225 206.495 ;
        RECT 65.395 205.950 70.740 206.495 ;
        RECT 70.915 205.950 76.260 206.495 ;
        RECT 76.435 205.950 81.780 206.495 ;
        RECT 81.955 205.950 87.300 206.495 ;
        RECT 59.600 204.380 59.950 205.630 ;
        RECT 61.715 205.205 62.925 205.725 ;
        RECT 63.095 205.035 64.305 205.555 ;
        RECT 66.980 205.120 67.320 205.950 ;
        RECT 39.635 203.945 44.980 204.380 ;
        RECT 45.155 203.945 50.500 204.380 ;
        RECT 50.675 203.945 56.020 204.380 ;
        RECT 56.195 203.945 61.540 204.380 ;
        RECT 61.715 203.945 64.305 205.035 ;
        RECT 64.935 203.945 65.225 205.110 ;
        RECT 68.800 204.380 69.150 205.630 ;
        RECT 72.500 205.120 72.840 205.950 ;
        RECT 74.320 204.380 74.670 205.630 ;
        RECT 78.020 205.120 78.360 205.950 ;
        RECT 79.840 204.380 80.190 205.630 ;
        RECT 83.540 205.120 83.880 205.950 ;
        RECT 87.475 205.725 90.065 206.495 ;
        RECT 90.695 205.770 90.985 206.495 ;
        RECT 91.155 205.950 96.500 206.495 ;
        RECT 96.675 205.950 102.020 206.495 ;
        RECT 102.195 205.950 107.540 206.495 ;
        RECT 107.715 205.950 113.060 206.495 ;
        RECT 85.360 204.380 85.710 205.630 ;
        RECT 87.475 205.205 88.685 205.725 ;
        RECT 88.855 205.035 90.065 205.555 ;
        RECT 92.740 205.120 93.080 205.950 ;
        RECT 65.395 203.945 70.740 204.380 ;
        RECT 70.915 203.945 76.260 204.380 ;
        RECT 76.435 203.945 81.780 204.380 ;
        RECT 81.955 203.945 87.300 204.380 ;
        RECT 87.475 203.945 90.065 205.035 ;
        RECT 90.695 203.945 90.985 205.110 ;
        RECT 94.560 204.380 94.910 205.630 ;
        RECT 98.260 205.120 98.600 205.950 ;
        RECT 100.080 204.380 100.430 205.630 ;
        RECT 103.780 205.120 104.120 205.950 ;
        RECT 105.600 204.380 105.950 205.630 ;
        RECT 109.300 205.120 109.640 205.950 ;
        RECT 113.235 205.725 115.825 206.495 ;
        RECT 116.455 205.770 116.745 206.495 ;
        RECT 116.915 205.950 122.260 206.495 ;
        RECT 122.435 205.950 127.780 206.495 ;
        RECT 127.955 205.950 133.300 206.495 ;
        RECT 111.120 204.380 111.470 205.630 ;
        RECT 113.235 205.205 114.445 205.725 ;
        RECT 114.615 205.035 115.825 205.555 ;
        RECT 118.500 205.120 118.840 205.950 ;
        RECT 91.155 203.945 96.500 204.380 ;
        RECT 96.675 203.945 102.020 204.380 ;
        RECT 102.195 203.945 107.540 204.380 ;
        RECT 107.715 203.945 113.060 204.380 ;
        RECT 113.235 203.945 115.825 205.035 ;
        RECT 116.455 203.945 116.745 205.110 ;
        RECT 120.320 204.380 120.670 205.630 ;
        RECT 124.020 205.120 124.360 205.950 ;
        RECT 125.840 204.380 126.190 205.630 ;
        RECT 129.540 205.120 129.880 205.950 ;
        RECT 133.475 205.725 136.985 206.495 ;
        RECT 137.615 205.745 138.825 206.495 ;
        RECT 131.360 204.380 131.710 205.630 ;
        RECT 133.475 205.205 135.125 205.725 ;
        RECT 135.295 205.035 136.985 205.555 ;
        RECT 116.915 203.945 122.260 204.380 ;
        RECT 122.435 203.945 127.780 204.380 ;
        RECT 127.955 203.945 133.300 204.380 ;
        RECT 133.475 203.945 136.985 205.035 ;
        RECT 137.615 205.035 138.135 205.575 ;
        RECT 138.305 205.205 138.825 205.745 ;
        RECT 137.615 203.945 138.825 205.035 ;
        RECT 13.330 203.775 138.910 203.945 ;
        RECT 13.415 202.685 14.625 203.775 ;
        RECT 14.795 203.340 20.140 203.775 ;
        RECT 20.315 203.340 25.660 203.775 ;
        RECT 13.415 201.975 13.935 202.515 ;
        RECT 14.105 202.145 14.625 202.685 ;
        RECT 13.415 201.225 14.625 201.975 ;
        RECT 16.380 201.770 16.720 202.600 ;
        RECT 18.200 202.090 18.550 203.340 ;
        RECT 21.900 201.770 22.240 202.600 ;
        RECT 23.720 202.090 24.070 203.340 ;
        RECT 26.295 202.610 26.585 203.775 ;
        RECT 26.755 203.340 32.100 203.775 ;
        RECT 32.275 203.340 37.620 203.775 ;
        RECT 37.795 203.340 43.140 203.775 ;
        RECT 43.315 203.340 48.660 203.775 ;
        RECT 14.795 201.225 20.140 201.770 ;
        RECT 20.315 201.225 25.660 201.770 ;
        RECT 26.295 201.225 26.585 201.950 ;
        RECT 28.340 201.770 28.680 202.600 ;
        RECT 30.160 202.090 30.510 203.340 ;
        RECT 33.860 201.770 34.200 202.600 ;
        RECT 35.680 202.090 36.030 203.340 ;
        RECT 39.380 201.770 39.720 202.600 ;
        RECT 41.200 202.090 41.550 203.340 ;
        RECT 44.900 201.770 45.240 202.600 ;
        RECT 46.720 202.090 47.070 203.340 ;
        RECT 48.835 202.685 51.425 203.775 ;
        RECT 48.835 201.995 50.045 202.515 ;
        RECT 50.215 202.165 51.425 202.685 ;
        RECT 52.055 202.610 52.345 203.775 ;
        RECT 52.515 203.340 57.860 203.775 ;
        RECT 58.035 203.340 63.380 203.775 ;
        RECT 63.555 203.340 68.900 203.775 ;
        RECT 69.075 203.340 74.420 203.775 ;
        RECT 26.755 201.225 32.100 201.770 ;
        RECT 32.275 201.225 37.620 201.770 ;
        RECT 37.795 201.225 43.140 201.770 ;
        RECT 43.315 201.225 48.660 201.770 ;
        RECT 48.835 201.225 51.425 201.995 ;
        RECT 52.055 201.225 52.345 201.950 ;
        RECT 54.100 201.770 54.440 202.600 ;
        RECT 55.920 202.090 56.270 203.340 ;
        RECT 59.620 201.770 59.960 202.600 ;
        RECT 61.440 202.090 61.790 203.340 ;
        RECT 65.140 201.770 65.480 202.600 ;
        RECT 66.960 202.090 67.310 203.340 ;
        RECT 70.660 201.770 71.000 202.600 ;
        RECT 72.480 202.090 72.830 203.340 ;
        RECT 74.595 202.685 77.185 203.775 ;
        RECT 74.595 201.995 75.805 202.515 ;
        RECT 75.975 202.165 77.185 202.685 ;
        RECT 77.815 202.610 78.105 203.775 ;
        RECT 78.275 203.340 83.620 203.775 ;
        RECT 83.795 203.340 89.140 203.775 ;
        RECT 89.315 203.340 94.660 203.775 ;
        RECT 94.835 203.340 100.180 203.775 ;
        RECT 52.515 201.225 57.860 201.770 ;
        RECT 58.035 201.225 63.380 201.770 ;
        RECT 63.555 201.225 68.900 201.770 ;
        RECT 69.075 201.225 74.420 201.770 ;
        RECT 74.595 201.225 77.185 201.995 ;
        RECT 77.815 201.225 78.105 201.950 ;
        RECT 79.860 201.770 80.200 202.600 ;
        RECT 81.680 202.090 82.030 203.340 ;
        RECT 85.380 201.770 85.720 202.600 ;
        RECT 87.200 202.090 87.550 203.340 ;
        RECT 90.900 201.770 91.240 202.600 ;
        RECT 92.720 202.090 93.070 203.340 ;
        RECT 96.420 201.770 96.760 202.600 ;
        RECT 98.240 202.090 98.590 203.340 ;
        RECT 100.355 202.685 102.945 203.775 ;
        RECT 100.355 201.995 101.565 202.515 ;
        RECT 101.735 202.165 102.945 202.685 ;
        RECT 103.575 202.610 103.865 203.775 ;
        RECT 104.035 203.340 109.380 203.775 ;
        RECT 109.555 203.340 114.900 203.775 ;
        RECT 115.075 203.340 120.420 203.775 ;
        RECT 120.595 203.340 125.940 203.775 ;
        RECT 78.275 201.225 83.620 201.770 ;
        RECT 83.795 201.225 89.140 201.770 ;
        RECT 89.315 201.225 94.660 201.770 ;
        RECT 94.835 201.225 100.180 201.770 ;
        RECT 100.355 201.225 102.945 201.995 ;
        RECT 103.575 201.225 103.865 201.950 ;
        RECT 105.620 201.770 105.960 202.600 ;
        RECT 107.440 202.090 107.790 203.340 ;
        RECT 111.140 201.770 111.480 202.600 ;
        RECT 112.960 202.090 113.310 203.340 ;
        RECT 116.660 201.770 117.000 202.600 ;
        RECT 118.480 202.090 118.830 203.340 ;
        RECT 122.180 201.770 122.520 202.600 ;
        RECT 124.000 202.090 124.350 203.340 ;
        RECT 126.115 202.685 128.705 203.775 ;
        RECT 126.115 201.995 127.325 202.515 ;
        RECT 127.495 202.165 128.705 202.685 ;
        RECT 129.335 202.610 129.625 203.775 ;
        RECT 129.795 203.340 135.140 203.775 ;
        RECT 104.035 201.225 109.380 201.770 ;
        RECT 109.555 201.225 114.900 201.770 ;
        RECT 115.075 201.225 120.420 201.770 ;
        RECT 120.595 201.225 125.940 201.770 ;
        RECT 126.115 201.225 128.705 201.995 ;
        RECT 129.335 201.225 129.625 201.950 ;
        RECT 131.380 201.770 131.720 202.600 ;
        RECT 133.200 202.090 133.550 203.340 ;
        RECT 135.315 202.685 136.985 203.775 ;
        RECT 135.315 201.995 136.065 202.515 ;
        RECT 136.235 202.165 136.985 202.685 ;
        RECT 137.615 202.685 138.825 203.775 ;
        RECT 137.615 202.145 138.135 202.685 ;
        RECT 129.795 201.225 135.140 201.770 ;
        RECT 135.315 201.225 136.985 201.995 ;
        RECT 138.305 201.975 138.825 202.515 ;
        RECT 137.615 201.225 138.825 201.975 ;
        RECT 13.330 201.055 138.910 201.225 ;
        RECT 13.415 200.305 14.625 201.055 ;
        RECT 14.795 200.510 20.140 201.055 ;
        RECT 20.315 200.510 25.660 201.055 ;
        RECT 25.835 200.510 31.180 201.055 ;
        RECT 31.355 200.510 36.700 201.055 ;
        RECT 13.415 199.765 13.935 200.305 ;
        RECT 14.105 199.595 14.625 200.135 ;
        RECT 16.380 199.680 16.720 200.510 ;
        RECT 13.415 198.505 14.625 199.595 ;
        RECT 18.200 198.940 18.550 200.190 ;
        RECT 21.900 199.680 22.240 200.510 ;
        RECT 23.720 198.940 24.070 200.190 ;
        RECT 27.420 199.680 27.760 200.510 ;
        RECT 29.240 198.940 29.590 200.190 ;
        RECT 32.940 199.680 33.280 200.510 ;
        RECT 36.875 200.285 38.545 201.055 ;
        RECT 39.175 200.330 39.465 201.055 ;
        RECT 39.635 200.510 44.980 201.055 ;
        RECT 45.155 200.510 50.500 201.055 ;
        RECT 50.675 200.510 56.020 201.055 ;
        RECT 56.195 200.510 61.540 201.055 ;
        RECT 34.760 198.940 35.110 200.190 ;
        RECT 36.875 199.765 37.625 200.285 ;
        RECT 37.795 199.595 38.545 200.115 ;
        RECT 41.220 199.680 41.560 200.510 ;
        RECT 14.795 198.505 20.140 198.940 ;
        RECT 20.315 198.505 25.660 198.940 ;
        RECT 25.835 198.505 31.180 198.940 ;
        RECT 31.355 198.505 36.700 198.940 ;
        RECT 36.875 198.505 38.545 199.595 ;
        RECT 39.175 198.505 39.465 199.670 ;
        RECT 43.040 198.940 43.390 200.190 ;
        RECT 46.740 199.680 47.080 200.510 ;
        RECT 48.560 198.940 48.910 200.190 ;
        RECT 52.260 199.680 52.600 200.510 ;
        RECT 54.080 198.940 54.430 200.190 ;
        RECT 57.780 199.680 58.120 200.510 ;
        RECT 61.715 200.305 62.925 201.055 ;
        RECT 63.095 200.380 63.355 200.885 ;
        RECT 63.535 200.675 63.865 201.055 ;
        RECT 64.045 200.505 64.215 200.885 ;
        RECT 59.600 198.940 59.950 200.190 ;
        RECT 61.715 199.765 62.235 200.305 ;
        RECT 62.405 199.595 62.925 200.135 ;
        RECT 39.635 198.505 44.980 198.940 ;
        RECT 45.155 198.505 50.500 198.940 ;
        RECT 50.675 198.505 56.020 198.940 ;
        RECT 56.195 198.505 61.540 198.940 ;
        RECT 61.715 198.505 62.925 199.595 ;
        RECT 63.095 199.580 63.265 200.380 ;
        RECT 63.550 200.335 64.215 200.505 ;
        RECT 63.550 200.080 63.720 200.335 ;
        RECT 64.935 200.330 65.225 201.055 ;
        RECT 65.455 200.235 65.665 201.055 ;
        RECT 65.835 200.255 66.165 200.885 ;
        RECT 63.435 199.750 63.720 200.080 ;
        RECT 63.955 199.785 64.285 200.155 ;
        RECT 63.550 199.605 63.720 199.750 ;
        RECT 63.095 198.675 63.365 199.580 ;
        RECT 63.550 199.435 64.215 199.605 ;
        RECT 63.535 198.505 63.865 199.265 ;
        RECT 64.045 198.675 64.215 199.435 ;
        RECT 64.935 198.505 65.225 199.670 ;
        RECT 65.835 199.655 66.085 200.255 ;
        RECT 66.335 200.235 66.565 201.055 ;
        RECT 66.865 200.505 67.035 200.795 ;
        RECT 67.205 200.675 67.535 201.055 ;
        RECT 66.865 200.335 67.530 200.505 ;
        RECT 66.255 199.815 66.585 200.065 ;
        RECT 65.455 198.505 65.665 199.645 ;
        RECT 65.835 198.675 66.165 199.655 ;
        RECT 66.335 198.505 66.565 199.645 ;
        RECT 66.780 199.515 67.130 200.165 ;
        RECT 67.300 199.345 67.530 200.335 ;
        RECT 66.865 199.175 67.530 199.345 ;
        RECT 66.865 198.675 67.035 199.175 ;
        RECT 67.205 198.505 67.535 199.005 ;
        RECT 67.705 198.675 67.890 200.795 ;
        RECT 68.145 200.595 68.395 201.055 ;
        RECT 68.565 200.605 68.900 200.775 ;
        RECT 69.095 200.605 69.770 200.775 ;
        RECT 68.565 200.465 68.735 200.605 ;
        RECT 68.060 199.475 68.340 200.425 ;
        RECT 68.510 200.335 68.735 200.465 ;
        RECT 68.510 199.230 68.680 200.335 ;
        RECT 68.905 200.185 69.430 200.405 ;
        RECT 68.850 199.420 69.090 200.015 ;
        RECT 69.260 199.485 69.430 200.185 ;
        RECT 69.600 199.825 69.770 200.605 ;
        RECT 70.090 200.555 70.460 201.055 ;
        RECT 70.640 200.605 71.045 200.775 ;
        RECT 71.215 200.605 72.000 200.775 ;
        RECT 70.640 200.375 70.810 200.605 ;
        RECT 69.980 200.075 70.810 200.375 ;
        RECT 71.195 200.105 71.660 200.435 ;
        RECT 69.980 200.045 70.180 200.075 ;
        RECT 70.300 199.825 70.470 199.895 ;
        RECT 69.600 199.655 70.470 199.825 ;
        RECT 69.960 199.565 70.470 199.655 ;
        RECT 68.510 199.100 68.815 199.230 ;
        RECT 69.260 199.120 69.790 199.485 ;
        RECT 68.130 198.505 68.395 198.965 ;
        RECT 68.565 198.675 68.815 199.100 ;
        RECT 69.960 198.950 70.130 199.565 ;
        RECT 69.025 198.780 70.130 198.950 ;
        RECT 70.300 198.505 70.470 199.305 ;
        RECT 70.640 199.005 70.810 200.075 ;
        RECT 70.980 199.175 71.170 199.895 ;
        RECT 71.340 199.145 71.660 200.105 ;
        RECT 71.830 200.145 72.000 200.605 ;
        RECT 72.275 200.525 72.485 201.055 ;
        RECT 72.745 200.315 73.075 200.840 ;
        RECT 73.245 200.445 73.415 201.055 ;
        RECT 73.585 200.400 73.915 200.835 ;
        RECT 73.585 200.315 73.965 200.400 ;
        RECT 72.875 200.145 73.075 200.315 ;
        RECT 73.740 200.275 73.965 200.315 ;
        RECT 71.830 199.815 72.705 200.145 ;
        RECT 72.875 199.815 73.625 200.145 ;
        RECT 70.640 198.675 70.890 199.005 ;
        RECT 71.830 198.975 72.000 199.815 ;
        RECT 72.875 199.610 73.065 199.815 ;
        RECT 73.795 199.695 73.965 200.275 ;
        RECT 73.750 199.645 73.965 199.695 ;
        RECT 72.170 199.235 73.065 199.610 ;
        RECT 73.575 199.565 73.965 199.645 ;
        RECT 74.135 200.315 74.520 200.885 ;
        RECT 74.690 200.595 75.015 201.055 ;
        RECT 75.535 200.425 75.815 200.885 ;
        RECT 74.135 199.645 74.415 200.315 ;
        RECT 74.690 200.255 75.815 200.425 ;
        RECT 74.690 200.145 75.140 200.255 ;
        RECT 74.585 199.815 75.140 200.145 ;
        RECT 76.005 200.085 76.405 200.885 ;
        RECT 76.805 200.595 77.075 201.055 ;
        RECT 77.245 200.425 77.530 200.885 ;
        RECT 77.875 200.575 78.155 201.055 ;
        RECT 71.115 198.805 72.000 198.975 ;
        RECT 72.180 198.505 72.495 199.005 ;
        RECT 72.725 198.675 73.065 199.235 ;
        RECT 73.235 198.505 73.405 199.515 ;
        RECT 73.575 198.720 73.905 199.565 ;
        RECT 74.135 198.675 74.520 199.645 ;
        RECT 74.690 199.355 75.140 199.815 ;
        RECT 75.310 199.525 76.405 200.085 ;
        RECT 74.690 199.135 75.815 199.355 ;
        RECT 74.690 198.505 75.015 198.965 ;
        RECT 75.535 198.675 75.815 199.135 ;
        RECT 76.005 198.675 76.405 199.525 ;
        RECT 76.575 200.255 77.530 200.425 ;
        RECT 78.325 200.405 78.585 200.795 ;
        RECT 78.760 200.575 79.015 201.055 ;
        RECT 79.185 200.405 79.480 200.795 ;
        RECT 79.660 200.575 79.935 201.055 ;
        RECT 80.105 200.555 80.405 200.885 ;
        RECT 76.575 199.355 76.785 200.255 ;
        RECT 77.830 200.235 79.480 200.405 ;
        RECT 76.955 199.525 77.645 200.085 ;
        RECT 77.830 199.725 78.235 200.235 ;
        RECT 78.405 199.895 79.545 200.065 ;
        RECT 77.830 199.555 78.585 199.725 ;
        RECT 76.575 199.135 77.530 199.355 ;
        RECT 76.805 198.505 77.075 198.965 ;
        RECT 77.245 198.675 77.530 199.135 ;
        RECT 77.870 198.505 78.155 199.375 ;
        RECT 78.325 199.305 78.585 199.555 ;
        RECT 79.375 199.645 79.545 199.895 ;
        RECT 79.715 199.815 80.065 200.385 ;
        RECT 80.235 199.645 80.405 200.555 ;
        RECT 80.575 200.510 85.920 201.055 ;
        RECT 82.160 199.680 82.500 200.510 ;
        RECT 86.095 200.285 89.605 201.055 ;
        RECT 90.695 200.330 90.985 201.055 ;
        RECT 91.155 200.510 96.500 201.055 ;
        RECT 96.675 200.510 102.020 201.055 ;
        RECT 102.195 200.510 107.540 201.055 ;
        RECT 107.715 200.510 113.060 201.055 ;
        RECT 79.375 199.475 80.405 199.645 ;
        RECT 78.325 199.135 79.445 199.305 ;
        RECT 78.325 198.675 78.585 199.135 ;
        RECT 78.760 198.505 79.015 198.965 ;
        RECT 79.185 198.675 79.445 199.135 ;
        RECT 79.615 198.505 79.925 199.305 ;
        RECT 80.095 198.675 80.405 199.475 ;
        RECT 83.980 198.940 84.330 200.190 ;
        RECT 86.095 199.765 87.745 200.285 ;
        RECT 87.915 199.595 89.605 200.115 ;
        RECT 92.740 199.680 93.080 200.510 ;
        RECT 80.575 198.505 85.920 198.940 ;
        RECT 86.095 198.505 89.605 199.595 ;
        RECT 90.695 198.505 90.985 199.670 ;
        RECT 94.560 198.940 94.910 200.190 ;
        RECT 98.260 199.680 98.600 200.510 ;
        RECT 100.080 198.940 100.430 200.190 ;
        RECT 103.780 199.680 104.120 200.510 ;
        RECT 105.600 198.940 105.950 200.190 ;
        RECT 109.300 199.680 109.640 200.510 ;
        RECT 113.240 200.215 113.500 201.055 ;
        RECT 113.675 200.310 113.930 200.885 ;
        RECT 114.100 200.675 114.430 201.055 ;
        RECT 114.645 200.505 114.815 200.885 ;
        RECT 114.100 200.335 114.815 200.505 ;
        RECT 111.120 198.940 111.470 200.190 ;
        RECT 91.155 198.505 96.500 198.940 ;
        RECT 96.675 198.505 102.020 198.940 ;
        RECT 102.195 198.505 107.540 198.940 ;
        RECT 107.715 198.505 113.060 198.940 ;
        RECT 113.240 198.505 113.500 199.655 ;
        RECT 113.675 199.580 113.845 200.310 ;
        RECT 114.100 200.145 114.270 200.335 ;
        RECT 115.075 200.305 116.285 201.055 ;
        RECT 116.455 200.330 116.745 201.055 ;
        RECT 116.915 200.510 122.260 201.055 ;
        RECT 122.435 200.510 127.780 201.055 ;
        RECT 127.955 200.510 133.300 201.055 ;
        RECT 114.015 199.815 114.270 200.145 ;
        RECT 114.100 199.605 114.270 199.815 ;
        RECT 114.550 199.785 114.905 200.155 ;
        RECT 115.075 199.765 115.595 200.305 ;
        RECT 113.675 198.675 113.930 199.580 ;
        RECT 114.100 199.435 114.815 199.605 ;
        RECT 115.765 199.595 116.285 200.135 ;
        RECT 118.500 199.680 118.840 200.510 ;
        RECT 114.100 198.505 114.430 199.265 ;
        RECT 114.645 198.675 114.815 199.435 ;
        RECT 115.075 198.505 116.285 199.595 ;
        RECT 116.455 198.505 116.745 199.670 ;
        RECT 120.320 198.940 120.670 200.190 ;
        RECT 124.020 199.680 124.360 200.510 ;
        RECT 125.840 198.940 126.190 200.190 ;
        RECT 129.540 199.680 129.880 200.510 ;
        RECT 133.475 200.285 136.985 201.055 ;
        RECT 137.615 200.305 138.825 201.055 ;
        RECT 131.360 198.940 131.710 200.190 ;
        RECT 133.475 199.765 135.125 200.285 ;
        RECT 135.295 199.595 136.985 200.115 ;
        RECT 116.915 198.505 122.260 198.940 ;
        RECT 122.435 198.505 127.780 198.940 ;
        RECT 127.955 198.505 133.300 198.940 ;
        RECT 133.475 198.505 136.985 199.595 ;
        RECT 137.615 199.595 138.135 200.135 ;
        RECT 138.305 199.765 138.825 200.305 ;
        RECT 137.615 198.505 138.825 199.595 ;
        RECT 13.330 198.335 138.910 198.505 ;
        RECT 13.415 197.245 14.625 198.335 ;
        RECT 14.795 197.900 20.140 198.335 ;
        RECT 20.315 197.900 25.660 198.335 ;
        RECT 13.415 196.535 13.935 197.075 ;
        RECT 14.105 196.705 14.625 197.245 ;
        RECT 13.415 195.785 14.625 196.535 ;
        RECT 16.380 196.330 16.720 197.160 ;
        RECT 18.200 196.650 18.550 197.900 ;
        RECT 21.900 196.330 22.240 197.160 ;
        RECT 23.720 196.650 24.070 197.900 ;
        RECT 26.295 197.170 26.585 198.335 ;
        RECT 26.755 197.900 32.100 198.335 ;
        RECT 32.275 197.900 37.620 198.335 ;
        RECT 37.795 197.900 43.140 198.335 ;
        RECT 43.315 197.900 48.660 198.335 ;
        RECT 14.795 195.785 20.140 196.330 ;
        RECT 20.315 195.785 25.660 196.330 ;
        RECT 26.295 195.785 26.585 196.510 ;
        RECT 28.340 196.330 28.680 197.160 ;
        RECT 30.160 196.650 30.510 197.900 ;
        RECT 33.860 196.330 34.200 197.160 ;
        RECT 35.680 196.650 36.030 197.900 ;
        RECT 39.380 196.330 39.720 197.160 ;
        RECT 41.200 196.650 41.550 197.900 ;
        RECT 44.900 196.330 45.240 197.160 ;
        RECT 46.720 196.650 47.070 197.900 ;
        RECT 48.835 197.245 51.425 198.335 ;
        RECT 48.835 196.555 50.045 197.075 ;
        RECT 50.215 196.725 51.425 197.245 ;
        RECT 52.055 197.170 52.345 198.335 ;
        RECT 52.515 197.900 57.860 198.335 ;
        RECT 26.755 195.785 32.100 196.330 ;
        RECT 32.275 195.785 37.620 196.330 ;
        RECT 37.795 195.785 43.140 196.330 ;
        RECT 43.315 195.785 48.660 196.330 ;
        RECT 48.835 195.785 51.425 196.555 ;
        RECT 52.055 195.785 52.345 196.510 ;
        RECT 54.100 196.330 54.440 197.160 ;
        RECT 55.920 196.650 56.270 197.900 ;
        RECT 58.035 197.245 60.625 198.335 ;
        RECT 58.035 196.555 59.245 197.075 ;
        RECT 59.415 196.725 60.625 197.245 ;
        RECT 61.255 197.195 61.640 198.165 ;
        RECT 61.810 197.875 62.135 198.335 ;
        RECT 62.655 197.705 62.935 198.165 ;
        RECT 61.810 197.485 62.935 197.705 ;
        RECT 52.515 195.785 57.860 196.330 ;
        RECT 58.035 195.785 60.625 196.555 ;
        RECT 61.255 196.525 61.535 197.195 ;
        RECT 61.810 197.025 62.260 197.485 ;
        RECT 63.125 197.315 63.525 198.165 ;
        RECT 63.925 197.875 64.195 198.335 ;
        RECT 64.365 197.705 64.650 198.165 ;
        RECT 61.705 196.695 62.260 197.025 ;
        RECT 62.430 196.755 63.525 197.315 ;
        RECT 61.810 196.585 62.260 196.695 ;
        RECT 61.255 195.955 61.640 196.525 ;
        RECT 61.810 196.415 62.935 196.585 ;
        RECT 61.810 195.785 62.135 196.245 ;
        RECT 62.655 195.955 62.935 196.415 ;
        RECT 63.125 195.955 63.525 196.755 ;
        RECT 63.695 197.485 64.650 197.705 ;
        RECT 63.695 196.585 63.905 197.485 ;
        RECT 64.075 196.755 64.765 197.315 ;
        RECT 65.865 197.195 66.195 198.335 ;
        RECT 66.725 197.365 67.055 198.150 ;
        RECT 67.235 197.825 67.535 198.335 ;
        RECT 67.705 197.655 68.035 198.165 ;
        RECT 68.205 197.825 68.835 198.335 ;
        RECT 69.415 197.825 69.795 197.995 ;
        RECT 69.965 197.825 70.265 198.335 ;
        RECT 69.625 197.655 69.795 197.825 ;
        RECT 70.545 197.665 70.715 198.165 ;
        RECT 70.885 197.835 71.215 198.335 ;
        RECT 66.375 197.195 67.055 197.365 ;
        RECT 67.235 197.485 69.455 197.655 ;
        RECT 65.855 196.775 66.205 197.025 ;
        RECT 66.375 196.595 66.545 197.195 ;
        RECT 66.715 196.775 67.065 197.025 ;
        RECT 63.695 196.415 64.650 196.585 ;
        RECT 63.925 195.785 64.195 196.245 ;
        RECT 64.365 195.955 64.650 196.415 ;
        RECT 65.865 195.785 66.135 196.595 ;
        RECT 66.305 195.955 66.635 196.595 ;
        RECT 66.805 195.785 67.045 196.595 ;
        RECT 67.235 196.525 67.405 197.485 ;
        RECT 67.575 197.145 69.115 197.315 ;
        RECT 67.575 196.695 67.820 197.145 ;
        RECT 68.080 196.775 68.775 196.975 ;
        RECT 68.945 196.945 69.115 197.145 ;
        RECT 69.285 197.285 69.455 197.485 ;
        RECT 69.625 197.455 70.285 197.655 ;
        RECT 70.545 197.495 71.210 197.665 ;
        RECT 69.285 197.115 69.945 197.285 ;
        RECT 68.945 196.775 69.545 196.945 ;
        RECT 69.775 196.695 69.945 197.115 ;
        RECT 67.235 195.980 67.700 196.525 ;
        RECT 68.205 195.785 68.375 196.605 ;
        RECT 68.545 196.525 69.455 196.605 ;
        RECT 70.115 196.525 70.285 197.455 ;
        RECT 70.460 196.675 70.810 197.325 ;
        RECT 68.545 196.435 69.795 196.525 ;
        RECT 68.545 195.955 68.875 196.435 ;
        RECT 69.285 196.355 69.795 196.435 ;
        RECT 69.045 195.785 69.395 196.175 ;
        RECT 69.565 195.955 69.795 196.355 ;
        RECT 69.965 196.045 70.285 196.525 ;
        RECT 70.980 196.505 71.210 197.495 ;
        RECT 70.545 196.335 71.210 196.505 ;
        RECT 70.545 196.045 70.715 196.335 ;
        RECT 70.885 195.785 71.215 196.165 ;
        RECT 71.385 196.045 71.570 198.165 ;
        RECT 71.810 197.875 72.075 198.335 ;
        RECT 72.245 197.740 72.495 198.165 ;
        RECT 72.705 197.890 73.810 198.060 ;
        RECT 72.190 197.610 72.495 197.740 ;
        RECT 71.740 196.415 72.020 197.365 ;
        RECT 72.190 196.505 72.360 197.610 ;
        RECT 72.530 196.825 72.770 197.420 ;
        RECT 72.940 197.355 73.470 197.720 ;
        RECT 72.940 196.655 73.110 197.355 ;
        RECT 73.640 197.275 73.810 197.890 ;
        RECT 73.980 197.535 74.150 198.335 ;
        RECT 74.320 197.835 74.570 198.165 ;
        RECT 74.795 197.865 75.680 198.035 ;
        RECT 73.640 197.185 74.150 197.275 ;
        RECT 72.190 196.375 72.415 196.505 ;
        RECT 72.585 196.435 73.110 196.655 ;
        RECT 73.280 197.015 74.150 197.185 ;
        RECT 71.825 195.785 72.075 196.245 ;
        RECT 72.245 196.235 72.415 196.375 ;
        RECT 73.280 196.235 73.450 197.015 ;
        RECT 73.980 196.945 74.150 197.015 ;
        RECT 73.660 196.765 73.860 196.795 ;
        RECT 74.320 196.765 74.490 197.835 ;
        RECT 74.660 196.945 74.850 197.665 ;
        RECT 73.660 196.465 74.490 196.765 ;
        RECT 75.020 196.735 75.340 197.695 ;
        RECT 72.245 196.065 72.580 196.235 ;
        RECT 72.775 196.065 73.450 196.235 ;
        RECT 73.770 195.785 74.140 196.285 ;
        RECT 74.320 196.235 74.490 196.465 ;
        RECT 74.875 196.405 75.340 196.735 ;
        RECT 75.510 197.025 75.680 197.865 ;
        RECT 75.860 197.835 76.175 198.335 ;
        RECT 76.405 197.605 76.745 198.165 ;
        RECT 75.850 197.230 76.745 197.605 ;
        RECT 76.915 197.325 77.085 198.335 ;
        RECT 76.555 197.025 76.745 197.230 ;
        RECT 77.255 197.275 77.585 198.120 ;
        RECT 77.255 197.195 77.645 197.275 ;
        RECT 77.430 197.145 77.645 197.195 ;
        RECT 77.815 197.170 78.105 198.335 ;
        RECT 78.460 197.365 78.850 197.540 ;
        RECT 79.335 197.535 79.665 198.335 ;
        RECT 79.835 197.545 80.370 198.165 ;
        RECT 80.575 197.900 85.920 198.335 ;
        RECT 78.460 197.195 79.885 197.365 ;
        RECT 75.510 196.695 76.385 197.025 ;
        RECT 76.555 196.695 77.305 197.025 ;
        RECT 75.510 196.235 75.680 196.695 ;
        RECT 76.555 196.525 76.755 196.695 ;
        RECT 77.475 196.565 77.645 197.145 ;
        RECT 77.420 196.525 77.645 196.565 ;
        RECT 74.320 196.065 74.725 196.235 ;
        RECT 74.895 196.065 75.680 196.235 ;
        RECT 75.955 195.785 76.165 196.315 ;
        RECT 76.425 196.000 76.755 196.525 ;
        RECT 77.265 196.440 77.645 196.525 ;
        RECT 76.925 195.785 77.095 196.395 ;
        RECT 77.265 196.005 77.595 196.440 ;
        RECT 77.815 195.785 78.105 196.510 ;
        RECT 78.335 196.465 78.690 197.025 ;
        RECT 78.860 196.295 79.030 197.195 ;
        RECT 79.200 196.465 79.465 197.025 ;
        RECT 79.715 196.695 79.885 197.195 ;
        RECT 80.055 196.525 80.370 197.545 ;
        RECT 78.440 195.785 78.680 196.295 ;
        RECT 78.860 195.965 79.140 196.295 ;
        RECT 79.370 195.785 79.585 196.295 ;
        RECT 79.755 195.955 80.370 196.525 ;
        RECT 82.160 196.330 82.500 197.160 ;
        RECT 83.980 196.650 84.330 197.900 ;
        RECT 86.095 197.245 88.685 198.335 ;
        RECT 86.095 196.555 87.305 197.075 ;
        RECT 87.475 196.725 88.685 197.245 ;
        RECT 89.325 197.195 89.655 198.335 ;
        RECT 90.185 197.365 90.515 198.150 ;
        RECT 89.835 197.195 90.515 197.365 ;
        RECT 91.675 197.275 92.005 198.120 ;
        RECT 92.175 197.325 92.345 198.335 ;
        RECT 92.515 197.605 92.855 198.165 ;
        RECT 93.085 197.835 93.400 198.335 ;
        RECT 93.580 197.865 94.465 198.035 ;
        RECT 91.615 197.195 92.005 197.275 ;
        RECT 92.515 197.230 93.410 197.605 ;
        RECT 89.315 196.775 89.665 197.025 ;
        RECT 89.835 196.595 90.005 197.195 ;
        RECT 91.615 197.145 91.830 197.195 ;
        RECT 90.175 196.775 90.525 197.025 ;
        RECT 80.575 195.785 85.920 196.330 ;
        RECT 86.095 195.785 88.685 196.555 ;
        RECT 89.325 195.785 89.595 196.595 ;
        RECT 89.765 195.955 90.095 196.595 ;
        RECT 90.265 195.785 90.505 196.595 ;
        RECT 91.615 196.565 91.785 197.145 ;
        RECT 92.515 197.025 92.705 197.230 ;
        RECT 93.580 197.025 93.750 197.865 ;
        RECT 94.690 197.835 94.940 198.165 ;
        RECT 91.955 196.695 92.705 197.025 ;
        RECT 92.875 196.695 93.750 197.025 ;
        RECT 91.615 196.525 91.840 196.565 ;
        RECT 92.505 196.525 92.705 196.695 ;
        RECT 91.615 196.440 91.995 196.525 ;
        RECT 91.665 196.005 91.995 196.440 ;
        RECT 92.165 195.785 92.335 196.395 ;
        RECT 92.505 196.000 92.835 196.525 ;
        RECT 93.095 195.785 93.305 196.315 ;
        RECT 93.580 196.235 93.750 196.695 ;
        RECT 93.920 196.735 94.240 197.695 ;
        RECT 94.410 196.945 94.600 197.665 ;
        RECT 94.770 196.765 94.940 197.835 ;
        RECT 95.110 197.535 95.280 198.335 ;
        RECT 95.450 197.890 96.555 198.060 ;
        RECT 95.450 197.275 95.620 197.890 ;
        RECT 96.765 197.740 97.015 198.165 ;
        RECT 97.185 197.875 97.450 198.335 ;
        RECT 95.790 197.355 96.320 197.720 ;
        RECT 96.765 197.610 97.070 197.740 ;
        RECT 95.110 197.185 95.620 197.275 ;
        RECT 95.110 197.015 95.980 197.185 ;
        RECT 95.110 196.945 95.280 197.015 ;
        RECT 95.400 196.765 95.600 196.795 ;
        RECT 93.920 196.405 94.385 196.735 ;
        RECT 94.770 196.465 95.600 196.765 ;
        RECT 94.770 196.235 94.940 196.465 ;
        RECT 93.580 196.065 94.365 196.235 ;
        RECT 94.535 196.065 94.940 196.235 ;
        RECT 95.120 195.785 95.490 196.285 ;
        RECT 95.810 196.235 95.980 197.015 ;
        RECT 96.150 196.655 96.320 197.355 ;
        RECT 96.490 196.825 96.730 197.420 ;
        RECT 96.150 196.435 96.675 196.655 ;
        RECT 96.900 196.505 97.070 197.610 ;
        RECT 96.845 196.375 97.070 196.505 ;
        RECT 97.240 196.415 97.520 197.365 ;
        RECT 96.845 196.235 97.015 196.375 ;
        RECT 95.810 196.065 96.485 196.235 ;
        RECT 96.680 196.065 97.015 196.235 ;
        RECT 97.185 195.785 97.435 196.245 ;
        RECT 97.690 196.045 97.875 198.165 ;
        RECT 98.045 197.835 98.375 198.335 ;
        RECT 98.545 197.665 98.715 198.165 ;
        RECT 99.025 197.875 99.235 198.335 ;
        RECT 99.725 197.745 100.225 198.165 ;
        RECT 98.050 197.495 98.715 197.665 ;
        RECT 98.050 196.505 98.280 197.495 ;
        RECT 98.450 196.675 98.800 197.325 ;
        RECT 98.050 196.335 98.715 196.505 ;
        RECT 98.975 196.365 99.215 197.690 ;
        RECT 99.385 197.535 100.225 197.745 ;
        RECT 99.385 196.525 99.555 197.535 ;
        RECT 99.725 197.115 100.125 197.365 ;
        RECT 100.415 197.315 100.615 198.105 ;
        RECT 100.295 197.145 100.615 197.315 ;
        RECT 100.785 197.155 101.105 198.335 ;
        RECT 101.280 197.195 101.600 198.335 ;
        RECT 99.725 196.695 99.895 197.115 ;
        RECT 100.295 196.945 100.475 197.145 ;
        RECT 101.780 197.025 101.975 198.075 ;
        RECT 102.155 197.485 102.485 198.165 ;
        RECT 102.685 197.535 102.940 198.335 ;
        RECT 102.155 197.205 102.505 197.485 ;
        RECT 101.340 196.975 101.600 197.025 ;
        RECT 100.110 196.775 100.475 196.945 ;
        RECT 100.645 196.775 101.105 196.975 ;
        RECT 101.335 196.805 101.600 196.975 ;
        RECT 101.340 196.695 101.600 196.805 ;
        RECT 101.780 196.695 102.165 197.025 ;
        RECT 102.335 196.825 102.505 197.205 ;
        RECT 102.695 196.995 102.940 197.355 ;
        RECT 103.575 197.170 103.865 198.335 ;
        RECT 104.035 197.245 107.545 198.335 ;
        RECT 108.695 197.275 109.025 198.120 ;
        RECT 109.195 197.325 109.365 198.335 ;
        RECT 109.535 197.605 109.875 198.165 ;
        RECT 110.105 197.835 110.420 198.335 ;
        RECT 110.600 197.865 111.485 198.035 ;
        RECT 102.335 196.655 102.855 196.825 ;
        RECT 100.075 196.525 101.105 196.565 ;
        RECT 99.385 196.345 99.735 196.525 ;
        RECT 99.905 196.395 101.105 196.525 ;
        RECT 98.045 195.785 98.375 196.165 ;
        RECT 98.545 196.045 98.715 196.335 ;
        RECT 99.905 196.175 100.235 196.395 ;
        RECT 98.975 195.995 100.235 196.175 ;
        RECT 100.425 195.785 100.595 196.225 ;
        RECT 100.765 195.980 101.105 196.395 ;
        RECT 101.280 196.315 102.495 196.485 ;
        RECT 101.280 195.965 101.570 196.315 ;
        RECT 101.765 195.785 102.095 196.145 ;
        RECT 102.265 196.010 102.495 196.315 ;
        RECT 102.685 196.295 102.855 196.655 ;
        RECT 104.035 196.555 105.685 197.075 ;
        RECT 105.855 196.725 107.545 197.245 ;
        RECT 108.635 197.195 109.025 197.275 ;
        RECT 109.535 197.230 110.430 197.605 ;
        RECT 108.635 197.145 108.850 197.195 ;
        RECT 108.635 196.565 108.805 197.145 ;
        RECT 109.535 197.025 109.725 197.230 ;
        RECT 110.600 197.025 110.770 197.865 ;
        RECT 111.710 197.835 111.960 198.165 ;
        RECT 108.975 196.695 109.725 197.025 ;
        RECT 109.895 196.695 110.770 197.025 ;
        RECT 102.685 196.125 102.885 196.295 ;
        RECT 102.685 196.090 102.855 196.125 ;
        RECT 103.575 195.785 103.865 196.510 ;
        RECT 104.035 195.785 107.545 196.555 ;
        RECT 108.635 196.525 108.860 196.565 ;
        RECT 109.525 196.525 109.725 196.695 ;
        RECT 108.635 196.440 109.015 196.525 ;
        RECT 108.685 196.005 109.015 196.440 ;
        RECT 109.185 195.785 109.355 196.395 ;
        RECT 109.525 196.000 109.855 196.525 ;
        RECT 110.115 195.785 110.325 196.315 ;
        RECT 110.600 196.235 110.770 196.695 ;
        RECT 110.940 196.735 111.260 197.695 ;
        RECT 111.430 196.945 111.620 197.665 ;
        RECT 111.790 196.765 111.960 197.835 ;
        RECT 112.130 197.535 112.300 198.335 ;
        RECT 112.470 197.890 113.575 198.060 ;
        RECT 112.470 197.275 112.640 197.890 ;
        RECT 113.785 197.740 114.035 198.165 ;
        RECT 114.205 197.875 114.470 198.335 ;
        RECT 112.810 197.355 113.340 197.720 ;
        RECT 113.785 197.610 114.090 197.740 ;
        RECT 112.130 197.185 112.640 197.275 ;
        RECT 112.130 197.015 113.000 197.185 ;
        RECT 112.130 196.945 112.300 197.015 ;
        RECT 112.420 196.765 112.620 196.795 ;
        RECT 110.940 196.405 111.405 196.735 ;
        RECT 111.790 196.465 112.620 196.765 ;
        RECT 111.790 196.235 111.960 196.465 ;
        RECT 110.600 196.065 111.385 196.235 ;
        RECT 111.555 196.065 111.960 196.235 ;
        RECT 112.140 195.785 112.510 196.285 ;
        RECT 112.830 196.235 113.000 197.015 ;
        RECT 113.170 196.655 113.340 197.355 ;
        RECT 113.510 196.825 113.750 197.420 ;
        RECT 113.170 196.435 113.695 196.655 ;
        RECT 113.920 196.505 114.090 197.610 ;
        RECT 113.865 196.375 114.090 196.505 ;
        RECT 114.260 196.415 114.540 197.365 ;
        RECT 113.865 196.235 114.035 196.375 ;
        RECT 112.830 196.065 113.505 196.235 ;
        RECT 113.700 196.065 114.035 196.235 ;
        RECT 114.205 195.785 114.455 196.245 ;
        RECT 114.710 196.045 114.895 198.165 ;
        RECT 115.065 197.835 115.395 198.335 ;
        RECT 115.565 197.665 115.735 198.165 ;
        RECT 115.070 197.495 115.735 197.665 ;
        RECT 115.070 196.505 115.300 197.495 ;
        RECT 115.470 196.675 115.820 197.325 ;
        RECT 116.055 197.275 116.385 198.120 ;
        RECT 116.555 197.325 116.725 198.335 ;
        RECT 116.895 197.605 117.235 198.165 ;
        RECT 117.465 197.835 117.780 198.335 ;
        RECT 117.960 197.865 118.845 198.035 ;
        RECT 115.995 197.195 116.385 197.275 ;
        RECT 116.895 197.230 117.790 197.605 ;
        RECT 115.995 197.145 116.210 197.195 ;
        RECT 115.995 196.565 116.165 197.145 ;
        RECT 116.895 197.025 117.085 197.230 ;
        RECT 117.960 197.025 118.130 197.865 ;
        RECT 119.070 197.835 119.320 198.165 ;
        RECT 116.335 196.695 117.085 197.025 ;
        RECT 117.255 196.695 118.130 197.025 ;
        RECT 115.995 196.525 116.220 196.565 ;
        RECT 116.885 196.525 117.085 196.695 ;
        RECT 115.070 196.335 115.735 196.505 ;
        RECT 115.995 196.440 116.375 196.525 ;
        RECT 115.065 195.785 115.395 196.165 ;
        RECT 115.565 196.045 115.735 196.335 ;
        RECT 116.045 196.005 116.375 196.440 ;
        RECT 116.545 195.785 116.715 196.395 ;
        RECT 116.885 196.000 117.215 196.525 ;
        RECT 117.475 195.785 117.685 196.315 ;
        RECT 117.960 196.235 118.130 196.695 ;
        RECT 118.300 196.735 118.620 197.695 ;
        RECT 118.790 196.945 118.980 197.665 ;
        RECT 119.150 196.765 119.320 197.835 ;
        RECT 119.490 197.535 119.660 198.335 ;
        RECT 119.830 197.890 120.935 198.060 ;
        RECT 119.830 197.275 120.000 197.890 ;
        RECT 121.145 197.740 121.395 198.165 ;
        RECT 121.565 197.875 121.830 198.335 ;
        RECT 120.170 197.355 120.700 197.720 ;
        RECT 121.145 197.610 121.450 197.740 ;
        RECT 119.490 197.185 120.000 197.275 ;
        RECT 119.490 197.015 120.360 197.185 ;
        RECT 119.490 196.945 119.660 197.015 ;
        RECT 119.780 196.765 119.980 196.795 ;
        RECT 118.300 196.405 118.765 196.735 ;
        RECT 119.150 196.465 119.980 196.765 ;
        RECT 119.150 196.235 119.320 196.465 ;
        RECT 117.960 196.065 118.745 196.235 ;
        RECT 118.915 196.065 119.320 196.235 ;
        RECT 119.500 195.785 119.870 196.285 ;
        RECT 120.190 196.235 120.360 197.015 ;
        RECT 120.530 196.655 120.700 197.355 ;
        RECT 120.870 196.825 121.110 197.420 ;
        RECT 120.530 196.435 121.055 196.655 ;
        RECT 121.280 196.505 121.450 197.610 ;
        RECT 121.225 196.375 121.450 196.505 ;
        RECT 121.620 196.415 121.900 197.365 ;
        RECT 121.225 196.235 121.395 196.375 ;
        RECT 120.190 196.065 120.865 196.235 ;
        RECT 121.060 196.065 121.395 196.235 ;
        RECT 121.565 195.785 121.815 196.245 ;
        RECT 122.070 196.045 122.255 198.165 ;
        RECT 122.425 197.835 122.755 198.335 ;
        RECT 122.925 197.665 123.095 198.165 ;
        RECT 123.355 197.900 128.700 198.335 ;
        RECT 122.430 197.495 123.095 197.665 ;
        RECT 122.430 196.505 122.660 197.495 ;
        RECT 122.830 196.675 123.180 197.325 ;
        RECT 122.430 196.335 123.095 196.505 ;
        RECT 122.425 195.785 122.755 196.165 ;
        RECT 122.925 196.045 123.095 196.335 ;
        RECT 124.940 196.330 125.280 197.160 ;
        RECT 126.760 196.650 127.110 197.900 ;
        RECT 129.335 197.170 129.625 198.335 ;
        RECT 129.795 197.900 135.140 198.335 ;
        RECT 123.355 195.785 128.700 196.330 ;
        RECT 129.335 195.785 129.625 196.510 ;
        RECT 131.380 196.330 131.720 197.160 ;
        RECT 133.200 196.650 133.550 197.900 ;
        RECT 135.315 197.245 136.985 198.335 ;
        RECT 135.315 196.555 136.065 197.075 ;
        RECT 136.235 196.725 136.985 197.245 ;
        RECT 137.615 197.245 138.825 198.335 ;
        RECT 137.615 196.705 138.135 197.245 ;
        RECT 129.795 195.785 135.140 196.330 ;
        RECT 135.315 195.785 136.985 196.555 ;
        RECT 138.305 196.535 138.825 197.075 ;
        RECT 137.615 195.785 138.825 196.535 ;
        RECT 13.330 195.615 138.910 195.785 ;
        RECT 13.415 194.865 14.625 195.615 ;
        RECT 14.795 195.070 20.140 195.615 ;
        RECT 20.315 195.070 25.660 195.615 ;
        RECT 25.835 195.070 31.180 195.615 ;
        RECT 13.415 194.325 13.935 194.865 ;
        RECT 14.105 194.155 14.625 194.695 ;
        RECT 16.380 194.240 16.720 195.070 ;
        RECT 13.415 193.065 14.625 194.155 ;
        RECT 18.200 193.500 18.550 194.750 ;
        RECT 21.900 194.240 22.240 195.070 ;
        RECT 23.720 193.500 24.070 194.750 ;
        RECT 27.420 194.240 27.760 195.070 ;
        RECT 32.360 195.045 32.535 195.445 ;
        RECT 32.705 195.235 33.035 195.615 ;
        RECT 33.280 195.115 33.510 195.445 ;
        RECT 32.360 194.875 32.990 195.045 ;
        RECT 29.240 193.500 29.590 194.750 ;
        RECT 32.820 194.705 32.990 194.875 ;
        RECT 32.275 194.025 32.640 194.705 ;
        RECT 32.820 194.375 33.170 194.705 ;
        RECT 32.820 193.855 32.990 194.375 ;
        RECT 32.360 193.685 32.990 193.855 ;
        RECT 33.340 193.825 33.510 195.115 ;
        RECT 33.710 194.005 33.990 195.280 ;
        RECT 34.215 194.255 34.485 195.280 ;
        RECT 34.945 195.235 35.275 195.615 ;
        RECT 35.445 195.360 35.780 195.405 ;
        RECT 34.175 194.085 34.485 194.255 ;
        RECT 34.215 194.005 34.485 194.085 ;
        RECT 34.675 194.005 35.015 195.035 ;
        RECT 35.445 194.895 35.785 195.360 ;
        RECT 35.185 194.375 35.445 194.705 ;
        RECT 35.185 193.825 35.355 194.375 ;
        RECT 35.615 194.205 35.785 194.895 ;
        RECT 35.955 194.845 38.545 195.615 ;
        RECT 39.175 194.890 39.465 195.615 ;
        RECT 39.635 195.070 44.980 195.615 ;
        RECT 45.155 195.070 50.500 195.615 ;
        RECT 50.680 195.215 51.015 195.615 ;
        RECT 35.955 194.325 37.165 194.845 ;
        RECT 14.795 193.065 20.140 193.500 ;
        RECT 20.315 193.065 25.660 193.500 ;
        RECT 25.835 193.065 31.180 193.500 ;
        RECT 32.360 193.235 32.535 193.685 ;
        RECT 33.340 193.655 35.355 193.825 ;
        RECT 32.705 193.065 33.035 193.505 ;
        RECT 33.340 193.235 33.510 193.655 ;
        RECT 33.745 193.065 34.415 193.475 ;
        RECT 34.630 193.235 34.800 193.655 ;
        RECT 35.000 193.065 35.330 193.475 ;
        RECT 35.525 193.235 35.785 194.205 ;
        RECT 37.335 194.155 38.545 194.675 ;
        RECT 41.220 194.240 41.560 195.070 ;
        RECT 35.955 193.065 38.545 194.155 ;
        RECT 39.175 193.065 39.465 194.230 ;
        RECT 43.040 193.500 43.390 194.750 ;
        RECT 46.740 194.240 47.080 195.070 ;
        RECT 51.185 195.045 51.390 195.445 ;
        RECT 51.600 195.135 51.875 195.615 ;
        RECT 52.085 195.115 52.345 195.445 ;
        RECT 50.705 194.875 51.390 195.045 ;
        RECT 48.560 193.500 48.910 194.750 ;
        RECT 50.705 193.845 51.045 194.875 ;
        RECT 51.215 194.205 51.465 194.705 ;
        RECT 51.645 194.375 52.005 194.955 ;
        RECT 52.175 194.205 52.345 195.115 ;
        RECT 52.515 194.845 54.185 195.615 ;
        RECT 54.865 194.960 55.195 195.395 ;
        RECT 55.365 195.005 55.535 195.615 ;
        RECT 54.815 194.875 55.195 194.960 ;
        RECT 55.705 194.875 56.035 195.400 ;
        RECT 56.295 195.085 56.505 195.615 ;
        RECT 56.780 195.165 57.565 195.335 ;
        RECT 57.735 195.165 58.140 195.335 ;
        RECT 52.515 194.325 53.265 194.845 ;
        RECT 54.815 194.835 55.040 194.875 ;
        RECT 51.215 194.035 52.345 194.205 ;
        RECT 53.435 194.155 54.185 194.675 ;
        RECT 50.705 193.670 51.370 193.845 ;
        RECT 39.635 193.065 44.980 193.500 ;
        RECT 45.155 193.065 50.500 193.500 ;
        RECT 50.680 193.065 51.015 193.490 ;
        RECT 51.185 193.265 51.370 193.670 ;
        RECT 51.575 193.065 51.905 193.845 ;
        RECT 52.075 193.265 52.345 194.035 ;
        RECT 52.515 193.065 54.185 194.155 ;
        RECT 54.815 194.255 54.985 194.835 ;
        RECT 55.705 194.705 55.905 194.875 ;
        RECT 56.780 194.705 56.950 195.165 ;
        RECT 55.155 194.375 55.905 194.705 ;
        RECT 56.075 194.375 56.950 194.705 ;
        RECT 54.815 194.205 55.030 194.255 ;
        RECT 54.815 194.125 55.205 194.205 ;
        RECT 54.875 193.280 55.205 194.125 ;
        RECT 55.715 194.170 55.905 194.375 ;
        RECT 55.375 193.065 55.545 194.075 ;
        RECT 55.715 193.795 56.610 194.170 ;
        RECT 55.715 193.235 56.055 193.795 ;
        RECT 56.285 193.065 56.600 193.565 ;
        RECT 56.780 193.535 56.950 194.375 ;
        RECT 57.120 194.665 57.585 194.995 ;
        RECT 57.970 194.935 58.140 195.165 ;
        RECT 58.320 195.115 58.690 195.615 ;
        RECT 59.010 195.165 59.685 195.335 ;
        RECT 59.880 195.165 60.215 195.335 ;
        RECT 57.120 193.705 57.440 194.665 ;
        RECT 57.970 194.635 58.800 194.935 ;
        RECT 57.610 193.735 57.800 194.455 ;
        RECT 57.970 193.565 58.140 194.635 ;
        RECT 58.600 194.605 58.800 194.635 ;
        RECT 58.310 194.385 58.480 194.455 ;
        RECT 59.010 194.385 59.180 195.165 ;
        RECT 60.045 195.025 60.215 195.165 ;
        RECT 60.385 195.155 60.635 195.615 ;
        RECT 58.310 194.215 59.180 194.385 ;
        RECT 59.350 194.745 59.875 194.965 ;
        RECT 60.045 194.895 60.270 195.025 ;
        RECT 58.310 194.125 58.820 194.215 ;
        RECT 56.780 193.365 57.665 193.535 ;
        RECT 57.890 193.235 58.140 193.565 ;
        RECT 58.310 193.065 58.480 193.865 ;
        RECT 58.650 193.510 58.820 194.125 ;
        RECT 59.350 194.045 59.520 194.745 ;
        RECT 58.990 193.680 59.520 194.045 ;
        RECT 59.690 193.980 59.930 194.575 ;
        RECT 60.100 193.790 60.270 194.895 ;
        RECT 60.440 194.035 60.720 194.985 ;
        RECT 59.965 193.660 60.270 193.790 ;
        RECT 58.650 193.340 59.755 193.510 ;
        RECT 59.965 193.235 60.215 193.660 ;
        RECT 60.385 193.065 60.650 193.525 ;
        RECT 60.890 193.235 61.075 195.355 ;
        RECT 61.245 195.235 61.575 195.615 ;
        RECT 61.745 195.065 61.915 195.355 ;
        RECT 61.250 194.895 61.915 195.065 ;
        RECT 62.185 195.085 62.515 195.445 ;
        RECT 62.685 195.255 63.015 195.615 ;
        RECT 63.215 195.085 63.545 195.445 ;
        RECT 61.250 193.905 61.480 194.895 ;
        RECT 62.185 194.875 63.545 195.085 ;
        RECT 64.055 194.855 64.765 195.445 ;
        RECT 64.935 194.890 65.225 195.615 ;
        RECT 65.485 195.065 65.655 195.355 ;
        RECT 65.825 195.235 66.155 195.615 ;
        RECT 65.485 194.895 66.150 195.065 ;
        RECT 61.650 194.075 62.000 194.725 ;
        RECT 62.175 194.375 62.485 194.705 ;
        RECT 62.695 194.375 63.070 194.705 ;
        RECT 63.390 194.375 63.885 194.705 ;
        RECT 61.250 193.735 61.915 193.905 ;
        RECT 61.245 193.065 61.575 193.565 ;
        RECT 61.745 193.235 61.915 193.735 ;
        RECT 62.185 193.065 62.515 194.125 ;
        RECT 62.695 193.450 62.865 194.375 ;
        RECT 63.035 193.885 63.365 194.105 ;
        RECT 63.560 194.085 63.885 194.375 ;
        RECT 64.060 194.085 64.390 194.625 ;
        RECT 64.560 193.885 64.765 194.855 ;
        RECT 63.035 193.655 64.765 193.885 ;
        RECT 63.035 193.255 63.365 193.655 ;
        RECT 63.535 193.065 63.865 193.425 ;
        RECT 64.065 193.235 64.765 193.655 ;
        RECT 64.935 193.065 65.225 194.230 ;
        RECT 65.400 194.075 65.750 194.725 ;
        RECT 65.920 193.905 66.150 194.895 ;
        RECT 65.485 193.735 66.150 193.905 ;
        RECT 65.485 193.235 65.655 193.735 ;
        RECT 65.825 193.065 66.155 193.565 ;
        RECT 66.325 193.235 66.510 195.355 ;
        RECT 66.765 195.155 67.015 195.615 ;
        RECT 67.185 195.165 67.520 195.335 ;
        RECT 67.715 195.165 68.390 195.335 ;
        RECT 67.185 195.025 67.355 195.165 ;
        RECT 66.680 194.035 66.960 194.985 ;
        RECT 67.130 194.895 67.355 195.025 ;
        RECT 67.130 193.790 67.300 194.895 ;
        RECT 67.525 194.745 68.050 194.965 ;
        RECT 67.470 193.980 67.710 194.575 ;
        RECT 67.880 194.045 68.050 194.745 ;
        RECT 68.220 194.385 68.390 195.165 ;
        RECT 68.710 195.115 69.080 195.615 ;
        RECT 69.260 195.165 69.665 195.335 ;
        RECT 69.835 195.165 70.620 195.335 ;
        RECT 69.260 194.935 69.430 195.165 ;
        RECT 68.600 194.635 69.430 194.935 ;
        RECT 69.815 194.665 70.280 194.995 ;
        RECT 68.600 194.605 68.800 194.635 ;
        RECT 68.920 194.385 69.090 194.455 ;
        RECT 68.220 194.215 69.090 194.385 ;
        RECT 68.580 194.125 69.090 194.215 ;
        RECT 67.130 193.660 67.435 193.790 ;
        RECT 67.880 193.680 68.410 194.045 ;
        RECT 66.750 193.065 67.015 193.525 ;
        RECT 67.185 193.235 67.435 193.660 ;
        RECT 68.580 193.510 68.750 194.125 ;
        RECT 67.645 193.340 68.750 193.510 ;
        RECT 68.920 193.065 69.090 193.865 ;
        RECT 69.260 193.565 69.430 194.635 ;
        RECT 69.600 193.735 69.790 194.455 ;
        RECT 69.960 193.705 70.280 194.665 ;
        RECT 70.450 194.705 70.620 195.165 ;
        RECT 70.895 195.085 71.105 195.615 ;
        RECT 71.365 194.875 71.695 195.400 ;
        RECT 71.865 195.005 72.035 195.615 ;
        RECT 72.205 194.960 72.535 195.395 ;
        RECT 72.205 194.875 72.585 194.960 ;
        RECT 71.495 194.705 71.695 194.875 ;
        RECT 72.360 194.835 72.585 194.875 ;
        RECT 70.450 194.375 71.325 194.705 ;
        RECT 71.495 194.375 72.245 194.705 ;
        RECT 69.260 193.235 69.510 193.565 ;
        RECT 70.450 193.535 70.620 194.375 ;
        RECT 71.495 194.170 71.685 194.375 ;
        RECT 72.415 194.255 72.585 194.835 ;
        RECT 72.370 194.205 72.585 194.255 ;
        RECT 70.790 193.795 71.685 194.170 ;
        RECT 72.195 194.125 72.585 194.205 ;
        RECT 72.755 194.890 73.015 195.445 ;
        RECT 73.185 195.170 73.615 195.615 ;
        RECT 73.850 195.045 74.020 195.445 ;
        RECT 74.190 195.215 74.910 195.615 ;
        RECT 72.755 194.175 72.930 194.890 ;
        RECT 73.850 194.875 74.730 195.045 ;
        RECT 75.080 195.000 75.250 195.445 ;
        RECT 75.825 195.105 76.225 195.615 ;
        RECT 73.100 194.375 73.355 194.705 ;
        RECT 69.735 193.365 70.620 193.535 ;
        RECT 70.800 193.065 71.115 193.565 ;
        RECT 71.345 193.235 71.685 193.795 ;
        RECT 71.855 193.065 72.025 194.075 ;
        RECT 72.195 193.280 72.525 194.125 ;
        RECT 72.755 193.235 73.015 194.175 ;
        RECT 73.185 193.895 73.355 194.375 ;
        RECT 73.580 194.085 73.910 194.705 ;
        RECT 74.080 194.325 74.370 194.705 ;
        RECT 74.560 194.155 74.730 194.875 ;
        RECT 74.210 193.985 74.730 194.155 ;
        RECT 74.900 194.830 75.250 195.000 ;
        RECT 73.185 193.725 73.945 193.895 ;
        RECT 74.210 193.795 74.380 193.985 ;
        RECT 74.900 193.805 75.070 194.830 ;
        RECT 75.490 194.345 75.750 194.935 ;
        RECT 75.270 194.045 75.750 194.345 ;
        RECT 75.950 194.045 76.210 194.935 ;
        RECT 76.435 194.875 76.820 195.445 ;
        RECT 76.990 195.155 77.315 195.615 ;
        RECT 77.835 194.985 78.115 195.445 ;
        RECT 76.435 194.205 76.715 194.875 ;
        RECT 76.990 194.815 78.115 194.985 ;
        RECT 76.990 194.705 77.440 194.815 ;
        RECT 76.885 194.375 77.440 194.705 ;
        RECT 78.305 194.645 78.705 195.445 ;
        RECT 79.105 195.155 79.375 195.615 ;
        RECT 79.545 194.985 79.830 195.445 ;
        RECT 73.775 193.500 73.945 193.725 ;
        RECT 74.660 193.635 75.070 193.805 ;
        RECT 75.245 193.695 76.185 193.865 ;
        RECT 74.660 193.500 74.915 193.635 ;
        RECT 73.185 193.065 73.515 193.465 ;
        RECT 73.775 193.330 74.915 193.500 ;
        RECT 75.245 193.445 75.415 193.695 ;
        RECT 74.660 193.235 74.915 193.330 ;
        RECT 75.085 193.275 75.415 193.445 ;
        RECT 75.585 193.065 75.835 193.525 ;
        RECT 76.005 193.235 76.185 193.695 ;
        RECT 76.435 193.235 76.820 194.205 ;
        RECT 76.990 193.915 77.440 194.375 ;
        RECT 77.610 194.085 78.705 194.645 ;
        RECT 76.990 193.695 78.115 193.915 ;
        RECT 76.990 193.065 77.315 193.525 ;
        RECT 77.835 193.235 78.115 193.695 ;
        RECT 78.305 193.235 78.705 194.085 ;
        RECT 78.875 194.815 79.830 194.985 ;
        RECT 78.875 193.915 79.085 194.815 ;
        RECT 80.585 194.805 80.855 195.615 ;
        RECT 81.025 194.805 81.355 195.445 ;
        RECT 81.525 194.805 81.765 195.615 ;
        RECT 81.955 194.845 85.465 195.615 ;
        RECT 86.095 194.875 86.480 195.445 ;
        RECT 86.650 195.155 86.975 195.615 ;
        RECT 87.495 194.985 87.775 195.445 ;
        RECT 79.255 194.085 79.945 194.645 ;
        RECT 80.575 194.375 80.925 194.625 ;
        RECT 81.095 194.205 81.265 194.805 ;
        RECT 81.435 194.375 81.785 194.625 ;
        RECT 81.955 194.325 83.605 194.845 ;
        RECT 78.875 193.695 79.830 193.915 ;
        RECT 79.105 193.065 79.375 193.525 ;
        RECT 79.545 193.235 79.830 193.695 ;
        RECT 80.585 193.065 80.915 194.205 ;
        RECT 81.095 194.035 81.775 194.205 ;
        RECT 83.775 194.155 85.465 194.675 ;
        RECT 81.445 193.250 81.775 194.035 ;
        RECT 81.955 193.065 85.465 194.155 ;
        RECT 86.095 194.205 86.375 194.875 ;
        RECT 86.650 194.815 87.775 194.985 ;
        RECT 86.650 194.705 87.100 194.815 ;
        RECT 86.545 194.375 87.100 194.705 ;
        RECT 87.965 194.645 88.365 195.445 ;
        RECT 88.765 195.155 89.035 195.615 ;
        RECT 89.205 194.985 89.490 195.445 ;
        RECT 86.095 193.235 86.480 194.205 ;
        RECT 86.650 193.915 87.100 194.375 ;
        RECT 87.270 194.085 88.365 194.645 ;
        RECT 86.650 193.695 87.775 193.915 ;
        RECT 86.650 193.065 86.975 193.525 ;
        RECT 87.495 193.235 87.775 193.695 ;
        RECT 87.965 193.235 88.365 194.085 ;
        RECT 88.535 194.815 89.490 194.985 ;
        RECT 90.695 194.890 90.985 195.615 ;
        RECT 91.205 194.960 91.535 195.395 ;
        RECT 91.705 195.005 91.875 195.615 ;
        RECT 91.155 194.875 91.535 194.960 ;
        RECT 92.045 194.875 92.375 195.400 ;
        RECT 92.635 195.085 92.845 195.615 ;
        RECT 93.120 195.165 93.905 195.335 ;
        RECT 94.075 195.165 94.480 195.335 ;
        RECT 91.155 194.835 91.380 194.875 ;
        RECT 88.535 193.915 88.745 194.815 ;
        RECT 88.915 194.085 89.605 194.645 ;
        RECT 91.155 194.255 91.325 194.835 ;
        RECT 92.045 194.705 92.245 194.875 ;
        RECT 93.120 194.705 93.290 195.165 ;
        RECT 91.495 194.375 92.245 194.705 ;
        RECT 92.415 194.375 93.290 194.705 ;
        RECT 88.535 193.695 89.490 193.915 ;
        RECT 88.765 193.065 89.035 193.525 ;
        RECT 89.205 193.235 89.490 193.695 ;
        RECT 90.695 193.065 90.985 194.230 ;
        RECT 91.155 194.205 91.370 194.255 ;
        RECT 91.155 194.125 91.545 194.205 ;
        RECT 91.215 193.280 91.545 194.125 ;
        RECT 92.055 194.170 92.245 194.375 ;
        RECT 91.715 193.065 91.885 194.075 ;
        RECT 92.055 193.795 92.950 194.170 ;
        RECT 92.055 193.235 92.395 193.795 ;
        RECT 92.625 193.065 92.940 193.565 ;
        RECT 93.120 193.535 93.290 194.375 ;
        RECT 93.460 194.665 93.925 194.995 ;
        RECT 94.310 194.935 94.480 195.165 ;
        RECT 94.660 195.115 95.030 195.615 ;
        RECT 95.350 195.165 96.025 195.335 ;
        RECT 96.220 195.165 96.555 195.335 ;
        RECT 93.460 193.705 93.780 194.665 ;
        RECT 94.310 194.635 95.140 194.935 ;
        RECT 93.950 193.735 94.140 194.455 ;
        RECT 94.310 193.565 94.480 194.635 ;
        RECT 94.940 194.605 95.140 194.635 ;
        RECT 94.650 194.385 94.820 194.455 ;
        RECT 95.350 194.385 95.520 195.165 ;
        RECT 96.385 195.025 96.555 195.165 ;
        RECT 96.725 195.155 96.975 195.615 ;
        RECT 94.650 194.215 95.520 194.385 ;
        RECT 95.690 194.745 96.215 194.965 ;
        RECT 96.385 194.895 96.610 195.025 ;
        RECT 94.650 194.125 95.160 194.215 ;
        RECT 93.120 193.365 94.005 193.535 ;
        RECT 94.230 193.235 94.480 193.565 ;
        RECT 94.650 193.065 94.820 193.865 ;
        RECT 94.990 193.510 95.160 194.125 ;
        RECT 95.690 194.045 95.860 194.745 ;
        RECT 95.330 193.680 95.860 194.045 ;
        RECT 96.030 193.980 96.270 194.575 ;
        RECT 96.440 193.790 96.610 194.895 ;
        RECT 96.780 194.035 97.060 194.985 ;
        RECT 96.305 193.660 96.610 193.790 ;
        RECT 94.990 193.340 96.095 193.510 ;
        RECT 96.305 193.235 96.555 193.660 ;
        RECT 96.725 193.065 96.990 193.525 ;
        RECT 97.230 193.235 97.415 195.355 ;
        RECT 97.585 195.235 97.915 195.615 ;
        RECT 98.085 195.065 98.255 195.355 ;
        RECT 97.590 194.895 98.255 195.065 ;
        RECT 98.630 194.985 98.915 195.445 ;
        RECT 99.085 195.155 99.355 195.615 ;
        RECT 97.590 193.905 97.820 194.895 ;
        RECT 98.630 194.815 99.585 194.985 ;
        RECT 97.990 194.075 98.340 194.725 ;
        RECT 98.515 194.085 99.205 194.645 ;
        RECT 99.375 193.915 99.585 194.815 ;
        RECT 97.590 193.735 98.255 193.905 ;
        RECT 97.585 193.065 97.915 193.565 ;
        RECT 98.085 193.235 98.255 193.735 ;
        RECT 98.630 193.695 99.585 193.915 ;
        RECT 99.755 194.645 100.155 195.445 ;
        RECT 100.345 194.985 100.625 195.445 ;
        RECT 101.145 195.155 101.470 195.615 ;
        RECT 100.345 194.815 101.470 194.985 ;
        RECT 101.640 194.875 102.025 195.445 ;
        RECT 103.205 195.065 103.375 195.355 ;
        RECT 103.545 195.235 103.875 195.615 ;
        RECT 103.205 194.895 103.870 195.065 ;
        RECT 101.020 194.705 101.470 194.815 ;
        RECT 99.755 194.085 100.850 194.645 ;
        RECT 101.020 194.375 101.575 194.705 ;
        RECT 98.630 193.235 98.915 193.695 ;
        RECT 99.085 193.065 99.355 193.525 ;
        RECT 99.755 193.235 100.155 194.085 ;
        RECT 101.020 193.915 101.470 194.375 ;
        RECT 101.745 194.205 102.025 194.875 ;
        RECT 100.345 193.695 101.470 193.915 ;
        RECT 100.345 193.235 100.625 193.695 ;
        RECT 101.145 193.065 101.470 193.525 ;
        RECT 101.640 193.235 102.025 194.205 ;
        RECT 103.120 194.075 103.470 194.725 ;
        RECT 103.640 193.905 103.870 194.895 ;
        RECT 103.205 193.735 103.870 193.905 ;
        RECT 103.205 193.235 103.375 193.735 ;
        RECT 103.545 193.065 103.875 193.565 ;
        RECT 104.045 193.235 104.230 195.355 ;
        RECT 104.485 195.155 104.735 195.615 ;
        RECT 104.905 195.165 105.240 195.335 ;
        RECT 105.435 195.165 106.110 195.335 ;
        RECT 104.905 195.025 105.075 195.165 ;
        RECT 104.400 194.035 104.680 194.985 ;
        RECT 104.850 194.895 105.075 195.025 ;
        RECT 104.850 193.790 105.020 194.895 ;
        RECT 105.245 194.745 105.770 194.965 ;
        RECT 105.190 193.980 105.430 194.575 ;
        RECT 105.600 194.045 105.770 194.745 ;
        RECT 105.940 194.385 106.110 195.165 ;
        RECT 106.430 195.115 106.800 195.615 ;
        RECT 106.980 195.165 107.385 195.335 ;
        RECT 107.555 195.165 108.340 195.335 ;
        RECT 106.980 194.935 107.150 195.165 ;
        RECT 106.320 194.635 107.150 194.935 ;
        RECT 107.535 194.665 108.000 194.995 ;
        RECT 106.320 194.605 106.520 194.635 ;
        RECT 106.640 194.385 106.810 194.455 ;
        RECT 105.940 194.215 106.810 194.385 ;
        RECT 106.300 194.125 106.810 194.215 ;
        RECT 104.850 193.660 105.155 193.790 ;
        RECT 105.600 193.680 106.130 194.045 ;
        RECT 104.470 193.065 104.735 193.525 ;
        RECT 104.905 193.235 105.155 193.660 ;
        RECT 106.300 193.510 106.470 194.125 ;
        RECT 105.365 193.340 106.470 193.510 ;
        RECT 106.640 193.065 106.810 193.865 ;
        RECT 106.980 193.565 107.150 194.635 ;
        RECT 107.320 193.735 107.510 194.455 ;
        RECT 107.680 193.705 108.000 194.665 ;
        RECT 108.170 194.705 108.340 195.165 ;
        RECT 108.615 195.085 108.825 195.615 ;
        RECT 109.085 194.875 109.415 195.400 ;
        RECT 109.585 195.005 109.755 195.615 ;
        RECT 109.925 194.960 110.255 195.395 ;
        RECT 109.925 194.875 110.305 194.960 ;
        RECT 109.215 194.705 109.415 194.875 ;
        RECT 110.080 194.835 110.305 194.875 ;
        RECT 108.170 194.375 109.045 194.705 ;
        RECT 109.215 194.375 109.965 194.705 ;
        RECT 106.980 193.235 107.230 193.565 ;
        RECT 108.170 193.535 108.340 194.375 ;
        RECT 109.215 194.170 109.405 194.375 ;
        RECT 110.135 194.255 110.305 194.835 ;
        RECT 111.210 194.805 111.455 195.410 ;
        RECT 111.675 195.080 112.185 195.615 ;
        RECT 110.090 194.205 110.305 194.255 ;
        RECT 108.510 193.795 109.405 194.170 ;
        RECT 109.915 194.125 110.305 194.205 ;
        RECT 110.935 194.635 112.165 194.805 ;
        RECT 107.455 193.365 108.340 193.535 ;
        RECT 108.520 193.065 108.835 193.565 ;
        RECT 109.065 193.235 109.405 193.795 ;
        RECT 109.575 193.065 109.745 194.075 ;
        RECT 109.915 193.280 110.245 194.125 ;
        RECT 110.935 193.825 111.275 194.635 ;
        RECT 111.445 194.070 112.195 194.260 ;
        RECT 110.935 193.415 111.450 193.825 ;
        RECT 111.685 193.065 111.855 193.825 ;
        RECT 112.025 193.405 112.195 194.070 ;
        RECT 112.365 194.085 112.555 195.445 ;
        RECT 112.725 194.595 113.000 195.445 ;
        RECT 113.190 195.080 113.720 195.445 ;
        RECT 114.145 195.215 114.475 195.615 ;
        RECT 113.545 195.045 113.720 195.080 ;
        RECT 112.725 194.425 113.005 194.595 ;
        RECT 112.725 194.285 113.000 194.425 ;
        RECT 113.205 194.085 113.375 194.885 ;
        RECT 112.365 193.915 113.375 194.085 ;
        RECT 113.545 194.875 114.475 195.045 ;
        RECT 114.645 194.875 114.900 195.445 ;
        RECT 113.545 193.745 113.715 194.875 ;
        RECT 114.305 194.705 114.475 194.875 ;
        RECT 112.590 193.575 113.715 193.745 ;
        RECT 113.885 194.375 114.080 194.705 ;
        RECT 114.305 194.375 114.560 194.705 ;
        RECT 113.885 193.405 114.055 194.375 ;
        RECT 114.730 194.205 114.900 194.875 ;
        RECT 115.075 194.865 116.285 195.615 ;
        RECT 116.455 194.890 116.745 195.615 ;
        RECT 116.915 195.070 122.260 195.615 ;
        RECT 122.435 195.070 127.780 195.615 ;
        RECT 127.955 195.070 133.300 195.615 ;
        RECT 115.075 194.325 115.595 194.865 ;
        RECT 112.025 193.235 114.055 193.405 ;
        RECT 114.225 193.065 114.395 194.205 ;
        RECT 114.565 193.235 114.900 194.205 ;
        RECT 115.765 194.155 116.285 194.695 ;
        RECT 118.500 194.240 118.840 195.070 ;
        RECT 115.075 193.065 116.285 194.155 ;
        RECT 116.455 193.065 116.745 194.230 ;
        RECT 120.320 193.500 120.670 194.750 ;
        RECT 124.020 194.240 124.360 195.070 ;
        RECT 125.840 193.500 126.190 194.750 ;
        RECT 129.540 194.240 129.880 195.070 ;
        RECT 133.475 194.845 136.985 195.615 ;
        RECT 137.615 194.865 138.825 195.615 ;
        RECT 131.360 193.500 131.710 194.750 ;
        RECT 133.475 194.325 135.125 194.845 ;
        RECT 135.295 194.155 136.985 194.675 ;
        RECT 116.915 193.065 122.260 193.500 ;
        RECT 122.435 193.065 127.780 193.500 ;
        RECT 127.955 193.065 133.300 193.500 ;
        RECT 133.475 193.065 136.985 194.155 ;
        RECT 137.615 194.155 138.135 194.695 ;
        RECT 138.305 194.325 138.825 194.865 ;
        RECT 137.615 193.065 138.825 194.155 ;
        RECT 13.330 192.895 138.910 193.065 ;
        RECT 13.415 191.805 14.625 192.895 ;
        RECT 14.795 191.805 18.305 192.895 ;
        RECT 19.025 192.225 19.195 192.725 ;
        RECT 19.365 192.395 19.695 192.895 ;
        RECT 19.025 192.055 19.690 192.225 ;
        RECT 13.415 191.095 13.935 191.635 ;
        RECT 14.105 191.265 14.625 191.805 ;
        RECT 14.795 191.115 16.445 191.635 ;
        RECT 16.615 191.285 18.305 191.805 ;
        RECT 18.940 191.235 19.290 191.885 ;
        RECT 13.415 190.345 14.625 191.095 ;
        RECT 14.795 190.345 18.305 191.115 ;
        RECT 19.460 191.065 19.690 192.055 ;
        RECT 19.025 190.895 19.690 191.065 ;
        RECT 19.025 190.605 19.195 190.895 ;
        RECT 19.365 190.345 19.695 190.725 ;
        RECT 19.865 190.605 20.050 192.725 ;
        RECT 20.290 192.435 20.555 192.895 ;
        RECT 20.725 192.300 20.975 192.725 ;
        RECT 21.185 192.450 22.290 192.620 ;
        RECT 20.670 192.170 20.975 192.300 ;
        RECT 20.220 190.975 20.500 191.925 ;
        RECT 20.670 191.065 20.840 192.170 ;
        RECT 21.010 191.385 21.250 191.980 ;
        RECT 21.420 191.915 21.950 192.280 ;
        RECT 21.420 191.215 21.590 191.915 ;
        RECT 22.120 191.835 22.290 192.450 ;
        RECT 22.460 192.095 22.630 192.895 ;
        RECT 22.800 192.395 23.050 192.725 ;
        RECT 23.275 192.425 24.160 192.595 ;
        RECT 22.120 191.745 22.630 191.835 ;
        RECT 20.670 190.935 20.895 191.065 ;
        RECT 21.065 190.995 21.590 191.215 ;
        RECT 21.760 191.575 22.630 191.745 ;
        RECT 20.305 190.345 20.555 190.805 ;
        RECT 20.725 190.795 20.895 190.935 ;
        RECT 21.760 190.795 21.930 191.575 ;
        RECT 22.460 191.505 22.630 191.575 ;
        RECT 22.140 191.325 22.340 191.355 ;
        RECT 22.800 191.325 22.970 192.395 ;
        RECT 23.140 191.505 23.330 192.225 ;
        RECT 22.140 191.025 22.970 191.325 ;
        RECT 23.500 191.295 23.820 192.255 ;
        RECT 20.725 190.625 21.060 190.795 ;
        RECT 21.255 190.625 21.930 190.795 ;
        RECT 22.250 190.345 22.620 190.845 ;
        RECT 22.800 190.795 22.970 191.025 ;
        RECT 23.355 190.965 23.820 191.295 ;
        RECT 23.990 191.585 24.160 192.425 ;
        RECT 24.340 192.395 24.655 192.895 ;
        RECT 24.885 192.165 25.225 192.725 ;
        RECT 24.330 191.790 25.225 192.165 ;
        RECT 25.395 191.885 25.565 192.895 ;
        RECT 25.035 191.585 25.225 191.790 ;
        RECT 25.735 191.835 26.065 192.680 ;
        RECT 25.735 191.755 26.125 191.835 ;
        RECT 25.910 191.705 26.125 191.755 ;
        RECT 26.295 191.730 26.585 192.895 ;
        RECT 26.755 191.805 28.425 192.895 ;
        RECT 29.140 192.275 29.315 192.725 ;
        RECT 29.485 192.455 29.815 192.895 ;
        RECT 30.120 192.305 30.290 192.725 ;
        RECT 30.525 192.485 31.195 192.895 ;
        RECT 31.410 192.305 31.580 192.725 ;
        RECT 31.780 192.485 32.110 192.895 ;
        RECT 29.140 192.105 29.770 192.275 ;
        RECT 23.990 191.255 24.865 191.585 ;
        RECT 25.035 191.255 25.785 191.585 ;
        RECT 23.990 190.795 24.160 191.255 ;
        RECT 25.035 191.085 25.235 191.255 ;
        RECT 25.955 191.125 26.125 191.705 ;
        RECT 25.900 191.085 26.125 191.125 ;
        RECT 22.800 190.625 23.205 190.795 ;
        RECT 23.375 190.625 24.160 190.795 ;
        RECT 24.435 190.345 24.645 190.875 ;
        RECT 24.905 190.560 25.235 191.085 ;
        RECT 25.745 191.000 26.125 191.085 ;
        RECT 26.755 191.115 27.505 191.635 ;
        RECT 27.675 191.285 28.425 191.805 ;
        RECT 29.055 191.255 29.420 191.935 ;
        RECT 29.600 191.585 29.770 192.105 ;
        RECT 30.120 192.135 32.135 192.305 ;
        RECT 29.600 191.255 29.950 191.585 ;
        RECT 25.405 190.345 25.575 190.955 ;
        RECT 25.745 190.565 26.075 191.000 ;
        RECT 26.295 190.345 26.585 191.070 ;
        RECT 26.755 190.345 28.425 191.115 ;
        RECT 29.600 191.085 29.770 191.255 ;
        RECT 29.140 190.915 29.770 191.085 ;
        RECT 29.140 190.515 29.315 190.915 ;
        RECT 30.120 190.845 30.290 192.135 ;
        RECT 29.485 190.345 29.815 190.725 ;
        RECT 30.060 190.515 30.290 190.845 ;
        RECT 30.490 190.680 30.770 191.955 ;
        RECT 30.995 191.875 31.265 191.955 ;
        RECT 30.955 191.705 31.265 191.875 ;
        RECT 30.995 190.680 31.265 191.705 ;
        RECT 31.455 190.925 31.795 191.955 ;
        RECT 31.965 191.585 32.135 192.135 ;
        RECT 32.305 191.755 32.565 192.725 ;
        RECT 32.825 192.225 32.995 192.725 ;
        RECT 33.165 192.395 33.495 192.895 ;
        RECT 32.825 192.055 33.490 192.225 ;
        RECT 31.965 191.255 32.225 191.585 ;
        RECT 32.395 191.065 32.565 191.755 ;
        RECT 32.740 191.235 33.090 191.885 ;
        RECT 33.260 191.065 33.490 192.055 ;
        RECT 31.725 190.345 32.055 190.725 ;
        RECT 32.225 190.600 32.565 191.065 ;
        RECT 32.825 190.895 33.490 191.065 ;
        RECT 32.825 190.605 32.995 190.895 ;
        RECT 32.225 190.555 32.560 190.600 ;
        RECT 33.165 190.345 33.495 190.725 ;
        RECT 33.665 190.605 33.850 192.725 ;
        RECT 34.090 192.435 34.355 192.895 ;
        RECT 34.525 192.300 34.775 192.725 ;
        RECT 34.985 192.450 36.090 192.620 ;
        RECT 34.470 192.170 34.775 192.300 ;
        RECT 34.020 190.975 34.300 191.925 ;
        RECT 34.470 191.065 34.640 192.170 ;
        RECT 34.810 191.385 35.050 191.980 ;
        RECT 35.220 191.915 35.750 192.280 ;
        RECT 35.220 191.215 35.390 191.915 ;
        RECT 35.920 191.835 36.090 192.450 ;
        RECT 36.260 192.095 36.430 192.895 ;
        RECT 36.600 192.395 36.850 192.725 ;
        RECT 37.075 192.425 37.960 192.595 ;
        RECT 35.920 191.745 36.430 191.835 ;
        RECT 34.470 190.935 34.695 191.065 ;
        RECT 34.865 190.995 35.390 191.215 ;
        RECT 35.560 191.575 36.430 191.745 ;
        RECT 34.105 190.345 34.355 190.805 ;
        RECT 34.525 190.795 34.695 190.935 ;
        RECT 35.560 190.795 35.730 191.575 ;
        RECT 36.260 191.505 36.430 191.575 ;
        RECT 35.940 191.325 36.140 191.355 ;
        RECT 36.600 191.325 36.770 192.395 ;
        RECT 36.940 191.505 37.130 192.225 ;
        RECT 35.940 191.025 36.770 191.325 ;
        RECT 37.300 191.295 37.620 192.255 ;
        RECT 34.525 190.625 34.860 190.795 ;
        RECT 35.055 190.625 35.730 190.795 ;
        RECT 36.050 190.345 36.420 190.845 ;
        RECT 36.600 190.795 36.770 191.025 ;
        RECT 37.155 190.965 37.620 191.295 ;
        RECT 37.790 191.585 37.960 192.425 ;
        RECT 38.140 192.395 38.455 192.895 ;
        RECT 38.685 192.165 39.025 192.725 ;
        RECT 38.130 191.790 39.025 192.165 ;
        RECT 39.195 191.885 39.365 192.895 ;
        RECT 38.835 191.585 39.025 191.790 ;
        RECT 39.535 191.835 39.865 192.680 ;
        RECT 39.535 191.755 39.925 191.835 ;
        RECT 40.095 191.805 43.605 192.895 ;
        RECT 43.865 192.225 44.035 192.725 ;
        RECT 44.205 192.395 44.535 192.895 ;
        RECT 43.865 192.055 44.530 192.225 ;
        RECT 39.710 191.705 39.925 191.755 ;
        RECT 37.790 191.255 38.665 191.585 ;
        RECT 38.835 191.255 39.585 191.585 ;
        RECT 37.790 190.795 37.960 191.255 ;
        RECT 38.835 191.085 39.035 191.255 ;
        RECT 39.755 191.125 39.925 191.705 ;
        RECT 39.700 191.085 39.925 191.125 ;
        RECT 36.600 190.625 37.005 190.795 ;
        RECT 37.175 190.625 37.960 190.795 ;
        RECT 38.235 190.345 38.445 190.875 ;
        RECT 38.705 190.560 39.035 191.085 ;
        RECT 39.545 191.000 39.925 191.085 ;
        RECT 40.095 191.115 41.745 191.635 ;
        RECT 41.915 191.285 43.605 191.805 ;
        RECT 43.780 191.235 44.130 191.885 ;
        RECT 39.205 190.345 39.375 190.955 ;
        RECT 39.545 190.565 39.875 191.000 ;
        RECT 40.095 190.345 43.605 191.115 ;
        RECT 44.300 191.065 44.530 192.055 ;
        RECT 43.865 190.895 44.530 191.065 ;
        RECT 43.865 190.605 44.035 190.895 ;
        RECT 44.205 190.345 44.535 190.725 ;
        RECT 44.705 190.605 44.890 192.725 ;
        RECT 45.130 192.435 45.395 192.895 ;
        RECT 45.565 192.300 45.815 192.725 ;
        RECT 46.025 192.450 47.130 192.620 ;
        RECT 45.510 192.170 45.815 192.300 ;
        RECT 45.060 190.975 45.340 191.925 ;
        RECT 45.510 191.065 45.680 192.170 ;
        RECT 45.850 191.385 46.090 191.980 ;
        RECT 46.260 191.915 46.790 192.280 ;
        RECT 46.260 191.215 46.430 191.915 ;
        RECT 46.960 191.835 47.130 192.450 ;
        RECT 47.300 192.095 47.470 192.895 ;
        RECT 47.640 192.395 47.890 192.725 ;
        RECT 48.115 192.425 49.000 192.595 ;
        RECT 46.960 191.745 47.470 191.835 ;
        RECT 45.510 190.935 45.735 191.065 ;
        RECT 45.905 190.995 46.430 191.215 ;
        RECT 46.600 191.575 47.470 191.745 ;
        RECT 45.145 190.345 45.395 190.805 ;
        RECT 45.565 190.795 45.735 190.935 ;
        RECT 46.600 190.795 46.770 191.575 ;
        RECT 47.300 191.505 47.470 191.575 ;
        RECT 46.980 191.325 47.180 191.355 ;
        RECT 47.640 191.325 47.810 192.395 ;
        RECT 47.980 191.505 48.170 192.225 ;
        RECT 46.980 191.025 47.810 191.325 ;
        RECT 48.340 191.295 48.660 192.255 ;
        RECT 45.565 190.625 45.900 190.795 ;
        RECT 46.095 190.625 46.770 190.795 ;
        RECT 47.090 190.345 47.460 190.845 ;
        RECT 47.640 190.795 47.810 191.025 ;
        RECT 48.195 190.965 48.660 191.295 ;
        RECT 48.830 191.585 49.000 192.425 ;
        RECT 49.180 192.395 49.495 192.895 ;
        RECT 49.725 192.165 50.065 192.725 ;
        RECT 49.170 191.790 50.065 192.165 ;
        RECT 50.235 191.885 50.405 192.895 ;
        RECT 49.875 191.585 50.065 191.790 ;
        RECT 50.575 191.835 50.905 192.680 ;
        RECT 50.575 191.755 50.965 191.835 ;
        RECT 50.750 191.705 50.965 191.755 ;
        RECT 52.055 191.730 52.345 192.895 ;
        RECT 52.605 192.225 52.775 192.725 ;
        RECT 52.945 192.395 53.275 192.895 ;
        RECT 52.605 192.055 53.270 192.225 ;
        RECT 48.830 191.255 49.705 191.585 ;
        RECT 49.875 191.255 50.625 191.585 ;
        RECT 48.830 190.795 49.000 191.255 ;
        RECT 49.875 191.085 50.075 191.255 ;
        RECT 50.795 191.125 50.965 191.705 ;
        RECT 52.520 191.235 52.870 191.885 ;
        RECT 50.740 191.085 50.965 191.125 ;
        RECT 47.640 190.625 48.045 190.795 ;
        RECT 48.215 190.625 49.000 190.795 ;
        RECT 49.275 190.345 49.485 190.875 ;
        RECT 49.745 190.560 50.075 191.085 ;
        RECT 50.585 191.000 50.965 191.085 ;
        RECT 50.245 190.345 50.415 190.955 ;
        RECT 50.585 190.565 50.915 191.000 ;
        RECT 52.055 190.345 52.345 191.070 ;
        RECT 53.040 191.065 53.270 192.055 ;
        RECT 52.605 190.895 53.270 191.065 ;
        RECT 52.605 190.605 52.775 190.895 ;
        RECT 52.945 190.345 53.275 190.725 ;
        RECT 53.445 190.605 53.630 192.725 ;
        RECT 53.870 192.435 54.135 192.895 ;
        RECT 54.305 192.300 54.555 192.725 ;
        RECT 54.765 192.450 55.870 192.620 ;
        RECT 54.250 192.170 54.555 192.300 ;
        RECT 53.800 190.975 54.080 191.925 ;
        RECT 54.250 191.065 54.420 192.170 ;
        RECT 54.590 191.385 54.830 191.980 ;
        RECT 55.000 191.915 55.530 192.280 ;
        RECT 55.000 191.215 55.170 191.915 ;
        RECT 55.700 191.835 55.870 192.450 ;
        RECT 56.040 192.095 56.210 192.895 ;
        RECT 56.380 192.395 56.630 192.725 ;
        RECT 56.855 192.425 57.740 192.595 ;
        RECT 55.700 191.745 56.210 191.835 ;
        RECT 54.250 190.935 54.475 191.065 ;
        RECT 54.645 190.995 55.170 191.215 ;
        RECT 55.340 191.575 56.210 191.745 ;
        RECT 53.885 190.345 54.135 190.805 ;
        RECT 54.305 190.795 54.475 190.935 ;
        RECT 55.340 190.795 55.510 191.575 ;
        RECT 56.040 191.505 56.210 191.575 ;
        RECT 55.720 191.325 55.920 191.355 ;
        RECT 56.380 191.325 56.550 192.395 ;
        RECT 56.720 191.505 56.910 192.225 ;
        RECT 55.720 191.025 56.550 191.325 ;
        RECT 57.080 191.295 57.400 192.255 ;
        RECT 54.305 190.625 54.640 190.795 ;
        RECT 54.835 190.625 55.510 190.795 ;
        RECT 55.830 190.345 56.200 190.845 ;
        RECT 56.380 190.795 56.550 191.025 ;
        RECT 56.935 190.965 57.400 191.295 ;
        RECT 57.570 191.585 57.740 192.425 ;
        RECT 57.920 192.395 58.235 192.895 ;
        RECT 58.465 192.165 58.805 192.725 ;
        RECT 57.910 191.790 58.805 192.165 ;
        RECT 58.975 191.885 59.145 192.895 ;
        RECT 58.615 191.585 58.805 191.790 ;
        RECT 59.315 191.835 59.645 192.680 ;
        RECT 59.315 191.755 59.705 191.835 ;
        RECT 59.490 191.705 59.705 191.755 ;
        RECT 57.570 191.255 58.445 191.585 ;
        RECT 58.615 191.255 59.365 191.585 ;
        RECT 57.570 190.795 57.740 191.255 ;
        RECT 58.615 191.085 58.815 191.255 ;
        RECT 59.535 191.125 59.705 191.705 ;
        RECT 59.480 191.085 59.705 191.125 ;
        RECT 56.380 190.625 56.785 190.795 ;
        RECT 56.955 190.625 57.740 190.795 ;
        RECT 58.015 190.345 58.225 190.875 ;
        RECT 58.485 190.560 58.815 191.085 ;
        RECT 59.325 191.000 59.705 191.085 ;
        RECT 60.335 191.785 60.595 192.725 ;
        RECT 60.765 192.495 61.095 192.895 ;
        RECT 62.240 192.630 62.495 192.725 ;
        RECT 61.355 192.460 62.495 192.630 ;
        RECT 62.665 192.515 62.995 192.685 ;
        RECT 61.355 192.235 61.525 192.460 ;
        RECT 60.765 192.065 61.525 192.235 ;
        RECT 62.240 192.325 62.495 192.460 ;
        RECT 60.335 191.070 60.510 191.785 ;
        RECT 60.765 191.585 60.935 192.065 ;
        RECT 61.790 191.975 61.960 192.165 ;
        RECT 62.240 192.155 62.650 192.325 ;
        RECT 60.680 191.255 60.935 191.585 ;
        RECT 61.160 191.255 61.490 191.875 ;
        RECT 61.790 191.805 62.310 191.975 ;
        RECT 61.660 191.255 61.950 191.635 ;
        RECT 62.140 191.085 62.310 191.805 ;
        RECT 58.985 190.345 59.155 190.955 ;
        RECT 59.325 190.565 59.655 191.000 ;
        RECT 60.335 190.515 60.595 191.070 ;
        RECT 61.430 190.915 62.310 191.085 ;
        RECT 62.480 191.130 62.650 192.155 ;
        RECT 62.825 192.265 62.995 192.515 ;
        RECT 63.165 192.435 63.415 192.895 ;
        RECT 63.585 192.265 63.765 192.725 ;
        RECT 62.825 192.095 63.765 192.265 ;
        RECT 62.850 191.615 63.330 191.915 ;
        RECT 62.480 190.960 62.830 191.130 ;
        RECT 63.070 191.025 63.330 191.615 ;
        RECT 63.530 191.025 63.790 191.915 ;
        RECT 64.015 191.755 64.295 192.895 ;
        RECT 64.465 191.745 64.795 192.725 ;
        RECT 64.965 191.755 65.225 192.895 ;
        RECT 65.510 192.265 65.795 192.725 ;
        RECT 65.965 192.435 66.235 192.895 ;
        RECT 65.510 192.045 66.465 192.265 ;
        RECT 64.025 191.315 64.360 191.585 ;
        RECT 64.530 191.145 64.700 191.745 ;
        RECT 64.870 191.335 65.205 191.585 ;
        RECT 65.395 191.315 66.085 191.875 ;
        RECT 66.255 191.145 66.465 192.045 ;
        RECT 60.765 190.345 61.195 190.790 ;
        RECT 61.430 190.515 61.600 190.915 ;
        RECT 61.770 190.345 62.490 190.745 ;
        RECT 62.660 190.515 62.830 190.960 ;
        RECT 63.405 190.345 63.805 190.855 ;
        RECT 64.015 190.345 64.325 191.145 ;
        RECT 64.530 190.515 65.225 191.145 ;
        RECT 65.510 190.975 66.465 191.145 ;
        RECT 66.635 191.875 67.035 192.725 ;
        RECT 67.225 192.265 67.505 192.725 ;
        RECT 68.025 192.435 68.350 192.895 ;
        RECT 67.225 192.045 68.350 192.265 ;
        RECT 66.635 191.315 67.730 191.875 ;
        RECT 67.900 191.585 68.350 192.045 ;
        RECT 68.520 191.755 68.905 192.725 ;
        RECT 65.510 190.515 65.795 190.975 ;
        RECT 65.965 190.345 66.235 190.805 ;
        RECT 66.635 190.515 67.035 191.315 ;
        RECT 67.900 191.255 68.455 191.585 ;
        RECT 67.900 191.145 68.350 191.255 ;
        RECT 67.225 190.975 68.350 191.145 ;
        RECT 68.625 191.085 68.905 191.755 ;
        RECT 67.225 190.515 67.505 190.975 ;
        RECT 68.025 190.345 68.350 190.805 ;
        RECT 68.520 190.515 68.905 191.085 ;
        RECT 69.075 191.330 69.425 192.725 ;
        RECT 69.595 192.095 70.000 192.895 ;
        RECT 70.170 192.555 71.705 192.725 ;
        RECT 70.170 191.925 70.340 192.555 ;
        RECT 69.595 191.755 70.340 191.925 ;
        RECT 69.075 190.515 69.345 191.330 ;
        RECT 69.595 191.255 69.765 191.755 ;
        RECT 70.510 191.585 70.780 192.330 ;
        RECT 69.935 191.255 70.270 191.585 ;
        RECT 70.440 191.255 70.780 191.585 ;
        RECT 70.970 191.585 71.205 192.330 ;
        RECT 71.375 191.925 71.705 192.555 ;
        RECT 71.890 192.095 72.125 192.895 ;
        RECT 72.295 191.925 72.585 192.725 ;
        RECT 71.375 191.755 72.585 191.925 ;
        RECT 72.755 191.805 73.965 192.895 ;
        RECT 74.135 192.385 75.325 192.675 ;
        RECT 70.970 191.255 71.260 191.585 ;
        RECT 71.430 191.255 71.830 191.585 ;
        RECT 72.000 191.085 72.170 191.755 ;
        RECT 72.340 191.255 72.585 191.585 ;
        RECT 72.755 191.095 73.275 191.635 ;
        RECT 73.445 191.265 73.965 191.805 ;
        RECT 74.155 192.045 75.325 192.215 ;
        RECT 75.495 192.095 75.775 192.895 ;
        RECT 74.155 191.755 74.480 192.045 ;
        RECT 75.155 191.925 75.325 192.045 ;
        RECT 74.650 191.585 74.845 191.875 ;
        RECT 75.155 191.755 75.815 191.925 ;
        RECT 75.985 191.755 76.260 192.725 ;
        RECT 76.435 191.755 76.695 192.895 ;
        RECT 75.645 191.585 75.815 191.755 ;
        RECT 74.135 191.255 74.480 191.585 ;
        RECT 74.650 191.255 75.475 191.585 ;
        RECT 75.645 191.255 75.920 191.585 ;
        RECT 69.515 190.345 70.185 191.085 ;
        RECT 70.355 190.915 71.750 191.085 ;
        RECT 70.355 190.570 70.650 190.915 ;
        RECT 70.830 190.345 71.205 190.745 ;
        RECT 71.420 190.570 71.750 190.915 ;
        RECT 72.000 190.515 72.585 191.085 ;
        RECT 72.755 190.345 73.965 191.095 ;
        RECT 75.645 191.085 75.815 191.255 ;
        RECT 74.150 190.915 75.815 191.085 ;
        RECT 76.090 191.020 76.260 191.755 ;
        RECT 76.865 191.745 77.195 192.725 ;
        RECT 77.365 191.755 77.645 192.895 ;
        RECT 76.455 191.335 76.790 191.585 ;
        RECT 76.960 191.145 77.130 191.745 ;
        RECT 77.815 191.730 78.105 192.895 ;
        RECT 79.255 191.835 79.585 192.680 ;
        RECT 79.755 191.885 79.925 192.895 ;
        RECT 80.095 192.165 80.435 192.725 ;
        RECT 80.665 192.395 80.980 192.895 ;
        RECT 81.160 192.425 82.045 192.595 ;
        RECT 79.195 191.755 79.585 191.835 ;
        RECT 80.095 191.790 80.990 192.165 ;
        RECT 79.195 191.705 79.410 191.755 ;
        RECT 77.300 191.315 77.635 191.585 ;
        RECT 74.150 190.565 74.405 190.915 ;
        RECT 74.575 190.345 74.905 190.745 ;
        RECT 75.075 190.565 75.245 190.915 ;
        RECT 75.415 190.345 75.795 190.745 ;
        RECT 75.985 190.675 76.260 191.020 ;
        RECT 76.435 190.515 77.130 191.145 ;
        RECT 77.335 190.345 77.645 191.145 ;
        RECT 79.195 191.125 79.365 191.705 ;
        RECT 80.095 191.585 80.285 191.790 ;
        RECT 81.160 191.585 81.330 192.425 ;
        RECT 82.270 192.395 82.520 192.725 ;
        RECT 79.535 191.255 80.285 191.585 ;
        RECT 80.455 191.255 81.330 191.585 ;
        RECT 79.195 191.085 79.420 191.125 ;
        RECT 80.085 191.085 80.285 191.255 ;
        RECT 77.815 190.345 78.105 191.070 ;
        RECT 79.195 191.000 79.575 191.085 ;
        RECT 79.245 190.565 79.575 191.000 ;
        RECT 79.745 190.345 79.915 190.955 ;
        RECT 80.085 190.560 80.415 191.085 ;
        RECT 80.675 190.345 80.885 190.875 ;
        RECT 81.160 190.795 81.330 191.255 ;
        RECT 81.500 191.295 81.820 192.255 ;
        RECT 81.990 191.505 82.180 192.225 ;
        RECT 82.350 191.325 82.520 192.395 ;
        RECT 82.690 192.095 82.860 192.895 ;
        RECT 83.030 192.450 84.135 192.620 ;
        RECT 83.030 191.835 83.200 192.450 ;
        RECT 84.345 192.300 84.595 192.725 ;
        RECT 84.765 192.435 85.030 192.895 ;
        RECT 83.370 191.915 83.900 192.280 ;
        RECT 84.345 192.170 84.650 192.300 ;
        RECT 82.690 191.745 83.200 191.835 ;
        RECT 82.690 191.575 83.560 191.745 ;
        RECT 82.690 191.505 82.860 191.575 ;
        RECT 82.980 191.325 83.180 191.355 ;
        RECT 81.500 190.965 81.965 191.295 ;
        RECT 82.350 191.025 83.180 191.325 ;
        RECT 82.350 190.795 82.520 191.025 ;
        RECT 81.160 190.625 81.945 190.795 ;
        RECT 82.115 190.625 82.520 190.795 ;
        RECT 82.700 190.345 83.070 190.845 ;
        RECT 83.390 190.795 83.560 191.575 ;
        RECT 83.730 191.215 83.900 191.915 ;
        RECT 84.070 191.385 84.310 191.980 ;
        RECT 83.730 190.995 84.255 191.215 ;
        RECT 84.480 191.065 84.650 192.170 ;
        RECT 84.425 190.935 84.650 191.065 ;
        RECT 84.820 190.975 85.100 191.925 ;
        RECT 84.425 190.795 84.595 190.935 ;
        RECT 83.390 190.625 84.065 190.795 ;
        RECT 84.260 190.625 84.595 190.795 ;
        RECT 84.765 190.345 85.015 190.805 ;
        RECT 85.270 190.605 85.455 192.725 ;
        RECT 85.625 192.395 85.955 192.895 ;
        RECT 86.125 192.225 86.295 192.725 ;
        RECT 85.630 192.055 86.295 192.225 ;
        RECT 86.670 192.265 86.955 192.725 ;
        RECT 87.125 192.435 87.395 192.895 ;
        RECT 85.630 191.065 85.860 192.055 ;
        RECT 86.670 192.045 87.625 192.265 ;
        RECT 86.030 191.235 86.380 191.885 ;
        RECT 86.555 191.315 87.245 191.875 ;
        RECT 87.415 191.145 87.625 192.045 ;
        RECT 85.630 190.895 86.295 191.065 ;
        RECT 85.625 190.345 85.955 190.725 ;
        RECT 86.125 190.605 86.295 190.895 ;
        RECT 86.670 190.975 87.625 191.145 ;
        RECT 87.795 191.875 88.195 192.725 ;
        RECT 88.385 192.265 88.665 192.725 ;
        RECT 89.185 192.435 89.510 192.895 ;
        RECT 88.385 192.045 89.510 192.265 ;
        RECT 87.795 191.315 88.890 191.875 ;
        RECT 89.060 191.585 89.510 192.045 ;
        RECT 89.680 191.755 90.065 192.725 ;
        RECT 90.325 192.225 90.495 192.725 ;
        RECT 90.665 192.395 90.995 192.895 ;
        RECT 90.325 192.055 90.990 192.225 ;
        RECT 86.670 190.515 86.955 190.975 ;
        RECT 87.125 190.345 87.395 190.805 ;
        RECT 87.795 190.515 88.195 191.315 ;
        RECT 89.060 191.255 89.615 191.585 ;
        RECT 89.060 191.145 89.510 191.255 ;
        RECT 88.385 190.975 89.510 191.145 ;
        RECT 89.785 191.085 90.065 191.755 ;
        RECT 90.240 191.235 90.590 191.885 ;
        RECT 88.385 190.515 88.665 190.975 ;
        RECT 89.185 190.345 89.510 190.805 ;
        RECT 89.680 190.515 90.065 191.085 ;
        RECT 90.760 191.065 90.990 192.055 ;
        RECT 90.325 190.895 90.990 191.065 ;
        RECT 90.325 190.605 90.495 190.895 ;
        RECT 90.665 190.345 90.995 190.725 ;
        RECT 91.165 190.605 91.350 192.725 ;
        RECT 91.590 192.435 91.855 192.895 ;
        RECT 92.025 192.300 92.275 192.725 ;
        RECT 92.485 192.450 93.590 192.620 ;
        RECT 91.970 192.170 92.275 192.300 ;
        RECT 91.520 190.975 91.800 191.925 ;
        RECT 91.970 191.065 92.140 192.170 ;
        RECT 92.310 191.385 92.550 191.980 ;
        RECT 92.720 191.915 93.250 192.280 ;
        RECT 92.720 191.215 92.890 191.915 ;
        RECT 93.420 191.835 93.590 192.450 ;
        RECT 93.760 192.095 93.930 192.895 ;
        RECT 94.100 192.395 94.350 192.725 ;
        RECT 94.575 192.425 95.460 192.595 ;
        RECT 93.420 191.745 93.930 191.835 ;
        RECT 91.970 190.935 92.195 191.065 ;
        RECT 92.365 190.995 92.890 191.215 ;
        RECT 93.060 191.575 93.930 191.745 ;
        RECT 91.605 190.345 91.855 190.805 ;
        RECT 92.025 190.795 92.195 190.935 ;
        RECT 93.060 190.795 93.230 191.575 ;
        RECT 93.760 191.505 93.930 191.575 ;
        RECT 93.440 191.325 93.640 191.355 ;
        RECT 94.100 191.325 94.270 192.395 ;
        RECT 94.440 191.505 94.630 192.225 ;
        RECT 93.440 191.025 94.270 191.325 ;
        RECT 94.800 191.295 95.120 192.255 ;
        RECT 92.025 190.625 92.360 190.795 ;
        RECT 92.555 190.625 93.230 190.795 ;
        RECT 93.550 190.345 93.920 190.845 ;
        RECT 94.100 190.795 94.270 191.025 ;
        RECT 94.655 190.965 95.120 191.295 ;
        RECT 95.290 191.585 95.460 192.425 ;
        RECT 95.640 192.395 95.955 192.895 ;
        RECT 96.185 192.165 96.525 192.725 ;
        RECT 95.630 191.790 96.525 192.165 ;
        RECT 96.695 191.885 96.865 192.895 ;
        RECT 96.335 191.585 96.525 191.790 ;
        RECT 97.035 191.835 97.365 192.680 ;
        RECT 97.035 191.755 97.425 191.835 ;
        RECT 97.210 191.705 97.425 191.755 ;
        RECT 95.290 191.255 96.165 191.585 ;
        RECT 96.335 191.255 97.085 191.585 ;
        RECT 95.290 190.795 95.460 191.255 ;
        RECT 96.335 191.085 96.535 191.255 ;
        RECT 97.255 191.125 97.425 191.705 ;
        RECT 97.200 191.085 97.425 191.125 ;
        RECT 94.100 190.625 94.505 190.795 ;
        RECT 94.675 190.625 95.460 190.795 ;
        RECT 95.735 190.345 95.945 190.875 ;
        RECT 96.205 190.560 96.535 191.085 ;
        RECT 97.045 191.000 97.425 191.085 ;
        RECT 97.595 191.755 97.980 192.725 ;
        RECT 98.150 192.435 98.475 192.895 ;
        RECT 98.995 192.265 99.275 192.725 ;
        RECT 98.150 192.045 99.275 192.265 ;
        RECT 97.595 191.085 97.875 191.755 ;
        RECT 98.150 191.585 98.600 192.045 ;
        RECT 99.465 191.875 99.865 192.725 ;
        RECT 100.265 192.435 100.535 192.895 ;
        RECT 100.705 192.265 100.990 192.725 ;
        RECT 101.275 192.385 102.465 192.675 ;
        RECT 98.045 191.255 98.600 191.585 ;
        RECT 98.770 191.315 99.865 191.875 ;
        RECT 98.150 191.145 98.600 191.255 ;
        RECT 96.705 190.345 96.875 190.955 ;
        RECT 97.045 190.565 97.375 191.000 ;
        RECT 97.595 190.515 97.980 191.085 ;
        RECT 98.150 190.975 99.275 191.145 ;
        RECT 98.150 190.345 98.475 190.805 ;
        RECT 98.995 190.515 99.275 190.975 ;
        RECT 99.465 190.515 99.865 191.315 ;
        RECT 100.035 192.045 100.990 192.265 ;
        RECT 101.295 192.045 102.465 192.215 ;
        RECT 102.635 192.095 102.915 192.895 ;
        RECT 100.035 191.145 100.245 192.045 ;
        RECT 100.415 191.315 101.105 191.875 ;
        RECT 101.295 191.755 101.620 192.045 ;
        RECT 102.295 191.925 102.465 192.045 ;
        RECT 101.790 191.585 101.985 191.875 ;
        RECT 102.295 191.755 102.955 191.925 ;
        RECT 103.125 191.755 103.400 192.725 ;
        RECT 102.785 191.585 102.955 191.755 ;
        RECT 101.275 191.255 101.620 191.585 ;
        RECT 101.790 191.255 102.615 191.585 ;
        RECT 102.785 191.255 103.060 191.585 ;
        RECT 100.035 190.975 100.990 191.145 ;
        RECT 102.785 191.085 102.955 191.255 ;
        RECT 100.265 190.345 100.535 190.805 ;
        RECT 100.705 190.515 100.990 190.975 ;
        RECT 101.290 190.915 102.955 191.085 ;
        RECT 103.230 191.020 103.400 191.755 ;
        RECT 103.575 191.730 103.865 192.895 ;
        RECT 104.040 191.945 104.305 192.715 ;
        RECT 104.475 192.175 104.805 192.895 ;
        RECT 104.995 192.355 105.255 192.715 ;
        RECT 105.425 192.525 105.755 192.895 ;
        RECT 105.925 192.355 106.185 192.715 ;
        RECT 104.995 192.125 106.185 192.355 ;
        RECT 106.755 191.945 107.045 192.715 ;
        RECT 101.290 190.565 101.545 190.915 ;
        RECT 101.715 190.345 102.045 190.745 ;
        RECT 102.215 190.565 102.385 190.915 ;
        RECT 102.555 190.345 102.935 190.745 ;
        RECT 103.125 190.675 103.400 191.020 ;
        RECT 103.575 190.345 103.865 191.070 ;
        RECT 104.040 190.525 104.375 191.945 ;
        RECT 104.550 191.765 107.045 191.945 ;
        RECT 104.550 191.075 104.775 191.765 ;
        RECT 107.255 191.755 107.515 192.895 ;
        RECT 107.685 191.925 108.015 192.725 ;
        RECT 108.185 192.095 108.355 192.895 ;
        RECT 108.525 191.925 108.855 192.725 ;
        RECT 109.025 192.095 109.280 192.895 ;
        RECT 110.105 192.555 111.265 192.725 ;
        RECT 110.105 192.055 110.275 192.555 ;
        RECT 110.535 191.925 110.705 192.385 ;
        RECT 110.935 192.305 111.265 192.555 ;
        RECT 111.490 192.475 111.820 192.895 ;
        RECT 112.075 192.305 112.360 192.725 ;
        RECT 110.935 192.135 112.360 192.305 ;
        RECT 112.605 192.095 112.935 192.895 ;
        RECT 113.185 192.175 113.520 192.685 ;
        RECT 107.685 191.755 109.385 191.925 ;
        RECT 104.975 191.255 105.255 191.585 ;
        RECT 105.435 191.255 106.010 191.585 ;
        RECT 106.190 191.255 106.625 191.585 ;
        RECT 106.805 191.255 107.075 191.585 ;
        RECT 107.255 191.335 108.015 191.585 ;
        RECT 108.185 191.335 108.935 191.585 ;
        RECT 109.105 191.165 109.385 191.755 ;
        RECT 110.080 191.585 110.285 191.875 ;
        RECT 110.535 191.755 112.905 191.925 ;
        RECT 112.735 191.585 112.905 191.755 ;
        RECT 110.080 191.535 110.430 191.585 ;
        RECT 110.075 191.365 110.430 191.535 ;
        RECT 110.080 191.255 110.430 191.365 ;
        RECT 104.550 190.885 107.035 191.075 ;
        RECT 104.555 190.345 105.300 190.715 ;
        RECT 105.865 190.525 106.120 190.885 ;
        RECT 106.300 190.345 106.630 190.715 ;
        RECT 106.810 190.525 107.035 190.885 ;
        RECT 107.255 190.975 108.355 191.145 ;
        RECT 107.255 190.515 107.595 190.975 ;
        RECT 107.765 190.345 107.935 190.805 ;
        RECT 108.105 190.725 108.355 190.975 ;
        RECT 108.525 190.915 109.385 191.165 ;
        RECT 108.945 190.725 109.275 190.745 ;
        RECT 108.105 190.515 109.275 190.725 ;
        RECT 110.025 190.345 110.355 191.065 ;
        RECT 110.740 190.920 111.160 191.585 ;
        RECT 111.330 191.195 111.620 191.585 ;
        RECT 111.810 191.195 112.080 191.585 ;
        RECT 112.290 191.535 112.540 191.585 ;
        RECT 112.290 191.365 112.545 191.535 ;
        RECT 112.290 191.255 112.540 191.365 ;
        RECT 112.735 191.255 113.040 191.585 ;
        RECT 111.330 191.025 111.625 191.195 ;
        RECT 111.810 191.025 112.085 191.195 ;
        RECT 112.735 191.085 112.905 191.255 ;
        RECT 111.330 190.925 111.620 191.025 ;
        RECT 111.810 190.925 112.080 191.025 ;
        RECT 112.345 190.915 112.905 191.085 ;
        RECT 112.345 190.745 112.515 190.915 ;
        RECT 113.265 190.820 113.520 192.175 ;
        RECT 110.900 190.575 112.515 190.745 ;
        RECT 112.685 190.345 113.015 190.745 ;
        RECT 113.185 190.560 113.520 190.820 ;
        RECT 113.730 192.105 114.265 192.725 ;
        RECT 113.730 191.085 114.045 192.105 ;
        RECT 114.435 192.095 114.765 192.895 ;
        RECT 115.250 191.925 115.640 192.100 ;
        RECT 114.215 191.755 115.640 191.925 ;
        RECT 116.005 191.925 116.335 192.710 ;
        RECT 116.005 191.755 116.685 191.925 ;
        RECT 116.865 191.755 117.195 192.895 ;
        RECT 117.375 191.755 117.635 192.895 ;
        RECT 114.215 191.255 114.385 191.755 ;
        RECT 113.730 190.515 114.345 191.085 ;
        RECT 114.635 191.025 114.900 191.585 ;
        RECT 115.070 190.855 115.240 191.755 ;
        RECT 115.410 191.025 115.765 191.585 ;
        RECT 115.995 191.335 116.345 191.585 ;
        RECT 116.515 191.155 116.685 191.755 ;
        RECT 117.805 191.745 118.135 192.725 ;
        RECT 118.305 191.755 118.585 192.895 ;
        RECT 118.755 192.460 124.100 192.895 ;
        RECT 116.855 191.335 117.205 191.585 ;
        RECT 117.395 191.335 117.730 191.585 ;
        RECT 114.515 190.345 114.730 190.855 ;
        RECT 114.960 190.525 115.240 190.855 ;
        RECT 115.420 190.345 115.660 190.855 ;
        RECT 116.015 190.345 116.255 191.155 ;
        RECT 116.425 190.515 116.755 191.155 ;
        RECT 116.925 190.345 117.195 191.155 ;
        RECT 117.900 191.145 118.070 191.745 ;
        RECT 118.240 191.315 118.575 191.585 ;
        RECT 117.375 190.515 118.070 191.145 ;
        RECT 118.275 190.345 118.585 191.145 ;
        RECT 120.340 190.890 120.680 191.720 ;
        RECT 122.160 191.210 122.510 192.460 ;
        RECT 124.275 191.805 127.785 192.895 ;
        RECT 127.955 191.805 129.165 192.895 ;
        RECT 124.275 191.115 125.925 191.635 ;
        RECT 126.095 191.285 127.785 191.805 ;
        RECT 118.755 190.345 124.100 190.890 ;
        RECT 124.275 190.345 127.785 191.115 ;
        RECT 127.955 191.095 128.475 191.635 ;
        RECT 128.645 191.265 129.165 191.805 ;
        RECT 129.335 191.730 129.625 192.895 ;
        RECT 129.795 191.805 133.305 192.895 ;
        RECT 129.795 191.115 131.445 191.635 ;
        RECT 131.615 191.285 133.305 191.805 ;
        RECT 134.025 191.965 134.195 192.725 ;
        RECT 134.375 192.135 134.705 192.895 ;
        RECT 134.025 191.795 134.690 191.965 ;
        RECT 134.875 191.820 135.145 192.725 ;
        RECT 134.520 191.650 134.690 191.795 ;
        RECT 133.955 191.245 134.285 191.615 ;
        RECT 134.520 191.320 134.805 191.650 ;
        RECT 127.955 190.345 129.165 191.095 ;
        RECT 129.335 190.345 129.625 191.070 ;
        RECT 129.795 190.345 133.305 191.115 ;
        RECT 134.520 191.065 134.690 191.320 ;
        RECT 134.025 190.895 134.690 191.065 ;
        RECT 134.975 191.020 135.145 191.820 ;
        RECT 134.025 190.515 134.195 190.895 ;
        RECT 134.375 190.345 134.705 190.725 ;
        RECT 134.885 190.515 135.145 191.020 ;
        RECT 136.235 191.820 136.505 192.725 ;
        RECT 136.675 192.135 137.005 192.895 ;
        RECT 137.185 191.965 137.365 192.725 ;
        RECT 136.235 191.020 136.415 191.820 ;
        RECT 136.690 191.795 137.365 191.965 ;
        RECT 137.615 191.805 138.825 192.895 ;
        RECT 136.690 191.650 136.860 191.795 ;
        RECT 136.585 191.320 136.860 191.650 ;
        RECT 136.690 191.065 136.860 191.320 ;
        RECT 137.085 191.245 137.425 191.615 ;
        RECT 137.615 191.265 138.135 191.805 ;
        RECT 138.305 191.095 138.825 191.635 ;
        RECT 136.235 190.515 136.495 191.020 ;
        RECT 136.690 190.895 137.355 191.065 ;
        RECT 136.675 190.345 137.005 190.725 ;
        RECT 137.185 190.515 137.355 190.895 ;
        RECT 137.615 190.345 138.825 191.095 ;
        RECT 13.330 190.175 138.910 190.345 ;
        RECT 13.415 189.425 14.625 190.175 ;
        RECT 14.795 189.630 20.140 190.175 ;
        RECT 20.320 189.920 20.655 189.965 ;
        RECT 13.415 188.885 13.935 189.425 ;
        RECT 14.105 188.715 14.625 189.255 ;
        RECT 16.380 188.800 16.720 189.630 ;
        RECT 20.315 189.455 20.655 189.920 ;
        RECT 20.825 189.795 21.155 190.175 ;
        RECT 13.415 187.625 14.625 188.715 ;
        RECT 18.200 188.060 18.550 189.310 ;
        RECT 20.315 188.765 20.485 189.455 ;
        RECT 20.655 188.935 20.915 189.265 ;
        RECT 14.795 187.625 20.140 188.060 ;
        RECT 20.315 187.795 20.575 188.765 ;
        RECT 20.745 188.385 20.915 188.935 ;
        RECT 21.085 188.565 21.425 189.595 ;
        RECT 21.615 188.815 21.885 189.840 ;
        RECT 21.615 188.645 21.925 188.815 ;
        RECT 21.615 188.565 21.885 188.645 ;
        RECT 22.110 188.565 22.390 189.840 ;
        RECT 22.590 189.675 22.820 190.005 ;
        RECT 23.065 189.795 23.395 190.175 ;
        RECT 22.590 188.385 22.760 189.675 ;
        RECT 23.565 189.605 23.740 190.005 ;
        RECT 23.110 189.435 23.740 189.605 ;
        RECT 23.110 189.265 23.280 189.435 ;
        RECT 23.995 189.340 24.285 190.175 ;
        RECT 24.455 189.775 25.410 189.945 ;
        RECT 25.825 189.785 26.155 190.175 ;
        RECT 22.930 188.935 23.280 189.265 ;
        RECT 20.745 188.215 22.760 188.385 ;
        RECT 23.110 188.415 23.280 188.935 ;
        RECT 23.460 188.585 23.825 189.265 ;
        RECT 24.455 188.895 24.625 189.775 ;
        RECT 26.325 189.605 26.495 189.925 ;
        RECT 26.665 189.785 26.995 190.175 ;
        RECT 24.795 189.435 27.045 189.605 ;
        RECT 24.795 188.935 25.025 189.435 ;
        RECT 25.195 189.015 25.570 189.185 ;
        RECT 23.995 188.725 24.625 188.895 ;
        RECT 25.400 188.815 25.570 189.015 ;
        RECT 25.740 188.985 26.290 189.185 ;
        RECT 26.460 188.815 26.705 189.265 ;
        RECT 23.110 188.245 23.740 188.415 ;
        RECT 20.770 187.625 21.100 188.035 ;
        RECT 21.300 187.795 21.470 188.215 ;
        RECT 21.685 187.625 22.355 188.035 ;
        RECT 22.590 187.795 22.760 188.215 ;
        RECT 23.065 187.625 23.395 188.065 ;
        RECT 23.565 187.795 23.740 188.245 ;
        RECT 23.995 187.795 24.315 188.725 ;
        RECT 25.400 188.645 26.705 188.815 ;
        RECT 26.875 188.475 27.045 189.435 ;
        RECT 27.215 189.425 28.425 190.175 ;
        RECT 28.595 189.795 29.485 189.965 ;
        RECT 27.215 188.885 27.735 189.425 ;
        RECT 27.905 188.715 28.425 189.255 ;
        RECT 28.595 189.240 29.145 189.625 ;
        RECT 29.315 189.070 29.485 189.795 ;
        RECT 24.495 188.305 25.735 188.475 ;
        RECT 24.495 187.795 24.895 188.305 ;
        RECT 25.065 187.625 25.235 188.135 ;
        RECT 25.405 187.795 25.735 188.305 ;
        RECT 25.905 187.625 26.075 188.475 ;
        RECT 26.665 187.795 27.045 188.475 ;
        RECT 27.215 187.625 28.425 188.715 ;
        RECT 28.595 189.000 29.485 189.070 ;
        RECT 29.655 189.470 29.875 189.955 ;
        RECT 30.045 189.635 30.295 190.175 ;
        RECT 30.465 189.525 30.725 190.005 ;
        RECT 29.655 189.045 29.985 189.470 ;
        RECT 28.595 188.975 29.490 189.000 ;
        RECT 28.595 188.960 29.500 188.975 ;
        RECT 28.595 188.945 29.505 188.960 ;
        RECT 28.595 188.940 29.515 188.945 ;
        RECT 28.595 188.930 29.520 188.940 ;
        RECT 28.595 188.920 29.525 188.930 ;
        RECT 28.595 188.915 29.535 188.920 ;
        RECT 28.595 188.905 29.545 188.915 ;
        RECT 28.595 188.900 29.555 188.905 ;
        RECT 28.595 188.450 28.855 188.900 ;
        RECT 29.220 188.895 29.555 188.900 ;
        RECT 29.220 188.890 29.570 188.895 ;
        RECT 29.220 188.880 29.585 188.890 ;
        RECT 29.220 188.875 29.610 188.880 ;
        RECT 30.155 188.875 30.385 189.270 ;
        RECT 29.220 188.870 30.385 188.875 ;
        RECT 29.250 188.835 30.385 188.870 ;
        RECT 29.285 188.810 30.385 188.835 ;
        RECT 29.315 188.780 30.385 188.810 ;
        RECT 29.335 188.750 30.385 188.780 ;
        RECT 29.355 188.720 30.385 188.750 ;
        RECT 29.425 188.710 30.385 188.720 ;
        RECT 29.450 188.700 30.385 188.710 ;
        RECT 29.470 188.685 30.385 188.700 ;
        RECT 29.490 188.670 30.385 188.685 ;
        RECT 29.495 188.660 30.280 188.670 ;
        RECT 29.510 188.625 30.280 188.660 ;
        RECT 29.025 188.305 29.355 188.550 ;
        RECT 29.525 188.375 30.280 188.625 ;
        RECT 30.555 188.495 30.725 189.525 ;
        RECT 30.985 189.625 31.155 189.915 ;
        RECT 31.325 189.795 31.655 190.175 ;
        RECT 30.985 189.455 31.650 189.625 ;
        RECT 30.900 188.635 31.250 189.285 ;
        RECT 29.025 188.280 29.210 188.305 ;
        RECT 28.595 188.180 29.210 188.280 ;
        RECT 28.595 187.625 29.200 188.180 ;
        RECT 29.375 187.795 29.855 188.135 ;
        RECT 30.025 187.625 30.280 188.170 ;
        RECT 30.450 187.795 30.725 188.495 ;
        RECT 31.420 188.465 31.650 189.455 ;
        RECT 30.985 188.295 31.650 188.465 ;
        RECT 30.985 187.795 31.155 188.295 ;
        RECT 31.325 187.625 31.655 188.125 ;
        RECT 31.825 187.795 32.010 189.915 ;
        RECT 32.265 189.715 32.515 190.175 ;
        RECT 32.685 189.725 33.020 189.895 ;
        RECT 33.215 189.725 33.890 189.895 ;
        RECT 32.685 189.585 32.855 189.725 ;
        RECT 32.180 188.595 32.460 189.545 ;
        RECT 32.630 189.455 32.855 189.585 ;
        RECT 32.630 188.350 32.800 189.455 ;
        RECT 33.025 189.305 33.550 189.525 ;
        RECT 32.970 188.540 33.210 189.135 ;
        RECT 33.380 188.605 33.550 189.305 ;
        RECT 33.720 188.945 33.890 189.725 ;
        RECT 34.210 189.675 34.580 190.175 ;
        RECT 34.760 189.725 35.165 189.895 ;
        RECT 35.335 189.725 36.120 189.895 ;
        RECT 34.760 189.495 34.930 189.725 ;
        RECT 34.100 189.195 34.930 189.495 ;
        RECT 35.315 189.225 35.780 189.555 ;
        RECT 34.100 189.165 34.300 189.195 ;
        RECT 34.420 188.945 34.590 189.015 ;
        RECT 33.720 188.775 34.590 188.945 ;
        RECT 34.080 188.685 34.590 188.775 ;
        RECT 32.630 188.220 32.935 188.350 ;
        RECT 33.380 188.240 33.910 188.605 ;
        RECT 32.250 187.625 32.515 188.085 ;
        RECT 32.685 187.795 32.935 188.220 ;
        RECT 34.080 188.070 34.250 188.685 ;
        RECT 33.145 187.900 34.250 188.070 ;
        RECT 34.420 187.625 34.590 188.425 ;
        RECT 34.760 188.125 34.930 189.195 ;
        RECT 35.100 188.295 35.290 189.015 ;
        RECT 35.460 188.265 35.780 189.225 ;
        RECT 35.950 189.265 36.120 189.725 ;
        RECT 36.395 189.645 36.605 190.175 ;
        RECT 36.865 189.435 37.195 189.960 ;
        RECT 37.365 189.565 37.535 190.175 ;
        RECT 37.705 189.520 38.035 189.955 ;
        RECT 37.705 189.435 38.085 189.520 ;
        RECT 39.175 189.450 39.465 190.175 ;
        RECT 39.685 189.785 40.015 190.175 ;
        RECT 40.185 189.605 40.355 189.925 ;
        RECT 40.525 189.785 40.855 190.175 ;
        RECT 41.270 189.775 42.225 189.945 ;
        RECT 36.995 189.265 37.195 189.435 ;
        RECT 37.860 189.395 38.085 189.435 ;
        RECT 35.950 188.935 36.825 189.265 ;
        RECT 36.995 188.935 37.745 189.265 ;
        RECT 34.760 187.795 35.010 188.125 ;
        RECT 35.950 188.095 36.120 188.935 ;
        RECT 36.995 188.730 37.185 188.935 ;
        RECT 37.915 188.815 38.085 189.395 ;
        RECT 37.870 188.765 38.085 188.815 ;
        RECT 39.635 189.435 41.885 189.605 ;
        RECT 36.290 188.355 37.185 188.730 ;
        RECT 37.695 188.685 38.085 188.765 ;
        RECT 35.235 187.925 36.120 188.095 ;
        RECT 36.300 187.625 36.615 188.125 ;
        RECT 36.845 187.795 37.185 188.355 ;
        RECT 37.355 187.625 37.525 188.635 ;
        RECT 37.695 187.840 38.025 188.685 ;
        RECT 39.175 187.625 39.465 188.790 ;
        RECT 39.635 188.475 39.805 189.435 ;
        RECT 39.975 188.815 40.220 189.265 ;
        RECT 40.390 188.985 40.940 189.185 ;
        RECT 41.110 189.015 41.485 189.185 ;
        RECT 41.110 188.815 41.280 189.015 ;
        RECT 41.655 188.935 41.885 189.435 ;
        RECT 39.975 188.645 41.280 188.815 ;
        RECT 42.055 188.895 42.225 189.775 ;
        RECT 42.395 189.340 42.685 190.175 ;
        RECT 42.860 189.920 43.195 189.965 ;
        RECT 42.855 189.455 43.195 189.920 ;
        RECT 43.365 189.795 43.695 190.175 ;
        RECT 42.055 188.725 42.685 188.895 ;
        RECT 39.635 187.795 40.015 188.475 ;
        RECT 40.605 187.625 40.775 188.475 ;
        RECT 40.945 188.305 42.185 188.475 ;
        RECT 40.945 187.795 41.275 188.305 ;
        RECT 41.445 187.625 41.615 188.135 ;
        RECT 41.785 187.795 42.185 188.305 ;
        RECT 42.365 187.795 42.685 188.725 ;
        RECT 42.855 188.765 43.025 189.455 ;
        RECT 43.195 188.935 43.455 189.265 ;
        RECT 42.855 187.795 43.115 188.765 ;
        RECT 43.285 188.385 43.455 188.935 ;
        RECT 43.625 188.565 43.965 189.595 ;
        RECT 44.155 189.495 44.425 189.840 ;
        RECT 44.155 189.325 44.465 189.495 ;
        RECT 44.155 188.565 44.425 189.325 ;
        RECT 44.650 188.565 44.930 189.840 ;
        RECT 45.130 189.675 45.360 190.005 ;
        RECT 45.605 189.795 45.935 190.175 ;
        RECT 45.130 188.385 45.300 189.675 ;
        RECT 46.105 189.605 46.280 190.005 ;
        RECT 45.650 189.435 46.280 189.605 ;
        RECT 45.650 189.265 45.820 189.435 ;
        RECT 46.535 189.405 50.045 190.175 ;
        RECT 50.225 189.445 50.525 190.175 ;
        RECT 45.470 188.935 45.820 189.265 ;
        RECT 43.285 188.215 45.300 188.385 ;
        RECT 45.650 188.415 45.820 188.935 ;
        RECT 46.000 188.585 46.365 189.265 ;
        RECT 46.535 188.885 48.185 189.405 ;
        RECT 50.705 189.265 50.935 189.885 ;
        RECT 51.135 189.615 51.360 189.995 ;
        RECT 51.530 189.785 51.860 190.175 ;
        RECT 52.055 189.630 57.400 190.175 ;
        RECT 57.575 189.630 62.920 190.175 ;
        RECT 51.135 189.435 51.465 189.615 ;
        RECT 48.355 188.715 50.045 189.235 ;
        RECT 50.230 188.935 50.525 189.265 ;
        RECT 50.705 188.935 51.120 189.265 ;
        RECT 51.290 188.765 51.465 189.435 ;
        RECT 51.635 188.935 51.875 189.585 ;
        RECT 53.640 188.800 53.980 189.630 ;
        RECT 45.650 188.245 46.280 188.415 ;
        RECT 43.310 187.625 43.640 188.035 ;
        RECT 43.840 187.795 44.010 188.215 ;
        RECT 44.225 187.625 44.895 188.035 ;
        RECT 45.130 187.795 45.300 188.215 ;
        RECT 45.605 187.625 45.935 188.065 ;
        RECT 46.105 187.795 46.280 188.245 ;
        RECT 46.535 187.625 50.045 188.715 ;
        RECT 50.225 188.405 51.120 188.735 ;
        RECT 51.290 188.575 51.875 188.765 ;
        RECT 50.225 188.235 51.430 188.405 ;
        RECT 50.225 187.805 50.555 188.235 ;
        RECT 50.735 187.625 50.930 188.065 ;
        RECT 51.100 187.805 51.430 188.235 ;
        RECT 51.600 187.805 51.875 188.575 ;
        RECT 55.460 188.060 55.810 189.310 ;
        RECT 59.160 188.800 59.500 189.630 ;
        RECT 63.615 189.355 63.825 190.175 ;
        RECT 63.995 189.375 64.325 190.005 ;
        RECT 60.980 188.060 61.330 189.310 ;
        RECT 63.995 188.775 64.245 189.375 ;
        RECT 64.495 189.355 64.725 190.175 ;
        RECT 64.935 189.450 65.225 190.175 ;
        RECT 65.400 189.500 65.675 189.845 ;
        RECT 65.865 189.775 66.245 190.175 ;
        RECT 66.415 189.605 66.585 189.955 ;
        RECT 66.755 189.775 67.085 190.175 ;
        RECT 67.255 189.605 67.510 189.955 ;
        RECT 67.860 189.665 68.100 190.175 ;
        RECT 68.280 189.665 68.560 189.995 ;
        RECT 68.790 189.665 69.005 190.175 ;
        RECT 64.415 188.935 64.745 189.185 ;
        RECT 52.055 187.625 57.400 188.060 ;
        RECT 57.575 187.625 62.920 188.060 ;
        RECT 63.615 187.625 63.825 188.765 ;
        RECT 63.995 187.795 64.325 188.775 ;
        RECT 64.495 187.625 64.725 188.765 ;
        RECT 64.935 187.625 65.225 188.790 ;
        RECT 65.400 188.765 65.570 189.500 ;
        RECT 65.845 189.435 67.510 189.605 ;
        RECT 65.845 189.265 66.015 189.435 ;
        RECT 65.740 188.935 66.015 189.265 ;
        RECT 66.185 188.935 67.010 189.265 ;
        RECT 67.180 188.935 67.525 189.265 ;
        RECT 67.755 188.935 68.110 189.495 ;
        RECT 65.845 188.765 66.015 188.935 ;
        RECT 65.400 187.795 65.675 188.765 ;
        RECT 65.845 188.595 66.505 188.765 ;
        RECT 66.815 188.645 67.010 188.935 ;
        RECT 68.280 188.765 68.450 189.665 ;
        RECT 68.620 188.935 68.885 189.495 ;
        RECT 69.175 189.435 69.790 190.005 ;
        RECT 69.995 189.630 75.340 190.175 ;
        RECT 69.135 188.765 69.305 189.265 ;
        RECT 66.335 188.475 66.505 188.595 ;
        RECT 67.180 188.475 67.505 188.765 ;
        RECT 65.885 187.625 66.165 188.425 ;
        RECT 66.335 188.305 67.505 188.475 ;
        RECT 67.880 188.595 69.305 188.765 ;
        RECT 67.880 188.420 68.270 188.595 ;
        RECT 66.335 187.845 67.525 188.135 ;
        RECT 68.755 187.625 69.085 188.425 ;
        RECT 69.475 188.415 69.790 189.435 ;
        RECT 71.580 188.800 71.920 189.630 ;
        RECT 75.605 189.625 75.775 189.915 ;
        RECT 75.945 189.795 76.275 190.175 ;
        RECT 75.605 189.455 76.270 189.625 ;
        RECT 69.255 187.795 69.790 188.415 ;
        RECT 73.400 188.060 73.750 189.310 ;
        RECT 75.520 188.635 75.870 189.285 ;
        RECT 76.040 188.465 76.270 189.455 ;
        RECT 75.605 188.295 76.270 188.465 ;
        RECT 69.995 187.625 75.340 188.060 ;
        RECT 75.605 187.795 75.775 188.295 ;
        RECT 75.945 187.625 76.275 188.125 ;
        RECT 76.445 187.795 76.630 189.915 ;
        RECT 76.885 189.715 77.135 190.175 ;
        RECT 77.305 189.725 77.640 189.895 ;
        RECT 77.835 189.725 78.510 189.895 ;
        RECT 77.305 189.585 77.475 189.725 ;
        RECT 76.800 188.595 77.080 189.545 ;
        RECT 77.250 189.455 77.475 189.585 ;
        RECT 77.250 188.350 77.420 189.455 ;
        RECT 77.645 189.305 78.170 189.525 ;
        RECT 77.590 188.540 77.830 189.135 ;
        RECT 78.000 188.605 78.170 189.305 ;
        RECT 78.340 188.945 78.510 189.725 ;
        RECT 78.830 189.675 79.200 190.175 ;
        RECT 79.380 189.725 79.785 189.895 ;
        RECT 79.955 189.725 80.740 189.895 ;
        RECT 79.380 189.495 79.550 189.725 ;
        RECT 78.720 189.195 79.550 189.495 ;
        RECT 79.935 189.225 80.400 189.555 ;
        RECT 78.720 189.165 78.920 189.195 ;
        RECT 79.040 188.945 79.210 189.015 ;
        RECT 78.340 188.775 79.210 188.945 ;
        RECT 78.700 188.685 79.210 188.775 ;
        RECT 77.250 188.220 77.555 188.350 ;
        RECT 78.000 188.240 78.530 188.605 ;
        RECT 76.870 187.625 77.135 188.085 ;
        RECT 77.305 187.795 77.555 188.220 ;
        RECT 78.700 188.070 78.870 188.685 ;
        RECT 77.765 187.900 78.870 188.070 ;
        RECT 79.040 187.625 79.210 188.425 ;
        RECT 79.380 188.125 79.550 189.195 ;
        RECT 79.720 188.295 79.910 189.015 ;
        RECT 80.080 188.265 80.400 189.225 ;
        RECT 80.570 189.265 80.740 189.725 ;
        RECT 81.015 189.645 81.225 190.175 ;
        RECT 81.485 189.435 81.815 189.960 ;
        RECT 81.985 189.565 82.155 190.175 ;
        RECT 82.325 189.520 82.655 189.955 ;
        RECT 82.325 189.435 82.705 189.520 ;
        RECT 81.615 189.265 81.815 189.435 ;
        RECT 82.480 189.395 82.705 189.435 ;
        RECT 80.570 188.935 81.445 189.265 ;
        RECT 81.615 188.935 82.365 189.265 ;
        RECT 79.380 187.795 79.630 188.125 ;
        RECT 80.570 188.095 80.740 188.935 ;
        RECT 81.615 188.730 81.805 188.935 ;
        RECT 82.535 188.815 82.705 189.395 ;
        RECT 82.875 189.405 86.385 190.175 ;
        RECT 82.875 188.885 84.525 189.405 ;
        RECT 86.555 189.375 86.895 190.005 ;
        RECT 87.065 189.375 87.315 190.175 ;
        RECT 87.505 189.525 87.835 190.005 ;
        RECT 88.005 189.715 88.230 190.175 ;
        RECT 88.400 189.525 88.730 190.005 ;
        RECT 82.490 188.765 82.705 188.815 ;
        RECT 80.910 188.355 81.805 188.730 ;
        RECT 82.315 188.685 82.705 188.765 ;
        RECT 84.695 188.715 86.385 189.235 ;
        RECT 79.855 187.925 80.740 188.095 ;
        RECT 80.920 187.625 81.235 188.125 ;
        RECT 81.465 187.795 81.805 188.355 ;
        RECT 81.975 187.625 82.145 188.635 ;
        RECT 82.315 187.840 82.645 188.685 ;
        RECT 82.875 187.625 86.385 188.715 ;
        RECT 86.555 188.765 86.730 189.375 ;
        RECT 87.505 189.355 88.730 189.525 ;
        RECT 89.360 189.395 89.860 190.005 ;
        RECT 90.695 189.450 90.985 190.175 ;
        RECT 91.700 189.605 91.875 190.005 ;
        RECT 92.045 189.795 92.375 190.175 ;
        RECT 92.620 189.675 92.850 190.005 ;
        RECT 91.700 189.435 92.330 189.605 ;
        RECT 86.900 189.015 87.595 189.185 ;
        RECT 87.425 188.765 87.595 189.015 ;
        RECT 87.770 188.985 88.190 189.185 ;
        RECT 88.360 188.985 88.690 189.185 ;
        RECT 88.860 188.985 89.190 189.185 ;
        RECT 89.360 188.765 89.530 189.395 ;
        RECT 92.160 189.265 92.330 189.435 ;
        RECT 89.715 188.935 90.065 189.185 ;
        RECT 86.555 187.795 86.895 188.765 ;
        RECT 87.065 187.625 87.235 188.765 ;
        RECT 87.425 188.595 89.860 188.765 ;
        RECT 87.505 187.625 87.755 188.425 ;
        RECT 88.400 187.795 88.730 188.595 ;
        RECT 89.030 187.625 89.360 188.425 ;
        RECT 89.530 187.795 89.860 188.595 ;
        RECT 90.695 187.625 90.985 188.790 ;
        RECT 91.615 188.585 91.980 189.265 ;
        RECT 92.160 188.935 92.510 189.265 ;
        RECT 92.160 188.415 92.330 188.935 ;
        RECT 91.700 188.245 92.330 188.415 ;
        RECT 92.680 188.385 92.850 189.675 ;
        RECT 93.050 188.565 93.330 189.840 ;
        RECT 93.555 189.495 93.825 189.840 ;
        RECT 94.285 189.795 94.615 190.175 ;
        RECT 94.785 189.920 95.120 189.965 ;
        RECT 93.515 189.325 93.825 189.495 ;
        RECT 93.555 188.565 93.825 189.325 ;
        RECT 94.015 188.565 94.355 189.595 ;
        RECT 94.785 189.455 95.125 189.920 ;
        RECT 94.525 188.935 94.785 189.265 ;
        RECT 94.525 188.385 94.695 188.935 ;
        RECT 94.955 188.765 95.125 189.455 ;
        RECT 95.295 189.355 95.555 190.175 ;
        RECT 95.725 189.355 96.055 189.775 ;
        RECT 96.235 189.690 97.025 189.955 ;
        RECT 95.805 189.265 96.055 189.355 ;
        RECT 91.700 187.795 91.875 188.245 ;
        RECT 92.680 188.215 94.695 188.385 ;
        RECT 92.045 187.625 92.375 188.065 ;
        RECT 92.680 187.795 92.850 188.215 ;
        RECT 93.085 187.625 93.755 188.035 ;
        RECT 93.970 187.795 94.140 188.215 ;
        RECT 94.340 187.625 94.670 188.035 ;
        RECT 94.865 187.795 95.125 188.765 ;
        RECT 95.295 188.305 95.635 189.185 ;
        RECT 95.805 189.015 96.600 189.265 ;
        RECT 95.295 187.625 95.555 188.135 ;
        RECT 95.805 187.795 95.975 189.015 ;
        RECT 96.770 188.835 97.025 189.690 ;
        RECT 97.195 189.535 97.395 189.955 ;
        RECT 97.585 189.715 97.915 190.175 ;
        RECT 97.195 189.015 97.605 189.535 ;
        RECT 98.085 189.525 98.345 190.005 ;
        RECT 97.775 188.835 98.005 189.265 ;
        RECT 96.215 188.665 98.005 188.835 ;
        RECT 96.215 188.300 96.465 188.665 ;
        RECT 96.635 188.305 96.965 188.495 ;
        RECT 97.185 188.370 97.900 188.665 ;
        RECT 98.175 188.495 98.345 189.525 ;
        RECT 96.635 188.130 96.830 188.305 ;
        RECT 96.215 187.625 96.830 188.130 ;
        RECT 97.000 187.795 97.475 188.135 ;
        RECT 97.645 187.625 97.860 188.170 ;
        RECT 98.070 187.795 98.345 188.495 ;
        RECT 98.515 189.675 98.775 190.005 ;
        RECT 98.945 189.815 99.275 190.175 ;
        RECT 99.530 189.795 100.830 190.005 ;
        RECT 98.515 189.665 98.745 189.675 ;
        RECT 98.515 188.475 98.685 189.665 ;
        RECT 99.530 189.645 99.700 189.795 ;
        RECT 98.945 189.520 99.700 189.645 ;
        RECT 98.855 189.475 99.700 189.520 ;
        RECT 98.855 189.355 99.125 189.475 ;
        RECT 98.855 188.780 99.025 189.355 ;
        RECT 99.255 188.915 99.665 189.220 ;
        RECT 99.955 189.185 100.165 189.585 ;
        RECT 99.835 188.975 100.165 189.185 ;
        RECT 100.410 189.185 100.630 189.585 ;
        RECT 101.105 189.410 101.560 190.175 ;
        RECT 101.735 189.230 102.075 190.005 ;
        RECT 102.245 189.715 102.415 190.175 ;
        RECT 102.655 189.740 103.015 190.005 ;
        RECT 102.655 189.735 103.010 189.740 ;
        RECT 102.655 189.725 103.005 189.735 ;
        RECT 102.655 189.720 103.000 189.725 ;
        RECT 102.655 189.710 102.995 189.720 ;
        RECT 103.645 189.715 103.815 190.175 ;
        RECT 102.655 189.705 102.990 189.710 ;
        RECT 102.655 189.695 102.980 189.705 ;
        RECT 102.655 189.685 102.970 189.695 ;
        RECT 102.655 189.545 102.955 189.685 ;
        RECT 102.245 189.355 102.955 189.545 ;
        RECT 103.145 189.545 103.475 189.625 ;
        RECT 103.985 189.545 104.325 190.005 ;
        RECT 103.145 189.355 104.325 189.545 ;
        RECT 104.495 189.545 104.835 190.005 ;
        RECT 105.005 189.715 105.175 190.175 ;
        RECT 105.345 189.795 106.515 190.005 ;
        RECT 105.345 189.545 105.595 189.795 ;
        RECT 106.185 189.775 106.515 189.795 ;
        RECT 104.495 189.375 105.595 189.545 ;
        RECT 105.765 189.355 106.625 189.605 ;
        RECT 100.410 188.975 100.885 189.185 ;
        RECT 101.075 188.985 101.565 189.185 ;
        RECT 98.855 188.745 99.055 188.780 ;
        RECT 100.385 188.745 101.560 188.805 ;
        RECT 98.855 188.635 101.560 188.745 ;
        RECT 98.915 188.575 100.715 188.635 ;
        RECT 100.385 188.545 100.715 188.575 ;
        RECT 98.515 187.795 98.775 188.475 ;
        RECT 98.945 187.625 99.195 188.405 ;
        RECT 99.445 188.375 100.280 188.385 ;
        RECT 100.870 188.375 101.055 188.465 ;
        RECT 99.445 188.175 101.055 188.375 ;
        RECT 99.445 187.795 99.695 188.175 ;
        RECT 100.825 188.135 101.055 188.175 ;
        RECT 101.305 188.015 101.560 188.635 ;
        RECT 99.865 187.625 100.220 188.005 ;
        RECT 101.225 187.795 101.560 188.015 ;
        RECT 101.735 187.795 102.015 189.230 ;
        RECT 102.245 188.785 102.530 189.355 ;
        RECT 102.715 188.955 103.185 189.185 ;
        RECT 103.355 189.165 103.685 189.185 ;
        RECT 103.355 188.985 103.805 189.165 ;
        RECT 103.995 188.985 104.325 189.185 ;
        RECT 102.245 188.570 103.395 188.785 ;
        RECT 102.185 187.625 102.895 188.400 ;
        RECT 103.065 187.795 103.395 188.570 ;
        RECT 103.590 187.870 103.805 188.985 ;
        RECT 104.095 188.645 104.325 188.985 ;
        RECT 104.495 188.935 105.255 189.185 ;
        RECT 105.425 188.935 106.175 189.185 ;
        RECT 106.345 188.765 106.625 189.355 ;
        RECT 103.985 187.625 104.315 188.345 ;
        RECT 104.495 187.625 104.755 188.765 ;
        RECT 104.925 188.595 106.625 188.765 ;
        RECT 106.795 189.525 107.055 190.005 ;
        RECT 107.225 189.635 107.475 190.175 ;
        RECT 104.925 187.795 105.255 188.595 ;
        RECT 105.425 187.625 105.595 188.425 ;
        RECT 105.765 187.795 106.095 188.595 ;
        RECT 106.795 188.495 106.965 189.525 ;
        RECT 107.645 189.470 107.865 189.955 ;
        RECT 107.135 188.875 107.365 189.270 ;
        RECT 107.535 189.045 107.865 189.470 ;
        RECT 108.035 189.795 108.925 189.965 ;
        RECT 110.015 189.795 110.905 189.965 ;
        RECT 108.035 189.070 108.205 189.795 ;
        RECT 108.375 189.240 108.925 189.625 ;
        RECT 110.015 189.240 110.565 189.625 ;
        RECT 110.735 189.070 110.905 189.795 ;
        RECT 108.035 189.000 108.925 189.070 ;
        RECT 108.030 188.975 108.925 189.000 ;
        RECT 108.020 188.960 108.925 188.975 ;
        RECT 108.015 188.945 108.925 188.960 ;
        RECT 108.005 188.940 108.925 188.945 ;
        RECT 108.000 188.930 108.925 188.940 ;
        RECT 107.995 188.920 108.925 188.930 ;
        RECT 107.985 188.915 108.925 188.920 ;
        RECT 107.975 188.905 108.925 188.915 ;
        RECT 107.965 188.900 108.925 188.905 ;
        RECT 107.965 188.895 108.300 188.900 ;
        RECT 107.950 188.890 108.300 188.895 ;
        RECT 107.935 188.880 108.300 188.890 ;
        RECT 107.910 188.875 108.300 188.880 ;
        RECT 107.135 188.870 108.300 188.875 ;
        RECT 107.135 188.835 108.270 188.870 ;
        RECT 107.135 188.810 108.235 188.835 ;
        RECT 107.135 188.780 108.205 188.810 ;
        RECT 107.135 188.750 108.185 188.780 ;
        RECT 107.135 188.720 108.165 188.750 ;
        RECT 107.135 188.710 108.095 188.720 ;
        RECT 107.135 188.700 108.070 188.710 ;
        RECT 107.135 188.685 108.050 188.700 ;
        RECT 107.135 188.670 108.030 188.685 ;
        RECT 107.240 188.660 108.025 188.670 ;
        RECT 107.240 188.625 108.010 188.660 ;
        RECT 106.265 187.625 106.520 188.425 ;
        RECT 106.795 187.795 107.070 188.495 ;
        RECT 107.240 188.375 107.995 188.625 ;
        RECT 108.165 188.305 108.495 188.550 ;
        RECT 108.665 188.450 108.925 188.900 ;
        RECT 110.015 189.000 110.905 189.070 ;
        RECT 111.075 189.470 111.295 189.955 ;
        RECT 111.465 189.635 111.715 190.175 ;
        RECT 111.885 189.525 112.145 190.005 ;
        RECT 111.075 189.045 111.405 189.470 ;
        RECT 110.015 188.975 110.910 189.000 ;
        RECT 110.015 188.960 110.920 188.975 ;
        RECT 110.015 188.945 110.925 188.960 ;
        RECT 110.015 188.940 110.935 188.945 ;
        RECT 110.015 188.930 110.940 188.940 ;
        RECT 110.015 188.920 110.945 188.930 ;
        RECT 110.015 188.915 110.955 188.920 ;
        RECT 110.015 188.905 110.965 188.915 ;
        RECT 110.015 188.900 110.975 188.905 ;
        RECT 110.015 188.450 110.275 188.900 ;
        RECT 110.640 188.895 110.975 188.900 ;
        RECT 110.640 188.890 110.990 188.895 ;
        RECT 110.640 188.880 111.005 188.890 ;
        RECT 110.640 188.875 111.030 188.880 ;
        RECT 111.575 188.875 111.805 189.270 ;
        RECT 110.640 188.870 111.805 188.875 ;
        RECT 110.670 188.835 111.805 188.870 ;
        RECT 110.705 188.810 111.805 188.835 ;
        RECT 110.735 188.780 111.805 188.810 ;
        RECT 110.755 188.750 111.805 188.780 ;
        RECT 110.775 188.720 111.805 188.750 ;
        RECT 110.845 188.710 111.805 188.720 ;
        RECT 110.870 188.700 111.805 188.710 ;
        RECT 110.890 188.685 111.805 188.700 ;
        RECT 110.910 188.670 111.805 188.685 ;
        RECT 110.915 188.660 111.700 188.670 ;
        RECT 110.930 188.625 111.700 188.660 ;
        RECT 108.310 188.280 108.495 188.305 ;
        RECT 110.445 188.305 110.775 188.550 ;
        RECT 110.945 188.375 111.700 188.625 ;
        RECT 111.975 188.495 112.145 189.525 ;
        RECT 112.315 189.355 112.575 190.175 ;
        RECT 112.745 189.355 113.075 189.775 ;
        RECT 113.255 189.690 114.045 189.955 ;
        RECT 112.825 189.265 113.075 189.355 ;
        RECT 110.445 188.280 110.630 188.305 ;
        RECT 108.310 188.180 108.925 188.280 ;
        RECT 107.240 187.625 107.495 188.170 ;
        RECT 107.665 187.795 108.145 188.135 ;
        RECT 108.320 187.625 108.925 188.180 ;
        RECT 110.015 188.180 110.630 188.280 ;
        RECT 110.015 187.625 110.620 188.180 ;
        RECT 110.795 187.795 111.275 188.135 ;
        RECT 111.445 187.625 111.700 188.170 ;
        RECT 111.870 187.795 112.145 188.495 ;
        RECT 112.315 188.305 112.655 189.185 ;
        RECT 112.825 189.015 113.620 189.265 ;
        RECT 112.315 187.625 112.575 188.135 ;
        RECT 112.825 187.795 112.995 189.015 ;
        RECT 113.790 188.835 114.045 189.690 ;
        RECT 114.215 189.535 114.415 189.955 ;
        RECT 114.605 189.715 114.935 190.175 ;
        RECT 114.215 189.015 114.625 189.535 ;
        RECT 115.105 189.525 115.365 190.005 ;
        RECT 114.795 188.835 115.025 189.265 ;
        RECT 113.235 188.665 115.025 188.835 ;
        RECT 113.235 188.300 113.485 188.665 ;
        RECT 113.655 188.305 113.985 188.495 ;
        RECT 114.205 188.370 114.920 188.665 ;
        RECT 115.195 188.495 115.365 189.525 ;
        RECT 116.455 189.450 116.745 190.175 ;
        RECT 116.915 189.630 122.260 190.175 ;
        RECT 118.500 188.800 118.840 189.630 ;
        RECT 122.435 189.405 124.105 190.175 ;
        RECT 124.825 189.625 124.995 189.915 ;
        RECT 125.165 189.795 125.495 190.175 ;
        RECT 124.825 189.455 125.490 189.625 ;
        RECT 113.655 188.130 113.850 188.305 ;
        RECT 113.235 187.625 113.850 188.130 ;
        RECT 114.020 187.795 114.495 188.135 ;
        RECT 114.665 187.625 114.880 188.170 ;
        RECT 115.090 187.795 115.365 188.495 ;
        RECT 116.455 187.625 116.745 188.790 ;
        RECT 120.320 188.060 120.670 189.310 ;
        RECT 122.435 188.885 123.185 189.405 ;
        RECT 123.355 188.715 124.105 189.235 ;
        RECT 116.915 187.625 122.260 188.060 ;
        RECT 122.435 187.625 124.105 188.715 ;
        RECT 124.740 188.635 125.090 189.285 ;
        RECT 125.260 188.465 125.490 189.455 ;
        RECT 124.825 188.295 125.490 188.465 ;
        RECT 124.825 187.795 124.995 188.295 ;
        RECT 125.165 187.625 125.495 188.125 ;
        RECT 125.665 187.795 125.850 189.915 ;
        RECT 126.105 189.715 126.355 190.175 ;
        RECT 126.525 189.725 126.860 189.895 ;
        RECT 127.055 189.725 127.730 189.895 ;
        RECT 126.525 189.585 126.695 189.725 ;
        RECT 126.020 188.595 126.300 189.545 ;
        RECT 126.470 189.455 126.695 189.585 ;
        RECT 126.470 188.350 126.640 189.455 ;
        RECT 126.865 189.305 127.390 189.525 ;
        RECT 126.810 188.540 127.050 189.135 ;
        RECT 127.220 188.605 127.390 189.305 ;
        RECT 127.560 188.945 127.730 189.725 ;
        RECT 128.050 189.675 128.420 190.175 ;
        RECT 128.600 189.725 129.005 189.895 ;
        RECT 129.175 189.725 129.960 189.895 ;
        RECT 128.600 189.495 128.770 189.725 ;
        RECT 127.940 189.195 128.770 189.495 ;
        RECT 129.155 189.225 129.620 189.555 ;
        RECT 127.940 189.165 128.140 189.195 ;
        RECT 128.260 188.945 128.430 189.015 ;
        RECT 127.560 188.775 128.430 188.945 ;
        RECT 127.920 188.685 128.430 188.775 ;
        RECT 126.470 188.220 126.775 188.350 ;
        RECT 127.220 188.240 127.750 188.605 ;
        RECT 126.090 187.625 126.355 188.085 ;
        RECT 126.525 187.795 126.775 188.220 ;
        RECT 127.920 188.070 128.090 188.685 ;
        RECT 126.985 187.900 128.090 188.070 ;
        RECT 128.260 187.625 128.430 188.425 ;
        RECT 128.600 188.125 128.770 189.195 ;
        RECT 128.940 188.295 129.130 189.015 ;
        RECT 129.300 188.265 129.620 189.225 ;
        RECT 129.790 189.265 129.960 189.725 ;
        RECT 130.235 189.645 130.445 190.175 ;
        RECT 130.705 189.435 131.035 189.960 ;
        RECT 131.205 189.565 131.375 190.175 ;
        RECT 131.545 189.520 131.875 189.955 ;
        RECT 131.545 189.435 131.925 189.520 ;
        RECT 130.835 189.265 131.035 189.435 ;
        RECT 131.700 189.395 131.925 189.435 ;
        RECT 129.790 188.935 130.665 189.265 ;
        RECT 130.835 188.935 131.585 189.265 ;
        RECT 128.600 187.795 128.850 188.125 ;
        RECT 129.790 188.095 129.960 188.935 ;
        RECT 130.835 188.730 131.025 188.935 ;
        RECT 131.755 188.815 131.925 189.395 ;
        RECT 131.710 188.765 131.925 188.815 ;
        RECT 130.130 188.355 131.025 188.730 ;
        RECT 131.535 188.685 131.925 188.765 ;
        RECT 132.095 189.435 132.480 190.005 ;
        RECT 132.650 189.715 132.975 190.175 ;
        RECT 133.495 189.545 133.775 190.005 ;
        RECT 132.095 188.765 132.375 189.435 ;
        RECT 132.650 189.375 133.775 189.545 ;
        RECT 132.650 189.265 133.100 189.375 ;
        RECT 132.545 188.935 133.100 189.265 ;
        RECT 133.965 189.205 134.365 190.005 ;
        RECT 134.765 189.715 135.035 190.175 ;
        RECT 135.205 189.545 135.490 190.005 ;
        RECT 129.075 187.925 129.960 188.095 ;
        RECT 130.140 187.625 130.455 188.125 ;
        RECT 130.685 187.795 131.025 188.355 ;
        RECT 131.195 187.625 131.365 188.635 ;
        RECT 131.535 187.840 131.865 188.685 ;
        RECT 132.095 187.795 132.480 188.765 ;
        RECT 132.650 188.475 133.100 188.935 ;
        RECT 133.270 188.645 134.365 189.205 ;
        RECT 132.650 188.255 133.775 188.475 ;
        RECT 132.650 187.625 132.975 188.085 ;
        RECT 133.495 187.795 133.775 188.255 ;
        RECT 133.965 187.795 134.365 188.645 ;
        RECT 134.535 189.375 135.490 189.545 ;
        RECT 135.865 189.625 136.035 190.005 ;
        RECT 136.250 189.795 136.580 190.175 ;
        RECT 135.865 189.455 136.580 189.625 ;
        RECT 134.535 188.475 134.745 189.375 ;
        RECT 134.915 188.645 135.605 189.205 ;
        RECT 135.775 188.905 136.130 189.275 ;
        RECT 136.410 189.265 136.580 189.455 ;
        RECT 136.750 189.430 137.005 190.005 ;
        RECT 136.410 188.935 136.665 189.265 ;
        RECT 136.410 188.725 136.580 188.935 ;
        RECT 135.865 188.555 136.580 188.725 ;
        RECT 136.835 188.700 137.005 189.430 ;
        RECT 137.180 189.335 137.440 190.175 ;
        RECT 137.615 189.425 138.825 190.175 ;
        RECT 134.535 188.255 135.490 188.475 ;
        RECT 134.765 187.625 135.035 188.085 ;
        RECT 135.205 187.795 135.490 188.255 ;
        RECT 135.865 187.795 136.035 188.555 ;
        RECT 136.250 187.625 136.580 188.385 ;
        RECT 136.750 187.795 137.005 188.700 ;
        RECT 137.180 187.625 137.440 188.775 ;
        RECT 137.615 188.715 138.135 189.255 ;
        RECT 138.305 188.885 138.825 189.425 ;
        RECT 137.615 187.625 138.825 188.715 ;
        RECT 13.330 187.455 138.910 187.625 ;
        RECT 13.415 186.365 14.625 187.455 ;
        RECT 14.795 186.365 18.305 187.455 ;
        RECT 13.415 185.655 13.935 186.195 ;
        RECT 14.105 185.825 14.625 186.365 ;
        RECT 14.795 185.675 16.445 186.195 ;
        RECT 16.615 185.845 18.305 186.365 ;
        RECT 18.475 186.315 18.735 187.285 ;
        RECT 18.930 187.045 19.260 187.455 ;
        RECT 19.460 186.865 19.630 187.285 ;
        RECT 19.845 187.045 20.515 187.455 ;
        RECT 20.750 186.865 20.920 187.285 ;
        RECT 21.225 187.015 21.555 187.455 ;
        RECT 18.905 186.695 20.920 186.865 ;
        RECT 21.725 186.835 21.900 187.285 ;
        RECT 13.415 184.905 14.625 185.655 ;
        RECT 14.795 184.905 18.305 185.675 ;
        RECT 18.475 185.625 18.645 186.315 ;
        RECT 18.905 186.145 19.075 186.695 ;
        RECT 18.815 185.815 19.075 186.145 ;
        RECT 18.475 185.160 18.815 185.625 ;
        RECT 19.245 185.485 19.585 186.515 ;
        RECT 19.775 186.095 20.045 186.515 ;
        RECT 19.775 185.925 20.085 186.095 ;
        RECT 18.480 185.115 18.815 185.160 ;
        RECT 18.985 184.905 19.315 185.285 ;
        RECT 19.775 185.240 20.045 185.925 ;
        RECT 20.270 185.240 20.550 186.515 ;
        RECT 20.750 185.405 20.920 186.695 ;
        RECT 21.270 186.665 21.900 186.835 ;
        RECT 21.270 186.145 21.440 186.665 ;
        RECT 21.090 185.815 21.440 186.145 ;
        RECT 21.620 185.815 21.985 186.495 ;
        RECT 22.155 186.365 25.665 187.455 ;
        RECT 21.270 185.645 21.440 185.815 ;
        RECT 22.155 185.675 23.805 186.195 ;
        RECT 23.975 185.845 25.665 186.365 ;
        RECT 26.295 186.290 26.585 187.455 ;
        RECT 26.755 186.365 30.265 187.455 ;
        RECT 26.755 185.675 28.405 186.195 ;
        RECT 28.575 185.845 30.265 186.365 ;
        RECT 30.905 186.315 31.235 187.455 ;
        RECT 31.765 186.485 32.095 187.270 ;
        RECT 31.415 186.315 32.095 186.485 ;
        RECT 32.285 186.505 32.560 187.275 ;
        RECT 32.730 186.845 33.060 187.275 ;
        RECT 33.230 187.015 33.425 187.455 ;
        RECT 33.605 186.845 33.935 187.275 ;
        RECT 34.120 187.075 34.455 187.455 ;
        RECT 32.730 186.675 33.935 186.845 ;
        RECT 32.285 186.315 32.870 186.505 ;
        RECT 33.040 186.345 33.935 186.675 ;
        RECT 30.895 185.895 31.245 186.145 ;
        RECT 31.415 185.715 31.585 186.315 ;
        RECT 31.755 185.895 32.105 186.145 ;
        RECT 21.270 185.475 21.900 185.645 ;
        RECT 20.750 185.075 20.980 185.405 ;
        RECT 21.225 184.905 21.555 185.285 ;
        RECT 21.725 185.075 21.900 185.475 ;
        RECT 22.155 184.905 25.665 185.675 ;
        RECT 26.295 184.905 26.585 185.630 ;
        RECT 26.755 184.905 30.265 185.675 ;
        RECT 30.905 184.905 31.175 185.715 ;
        RECT 31.345 185.075 31.675 185.715 ;
        RECT 31.845 184.905 32.085 185.715 ;
        RECT 32.285 185.495 32.525 186.145 ;
        RECT 32.695 185.645 32.870 186.315 ;
        RECT 33.040 185.815 33.455 186.145 ;
        RECT 33.635 185.815 33.930 186.145 ;
        RECT 32.695 185.465 33.025 185.645 ;
        RECT 32.300 184.905 32.630 185.295 ;
        RECT 32.800 185.085 33.025 185.465 ;
        RECT 33.225 185.195 33.455 185.815 ;
        RECT 33.635 184.905 33.935 185.635 ;
        RECT 34.115 185.585 34.355 186.895 ;
        RECT 34.625 186.485 34.875 187.285 ;
        RECT 35.095 186.735 35.425 187.455 ;
        RECT 35.610 186.485 35.860 187.285 ;
        RECT 36.325 186.655 36.655 187.455 ;
        RECT 36.825 187.025 37.165 187.285 ;
        RECT 34.525 186.315 36.715 186.485 ;
        RECT 34.525 185.405 34.695 186.315 ;
        RECT 36.400 186.145 36.715 186.315 ;
        RECT 34.200 185.075 34.695 185.405 ;
        RECT 34.915 185.180 35.265 186.145 ;
        RECT 35.445 185.175 35.745 186.145 ;
        RECT 35.925 185.175 36.205 186.145 ;
        RECT 36.400 185.895 36.730 186.145 ;
        RECT 36.385 184.905 36.655 185.705 ;
        RECT 36.905 185.625 37.165 187.025 ;
        RECT 37.345 186.315 37.675 187.455 ;
        RECT 38.205 186.485 38.535 187.270 ;
        RECT 37.855 186.315 38.535 186.485 ;
        RECT 38.725 186.485 39.055 187.270 ;
        RECT 38.725 186.315 39.405 186.485 ;
        RECT 39.585 186.315 39.915 187.455 ;
        RECT 40.095 187.020 45.440 187.455 ;
        RECT 37.335 185.895 37.685 186.145 ;
        RECT 37.855 185.715 38.025 186.315 ;
        RECT 38.195 185.895 38.545 186.145 ;
        RECT 38.715 185.895 39.065 186.145 ;
        RECT 39.235 185.715 39.405 186.315 ;
        RECT 39.575 185.895 39.925 186.145 ;
        RECT 36.825 185.115 37.165 185.625 ;
        RECT 37.345 184.905 37.615 185.715 ;
        RECT 37.785 185.075 38.115 185.715 ;
        RECT 38.285 184.905 38.525 185.715 ;
        RECT 38.735 184.905 38.975 185.715 ;
        RECT 39.145 185.075 39.475 185.715 ;
        RECT 39.645 184.905 39.915 185.715 ;
        RECT 41.680 185.450 42.020 186.280 ;
        RECT 43.500 185.770 43.850 187.020 ;
        RECT 45.700 186.835 45.875 187.285 ;
        RECT 46.045 187.015 46.375 187.455 ;
        RECT 46.680 186.865 46.850 187.285 ;
        RECT 47.085 187.045 47.755 187.455 ;
        RECT 47.970 186.865 48.140 187.285 ;
        RECT 48.340 187.045 48.670 187.455 ;
        RECT 45.700 186.665 46.330 186.835 ;
        RECT 45.615 185.815 45.980 186.495 ;
        RECT 46.160 186.145 46.330 186.665 ;
        RECT 46.680 186.695 48.695 186.865 ;
        RECT 46.160 185.815 46.510 186.145 ;
        RECT 46.160 185.645 46.330 185.815 ;
        RECT 45.700 185.475 46.330 185.645 ;
        RECT 40.095 184.905 45.440 185.450 ;
        RECT 45.700 185.075 45.875 185.475 ;
        RECT 46.680 185.405 46.850 186.695 ;
        RECT 46.045 184.905 46.375 185.285 ;
        RECT 46.620 185.075 46.850 185.405 ;
        RECT 47.050 185.240 47.330 186.515 ;
        RECT 47.555 185.415 47.825 186.515 ;
        RECT 48.015 185.485 48.355 186.515 ;
        RECT 48.525 186.145 48.695 186.695 ;
        RECT 48.865 186.315 49.125 187.285 ;
        RECT 49.305 186.485 49.635 187.270 ;
        RECT 49.305 186.315 49.985 186.485 ;
        RECT 50.165 186.315 50.495 187.455 ;
        RECT 50.675 186.365 51.885 187.455 ;
        RECT 48.525 185.815 48.785 186.145 ;
        RECT 48.955 185.625 49.125 186.315 ;
        RECT 49.295 185.895 49.645 186.145 ;
        RECT 49.815 185.715 49.985 186.315 ;
        RECT 50.155 185.895 50.505 186.145 ;
        RECT 47.515 185.245 47.825 185.415 ;
        RECT 47.555 185.240 47.825 185.245 ;
        RECT 48.285 184.905 48.615 185.285 ;
        RECT 48.785 185.160 49.125 185.625 ;
        RECT 48.785 185.115 49.120 185.160 ;
        RECT 49.315 184.905 49.555 185.715 ;
        RECT 49.725 185.075 50.055 185.715 ;
        RECT 50.225 184.905 50.495 185.715 ;
        RECT 50.675 185.655 51.195 186.195 ;
        RECT 51.365 185.825 51.885 186.365 ;
        RECT 52.055 186.290 52.345 187.455 ;
        RECT 52.515 187.020 57.860 187.455 ;
        RECT 50.675 184.905 51.885 185.655 ;
        RECT 52.055 184.905 52.345 185.630 ;
        RECT 54.100 185.450 54.440 186.280 ;
        RECT 55.920 185.770 56.270 187.020 ;
        RECT 58.965 186.395 59.295 187.245 ;
        RECT 58.965 185.630 59.155 186.395 ;
        RECT 59.465 186.315 59.715 187.455 ;
        RECT 59.905 186.815 60.155 187.235 ;
        RECT 60.385 186.985 60.715 187.455 ;
        RECT 60.945 186.815 61.195 187.235 ;
        RECT 59.905 186.645 61.195 186.815 ;
        RECT 61.375 186.815 61.705 187.245 ;
        RECT 61.375 186.645 61.830 186.815 ;
        RECT 59.895 186.145 60.110 186.475 ;
        RECT 59.325 185.815 59.635 186.145 ;
        RECT 59.805 185.815 60.110 186.145 ;
        RECT 60.285 185.815 60.570 186.475 ;
        RECT 60.765 185.815 61.030 186.475 ;
        RECT 61.245 185.815 61.490 186.475 ;
        RECT 59.465 185.645 59.635 185.815 ;
        RECT 61.660 185.645 61.830 186.645 ;
        RECT 52.515 184.905 57.860 185.450 ;
        RECT 58.965 185.120 59.295 185.630 ;
        RECT 59.465 185.475 61.830 185.645 ;
        RECT 62.175 186.315 62.560 187.285 ;
        RECT 62.730 186.995 63.055 187.455 ;
        RECT 63.575 186.825 63.855 187.285 ;
        RECT 62.730 186.605 63.855 186.825 ;
        RECT 62.175 185.645 62.455 186.315 ;
        RECT 62.730 186.145 63.180 186.605 ;
        RECT 64.045 186.435 64.445 187.285 ;
        RECT 64.845 186.995 65.115 187.455 ;
        RECT 65.285 186.825 65.570 187.285 ;
        RECT 62.625 185.815 63.180 186.145 ;
        RECT 63.350 185.875 64.445 186.435 ;
        RECT 62.730 185.705 63.180 185.815 ;
        RECT 59.465 184.905 59.795 185.305 ;
        RECT 60.845 185.135 61.175 185.475 ;
        RECT 61.345 184.905 61.675 185.305 ;
        RECT 62.175 185.075 62.560 185.645 ;
        RECT 62.730 185.535 63.855 185.705 ;
        RECT 62.730 184.905 63.055 185.365 ;
        RECT 63.575 185.075 63.855 185.535 ;
        RECT 64.045 185.075 64.445 185.875 ;
        RECT 64.615 186.605 65.570 186.825 ;
        RECT 64.615 185.705 64.825 186.605 ;
        RECT 64.995 185.875 65.685 186.435 ;
        RECT 65.855 186.315 66.240 187.285 ;
        RECT 66.410 186.995 66.735 187.455 ;
        RECT 67.255 186.825 67.535 187.285 ;
        RECT 66.410 186.605 67.535 186.825 ;
        RECT 64.615 185.535 65.570 185.705 ;
        RECT 64.845 184.905 65.115 185.365 ;
        RECT 65.285 185.075 65.570 185.535 ;
        RECT 65.855 185.645 66.135 186.315 ;
        RECT 66.410 186.145 66.860 186.605 ;
        RECT 67.725 186.435 68.125 187.285 ;
        RECT 68.525 186.995 68.795 187.455 ;
        RECT 68.965 186.825 69.250 187.285 ;
        RECT 66.305 185.815 66.860 186.145 ;
        RECT 67.030 185.875 68.125 186.435 ;
        RECT 66.410 185.705 66.860 185.815 ;
        RECT 65.855 185.075 66.240 185.645 ;
        RECT 66.410 185.535 67.535 185.705 ;
        RECT 66.410 184.905 66.735 185.365 ;
        RECT 67.255 185.075 67.535 185.535 ;
        RECT 67.725 185.075 68.125 185.875 ;
        RECT 68.295 186.605 69.250 186.825 ;
        RECT 68.295 185.705 68.505 186.605 ;
        RECT 68.675 185.875 69.365 186.435 ;
        RECT 69.535 186.315 69.815 187.455 ;
        RECT 69.985 186.305 70.315 187.285 ;
        RECT 70.485 186.315 70.745 187.455 ;
        RECT 70.915 186.315 71.175 187.455 ;
        RECT 71.345 186.305 71.675 187.285 ;
        RECT 71.845 186.315 72.125 187.455 ;
        RECT 72.295 187.020 77.640 187.455 ;
        RECT 69.545 185.875 69.880 186.145 ;
        RECT 70.050 185.755 70.220 186.305 ;
        RECT 70.390 185.895 70.725 186.145 ;
        RECT 70.935 185.895 71.270 186.145 ;
        RECT 70.050 185.705 70.225 185.755 ;
        RECT 71.440 185.705 71.610 186.305 ;
        RECT 71.780 185.875 72.115 186.145 ;
        RECT 68.295 185.535 69.250 185.705 ;
        RECT 68.525 184.905 68.795 185.365 ;
        RECT 68.965 185.075 69.250 185.535 ;
        RECT 69.535 184.905 69.845 185.705 ;
        RECT 70.050 185.075 70.745 185.705 ;
        RECT 70.915 185.075 71.610 185.705 ;
        RECT 71.815 184.905 72.125 185.705 ;
        RECT 73.880 185.450 74.220 186.280 ;
        RECT 75.700 185.770 76.050 187.020 ;
        RECT 77.815 186.290 78.105 187.455 ;
        RECT 78.390 186.825 78.675 187.285 ;
        RECT 78.845 186.995 79.115 187.455 ;
        RECT 78.390 186.605 79.345 186.825 ;
        RECT 78.275 185.875 78.965 186.435 ;
        RECT 79.135 185.705 79.345 186.605 ;
        RECT 72.295 184.905 77.640 185.450 ;
        RECT 77.815 184.905 78.105 185.630 ;
        RECT 78.390 185.535 79.345 185.705 ;
        RECT 79.515 186.435 79.915 187.285 ;
        RECT 80.105 186.825 80.385 187.285 ;
        RECT 80.905 186.995 81.230 187.455 ;
        RECT 80.105 186.605 81.230 186.825 ;
        RECT 79.515 185.875 80.610 186.435 ;
        RECT 80.780 186.145 81.230 186.605 ;
        RECT 81.400 186.315 81.785 187.285 ;
        RECT 81.955 187.020 87.300 187.455 ;
        RECT 78.390 185.075 78.675 185.535 ;
        RECT 78.845 184.905 79.115 185.365 ;
        RECT 79.515 185.075 79.915 185.875 ;
        RECT 80.780 185.815 81.335 186.145 ;
        RECT 80.780 185.705 81.230 185.815 ;
        RECT 80.105 185.535 81.230 185.705 ;
        RECT 81.505 185.645 81.785 186.315 ;
        RECT 80.105 185.075 80.385 185.535 ;
        RECT 80.905 184.905 81.230 185.365 ;
        RECT 81.400 185.075 81.785 185.645 ;
        RECT 83.540 185.450 83.880 186.280 ;
        RECT 85.360 185.770 85.710 187.020 ;
        RECT 87.935 186.315 88.195 187.455 ;
        RECT 88.365 186.305 88.695 187.285 ;
        RECT 88.865 186.315 89.145 187.455 ;
        RECT 89.325 186.315 89.655 187.455 ;
        RECT 90.185 186.485 90.515 187.270 ;
        RECT 89.835 186.315 90.515 186.485 ;
        RECT 90.695 186.365 92.365 187.455 ;
        RECT 92.625 186.835 92.795 187.265 ;
        RECT 92.965 187.005 93.295 187.455 ;
        RECT 92.625 186.605 93.300 186.835 ;
        RECT 87.955 185.895 88.290 186.145 ;
        RECT 88.460 185.705 88.630 186.305 ;
        RECT 88.800 185.875 89.135 186.145 ;
        RECT 89.315 185.895 89.665 186.145 ;
        RECT 89.835 185.715 90.005 186.315 ;
        RECT 90.175 185.895 90.525 186.145 ;
        RECT 81.955 184.905 87.300 185.450 ;
        RECT 87.935 185.075 88.630 185.705 ;
        RECT 88.835 184.905 89.145 185.705 ;
        RECT 89.325 184.905 89.595 185.715 ;
        RECT 89.765 185.075 90.095 185.715 ;
        RECT 90.265 184.905 90.505 185.715 ;
        RECT 90.695 185.675 91.445 186.195 ;
        RECT 91.615 185.845 92.365 186.365 ;
        RECT 90.695 184.905 92.365 185.675 ;
        RECT 92.595 185.585 92.895 186.435 ;
        RECT 93.065 185.955 93.300 186.605 ;
        RECT 93.470 186.295 93.755 187.240 ;
        RECT 93.935 186.985 94.620 187.455 ;
        RECT 93.930 186.465 94.625 186.775 ;
        RECT 94.800 186.400 95.105 187.185 ;
        RECT 93.470 186.145 94.330 186.295 ;
        RECT 93.470 186.125 94.755 186.145 ;
        RECT 93.065 185.625 93.600 185.955 ;
        RECT 93.770 185.765 94.755 186.125 ;
        RECT 93.065 185.475 93.285 185.625 ;
        RECT 92.540 184.905 92.875 185.410 ;
        RECT 93.045 185.100 93.285 185.475 ;
        RECT 93.770 185.430 93.940 185.765 ;
        RECT 94.930 185.595 95.105 186.400 ;
        RECT 95.355 186.315 95.565 187.455 ;
        RECT 95.735 186.305 96.065 187.285 ;
        RECT 96.235 186.315 96.465 187.455 ;
        RECT 97.175 186.315 97.405 187.455 ;
        RECT 97.575 186.305 97.905 187.285 ;
        RECT 98.075 186.315 98.285 187.455 ;
        RECT 98.515 186.365 99.725 187.455 ;
        RECT 100.395 186.995 100.610 187.455 ;
        RECT 100.780 186.825 101.110 187.285 ;
        RECT 93.565 185.235 93.940 185.430 ;
        RECT 93.565 185.090 93.735 185.235 ;
        RECT 94.300 184.905 94.695 185.400 ;
        RECT 94.865 185.075 95.105 185.595 ;
        RECT 95.355 184.905 95.565 185.725 ;
        RECT 95.735 185.705 95.985 186.305 ;
        RECT 96.155 185.895 96.485 186.145 ;
        RECT 97.155 185.895 97.485 186.145 ;
        RECT 95.735 185.075 96.065 185.705 ;
        RECT 96.235 184.905 96.465 185.725 ;
        RECT 97.175 184.905 97.405 185.725 ;
        RECT 97.655 185.705 97.905 186.305 ;
        RECT 97.575 185.075 97.905 185.705 ;
        RECT 98.075 184.905 98.285 185.725 ;
        RECT 98.515 185.655 99.035 186.195 ;
        RECT 99.205 185.825 99.725 186.365 ;
        RECT 99.940 186.655 101.110 186.825 ;
        RECT 101.280 186.655 101.530 187.455 ;
        RECT 98.515 184.905 99.725 185.655 ;
        RECT 99.940 185.365 100.310 186.655 ;
        RECT 101.740 186.485 102.020 186.645 ;
        RECT 100.685 186.315 102.020 186.485 ;
        RECT 102.195 186.365 103.405 187.455 ;
        RECT 100.685 186.145 100.855 186.315 ;
        RECT 100.480 185.895 100.855 186.145 ;
        RECT 101.025 185.895 101.500 186.135 ;
        RECT 101.670 185.895 102.020 186.135 ;
        RECT 100.685 185.725 100.855 185.895 ;
        RECT 100.685 185.555 102.020 185.725 ;
        RECT 99.940 185.075 100.690 185.365 ;
        RECT 101.200 184.905 101.530 185.365 ;
        RECT 101.750 185.345 102.020 185.555 ;
        RECT 102.195 185.655 102.715 186.195 ;
        RECT 102.885 185.825 103.405 186.365 ;
        RECT 103.575 186.290 103.865 187.455 ;
        RECT 104.035 186.365 106.625 187.455 ;
        RECT 104.035 185.675 105.245 186.195 ;
        RECT 105.415 185.845 106.625 186.365 ;
        RECT 107.255 186.585 107.530 187.285 ;
        RECT 107.700 186.910 107.955 187.455 ;
        RECT 108.125 186.945 108.605 187.285 ;
        RECT 108.780 186.900 109.385 187.455 ;
        RECT 108.770 186.800 109.385 186.900 ;
        RECT 109.645 186.835 109.815 187.265 ;
        RECT 109.985 187.005 110.315 187.455 ;
        RECT 108.770 186.775 108.955 186.800 ;
        RECT 102.195 184.905 103.405 185.655 ;
        RECT 103.575 184.905 103.865 185.630 ;
        RECT 104.035 184.905 106.625 185.675 ;
        RECT 107.255 185.555 107.425 186.585 ;
        RECT 107.700 186.455 108.455 186.705 ;
        RECT 108.625 186.530 108.955 186.775 ;
        RECT 107.700 186.420 108.470 186.455 ;
        RECT 107.700 186.410 108.485 186.420 ;
        RECT 107.595 186.395 108.490 186.410 ;
        RECT 107.595 186.380 108.510 186.395 ;
        RECT 107.595 186.370 108.530 186.380 ;
        RECT 107.595 186.360 108.555 186.370 ;
        RECT 107.595 186.330 108.625 186.360 ;
        RECT 107.595 186.300 108.645 186.330 ;
        RECT 107.595 186.270 108.665 186.300 ;
        RECT 107.595 186.245 108.695 186.270 ;
        RECT 107.595 186.210 108.730 186.245 ;
        RECT 107.595 186.205 108.760 186.210 ;
        RECT 107.595 185.810 107.825 186.205 ;
        RECT 108.370 186.200 108.760 186.205 ;
        RECT 108.395 186.190 108.760 186.200 ;
        RECT 108.410 186.185 108.760 186.190 ;
        RECT 108.425 186.180 108.760 186.185 ;
        RECT 109.125 186.180 109.385 186.630 ;
        RECT 109.645 186.605 110.320 186.835 ;
        RECT 108.425 186.175 109.385 186.180 ;
        RECT 108.435 186.165 109.385 186.175 ;
        RECT 108.445 186.160 109.385 186.165 ;
        RECT 108.455 186.150 109.385 186.160 ;
        RECT 108.460 186.140 109.385 186.150 ;
        RECT 108.465 186.135 109.385 186.140 ;
        RECT 108.475 186.120 109.385 186.135 ;
        RECT 108.480 186.105 109.385 186.120 ;
        RECT 108.490 186.080 109.385 186.105 ;
        RECT 107.995 185.610 108.325 186.035 ;
        RECT 107.255 185.075 107.515 185.555 ;
        RECT 107.685 184.905 107.935 185.445 ;
        RECT 108.105 185.125 108.325 185.610 ;
        RECT 108.495 186.010 109.385 186.080 ;
        RECT 108.495 185.285 108.665 186.010 ;
        RECT 108.835 185.455 109.385 185.840 ;
        RECT 109.615 185.585 109.915 186.435 ;
        RECT 110.085 185.955 110.320 186.605 ;
        RECT 110.490 186.295 110.775 187.240 ;
        RECT 110.955 186.985 111.640 187.455 ;
        RECT 110.950 186.465 111.645 186.775 ;
        RECT 111.820 186.400 112.125 187.185 ;
        RECT 110.490 186.145 111.350 186.295 ;
        RECT 110.490 186.125 111.775 186.145 ;
        RECT 110.085 185.625 110.620 185.955 ;
        RECT 110.790 185.765 111.775 186.125 ;
        RECT 110.085 185.475 110.305 185.625 ;
        RECT 108.495 185.115 109.385 185.285 ;
        RECT 109.560 184.905 109.895 185.410 ;
        RECT 110.065 185.100 110.305 185.475 ;
        RECT 110.790 185.430 110.960 185.765 ;
        RECT 111.950 185.595 112.125 186.400 ;
        RECT 110.585 185.235 110.960 185.430 ;
        RECT 110.585 185.090 110.755 185.235 ;
        RECT 111.320 184.905 111.715 185.400 ;
        RECT 111.885 185.075 112.125 185.595 ;
        RECT 112.335 186.400 112.640 187.185 ;
        RECT 112.820 186.985 113.505 187.455 ;
        RECT 112.815 186.465 113.510 186.775 ;
        RECT 112.335 185.595 112.510 186.400 ;
        RECT 113.685 186.295 113.970 187.240 ;
        RECT 114.145 187.005 114.475 187.455 ;
        RECT 114.645 186.835 114.815 187.265 ;
        RECT 115.075 186.945 116.265 187.235 ;
        RECT 113.110 186.145 113.970 186.295 ;
        RECT 112.685 186.125 113.970 186.145 ;
        RECT 114.140 186.605 114.815 186.835 ;
        RECT 115.095 186.605 116.265 186.775 ;
        RECT 116.435 186.655 116.715 187.455 ;
        RECT 112.685 185.765 113.670 186.125 ;
        RECT 114.140 185.955 114.375 186.605 ;
        RECT 112.335 185.075 112.575 185.595 ;
        RECT 113.500 185.430 113.670 185.765 ;
        RECT 113.840 185.625 114.375 185.955 ;
        RECT 114.155 185.475 114.375 185.625 ;
        RECT 114.545 185.585 114.845 186.435 ;
        RECT 115.095 186.315 115.420 186.605 ;
        RECT 116.095 186.485 116.265 186.605 ;
        RECT 115.590 186.145 115.785 186.435 ;
        RECT 116.095 186.315 116.755 186.485 ;
        RECT 116.925 186.315 117.200 187.285 ;
        RECT 117.380 186.315 117.700 187.455 ;
        RECT 116.585 186.145 116.755 186.315 ;
        RECT 115.075 185.815 115.420 186.145 ;
        RECT 115.590 185.815 116.415 186.145 ;
        RECT 116.585 185.815 116.860 186.145 ;
        RECT 116.585 185.645 116.755 185.815 ;
        RECT 115.090 185.475 116.755 185.645 ;
        RECT 117.030 185.580 117.200 186.315 ;
        RECT 117.880 186.145 118.075 187.195 ;
        RECT 118.255 186.605 118.585 187.285 ;
        RECT 118.785 186.655 119.040 187.455 ;
        RECT 118.255 186.325 118.605 186.605 ;
        RECT 119.305 186.525 119.475 187.285 ;
        RECT 119.690 186.695 120.020 187.455 ;
        RECT 117.440 186.095 117.700 186.145 ;
        RECT 117.435 185.925 117.700 186.095 ;
        RECT 117.440 185.815 117.700 185.925 ;
        RECT 117.880 185.815 118.265 186.145 ;
        RECT 118.435 185.945 118.605 186.325 ;
        RECT 118.795 186.115 119.040 186.475 ;
        RECT 119.305 186.355 120.020 186.525 ;
        RECT 120.190 186.380 120.445 187.285 ;
        RECT 118.435 185.775 118.955 185.945 ;
        RECT 119.215 185.805 119.570 186.175 ;
        RECT 119.850 186.145 120.020 186.355 ;
        RECT 119.850 185.815 120.105 186.145 ;
        RECT 112.745 184.905 113.140 185.400 ;
        RECT 113.500 185.235 113.875 185.430 ;
        RECT 113.705 185.090 113.875 185.235 ;
        RECT 114.155 185.100 114.395 185.475 ;
        RECT 114.565 184.905 114.900 185.410 ;
        RECT 115.090 185.125 115.345 185.475 ;
        RECT 115.515 184.905 115.845 185.305 ;
        RECT 116.015 185.125 116.185 185.475 ;
        RECT 116.355 184.905 116.735 185.305 ;
        RECT 116.925 185.235 117.200 185.580 ;
        RECT 117.380 185.435 118.595 185.605 ;
        RECT 117.380 185.085 117.670 185.435 ;
        RECT 117.865 184.905 118.195 185.265 ;
        RECT 118.365 185.130 118.595 185.435 ;
        RECT 118.785 185.415 118.955 185.775 ;
        RECT 119.850 185.625 120.020 185.815 ;
        RECT 120.275 185.650 120.445 186.380 ;
        RECT 120.620 186.305 120.880 187.455 ;
        RECT 121.055 187.020 126.400 187.455 ;
        RECT 119.305 185.455 120.020 185.625 ;
        RECT 118.785 185.245 118.985 185.415 ;
        RECT 118.785 185.210 118.955 185.245 ;
        RECT 119.305 185.075 119.475 185.455 ;
        RECT 119.690 184.905 120.020 185.285 ;
        RECT 120.190 185.075 120.445 185.650 ;
        RECT 120.620 184.905 120.880 185.745 ;
        RECT 122.640 185.450 122.980 186.280 ;
        RECT 124.460 185.770 124.810 187.020 ;
        RECT 126.575 186.365 129.165 187.455 ;
        RECT 126.575 185.675 127.785 186.195 ;
        RECT 127.955 185.845 129.165 186.365 ;
        RECT 129.335 186.290 129.625 187.455 ;
        RECT 129.800 186.315 130.135 187.285 ;
        RECT 130.305 186.315 130.475 187.455 ;
        RECT 130.645 187.115 132.675 187.285 ;
        RECT 121.055 184.905 126.400 185.450 ;
        RECT 126.575 184.905 129.165 185.675 ;
        RECT 129.800 185.645 129.970 186.315 ;
        RECT 130.645 186.145 130.815 187.115 ;
        RECT 130.140 185.815 130.395 186.145 ;
        RECT 130.620 185.815 130.815 186.145 ;
        RECT 130.985 186.775 132.110 186.945 ;
        RECT 130.225 185.645 130.395 185.815 ;
        RECT 130.985 185.645 131.155 186.775 ;
        RECT 129.335 184.905 129.625 185.630 ;
        RECT 129.800 185.075 130.055 185.645 ;
        RECT 130.225 185.475 131.155 185.645 ;
        RECT 131.325 186.435 132.335 186.605 ;
        RECT 131.325 185.635 131.495 186.435 ;
        RECT 131.700 186.095 131.975 186.235 ;
        RECT 131.695 185.925 131.975 186.095 ;
        RECT 130.980 185.440 131.155 185.475 ;
        RECT 130.225 184.905 130.555 185.305 ;
        RECT 130.980 185.075 131.510 185.440 ;
        RECT 131.700 185.075 131.975 185.925 ;
        RECT 132.145 185.075 132.335 186.435 ;
        RECT 132.505 186.450 132.675 187.115 ;
        RECT 132.845 186.695 133.015 187.455 ;
        RECT 133.250 186.695 133.765 187.105 ;
        RECT 132.505 186.260 133.255 186.450 ;
        RECT 133.425 185.885 133.765 186.695 ;
        RECT 134.025 186.525 134.195 187.285 ;
        RECT 134.410 186.695 134.740 187.455 ;
        RECT 134.025 186.355 134.740 186.525 ;
        RECT 134.910 186.380 135.165 187.285 ;
        RECT 132.535 185.715 133.765 185.885 ;
        RECT 133.935 185.805 134.290 186.175 ;
        RECT 134.570 186.145 134.740 186.355 ;
        RECT 134.570 185.815 134.825 186.145 ;
        RECT 132.515 184.905 133.025 185.440 ;
        RECT 133.245 185.110 133.490 185.715 ;
        RECT 134.570 185.625 134.740 185.815 ;
        RECT 134.995 185.650 135.165 186.380 ;
        RECT 135.340 186.305 135.600 187.455 ;
        RECT 135.865 186.525 136.035 187.285 ;
        RECT 136.250 186.695 136.580 187.455 ;
        RECT 135.865 186.355 136.580 186.525 ;
        RECT 136.750 186.380 137.005 187.285 ;
        RECT 135.775 185.805 136.130 186.175 ;
        RECT 136.410 186.145 136.580 186.355 ;
        RECT 136.410 185.815 136.665 186.145 ;
        RECT 134.025 185.455 134.740 185.625 ;
        RECT 134.025 185.075 134.195 185.455 ;
        RECT 134.410 184.905 134.740 185.285 ;
        RECT 134.910 185.075 135.165 185.650 ;
        RECT 135.340 184.905 135.600 185.745 ;
        RECT 136.410 185.625 136.580 185.815 ;
        RECT 136.835 185.650 137.005 186.380 ;
        RECT 137.180 186.305 137.440 187.455 ;
        RECT 137.615 186.365 138.825 187.455 ;
        RECT 137.615 185.825 138.135 186.365 ;
        RECT 135.865 185.455 136.580 185.625 ;
        RECT 135.865 185.075 136.035 185.455 ;
        RECT 136.250 184.905 136.580 185.285 ;
        RECT 136.750 185.075 137.005 185.650 ;
        RECT 137.180 184.905 137.440 185.745 ;
        RECT 138.305 185.655 138.825 186.195 ;
        RECT 137.615 184.905 138.825 185.655 ;
        RECT 13.330 184.735 138.910 184.905 ;
        RECT 13.415 183.985 14.625 184.735 ;
        RECT 14.885 184.185 15.055 184.565 ;
        RECT 15.235 184.355 15.565 184.735 ;
        RECT 14.885 184.015 15.550 184.185 ;
        RECT 15.745 184.060 16.005 184.565 ;
        RECT 13.415 183.445 13.935 183.985 ;
        RECT 14.105 183.275 14.625 183.815 ;
        RECT 14.815 183.465 15.145 183.835 ;
        RECT 15.380 183.760 15.550 184.015 ;
        RECT 15.380 183.430 15.665 183.760 ;
        RECT 15.380 183.285 15.550 183.430 ;
        RECT 13.415 182.185 14.625 183.275 ;
        RECT 14.885 183.115 15.550 183.285 ;
        RECT 15.835 183.260 16.005 184.060 ;
        RECT 16.175 183.965 17.845 184.735 ;
        RECT 18.105 184.185 18.275 184.475 ;
        RECT 18.445 184.355 18.775 184.735 ;
        RECT 18.105 184.015 18.770 184.185 ;
        RECT 16.175 183.445 16.925 183.965 ;
        RECT 17.095 183.275 17.845 183.795 ;
        RECT 14.885 182.355 15.055 183.115 ;
        RECT 15.235 182.185 15.565 182.945 ;
        RECT 15.735 182.355 16.005 183.260 ;
        RECT 16.175 182.185 17.845 183.275 ;
        RECT 18.020 183.195 18.370 183.845 ;
        RECT 18.540 183.025 18.770 184.015 ;
        RECT 18.105 182.855 18.770 183.025 ;
        RECT 18.105 182.355 18.275 182.855 ;
        RECT 18.445 182.185 18.775 182.685 ;
        RECT 18.945 182.355 19.130 184.475 ;
        RECT 19.385 184.275 19.635 184.735 ;
        RECT 19.805 184.285 20.140 184.455 ;
        RECT 20.335 184.285 21.010 184.455 ;
        RECT 19.805 184.145 19.975 184.285 ;
        RECT 19.300 183.155 19.580 184.105 ;
        RECT 19.750 184.015 19.975 184.145 ;
        RECT 19.750 182.910 19.920 184.015 ;
        RECT 20.145 183.865 20.670 184.085 ;
        RECT 20.090 183.100 20.330 183.695 ;
        RECT 20.500 183.165 20.670 183.865 ;
        RECT 20.840 183.505 21.010 184.285 ;
        RECT 21.330 184.235 21.700 184.735 ;
        RECT 21.880 184.285 22.285 184.455 ;
        RECT 22.455 184.285 23.240 184.455 ;
        RECT 21.880 184.055 22.050 184.285 ;
        RECT 21.220 183.755 22.050 184.055 ;
        RECT 22.435 183.785 22.900 184.115 ;
        RECT 21.220 183.725 21.420 183.755 ;
        RECT 21.540 183.505 21.710 183.575 ;
        RECT 20.840 183.335 21.710 183.505 ;
        RECT 21.200 183.245 21.710 183.335 ;
        RECT 19.750 182.780 20.055 182.910 ;
        RECT 20.500 182.800 21.030 183.165 ;
        RECT 19.370 182.185 19.635 182.645 ;
        RECT 19.805 182.355 20.055 182.780 ;
        RECT 21.200 182.630 21.370 183.245 ;
        RECT 20.265 182.460 21.370 182.630 ;
        RECT 21.540 182.185 21.710 182.985 ;
        RECT 21.880 182.685 22.050 183.755 ;
        RECT 22.220 182.855 22.410 183.575 ;
        RECT 22.580 182.825 22.900 183.785 ;
        RECT 23.070 183.825 23.240 184.285 ;
        RECT 23.515 184.205 23.725 184.735 ;
        RECT 23.985 183.995 24.315 184.520 ;
        RECT 24.485 184.125 24.655 184.735 ;
        RECT 24.825 184.080 25.155 184.515 ;
        RECT 24.825 183.995 25.205 184.080 ;
        RECT 24.115 183.825 24.315 183.995 ;
        RECT 24.980 183.955 25.205 183.995 ;
        RECT 23.070 183.495 23.945 183.825 ;
        RECT 24.115 183.495 24.865 183.825 ;
        RECT 21.880 182.355 22.130 182.685 ;
        RECT 23.070 182.655 23.240 183.495 ;
        RECT 24.115 183.290 24.305 183.495 ;
        RECT 25.035 183.375 25.205 183.955 ;
        RECT 25.395 183.925 25.635 184.735 ;
        RECT 25.805 183.925 26.135 184.565 ;
        RECT 26.305 183.925 26.575 184.735 ;
        RECT 26.755 184.190 32.100 184.735 ;
        RECT 32.275 184.190 37.620 184.735 ;
        RECT 25.375 183.495 25.725 183.745 ;
        RECT 24.990 183.325 25.205 183.375 ;
        RECT 25.895 183.325 26.065 183.925 ;
        RECT 26.235 183.495 26.585 183.745 ;
        RECT 28.340 183.360 28.680 184.190 ;
        RECT 23.410 182.915 24.305 183.290 ;
        RECT 24.815 183.245 25.205 183.325 ;
        RECT 22.355 182.485 23.240 182.655 ;
        RECT 23.420 182.185 23.735 182.685 ;
        RECT 23.965 182.355 24.305 182.915 ;
        RECT 24.475 182.185 24.645 183.195 ;
        RECT 24.815 182.400 25.145 183.245 ;
        RECT 25.385 183.155 26.065 183.325 ;
        RECT 25.385 182.370 25.715 183.155 ;
        RECT 26.245 182.185 26.575 183.325 ;
        RECT 30.160 182.620 30.510 183.870 ;
        RECT 33.860 183.360 34.200 184.190 ;
        RECT 37.795 183.985 39.005 184.735 ;
        RECT 39.175 184.010 39.465 184.735 ;
        RECT 35.680 182.620 36.030 183.870 ;
        RECT 37.795 183.445 38.315 183.985 ;
        RECT 39.635 183.965 41.305 184.735 ;
        RECT 41.945 184.005 42.245 184.735 ;
        RECT 38.485 183.275 39.005 183.815 ;
        RECT 39.635 183.445 40.385 183.965 ;
        RECT 42.425 183.825 42.655 184.445 ;
        RECT 42.855 184.175 43.080 184.555 ;
        RECT 43.250 184.345 43.580 184.735 ;
        RECT 43.775 184.355 44.665 184.525 ;
        RECT 42.855 183.995 43.185 184.175 ;
        RECT 26.755 182.185 32.100 182.620 ;
        RECT 32.275 182.185 37.620 182.620 ;
        RECT 37.795 182.185 39.005 183.275 ;
        RECT 39.175 182.185 39.465 183.350 ;
        RECT 40.555 183.275 41.305 183.795 ;
        RECT 41.950 183.495 42.245 183.825 ;
        RECT 42.425 183.495 42.840 183.825 ;
        RECT 43.010 183.325 43.185 183.995 ;
        RECT 43.355 183.495 43.595 184.145 ;
        RECT 43.775 183.800 44.325 184.185 ;
        RECT 44.495 183.630 44.665 184.355 ;
        RECT 43.775 183.560 44.665 183.630 ;
        RECT 44.835 184.030 45.055 184.515 ;
        RECT 45.225 184.195 45.475 184.735 ;
        RECT 45.645 184.085 45.905 184.565 ;
        RECT 44.835 183.605 45.165 184.030 ;
        RECT 43.775 183.535 44.670 183.560 ;
        RECT 43.775 183.520 44.680 183.535 ;
        RECT 43.775 183.505 44.685 183.520 ;
        RECT 43.775 183.500 44.695 183.505 ;
        RECT 43.775 183.490 44.700 183.500 ;
        RECT 43.775 183.480 44.705 183.490 ;
        RECT 43.775 183.475 44.715 183.480 ;
        RECT 43.775 183.465 44.725 183.475 ;
        RECT 43.775 183.460 44.735 183.465 ;
        RECT 39.635 182.185 41.305 183.275 ;
        RECT 41.945 182.965 42.840 183.295 ;
        RECT 43.010 183.135 43.595 183.325 ;
        RECT 41.945 182.795 43.150 182.965 ;
        RECT 41.945 182.365 42.275 182.795 ;
        RECT 42.455 182.185 42.650 182.625 ;
        RECT 42.820 182.365 43.150 182.795 ;
        RECT 43.320 182.365 43.595 183.135 ;
        RECT 43.775 183.010 44.035 183.460 ;
        RECT 44.400 183.455 44.735 183.460 ;
        RECT 44.400 183.450 44.750 183.455 ;
        RECT 44.400 183.440 44.765 183.450 ;
        RECT 44.400 183.435 44.790 183.440 ;
        RECT 45.335 183.435 45.565 183.830 ;
        RECT 44.400 183.430 45.565 183.435 ;
        RECT 44.430 183.395 45.565 183.430 ;
        RECT 44.465 183.370 45.565 183.395 ;
        RECT 44.495 183.340 45.565 183.370 ;
        RECT 44.515 183.310 45.565 183.340 ;
        RECT 44.535 183.280 45.565 183.310 ;
        RECT 44.605 183.270 45.565 183.280 ;
        RECT 44.630 183.260 45.565 183.270 ;
        RECT 44.650 183.245 45.565 183.260 ;
        RECT 44.670 183.230 45.565 183.245 ;
        RECT 44.675 183.220 45.460 183.230 ;
        RECT 44.690 183.185 45.460 183.220 ;
        RECT 44.205 182.865 44.535 183.110 ;
        RECT 44.705 182.935 45.460 183.185 ;
        RECT 45.735 183.055 45.905 184.085 ;
        RECT 46.165 184.185 46.335 184.475 ;
        RECT 46.505 184.355 46.835 184.735 ;
        RECT 46.165 184.015 46.830 184.185 ;
        RECT 46.080 183.195 46.430 183.845 ;
        RECT 44.205 182.840 44.390 182.865 ;
        RECT 43.775 182.740 44.390 182.840 ;
        RECT 43.775 182.185 44.380 182.740 ;
        RECT 44.555 182.355 45.035 182.695 ;
        RECT 45.205 182.185 45.460 182.730 ;
        RECT 45.630 182.355 45.905 183.055 ;
        RECT 46.600 183.025 46.830 184.015 ;
        RECT 46.165 182.855 46.830 183.025 ;
        RECT 46.165 182.355 46.335 182.855 ;
        RECT 46.505 182.185 46.835 182.685 ;
        RECT 47.005 182.355 47.190 184.475 ;
        RECT 47.445 184.275 47.695 184.735 ;
        RECT 47.865 184.285 48.200 184.455 ;
        RECT 48.395 184.285 49.070 184.455 ;
        RECT 47.865 184.145 48.035 184.285 ;
        RECT 47.360 183.155 47.640 184.105 ;
        RECT 47.810 184.015 48.035 184.145 ;
        RECT 47.810 182.910 47.980 184.015 ;
        RECT 48.205 183.865 48.730 184.085 ;
        RECT 48.150 183.100 48.390 183.695 ;
        RECT 48.560 183.165 48.730 183.865 ;
        RECT 48.900 183.505 49.070 184.285 ;
        RECT 49.390 184.235 49.760 184.735 ;
        RECT 49.940 184.285 50.345 184.455 ;
        RECT 50.515 184.285 51.300 184.455 ;
        RECT 49.940 184.055 50.110 184.285 ;
        RECT 49.280 183.755 50.110 184.055 ;
        RECT 50.495 183.785 50.960 184.115 ;
        RECT 49.280 183.725 49.480 183.755 ;
        RECT 49.600 183.505 49.770 183.575 ;
        RECT 48.900 183.335 49.770 183.505 ;
        RECT 49.260 183.245 49.770 183.335 ;
        RECT 47.810 182.780 48.115 182.910 ;
        RECT 48.560 182.800 49.090 183.165 ;
        RECT 47.430 182.185 47.695 182.645 ;
        RECT 47.865 182.355 48.115 182.780 ;
        RECT 49.260 182.630 49.430 183.245 ;
        RECT 48.325 182.460 49.430 182.630 ;
        RECT 49.600 182.185 49.770 182.985 ;
        RECT 49.940 182.685 50.110 183.755 ;
        RECT 50.280 182.855 50.470 183.575 ;
        RECT 50.640 182.825 50.960 183.785 ;
        RECT 51.130 183.825 51.300 184.285 ;
        RECT 51.575 184.205 51.785 184.735 ;
        RECT 52.045 183.995 52.375 184.520 ;
        RECT 52.545 184.125 52.715 184.735 ;
        RECT 52.885 184.080 53.215 184.515 ;
        RECT 52.885 183.995 53.265 184.080 ;
        RECT 52.175 183.825 52.375 183.995 ;
        RECT 53.040 183.955 53.265 183.995 ;
        RECT 51.130 183.495 52.005 183.825 ;
        RECT 52.175 183.495 52.925 183.825 ;
        RECT 49.940 182.355 50.190 182.685 ;
        RECT 51.130 182.655 51.300 183.495 ;
        RECT 52.175 183.290 52.365 183.495 ;
        RECT 53.095 183.375 53.265 183.955 ;
        RECT 53.435 183.965 56.945 184.735 ;
        RECT 57.665 184.185 57.835 184.475 ;
        RECT 58.005 184.355 58.335 184.735 ;
        RECT 57.665 184.015 58.330 184.185 ;
        RECT 53.435 183.445 55.085 183.965 ;
        RECT 53.050 183.325 53.265 183.375 ;
        RECT 51.470 182.915 52.365 183.290 ;
        RECT 52.875 183.245 53.265 183.325 ;
        RECT 55.255 183.275 56.945 183.795 ;
        RECT 50.415 182.485 51.300 182.655 ;
        RECT 51.480 182.185 51.795 182.685 ;
        RECT 52.025 182.355 52.365 182.915 ;
        RECT 52.535 182.185 52.705 183.195 ;
        RECT 52.875 182.400 53.205 183.245 ;
        RECT 53.435 182.185 56.945 183.275 ;
        RECT 57.580 183.195 57.930 183.845 ;
        RECT 58.100 183.025 58.330 184.015 ;
        RECT 57.665 182.855 58.330 183.025 ;
        RECT 57.665 182.355 57.835 182.855 ;
        RECT 58.005 182.185 58.335 182.685 ;
        RECT 58.505 182.355 58.690 184.475 ;
        RECT 58.945 184.275 59.195 184.735 ;
        RECT 59.365 184.285 59.700 184.455 ;
        RECT 59.895 184.285 60.570 184.455 ;
        RECT 59.365 184.145 59.535 184.285 ;
        RECT 58.860 183.155 59.140 184.105 ;
        RECT 59.310 184.015 59.535 184.145 ;
        RECT 59.310 182.910 59.480 184.015 ;
        RECT 59.705 183.865 60.230 184.085 ;
        RECT 59.650 183.100 59.890 183.695 ;
        RECT 60.060 183.165 60.230 183.865 ;
        RECT 60.400 183.505 60.570 184.285 ;
        RECT 60.890 184.235 61.260 184.735 ;
        RECT 61.440 184.285 61.845 184.455 ;
        RECT 62.015 184.285 62.800 184.455 ;
        RECT 61.440 184.055 61.610 184.285 ;
        RECT 60.780 183.755 61.610 184.055 ;
        RECT 61.995 183.785 62.460 184.115 ;
        RECT 60.780 183.725 60.980 183.755 ;
        RECT 61.100 183.505 61.270 183.575 ;
        RECT 60.400 183.335 61.270 183.505 ;
        RECT 60.760 183.245 61.270 183.335 ;
        RECT 59.310 182.780 59.615 182.910 ;
        RECT 60.060 182.800 60.590 183.165 ;
        RECT 58.930 182.185 59.195 182.645 ;
        RECT 59.365 182.355 59.615 182.780 ;
        RECT 60.760 182.630 60.930 183.245 ;
        RECT 59.825 182.460 60.930 182.630 ;
        RECT 61.100 182.185 61.270 182.985 ;
        RECT 61.440 182.685 61.610 183.755 ;
        RECT 61.780 182.855 61.970 183.575 ;
        RECT 62.140 182.825 62.460 183.785 ;
        RECT 62.630 183.825 62.800 184.285 ;
        RECT 63.075 184.205 63.285 184.735 ;
        RECT 63.545 183.995 63.875 184.520 ;
        RECT 64.045 184.125 64.215 184.735 ;
        RECT 64.385 184.080 64.715 184.515 ;
        RECT 64.385 183.995 64.765 184.080 ;
        RECT 64.935 184.010 65.225 184.735 ;
        RECT 63.675 183.825 63.875 183.995 ;
        RECT 64.540 183.955 64.765 183.995 ;
        RECT 62.630 183.495 63.505 183.825 ;
        RECT 63.675 183.495 64.425 183.825 ;
        RECT 61.440 182.355 61.690 182.685 ;
        RECT 62.630 182.655 62.800 183.495 ;
        RECT 63.675 183.290 63.865 183.495 ;
        RECT 64.595 183.375 64.765 183.955 ;
        RECT 64.550 183.325 64.765 183.375 ;
        RECT 62.970 182.915 63.865 183.290 ;
        RECT 64.375 183.245 64.765 183.325 ;
        RECT 61.915 182.485 62.800 182.655 ;
        RECT 62.980 182.185 63.295 182.685 ;
        RECT 63.525 182.355 63.865 182.915 ;
        RECT 64.035 182.185 64.205 183.195 ;
        RECT 64.375 182.400 64.705 183.245 ;
        RECT 64.935 182.185 65.225 183.350 ;
        RECT 65.405 182.365 65.665 184.555 ;
        RECT 65.925 184.365 66.595 184.735 ;
        RECT 66.775 184.185 67.085 184.555 ;
        RECT 65.855 183.985 67.085 184.185 ;
        RECT 65.855 183.315 66.145 183.985 ;
        RECT 67.265 183.805 67.495 184.445 ;
        RECT 67.675 184.005 67.965 184.735 ;
        RECT 68.245 184.185 68.415 184.475 ;
        RECT 68.585 184.355 68.915 184.735 ;
        RECT 68.245 184.015 68.910 184.185 ;
        RECT 66.325 183.495 66.790 183.805 ;
        RECT 66.970 183.495 67.495 183.805 ;
        RECT 67.675 183.495 67.975 183.825 ;
        RECT 65.855 183.095 66.625 183.315 ;
        RECT 65.835 182.185 66.175 182.915 ;
        RECT 66.355 182.365 66.625 183.095 ;
        RECT 66.805 183.075 67.965 183.315 ;
        RECT 68.160 183.195 68.510 183.845 ;
        RECT 66.805 182.365 67.035 183.075 ;
        RECT 67.205 182.185 67.535 182.895 ;
        RECT 67.705 182.365 67.965 183.075 ;
        RECT 68.680 183.025 68.910 184.015 ;
        RECT 68.245 182.855 68.910 183.025 ;
        RECT 68.245 182.355 68.415 182.855 ;
        RECT 68.585 182.185 68.915 182.685 ;
        RECT 69.085 182.355 69.270 184.475 ;
        RECT 69.525 184.275 69.775 184.735 ;
        RECT 69.945 184.285 70.280 184.455 ;
        RECT 70.475 184.285 71.150 184.455 ;
        RECT 69.945 184.145 70.115 184.285 ;
        RECT 69.440 183.155 69.720 184.105 ;
        RECT 69.890 184.015 70.115 184.145 ;
        RECT 69.890 182.910 70.060 184.015 ;
        RECT 70.285 183.865 70.810 184.085 ;
        RECT 70.230 183.100 70.470 183.695 ;
        RECT 70.640 183.165 70.810 183.865 ;
        RECT 70.980 183.505 71.150 184.285 ;
        RECT 71.470 184.235 71.840 184.735 ;
        RECT 72.020 184.285 72.425 184.455 ;
        RECT 72.595 184.285 73.380 184.455 ;
        RECT 72.020 184.055 72.190 184.285 ;
        RECT 71.360 183.755 72.190 184.055 ;
        RECT 72.575 183.785 73.040 184.115 ;
        RECT 71.360 183.725 71.560 183.755 ;
        RECT 71.680 183.505 71.850 183.575 ;
        RECT 70.980 183.335 71.850 183.505 ;
        RECT 71.340 183.245 71.850 183.335 ;
        RECT 69.890 182.780 70.195 182.910 ;
        RECT 70.640 182.800 71.170 183.165 ;
        RECT 69.510 182.185 69.775 182.645 ;
        RECT 69.945 182.355 70.195 182.780 ;
        RECT 71.340 182.630 71.510 183.245 ;
        RECT 70.405 182.460 71.510 182.630 ;
        RECT 71.680 182.185 71.850 182.985 ;
        RECT 72.020 182.685 72.190 183.755 ;
        RECT 72.360 182.855 72.550 183.575 ;
        RECT 72.720 182.825 73.040 183.785 ;
        RECT 73.210 183.825 73.380 184.285 ;
        RECT 73.655 184.205 73.865 184.735 ;
        RECT 74.125 183.995 74.455 184.520 ;
        RECT 74.625 184.125 74.795 184.735 ;
        RECT 74.965 184.080 75.295 184.515 ;
        RECT 75.565 184.080 75.895 184.515 ;
        RECT 76.065 184.125 76.235 184.735 ;
        RECT 74.965 183.995 75.345 184.080 ;
        RECT 74.255 183.825 74.455 183.995 ;
        RECT 75.120 183.955 75.345 183.995 ;
        RECT 73.210 183.495 74.085 183.825 ;
        RECT 74.255 183.495 75.005 183.825 ;
        RECT 72.020 182.355 72.270 182.685 ;
        RECT 73.210 182.655 73.380 183.495 ;
        RECT 74.255 183.290 74.445 183.495 ;
        RECT 75.175 183.375 75.345 183.955 ;
        RECT 75.130 183.325 75.345 183.375 ;
        RECT 73.550 182.915 74.445 183.290 ;
        RECT 74.955 183.245 75.345 183.325 ;
        RECT 75.515 183.995 75.895 184.080 ;
        RECT 76.405 183.995 76.735 184.520 ;
        RECT 76.995 184.205 77.205 184.735 ;
        RECT 77.480 184.285 78.265 184.455 ;
        RECT 78.435 184.285 78.840 184.455 ;
        RECT 75.515 183.955 75.740 183.995 ;
        RECT 75.515 183.375 75.685 183.955 ;
        RECT 76.405 183.825 76.605 183.995 ;
        RECT 77.480 183.825 77.650 184.285 ;
        RECT 75.855 183.495 76.605 183.825 ;
        RECT 76.775 183.495 77.650 183.825 ;
        RECT 75.515 183.325 75.730 183.375 ;
        RECT 75.515 183.245 75.905 183.325 ;
        RECT 72.495 182.485 73.380 182.655 ;
        RECT 73.560 182.185 73.875 182.685 ;
        RECT 74.105 182.355 74.445 182.915 ;
        RECT 74.615 182.185 74.785 183.195 ;
        RECT 74.955 182.400 75.285 183.245 ;
        RECT 75.575 182.400 75.905 183.245 ;
        RECT 76.415 183.290 76.605 183.495 ;
        RECT 76.075 182.185 76.245 183.195 ;
        RECT 76.415 182.915 77.310 183.290 ;
        RECT 76.415 182.355 76.755 182.915 ;
        RECT 76.985 182.185 77.300 182.685 ;
        RECT 77.480 182.655 77.650 183.495 ;
        RECT 77.820 183.785 78.285 184.115 ;
        RECT 78.670 184.055 78.840 184.285 ;
        RECT 79.020 184.235 79.390 184.735 ;
        RECT 79.710 184.285 80.385 184.455 ;
        RECT 80.580 184.285 80.915 184.455 ;
        RECT 77.820 182.825 78.140 183.785 ;
        RECT 78.670 183.755 79.500 184.055 ;
        RECT 78.310 182.855 78.500 183.575 ;
        RECT 78.670 182.685 78.840 183.755 ;
        RECT 79.300 183.725 79.500 183.755 ;
        RECT 79.010 183.505 79.180 183.575 ;
        RECT 79.710 183.505 79.880 184.285 ;
        RECT 80.745 184.145 80.915 184.285 ;
        RECT 81.085 184.275 81.335 184.735 ;
        RECT 79.010 183.335 79.880 183.505 ;
        RECT 80.050 183.865 80.575 184.085 ;
        RECT 80.745 184.015 80.970 184.145 ;
        RECT 79.010 183.245 79.520 183.335 ;
        RECT 77.480 182.485 78.365 182.655 ;
        RECT 78.590 182.355 78.840 182.685 ;
        RECT 79.010 182.185 79.180 182.985 ;
        RECT 79.350 182.630 79.520 183.245 ;
        RECT 80.050 183.165 80.220 183.865 ;
        RECT 79.690 182.800 80.220 183.165 ;
        RECT 80.390 183.100 80.630 183.695 ;
        RECT 80.800 182.910 80.970 184.015 ;
        RECT 81.140 183.155 81.420 184.105 ;
        RECT 80.665 182.780 80.970 182.910 ;
        RECT 79.350 182.460 80.455 182.630 ;
        RECT 80.665 182.355 80.915 182.780 ;
        RECT 81.085 182.185 81.350 182.645 ;
        RECT 81.590 182.355 81.775 184.475 ;
        RECT 81.945 184.355 82.275 184.735 ;
        RECT 82.445 184.185 82.615 184.475 ;
        RECT 81.950 184.015 82.615 184.185 ;
        RECT 81.950 183.025 82.180 184.015 ;
        RECT 82.875 183.995 83.260 184.565 ;
        RECT 83.430 184.275 83.755 184.735 ;
        RECT 84.275 184.105 84.555 184.565 ;
        RECT 82.350 183.195 82.700 183.845 ;
        RECT 82.875 183.325 83.155 183.995 ;
        RECT 83.430 183.935 84.555 184.105 ;
        RECT 83.430 183.825 83.880 183.935 ;
        RECT 83.325 183.495 83.880 183.825 ;
        RECT 84.745 183.765 85.145 184.565 ;
        RECT 85.545 184.275 85.815 184.735 ;
        RECT 85.985 184.105 86.270 184.565 ;
        RECT 81.950 182.855 82.615 183.025 ;
        RECT 81.945 182.185 82.275 182.685 ;
        RECT 82.445 182.355 82.615 182.855 ;
        RECT 82.875 182.355 83.260 183.325 ;
        RECT 83.430 183.035 83.880 183.495 ;
        RECT 84.050 183.205 85.145 183.765 ;
        RECT 83.430 182.815 84.555 183.035 ;
        RECT 83.430 182.185 83.755 182.645 ;
        RECT 84.275 182.355 84.555 182.815 ;
        RECT 84.745 182.355 85.145 183.205 ;
        RECT 85.315 183.935 86.270 184.105 ;
        RECT 86.555 183.965 90.065 184.735 ;
        RECT 90.695 184.010 90.985 184.735 ;
        RECT 91.155 184.190 96.500 184.735 ;
        RECT 96.675 184.190 102.020 184.735 ;
        RECT 85.315 183.035 85.525 183.935 ;
        RECT 85.695 183.205 86.385 183.765 ;
        RECT 86.555 183.445 88.205 183.965 ;
        RECT 88.375 183.275 90.065 183.795 ;
        RECT 92.740 183.360 93.080 184.190 ;
        RECT 85.315 182.815 86.270 183.035 ;
        RECT 85.545 182.185 85.815 182.645 ;
        RECT 85.985 182.355 86.270 182.815 ;
        RECT 86.555 182.185 90.065 183.275 ;
        RECT 90.695 182.185 90.985 183.350 ;
        RECT 94.560 182.620 94.910 183.870 ;
        RECT 98.260 183.360 98.600 184.190 ;
        RECT 102.195 183.965 105.705 184.735 ;
        RECT 106.335 183.995 106.825 184.565 ;
        RECT 106.995 184.165 107.225 184.565 ;
        RECT 107.395 184.335 107.815 184.735 ;
        RECT 107.985 184.165 108.155 184.565 ;
        RECT 106.995 183.995 108.155 184.165 ;
        RECT 108.325 183.995 108.775 184.735 ;
        RECT 108.945 183.995 109.385 184.555 ;
        RECT 109.575 184.225 109.815 184.735 ;
        RECT 109.985 184.225 110.275 184.565 ;
        RECT 110.505 184.225 110.820 184.735 ;
        RECT 100.080 182.620 100.430 183.870 ;
        RECT 102.195 183.445 103.845 183.965 ;
        RECT 104.015 183.275 105.705 183.795 ;
        RECT 91.155 182.185 96.500 182.620 ;
        RECT 96.675 182.185 102.020 182.620 ;
        RECT 102.195 182.185 105.705 183.275 ;
        RECT 106.335 183.325 106.505 183.995 ;
        RECT 106.675 183.495 107.080 183.825 ;
        RECT 106.335 183.155 107.105 183.325 ;
        RECT 106.345 182.185 106.675 182.985 ;
        RECT 106.855 182.525 107.105 183.155 ;
        RECT 107.295 182.695 107.545 183.825 ;
        RECT 107.745 183.495 107.990 183.825 ;
        RECT 108.175 183.545 108.565 183.825 ;
        RECT 107.745 182.695 107.945 183.495 ;
        RECT 108.735 183.375 108.905 183.825 ;
        RECT 108.115 183.205 108.905 183.375 ;
        RECT 108.115 182.525 108.285 183.205 ;
        RECT 106.855 182.355 108.285 182.525 ;
        RECT 108.455 182.185 108.770 183.035 ;
        RECT 109.075 182.985 109.385 183.995 ;
        RECT 109.615 183.885 109.815 184.055 ;
        RECT 109.620 183.495 109.815 183.885 ;
        RECT 109.985 183.325 110.165 184.225 ;
        RECT 110.990 184.165 111.160 184.435 ;
        RECT 111.330 184.335 111.660 184.735 ;
        RECT 111.860 184.205 112.150 184.555 ;
        RECT 112.345 184.375 112.675 184.735 ;
        RECT 112.845 184.205 113.075 184.510 ;
        RECT 110.335 183.495 110.745 184.055 ;
        RECT 110.990 183.995 111.685 184.165 ;
        RECT 111.860 184.035 113.075 184.205 ;
        RECT 110.915 183.325 111.085 183.825 ;
        RECT 108.945 182.355 109.385 182.985 ;
        RECT 109.625 183.155 111.085 183.325 ;
        RECT 109.625 182.980 109.985 183.155 ;
        RECT 111.255 182.985 111.685 183.995 ;
        RECT 113.265 183.865 113.435 184.430 ;
        RECT 113.720 184.335 114.050 184.735 ;
        RECT 114.220 184.165 114.390 184.435 ;
        RECT 114.560 184.225 114.875 184.735 ;
        RECT 115.105 184.225 115.395 184.565 ;
        RECT 115.565 184.225 115.805 184.735 ;
        RECT 111.920 183.715 112.180 183.825 ;
        RECT 111.915 183.545 112.180 183.715 ;
        RECT 111.920 183.495 112.180 183.545 ;
        RECT 112.360 183.495 112.745 183.825 ;
        RECT 112.915 183.695 113.435 183.865 ;
        RECT 113.695 183.995 114.390 184.165 ;
        RECT 110.570 182.185 110.740 182.985 ;
        RECT 110.910 182.815 111.685 182.985 ;
        RECT 110.910 182.355 111.240 182.815 ;
        RECT 111.410 182.185 111.580 182.645 ;
        RECT 111.860 182.185 112.180 183.325 ;
        RECT 112.360 182.445 112.555 183.495 ;
        RECT 112.915 183.315 113.085 183.695 ;
        RECT 112.735 183.035 113.085 183.315 ;
        RECT 113.275 183.165 113.520 183.525 ;
        RECT 112.735 182.355 113.065 183.035 ;
        RECT 113.695 182.985 114.125 183.995 ;
        RECT 114.295 183.325 114.465 183.825 ;
        RECT 114.635 183.495 115.045 184.055 ;
        RECT 115.215 183.325 115.395 184.225 ;
        RECT 115.565 183.885 115.765 184.055 ;
        RECT 116.455 184.010 116.745 184.735 ;
        RECT 117.120 183.955 117.620 184.565 ;
        RECT 115.565 183.495 115.760 183.885 ;
        RECT 116.915 183.495 117.265 183.745 ;
        RECT 114.295 183.155 115.755 183.325 ;
        RECT 113.265 182.185 113.520 182.985 ;
        RECT 113.695 182.815 114.470 182.985 ;
        RECT 113.800 182.185 113.970 182.645 ;
        RECT 114.140 182.355 114.470 182.815 ;
        RECT 114.640 182.185 114.810 182.985 ;
        RECT 115.395 182.980 115.755 183.155 ;
        RECT 116.455 182.185 116.745 183.350 ;
        RECT 117.450 183.325 117.620 183.955 ;
        RECT 118.250 184.085 118.580 184.565 ;
        RECT 118.750 184.275 118.975 184.735 ;
        RECT 119.145 184.085 119.475 184.565 ;
        RECT 118.250 183.915 119.475 184.085 ;
        RECT 119.665 183.935 119.915 184.735 ;
        RECT 120.085 183.935 120.425 184.565 ;
        RECT 117.790 183.545 118.120 183.745 ;
        RECT 118.290 183.545 118.620 183.745 ;
        RECT 118.790 183.545 119.210 183.745 ;
        RECT 119.385 183.575 120.080 183.745 ;
        RECT 119.385 183.325 119.555 183.575 ;
        RECT 120.250 183.325 120.425 183.935 ;
        RECT 120.600 183.915 120.875 184.735 ;
        RECT 121.045 184.095 121.375 184.565 ;
        RECT 121.545 184.265 121.715 184.735 ;
        RECT 121.885 184.095 122.215 184.565 ;
        RECT 122.385 184.265 122.675 184.735 ;
        RECT 121.045 184.085 122.215 184.095 ;
        RECT 121.045 183.915 122.645 184.085 ;
        RECT 120.600 183.545 121.320 183.745 ;
        RECT 121.490 183.545 122.260 183.745 ;
        RECT 122.430 183.375 122.645 183.915 ;
        RECT 122.895 183.965 124.565 184.735 ;
        RECT 125.285 184.185 125.455 184.565 ;
        RECT 125.635 184.355 125.965 184.735 ;
        RECT 125.285 184.015 125.950 184.185 ;
        RECT 126.145 184.060 126.405 184.565 ;
        RECT 122.895 183.445 123.645 183.965 ;
        RECT 117.120 183.155 119.555 183.325 ;
        RECT 117.120 182.355 117.450 183.155 ;
        RECT 117.620 182.185 117.950 182.985 ;
        RECT 118.250 182.355 118.580 183.155 ;
        RECT 119.225 182.185 119.475 182.985 ;
        RECT 119.745 182.185 119.915 183.325 ;
        RECT 120.085 182.355 120.425 183.325 ;
        RECT 120.600 183.155 121.715 183.365 ;
        RECT 120.600 182.355 120.875 183.155 ;
        RECT 121.045 182.185 121.375 182.985 ;
        RECT 121.545 182.525 121.715 183.155 ;
        RECT 121.885 183.205 122.665 183.375 ;
        RECT 123.815 183.275 124.565 183.795 ;
        RECT 125.215 183.465 125.545 183.835 ;
        RECT 125.780 183.760 125.950 184.015 ;
        RECT 125.780 183.430 126.065 183.760 ;
        RECT 125.780 183.285 125.950 183.430 ;
        RECT 121.885 183.155 122.645 183.205 ;
        RECT 121.885 182.695 122.215 183.155 ;
        RECT 122.385 182.525 122.685 182.985 ;
        RECT 121.545 182.355 122.685 182.525 ;
        RECT 122.895 182.185 124.565 183.275 ;
        RECT 125.285 183.115 125.950 183.285 ;
        RECT 126.235 183.260 126.405 184.060 ;
        RECT 126.665 184.185 126.835 184.475 ;
        RECT 127.005 184.355 127.335 184.735 ;
        RECT 126.665 184.015 127.330 184.185 ;
        RECT 125.285 182.355 125.455 183.115 ;
        RECT 125.635 182.185 125.965 182.945 ;
        RECT 126.135 182.355 126.405 183.260 ;
        RECT 126.580 183.195 126.930 183.845 ;
        RECT 127.100 183.025 127.330 184.015 ;
        RECT 126.665 182.855 127.330 183.025 ;
        RECT 126.665 182.355 126.835 182.855 ;
        RECT 127.005 182.185 127.335 182.685 ;
        RECT 127.505 182.355 127.690 184.475 ;
        RECT 127.945 184.275 128.195 184.735 ;
        RECT 128.365 184.285 128.700 184.455 ;
        RECT 128.895 184.285 129.570 184.455 ;
        RECT 128.365 184.145 128.535 184.285 ;
        RECT 127.860 183.155 128.140 184.105 ;
        RECT 128.310 184.015 128.535 184.145 ;
        RECT 128.310 182.910 128.480 184.015 ;
        RECT 128.705 183.865 129.230 184.085 ;
        RECT 128.650 183.100 128.890 183.695 ;
        RECT 129.060 183.165 129.230 183.865 ;
        RECT 129.400 183.505 129.570 184.285 ;
        RECT 129.890 184.235 130.260 184.735 ;
        RECT 130.440 184.285 130.845 184.455 ;
        RECT 131.015 184.285 131.800 184.455 ;
        RECT 130.440 184.055 130.610 184.285 ;
        RECT 129.780 183.755 130.610 184.055 ;
        RECT 130.995 183.785 131.460 184.115 ;
        RECT 129.780 183.725 129.980 183.755 ;
        RECT 130.100 183.505 130.270 183.575 ;
        RECT 129.400 183.335 130.270 183.505 ;
        RECT 129.760 183.245 130.270 183.335 ;
        RECT 128.310 182.780 128.615 182.910 ;
        RECT 129.060 182.800 129.590 183.165 ;
        RECT 127.930 182.185 128.195 182.645 ;
        RECT 128.365 182.355 128.615 182.780 ;
        RECT 129.760 182.630 129.930 183.245 ;
        RECT 128.825 182.460 129.930 182.630 ;
        RECT 130.100 182.185 130.270 182.985 ;
        RECT 130.440 182.685 130.610 183.755 ;
        RECT 130.780 182.855 130.970 183.575 ;
        RECT 131.140 182.825 131.460 183.785 ;
        RECT 131.630 183.825 131.800 184.285 ;
        RECT 132.075 184.205 132.285 184.735 ;
        RECT 132.545 183.995 132.875 184.520 ;
        RECT 133.045 184.125 133.215 184.735 ;
        RECT 133.385 184.080 133.715 184.515 ;
        RECT 133.385 183.995 133.765 184.080 ;
        RECT 132.675 183.825 132.875 183.995 ;
        RECT 133.540 183.955 133.765 183.995 ;
        RECT 131.630 183.495 132.505 183.825 ;
        RECT 132.675 183.495 133.425 183.825 ;
        RECT 130.440 182.355 130.690 182.685 ;
        RECT 131.630 182.655 131.800 183.495 ;
        RECT 132.675 183.290 132.865 183.495 ;
        RECT 133.595 183.375 133.765 183.955 ;
        RECT 133.550 183.325 133.765 183.375 ;
        RECT 131.970 182.915 132.865 183.290 ;
        RECT 133.375 183.245 133.765 183.325 ;
        RECT 133.935 183.995 134.320 184.565 ;
        RECT 134.490 184.275 134.815 184.735 ;
        RECT 135.335 184.105 135.615 184.565 ;
        RECT 133.935 183.325 134.215 183.995 ;
        RECT 134.490 183.935 135.615 184.105 ;
        RECT 134.490 183.825 134.940 183.935 ;
        RECT 134.385 183.495 134.940 183.825 ;
        RECT 135.805 183.765 136.205 184.565 ;
        RECT 136.605 184.275 136.875 184.735 ;
        RECT 137.045 184.105 137.330 184.565 ;
        RECT 130.915 182.485 131.800 182.655 ;
        RECT 131.980 182.185 132.295 182.685 ;
        RECT 132.525 182.355 132.865 182.915 ;
        RECT 133.035 182.185 133.205 183.195 ;
        RECT 133.375 182.400 133.705 183.245 ;
        RECT 133.935 182.355 134.320 183.325 ;
        RECT 134.490 183.035 134.940 183.495 ;
        RECT 135.110 183.205 136.205 183.765 ;
        RECT 134.490 182.815 135.615 183.035 ;
        RECT 134.490 182.185 134.815 182.645 ;
        RECT 135.335 182.355 135.615 182.815 ;
        RECT 135.805 182.355 136.205 183.205 ;
        RECT 136.375 183.935 137.330 184.105 ;
        RECT 137.615 183.985 138.825 184.735 ;
        RECT 136.375 183.035 136.585 183.935 ;
        RECT 136.755 183.205 137.445 183.765 ;
        RECT 137.615 183.275 138.135 183.815 ;
        RECT 138.305 183.445 138.825 183.985 ;
        RECT 136.375 182.815 137.330 183.035 ;
        RECT 136.605 182.185 136.875 182.645 ;
        RECT 137.045 182.355 137.330 182.815 ;
        RECT 137.615 182.185 138.825 183.275 ;
        RECT 13.330 182.015 138.910 182.185 ;
        RECT 13.415 180.925 14.625 182.015 ;
        RECT 14.795 180.925 16.465 182.015 ;
        RECT 17.185 181.345 17.355 181.845 ;
        RECT 17.525 181.515 17.855 182.015 ;
        RECT 17.185 181.175 17.850 181.345 ;
        RECT 13.415 180.215 13.935 180.755 ;
        RECT 14.105 180.385 14.625 180.925 ;
        RECT 14.795 180.235 15.545 180.755 ;
        RECT 15.715 180.405 16.465 180.925 ;
        RECT 17.100 180.355 17.450 181.005 ;
        RECT 13.415 179.465 14.625 180.215 ;
        RECT 14.795 179.465 16.465 180.235 ;
        RECT 17.620 180.185 17.850 181.175 ;
        RECT 17.185 180.015 17.850 180.185 ;
        RECT 17.185 179.725 17.355 180.015 ;
        RECT 17.525 179.465 17.855 179.845 ;
        RECT 18.025 179.725 18.210 181.845 ;
        RECT 18.450 181.555 18.715 182.015 ;
        RECT 18.885 181.420 19.135 181.845 ;
        RECT 19.345 181.570 20.450 181.740 ;
        RECT 18.830 181.290 19.135 181.420 ;
        RECT 18.380 180.095 18.660 181.045 ;
        RECT 18.830 180.185 19.000 181.290 ;
        RECT 19.170 180.505 19.410 181.100 ;
        RECT 19.580 181.035 20.110 181.400 ;
        RECT 19.580 180.335 19.750 181.035 ;
        RECT 20.280 180.955 20.450 181.570 ;
        RECT 20.620 181.215 20.790 182.015 ;
        RECT 20.960 181.515 21.210 181.845 ;
        RECT 21.435 181.545 22.320 181.715 ;
        RECT 20.280 180.865 20.790 180.955 ;
        RECT 18.830 180.055 19.055 180.185 ;
        RECT 19.225 180.115 19.750 180.335 ;
        RECT 19.920 180.695 20.790 180.865 ;
        RECT 18.465 179.465 18.715 179.925 ;
        RECT 18.885 179.915 19.055 180.055 ;
        RECT 19.920 179.915 20.090 180.695 ;
        RECT 20.620 180.625 20.790 180.695 ;
        RECT 20.300 180.445 20.500 180.475 ;
        RECT 20.960 180.445 21.130 181.515 ;
        RECT 21.300 180.625 21.490 181.345 ;
        RECT 20.300 180.145 21.130 180.445 ;
        RECT 21.660 180.415 21.980 181.375 ;
        RECT 18.885 179.745 19.220 179.915 ;
        RECT 19.415 179.745 20.090 179.915 ;
        RECT 20.410 179.465 20.780 179.965 ;
        RECT 20.960 179.915 21.130 180.145 ;
        RECT 21.515 180.085 21.980 180.415 ;
        RECT 22.150 180.705 22.320 181.545 ;
        RECT 22.500 181.515 22.815 182.015 ;
        RECT 23.045 181.285 23.385 181.845 ;
        RECT 22.490 180.910 23.385 181.285 ;
        RECT 23.555 181.005 23.725 182.015 ;
        RECT 23.195 180.705 23.385 180.910 ;
        RECT 23.895 180.955 24.225 181.800 ;
        RECT 24.465 181.045 24.795 181.830 ;
        RECT 23.895 180.875 24.285 180.955 ;
        RECT 24.465 180.875 25.145 181.045 ;
        RECT 25.325 180.875 25.655 182.015 ;
        RECT 24.070 180.825 24.285 180.875 ;
        RECT 22.150 180.375 23.025 180.705 ;
        RECT 23.195 180.375 23.945 180.705 ;
        RECT 22.150 179.915 22.320 180.375 ;
        RECT 23.195 180.205 23.395 180.375 ;
        RECT 24.115 180.245 24.285 180.825 ;
        RECT 24.455 180.455 24.805 180.705 ;
        RECT 24.975 180.275 25.145 180.875 ;
        RECT 26.295 180.850 26.585 182.015 ;
        RECT 26.755 180.925 28.425 182.015 ;
        RECT 25.315 180.455 25.665 180.705 ;
        RECT 24.060 180.205 24.285 180.245 ;
        RECT 20.960 179.745 21.365 179.915 ;
        RECT 21.535 179.745 22.320 179.915 ;
        RECT 22.595 179.465 22.805 179.995 ;
        RECT 23.065 179.680 23.395 180.205 ;
        RECT 23.905 180.120 24.285 180.205 ;
        RECT 23.565 179.465 23.735 180.075 ;
        RECT 23.905 179.685 24.235 180.120 ;
        RECT 24.475 179.465 24.715 180.275 ;
        RECT 24.885 179.635 25.215 180.275 ;
        RECT 25.385 179.465 25.655 180.275 ;
        RECT 26.755 180.235 27.505 180.755 ;
        RECT 27.675 180.405 28.425 180.925 ;
        RECT 29.145 181.085 29.315 181.845 ;
        RECT 29.530 181.255 29.860 182.015 ;
        RECT 29.145 180.915 29.860 181.085 ;
        RECT 30.030 180.940 30.285 181.845 ;
        RECT 29.055 180.365 29.410 180.735 ;
        RECT 29.690 180.705 29.860 180.915 ;
        RECT 29.690 180.375 29.945 180.705 ;
        RECT 26.295 179.465 26.585 180.190 ;
        RECT 26.755 179.465 28.425 180.235 ;
        RECT 29.690 180.185 29.860 180.375 ;
        RECT 30.115 180.210 30.285 180.940 ;
        RECT 30.460 180.865 30.720 182.015 ;
        RECT 31.395 181.555 31.610 182.015 ;
        RECT 31.780 181.385 32.110 181.845 ;
        RECT 30.940 181.215 32.110 181.385 ;
        RECT 32.280 181.215 32.530 182.015 ;
        RECT 33.205 181.295 33.535 182.015 ;
        RECT 29.145 180.015 29.860 180.185 ;
        RECT 29.145 179.635 29.315 180.015 ;
        RECT 29.530 179.465 29.860 179.845 ;
        RECT 30.030 179.635 30.285 180.210 ;
        RECT 30.460 179.465 30.720 180.305 ;
        RECT 30.940 179.925 31.310 181.215 ;
        RECT 32.740 181.045 33.020 181.205 ;
        RECT 31.685 180.875 33.020 181.045 ;
        RECT 31.685 180.705 31.855 180.875 ;
        RECT 31.480 180.455 31.855 180.705 ;
        RECT 32.025 180.455 32.500 180.695 ;
        RECT 32.670 180.455 33.020 180.695 ;
        RECT 33.195 180.655 33.425 180.995 ;
        RECT 33.715 180.655 33.930 181.770 ;
        RECT 34.125 181.070 34.455 181.845 ;
        RECT 34.625 181.240 35.335 182.015 ;
        RECT 34.125 180.855 35.275 181.070 ;
        RECT 33.195 180.455 33.525 180.655 ;
        RECT 33.715 180.475 34.165 180.655 ;
        RECT 33.835 180.455 34.165 180.475 ;
        RECT 34.335 180.455 34.805 180.685 ;
        RECT 31.685 180.285 31.855 180.455 ;
        RECT 34.990 180.285 35.275 180.855 ;
        RECT 35.505 180.410 35.785 181.845 ;
        RECT 31.685 180.115 33.020 180.285 ;
        RECT 30.940 179.635 31.690 179.925 ;
        RECT 32.200 179.465 32.530 179.925 ;
        RECT 32.750 179.905 33.020 180.115 ;
        RECT 33.195 180.095 34.375 180.285 ;
        RECT 33.195 179.635 33.535 180.095 ;
        RECT 34.045 180.015 34.375 180.095 ;
        RECT 34.565 180.095 35.275 180.285 ;
        RECT 34.565 179.955 34.865 180.095 ;
        RECT 34.550 179.945 34.865 179.955 ;
        RECT 34.540 179.935 34.865 179.945 ;
        RECT 34.530 179.930 34.865 179.935 ;
        RECT 33.705 179.465 33.875 179.925 ;
        RECT 34.525 179.920 34.865 179.930 ;
        RECT 34.520 179.915 34.865 179.920 ;
        RECT 34.515 179.905 34.865 179.915 ;
        RECT 34.510 179.900 34.865 179.905 ;
        RECT 34.505 179.635 34.865 179.900 ;
        RECT 35.105 179.465 35.275 179.925 ;
        RECT 35.445 179.635 35.785 180.410 ;
        RECT 35.955 179.745 36.235 181.845 ;
        RECT 36.425 181.255 37.210 182.015 ;
        RECT 37.605 181.185 37.990 181.845 ;
        RECT 37.605 181.085 38.015 181.185 ;
        RECT 36.405 180.875 38.015 181.085 ;
        RECT 38.315 180.995 38.515 181.785 ;
        RECT 36.405 180.275 36.680 180.875 ;
        RECT 38.185 180.825 38.515 180.995 ;
        RECT 38.685 180.835 39.005 182.015 ;
        RECT 39.230 181.145 39.515 182.015 ;
        RECT 39.685 181.385 39.945 181.845 ;
        RECT 40.120 181.555 40.375 182.015 ;
        RECT 40.545 181.385 40.805 181.845 ;
        RECT 39.685 181.215 40.805 181.385 ;
        RECT 40.975 181.215 41.285 182.015 ;
        RECT 39.685 180.965 39.945 181.215 ;
        RECT 41.455 181.045 41.765 181.845 ;
        RECT 38.185 180.705 38.365 180.825 ;
        RECT 36.850 180.455 37.205 180.705 ;
        RECT 37.400 180.655 37.865 180.705 ;
        RECT 37.395 180.485 37.865 180.655 ;
        RECT 37.400 180.455 37.865 180.485 ;
        RECT 38.035 180.455 38.365 180.705 ;
        RECT 39.190 180.795 39.945 180.965 ;
        RECT 40.735 180.875 41.765 181.045 ;
        RECT 38.540 180.455 39.005 180.655 ;
        RECT 39.190 180.285 39.595 180.795 ;
        RECT 40.735 180.625 40.905 180.875 ;
        RECT 39.765 180.455 40.905 180.625 ;
        RECT 36.405 180.095 37.655 180.275 ;
        RECT 37.290 180.025 37.655 180.095 ;
        RECT 37.825 180.075 39.005 180.245 ;
        RECT 39.190 180.115 40.840 180.285 ;
        RECT 41.075 180.135 41.425 180.705 ;
        RECT 36.465 179.465 36.635 179.925 ;
        RECT 37.825 179.855 38.155 180.075 ;
        RECT 36.905 179.675 38.155 179.855 ;
        RECT 38.325 179.465 38.495 179.905 ;
        RECT 38.665 179.660 39.005 180.075 ;
        RECT 39.235 179.465 39.515 179.945 ;
        RECT 39.685 179.725 39.945 180.115 ;
        RECT 40.120 179.465 40.375 179.945 ;
        RECT 40.545 179.725 40.840 180.115 ;
        RECT 41.595 179.965 41.765 180.875 ;
        RECT 41.020 179.465 41.295 179.945 ;
        RECT 41.465 179.635 41.765 179.965 ;
        RECT 41.935 181.295 42.395 181.845 ;
        RECT 42.585 181.295 42.915 182.015 ;
        RECT 41.935 179.925 42.185 181.295 ;
        RECT 43.115 181.125 43.415 181.675 ;
        RECT 43.585 181.345 43.865 182.015 ;
        RECT 42.475 180.955 43.415 181.125 ;
        RECT 42.475 180.705 42.645 180.955 ;
        RECT 43.785 180.705 44.050 181.065 ;
        RECT 44.755 180.955 45.085 181.800 ;
        RECT 45.255 181.005 45.425 182.015 ;
        RECT 45.595 181.285 45.935 181.845 ;
        RECT 46.165 181.515 46.480 182.015 ;
        RECT 46.660 181.545 47.545 181.715 ;
        RECT 42.355 180.375 42.645 180.705 ;
        RECT 42.815 180.455 43.155 180.705 ;
        RECT 43.375 180.455 44.050 180.705 ;
        RECT 44.695 180.875 45.085 180.955 ;
        RECT 45.595 180.910 46.490 181.285 ;
        RECT 44.695 180.825 44.910 180.875 ;
        RECT 42.475 180.285 42.645 180.375 ;
        RECT 42.475 180.095 43.865 180.285 ;
        RECT 44.695 180.245 44.865 180.825 ;
        RECT 45.595 180.705 45.785 180.910 ;
        RECT 46.660 180.705 46.830 181.545 ;
        RECT 47.770 181.515 48.020 181.845 ;
        RECT 45.035 180.375 45.785 180.705 ;
        RECT 45.955 180.375 46.830 180.705 ;
        RECT 44.695 180.205 44.920 180.245 ;
        RECT 45.585 180.205 45.785 180.375 ;
        RECT 44.695 180.120 45.075 180.205 ;
        RECT 41.935 179.635 42.495 179.925 ;
        RECT 42.665 179.465 42.915 179.925 ;
        RECT 43.535 179.735 43.865 180.095 ;
        RECT 44.745 179.685 45.075 180.120 ;
        RECT 45.245 179.465 45.415 180.075 ;
        RECT 45.585 179.680 45.915 180.205 ;
        RECT 46.175 179.465 46.385 179.995 ;
        RECT 46.660 179.915 46.830 180.375 ;
        RECT 47.000 180.415 47.320 181.375 ;
        RECT 47.490 180.625 47.680 181.345 ;
        RECT 47.850 180.445 48.020 181.515 ;
        RECT 48.190 181.215 48.360 182.015 ;
        RECT 48.530 181.570 49.635 181.740 ;
        RECT 48.530 180.955 48.700 181.570 ;
        RECT 49.845 181.420 50.095 181.845 ;
        RECT 50.265 181.555 50.530 182.015 ;
        RECT 48.870 181.035 49.400 181.400 ;
        RECT 49.845 181.290 50.150 181.420 ;
        RECT 48.190 180.865 48.700 180.955 ;
        RECT 48.190 180.695 49.060 180.865 ;
        RECT 48.190 180.625 48.360 180.695 ;
        RECT 48.480 180.445 48.680 180.475 ;
        RECT 47.000 180.085 47.465 180.415 ;
        RECT 47.850 180.145 48.680 180.445 ;
        RECT 47.850 179.915 48.020 180.145 ;
        RECT 46.660 179.745 47.445 179.915 ;
        RECT 47.615 179.745 48.020 179.915 ;
        RECT 48.200 179.465 48.570 179.965 ;
        RECT 48.890 179.915 49.060 180.695 ;
        RECT 49.230 180.335 49.400 181.035 ;
        RECT 49.570 180.505 49.810 181.100 ;
        RECT 49.230 180.115 49.755 180.335 ;
        RECT 49.980 180.185 50.150 181.290 ;
        RECT 49.925 180.055 50.150 180.185 ;
        RECT 50.320 180.095 50.600 181.045 ;
        RECT 49.925 179.915 50.095 180.055 ;
        RECT 48.890 179.745 49.565 179.915 ;
        RECT 49.760 179.745 50.095 179.915 ;
        RECT 50.265 179.465 50.515 179.925 ;
        RECT 50.770 179.725 50.955 181.845 ;
        RECT 51.125 181.515 51.455 182.015 ;
        RECT 51.625 181.345 51.795 181.845 ;
        RECT 51.130 181.175 51.795 181.345 ;
        RECT 51.130 180.185 51.360 181.175 ;
        RECT 51.530 180.355 51.880 181.005 ;
        RECT 52.055 180.850 52.345 182.015 ;
        RECT 52.515 181.585 52.855 181.845 ;
        RECT 51.130 180.015 51.795 180.185 ;
        RECT 51.125 179.465 51.455 179.845 ;
        RECT 51.625 179.725 51.795 180.015 ;
        RECT 52.055 179.465 52.345 180.190 ;
        RECT 52.515 180.185 52.775 181.585 ;
        RECT 53.025 181.215 53.355 182.015 ;
        RECT 53.820 181.045 54.070 181.845 ;
        RECT 54.255 181.295 54.585 182.015 ;
        RECT 54.805 181.045 55.055 181.845 ;
        RECT 55.225 181.635 55.560 182.015 ;
        RECT 52.965 180.875 55.155 181.045 ;
        RECT 52.965 180.705 53.280 180.875 ;
        RECT 52.950 180.455 53.280 180.705 ;
        RECT 52.515 179.675 52.855 180.185 ;
        RECT 53.025 179.465 53.295 180.265 ;
        RECT 53.475 179.735 53.755 180.705 ;
        RECT 53.935 179.735 54.235 180.705 ;
        RECT 54.415 179.740 54.765 180.705 ;
        RECT 54.985 179.965 55.155 180.875 ;
        RECT 55.325 180.145 55.565 181.455 ;
        RECT 55.735 180.925 56.945 182.015 ;
        RECT 57.205 181.345 57.375 181.845 ;
        RECT 57.545 181.515 57.875 182.015 ;
        RECT 57.205 181.175 57.870 181.345 ;
        RECT 55.735 180.215 56.255 180.755 ;
        RECT 56.425 180.385 56.945 180.925 ;
        RECT 57.120 180.355 57.470 181.005 ;
        RECT 54.985 179.635 55.480 179.965 ;
        RECT 55.735 179.465 56.945 180.215 ;
        RECT 57.640 180.185 57.870 181.175 ;
        RECT 57.205 180.015 57.870 180.185 ;
        RECT 57.205 179.725 57.375 180.015 ;
        RECT 57.545 179.465 57.875 179.845 ;
        RECT 58.045 179.725 58.230 181.845 ;
        RECT 58.470 181.555 58.735 182.015 ;
        RECT 58.905 181.420 59.155 181.845 ;
        RECT 59.365 181.570 60.470 181.740 ;
        RECT 58.850 181.290 59.155 181.420 ;
        RECT 58.400 180.095 58.680 181.045 ;
        RECT 58.850 180.185 59.020 181.290 ;
        RECT 59.190 180.505 59.430 181.100 ;
        RECT 59.600 181.035 60.130 181.400 ;
        RECT 59.600 180.335 59.770 181.035 ;
        RECT 60.300 180.955 60.470 181.570 ;
        RECT 60.640 181.215 60.810 182.015 ;
        RECT 60.980 181.515 61.230 181.845 ;
        RECT 61.455 181.545 62.340 181.715 ;
        RECT 60.300 180.865 60.810 180.955 ;
        RECT 58.850 180.055 59.075 180.185 ;
        RECT 59.245 180.115 59.770 180.335 ;
        RECT 59.940 180.695 60.810 180.865 ;
        RECT 58.485 179.465 58.735 179.925 ;
        RECT 58.905 179.915 59.075 180.055 ;
        RECT 59.940 179.915 60.110 180.695 ;
        RECT 60.640 180.625 60.810 180.695 ;
        RECT 60.320 180.445 60.520 180.475 ;
        RECT 60.980 180.445 61.150 181.515 ;
        RECT 61.320 180.625 61.510 181.345 ;
        RECT 60.320 180.145 61.150 180.445 ;
        RECT 61.680 180.415 62.000 181.375 ;
        RECT 58.905 179.745 59.240 179.915 ;
        RECT 59.435 179.745 60.110 179.915 ;
        RECT 60.430 179.465 60.800 179.965 ;
        RECT 60.980 179.915 61.150 180.145 ;
        RECT 61.535 180.085 62.000 180.415 ;
        RECT 62.170 180.705 62.340 181.545 ;
        RECT 62.520 181.515 62.835 182.015 ;
        RECT 63.065 181.285 63.405 181.845 ;
        RECT 62.510 180.910 63.405 181.285 ;
        RECT 63.575 181.005 63.745 182.015 ;
        RECT 63.215 180.705 63.405 180.910 ;
        RECT 63.915 180.955 64.245 181.800 ;
        RECT 63.915 180.875 64.305 180.955 ;
        RECT 64.475 180.875 64.755 182.015 ;
        RECT 64.090 180.825 64.305 180.875 ;
        RECT 64.925 180.865 65.255 181.845 ;
        RECT 65.425 180.875 65.685 182.015 ;
        RECT 65.855 180.925 67.065 182.015 ;
        RECT 62.170 180.375 63.045 180.705 ;
        RECT 63.215 180.375 63.965 180.705 ;
        RECT 62.170 179.915 62.340 180.375 ;
        RECT 63.215 180.205 63.415 180.375 ;
        RECT 64.135 180.245 64.305 180.825 ;
        RECT 64.485 180.435 64.820 180.705 ;
        RECT 64.990 180.265 65.160 180.865 ;
        RECT 65.330 180.455 65.665 180.705 ;
        RECT 64.080 180.205 64.305 180.245 ;
        RECT 60.980 179.745 61.385 179.915 ;
        RECT 61.555 179.745 62.340 179.915 ;
        RECT 62.615 179.465 62.825 179.995 ;
        RECT 63.085 179.680 63.415 180.205 ;
        RECT 63.925 180.120 64.305 180.205 ;
        RECT 63.585 179.465 63.755 180.075 ;
        RECT 63.925 179.685 64.255 180.120 ;
        RECT 64.475 179.465 64.785 180.265 ;
        RECT 64.990 179.635 65.685 180.265 ;
        RECT 65.855 180.215 66.375 180.755 ;
        RECT 66.545 180.385 67.065 180.925 ;
        RECT 67.235 180.875 67.620 181.845 ;
        RECT 67.790 181.555 68.115 182.015 ;
        RECT 68.635 181.385 68.915 181.845 ;
        RECT 67.790 181.165 68.915 181.385 ;
        RECT 65.855 179.465 67.065 180.215 ;
        RECT 67.235 180.205 67.515 180.875 ;
        RECT 67.790 180.705 68.240 181.165 ;
        RECT 69.105 180.995 69.505 181.845 ;
        RECT 69.905 181.555 70.175 182.015 ;
        RECT 70.345 181.385 70.630 181.845 ;
        RECT 67.685 180.375 68.240 180.705 ;
        RECT 68.410 180.435 69.505 180.995 ;
        RECT 67.790 180.265 68.240 180.375 ;
        RECT 67.235 179.635 67.620 180.205 ;
        RECT 67.790 180.095 68.915 180.265 ;
        RECT 67.790 179.465 68.115 179.925 ;
        RECT 68.635 179.635 68.915 180.095 ;
        RECT 69.105 179.635 69.505 180.435 ;
        RECT 69.675 181.165 70.630 181.385 ;
        RECT 69.675 180.265 69.885 181.165 ;
        RECT 70.055 180.435 70.745 180.995 ;
        RECT 70.915 180.875 71.300 181.835 ;
        RECT 71.515 181.215 71.805 182.015 ;
        RECT 71.975 181.675 73.340 181.845 ;
        RECT 71.975 181.045 72.145 181.675 ;
        RECT 71.470 180.875 72.145 181.045 ;
        RECT 69.675 180.095 70.630 180.265 ;
        RECT 69.905 179.465 70.175 179.925 ;
        RECT 70.345 179.635 70.630 180.095 ;
        RECT 70.915 180.205 71.090 180.875 ;
        RECT 71.470 180.705 71.640 180.875 ;
        RECT 72.315 180.705 72.640 181.505 ;
        RECT 73.010 181.465 73.340 181.675 ;
        RECT 73.010 181.215 73.965 181.465 ;
        RECT 71.275 180.455 71.640 180.705 ;
        RECT 71.835 180.455 72.085 180.705 ;
        RECT 71.275 180.375 71.465 180.455 ;
        RECT 71.835 180.375 72.005 180.455 ;
        RECT 72.295 180.375 72.640 180.705 ;
        RECT 72.810 180.375 73.085 181.040 ;
        RECT 73.270 180.375 73.625 181.040 ;
        RECT 73.795 180.205 73.965 181.215 ;
        RECT 74.135 180.875 74.425 182.015 ;
        RECT 74.595 180.875 74.870 181.845 ;
        RECT 75.080 181.215 75.360 182.015 ;
        RECT 75.530 181.505 77.145 181.835 ;
        RECT 75.530 181.165 76.705 181.335 ;
        RECT 75.530 181.045 75.700 181.165 ;
        RECT 75.040 180.875 75.700 181.045 ;
        RECT 74.150 180.375 74.425 180.705 ;
        RECT 70.915 179.635 71.425 180.205 ;
        RECT 71.970 180.035 73.370 180.205 ;
        RECT 71.595 179.465 71.765 180.025 ;
        RECT 71.970 179.635 72.300 180.035 ;
        RECT 72.475 179.465 72.805 179.865 ;
        RECT 73.040 179.845 73.370 180.035 ;
        RECT 73.540 180.015 73.965 180.205 ;
        RECT 74.595 180.140 74.765 180.875 ;
        RECT 75.040 180.705 75.210 180.875 ;
        RECT 75.960 180.705 76.205 180.995 ;
        RECT 76.375 180.875 76.705 181.165 ;
        RECT 76.965 180.705 77.135 181.265 ;
        RECT 77.385 180.875 77.645 182.015 ;
        RECT 77.815 180.850 78.105 182.015 ;
        RECT 78.735 181.255 79.250 181.665 ;
        RECT 79.485 181.255 79.655 182.015 ;
        RECT 79.825 181.675 81.855 181.845 ;
        RECT 74.935 180.375 75.210 180.705 ;
        RECT 75.380 180.375 76.205 180.705 ;
        RECT 76.420 180.375 77.135 180.705 ;
        RECT 77.305 180.455 77.640 180.705 ;
        RECT 75.040 180.205 75.210 180.375 ;
        RECT 76.885 180.285 77.135 180.375 ;
        RECT 78.735 180.445 79.075 181.255 ;
        RECT 79.825 181.010 79.995 181.675 ;
        RECT 80.390 181.335 81.515 181.505 ;
        RECT 79.245 180.820 79.995 181.010 ;
        RECT 80.165 180.995 81.175 181.165 ;
        RECT 74.135 179.845 74.425 180.115 ;
        RECT 73.040 179.635 74.425 179.845 ;
        RECT 74.595 179.795 74.870 180.140 ;
        RECT 75.040 180.035 76.705 180.205 ;
        RECT 75.060 179.465 75.435 179.865 ;
        RECT 75.605 179.685 75.775 180.035 ;
        RECT 75.945 179.465 76.275 179.865 ;
        RECT 76.445 179.635 76.705 180.035 ;
        RECT 76.885 179.865 77.215 180.285 ;
        RECT 77.385 179.465 77.645 180.285 ;
        RECT 78.735 180.275 79.965 180.445 ;
        RECT 77.815 179.465 78.105 180.190 ;
        RECT 79.010 179.670 79.255 180.275 ;
        RECT 79.475 179.465 79.985 180.000 ;
        RECT 80.165 179.635 80.355 180.995 ;
        RECT 80.525 180.315 80.800 180.795 ;
        RECT 80.525 180.145 80.805 180.315 ;
        RECT 81.005 180.195 81.175 180.995 ;
        RECT 81.345 180.205 81.515 181.335 ;
        RECT 81.685 180.705 81.855 181.675 ;
        RECT 82.025 180.875 82.195 182.015 ;
        RECT 82.365 180.875 82.700 181.845 ;
        RECT 82.885 181.045 83.215 181.830 ;
        RECT 82.885 180.875 83.565 181.045 ;
        RECT 83.745 180.875 84.075 182.015 ;
        RECT 84.255 181.580 89.600 182.015 ;
        RECT 81.685 180.375 81.880 180.705 ;
        RECT 82.105 180.375 82.360 180.705 ;
        RECT 82.105 180.205 82.275 180.375 ;
        RECT 82.530 180.205 82.700 180.875 ;
        RECT 82.875 180.455 83.225 180.705 ;
        RECT 83.395 180.275 83.565 180.875 ;
        RECT 83.735 180.455 84.085 180.705 ;
        RECT 80.525 179.635 80.800 180.145 ;
        RECT 81.345 180.035 82.275 180.205 ;
        RECT 81.345 180.000 81.520 180.035 ;
        RECT 80.990 179.635 81.520 180.000 ;
        RECT 81.945 179.465 82.275 179.865 ;
        RECT 82.445 179.635 82.700 180.205 ;
        RECT 82.895 179.465 83.135 180.275 ;
        RECT 83.305 179.635 83.635 180.275 ;
        RECT 83.805 179.465 84.075 180.275 ;
        RECT 85.840 180.010 86.180 180.840 ;
        RECT 87.660 180.330 88.010 181.580 ;
        RECT 89.775 180.925 90.985 182.015 ;
        RECT 89.775 180.215 90.295 180.755 ;
        RECT 90.465 180.385 90.985 180.925 ;
        RECT 91.160 180.875 91.495 181.845 ;
        RECT 91.665 180.875 91.835 182.015 ;
        RECT 92.005 181.675 94.035 181.845 ;
        RECT 84.255 179.465 89.600 180.010 ;
        RECT 89.775 179.465 90.985 180.215 ;
        RECT 91.160 180.205 91.330 180.875 ;
        RECT 92.005 180.705 92.175 181.675 ;
        RECT 91.500 180.375 91.755 180.705 ;
        RECT 91.980 180.375 92.175 180.705 ;
        RECT 92.345 181.335 93.470 181.505 ;
        RECT 91.585 180.205 91.755 180.375 ;
        RECT 92.345 180.205 92.515 181.335 ;
        RECT 91.160 179.635 91.415 180.205 ;
        RECT 91.585 180.035 92.515 180.205 ;
        RECT 92.685 180.995 93.695 181.165 ;
        RECT 92.685 180.195 92.855 180.995 ;
        RECT 93.060 180.655 93.335 180.795 ;
        RECT 93.055 180.485 93.335 180.655 ;
        RECT 92.340 180.000 92.515 180.035 ;
        RECT 91.585 179.465 91.915 179.865 ;
        RECT 92.340 179.635 92.870 180.000 ;
        RECT 93.060 179.635 93.335 180.485 ;
        RECT 93.505 179.635 93.695 180.995 ;
        RECT 93.865 181.010 94.035 181.675 ;
        RECT 94.205 181.255 94.375 182.015 ;
        RECT 94.610 181.255 95.125 181.665 ;
        RECT 93.865 180.820 94.615 181.010 ;
        RECT 94.785 180.445 95.125 181.255 ;
        RECT 93.895 180.275 95.125 180.445 ;
        RECT 95.295 180.875 95.680 181.845 ;
        RECT 95.850 181.555 96.175 182.015 ;
        RECT 96.695 181.385 96.975 181.845 ;
        RECT 95.850 181.165 96.975 181.385 ;
        RECT 93.875 179.465 94.385 180.000 ;
        RECT 94.605 179.670 94.850 180.275 ;
        RECT 95.295 180.205 95.575 180.875 ;
        RECT 95.850 180.705 96.300 181.165 ;
        RECT 97.165 180.995 97.565 181.845 ;
        RECT 97.965 181.555 98.235 182.015 ;
        RECT 98.405 181.385 98.690 181.845 ;
        RECT 95.745 180.375 96.300 180.705 ;
        RECT 96.470 180.435 97.565 180.995 ;
        RECT 95.850 180.265 96.300 180.375 ;
        RECT 95.295 179.635 95.680 180.205 ;
        RECT 95.850 180.095 96.975 180.265 ;
        RECT 95.850 179.465 96.175 179.925 ;
        RECT 96.695 179.635 96.975 180.095 ;
        RECT 97.165 179.635 97.565 180.435 ;
        RECT 97.735 181.165 98.690 181.385 ;
        RECT 99.090 181.385 99.375 181.845 ;
        RECT 99.545 181.555 99.815 182.015 ;
        RECT 99.090 181.165 100.045 181.385 ;
        RECT 97.735 180.265 97.945 181.165 ;
        RECT 98.115 180.435 98.805 180.995 ;
        RECT 98.975 180.435 99.665 180.995 ;
        RECT 99.835 180.265 100.045 181.165 ;
        RECT 97.735 180.095 98.690 180.265 ;
        RECT 97.965 179.465 98.235 179.925 ;
        RECT 98.405 179.635 98.690 180.095 ;
        RECT 99.090 180.095 100.045 180.265 ;
        RECT 100.215 180.995 100.615 181.845 ;
        RECT 100.805 181.385 101.085 181.845 ;
        RECT 101.605 181.555 101.930 182.015 ;
        RECT 100.805 181.165 101.930 181.385 ;
        RECT 100.215 180.435 101.310 180.995 ;
        RECT 101.480 180.705 101.930 181.165 ;
        RECT 102.100 180.875 102.485 181.845 ;
        RECT 99.090 179.635 99.375 180.095 ;
        RECT 99.545 179.465 99.815 179.925 ;
        RECT 100.215 179.635 100.615 180.435 ;
        RECT 101.480 180.375 102.035 180.705 ;
        RECT 101.480 180.265 101.930 180.375 ;
        RECT 100.805 180.095 101.930 180.265 ;
        RECT 102.205 180.205 102.485 180.875 ;
        RECT 103.575 180.850 103.865 182.015 ;
        RECT 104.075 181.675 105.215 181.845 ;
        RECT 104.075 181.215 104.375 181.675 ;
        RECT 104.545 181.045 104.875 181.505 ;
        RECT 100.805 179.635 101.085 180.095 ;
        RECT 101.605 179.465 101.930 179.925 ;
        RECT 102.100 179.635 102.485 180.205 ;
        RECT 104.115 180.825 104.875 181.045 ;
        RECT 105.045 181.045 105.215 181.675 ;
        RECT 105.385 181.215 105.715 182.015 ;
        RECT 105.885 181.045 106.160 181.845 ;
        RECT 105.045 180.835 106.160 181.045 ;
        RECT 106.345 181.045 106.675 181.830 ;
        RECT 106.345 180.875 107.025 181.045 ;
        RECT 107.205 180.875 107.535 182.015 ;
        RECT 107.715 180.875 107.975 182.015 ;
        RECT 104.115 180.285 104.330 180.825 ;
        RECT 104.500 180.455 105.270 180.655 ;
        RECT 105.440 180.455 106.160 180.655 ;
        RECT 106.335 180.455 106.685 180.705 ;
        RECT 103.575 179.465 103.865 180.190 ;
        RECT 104.115 180.115 105.715 180.285 ;
        RECT 104.545 180.105 105.715 180.115 ;
        RECT 104.085 179.465 104.375 179.935 ;
        RECT 104.545 179.635 104.875 180.105 ;
        RECT 105.045 179.465 105.215 179.935 ;
        RECT 105.385 179.635 105.715 180.105 ;
        RECT 105.885 179.465 106.160 180.285 ;
        RECT 106.855 180.275 107.025 180.875 ;
        RECT 108.145 180.865 108.475 181.845 ;
        RECT 108.645 180.875 108.925 182.015 ;
        RECT 109.555 181.505 110.745 181.795 ;
        RECT 109.575 181.165 110.745 181.335 ;
        RECT 110.915 181.215 111.195 182.015 ;
        RECT 109.575 180.875 109.900 181.165 ;
        RECT 110.575 181.045 110.745 181.165 ;
        RECT 107.195 180.455 107.545 180.705 ;
        RECT 107.735 180.455 108.070 180.705 ;
        RECT 106.355 179.465 106.595 180.275 ;
        RECT 106.765 179.635 107.095 180.275 ;
        RECT 107.265 179.465 107.535 180.275 ;
        RECT 108.240 180.265 108.410 180.865 ;
        RECT 110.070 180.705 110.265 180.995 ;
        RECT 110.575 180.875 111.235 181.045 ;
        RECT 111.405 180.875 111.680 181.845 ;
        RECT 111.065 180.705 111.235 180.875 ;
        RECT 108.580 180.435 108.915 180.705 ;
        RECT 109.555 180.375 109.900 180.705 ;
        RECT 110.070 180.375 110.895 180.705 ;
        RECT 111.065 180.375 111.340 180.705 ;
        RECT 107.715 179.635 108.410 180.265 ;
        RECT 108.615 179.465 108.925 180.265 ;
        RECT 111.065 180.205 111.235 180.375 ;
        RECT 109.570 180.035 111.235 180.205 ;
        RECT 111.510 180.140 111.680 180.875 ;
        RECT 112.010 181.005 112.310 181.845 ;
        RECT 112.505 181.175 112.755 182.015 ;
        RECT 113.345 181.425 114.150 181.845 ;
        RECT 112.925 181.255 114.490 181.425 ;
        RECT 112.925 181.005 113.095 181.255 ;
        RECT 112.010 180.835 113.095 181.005 ;
        RECT 111.855 180.375 112.185 180.665 ;
        RECT 112.355 180.205 112.525 180.835 ;
        RECT 113.265 180.705 113.585 181.085 ;
        RECT 113.775 180.995 114.150 181.085 ;
        RECT 113.755 180.825 114.150 180.995 ;
        RECT 114.320 181.005 114.490 181.255 ;
        RECT 114.660 181.175 114.990 182.015 ;
        RECT 115.160 181.255 115.825 181.845 ;
        RECT 115.995 181.505 117.185 181.795 ;
        RECT 114.320 180.835 115.240 181.005 ;
        RECT 112.695 180.455 113.025 180.665 ;
        RECT 113.205 180.455 113.585 180.705 ;
        RECT 113.775 180.665 114.150 180.825 ;
        RECT 115.070 180.665 115.240 180.835 ;
        RECT 113.775 180.455 114.260 180.665 ;
        RECT 114.450 180.455 114.900 180.665 ;
        RECT 115.070 180.455 115.405 180.665 ;
        RECT 115.575 180.285 115.825 181.255 ;
        RECT 116.015 181.165 117.185 181.335 ;
        RECT 117.355 181.215 117.635 182.015 ;
        RECT 116.015 180.875 116.340 181.165 ;
        RECT 117.015 181.045 117.185 181.165 ;
        RECT 116.510 180.705 116.705 180.995 ;
        RECT 117.015 180.875 117.675 181.045 ;
        RECT 117.845 180.875 118.120 181.845 ;
        RECT 118.480 181.045 118.870 181.220 ;
        RECT 119.355 181.215 119.685 182.015 ;
        RECT 119.855 181.225 120.390 181.845 ;
        RECT 118.480 180.875 119.905 181.045 ;
        RECT 117.505 180.705 117.675 180.875 ;
        RECT 115.995 180.375 116.340 180.705 ;
        RECT 116.510 180.375 117.335 180.705 ;
        RECT 117.505 180.375 117.780 180.705 ;
        RECT 109.570 179.685 109.825 180.035 ;
        RECT 109.995 179.465 110.325 179.865 ;
        RECT 110.495 179.685 110.665 180.035 ;
        RECT 110.835 179.465 111.215 179.865 ;
        RECT 111.405 179.795 111.680 180.140 ;
        RECT 112.015 180.025 112.525 180.205 ;
        RECT 112.930 180.115 114.630 180.285 ;
        RECT 112.930 180.025 113.315 180.115 ;
        RECT 112.015 179.635 112.345 180.025 ;
        RECT 112.515 179.685 113.700 179.855 ;
        RECT 113.960 179.465 114.130 179.935 ;
        RECT 114.300 179.650 114.630 180.115 ;
        RECT 114.800 179.465 114.970 180.285 ;
        RECT 115.140 179.645 115.825 180.285 ;
        RECT 117.505 180.205 117.675 180.375 ;
        RECT 116.010 180.035 117.675 180.205 ;
        RECT 117.950 180.140 118.120 180.875 ;
        RECT 118.355 180.145 118.710 180.705 ;
        RECT 116.010 179.685 116.265 180.035 ;
        RECT 116.435 179.465 116.765 179.865 ;
        RECT 116.935 179.685 117.105 180.035 ;
        RECT 117.275 179.465 117.655 179.865 ;
        RECT 117.845 179.795 118.120 180.140 ;
        RECT 118.880 179.975 119.050 180.875 ;
        RECT 119.220 180.145 119.485 180.705 ;
        RECT 119.735 180.375 119.905 180.875 ;
        RECT 120.075 180.205 120.390 181.225 ;
        RECT 120.595 180.925 121.805 182.015 ;
        RECT 118.460 179.465 118.700 179.975 ;
        RECT 118.880 179.645 119.160 179.975 ;
        RECT 119.390 179.465 119.605 179.975 ;
        RECT 119.775 179.635 120.390 180.205 ;
        RECT 120.595 180.215 121.115 180.755 ;
        RECT 121.285 180.385 121.805 180.925 ;
        RECT 121.980 181.625 122.315 181.845 ;
        RECT 123.320 181.635 123.675 182.015 ;
        RECT 121.980 181.005 122.235 181.625 ;
        RECT 122.485 181.465 122.715 181.505 ;
        RECT 123.845 181.465 124.095 181.845 ;
        RECT 122.485 181.265 124.095 181.465 ;
        RECT 122.485 181.175 122.670 181.265 ;
        RECT 123.260 181.255 124.095 181.265 ;
        RECT 124.345 181.235 124.595 182.015 ;
        RECT 124.765 181.165 125.025 181.845 ;
        RECT 122.825 181.065 123.155 181.095 ;
        RECT 122.825 181.005 124.625 181.065 ;
        RECT 121.980 180.895 124.685 181.005 ;
        RECT 121.980 180.835 123.155 180.895 ;
        RECT 124.485 180.860 124.685 180.895 ;
        RECT 121.975 180.455 122.465 180.655 ;
        RECT 122.655 180.455 123.130 180.665 ;
        RECT 120.595 179.465 121.805 180.215 ;
        RECT 121.980 179.465 122.435 180.230 ;
        RECT 122.910 180.055 123.130 180.455 ;
        RECT 123.375 180.455 123.705 180.665 ;
        RECT 123.375 180.055 123.585 180.455 ;
        RECT 123.875 180.420 124.285 180.725 ;
        RECT 124.515 180.285 124.685 180.860 ;
        RECT 124.415 180.165 124.685 180.285 ;
        RECT 123.840 180.120 124.685 180.165 ;
        RECT 123.840 179.995 124.595 180.120 ;
        RECT 123.840 179.845 124.010 179.995 ;
        RECT 124.855 179.965 125.025 181.165 ;
        RECT 125.195 181.255 125.710 181.665 ;
        RECT 125.945 181.255 126.115 182.015 ;
        RECT 126.285 181.675 128.315 181.845 ;
        RECT 125.195 180.445 125.535 181.255 ;
        RECT 126.285 181.010 126.455 181.675 ;
        RECT 126.850 181.335 127.975 181.505 ;
        RECT 125.705 180.820 126.455 181.010 ;
        RECT 126.625 180.995 127.635 181.165 ;
        RECT 125.195 180.275 126.425 180.445 ;
        RECT 122.710 179.635 124.010 179.845 ;
        RECT 124.265 179.465 124.595 179.825 ;
        RECT 124.765 179.635 125.025 179.965 ;
        RECT 125.470 179.670 125.715 180.275 ;
        RECT 125.935 179.465 126.445 180.000 ;
        RECT 126.625 179.635 126.815 180.995 ;
        RECT 126.985 180.655 127.260 180.795 ;
        RECT 126.985 180.485 127.265 180.655 ;
        RECT 126.985 179.635 127.260 180.485 ;
        RECT 127.465 180.195 127.635 180.995 ;
        RECT 127.805 180.205 127.975 181.335 ;
        RECT 128.145 180.705 128.315 181.675 ;
        RECT 128.485 180.875 128.655 182.015 ;
        RECT 128.825 180.875 129.160 181.845 ;
        RECT 128.145 180.375 128.340 180.705 ;
        RECT 128.565 180.375 128.820 180.705 ;
        RECT 128.565 180.205 128.735 180.375 ;
        RECT 128.990 180.205 129.160 180.875 ;
        RECT 129.335 180.850 129.625 182.015 ;
        RECT 129.885 181.345 130.055 181.845 ;
        RECT 130.225 181.515 130.555 182.015 ;
        RECT 129.885 181.175 130.550 181.345 ;
        RECT 129.800 180.355 130.150 181.005 ;
        RECT 127.805 180.035 128.735 180.205 ;
        RECT 127.805 180.000 127.980 180.035 ;
        RECT 127.450 179.635 127.980 180.000 ;
        RECT 128.405 179.465 128.735 179.865 ;
        RECT 128.905 179.635 129.160 180.205 ;
        RECT 129.335 179.465 129.625 180.190 ;
        RECT 130.320 180.185 130.550 181.175 ;
        RECT 129.885 180.015 130.550 180.185 ;
        RECT 129.885 179.725 130.055 180.015 ;
        RECT 130.225 179.465 130.555 179.845 ;
        RECT 130.725 179.725 130.910 181.845 ;
        RECT 131.150 181.555 131.415 182.015 ;
        RECT 131.585 181.420 131.835 181.845 ;
        RECT 132.045 181.570 133.150 181.740 ;
        RECT 131.530 181.290 131.835 181.420 ;
        RECT 131.080 180.095 131.360 181.045 ;
        RECT 131.530 180.185 131.700 181.290 ;
        RECT 131.870 180.505 132.110 181.100 ;
        RECT 132.280 181.035 132.810 181.400 ;
        RECT 132.280 180.335 132.450 181.035 ;
        RECT 132.980 180.955 133.150 181.570 ;
        RECT 133.320 181.215 133.490 182.015 ;
        RECT 133.660 181.515 133.910 181.845 ;
        RECT 134.135 181.545 135.020 181.715 ;
        RECT 132.980 180.865 133.490 180.955 ;
        RECT 131.530 180.055 131.755 180.185 ;
        RECT 131.925 180.115 132.450 180.335 ;
        RECT 132.620 180.695 133.490 180.865 ;
        RECT 131.165 179.465 131.415 179.925 ;
        RECT 131.585 179.915 131.755 180.055 ;
        RECT 132.620 179.915 132.790 180.695 ;
        RECT 133.320 180.625 133.490 180.695 ;
        RECT 133.000 180.445 133.200 180.475 ;
        RECT 133.660 180.445 133.830 181.515 ;
        RECT 134.000 180.625 134.190 181.345 ;
        RECT 133.000 180.145 133.830 180.445 ;
        RECT 134.360 180.415 134.680 181.375 ;
        RECT 131.585 179.745 131.920 179.915 ;
        RECT 132.115 179.745 132.790 179.915 ;
        RECT 133.110 179.465 133.480 179.965 ;
        RECT 133.660 179.915 133.830 180.145 ;
        RECT 134.215 180.085 134.680 180.415 ;
        RECT 134.850 180.705 135.020 181.545 ;
        RECT 135.200 181.515 135.515 182.015 ;
        RECT 135.745 181.285 136.085 181.845 ;
        RECT 135.190 180.910 136.085 181.285 ;
        RECT 136.255 181.005 136.425 182.015 ;
        RECT 135.895 180.705 136.085 180.910 ;
        RECT 136.595 180.955 136.925 181.800 ;
        RECT 136.595 180.875 136.985 180.955 ;
        RECT 136.770 180.825 136.985 180.875 ;
        RECT 134.850 180.375 135.725 180.705 ;
        RECT 135.895 180.375 136.645 180.705 ;
        RECT 134.850 179.915 135.020 180.375 ;
        RECT 135.895 180.205 136.095 180.375 ;
        RECT 136.815 180.245 136.985 180.825 ;
        RECT 137.615 180.925 138.825 182.015 ;
        RECT 137.615 180.385 138.135 180.925 ;
        RECT 136.760 180.205 136.985 180.245 ;
        RECT 138.305 180.215 138.825 180.755 ;
        RECT 133.660 179.745 134.065 179.915 ;
        RECT 134.235 179.745 135.020 179.915 ;
        RECT 135.295 179.465 135.505 179.995 ;
        RECT 135.765 179.680 136.095 180.205 ;
        RECT 136.605 180.120 136.985 180.205 ;
        RECT 136.265 179.465 136.435 180.075 ;
        RECT 136.605 179.685 136.935 180.120 ;
        RECT 137.615 179.465 138.825 180.215 ;
        RECT 13.330 179.295 138.910 179.465 ;
        RECT 13.415 178.545 14.625 179.295 ;
        RECT 13.415 178.005 13.935 178.545 ;
        RECT 14.795 178.525 16.465 179.295 ;
        RECT 14.105 177.835 14.625 178.375 ;
        RECT 14.795 178.005 15.545 178.525 ;
        RECT 16.645 178.485 16.915 179.295 ;
        RECT 17.085 178.485 17.415 179.125 ;
        RECT 17.585 178.485 17.825 179.295 ;
        RECT 18.020 179.040 18.355 179.085 ;
        RECT 18.015 178.575 18.355 179.040 ;
        RECT 18.525 178.915 18.855 179.295 ;
        RECT 19.315 178.955 19.585 178.960 ;
        RECT 19.315 178.785 19.625 178.955 ;
        RECT 15.715 177.835 16.465 178.355 ;
        RECT 16.635 178.055 16.985 178.305 ;
        RECT 17.155 177.885 17.325 178.485 ;
        RECT 17.495 178.055 17.845 178.305 ;
        RECT 18.015 177.885 18.185 178.575 ;
        RECT 18.355 178.055 18.615 178.385 ;
        RECT 13.415 176.745 14.625 177.835 ;
        RECT 14.795 176.745 16.465 177.835 ;
        RECT 16.645 176.745 16.975 177.885 ;
        RECT 17.155 177.715 17.835 177.885 ;
        RECT 17.505 176.930 17.835 177.715 ;
        RECT 18.015 176.915 18.275 177.885 ;
        RECT 18.445 177.505 18.615 178.055 ;
        RECT 18.785 177.685 19.125 178.715 ;
        RECT 19.315 177.685 19.585 178.785 ;
        RECT 19.810 177.685 20.090 178.960 ;
        RECT 20.290 178.795 20.520 179.125 ;
        RECT 20.765 178.915 21.095 179.295 ;
        RECT 20.290 177.505 20.460 178.795 ;
        RECT 21.265 178.725 21.440 179.125 ;
        RECT 20.810 178.555 21.440 178.725 ;
        RECT 21.695 178.645 21.955 179.125 ;
        RECT 22.125 178.755 22.375 179.295 ;
        RECT 20.810 178.385 20.980 178.555 ;
        RECT 20.630 178.055 20.980 178.385 ;
        RECT 18.445 177.335 20.460 177.505 ;
        RECT 20.810 177.535 20.980 178.055 ;
        RECT 21.160 177.705 21.525 178.385 ;
        RECT 21.695 177.615 21.865 178.645 ;
        RECT 22.545 178.615 22.765 179.075 ;
        RECT 22.515 178.590 22.765 178.615 ;
        RECT 22.035 177.995 22.265 178.390 ;
        RECT 22.435 178.165 22.765 178.590 ;
        RECT 22.935 178.915 23.825 179.085 ;
        RECT 22.935 178.190 23.105 178.915 ;
        RECT 24.080 178.795 24.575 179.125 ;
        RECT 23.275 178.360 23.825 178.745 ;
        RECT 22.935 178.120 23.825 178.190 ;
        RECT 22.930 178.095 23.825 178.120 ;
        RECT 22.920 178.080 23.825 178.095 ;
        RECT 22.915 178.065 23.825 178.080 ;
        RECT 22.905 178.060 23.825 178.065 ;
        RECT 22.900 178.050 23.825 178.060 ;
        RECT 22.895 178.040 23.825 178.050 ;
        RECT 22.885 178.035 23.825 178.040 ;
        RECT 22.875 178.025 23.825 178.035 ;
        RECT 22.865 178.020 23.825 178.025 ;
        RECT 22.865 178.015 23.200 178.020 ;
        RECT 22.850 178.010 23.200 178.015 ;
        RECT 22.835 178.000 23.200 178.010 ;
        RECT 22.810 177.995 23.200 178.000 ;
        RECT 22.035 177.990 23.200 177.995 ;
        RECT 22.035 177.955 23.170 177.990 ;
        RECT 22.035 177.930 23.135 177.955 ;
        RECT 22.035 177.900 23.105 177.930 ;
        RECT 22.035 177.870 23.085 177.900 ;
        RECT 22.035 177.840 23.065 177.870 ;
        RECT 22.035 177.830 22.995 177.840 ;
        RECT 22.035 177.820 22.970 177.830 ;
        RECT 22.035 177.805 22.950 177.820 ;
        RECT 22.035 177.790 22.930 177.805 ;
        RECT 22.140 177.780 22.925 177.790 ;
        RECT 22.140 177.745 22.910 177.780 ;
        RECT 20.810 177.365 21.440 177.535 ;
        RECT 18.470 176.745 18.800 177.155 ;
        RECT 19.000 176.915 19.170 177.335 ;
        RECT 19.385 176.745 20.055 177.155 ;
        RECT 20.290 176.915 20.460 177.335 ;
        RECT 20.765 176.745 21.095 177.185 ;
        RECT 21.265 176.915 21.440 177.365 ;
        RECT 21.695 176.915 21.970 177.615 ;
        RECT 22.140 177.495 22.895 177.745 ;
        RECT 23.065 177.425 23.395 177.670 ;
        RECT 23.565 177.570 23.825 178.020 ;
        RECT 23.210 177.400 23.395 177.425 ;
        RECT 23.210 177.300 23.825 177.400 ;
        RECT 23.995 177.305 24.235 178.615 ;
        RECT 24.405 177.885 24.575 178.795 ;
        RECT 24.795 178.055 25.145 179.020 ;
        RECT 25.325 178.055 25.625 179.025 ;
        RECT 25.805 178.055 26.085 179.025 ;
        RECT 26.265 178.495 26.535 179.295 ;
        RECT 26.705 178.575 27.045 179.085 ;
        RECT 26.280 178.055 26.610 178.305 ;
        RECT 26.280 177.885 26.595 178.055 ;
        RECT 24.405 177.715 26.595 177.885 ;
        RECT 22.140 176.745 22.395 177.290 ;
        RECT 22.565 176.915 23.045 177.255 ;
        RECT 23.220 176.745 23.825 177.300 ;
        RECT 24.000 176.745 24.335 177.125 ;
        RECT 24.505 176.915 24.755 177.715 ;
        RECT 24.975 176.745 25.305 177.465 ;
        RECT 25.490 176.915 25.740 177.715 ;
        RECT 26.205 176.745 26.535 177.545 ;
        RECT 26.785 177.175 27.045 178.575 ;
        RECT 27.215 178.525 29.805 179.295 ;
        RECT 27.215 178.005 28.425 178.525 ;
        RECT 30.180 178.515 30.680 179.125 ;
        RECT 28.595 177.835 29.805 178.355 ;
        RECT 29.975 178.055 30.325 178.305 ;
        RECT 30.510 177.885 30.680 178.515 ;
        RECT 31.310 178.645 31.640 179.125 ;
        RECT 31.810 178.835 32.035 179.295 ;
        RECT 32.205 178.645 32.535 179.125 ;
        RECT 31.310 178.475 32.535 178.645 ;
        RECT 32.725 178.495 32.975 179.295 ;
        RECT 33.145 178.495 33.485 179.125 ;
        RECT 34.360 178.815 34.660 179.295 ;
        RECT 34.830 178.645 35.090 179.100 ;
        RECT 35.260 178.815 35.520 179.295 ;
        RECT 35.690 178.645 35.950 179.100 ;
        RECT 36.120 178.815 36.380 179.295 ;
        RECT 36.550 178.645 36.810 179.100 ;
        RECT 36.980 178.815 37.240 179.295 ;
        RECT 37.410 178.645 37.670 179.100 ;
        RECT 37.840 178.770 38.100 179.295 ;
        RECT 30.850 178.105 31.180 178.305 ;
        RECT 31.350 178.105 31.680 178.305 ;
        RECT 31.850 178.105 32.270 178.305 ;
        RECT 32.445 178.135 33.140 178.305 ;
        RECT 32.445 177.885 32.615 178.135 ;
        RECT 33.310 177.885 33.485 178.495 ;
        RECT 26.705 176.915 27.045 177.175 ;
        RECT 27.215 176.745 29.805 177.835 ;
        RECT 30.180 177.715 32.615 177.885 ;
        RECT 30.180 176.915 30.510 177.715 ;
        RECT 30.680 176.745 31.010 177.545 ;
        RECT 31.310 176.915 31.640 177.715 ;
        RECT 32.285 176.745 32.535 177.545 ;
        RECT 32.805 176.745 32.975 177.885 ;
        RECT 33.145 176.915 33.485 177.885 ;
        RECT 34.360 178.475 37.670 178.645 ;
        RECT 34.360 177.885 35.330 178.475 ;
        RECT 38.270 178.305 38.520 179.115 ;
        RECT 38.700 178.835 38.945 179.295 ;
        RECT 35.500 178.055 38.520 178.305 ;
        RECT 38.690 178.055 39.005 178.665 ;
        RECT 39.175 178.570 39.465 179.295 ;
        RECT 39.645 178.645 39.975 179.120 ;
        RECT 40.145 178.815 40.315 179.295 ;
        RECT 40.485 178.645 40.815 179.120 ;
        RECT 40.985 178.815 41.155 179.295 ;
        RECT 41.325 178.645 41.655 179.120 ;
        RECT 41.825 178.815 41.995 179.295 ;
        RECT 42.165 178.645 42.495 179.120 ;
        RECT 42.665 178.815 42.835 179.295 ;
        RECT 43.005 178.645 43.335 179.120 ;
        RECT 43.505 178.815 43.675 179.295 ;
        RECT 43.845 179.120 44.095 179.125 ;
        RECT 43.845 178.645 44.175 179.120 ;
        RECT 44.345 178.815 44.515 179.295 ;
        RECT 44.765 179.120 44.935 179.125 ;
        RECT 44.685 178.645 45.015 179.120 ;
        RECT 45.185 178.815 45.355 179.295 ;
        RECT 45.605 179.120 45.775 179.125 ;
        RECT 45.525 178.645 45.855 179.120 ;
        RECT 46.025 178.815 46.195 179.295 ;
        RECT 46.365 178.645 46.695 179.120 ;
        RECT 46.865 178.815 47.035 179.295 ;
        RECT 47.205 178.645 47.535 179.120 ;
        RECT 47.705 178.815 47.875 179.295 ;
        RECT 48.045 178.645 48.375 179.120 ;
        RECT 48.545 178.815 48.715 179.295 ;
        RECT 48.885 178.645 49.215 179.120 ;
        RECT 49.385 178.815 49.555 179.295 ;
        RECT 49.725 178.645 50.055 179.120 ;
        RECT 50.225 178.815 50.395 179.295 ;
        RECT 50.920 178.815 51.220 179.295 ;
        RECT 51.390 178.645 51.650 179.100 ;
        RECT 51.820 178.815 52.080 179.295 ;
        RECT 52.250 178.645 52.510 179.100 ;
        RECT 52.680 178.815 52.940 179.295 ;
        RECT 53.110 178.645 53.370 179.100 ;
        RECT 53.540 178.815 53.800 179.295 ;
        RECT 53.970 178.645 54.230 179.100 ;
        RECT 54.400 178.770 54.660 179.295 ;
        RECT 39.645 178.475 41.155 178.645 ;
        RECT 41.325 178.475 43.675 178.645 ;
        RECT 43.845 178.475 50.505 178.645 ;
        RECT 40.985 178.305 41.155 178.475 ;
        RECT 43.500 178.305 43.675 178.475 ;
        RECT 39.640 178.105 40.815 178.305 ;
        RECT 40.985 178.105 43.295 178.305 ;
        RECT 43.500 178.105 50.060 178.305 ;
        RECT 34.360 177.645 37.670 177.885 ;
        RECT 34.365 176.745 34.660 177.475 ;
        RECT 34.830 176.920 35.090 177.645 ;
        RECT 35.260 176.745 35.520 177.475 ;
        RECT 35.690 176.920 35.950 177.645 ;
        RECT 36.120 176.745 36.380 177.475 ;
        RECT 36.550 176.920 36.810 177.645 ;
        RECT 36.980 176.745 37.240 177.475 ;
        RECT 37.410 176.920 37.670 177.645 ;
        RECT 37.840 176.745 38.100 177.855 ;
        RECT 38.270 176.920 38.520 178.055 ;
        RECT 40.985 177.935 41.155 178.105 ;
        RECT 43.500 177.935 43.675 178.105 ;
        RECT 50.230 177.935 50.505 178.475 ;
        RECT 38.700 176.745 38.995 177.855 ;
        RECT 39.175 176.745 39.465 177.910 ;
        RECT 39.645 177.765 41.155 177.935 ;
        RECT 41.325 177.765 43.675 177.935 ;
        RECT 43.845 177.765 50.505 177.935 ;
        RECT 50.920 178.475 54.230 178.645 ;
        RECT 50.920 177.885 51.890 178.475 ;
        RECT 54.830 178.305 55.080 179.115 ;
        RECT 55.260 178.835 55.505 179.295 ;
        RECT 52.060 178.055 55.080 178.305 ;
        RECT 55.250 178.055 55.565 178.665 ;
        RECT 55.755 178.485 55.995 179.295 ;
        RECT 56.165 178.485 56.495 179.125 ;
        RECT 56.665 178.485 56.935 179.295 ;
        RECT 57.115 178.750 62.460 179.295 ;
        RECT 55.735 178.055 56.085 178.305 ;
        RECT 39.645 176.915 39.975 177.765 ;
        RECT 40.145 176.745 40.315 177.595 ;
        RECT 40.485 176.915 40.815 177.765 ;
        RECT 40.985 176.745 41.155 177.595 ;
        RECT 41.325 176.915 41.655 177.765 ;
        RECT 41.825 176.745 41.995 177.545 ;
        RECT 42.165 176.915 42.495 177.765 ;
        RECT 42.665 176.745 42.835 177.545 ;
        RECT 43.005 176.915 43.335 177.765 ;
        RECT 43.505 176.745 43.675 177.545 ;
        RECT 43.845 176.915 44.175 177.765 ;
        RECT 44.345 176.745 44.515 177.545 ;
        RECT 44.685 176.915 45.015 177.765 ;
        RECT 45.185 176.745 45.355 177.545 ;
        RECT 45.525 176.915 45.855 177.765 ;
        RECT 46.025 176.745 46.195 177.545 ;
        RECT 46.365 176.915 46.695 177.765 ;
        RECT 46.865 176.745 47.035 177.545 ;
        RECT 47.205 176.915 47.535 177.765 ;
        RECT 47.705 176.745 47.875 177.545 ;
        RECT 48.045 176.915 48.375 177.765 ;
        RECT 48.545 176.745 48.715 177.545 ;
        RECT 48.885 176.915 49.215 177.765 ;
        RECT 49.385 176.745 49.555 177.545 ;
        RECT 49.725 176.915 50.055 177.765 ;
        RECT 50.920 177.645 54.230 177.885 ;
        RECT 50.225 176.745 50.395 177.545 ;
        RECT 50.925 176.745 51.220 177.475 ;
        RECT 51.390 176.920 51.650 177.645 ;
        RECT 51.820 176.745 52.080 177.475 ;
        RECT 52.250 176.920 52.510 177.645 ;
        RECT 52.680 176.745 52.940 177.475 ;
        RECT 53.110 176.920 53.370 177.645 ;
        RECT 53.540 176.745 53.800 177.475 ;
        RECT 53.970 176.920 54.230 177.645 ;
        RECT 54.400 176.745 54.660 177.855 ;
        RECT 54.830 176.920 55.080 178.055 ;
        RECT 56.255 177.885 56.425 178.485 ;
        RECT 56.595 178.055 56.945 178.305 ;
        RECT 58.700 177.920 59.040 178.750 ;
        RECT 62.635 178.525 64.305 179.295 ;
        RECT 64.935 178.570 65.225 179.295 ;
        RECT 65.445 178.640 65.775 179.075 ;
        RECT 65.945 178.685 66.115 179.295 ;
        RECT 65.395 178.555 65.775 178.640 ;
        RECT 66.285 178.555 66.615 179.080 ;
        RECT 66.875 178.765 67.085 179.295 ;
        RECT 67.360 178.845 68.145 179.015 ;
        RECT 68.315 178.845 68.720 179.015 ;
        RECT 55.260 176.745 55.555 177.855 ;
        RECT 55.745 177.715 56.425 177.885 ;
        RECT 55.745 176.930 56.075 177.715 ;
        RECT 56.605 176.745 56.935 177.885 ;
        RECT 60.520 177.180 60.870 178.430 ;
        RECT 62.635 178.005 63.385 178.525 ;
        RECT 65.395 178.515 65.620 178.555 ;
        RECT 63.555 177.835 64.305 178.355 ;
        RECT 65.395 177.935 65.565 178.515 ;
        RECT 66.285 178.385 66.485 178.555 ;
        RECT 67.360 178.385 67.530 178.845 ;
        RECT 65.735 178.055 66.485 178.385 ;
        RECT 66.655 178.055 67.530 178.385 ;
        RECT 57.115 176.745 62.460 177.180 ;
        RECT 62.635 176.745 64.305 177.835 ;
        RECT 64.935 176.745 65.225 177.910 ;
        RECT 65.395 177.885 65.610 177.935 ;
        RECT 65.395 177.805 65.785 177.885 ;
        RECT 65.455 176.960 65.785 177.805 ;
        RECT 66.295 177.850 66.485 178.055 ;
        RECT 65.955 176.745 66.125 177.755 ;
        RECT 66.295 177.475 67.190 177.850 ;
        RECT 66.295 176.915 66.635 177.475 ;
        RECT 66.865 176.745 67.180 177.245 ;
        RECT 67.360 177.215 67.530 178.055 ;
        RECT 67.700 178.345 68.165 178.675 ;
        RECT 68.550 178.615 68.720 178.845 ;
        RECT 68.900 178.795 69.270 179.295 ;
        RECT 69.590 178.845 70.265 179.015 ;
        RECT 70.460 178.845 70.795 179.015 ;
        RECT 67.700 177.385 68.020 178.345 ;
        RECT 68.550 178.315 69.380 178.615 ;
        RECT 68.190 177.415 68.380 178.135 ;
        RECT 68.550 177.245 68.720 178.315 ;
        RECT 69.180 178.285 69.380 178.315 ;
        RECT 68.890 178.065 69.060 178.135 ;
        RECT 69.590 178.065 69.760 178.845 ;
        RECT 70.625 178.705 70.795 178.845 ;
        RECT 70.965 178.835 71.215 179.295 ;
        RECT 68.890 177.895 69.760 178.065 ;
        RECT 69.930 178.425 70.455 178.645 ;
        RECT 70.625 178.575 70.850 178.705 ;
        RECT 68.890 177.805 69.400 177.895 ;
        RECT 67.360 177.045 68.245 177.215 ;
        RECT 68.470 176.915 68.720 177.245 ;
        RECT 68.890 176.745 69.060 177.545 ;
        RECT 69.230 177.190 69.400 177.805 ;
        RECT 69.930 177.725 70.100 178.425 ;
        RECT 69.570 177.360 70.100 177.725 ;
        RECT 70.270 177.660 70.510 178.255 ;
        RECT 70.680 177.470 70.850 178.575 ;
        RECT 71.020 177.715 71.300 178.665 ;
        RECT 70.545 177.340 70.850 177.470 ;
        RECT 69.230 177.020 70.335 177.190 ;
        RECT 70.545 176.915 70.795 177.340 ;
        RECT 70.965 176.745 71.230 177.205 ;
        RECT 71.470 176.915 71.655 179.035 ;
        RECT 71.825 178.915 72.155 179.295 ;
        RECT 72.325 178.745 72.495 179.035 ;
        RECT 71.830 178.575 72.495 178.745 ;
        RECT 71.830 177.585 72.060 178.575 ;
        RECT 72.230 177.755 72.580 178.405 ;
        RECT 71.830 177.415 72.495 177.585 ;
        RECT 71.825 176.745 72.155 177.245 ;
        RECT 72.325 176.915 72.495 177.415 ;
        RECT 72.765 176.925 73.025 179.115 ;
        RECT 73.285 178.925 73.955 179.295 ;
        RECT 74.135 178.745 74.445 179.115 ;
        RECT 73.215 178.545 74.445 178.745 ;
        RECT 73.215 177.875 73.505 178.545 ;
        RECT 74.625 178.365 74.855 179.005 ;
        RECT 75.035 178.565 75.325 179.295 ;
        RECT 75.550 178.555 76.165 179.125 ;
        RECT 76.335 178.785 76.550 179.295 ;
        RECT 76.780 178.785 77.060 179.115 ;
        RECT 77.240 178.785 77.480 179.295 ;
        RECT 77.815 178.835 78.375 179.125 ;
        RECT 78.545 178.835 78.795 179.295 ;
        RECT 73.685 178.055 74.150 178.365 ;
        RECT 74.330 178.055 74.855 178.365 ;
        RECT 75.035 178.055 75.335 178.385 ;
        RECT 73.215 177.655 73.985 177.875 ;
        RECT 73.195 176.745 73.535 177.475 ;
        RECT 73.715 176.925 73.985 177.655 ;
        RECT 74.165 177.635 75.325 177.875 ;
        RECT 74.165 176.925 74.395 177.635 ;
        RECT 74.565 176.745 74.895 177.455 ;
        RECT 75.065 176.925 75.325 177.635 ;
        RECT 75.550 177.535 75.865 178.555 ;
        RECT 76.035 177.885 76.205 178.385 ;
        RECT 76.455 178.055 76.720 178.615 ;
        RECT 76.890 177.885 77.060 178.785 ;
        RECT 77.230 178.055 77.585 178.615 ;
        RECT 76.035 177.715 77.460 177.885 ;
        RECT 75.550 176.915 76.085 177.535 ;
        RECT 76.255 176.745 76.585 177.545 ;
        RECT 77.070 177.540 77.460 177.715 ;
        RECT 77.815 177.465 78.065 178.835 ;
        RECT 79.415 178.665 79.745 179.025 ;
        RECT 78.355 178.475 79.745 178.665 ;
        RECT 80.230 178.665 80.515 179.125 ;
        RECT 80.685 178.835 80.955 179.295 ;
        RECT 80.230 178.495 81.185 178.665 ;
        RECT 78.355 178.385 78.525 178.475 ;
        RECT 78.235 178.055 78.525 178.385 ;
        RECT 78.695 178.055 79.035 178.305 ;
        RECT 79.255 178.055 79.930 178.305 ;
        RECT 78.355 177.805 78.525 178.055 ;
        RECT 78.355 177.635 79.295 177.805 ;
        RECT 79.665 177.695 79.930 178.055 ;
        RECT 80.115 177.765 80.805 178.325 ;
        RECT 77.815 176.915 78.275 177.465 ;
        RECT 78.465 176.745 78.795 177.465 ;
        RECT 78.995 177.085 79.295 177.635 ;
        RECT 80.975 177.595 81.185 178.495 ;
        RECT 79.465 176.745 79.745 177.415 ;
        RECT 80.230 177.375 81.185 177.595 ;
        RECT 81.355 178.325 81.755 179.125 ;
        RECT 81.945 178.665 82.225 179.125 ;
        RECT 82.745 178.835 83.070 179.295 ;
        RECT 81.945 178.495 83.070 178.665 ;
        RECT 83.240 178.555 83.625 179.125 ;
        RECT 82.620 178.385 83.070 178.495 ;
        RECT 81.355 177.765 82.450 178.325 ;
        RECT 82.620 178.055 83.175 178.385 ;
        RECT 80.230 176.915 80.515 177.375 ;
        RECT 80.685 176.745 80.955 177.205 ;
        RECT 81.355 176.915 81.755 177.765 ;
        RECT 82.620 177.595 83.070 178.055 ;
        RECT 83.345 177.885 83.625 178.555 ;
        RECT 81.945 177.375 83.070 177.595 ;
        RECT 81.945 176.915 82.225 177.375 ;
        RECT 82.745 176.745 83.070 177.205 ;
        RECT 83.240 176.915 83.625 177.885 ;
        RECT 83.800 178.555 84.055 179.125 ;
        RECT 84.225 178.895 84.555 179.295 ;
        RECT 84.980 178.760 85.510 179.125 ;
        RECT 84.980 178.725 85.155 178.760 ;
        RECT 84.225 178.555 85.155 178.725 ;
        RECT 83.800 177.885 83.970 178.555 ;
        RECT 84.225 178.385 84.395 178.555 ;
        RECT 84.140 178.055 84.395 178.385 ;
        RECT 84.620 178.055 84.815 178.385 ;
        RECT 83.800 176.915 84.135 177.885 ;
        RECT 84.305 176.745 84.475 177.885 ;
        RECT 84.645 177.085 84.815 178.055 ;
        RECT 84.985 177.425 85.155 178.555 ;
        RECT 85.325 177.765 85.495 178.565 ;
        RECT 85.700 178.275 85.975 179.125 ;
        RECT 85.695 178.105 85.975 178.275 ;
        RECT 85.700 177.965 85.975 178.105 ;
        RECT 86.145 177.765 86.335 179.125 ;
        RECT 86.515 178.760 87.025 179.295 ;
        RECT 87.245 178.485 87.490 179.090 ;
        RECT 87.935 178.525 90.525 179.295 ;
        RECT 90.695 178.570 90.985 179.295 ;
        RECT 91.205 178.640 91.535 179.075 ;
        RECT 91.705 178.685 91.875 179.295 ;
        RECT 91.155 178.555 91.535 178.640 ;
        RECT 92.045 178.555 92.375 179.080 ;
        RECT 92.635 178.765 92.845 179.295 ;
        RECT 93.120 178.845 93.905 179.015 ;
        RECT 94.075 178.845 94.480 179.015 ;
        RECT 86.535 178.315 87.765 178.485 ;
        RECT 85.325 177.595 86.335 177.765 ;
        RECT 86.505 177.750 87.255 177.940 ;
        RECT 84.985 177.255 86.110 177.425 ;
        RECT 86.505 177.085 86.675 177.750 ;
        RECT 87.425 177.505 87.765 178.315 ;
        RECT 87.935 178.005 89.145 178.525 ;
        RECT 91.155 178.515 91.380 178.555 ;
        RECT 89.315 177.835 90.525 178.355 ;
        RECT 91.155 177.935 91.325 178.515 ;
        RECT 92.045 178.385 92.245 178.555 ;
        RECT 93.120 178.385 93.290 178.845 ;
        RECT 91.495 178.055 92.245 178.385 ;
        RECT 92.415 178.055 93.290 178.385 ;
        RECT 84.645 176.915 86.675 177.085 ;
        RECT 86.845 176.745 87.015 177.505 ;
        RECT 87.250 177.095 87.765 177.505 ;
        RECT 87.935 176.745 90.525 177.835 ;
        RECT 90.695 176.745 90.985 177.910 ;
        RECT 91.155 177.885 91.370 177.935 ;
        RECT 91.155 177.805 91.545 177.885 ;
        RECT 91.215 176.960 91.545 177.805 ;
        RECT 92.055 177.850 92.245 178.055 ;
        RECT 91.715 176.745 91.885 177.755 ;
        RECT 92.055 177.475 92.950 177.850 ;
        RECT 92.055 176.915 92.395 177.475 ;
        RECT 92.625 176.745 92.940 177.245 ;
        RECT 93.120 177.215 93.290 178.055 ;
        RECT 93.460 178.345 93.925 178.675 ;
        RECT 94.310 178.615 94.480 178.845 ;
        RECT 94.660 178.795 95.030 179.295 ;
        RECT 95.350 178.845 96.025 179.015 ;
        RECT 96.220 178.845 96.555 179.015 ;
        RECT 93.460 177.385 93.780 178.345 ;
        RECT 94.310 178.315 95.140 178.615 ;
        RECT 93.950 177.415 94.140 178.135 ;
        RECT 94.310 177.245 94.480 178.315 ;
        RECT 94.940 178.285 95.140 178.315 ;
        RECT 94.650 178.065 94.820 178.135 ;
        RECT 95.350 178.065 95.520 178.845 ;
        RECT 96.385 178.705 96.555 178.845 ;
        RECT 96.725 178.835 96.975 179.295 ;
        RECT 94.650 177.895 95.520 178.065 ;
        RECT 95.690 178.425 96.215 178.645 ;
        RECT 96.385 178.575 96.610 178.705 ;
        RECT 94.650 177.805 95.160 177.895 ;
        RECT 93.120 177.045 94.005 177.215 ;
        RECT 94.230 176.915 94.480 177.245 ;
        RECT 94.650 176.745 94.820 177.545 ;
        RECT 94.990 177.190 95.160 177.805 ;
        RECT 95.690 177.725 95.860 178.425 ;
        RECT 95.330 177.360 95.860 177.725 ;
        RECT 96.030 177.660 96.270 178.255 ;
        RECT 96.440 177.470 96.610 178.575 ;
        RECT 96.780 177.715 97.060 178.665 ;
        RECT 96.305 177.340 96.610 177.470 ;
        RECT 94.990 177.020 96.095 177.190 ;
        RECT 96.305 176.915 96.555 177.340 ;
        RECT 96.725 176.745 96.990 177.205 ;
        RECT 97.230 176.915 97.415 179.035 ;
        RECT 97.585 178.915 97.915 179.295 ;
        RECT 98.085 178.745 98.255 179.035 ;
        RECT 97.590 178.575 98.255 178.745 ;
        RECT 98.515 178.795 98.775 179.125 ;
        RECT 98.945 178.935 99.275 179.295 ;
        RECT 99.530 178.915 100.830 179.125 ;
        RECT 98.515 178.785 98.745 178.795 ;
        RECT 97.590 177.585 97.820 178.575 ;
        RECT 97.990 177.755 98.340 178.405 ;
        RECT 98.515 177.595 98.685 178.785 ;
        RECT 99.530 178.765 99.700 178.915 ;
        RECT 98.945 178.640 99.700 178.765 ;
        RECT 98.855 178.595 99.700 178.640 ;
        RECT 98.855 178.475 99.125 178.595 ;
        RECT 98.855 177.900 99.025 178.475 ;
        RECT 99.255 178.035 99.665 178.340 ;
        RECT 99.955 178.305 100.165 178.705 ;
        RECT 99.835 178.095 100.165 178.305 ;
        RECT 100.410 178.305 100.630 178.705 ;
        RECT 101.105 178.530 101.560 179.295 ;
        RECT 100.410 178.095 100.885 178.305 ;
        RECT 101.075 178.105 101.565 178.305 ;
        RECT 98.855 177.865 99.055 177.900 ;
        RECT 100.385 177.865 101.560 177.925 ;
        RECT 98.855 177.755 101.560 177.865 ;
        RECT 98.915 177.695 100.715 177.755 ;
        RECT 100.385 177.665 100.715 177.695 ;
        RECT 97.590 177.415 98.255 177.585 ;
        RECT 97.585 176.745 97.915 177.245 ;
        RECT 98.085 176.915 98.255 177.415 ;
        RECT 98.515 176.915 98.775 177.595 ;
        RECT 98.945 176.745 99.195 177.525 ;
        RECT 99.445 177.495 100.280 177.505 ;
        RECT 100.870 177.495 101.055 177.585 ;
        RECT 99.445 177.295 101.055 177.495 ;
        RECT 99.445 176.915 99.695 177.295 ;
        RECT 100.825 177.255 101.055 177.295 ;
        RECT 101.305 177.135 101.560 177.755 ;
        RECT 99.865 176.745 100.220 177.125 ;
        RECT 101.225 176.915 101.560 177.135 ;
        RECT 101.740 177.695 102.075 179.115 ;
        RECT 102.255 178.925 103.000 179.295 ;
        RECT 103.565 178.755 103.820 179.115 ;
        RECT 104.000 178.925 104.330 179.295 ;
        RECT 104.510 178.755 104.735 179.115 ;
        RECT 102.250 178.565 104.735 178.755 ;
        RECT 102.250 177.875 102.475 178.565 ;
        RECT 104.955 178.525 108.465 179.295 ;
        RECT 102.675 178.055 102.955 178.385 ;
        RECT 103.135 178.055 103.710 178.385 ;
        RECT 103.890 178.055 104.325 178.385 ;
        RECT 104.505 178.055 104.775 178.385 ;
        RECT 104.955 178.005 106.605 178.525 ;
        RECT 102.250 177.695 104.745 177.875 ;
        RECT 106.775 177.835 108.465 178.355 ;
        RECT 101.740 176.925 102.005 177.695 ;
        RECT 102.175 176.745 102.505 177.465 ;
        RECT 102.695 177.285 103.885 177.515 ;
        RECT 102.695 176.925 102.955 177.285 ;
        RECT 103.125 176.745 103.455 177.115 ;
        RECT 103.625 176.925 103.885 177.285 ;
        RECT 104.455 176.925 104.745 177.695 ;
        RECT 104.955 176.745 108.465 177.835 ;
        RECT 109.555 176.915 109.835 179.015 ;
        RECT 110.065 178.835 110.235 179.295 ;
        RECT 110.505 178.905 111.755 179.085 ;
        RECT 110.890 178.665 111.255 178.735 ;
        RECT 110.005 178.485 111.255 178.665 ;
        RECT 111.425 178.685 111.755 178.905 ;
        RECT 111.925 178.855 112.095 179.295 ;
        RECT 112.265 178.685 112.605 179.100 ;
        RECT 111.425 178.515 112.605 178.685 ;
        RECT 110.005 177.885 110.280 178.485 ;
        RECT 110.450 178.055 110.805 178.305 ;
        RECT 111.000 178.275 111.465 178.305 ;
        RECT 110.995 178.105 111.465 178.275 ;
        RECT 111.000 178.055 111.465 178.105 ;
        RECT 111.635 178.055 111.965 178.305 ;
        RECT 112.140 178.105 112.605 178.305 ;
        RECT 111.785 177.935 111.965 178.055 ;
        RECT 110.005 177.675 111.615 177.885 ;
        RECT 111.785 177.765 112.115 177.935 ;
        RECT 111.205 177.575 111.615 177.675 ;
        RECT 110.025 176.745 110.810 177.505 ;
        RECT 111.205 176.915 111.590 177.575 ;
        RECT 111.915 176.975 112.115 177.765 ;
        RECT 112.285 176.745 112.605 177.925 ;
        RECT 112.785 176.925 113.045 179.115 ;
        RECT 113.305 178.925 113.975 179.295 ;
        RECT 114.155 178.745 114.465 179.115 ;
        RECT 113.235 178.545 114.465 178.745 ;
        RECT 113.235 177.875 113.525 178.545 ;
        RECT 114.645 178.365 114.875 179.005 ;
        RECT 115.055 178.565 115.345 179.295 ;
        RECT 116.455 178.570 116.745 179.295 ;
        RECT 117.075 178.735 117.405 179.125 ;
        RECT 117.575 178.905 118.760 179.075 ;
        RECT 119.020 178.825 119.190 179.295 ;
        RECT 117.075 178.555 117.585 178.735 ;
        RECT 113.705 178.055 114.170 178.365 ;
        RECT 114.350 178.055 114.875 178.365 ;
        RECT 115.055 178.055 115.355 178.385 ;
        RECT 116.915 178.095 117.245 178.385 ;
        RECT 117.415 177.925 117.585 178.555 ;
        RECT 117.990 178.645 118.375 178.735 ;
        RECT 119.360 178.645 119.690 179.110 ;
        RECT 117.990 178.475 119.690 178.645 ;
        RECT 119.860 178.475 120.030 179.295 ;
        RECT 120.200 178.475 120.885 179.115 ;
        RECT 121.060 178.530 121.515 179.295 ;
        RECT 121.790 178.915 123.090 179.125 ;
        RECT 123.345 178.935 123.675 179.295 ;
        RECT 122.920 178.765 123.090 178.915 ;
        RECT 123.845 178.795 124.105 179.125 ;
        RECT 117.755 178.095 118.085 178.305 ;
        RECT 118.265 178.055 118.645 178.305 ;
        RECT 113.235 177.655 114.005 177.875 ;
        RECT 113.215 176.745 113.555 177.475 ;
        RECT 113.735 176.925 114.005 177.655 ;
        RECT 114.185 177.635 115.345 177.875 ;
        RECT 114.185 176.925 114.415 177.635 ;
        RECT 114.585 176.745 114.915 177.455 ;
        RECT 115.085 176.925 115.345 177.635 ;
        RECT 116.455 176.745 116.745 177.910 ;
        RECT 117.070 177.755 118.155 177.925 ;
        RECT 117.070 176.915 117.370 177.755 ;
        RECT 117.565 176.745 117.815 177.585 ;
        RECT 117.985 177.505 118.155 177.755 ;
        RECT 118.325 177.675 118.645 178.055 ;
        RECT 118.835 178.095 119.320 178.305 ;
        RECT 119.510 178.095 119.960 178.305 ;
        RECT 120.130 178.095 120.465 178.305 ;
        RECT 118.835 177.935 119.210 178.095 ;
        RECT 118.815 177.765 119.210 177.935 ;
        RECT 120.130 177.925 120.300 178.095 ;
        RECT 118.835 177.675 119.210 177.765 ;
        RECT 119.380 177.755 120.300 177.925 ;
        RECT 119.380 177.505 119.550 177.755 ;
        RECT 117.985 177.335 119.550 177.505 ;
        RECT 118.405 176.915 119.210 177.335 ;
        RECT 119.720 176.745 120.050 177.585 ;
        RECT 120.635 177.505 120.885 178.475 ;
        RECT 121.990 178.305 122.210 178.705 ;
        RECT 121.055 178.105 121.545 178.305 ;
        RECT 121.735 178.095 122.210 178.305 ;
        RECT 122.455 178.305 122.665 178.705 ;
        RECT 122.920 178.640 123.675 178.765 ;
        RECT 122.920 178.595 123.765 178.640 ;
        RECT 123.495 178.475 123.765 178.595 ;
        RECT 122.455 178.095 122.785 178.305 ;
        RECT 122.955 178.035 123.365 178.340 ;
        RECT 120.220 176.915 120.885 177.505 ;
        RECT 121.060 177.865 122.235 177.925 ;
        RECT 123.595 177.900 123.765 178.475 ;
        RECT 123.565 177.865 123.765 177.900 ;
        RECT 121.060 177.755 123.765 177.865 ;
        RECT 121.060 177.135 121.315 177.755 ;
        RECT 121.905 177.695 123.705 177.755 ;
        RECT 121.905 177.665 122.235 177.695 ;
        RECT 123.935 177.595 124.105 178.795 ;
        RECT 124.280 178.530 124.735 179.295 ;
        RECT 125.010 178.915 126.310 179.125 ;
        RECT 126.565 178.935 126.895 179.295 ;
        RECT 126.140 178.765 126.310 178.915 ;
        RECT 127.065 178.795 127.325 179.125 ;
        RECT 127.095 178.785 127.325 178.795 ;
        RECT 125.210 178.305 125.430 178.705 ;
        RECT 124.275 178.105 124.765 178.305 ;
        RECT 124.955 178.095 125.430 178.305 ;
        RECT 125.675 178.305 125.885 178.705 ;
        RECT 126.140 178.640 126.895 178.765 ;
        RECT 126.140 178.595 126.985 178.640 ;
        RECT 126.715 178.475 126.985 178.595 ;
        RECT 125.675 178.095 126.005 178.305 ;
        RECT 126.175 178.035 126.585 178.340 ;
        RECT 121.565 177.495 121.750 177.585 ;
        RECT 122.340 177.495 123.175 177.505 ;
        RECT 121.565 177.295 123.175 177.495 ;
        RECT 121.565 177.255 121.795 177.295 ;
        RECT 121.060 176.915 121.395 177.135 ;
        RECT 122.400 176.745 122.755 177.125 ;
        RECT 122.925 176.915 123.175 177.295 ;
        RECT 123.425 176.745 123.675 177.525 ;
        RECT 123.845 176.915 124.105 177.595 ;
        RECT 124.280 177.865 125.455 177.925 ;
        RECT 126.815 177.900 126.985 178.475 ;
        RECT 126.785 177.865 126.985 177.900 ;
        RECT 124.280 177.755 126.985 177.865 ;
        RECT 124.280 177.135 124.535 177.755 ;
        RECT 125.125 177.695 126.925 177.755 ;
        RECT 125.125 177.665 125.455 177.695 ;
        RECT 127.155 177.595 127.325 178.785 ;
        RECT 127.770 178.485 128.015 179.090 ;
        RECT 128.235 178.760 128.745 179.295 ;
        RECT 124.785 177.495 124.970 177.585 ;
        RECT 125.560 177.495 126.395 177.505 ;
        RECT 124.785 177.295 126.395 177.495 ;
        RECT 124.785 177.255 125.015 177.295 ;
        RECT 124.280 176.915 124.615 177.135 ;
        RECT 125.620 176.745 125.975 177.125 ;
        RECT 126.145 176.915 126.395 177.295 ;
        RECT 126.645 176.745 126.895 177.525 ;
        RECT 127.065 176.915 127.325 177.595 ;
        RECT 127.495 178.315 128.725 178.485 ;
        RECT 127.495 177.505 127.835 178.315 ;
        RECT 128.005 177.750 128.755 177.940 ;
        RECT 127.495 177.095 128.010 177.505 ;
        RECT 128.245 176.745 128.415 177.505 ;
        RECT 128.585 177.085 128.755 177.750 ;
        RECT 128.925 177.765 129.115 179.125 ;
        RECT 129.285 178.615 129.560 179.125 ;
        RECT 129.750 178.760 130.280 179.125 ;
        RECT 130.705 178.895 131.035 179.295 ;
        RECT 130.105 178.725 130.280 178.760 ;
        RECT 129.285 178.445 129.565 178.615 ;
        RECT 129.285 177.965 129.560 178.445 ;
        RECT 129.765 177.765 129.935 178.565 ;
        RECT 128.925 177.595 129.935 177.765 ;
        RECT 130.105 178.555 131.035 178.725 ;
        RECT 131.205 178.555 131.460 179.125 ;
        RECT 131.725 178.745 131.895 179.125 ;
        RECT 132.075 178.915 132.405 179.295 ;
        RECT 131.725 178.575 132.390 178.745 ;
        RECT 132.585 178.620 132.845 179.125 ;
        RECT 130.105 177.425 130.275 178.555 ;
        RECT 130.865 178.385 131.035 178.555 ;
        RECT 129.150 177.255 130.275 177.425 ;
        RECT 130.445 178.055 130.640 178.385 ;
        RECT 130.865 178.055 131.120 178.385 ;
        RECT 130.445 177.085 130.615 178.055 ;
        RECT 131.290 177.885 131.460 178.555 ;
        RECT 131.655 178.025 131.985 178.395 ;
        RECT 132.220 178.320 132.390 178.575 ;
        RECT 128.585 176.915 130.615 177.085 ;
        RECT 130.785 176.745 130.955 177.885 ;
        RECT 131.125 176.915 131.460 177.885 ;
        RECT 132.220 177.990 132.505 178.320 ;
        RECT 132.220 177.845 132.390 177.990 ;
        RECT 131.725 177.675 132.390 177.845 ;
        RECT 132.675 177.820 132.845 178.620 ;
        RECT 131.725 176.915 131.895 177.675 ;
        RECT 132.075 176.745 132.405 177.505 ;
        RECT 132.575 176.915 132.845 177.820 ;
        RECT 133.015 178.555 133.400 179.125 ;
        RECT 133.570 178.835 133.895 179.295 ;
        RECT 134.415 178.665 134.695 179.125 ;
        RECT 133.015 177.885 133.295 178.555 ;
        RECT 133.570 178.495 134.695 178.665 ;
        RECT 133.570 178.385 134.020 178.495 ;
        RECT 133.465 178.055 134.020 178.385 ;
        RECT 134.885 178.325 135.285 179.125 ;
        RECT 135.685 178.835 135.955 179.295 ;
        RECT 136.125 178.665 136.410 179.125 ;
        RECT 133.015 176.915 133.400 177.885 ;
        RECT 133.570 177.595 134.020 178.055 ;
        RECT 134.190 177.765 135.285 178.325 ;
        RECT 133.570 177.375 134.695 177.595 ;
        RECT 133.570 176.745 133.895 177.205 ;
        RECT 134.415 176.915 134.695 177.375 ;
        RECT 134.885 176.915 135.285 177.765 ;
        RECT 135.455 178.495 136.410 178.665 ;
        RECT 137.615 178.545 138.825 179.295 ;
        RECT 135.455 177.595 135.665 178.495 ;
        RECT 135.835 177.765 136.525 178.325 ;
        RECT 137.615 177.835 138.135 178.375 ;
        RECT 138.305 178.005 138.825 178.545 ;
        RECT 135.455 177.375 136.410 177.595 ;
        RECT 135.685 176.745 135.955 177.205 ;
        RECT 136.125 176.915 136.410 177.375 ;
        RECT 137.615 176.745 138.825 177.835 ;
        RECT 13.330 176.575 138.910 176.745 ;
        RECT 13.415 175.485 14.625 176.575 ;
        RECT 14.795 176.140 20.140 176.575 ;
        RECT 13.415 174.775 13.935 175.315 ;
        RECT 14.105 174.945 14.625 175.485 ;
        RECT 13.415 174.025 14.625 174.775 ;
        RECT 16.380 174.570 16.720 175.400 ;
        RECT 18.200 174.890 18.550 176.140 ;
        RECT 21.245 175.965 21.575 176.395 ;
        RECT 21.755 176.135 21.950 176.575 ;
        RECT 22.120 175.965 22.450 176.395 ;
        RECT 21.245 175.795 22.450 175.965 ;
        RECT 21.245 175.465 22.140 175.795 ;
        RECT 22.620 175.625 22.895 176.395 ;
        RECT 22.310 175.435 22.895 175.625 ;
        RECT 23.075 175.485 25.665 176.575 ;
        RECT 21.250 174.935 21.545 175.265 ;
        RECT 21.725 174.935 22.140 175.265 ;
        RECT 14.795 174.025 20.140 174.570 ;
        RECT 21.245 174.025 21.545 174.755 ;
        RECT 21.725 174.315 21.955 174.935 ;
        RECT 22.310 174.765 22.485 175.435 ;
        RECT 22.155 174.585 22.485 174.765 ;
        RECT 22.655 174.615 22.895 175.265 ;
        RECT 23.075 174.795 24.285 175.315 ;
        RECT 24.455 174.965 25.665 175.485 ;
        RECT 26.295 175.410 26.585 176.575 ;
        RECT 26.755 175.485 28.425 176.575 ;
        RECT 29.055 176.065 30.245 176.355 ;
        RECT 26.755 174.795 27.505 175.315 ;
        RECT 27.675 174.965 28.425 175.485 ;
        RECT 29.075 175.725 30.245 175.895 ;
        RECT 30.415 175.775 30.695 176.575 ;
        RECT 29.075 175.435 29.400 175.725 ;
        RECT 30.075 175.605 30.245 175.725 ;
        RECT 29.570 175.265 29.765 175.555 ;
        RECT 30.075 175.435 30.735 175.605 ;
        RECT 30.905 175.435 31.180 176.405 ;
        RECT 32.275 175.435 32.555 176.575 ;
        RECT 30.565 175.265 30.735 175.435 ;
        RECT 29.055 174.935 29.400 175.265 ;
        RECT 29.570 174.935 30.395 175.265 ;
        RECT 30.565 174.935 30.840 175.265 ;
        RECT 22.155 174.205 22.380 174.585 ;
        RECT 22.550 174.025 22.880 174.415 ;
        RECT 23.075 174.025 25.665 174.795 ;
        RECT 26.295 174.025 26.585 174.750 ;
        RECT 26.755 174.025 28.425 174.795 ;
        RECT 30.565 174.765 30.735 174.935 ;
        RECT 29.070 174.595 30.735 174.765 ;
        RECT 31.010 174.700 31.180 175.435 ;
        RECT 32.725 175.425 33.055 176.405 ;
        RECT 33.225 175.435 33.485 176.575 ;
        RECT 33.860 175.605 34.190 176.405 ;
        RECT 34.360 175.775 34.690 176.575 ;
        RECT 34.990 175.605 35.320 176.405 ;
        RECT 35.965 175.775 36.215 176.575 ;
        RECT 33.860 175.435 36.295 175.605 ;
        RECT 36.485 175.435 36.655 176.575 ;
        RECT 36.825 175.435 37.165 176.405 ;
        RECT 32.285 174.995 32.620 175.265 ;
        RECT 32.790 174.825 32.960 175.425 ;
        RECT 33.130 175.015 33.465 175.265 ;
        RECT 33.655 175.015 34.005 175.265 ;
        RECT 29.070 174.245 29.325 174.595 ;
        RECT 29.495 174.025 29.825 174.425 ;
        RECT 29.995 174.245 30.165 174.595 ;
        RECT 30.335 174.025 30.715 174.425 ;
        RECT 30.905 174.355 31.180 174.700 ;
        RECT 32.275 174.025 32.585 174.825 ;
        RECT 32.790 174.195 33.485 174.825 ;
        RECT 34.190 174.805 34.360 175.435 ;
        RECT 34.530 175.015 34.860 175.215 ;
        RECT 35.030 175.015 35.360 175.215 ;
        RECT 35.530 175.015 35.950 175.215 ;
        RECT 36.125 175.185 36.295 175.435 ;
        RECT 36.125 175.015 36.820 175.185 ;
        RECT 33.860 174.195 34.360 174.805 ;
        RECT 34.990 174.675 36.215 174.845 ;
        RECT 36.990 174.825 37.165 175.435 ;
        RECT 34.990 174.195 35.320 174.675 ;
        RECT 35.490 174.025 35.715 174.485 ;
        RECT 35.885 174.195 36.215 174.675 ;
        RECT 36.405 174.025 36.655 174.825 ;
        RECT 36.825 174.195 37.165 174.825 ;
        RECT 37.335 175.435 37.610 176.405 ;
        RECT 37.820 175.775 38.100 176.575 ;
        RECT 38.270 176.065 39.885 176.395 ;
        RECT 38.270 175.725 39.445 175.895 ;
        RECT 38.270 175.605 38.440 175.725 ;
        RECT 37.780 175.435 38.440 175.605 ;
        RECT 37.335 174.700 37.505 175.435 ;
        RECT 37.780 175.265 37.950 175.435 ;
        RECT 38.700 175.265 38.945 175.555 ;
        RECT 39.115 175.435 39.445 175.725 ;
        RECT 39.705 175.265 39.875 175.825 ;
        RECT 40.125 175.435 40.385 176.575 ;
        RECT 40.740 175.605 41.130 175.780 ;
        RECT 41.615 175.775 41.945 176.575 ;
        RECT 42.115 175.785 42.650 176.405 ;
        RECT 40.740 175.435 42.165 175.605 ;
        RECT 37.675 174.935 37.950 175.265 ;
        RECT 38.120 174.935 38.945 175.265 ;
        RECT 39.160 174.935 39.875 175.265 ;
        RECT 40.045 175.015 40.380 175.265 ;
        RECT 37.780 174.765 37.950 174.935 ;
        RECT 39.625 174.845 39.875 174.935 ;
        RECT 37.335 174.355 37.610 174.700 ;
        RECT 37.780 174.595 39.445 174.765 ;
        RECT 37.800 174.025 38.175 174.425 ;
        RECT 38.345 174.245 38.515 174.595 ;
        RECT 38.685 174.025 39.015 174.425 ;
        RECT 39.185 174.195 39.445 174.595 ;
        RECT 39.625 174.425 39.955 174.845 ;
        RECT 40.125 174.025 40.385 174.845 ;
        RECT 40.615 174.705 40.970 175.265 ;
        RECT 41.140 174.535 41.310 175.435 ;
        RECT 41.480 174.705 41.745 175.265 ;
        RECT 41.995 174.935 42.165 175.435 ;
        RECT 42.335 174.765 42.650 175.785 ;
        RECT 42.855 175.485 46.365 176.575 ;
        RECT 46.620 175.955 46.795 176.405 ;
        RECT 46.965 176.135 47.295 176.575 ;
        RECT 47.600 175.985 47.770 176.405 ;
        RECT 48.005 176.165 48.675 176.575 ;
        RECT 48.890 175.985 49.060 176.405 ;
        RECT 49.260 176.165 49.590 176.575 ;
        RECT 46.620 175.785 47.250 175.955 ;
        RECT 40.720 174.025 40.960 174.535 ;
        RECT 41.140 174.205 41.420 174.535 ;
        RECT 41.650 174.025 41.865 174.535 ;
        RECT 42.035 174.195 42.650 174.765 ;
        RECT 42.855 174.795 44.505 175.315 ;
        RECT 44.675 174.965 46.365 175.485 ;
        RECT 46.535 174.935 46.900 175.615 ;
        RECT 47.080 175.265 47.250 175.785 ;
        RECT 47.600 175.815 49.615 175.985 ;
        RECT 47.080 174.935 47.430 175.265 ;
        RECT 42.855 174.025 46.365 174.795 ;
        RECT 47.080 174.765 47.250 174.935 ;
        RECT 46.620 174.595 47.250 174.765 ;
        RECT 46.620 174.195 46.795 174.595 ;
        RECT 47.600 174.525 47.770 175.815 ;
        RECT 46.965 174.025 47.295 174.405 ;
        RECT 47.540 174.195 47.770 174.525 ;
        RECT 47.970 174.360 48.250 175.635 ;
        RECT 48.475 175.555 48.745 175.635 ;
        RECT 48.435 175.385 48.745 175.555 ;
        RECT 48.475 174.360 48.745 175.385 ;
        RECT 48.935 174.605 49.275 175.635 ;
        RECT 49.445 175.265 49.615 175.815 ;
        RECT 49.785 175.435 50.045 176.405 ;
        RECT 50.225 175.435 50.555 176.575 ;
        RECT 51.085 175.605 51.415 176.390 ;
        RECT 50.735 175.435 51.415 175.605 ;
        RECT 49.445 174.935 49.705 175.265 ;
        RECT 49.875 174.745 50.045 175.435 ;
        RECT 50.215 175.015 50.565 175.265 ;
        RECT 50.735 174.835 50.905 175.435 ;
        RECT 52.055 175.410 52.345 176.575 ;
        RECT 52.515 175.740 52.900 176.575 ;
        RECT 53.070 175.570 53.330 176.375 ;
        RECT 53.500 175.740 53.760 176.575 ;
        RECT 53.930 175.570 54.185 176.375 ;
        RECT 54.360 175.740 54.620 176.575 ;
        RECT 54.790 175.570 55.045 176.375 ;
        RECT 55.220 175.740 55.565 176.575 ;
        RECT 52.515 175.400 55.545 175.570 ;
        RECT 55.735 175.485 59.245 176.575 ;
        RECT 51.075 175.015 51.425 175.265 ;
        RECT 52.515 174.835 52.815 175.400 ;
        RECT 52.990 175.005 55.205 175.230 ;
        RECT 55.375 174.835 55.545 175.400 ;
        RECT 49.205 174.025 49.535 174.405 ;
        RECT 49.705 174.280 50.045 174.745 ;
        RECT 49.705 174.235 50.040 174.280 ;
        RECT 50.225 174.025 50.495 174.835 ;
        RECT 50.665 174.195 50.995 174.835 ;
        RECT 51.165 174.025 51.405 174.835 ;
        RECT 52.055 174.025 52.345 174.750 ;
        RECT 52.515 174.665 55.545 174.835 ;
        RECT 55.735 174.795 57.385 175.315 ;
        RECT 57.555 174.965 59.245 175.485 ;
        RECT 60.345 175.465 60.640 176.575 ;
        RECT 60.820 175.265 61.070 176.400 ;
        RECT 61.240 175.465 61.500 176.575 ;
        RECT 61.670 175.675 61.930 176.400 ;
        RECT 62.100 175.845 62.360 176.575 ;
        RECT 62.530 175.675 62.790 176.400 ;
        RECT 62.960 175.845 63.220 176.575 ;
        RECT 63.390 175.675 63.650 176.400 ;
        RECT 63.820 175.845 64.080 176.575 ;
        RECT 64.250 175.675 64.510 176.400 ;
        RECT 64.680 175.845 64.975 176.575 ;
        RECT 61.670 175.435 64.980 175.675 ;
        RECT 53.035 174.025 53.335 174.495 ;
        RECT 53.505 174.220 53.760 174.665 ;
        RECT 53.930 174.025 54.190 174.495 ;
        RECT 54.360 174.220 54.620 174.665 ;
        RECT 54.790 174.025 55.085 174.495 ;
        RECT 55.735 174.025 59.245 174.795 ;
        RECT 60.335 174.655 60.650 175.265 ;
        RECT 60.820 175.015 63.840 175.265 ;
        RECT 60.395 174.025 60.640 174.485 ;
        RECT 60.820 174.205 61.070 175.015 ;
        RECT 64.010 174.845 64.980 175.435 ;
        RECT 65.405 175.555 65.735 176.405 ;
        RECT 65.905 175.725 66.075 176.575 ;
        RECT 66.245 175.555 66.575 176.405 ;
        RECT 66.745 175.725 66.915 176.575 ;
        RECT 67.085 175.555 67.415 176.405 ;
        RECT 67.585 175.775 67.755 176.575 ;
        RECT 67.925 175.555 68.255 176.405 ;
        RECT 68.425 175.775 68.595 176.575 ;
        RECT 68.765 175.555 69.095 176.405 ;
        RECT 69.265 175.775 69.435 176.575 ;
        RECT 69.605 175.555 69.935 176.405 ;
        RECT 70.105 175.775 70.275 176.575 ;
        RECT 70.445 175.555 70.775 176.405 ;
        RECT 70.945 175.775 71.115 176.575 ;
        RECT 71.285 175.555 71.615 176.405 ;
        RECT 71.785 175.775 71.955 176.575 ;
        RECT 72.125 175.555 72.455 176.405 ;
        RECT 72.625 175.775 72.795 176.575 ;
        RECT 72.965 175.555 73.295 176.405 ;
        RECT 73.465 175.775 73.635 176.575 ;
        RECT 73.805 175.555 74.135 176.405 ;
        RECT 74.305 175.775 74.475 176.575 ;
        RECT 74.645 175.555 74.975 176.405 ;
        RECT 75.145 175.775 75.315 176.575 ;
        RECT 75.485 175.555 75.815 176.405 ;
        RECT 75.985 175.775 76.155 176.575 ;
        RECT 65.405 175.385 66.915 175.555 ;
        RECT 67.085 175.385 69.435 175.555 ;
        RECT 69.605 175.385 76.265 175.555 ;
        RECT 76.435 175.435 76.695 176.575 ;
        RECT 76.865 175.425 77.195 176.405 ;
        RECT 77.365 175.435 77.645 176.575 ;
        RECT 66.745 175.215 66.915 175.385 ;
        RECT 69.260 175.215 69.435 175.385 ;
        RECT 65.400 175.015 66.575 175.215 ;
        RECT 66.745 175.015 69.055 175.215 ;
        RECT 69.260 175.015 75.820 175.215 ;
        RECT 66.745 174.845 66.915 175.015 ;
        RECT 69.260 174.845 69.435 175.015 ;
        RECT 75.990 174.845 76.265 175.385 ;
        RECT 76.455 175.015 76.790 175.265 ;
        RECT 61.670 174.675 64.980 174.845 ;
        RECT 65.405 174.675 66.915 174.845 ;
        RECT 67.085 174.675 69.435 174.845 ;
        RECT 69.605 174.675 76.265 174.845 ;
        RECT 76.960 174.825 77.130 175.425 ;
        RECT 77.815 175.410 78.105 176.575 ;
        RECT 78.795 175.515 79.125 176.360 ;
        RECT 79.295 175.565 79.465 176.575 ;
        RECT 79.635 175.845 79.975 176.405 ;
        RECT 80.205 176.075 80.520 176.575 ;
        RECT 80.700 176.105 81.585 176.275 ;
        RECT 78.735 175.435 79.125 175.515 ;
        RECT 79.635 175.470 80.530 175.845 ;
        RECT 78.735 175.385 78.950 175.435 ;
        RECT 77.300 174.995 77.635 175.265 ;
        RECT 61.240 174.025 61.500 174.550 ;
        RECT 61.670 174.220 61.930 174.675 ;
        RECT 62.100 174.025 62.360 174.505 ;
        RECT 62.530 174.220 62.790 174.675 ;
        RECT 62.960 174.025 63.220 174.505 ;
        RECT 63.390 174.220 63.650 174.675 ;
        RECT 63.820 174.025 64.080 174.505 ;
        RECT 64.250 174.220 64.510 174.675 ;
        RECT 64.680 174.025 64.980 174.505 ;
        RECT 65.405 174.200 65.735 174.675 ;
        RECT 65.905 174.025 66.075 174.505 ;
        RECT 66.245 174.200 66.575 174.675 ;
        RECT 66.745 174.025 66.915 174.505 ;
        RECT 67.085 174.200 67.415 174.675 ;
        RECT 67.585 174.025 67.755 174.505 ;
        RECT 67.925 174.200 68.255 174.675 ;
        RECT 68.425 174.025 68.595 174.505 ;
        RECT 68.765 174.200 69.095 174.675 ;
        RECT 69.265 174.025 69.435 174.505 ;
        RECT 69.605 174.200 69.935 174.675 ;
        RECT 69.605 174.195 69.855 174.200 ;
        RECT 70.105 174.025 70.275 174.505 ;
        RECT 70.445 174.200 70.775 174.675 ;
        RECT 70.525 174.195 70.695 174.200 ;
        RECT 70.945 174.025 71.115 174.505 ;
        RECT 71.285 174.200 71.615 174.675 ;
        RECT 71.365 174.195 71.535 174.200 ;
        RECT 71.785 174.025 71.955 174.505 ;
        RECT 72.125 174.200 72.455 174.675 ;
        RECT 72.625 174.025 72.795 174.505 ;
        RECT 72.965 174.200 73.295 174.675 ;
        RECT 73.465 174.025 73.635 174.505 ;
        RECT 73.805 174.200 74.135 174.675 ;
        RECT 74.305 174.025 74.475 174.505 ;
        RECT 74.645 174.200 74.975 174.675 ;
        RECT 75.145 174.025 75.315 174.505 ;
        RECT 75.485 174.200 75.815 174.675 ;
        RECT 75.985 174.025 76.155 174.505 ;
        RECT 76.435 174.195 77.130 174.825 ;
        RECT 77.335 174.025 77.645 174.825 ;
        RECT 78.735 174.805 78.905 175.385 ;
        RECT 79.635 175.265 79.825 175.470 ;
        RECT 80.700 175.265 80.870 176.105 ;
        RECT 81.810 176.075 82.060 176.405 ;
        RECT 79.075 174.935 79.825 175.265 ;
        RECT 79.995 174.935 80.870 175.265 ;
        RECT 78.735 174.765 78.960 174.805 ;
        RECT 79.625 174.765 79.825 174.935 ;
        RECT 77.815 174.025 78.105 174.750 ;
        RECT 78.735 174.680 79.115 174.765 ;
        RECT 78.785 174.245 79.115 174.680 ;
        RECT 79.285 174.025 79.455 174.635 ;
        RECT 79.625 174.240 79.955 174.765 ;
        RECT 80.215 174.025 80.425 174.555 ;
        RECT 80.700 174.475 80.870 174.935 ;
        RECT 81.040 174.975 81.360 175.935 ;
        RECT 81.530 175.185 81.720 175.905 ;
        RECT 81.890 175.005 82.060 176.075 ;
        RECT 82.230 175.775 82.400 176.575 ;
        RECT 82.570 176.130 83.675 176.300 ;
        RECT 82.570 175.515 82.740 176.130 ;
        RECT 83.885 175.980 84.135 176.405 ;
        RECT 84.305 176.115 84.570 176.575 ;
        RECT 82.910 175.595 83.440 175.960 ;
        RECT 83.885 175.850 84.190 175.980 ;
        RECT 82.230 175.425 82.740 175.515 ;
        RECT 82.230 175.255 83.100 175.425 ;
        RECT 82.230 175.185 82.400 175.255 ;
        RECT 82.520 175.005 82.720 175.035 ;
        RECT 81.040 174.645 81.505 174.975 ;
        RECT 81.890 174.705 82.720 175.005 ;
        RECT 81.890 174.475 82.060 174.705 ;
        RECT 80.700 174.305 81.485 174.475 ;
        RECT 81.655 174.305 82.060 174.475 ;
        RECT 82.240 174.025 82.610 174.525 ;
        RECT 82.930 174.475 83.100 175.255 ;
        RECT 83.270 174.895 83.440 175.595 ;
        RECT 83.610 175.065 83.850 175.660 ;
        RECT 83.270 174.675 83.795 174.895 ;
        RECT 84.020 174.745 84.190 175.850 ;
        RECT 83.965 174.615 84.190 174.745 ;
        RECT 84.360 174.655 84.640 175.605 ;
        RECT 83.965 174.475 84.135 174.615 ;
        RECT 82.930 174.305 83.605 174.475 ;
        RECT 83.800 174.305 84.135 174.475 ;
        RECT 84.305 174.025 84.555 174.485 ;
        RECT 84.810 174.285 84.995 176.405 ;
        RECT 85.165 176.075 85.495 176.575 ;
        RECT 85.665 175.905 85.835 176.405 ;
        RECT 85.170 175.735 85.835 175.905 ;
        RECT 86.185 175.905 86.355 176.405 ;
        RECT 86.525 176.075 86.855 176.575 ;
        RECT 86.185 175.735 86.850 175.905 ;
        RECT 85.170 174.745 85.400 175.735 ;
        RECT 85.570 174.915 85.920 175.565 ;
        RECT 86.100 174.915 86.450 175.565 ;
        RECT 86.620 174.745 86.850 175.735 ;
        RECT 85.170 174.575 85.835 174.745 ;
        RECT 85.165 174.025 85.495 174.405 ;
        RECT 85.665 174.285 85.835 174.575 ;
        RECT 86.185 174.575 86.850 174.745 ;
        RECT 86.185 174.285 86.355 174.575 ;
        RECT 86.525 174.025 86.855 174.405 ;
        RECT 87.025 174.285 87.210 176.405 ;
        RECT 87.450 176.115 87.715 176.575 ;
        RECT 87.885 175.980 88.135 176.405 ;
        RECT 88.345 176.130 89.450 176.300 ;
        RECT 87.830 175.850 88.135 175.980 ;
        RECT 87.380 174.655 87.660 175.605 ;
        RECT 87.830 174.745 88.000 175.850 ;
        RECT 88.170 175.065 88.410 175.660 ;
        RECT 88.580 175.595 89.110 175.960 ;
        RECT 88.580 174.895 88.750 175.595 ;
        RECT 89.280 175.515 89.450 176.130 ;
        RECT 89.620 175.775 89.790 176.575 ;
        RECT 89.960 176.075 90.210 176.405 ;
        RECT 90.435 176.105 91.320 176.275 ;
        RECT 89.280 175.425 89.790 175.515 ;
        RECT 87.830 174.615 88.055 174.745 ;
        RECT 88.225 174.675 88.750 174.895 ;
        RECT 88.920 175.255 89.790 175.425 ;
        RECT 87.465 174.025 87.715 174.485 ;
        RECT 87.885 174.475 88.055 174.615 ;
        RECT 88.920 174.475 89.090 175.255 ;
        RECT 89.620 175.185 89.790 175.255 ;
        RECT 89.300 175.005 89.500 175.035 ;
        RECT 89.960 175.005 90.130 176.075 ;
        RECT 90.300 175.185 90.490 175.905 ;
        RECT 89.300 174.705 90.130 175.005 ;
        RECT 90.660 174.975 90.980 175.935 ;
        RECT 87.885 174.305 88.220 174.475 ;
        RECT 88.415 174.305 89.090 174.475 ;
        RECT 89.410 174.025 89.780 174.525 ;
        RECT 89.960 174.475 90.130 174.705 ;
        RECT 90.515 174.645 90.980 174.975 ;
        RECT 91.150 175.265 91.320 176.105 ;
        RECT 91.500 176.075 91.815 176.575 ;
        RECT 92.045 175.845 92.385 176.405 ;
        RECT 91.490 175.470 92.385 175.845 ;
        RECT 92.555 175.565 92.725 176.575 ;
        RECT 92.195 175.265 92.385 175.470 ;
        RECT 92.895 175.515 93.225 176.360 ;
        RECT 92.895 175.435 93.285 175.515 ;
        RECT 93.455 175.485 95.125 176.575 ;
        RECT 95.355 175.515 95.685 176.360 ;
        RECT 95.855 175.565 96.025 176.575 ;
        RECT 96.195 175.845 96.535 176.405 ;
        RECT 96.765 176.075 97.080 176.575 ;
        RECT 97.260 176.105 98.145 176.275 ;
        RECT 93.070 175.385 93.285 175.435 ;
        RECT 91.150 174.935 92.025 175.265 ;
        RECT 92.195 174.935 92.945 175.265 ;
        RECT 91.150 174.475 91.320 174.935 ;
        RECT 92.195 174.765 92.395 174.935 ;
        RECT 93.115 174.805 93.285 175.385 ;
        RECT 93.060 174.765 93.285 174.805 ;
        RECT 89.960 174.305 90.365 174.475 ;
        RECT 90.535 174.305 91.320 174.475 ;
        RECT 91.595 174.025 91.805 174.555 ;
        RECT 92.065 174.240 92.395 174.765 ;
        RECT 92.905 174.680 93.285 174.765 ;
        RECT 93.455 174.795 94.205 175.315 ;
        RECT 94.375 174.965 95.125 175.485 ;
        RECT 95.295 175.435 95.685 175.515 ;
        RECT 96.195 175.470 97.090 175.845 ;
        RECT 95.295 175.385 95.510 175.435 ;
        RECT 95.295 174.805 95.465 175.385 ;
        RECT 96.195 175.265 96.385 175.470 ;
        RECT 97.260 175.265 97.430 176.105 ;
        RECT 98.370 176.075 98.620 176.405 ;
        RECT 95.635 174.935 96.385 175.265 ;
        RECT 96.555 174.935 97.430 175.265 ;
        RECT 92.565 174.025 92.735 174.635 ;
        RECT 92.905 174.245 93.235 174.680 ;
        RECT 93.455 174.025 95.125 174.795 ;
        RECT 95.295 174.765 95.520 174.805 ;
        RECT 96.185 174.765 96.385 174.935 ;
        RECT 95.295 174.680 95.675 174.765 ;
        RECT 95.345 174.245 95.675 174.680 ;
        RECT 95.845 174.025 96.015 174.635 ;
        RECT 96.185 174.240 96.515 174.765 ;
        RECT 96.775 174.025 96.985 174.555 ;
        RECT 97.260 174.475 97.430 174.935 ;
        RECT 97.600 174.975 97.920 175.935 ;
        RECT 98.090 175.185 98.280 175.905 ;
        RECT 98.450 175.005 98.620 176.075 ;
        RECT 98.790 175.775 98.960 176.575 ;
        RECT 99.130 176.130 100.235 176.300 ;
        RECT 99.130 175.515 99.300 176.130 ;
        RECT 100.445 175.980 100.695 176.405 ;
        RECT 100.865 176.115 101.130 176.575 ;
        RECT 99.470 175.595 100.000 175.960 ;
        RECT 100.445 175.850 100.750 175.980 ;
        RECT 98.790 175.425 99.300 175.515 ;
        RECT 98.790 175.255 99.660 175.425 ;
        RECT 98.790 175.185 98.960 175.255 ;
        RECT 99.080 175.005 99.280 175.035 ;
        RECT 97.600 174.645 98.065 174.975 ;
        RECT 98.450 174.705 99.280 175.005 ;
        RECT 98.450 174.475 98.620 174.705 ;
        RECT 97.260 174.305 98.045 174.475 ;
        RECT 98.215 174.305 98.620 174.475 ;
        RECT 98.800 174.025 99.170 174.525 ;
        RECT 99.490 174.475 99.660 175.255 ;
        RECT 99.830 174.895 100.000 175.595 ;
        RECT 100.170 175.065 100.410 175.660 ;
        RECT 99.830 174.675 100.355 174.895 ;
        RECT 100.580 174.745 100.750 175.850 ;
        RECT 100.525 174.615 100.750 174.745 ;
        RECT 100.920 174.655 101.200 175.605 ;
        RECT 100.525 174.475 100.695 174.615 ;
        RECT 99.490 174.305 100.165 174.475 ;
        RECT 100.360 174.305 100.695 174.475 ;
        RECT 100.865 174.025 101.115 174.485 ;
        RECT 101.370 174.285 101.555 176.405 ;
        RECT 101.725 176.075 102.055 176.575 ;
        RECT 102.225 175.905 102.395 176.405 ;
        RECT 101.730 175.735 102.395 175.905 ;
        RECT 101.730 174.745 101.960 175.735 ;
        RECT 102.130 174.915 102.480 175.565 ;
        RECT 103.575 175.410 103.865 176.575 ;
        RECT 104.150 175.945 104.435 176.405 ;
        RECT 104.605 176.115 104.875 176.575 ;
        RECT 104.150 175.725 105.105 175.945 ;
        RECT 104.035 174.995 104.725 175.555 ;
        RECT 104.895 174.825 105.105 175.725 ;
        RECT 101.730 174.575 102.395 174.745 ;
        RECT 101.725 174.025 102.055 174.405 ;
        RECT 102.225 174.285 102.395 174.575 ;
        RECT 103.575 174.025 103.865 174.750 ;
        RECT 104.150 174.655 105.105 174.825 ;
        RECT 105.275 175.555 105.675 176.405 ;
        RECT 105.865 175.945 106.145 176.405 ;
        RECT 106.665 176.115 106.990 176.575 ;
        RECT 105.865 175.725 106.990 175.945 ;
        RECT 105.275 174.995 106.370 175.555 ;
        RECT 106.540 175.265 106.990 175.725 ;
        RECT 107.160 175.435 107.545 176.405 ;
        RECT 104.150 174.195 104.435 174.655 ;
        RECT 104.605 174.025 104.875 174.485 ;
        RECT 105.275 174.195 105.675 174.995 ;
        RECT 106.540 174.935 107.095 175.265 ;
        RECT 106.540 174.825 106.990 174.935 ;
        RECT 105.865 174.655 106.990 174.825 ;
        RECT 107.265 174.765 107.545 175.435 ;
        RECT 105.865 174.195 106.145 174.655 ;
        RECT 106.665 174.025 106.990 174.485 ;
        RECT 107.160 174.195 107.545 174.765 ;
        RECT 107.715 175.775 108.155 176.405 ;
        RECT 107.715 174.765 108.025 175.775 ;
        RECT 108.330 175.725 108.645 176.575 ;
        RECT 108.815 176.235 110.245 176.405 ;
        RECT 108.815 175.555 108.985 176.235 ;
        RECT 108.195 175.385 108.985 175.555 ;
        RECT 108.195 174.935 108.365 175.385 ;
        RECT 109.155 175.265 109.355 176.065 ;
        RECT 108.535 174.935 108.925 175.215 ;
        RECT 109.110 174.935 109.355 175.265 ;
        RECT 109.555 174.935 109.805 176.065 ;
        RECT 109.995 175.605 110.245 176.235 ;
        RECT 110.425 175.775 110.755 176.575 ;
        RECT 109.995 175.435 110.765 175.605 ;
        RECT 110.020 174.935 110.425 175.265 ;
        RECT 110.595 174.765 110.765 175.435 ;
        RECT 107.715 174.205 108.155 174.765 ;
        RECT 108.325 174.025 108.775 174.765 ;
        RECT 108.945 174.595 110.105 174.765 ;
        RECT 108.945 174.195 109.115 174.595 ;
        RECT 109.285 174.025 109.705 174.425 ;
        RECT 109.875 174.195 110.105 174.595 ;
        RECT 110.275 174.195 110.765 174.765 ;
        RECT 110.945 175.515 111.275 176.365 ;
        RECT 110.945 175.385 111.165 175.515 ;
        RECT 111.445 175.435 111.695 176.575 ;
        RECT 111.885 175.935 112.135 176.355 ;
        RECT 112.365 176.105 112.695 176.575 ;
        RECT 112.925 175.935 113.175 176.355 ;
        RECT 111.885 175.765 113.175 175.935 ;
        RECT 113.355 175.935 113.685 176.365 ;
        RECT 113.355 175.765 113.810 175.935 ;
        RECT 110.945 174.750 111.135 175.385 ;
        RECT 111.875 175.265 112.090 175.595 ;
        RECT 111.305 174.935 111.615 175.265 ;
        RECT 111.785 174.935 112.090 175.265 ;
        RECT 112.265 174.935 112.550 175.595 ;
        RECT 112.745 174.935 113.010 175.595 ;
        RECT 113.225 174.935 113.470 175.595 ;
        RECT 111.445 174.765 111.615 174.935 ;
        RECT 113.640 174.765 113.810 175.765 ;
        RECT 114.155 175.485 115.825 176.575 ;
        RECT 110.945 174.240 111.275 174.750 ;
        RECT 111.445 174.595 113.810 174.765 ;
        RECT 114.155 174.795 114.905 175.315 ;
        RECT 115.075 174.965 115.825 175.485 ;
        RECT 116.015 175.685 116.275 176.395 ;
        RECT 116.445 175.865 116.775 176.575 ;
        RECT 116.945 175.685 117.175 176.395 ;
        RECT 116.015 175.445 117.175 175.685 ;
        RECT 117.355 175.665 117.625 176.395 ;
        RECT 117.805 175.845 118.145 176.575 ;
        RECT 117.355 175.445 118.125 175.665 ;
        RECT 116.005 174.935 116.305 175.265 ;
        RECT 116.485 174.955 117.010 175.265 ;
        RECT 117.190 174.955 117.655 175.265 ;
        RECT 111.445 174.025 111.775 174.425 ;
        RECT 112.825 174.255 113.155 174.595 ;
        RECT 113.325 174.025 113.655 174.425 ;
        RECT 114.155 174.025 115.825 174.795 ;
        RECT 116.015 174.025 116.305 174.755 ;
        RECT 116.485 174.315 116.715 174.955 ;
        RECT 117.835 174.775 118.125 175.445 ;
        RECT 116.895 174.575 118.125 174.775 ;
        RECT 116.895 174.205 117.205 174.575 ;
        RECT 117.385 174.025 118.055 174.395 ;
        RECT 118.315 174.205 118.575 176.395 ;
        RECT 118.790 175.785 119.325 176.405 ;
        RECT 118.790 174.765 119.105 175.785 ;
        RECT 119.495 175.775 119.825 176.575 ;
        RECT 121.055 176.140 126.400 176.575 ;
        RECT 120.310 175.605 120.700 175.780 ;
        RECT 119.275 175.435 120.700 175.605 ;
        RECT 119.275 174.935 119.445 175.435 ;
        RECT 118.790 174.195 119.405 174.765 ;
        RECT 119.695 174.705 119.960 175.265 ;
        RECT 120.130 174.535 120.300 175.435 ;
        RECT 120.470 174.705 120.825 175.265 ;
        RECT 122.640 174.570 122.980 175.400 ;
        RECT 124.460 174.890 124.810 176.140 ;
        RECT 127.585 175.645 127.755 176.405 ;
        RECT 127.970 175.815 128.300 176.575 ;
        RECT 127.585 175.475 128.300 175.645 ;
        RECT 128.470 175.500 128.725 176.405 ;
        RECT 127.495 174.925 127.850 175.295 ;
        RECT 128.130 175.265 128.300 175.475 ;
        RECT 128.130 174.935 128.385 175.265 ;
        RECT 128.130 174.745 128.300 174.935 ;
        RECT 128.555 174.770 128.725 175.500 ;
        RECT 128.900 175.425 129.160 176.575 ;
        RECT 129.335 175.410 129.625 176.575 ;
        RECT 129.800 175.435 130.135 176.405 ;
        RECT 130.305 175.435 130.475 176.575 ;
        RECT 130.645 176.235 132.675 176.405 ;
        RECT 127.585 174.575 128.300 174.745 ;
        RECT 119.575 174.025 119.790 174.535 ;
        RECT 120.020 174.205 120.300 174.535 ;
        RECT 120.480 174.025 120.720 174.535 ;
        RECT 121.055 174.025 126.400 174.570 ;
        RECT 127.585 174.195 127.755 174.575 ;
        RECT 127.970 174.025 128.300 174.405 ;
        RECT 128.470 174.195 128.725 174.770 ;
        RECT 128.900 174.025 129.160 174.865 ;
        RECT 129.800 174.765 129.970 175.435 ;
        RECT 130.645 175.265 130.815 176.235 ;
        RECT 130.140 174.935 130.395 175.265 ;
        RECT 130.620 174.935 130.815 175.265 ;
        RECT 130.985 175.895 132.110 176.065 ;
        RECT 130.225 174.765 130.395 174.935 ;
        RECT 130.985 174.765 131.155 175.895 ;
        RECT 129.335 174.025 129.625 174.750 ;
        RECT 129.800 174.195 130.055 174.765 ;
        RECT 130.225 174.595 131.155 174.765 ;
        RECT 131.325 175.555 132.335 175.725 ;
        RECT 131.325 174.755 131.495 175.555 ;
        RECT 131.700 174.875 131.975 175.355 ;
        RECT 131.695 174.705 131.975 174.875 ;
        RECT 130.980 174.560 131.155 174.595 ;
        RECT 130.225 174.025 130.555 174.425 ;
        RECT 130.980 174.195 131.510 174.560 ;
        RECT 131.700 174.195 131.975 174.705 ;
        RECT 132.145 174.195 132.335 175.555 ;
        RECT 132.505 175.570 132.675 176.235 ;
        RECT 132.845 175.815 133.015 176.575 ;
        RECT 133.250 175.815 133.765 176.225 ;
        RECT 132.505 175.380 133.255 175.570 ;
        RECT 133.425 175.005 133.765 175.815 ;
        RECT 132.535 174.835 133.765 175.005 ;
        RECT 133.935 175.435 134.320 176.405 ;
        RECT 134.490 176.115 134.815 176.575 ;
        RECT 135.335 175.945 135.615 176.405 ;
        RECT 134.490 175.725 135.615 175.945 ;
        RECT 132.515 174.025 133.025 174.560 ;
        RECT 133.245 174.230 133.490 174.835 ;
        RECT 133.935 174.765 134.215 175.435 ;
        RECT 134.490 175.265 134.940 175.725 ;
        RECT 135.805 175.555 136.205 176.405 ;
        RECT 136.605 176.115 136.875 176.575 ;
        RECT 137.045 175.945 137.330 176.405 ;
        RECT 134.385 174.935 134.940 175.265 ;
        RECT 135.110 174.995 136.205 175.555 ;
        RECT 134.490 174.825 134.940 174.935 ;
        RECT 133.935 174.195 134.320 174.765 ;
        RECT 134.490 174.655 135.615 174.825 ;
        RECT 134.490 174.025 134.815 174.485 ;
        RECT 135.335 174.195 135.615 174.655 ;
        RECT 135.805 174.195 136.205 174.995 ;
        RECT 136.375 175.725 137.330 175.945 ;
        RECT 136.375 174.825 136.585 175.725 ;
        RECT 136.755 174.995 137.445 175.555 ;
        RECT 137.615 175.485 138.825 176.575 ;
        RECT 137.615 174.945 138.135 175.485 ;
        RECT 136.375 174.655 137.330 174.825 ;
        RECT 138.305 174.775 138.825 175.315 ;
        RECT 136.605 174.025 136.875 174.485 ;
        RECT 137.045 174.195 137.330 174.655 ;
        RECT 137.615 174.025 138.825 174.775 ;
        RECT 13.330 173.855 138.910 174.025 ;
        RECT 13.415 173.105 14.625 173.855 ;
        RECT 13.415 172.565 13.935 173.105 ;
        RECT 14.795 173.085 17.385 173.855 ;
        RECT 18.065 173.465 18.395 173.855 ;
        RECT 18.565 173.285 18.735 173.605 ;
        RECT 18.905 173.465 19.235 173.855 ;
        RECT 19.650 173.455 20.605 173.625 ;
        RECT 18.015 173.115 20.265 173.285 ;
        RECT 14.105 172.395 14.625 172.935 ;
        RECT 14.795 172.565 16.005 173.085 ;
        RECT 16.175 172.395 17.385 172.915 ;
        RECT 13.415 171.305 14.625 172.395 ;
        RECT 14.795 171.305 17.385 172.395 ;
        RECT 18.015 172.155 18.185 173.115 ;
        RECT 18.355 172.495 18.600 172.945 ;
        RECT 18.770 172.665 19.320 172.865 ;
        RECT 19.490 172.695 19.865 172.865 ;
        RECT 19.490 172.495 19.660 172.695 ;
        RECT 20.035 172.615 20.265 173.115 ;
        RECT 18.355 172.325 19.660 172.495 ;
        RECT 20.435 172.575 20.605 173.455 ;
        RECT 20.775 173.020 21.065 173.855 ;
        RECT 21.240 173.455 21.575 173.855 ;
        RECT 21.745 173.285 21.950 173.685 ;
        RECT 22.160 173.375 22.435 173.855 ;
        RECT 22.645 173.355 22.905 173.685 ;
        RECT 21.265 173.115 21.950 173.285 ;
        RECT 20.435 172.405 21.065 172.575 ;
        RECT 18.015 171.475 18.395 172.155 ;
        RECT 18.985 171.305 19.155 172.155 ;
        RECT 19.325 171.985 20.565 172.155 ;
        RECT 19.325 171.475 19.655 171.985 ;
        RECT 19.825 171.305 19.995 171.815 ;
        RECT 20.165 171.475 20.565 171.985 ;
        RECT 20.745 171.475 21.065 172.405 ;
        RECT 21.265 172.085 21.605 173.115 ;
        RECT 21.775 172.445 22.025 172.945 ;
        RECT 22.205 172.615 22.565 173.195 ;
        RECT 22.735 172.445 22.905 173.355 ;
        RECT 23.075 173.085 25.665 173.855 ;
        RECT 25.835 173.115 26.300 173.660 ;
        RECT 23.075 172.565 24.285 173.085 ;
        RECT 21.775 172.275 22.905 172.445 ;
        RECT 24.455 172.395 25.665 172.915 ;
        RECT 21.265 171.910 21.930 172.085 ;
        RECT 21.240 171.305 21.575 171.730 ;
        RECT 21.745 171.505 21.930 171.910 ;
        RECT 22.135 171.305 22.465 172.085 ;
        RECT 22.635 171.505 22.905 172.275 ;
        RECT 23.075 171.305 25.665 172.395 ;
        RECT 25.835 172.155 26.005 173.115 ;
        RECT 26.805 173.035 26.975 173.855 ;
        RECT 27.145 173.205 27.475 173.685 ;
        RECT 27.645 173.465 27.995 173.855 ;
        RECT 28.165 173.285 28.395 173.685 ;
        RECT 27.885 173.205 28.395 173.285 ;
        RECT 27.145 173.115 28.395 173.205 ;
        RECT 28.565 173.115 28.885 173.595 ;
        RECT 27.145 173.035 28.055 173.115 ;
        RECT 26.175 172.495 26.420 172.945 ;
        RECT 26.680 172.665 27.375 172.865 ;
        RECT 27.545 172.695 28.145 172.865 ;
        RECT 27.545 172.495 27.715 172.695 ;
        RECT 28.375 172.525 28.545 172.945 ;
        RECT 26.175 172.325 27.715 172.495 ;
        RECT 27.885 172.355 28.545 172.525 ;
        RECT 27.885 172.155 28.055 172.355 ;
        RECT 28.715 172.185 28.885 173.115 ;
        RECT 25.835 171.985 28.055 172.155 ;
        RECT 28.225 171.985 28.885 172.185 ;
        RECT 29.055 173.115 29.520 173.660 ;
        RECT 29.055 172.155 29.225 173.115 ;
        RECT 30.025 173.035 30.195 173.855 ;
        RECT 30.365 173.205 30.695 173.685 ;
        RECT 30.865 173.465 31.215 173.855 ;
        RECT 31.385 173.285 31.615 173.685 ;
        RECT 31.105 173.205 31.615 173.285 ;
        RECT 30.365 173.115 31.615 173.205 ;
        RECT 31.785 173.115 32.105 173.595 ;
        RECT 30.365 173.035 31.275 173.115 ;
        RECT 29.395 172.495 29.640 172.945 ;
        RECT 29.900 172.665 30.595 172.865 ;
        RECT 30.765 172.695 31.365 172.865 ;
        RECT 30.765 172.495 30.935 172.695 ;
        RECT 31.595 172.525 31.765 172.945 ;
        RECT 29.395 172.325 30.935 172.495 ;
        RECT 31.105 172.355 31.765 172.525 ;
        RECT 31.105 172.155 31.275 172.355 ;
        RECT 31.935 172.185 32.105 173.115 ;
        RECT 32.275 173.085 34.865 173.855 ;
        RECT 35.510 173.285 35.765 173.635 ;
        RECT 35.935 173.455 36.265 173.855 ;
        RECT 36.435 173.285 36.605 173.635 ;
        RECT 36.775 173.455 37.155 173.855 ;
        RECT 35.510 173.115 37.175 173.285 ;
        RECT 37.345 173.180 37.620 173.525 ;
        RECT 32.275 172.565 33.485 173.085 ;
        RECT 37.005 172.945 37.175 173.115 ;
        RECT 33.655 172.395 34.865 172.915 ;
        RECT 35.495 172.615 35.840 172.945 ;
        RECT 36.010 172.615 36.835 172.945 ;
        RECT 37.005 172.615 37.280 172.945 ;
        RECT 29.055 171.985 31.275 172.155 ;
        RECT 31.445 171.985 32.105 172.185 ;
        RECT 25.835 171.305 26.135 171.815 ;
        RECT 26.305 171.475 26.635 171.985 ;
        RECT 28.225 171.815 28.395 171.985 ;
        RECT 26.805 171.305 27.435 171.815 ;
        RECT 28.015 171.645 28.395 171.815 ;
        RECT 28.565 171.305 28.865 171.815 ;
        RECT 29.055 171.305 29.355 171.815 ;
        RECT 29.525 171.475 29.855 171.985 ;
        RECT 31.445 171.815 31.615 171.985 ;
        RECT 30.025 171.305 30.655 171.815 ;
        RECT 31.235 171.645 31.615 171.815 ;
        RECT 31.785 171.305 32.085 171.815 ;
        RECT 32.275 171.305 34.865 172.395 ;
        RECT 35.515 172.155 35.840 172.445 ;
        RECT 36.010 172.325 36.205 172.615 ;
        RECT 37.005 172.445 37.175 172.615 ;
        RECT 37.450 172.445 37.620 173.180 ;
        RECT 37.795 173.105 39.005 173.855 ;
        RECT 39.175 173.130 39.465 173.855 ;
        RECT 39.725 173.205 39.895 173.685 ;
        RECT 40.065 173.375 40.395 173.855 ;
        RECT 40.620 173.435 42.155 173.685 ;
        RECT 40.620 173.205 40.790 173.435 ;
        RECT 37.795 172.565 38.315 173.105 ;
        RECT 39.725 173.035 40.790 173.205 ;
        RECT 36.515 172.275 37.175 172.445 ;
        RECT 36.515 172.155 36.685 172.275 ;
        RECT 35.515 171.985 36.685 172.155 ;
        RECT 35.495 171.525 36.685 171.815 ;
        RECT 36.855 171.305 37.135 172.105 ;
        RECT 37.345 171.475 37.620 172.445 ;
        RECT 38.485 172.395 39.005 172.935 ;
        RECT 40.970 172.865 41.250 173.265 ;
        RECT 39.640 172.655 39.990 172.865 ;
        RECT 40.160 172.665 40.605 172.865 ;
        RECT 40.775 172.665 41.250 172.865 ;
        RECT 41.520 172.865 41.805 173.265 ;
        RECT 41.985 173.205 42.155 173.435 ;
        RECT 42.325 173.375 42.655 173.855 ;
        RECT 42.870 173.355 43.125 173.685 ;
        RECT 42.940 173.275 43.125 173.355 ;
        RECT 43.315 173.310 48.660 173.855 ;
        RECT 48.885 173.465 49.215 173.855 ;
        RECT 41.985 173.035 42.785 173.205 ;
        RECT 41.520 172.665 41.850 172.865 ;
        RECT 42.020 172.835 42.385 172.865 ;
        RECT 42.020 172.665 42.395 172.835 ;
        RECT 42.615 172.485 42.785 173.035 ;
        RECT 37.795 171.305 39.005 172.395 ;
        RECT 39.175 171.305 39.465 172.470 ;
        RECT 39.725 172.315 42.785 172.485 ;
        RECT 39.725 171.475 39.895 172.315 ;
        RECT 42.955 172.145 43.125 173.275 ;
        RECT 44.900 172.480 45.240 173.310 ;
        RECT 49.385 173.285 49.555 173.605 ;
        RECT 49.725 173.465 50.055 173.855 ;
        RECT 50.470 173.455 51.425 173.625 ;
        RECT 48.835 173.115 51.085 173.285 ;
        RECT 40.065 171.645 40.395 172.145 ;
        RECT 40.565 171.905 42.200 172.145 ;
        RECT 40.565 171.815 40.795 171.905 ;
        RECT 40.905 171.645 41.235 171.685 ;
        RECT 40.065 171.475 41.235 171.645 ;
        RECT 41.425 171.305 41.780 171.725 ;
        RECT 41.950 171.475 42.200 171.905 ;
        RECT 42.370 171.305 42.700 172.065 ;
        RECT 42.870 171.475 43.125 172.145 ;
        RECT 46.720 171.740 47.070 172.990 ;
        RECT 48.835 172.155 49.005 173.115 ;
        RECT 49.175 172.495 49.420 172.945 ;
        RECT 49.590 172.665 50.140 172.865 ;
        RECT 50.310 172.695 50.685 172.865 ;
        RECT 50.310 172.495 50.480 172.695 ;
        RECT 50.855 172.615 51.085 173.115 ;
        RECT 49.175 172.325 50.480 172.495 ;
        RECT 51.255 172.575 51.425 173.455 ;
        RECT 51.595 173.020 51.885 173.855 ;
        RECT 52.060 173.455 52.395 173.855 ;
        RECT 52.565 173.285 52.770 173.685 ;
        RECT 52.980 173.375 53.255 173.855 ;
        RECT 53.465 173.355 53.725 173.685 ;
        RECT 52.085 173.115 52.770 173.285 ;
        RECT 51.255 172.405 51.885 172.575 ;
        RECT 43.315 171.305 48.660 171.740 ;
        RECT 48.835 171.475 49.215 172.155 ;
        RECT 49.805 171.305 49.975 172.155 ;
        RECT 50.145 171.985 51.385 172.155 ;
        RECT 50.145 171.475 50.475 171.985 ;
        RECT 50.645 171.305 50.815 171.815 ;
        RECT 50.985 171.475 51.385 171.985 ;
        RECT 51.565 171.475 51.885 172.405 ;
        RECT 52.085 172.085 52.425 173.115 ;
        RECT 52.595 172.445 52.845 172.945 ;
        RECT 53.025 172.615 53.385 173.195 ;
        RECT 53.555 172.445 53.725 173.355 ;
        RECT 53.895 173.310 59.240 173.855 ;
        RECT 55.480 172.480 55.820 173.310 ;
        RECT 59.415 173.085 61.085 173.855 ;
        RECT 61.260 173.325 61.550 173.675 ;
        RECT 61.745 173.495 62.075 173.855 ;
        RECT 62.245 173.325 62.475 173.630 ;
        RECT 61.260 173.155 62.475 173.325 ;
        RECT 62.665 173.175 62.835 173.550 ;
        RECT 52.595 172.275 53.725 172.445 ;
        RECT 52.085 171.910 52.750 172.085 ;
        RECT 52.060 171.305 52.395 171.730 ;
        RECT 52.565 171.505 52.750 171.910 ;
        RECT 52.955 171.305 53.285 172.085 ;
        RECT 53.455 171.505 53.725 172.275 ;
        RECT 57.300 171.740 57.650 172.990 ;
        RECT 59.415 172.565 60.165 173.085 ;
        RECT 62.665 173.005 62.865 173.175 ;
        RECT 63.095 173.085 64.765 173.855 ;
        RECT 64.935 173.130 65.225 173.855 ;
        RECT 65.485 173.305 65.655 173.595 ;
        RECT 65.825 173.475 66.155 173.855 ;
        RECT 65.485 173.135 66.150 173.305 ;
        RECT 62.665 172.985 62.835 173.005 ;
        RECT 60.335 172.395 61.085 172.915 ;
        RECT 61.320 172.835 61.580 172.945 ;
        RECT 61.315 172.665 61.580 172.835 ;
        RECT 61.320 172.615 61.580 172.665 ;
        RECT 61.760 172.615 62.145 172.945 ;
        RECT 62.315 172.815 62.835 172.985 ;
        RECT 53.895 171.305 59.240 171.740 ;
        RECT 59.415 171.305 61.085 172.395 ;
        RECT 61.260 171.305 61.580 172.445 ;
        RECT 61.760 171.565 61.955 172.615 ;
        RECT 62.315 172.435 62.485 172.815 ;
        RECT 62.135 172.155 62.485 172.435 ;
        RECT 62.675 172.285 62.920 172.645 ;
        RECT 63.095 172.565 63.845 173.085 ;
        RECT 64.015 172.395 64.765 172.915 ;
        RECT 62.135 171.475 62.465 172.155 ;
        RECT 62.665 171.305 62.920 172.105 ;
        RECT 63.095 171.305 64.765 172.395 ;
        RECT 64.935 171.305 65.225 172.470 ;
        RECT 65.400 172.315 65.750 172.965 ;
        RECT 65.920 172.145 66.150 173.135 ;
        RECT 65.485 171.975 66.150 172.145 ;
        RECT 65.485 171.475 65.655 171.975 ;
        RECT 65.825 171.305 66.155 171.805 ;
        RECT 66.325 171.475 66.510 173.595 ;
        RECT 66.765 173.395 67.015 173.855 ;
        RECT 67.185 173.405 67.520 173.575 ;
        RECT 67.715 173.405 68.390 173.575 ;
        RECT 67.185 173.265 67.355 173.405 ;
        RECT 66.680 172.275 66.960 173.225 ;
        RECT 67.130 173.135 67.355 173.265 ;
        RECT 67.130 172.030 67.300 173.135 ;
        RECT 67.525 172.985 68.050 173.205 ;
        RECT 67.470 172.220 67.710 172.815 ;
        RECT 67.880 172.285 68.050 172.985 ;
        RECT 68.220 172.625 68.390 173.405 ;
        RECT 68.710 173.355 69.080 173.855 ;
        RECT 69.260 173.405 69.665 173.575 ;
        RECT 69.835 173.405 70.620 173.575 ;
        RECT 69.260 173.175 69.430 173.405 ;
        RECT 68.600 172.875 69.430 173.175 ;
        RECT 69.815 172.905 70.280 173.235 ;
        RECT 68.600 172.845 68.800 172.875 ;
        RECT 68.920 172.625 69.090 172.695 ;
        RECT 68.220 172.455 69.090 172.625 ;
        RECT 68.580 172.365 69.090 172.455 ;
        RECT 67.130 171.900 67.435 172.030 ;
        RECT 67.880 171.920 68.410 172.285 ;
        RECT 66.750 171.305 67.015 171.765 ;
        RECT 67.185 171.475 67.435 171.900 ;
        RECT 68.580 171.750 68.750 172.365 ;
        RECT 67.645 171.580 68.750 171.750 ;
        RECT 68.920 171.305 69.090 172.105 ;
        RECT 69.260 171.805 69.430 172.875 ;
        RECT 69.600 171.975 69.790 172.695 ;
        RECT 69.960 171.945 70.280 172.905 ;
        RECT 70.450 172.945 70.620 173.405 ;
        RECT 70.895 173.325 71.105 173.855 ;
        RECT 71.365 173.115 71.695 173.640 ;
        RECT 71.865 173.245 72.035 173.855 ;
        RECT 72.205 173.200 72.535 173.635 ;
        RECT 72.205 173.115 72.585 173.200 ;
        RECT 71.495 172.945 71.695 173.115 ;
        RECT 72.360 173.075 72.585 173.115 ;
        RECT 70.450 172.615 71.325 172.945 ;
        RECT 71.495 172.615 72.245 172.945 ;
        RECT 69.260 171.475 69.510 171.805 ;
        RECT 70.450 171.775 70.620 172.615 ;
        RECT 71.495 172.410 71.685 172.615 ;
        RECT 72.415 172.495 72.585 173.075 ;
        RECT 72.755 173.105 73.965 173.855 ;
        RECT 74.250 173.225 74.535 173.685 ;
        RECT 74.705 173.395 74.975 173.855 ;
        RECT 72.755 172.565 73.275 173.105 ;
        RECT 74.250 173.055 75.205 173.225 ;
        RECT 72.370 172.445 72.585 172.495 ;
        RECT 70.790 172.035 71.685 172.410 ;
        RECT 72.195 172.365 72.585 172.445 ;
        RECT 73.445 172.395 73.965 172.935 ;
        RECT 69.735 171.605 70.620 171.775 ;
        RECT 70.800 171.305 71.115 171.805 ;
        RECT 71.345 171.475 71.685 172.035 ;
        RECT 71.855 171.305 72.025 172.315 ;
        RECT 72.195 171.520 72.525 172.365 ;
        RECT 72.755 171.305 73.965 172.395 ;
        RECT 74.135 172.325 74.825 172.885 ;
        RECT 74.995 172.155 75.205 173.055 ;
        RECT 74.250 171.935 75.205 172.155 ;
        RECT 75.375 172.885 75.775 173.685 ;
        RECT 75.965 173.225 76.245 173.685 ;
        RECT 76.765 173.395 77.090 173.855 ;
        RECT 75.965 173.055 77.090 173.225 ;
        RECT 77.260 173.115 77.645 173.685 ;
        RECT 76.640 172.945 77.090 173.055 ;
        RECT 75.375 172.325 76.470 172.885 ;
        RECT 76.640 172.615 77.195 172.945 ;
        RECT 74.250 171.475 74.535 171.935 ;
        RECT 74.705 171.305 74.975 171.765 ;
        RECT 75.375 171.475 75.775 172.325 ;
        RECT 76.640 172.155 77.090 172.615 ;
        RECT 77.365 172.445 77.645 173.115 ;
        RECT 75.965 171.935 77.090 172.155 ;
        RECT 75.965 171.475 76.245 171.935 ;
        RECT 76.765 171.305 77.090 171.765 ;
        RECT 77.260 171.475 77.645 172.445 ;
        RECT 77.820 173.115 78.075 173.685 ;
        RECT 78.245 173.455 78.575 173.855 ;
        RECT 79.000 173.320 79.530 173.685 ;
        RECT 79.720 173.515 79.995 173.685 ;
        RECT 79.715 173.345 79.995 173.515 ;
        RECT 79.000 173.285 79.175 173.320 ;
        RECT 78.245 173.115 79.175 173.285 ;
        RECT 77.820 172.445 77.990 173.115 ;
        RECT 78.245 172.945 78.415 173.115 ;
        RECT 78.160 172.615 78.415 172.945 ;
        RECT 78.640 172.615 78.835 172.945 ;
        RECT 77.820 171.475 78.155 172.445 ;
        RECT 78.325 171.305 78.495 172.445 ;
        RECT 78.665 171.645 78.835 172.615 ;
        RECT 79.005 171.985 79.175 173.115 ;
        RECT 79.345 172.325 79.515 173.125 ;
        RECT 79.720 172.525 79.995 173.345 ;
        RECT 80.165 172.325 80.355 173.685 ;
        RECT 80.535 173.320 81.045 173.855 ;
        RECT 81.265 173.045 81.510 173.650 ;
        RECT 81.960 173.115 82.215 173.685 ;
        RECT 82.385 173.455 82.715 173.855 ;
        RECT 83.140 173.320 83.670 173.685 ;
        RECT 83.140 173.285 83.315 173.320 ;
        RECT 82.385 173.115 83.315 173.285 ;
        RECT 80.555 172.875 81.785 173.045 ;
        RECT 79.345 172.155 80.355 172.325 ;
        RECT 80.525 172.310 81.275 172.500 ;
        RECT 79.005 171.815 80.130 171.985 ;
        RECT 80.525 171.645 80.695 172.310 ;
        RECT 81.445 172.065 81.785 172.875 ;
        RECT 78.665 171.475 80.695 171.645 ;
        RECT 80.865 171.305 81.035 172.065 ;
        RECT 81.270 171.655 81.785 172.065 ;
        RECT 81.960 172.445 82.130 173.115 ;
        RECT 82.385 172.945 82.555 173.115 ;
        RECT 82.300 172.615 82.555 172.945 ;
        RECT 82.780 172.615 82.975 172.945 ;
        RECT 81.960 171.475 82.295 172.445 ;
        RECT 82.465 171.305 82.635 172.445 ;
        RECT 82.805 171.645 82.975 172.615 ;
        RECT 83.145 171.985 83.315 173.115 ;
        RECT 83.485 172.325 83.655 173.125 ;
        RECT 83.860 172.835 84.135 173.685 ;
        RECT 83.855 172.665 84.135 172.835 ;
        RECT 83.860 172.525 84.135 172.665 ;
        RECT 84.305 172.325 84.495 173.685 ;
        RECT 84.675 173.320 85.185 173.855 ;
        RECT 85.405 173.045 85.650 173.650 ;
        RECT 86.095 173.085 89.605 173.855 ;
        RECT 90.695 173.130 90.985 173.855 ;
        RECT 91.155 173.085 93.745 173.855 ;
        RECT 93.975 173.395 94.220 173.855 ;
        RECT 84.695 172.875 85.925 173.045 ;
        RECT 83.485 172.155 84.495 172.325 ;
        RECT 84.665 172.310 85.415 172.500 ;
        RECT 83.145 171.815 84.270 171.985 ;
        RECT 84.665 171.645 84.835 172.310 ;
        RECT 85.585 172.065 85.925 172.875 ;
        RECT 86.095 172.565 87.745 173.085 ;
        RECT 87.915 172.395 89.605 172.915 ;
        RECT 91.155 172.565 92.365 173.085 ;
        RECT 82.805 171.475 84.835 171.645 ;
        RECT 85.005 171.305 85.175 172.065 ;
        RECT 85.410 171.655 85.925 172.065 ;
        RECT 86.095 171.305 89.605 172.395 ;
        RECT 90.695 171.305 90.985 172.470 ;
        RECT 92.535 172.395 93.745 172.915 ;
        RECT 93.915 172.615 94.230 173.225 ;
        RECT 94.400 172.865 94.650 173.675 ;
        RECT 94.820 173.330 95.080 173.855 ;
        RECT 95.250 173.205 95.510 173.660 ;
        RECT 95.680 173.375 95.940 173.855 ;
        RECT 96.110 173.205 96.370 173.660 ;
        RECT 96.540 173.375 96.800 173.855 ;
        RECT 96.970 173.205 97.230 173.660 ;
        RECT 97.400 173.375 97.660 173.855 ;
        RECT 97.830 173.205 98.090 173.660 ;
        RECT 98.260 173.375 98.560 173.855 ;
        RECT 95.250 173.035 98.560 173.205 ;
        RECT 94.400 172.615 97.420 172.865 ;
        RECT 91.155 171.305 93.745 172.395 ;
        RECT 93.925 171.305 94.220 172.415 ;
        RECT 94.400 171.480 94.650 172.615 ;
        RECT 97.590 172.445 98.560 173.035 ;
        RECT 98.975 173.085 101.565 173.855 ;
        RECT 98.975 172.565 100.185 173.085 ;
        RECT 102.195 173.055 102.505 173.855 ;
        RECT 102.710 173.055 103.405 173.685 ;
        RECT 103.575 173.310 108.920 173.855 ;
        RECT 94.820 171.305 95.080 172.415 ;
        RECT 95.250 172.205 98.560 172.445 ;
        RECT 100.355 172.395 101.565 172.915 ;
        RECT 102.205 172.615 102.540 172.885 ;
        RECT 102.710 172.455 102.880 173.055 ;
        RECT 103.050 172.615 103.385 172.865 ;
        RECT 105.160 172.480 105.500 173.310 ;
        RECT 109.095 173.085 112.605 173.855 ;
        RECT 113.235 173.205 113.495 173.685 ;
        RECT 113.665 173.315 113.915 173.855 ;
        RECT 95.250 171.480 95.510 172.205 ;
        RECT 95.680 171.305 95.940 172.035 ;
        RECT 96.110 171.480 96.370 172.205 ;
        RECT 96.540 171.305 96.800 172.035 ;
        RECT 96.970 171.480 97.230 172.205 ;
        RECT 97.400 171.305 97.660 172.035 ;
        RECT 97.830 171.480 98.090 172.205 ;
        RECT 98.260 171.305 98.555 172.035 ;
        RECT 98.975 171.305 101.565 172.395 ;
        RECT 102.195 171.305 102.475 172.445 ;
        RECT 102.645 171.475 102.975 172.455 ;
        RECT 103.145 171.305 103.405 172.445 ;
        RECT 106.980 171.740 107.330 172.990 ;
        RECT 109.095 172.565 110.745 173.085 ;
        RECT 110.915 172.395 112.605 172.915 ;
        RECT 103.575 171.305 108.920 171.740 ;
        RECT 109.095 171.305 112.605 172.395 ;
        RECT 113.235 172.175 113.405 173.205 ;
        RECT 114.085 173.150 114.305 173.635 ;
        RECT 113.575 172.555 113.805 172.950 ;
        RECT 113.975 172.725 114.305 173.150 ;
        RECT 114.475 173.475 115.365 173.645 ;
        RECT 114.475 172.750 114.645 173.475 ;
        RECT 114.815 172.920 115.365 173.305 ;
        RECT 116.455 173.130 116.745 173.855 ;
        RECT 117.120 173.075 117.620 173.685 ;
        RECT 114.475 172.680 115.365 172.750 ;
        RECT 114.470 172.655 115.365 172.680 ;
        RECT 114.460 172.640 115.365 172.655 ;
        RECT 114.455 172.625 115.365 172.640 ;
        RECT 114.445 172.620 115.365 172.625 ;
        RECT 114.440 172.610 115.365 172.620 ;
        RECT 116.915 172.615 117.265 172.865 ;
        RECT 114.435 172.600 115.365 172.610 ;
        RECT 114.425 172.595 115.365 172.600 ;
        RECT 114.415 172.585 115.365 172.595 ;
        RECT 114.405 172.580 115.365 172.585 ;
        RECT 114.405 172.575 114.740 172.580 ;
        RECT 114.390 172.570 114.740 172.575 ;
        RECT 114.375 172.560 114.740 172.570 ;
        RECT 114.350 172.555 114.740 172.560 ;
        RECT 113.575 172.550 114.740 172.555 ;
        RECT 113.575 172.515 114.710 172.550 ;
        RECT 113.575 172.490 114.675 172.515 ;
        RECT 113.575 172.460 114.645 172.490 ;
        RECT 113.575 172.430 114.625 172.460 ;
        RECT 113.575 172.400 114.605 172.430 ;
        RECT 113.575 172.390 114.535 172.400 ;
        RECT 113.575 172.380 114.510 172.390 ;
        RECT 113.575 172.365 114.490 172.380 ;
        RECT 113.575 172.350 114.470 172.365 ;
        RECT 113.680 172.340 114.465 172.350 ;
        RECT 113.680 172.305 114.450 172.340 ;
        RECT 113.235 171.475 113.510 172.175 ;
        RECT 113.680 172.055 114.435 172.305 ;
        RECT 114.605 171.985 114.935 172.230 ;
        RECT 115.105 172.130 115.365 172.580 ;
        RECT 114.750 171.960 114.935 171.985 ;
        RECT 114.750 171.860 115.365 171.960 ;
        RECT 113.680 171.305 113.935 171.850 ;
        RECT 114.105 171.475 114.585 171.815 ;
        RECT 114.760 171.305 115.365 171.860 ;
        RECT 116.455 171.305 116.745 172.470 ;
        RECT 117.450 172.445 117.620 173.075 ;
        RECT 118.250 173.205 118.580 173.685 ;
        RECT 118.750 173.395 118.975 173.855 ;
        RECT 119.145 173.205 119.475 173.685 ;
        RECT 118.250 173.035 119.475 173.205 ;
        RECT 119.665 173.055 119.915 173.855 ;
        RECT 120.085 173.055 120.425 173.685 ;
        RECT 117.790 172.665 118.120 172.865 ;
        RECT 118.290 172.665 118.620 172.865 ;
        RECT 118.790 172.665 119.210 172.865 ;
        RECT 119.385 172.695 120.080 172.865 ;
        RECT 119.385 172.445 119.555 172.695 ;
        RECT 120.250 172.445 120.425 173.055 ;
        RECT 120.595 173.085 124.105 173.855 ;
        RECT 124.275 173.105 125.485 173.855 ;
        RECT 125.745 173.305 125.915 173.685 ;
        RECT 126.095 173.475 126.425 173.855 ;
        RECT 125.745 173.135 126.410 173.305 ;
        RECT 126.605 173.180 126.865 173.685 ;
        RECT 120.595 172.565 122.245 173.085 ;
        RECT 117.120 172.275 119.555 172.445 ;
        RECT 117.120 171.475 117.450 172.275 ;
        RECT 117.620 171.305 117.950 172.105 ;
        RECT 118.250 171.475 118.580 172.275 ;
        RECT 119.225 171.305 119.475 172.105 ;
        RECT 119.745 171.305 119.915 172.445 ;
        RECT 120.085 171.475 120.425 172.445 ;
        RECT 122.415 172.395 124.105 172.915 ;
        RECT 124.275 172.565 124.795 173.105 ;
        RECT 124.965 172.395 125.485 172.935 ;
        RECT 125.675 172.585 126.005 172.955 ;
        RECT 126.240 172.880 126.410 173.135 ;
        RECT 126.240 172.550 126.525 172.880 ;
        RECT 126.240 172.405 126.410 172.550 ;
        RECT 120.595 171.305 124.105 172.395 ;
        RECT 124.275 171.305 125.485 172.395 ;
        RECT 125.745 172.235 126.410 172.405 ;
        RECT 126.695 172.380 126.865 173.180 ;
        RECT 127.125 173.305 127.295 173.595 ;
        RECT 127.465 173.475 127.795 173.855 ;
        RECT 127.125 173.135 127.790 173.305 ;
        RECT 125.745 171.475 125.915 172.235 ;
        RECT 126.095 171.305 126.425 172.065 ;
        RECT 126.595 171.475 126.865 172.380 ;
        RECT 127.040 172.315 127.390 172.965 ;
        RECT 127.560 172.145 127.790 173.135 ;
        RECT 127.125 171.975 127.790 172.145 ;
        RECT 127.125 171.475 127.295 171.975 ;
        RECT 127.465 171.305 127.795 171.805 ;
        RECT 127.965 171.475 128.150 173.595 ;
        RECT 128.405 173.395 128.655 173.855 ;
        RECT 128.825 173.405 129.160 173.575 ;
        RECT 129.355 173.405 130.030 173.575 ;
        RECT 128.825 173.265 128.995 173.405 ;
        RECT 128.320 172.275 128.600 173.225 ;
        RECT 128.770 173.135 128.995 173.265 ;
        RECT 128.770 172.030 128.940 173.135 ;
        RECT 129.165 172.985 129.690 173.205 ;
        RECT 129.110 172.220 129.350 172.815 ;
        RECT 129.520 172.285 129.690 172.985 ;
        RECT 129.860 172.625 130.030 173.405 ;
        RECT 130.350 173.355 130.720 173.855 ;
        RECT 130.900 173.405 131.305 173.575 ;
        RECT 131.475 173.405 132.260 173.575 ;
        RECT 130.900 173.175 131.070 173.405 ;
        RECT 130.240 172.875 131.070 173.175 ;
        RECT 131.455 172.905 131.920 173.235 ;
        RECT 130.240 172.845 130.440 172.875 ;
        RECT 130.560 172.625 130.730 172.695 ;
        RECT 129.860 172.455 130.730 172.625 ;
        RECT 130.220 172.365 130.730 172.455 ;
        RECT 128.770 171.900 129.075 172.030 ;
        RECT 129.520 171.920 130.050 172.285 ;
        RECT 128.390 171.305 128.655 171.765 ;
        RECT 128.825 171.475 129.075 171.900 ;
        RECT 130.220 171.750 130.390 172.365 ;
        RECT 129.285 171.580 130.390 171.750 ;
        RECT 130.560 171.305 130.730 172.105 ;
        RECT 130.900 171.805 131.070 172.875 ;
        RECT 131.240 171.975 131.430 172.695 ;
        RECT 131.600 171.945 131.920 172.905 ;
        RECT 132.090 172.945 132.260 173.405 ;
        RECT 132.535 173.325 132.745 173.855 ;
        RECT 133.005 173.115 133.335 173.640 ;
        RECT 133.505 173.245 133.675 173.855 ;
        RECT 133.845 173.200 134.175 173.635 ;
        RECT 133.845 173.115 134.225 173.200 ;
        RECT 133.135 172.945 133.335 173.115 ;
        RECT 134.000 173.075 134.225 173.115 ;
        RECT 132.090 172.615 132.965 172.945 ;
        RECT 133.135 172.615 133.885 172.945 ;
        RECT 130.900 171.475 131.150 171.805 ;
        RECT 132.090 171.775 132.260 172.615 ;
        RECT 133.135 172.410 133.325 172.615 ;
        RECT 134.055 172.495 134.225 173.075 ;
        RECT 134.010 172.445 134.225 172.495 ;
        RECT 132.430 172.035 133.325 172.410 ;
        RECT 133.835 172.365 134.225 172.445 ;
        RECT 134.395 173.180 134.655 173.685 ;
        RECT 134.835 173.475 135.165 173.855 ;
        RECT 135.345 173.305 135.515 173.685 ;
        RECT 134.395 172.380 134.565 173.180 ;
        RECT 134.850 173.135 135.515 173.305 ;
        RECT 135.865 173.305 136.035 173.685 ;
        RECT 136.250 173.475 136.580 173.855 ;
        RECT 135.865 173.135 136.580 173.305 ;
        RECT 134.850 172.880 135.020 173.135 ;
        RECT 134.735 172.550 135.020 172.880 ;
        RECT 135.255 172.585 135.585 172.955 ;
        RECT 135.775 172.585 136.130 172.955 ;
        RECT 136.410 172.945 136.580 173.135 ;
        RECT 136.750 173.110 137.005 173.685 ;
        RECT 136.410 172.615 136.665 172.945 ;
        RECT 134.850 172.405 135.020 172.550 ;
        RECT 136.410 172.405 136.580 172.615 ;
        RECT 131.375 171.605 132.260 171.775 ;
        RECT 132.440 171.305 132.755 171.805 ;
        RECT 132.985 171.475 133.325 172.035 ;
        RECT 133.495 171.305 133.665 172.315 ;
        RECT 133.835 171.520 134.165 172.365 ;
        RECT 134.395 171.475 134.665 172.380 ;
        RECT 134.850 172.235 135.515 172.405 ;
        RECT 134.835 171.305 135.165 172.065 ;
        RECT 135.345 171.475 135.515 172.235 ;
        RECT 135.865 172.235 136.580 172.405 ;
        RECT 136.835 172.380 137.005 173.110 ;
        RECT 137.180 173.015 137.440 173.855 ;
        RECT 137.615 173.105 138.825 173.855 ;
        RECT 135.865 171.475 136.035 172.235 ;
        RECT 136.250 171.305 136.580 172.065 ;
        RECT 136.750 171.475 137.005 172.380 ;
        RECT 137.180 171.305 137.440 172.455 ;
        RECT 137.615 172.395 138.135 172.935 ;
        RECT 138.305 172.565 138.825 173.105 ;
        RECT 137.615 171.305 138.825 172.395 ;
        RECT 13.330 171.135 138.910 171.305 ;
        RECT 13.415 170.045 14.625 171.135 ;
        RECT 13.415 169.335 13.935 169.875 ;
        RECT 14.105 169.505 14.625 170.045 ;
        RECT 14.875 170.205 15.055 170.965 ;
        RECT 15.235 170.375 15.565 171.135 ;
        RECT 14.875 170.035 15.550 170.205 ;
        RECT 15.735 170.060 16.005 170.965 ;
        RECT 15.380 169.890 15.550 170.035 ;
        RECT 14.815 169.485 15.155 169.855 ;
        RECT 15.380 169.560 15.655 169.890 ;
        RECT 13.415 168.585 14.625 169.335 ;
        RECT 15.380 169.305 15.550 169.560 ;
        RECT 14.885 169.135 15.550 169.305 ;
        RECT 15.825 169.260 16.005 170.060 ;
        RECT 16.175 170.045 17.385 171.135 ;
        RECT 14.885 168.755 15.055 169.135 ;
        RECT 15.235 168.585 15.565 168.965 ;
        RECT 15.745 168.755 16.005 169.260 ;
        RECT 16.175 169.335 16.695 169.875 ;
        RECT 16.865 169.505 17.385 170.045 ;
        RECT 16.175 168.585 17.385 169.335 ;
        RECT 17.555 168.755 17.815 170.965 ;
        RECT 17.985 170.755 18.315 171.135 ;
        RECT 18.740 170.585 18.910 170.965 ;
        RECT 19.170 170.755 19.500 171.135 ;
        RECT 19.695 170.585 19.865 170.965 ;
        RECT 20.075 170.755 20.405 171.135 ;
        RECT 20.655 170.585 20.845 170.965 ;
        RECT 21.085 170.755 21.415 171.135 ;
        RECT 21.725 170.635 21.985 170.965 ;
        RECT 17.985 170.415 19.935 170.585 ;
        RECT 17.985 169.495 18.155 170.415 ;
        RECT 18.525 169.825 18.720 170.135 ;
        RECT 18.990 169.825 19.175 170.135 ;
        RECT 18.465 169.495 18.720 169.825 ;
        RECT 18.945 169.495 19.175 169.825 ;
        RECT 17.985 168.585 18.315 168.965 ;
        RECT 18.525 168.920 18.720 169.495 ;
        RECT 18.990 168.915 19.175 169.495 ;
        RECT 19.425 168.925 19.595 169.825 ;
        RECT 19.765 169.425 19.935 170.415 ;
        RECT 20.105 170.415 20.845 170.585 ;
        RECT 20.105 169.905 20.275 170.415 ;
        RECT 20.445 170.075 21.025 170.245 ;
        RECT 21.295 170.125 21.645 170.455 ;
        RECT 20.855 169.955 21.025 170.075 ;
        RECT 21.815 169.955 21.985 170.635 ;
        RECT 20.105 169.735 20.675 169.905 ;
        RECT 20.855 169.785 21.985 169.955 ;
        RECT 19.765 169.095 20.315 169.425 ;
        RECT 20.505 169.255 20.675 169.735 ;
        RECT 20.845 169.445 21.465 169.615 ;
        RECT 21.255 169.265 21.465 169.445 ;
        RECT 20.505 168.925 20.905 169.255 ;
        RECT 21.815 169.085 21.985 169.785 ;
        RECT 19.425 168.755 20.905 168.925 ;
        RECT 21.085 168.585 21.415 168.965 ;
        RECT 21.725 168.755 21.985 169.085 ;
        RECT 22.155 169.995 22.415 170.965 ;
        RECT 22.610 170.725 22.940 171.135 ;
        RECT 23.140 170.545 23.310 170.965 ;
        RECT 23.525 170.725 24.195 171.135 ;
        RECT 24.430 170.545 24.600 170.965 ;
        RECT 24.905 170.695 25.235 171.135 ;
        RECT 22.585 170.375 24.600 170.545 ;
        RECT 25.405 170.515 25.580 170.965 ;
        RECT 22.155 169.305 22.325 169.995 ;
        RECT 22.585 169.825 22.755 170.375 ;
        RECT 22.495 169.495 22.755 169.825 ;
        RECT 22.155 168.840 22.495 169.305 ;
        RECT 22.925 169.165 23.265 170.195 ;
        RECT 23.455 170.115 23.725 170.195 ;
        RECT 23.455 169.945 23.765 170.115 ;
        RECT 22.160 168.795 22.495 168.840 ;
        RECT 22.665 168.585 22.995 168.965 ;
        RECT 23.455 168.920 23.725 169.945 ;
        RECT 23.950 168.920 24.230 170.195 ;
        RECT 24.430 169.085 24.600 170.375 ;
        RECT 24.950 170.345 25.580 170.515 ;
        RECT 24.950 169.825 25.120 170.345 ;
        RECT 24.770 169.495 25.120 169.825 ;
        RECT 25.300 169.495 25.665 170.175 ;
        RECT 26.295 169.970 26.585 171.135 ;
        RECT 27.225 169.995 27.555 171.135 ;
        RECT 28.085 170.165 28.415 170.950 ;
        RECT 27.735 169.995 28.415 170.165 ;
        RECT 28.595 170.045 31.185 171.135 ;
        RECT 27.215 169.575 27.565 169.825 ;
        RECT 24.950 169.325 25.120 169.495 ;
        RECT 27.735 169.395 27.905 169.995 ;
        RECT 28.075 169.575 28.425 169.825 ;
        RECT 24.950 169.155 25.580 169.325 ;
        RECT 24.430 168.755 24.660 169.085 ;
        RECT 24.905 168.585 25.235 168.965 ;
        RECT 25.405 168.755 25.580 169.155 ;
        RECT 26.295 168.585 26.585 169.310 ;
        RECT 27.225 168.585 27.495 169.395 ;
        RECT 27.665 168.755 27.995 169.395 ;
        RECT 28.165 168.585 28.405 169.395 ;
        RECT 28.595 169.355 29.805 169.875 ;
        RECT 29.975 169.525 31.185 170.045 ;
        RECT 31.395 170.185 31.685 170.955 ;
        RECT 32.255 170.595 32.515 170.955 ;
        RECT 32.685 170.765 33.015 171.135 ;
        RECT 33.185 170.595 33.445 170.955 ;
        RECT 32.255 170.365 33.445 170.595 ;
        RECT 33.635 170.415 33.965 171.135 ;
        RECT 34.135 170.185 34.400 170.955 ;
        RECT 31.395 170.005 33.890 170.185 ;
        RECT 31.365 169.495 31.635 169.825 ;
        RECT 31.815 169.495 32.250 169.825 ;
        RECT 32.430 169.495 33.005 169.825 ;
        RECT 33.185 169.495 33.465 169.825 ;
        RECT 28.595 168.585 31.185 169.355 ;
        RECT 33.665 169.315 33.890 170.005 ;
        RECT 31.405 169.125 33.890 169.315 ;
        RECT 31.405 168.765 31.630 169.125 ;
        RECT 31.810 168.585 32.140 168.955 ;
        RECT 32.320 168.765 32.575 169.125 ;
        RECT 33.140 168.585 33.885 168.955 ;
        RECT 34.065 168.765 34.400 170.185 ;
        RECT 34.575 170.060 34.915 171.135 ;
        RECT 35.100 170.795 37.150 170.915 ;
        RECT 35.095 170.625 37.150 170.795 ;
        RECT 35.085 169.825 35.325 170.420 ;
        RECT 35.520 170.285 37.150 170.455 ;
        RECT 37.320 170.335 37.600 171.135 ;
        RECT 35.520 169.995 35.840 170.285 ;
        RECT 36.980 170.165 37.150 170.285 ;
        RECT 34.575 169.255 34.915 169.825 ;
        RECT 35.085 169.495 35.740 169.825 ;
        RECT 36.010 169.495 36.750 170.115 ;
        RECT 36.980 169.995 37.640 170.165 ;
        RECT 37.810 169.995 38.085 170.965 ;
        RECT 37.470 169.825 37.640 169.995 ;
        RECT 36.920 169.495 37.300 169.825 ;
        RECT 37.470 169.495 37.745 169.825 ;
        RECT 34.575 168.585 34.915 169.085 ;
        RECT 35.085 168.805 35.330 169.495 ;
        RECT 37.470 169.325 37.640 169.495 ;
        RECT 36.055 169.155 37.640 169.325 ;
        RECT 37.915 169.260 38.085 169.995 ;
        RECT 35.525 168.585 35.855 169.085 ;
        RECT 36.055 168.805 36.225 169.155 ;
        RECT 36.400 168.585 36.730 168.985 ;
        RECT 36.900 168.805 37.070 169.155 ;
        RECT 37.240 168.585 37.620 168.985 ;
        RECT 37.810 168.915 38.085 169.260 ;
        RECT 39.210 170.345 39.745 170.965 ;
        RECT 39.210 169.325 39.525 170.345 ;
        RECT 39.915 170.335 40.245 171.135 ;
        RECT 40.730 170.165 41.120 170.340 ;
        RECT 39.695 169.995 41.120 170.165 ;
        RECT 41.475 170.045 44.985 171.135 ;
        RECT 39.695 169.495 39.865 169.995 ;
        RECT 39.210 168.755 39.825 169.325 ;
        RECT 40.115 169.265 40.380 169.825 ;
        RECT 40.550 169.095 40.720 169.995 ;
        RECT 40.890 169.265 41.245 169.825 ;
        RECT 41.475 169.355 43.125 169.875 ;
        RECT 43.295 169.525 44.985 170.045 ;
        RECT 39.995 168.585 40.210 169.095 ;
        RECT 40.440 168.765 40.720 169.095 ;
        RECT 40.900 168.585 41.140 169.095 ;
        RECT 41.475 168.585 44.985 169.355 ;
        RECT 45.625 168.765 45.885 170.955 ;
        RECT 46.055 170.405 46.395 171.135 ;
        RECT 46.575 170.225 46.845 170.955 ;
        RECT 46.075 170.005 46.845 170.225 ;
        RECT 47.025 170.245 47.255 170.955 ;
        RECT 47.425 170.425 47.755 171.135 ;
        RECT 47.925 170.245 48.185 170.955 ;
        RECT 49.135 170.495 49.465 170.925 ;
        RECT 47.025 170.005 48.185 170.245 ;
        RECT 49.010 170.325 49.465 170.495 ;
        RECT 49.645 170.495 49.895 170.915 ;
        RECT 50.125 170.665 50.455 171.135 ;
        RECT 50.685 170.495 50.935 170.915 ;
        RECT 49.645 170.325 50.935 170.495 ;
        RECT 46.075 169.335 46.365 170.005 ;
        RECT 46.545 169.515 47.010 169.825 ;
        RECT 47.190 169.515 47.715 169.825 ;
        RECT 46.075 169.135 47.305 169.335 ;
        RECT 46.145 168.585 46.815 168.955 ;
        RECT 46.995 168.765 47.305 169.135 ;
        RECT 47.485 168.875 47.715 169.515 ;
        RECT 47.895 169.495 48.195 169.825 ;
        RECT 49.010 169.325 49.180 170.325 ;
        RECT 49.350 169.495 49.595 170.155 ;
        RECT 49.810 169.495 50.075 170.155 ;
        RECT 50.270 169.495 50.555 170.155 ;
        RECT 50.730 169.825 50.945 170.155 ;
        RECT 51.125 169.995 51.375 171.135 ;
        RECT 51.545 170.075 51.875 170.925 ;
        RECT 50.730 169.495 51.035 169.825 ;
        RECT 51.205 169.495 51.515 169.825 ;
        RECT 51.205 169.325 51.375 169.495 ;
        RECT 47.895 168.585 48.185 169.315 ;
        RECT 49.010 169.155 51.375 169.325 ;
        RECT 51.685 169.310 51.875 170.075 ;
        RECT 52.055 169.970 52.345 171.135 ;
        RECT 52.575 170.075 52.905 170.920 ;
        RECT 53.075 170.125 53.245 171.135 ;
        RECT 53.415 170.405 53.755 170.965 ;
        RECT 53.985 170.635 54.300 171.135 ;
        RECT 54.480 170.665 55.365 170.835 ;
        RECT 52.515 169.995 52.905 170.075 ;
        RECT 53.415 170.030 54.310 170.405 ;
        RECT 52.515 169.945 52.730 169.995 ;
        RECT 52.515 169.365 52.685 169.945 ;
        RECT 53.415 169.825 53.605 170.030 ;
        RECT 54.480 169.825 54.650 170.665 ;
        RECT 55.590 170.635 55.840 170.965 ;
        RECT 52.855 169.495 53.605 169.825 ;
        RECT 53.775 169.495 54.650 169.825 ;
        RECT 52.515 169.325 52.740 169.365 ;
        RECT 53.405 169.325 53.605 169.495 ;
        RECT 49.165 168.585 49.495 168.985 ;
        RECT 49.665 168.815 49.995 169.155 ;
        RECT 51.045 168.585 51.375 168.985 ;
        RECT 51.545 168.800 51.875 169.310 ;
        RECT 52.055 168.585 52.345 169.310 ;
        RECT 52.515 169.240 52.895 169.325 ;
        RECT 52.565 168.805 52.895 169.240 ;
        RECT 53.065 168.585 53.235 169.195 ;
        RECT 53.405 168.800 53.735 169.325 ;
        RECT 53.995 168.585 54.205 169.115 ;
        RECT 54.480 169.035 54.650 169.495 ;
        RECT 54.820 169.535 55.140 170.495 ;
        RECT 55.310 169.745 55.500 170.465 ;
        RECT 55.670 169.565 55.840 170.635 ;
        RECT 56.010 170.335 56.180 171.135 ;
        RECT 56.350 170.690 57.455 170.860 ;
        RECT 56.350 170.075 56.520 170.690 ;
        RECT 57.665 170.540 57.915 170.965 ;
        RECT 58.085 170.675 58.350 171.135 ;
        RECT 56.690 170.155 57.220 170.520 ;
        RECT 57.665 170.410 57.970 170.540 ;
        RECT 56.010 169.985 56.520 170.075 ;
        RECT 56.010 169.815 56.880 169.985 ;
        RECT 56.010 169.745 56.180 169.815 ;
        RECT 56.300 169.565 56.500 169.595 ;
        RECT 54.820 169.205 55.285 169.535 ;
        RECT 55.670 169.265 56.500 169.565 ;
        RECT 55.670 169.035 55.840 169.265 ;
        RECT 54.480 168.865 55.265 169.035 ;
        RECT 55.435 168.865 55.840 169.035 ;
        RECT 56.020 168.585 56.390 169.085 ;
        RECT 56.710 169.035 56.880 169.815 ;
        RECT 57.050 169.455 57.220 170.155 ;
        RECT 57.390 169.625 57.630 170.220 ;
        RECT 57.050 169.235 57.575 169.455 ;
        RECT 57.800 169.305 57.970 170.410 ;
        RECT 57.745 169.175 57.970 169.305 ;
        RECT 58.140 169.215 58.420 170.165 ;
        RECT 57.745 169.035 57.915 169.175 ;
        RECT 56.710 168.865 57.385 169.035 ;
        RECT 57.580 168.865 57.915 169.035 ;
        RECT 58.085 168.585 58.335 169.045 ;
        RECT 58.590 168.845 58.775 170.965 ;
        RECT 58.945 170.635 59.275 171.135 ;
        RECT 59.445 170.465 59.615 170.965 ;
        RECT 59.875 170.700 65.220 171.135 ;
        RECT 58.950 170.295 59.615 170.465 ;
        RECT 58.950 169.305 59.180 170.295 ;
        RECT 59.350 169.475 59.700 170.125 ;
        RECT 58.950 169.135 59.615 169.305 ;
        RECT 58.945 168.585 59.275 168.965 ;
        RECT 59.445 168.845 59.615 169.135 ;
        RECT 61.460 169.130 61.800 169.960 ;
        RECT 63.280 169.450 63.630 170.700 ;
        RECT 65.395 170.580 66.000 171.135 ;
        RECT 66.175 170.625 66.655 170.965 ;
        RECT 66.825 170.590 67.080 171.135 ;
        RECT 65.395 170.480 66.010 170.580 ;
        RECT 65.825 170.455 66.010 170.480 ;
        RECT 65.395 169.860 65.655 170.310 ;
        RECT 65.825 170.210 66.155 170.455 ;
        RECT 66.325 170.135 67.080 170.385 ;
        RECT 67.250 170.265 67.525 170.965 ;
        RECT 68.155 170.580 68.760 171.135 ;
        RECT 68.935 170.625 69.415 170.965 ;
        RECT 69.585 170.590 69.840 171.135 ;
        RECT 68.155 170.480 68.770 170.580 ;
        RECT 68.585 170.455 68.770 170.480 ;
        RECT 66.310 170.100 67.080 170.135 ;
        RECT 66.295 170.090 67.080 170.100 ;
        RECT 66.290 170.075 67.185 170.090 ;
        RECT 66.270 170.060 67.185 170.075 ;
        RECT 66.250 170.050 67.185 170.060 ;
        RECT 66.225 170.040 67.185 170.050 ;
        RECT 66.155 170.010 67.185 170.040 ;
        RECT 66.135 169.980 67.185 170.010 ;
        RECT 66.115 169.950 67.185 169.980 ;
        RECT 66.085 169.925 67.185 169.950 ;
        RECT 66.050 169.890 67.185 169.925 ;
        RECT 66.020 169.885 67.185 169.890 ;
        RECT 66.020 169.880 66.410 169.885 ;
        RECT 66.020 169.870 66.385 169.880 ;
        RECT 66.020 169.865 66.370 169.870 ;
        RECT 66.020 169.860 66.355 169.865 ;
        RECT 65.395 169.855 66.355 169.860 ;
        RECT 65.395 169.845 66.345 169.855 ;
        RECT 65.395 169.840 66.335 169.845 ;
        RECT 65.395 169.830 66.325 169.840 ;
        RECT 65.395 169.820 66.320 169.830 ;
        RECT 65.395 169.815 66.315 169.820 ;
        RECT 65.395 169.800 66.305 169.815 ;
        RECT 65.395 169.785 66.300 169.800 ;
        RECT 65.395 169.760 66.290 169.785 ;
        RECT 65.395 169.690 66.285 169.760 ;
        RECT 65.395 169.135 65.945 169.520 ;
        RECT 59.875 168.585 65.220 169.130 ;
        RECT 66.115 168.965 66.285 169.690 ;
        RECT 65.395 168.795 66.285 168.965 ;
        RECT 66.455 169.290 66.785 169.715 ;
        RECT 66.955 169.490 67.185 169.885 ;
        RECT 66.455 168.805 66.675 169.290 ;
        RECT 67.355 169.235 67.525 170.265 ;
        RECT 68.155 169.860 68.415 170.310 ;
        RECT 68.585 170.210 68.915 170.455 ;
        RECT 69.085 170.135 69.840 170.385 ;
        RECT 70.010 170.265 70.285 170.965 ;
        RECT 69.070 170.100 69.840 170.135 ;
        RECT 69.055 170.090 69.840 170.100 ;
        RECT 69.050 170.075 69.945 170.090 ;
        RECT 69.030 170.060 69.945 170.075 ;
        RECT 69.010 170.050 69.945 170.060 ;
        RECT 68.985 170.040 69.945 170.050 ;
        RECT 68.915 170.010 69.945 170.040 ;
        RECT 68.895 169.980 69.945 170.010 ;
        RECT 68.875 169.950 69.945 169.980 ;
        RECT 68.845 169.925 69.945 169.950 ;
        RECT 68.810 169.890 69.945 169.925 ;
        RECT 68.780 169.885 69.945 169.890 ;
        RECT 68.780 169.880 69.170 169.885 ;
        RECT 68.780 169.870 69.145 169.880 ;
        RECT 68.780 169.865 69.130 169.870 ;
        RECT 68.780 169.860 69.115 169.865 ;
        RECT 68.155 169.855 69.115 169.860 ;
        RECT 68.155 169.845 69.105 169.855 ;
        RECT 68.155 169.840 69.095 169.845 ;
        RECT 68.155 169.830 69.085 169.840 ;
        RECT 68.155 169.820 69.080 169.830 ;
        RECT 68.155 169.815 69.075 169.820 ;
        RECT 68.155 169.800 69.065 169.815 ;
        RECT 68.155 169.785 69.060 169.800 ;
        RECT 68.155 169.760 69.050 169.785 ;
        RECT 68.155 169.690 69.045 169.760 ;
        RECT 66.845 168.585 67.095 169.125 ;
        RECT 67.265 168.755 67.525 169.235 ;
        RECT 68.155 169.135 68.705 169.520 ;
        RECT 68.875 168.965 69.045 169.690 ;
        RECT 68.155 168.795 69.045 168.965 ;
        RECT 69.215 169.290 69.545 169.715 ;
        RECT 69.715 169.490 69.945 169.885 ;
        RECT 69.215 168.805 69.435 169.290 ;
        RECT 70.115 169.235 70.285 170.265 ;
        RECT 69.605 168.585 69.855 169.125 ;
        RECT 70.025 168.755 70.285 169.235 ;
        RECT 70.455 169.995 70.795 170.965 ;
        RECT 70.965 169.995 71.135 171.135 ;
        RECT 71.405 170.335 71.655 171.135 ;
        RECT 72.300 170.165 72.630 170.965 ;
        RECT 72.930 170.335 73.260 171.135 ;
        RECT 73.430 170.165 73.760 170.965 ;
        RECT 71.325 169.995 73.760 170.165 ;
        RECT 74.135 169.995 74.410 170.965 ;
        RECT 74.620 170.335 74.900 171.135 ;
        RECT 75.070 170.795 77.120 170.915 ;
        RECT 75.070 170.625 77.125 170.795 ;
        RECT 75.070 170.285 76.700 170.455 ;
        RECT 75.070 170.165 75.240 170.285 ;
        RECT 74.580 169.995 75.240 170.165 ;
        RECT 70.455 169.385 70.630 169.995 ;
        RECT 71.325 169.745 71.495 169.995 ;
        RECT 70.800 169.575 71.495 169.745 ;
        RECT 71.670 169.575 72.090 169.775 ;
        RECT 72.260 169.575 72.590 169.775 ;
        RECT 72.760 169.575 73.090 169.775 ;
        RECT 70.455 168.755 70.795 169.385 ;
        RECT 70.965 168.585 71.215 169.385 ;
        RECT 71.405 169.235 72.630 169.405 ;
        RECT 71.405 168.755 71.735 169.235 ;
        RECT 71.905 168.585 72.130 169.045 ;
        RECT 72.300 168.755 72.630 169.235 ;
        RECT 73.260 169.365 73.430 169.995 ;
        RECT 73.615 169.575 73.965 169.825 ;
        RECT 73.260 168.755 73.760 169.365 ;
        RECT 74.135 169.260 74.305 169.995 ;
        RECT 74.580 169.825 74.750 169.995 ;
        RECT 74.475 169.495 74.750 169.825 ;
        RECT 74.920 169.495 75.300 169.825 ;
        RECT 75.470 169.495 76.210 170.115 ;
        RECT 76.380 169.995 76.700 170.285 ;
        RECT 76.895 169.825 77.135 170.420 ;
        RECT 77.305 170.060 77.645 171.135 ;
        RECT 77.815 169.970 78.105 171.135 ;
        RECT 79.310 170.505 79.595 170.965 ;
        RECT 79.765 170.675 80.035 171.135 ;
        RECT 79.310 170.285 80.265 170.505 ;
        RECT 76.480 169.495 77.135 169.825 ;
        RECT 74.580 169.325 74.750 169.495 ;
        RECT 74.135 168.915 74.410 169.260 ;
        RECT 74.580 169.155 76.165 169.325 ;
        RECT 74.600 168.585 74.980 168.985 ;
        RECT 75.150 168.805 75.320 169.155 ;
        RECT 75.490 168.585 75.820 168.985 ;
        RECT 75.995 168.805 76.165 169.155 ;
        RECT 76.365 168.585 76.695 169.085 ;
        RECT 76.890 168.805 77.135 169.495 ;
        RECT 77.305 169.255 77.645 169.825 ;
        RECT 79.195 169.555 79.885 170.115 ;
        RECT 80.055 169.385 80.265 170.285 ;
        RECT 77.305 168.585 77.645 169.085 ;
        RECT 77.815 168.585 78.105 169.310 ;
        RECT 79.310 169.215 80.265 169.385 ;
        RECT 80.435 170.115 80.835 170.965 ;
        RECT 81.025 170.505 81.305 170.965 ;
        RECT 81.825 170.675 82.150 171.135 ;
        RECT 81.025 170.285 82.150 170.505 ;
        RECT 80.435 169.555 81.530 170.115 ;
        RECT 81.700 169.825 82.150 170.285 ;
        RECT 82.320 169.995 82.705 170.965 ;
        RECT 79.310 168.755 79.595 169.215 ;
        RECT 79.765 168.585 80.035 169.045 ;
        RECT 80.435 168.755 80.835 169.555 ;
        RECT 81.700 169.495 82.255 169.825 ;
        RECT 81.700 169.385 82.150 169.495 ;
        RECT 81.025 169.215 82.150 169.385 ;
        RECT 82.425 169.325 82.705 169.995 ;
        RECT 82.875 170.375 83.390 170.785 ;
        RECT 83.625 170.375 83.795 171.135 ;
        RECT 83.965 170.795 85.995 170.965 ;
        RECT 82.875 169.565 83.215 170.375 ;
        RECT 83.965 170.130 84.135 170.795 ;
        RECT 84.530 170.455 85.655 170.625 ;
        RECT 83.385 169.940 84.135 170.130 ;
        RECT 84.305 170.115 85.315 170.285 ;
        RECT 82.875 169.395 84.105 169.565 ;
        RECT 81.025 168.755 81.305 169.215 ;
        RECT 81.825 168.585 82.150 169.045 ;
        RECT 82.320 168.755 82.705 169.325 ;
        RECT 83.150 168.790 83.395 169.395 ;
        RECT 83.615 168.585 84.125 169.120 ;
        RECT 84.305 168.755 84.495 170.115 ;
        RECT 84.665 169.435 84.940 169.915 ;
        RECT 84.665 169.265 84.945 169.435 ;
        RECT 85.145 169.315 85.315 170.115 ;
        RECT 85.485 169.325 85.655 170.455 ;
        RECT 85.825 169.825 85.995 170.795 ;
        RECT 86.165 169.995 86.335 171.135 ;
        RECT 86.505 169.995 86.840 170.965 ;
        RECT 87.130 170.505 87.415 170.965 ;
        RECT 87.585 170.675 87.855 171.135 ;
        RECT 87.130 170.285 88.085 170.505 ;
        RECT 85.825 169.495 86.020 169.825 ;
        RECT 86.245 169.495 86.500 169.825 ;
        RECT 86.245 169.325 86.415 169.495 ;
        RECT 86.670 169.325 86.840 169.995 ;
        RECT 87.015 169.555 87.705 170.115 ;
        RECT 87.875 169.385 88.085 170.285 ;
        RECT 84.665 168.755 84.940 169.265 ;
        RECT 85.485 169.155 86.415 169.325 ;
        RECT 85.485 169.120 85.660 169.155 ;
        RECT 85.130 168.755 85.660 169.120 ;
        RECT 86.085 168.585 86.415 168.985 ;
        RECT 86.585 168.755 86.840 169.325 ;
        RECT 87.130 169.215 88.085 169.385 ;
        RECT 88.255 170.115 88.655 170.965 ;
        RECT 88.845 170.505 89.125 170.965 ;
        RECT 89.645 170.675 89.970 171.135 ;
        RECT 88.845 170.285 89.970 170.505 ;
        RECT 88.255 169.555 89.350 170.115 ;
        RECT 89.520 169.825 89.970 170.285 ;
        RECT 90.140 169.995 90.525 170.965 ;
        RECT 87.130 168.755 87.415 169.215 ;
        RECT 87.585 168.585 87.855 169.045 ;
        RECT 88.255 168.755 88.655 169.555 ;
        RECT 89.520 169.495 90.075 169.825 ;
        RECT 89.520 169.385 89.970 169.495 ;
        RECT 88.845 169.215 89.970 169.385 ;
        RECT 90.245 169.325 90.525 169.995 ;
        RECT 88.845 168.755 89.125 169.215 ;
        RECT 89.645 168.585 89.970 169.045 ;
        RECT 90.140 168.755 90.525 169.325 ;
        RECT 91.160 169.995 91.495 170.965 ;
        RECT 91.665 169.995 91.835 171.135 ;
        RECT 92.005 170.795 94.035 170.965 ;
        RECT 91.160 169.325 91.330 169.995 ;
        RECT 92.005 169.825 92.175 170.795 ;
        RECT 91.500 169.495 91.755 169.825 ;
        RECT 91.980 169.495 92.175 169.825 ;
        RECT 92.345 170.455 93.470 170.625 ;
        RECT 91.585 169.325 91.755 169.495 ;
        RECT 92.345 169.325 92.515 170.455 ;
        RECT 91.160 168.755 91.415 169.325 ;
        RECT 91.585 169.155 92.515 169.325 ;
        RECT 92.685 170.115 93.695 170.285 ;
        RECT 92.685 169.315 92.855 170.115 ;
        RECT 92.340 169.120 92.515 169.155 ;
        RECT 91.585 168.585 91.915 168.985 ;
        RECT 92.340 168.755 92.870 169.120 ;
        RECT 93.060 169.095 93.335 169.915 ;
        RECT 93.055 168.925 93.335 169.095 ;
        RECT 93.060 168.755 93.335 168.925 ;
        RECT 93.505 168.755 93.695 170.115 ;
        RECT 93.865 170.130 94.035 170.795 ;
        RECT 94.205 170.375 94.375 171.135 ;
        RECT 94.610 170.375 95.125 170.785 ;
        RECT 93.865 169.940 94.615 170.130 ;
        RECT 94.785 169.565 95.125 170.375 ;
        RECT 95.295 170.045 96.505 171.135 ;
        RECT 96.790 170.505 97.075 170.965 ;
        RECT 97.245 170.675 97.515 171.135 ;
        RECT 96.790 170.285 97.745 170.505 ;
        RECT 93.895 169.395 95.125 169.565 ;
        RECT 93.875 168.585 94.385 169.120 ;
        RECT 94.605 168.790 94.850 169.395 ;
        RECT 95.295 169.335 95.815 169.875 ;
        RECT 95.985 169.505 96.505 170.045 ;
        RECT 96.675 169.555 97.365 170.115 ;
        RECT 97.535 169.385 97.745 170.285 ;
        RECT 95.295 168.585 96.505 169.335 ;
        RECT 96.790 169.215 97.745 169.385 ;
        RECT 97.915 170.115 98.315 170.965 ;
        RECT 98.505 170.505 98.785 170.965 ;
        RECT 99.305 170.675 99.630 171.135 ;
        RECT 98.505 170.285 99.630 170.505 ;
        RECT 97.915 169.555 99.010 170.115 ;
        RECT 99.180 169.825 99.630 170.285 ;
        RECT 99.800 169.995 100.185 170.965 ;
        RECT 100.355 170.045 102.945 171.135 ;
        RECT 96.790 168.755 97.075 169.215 ;
        RECT 97.245 168.585 97.515 169.045 ;
        RECT 97.915 168.755 98.315 169.555 ;
        RECT 99.180 169.495 99.735 169.825 ;
        RECT 99.180 169.385 99.630 169.495 ;
        RECT 98.505 169.215 99.630 169.385 ;
        RECT 99.905 169.325 100.185 169.995 ;
        RECT 98.505 168.755 98.785 169.215 ;
        RECT 99.305 168.585 99.630 169.045 ;
        RECT 99.800 168.755 100.185 169.325 ;
        RECT 100.355 169.355 101.565 169.875 ;
        RECT 101.735 169.525 102.945 170.045 ;
        RECT 103.575 169.970 103.865 171.135 ;
        RECT 104.035 170.700 109.380 171.135 ;
        RECT 100.355 168.585 102.945 169.355 ;
        RECT 103.575 168.585 103.865 169.310 ;
        RECT 105.620 169.130 105.960 169.960 ;
        RECT 107.440 169.450 107.790 170.700 ;
        RECT 109.555 170.045 113.065 171.135 ;
        RECT 113.895 170.465 114.175 171.135 ;
        RECT 114.345 170.245 114.645 170.795 ;
        RECT 114.845 170.415 115.175 171.135 ;
        RECT 115.365 170.415 115.825 170.965 ;
        RECT 109.555 169.355 111.205 169.875 ;
        RECT 111.375 169.525 113.065 170.045 ;
        RECT 113.710 169.825 113.975 170.185 ;
        RECT 114.345 170.075 115.285 170.245 ;
        RECT 115.115 169.825 115.285 170.075 ;
        RECT 113.710 169.575 114.385 169.825 ;
        RECT 114.605 169.575 114.945 169.825 ;
        RECT 115.115 169.495 115.405 169.825 ;
        RECT 115.115 169.405 115.285 169.495 ;
        RECT 104.035 168.585 109.380 169.130 ;
        RECT 109.555 168.585 113.065 169.355 ;
        RECT 113.895 169.215 115.285 169.405 ;
        RECT 113.895 168.855 114.225 169.215 ;
        RECT 115.575 169.045 115.825 170.415 ;
        RECT 114.845 168.585 115.095 169.045 ;
        RECT 115.265 168.755 115.825 169.045 ;
        RECT 115.995 170.025 116.255 170.965 ;
        RECT 116.425 170.735 116.755 171.135 ;
        RECT 117.900 170.870 118.155 170.965 ;
        RECT 117.015 170.700 118.155 170.870 ;
        RECT 118.325 170.755 118.655 170.925 ;
        RECT 117.015 170.475 117.185 170.700 ;
        RECT 116.425 170.305 117.185 170.475 ;
        RECT 117.900 170.565 118.155 170.700 ;
        RECT 115.995 169.310 116.170 170.025 ;
        RECT 116.425 169.825 116.595 170.305 ;
        RECT 117.450 170.215 117.620 170.405 ;
        RECT 117.900 170.395 118.310 170.565 ;
        RECT 116.340 169.495 116.595 169.825 ;
        RECT 116.820 169.495 117.150 170.115 ;
        RECT 117.450 170.045 117.970 170.215 ;
        RECT 117.320 169.495 117.610 169.875 ;
        RECT 117.800 169.325 117.970 170.045 ;
        RECT 115.995 168.755 116.255 169.310 ;
        RECT 117.090 169.155 117.970 169.325 ;
        RECT 118.140 169.370 118.310 170.395 ;
        RECT 118.485 170.505 118.655 170.755 ;
        RECT 118.825 170.675 119.075 171.135 ;
        RECT 119.245 170.505 119.425 170.965 ;
        RECT 118.485 170.335 119.425 170.505 ;
        RECT 119.880 170.165 120.210 170.965 ;
        RECT 120.380 170.335 120.710 171.135 ;
        RECT 121.010 170.165 121.340 170.965 ;
        RECT 121.985 170.335 122.235 171.135 ;
        RECT 118.510 169.855 118.990 170.155 ;
        RECT 118.140 169.200 118.490 169.370 ;
        RECT 118.730 169.265 118.990 169.855 ;
        RECT 119.190 169.265 119.450 170.155 ;
        RECT 119.880 169.995 122.315 170.165 ;
        RECT 122.505 169.995 122.675 171.135 ;
        RECT 122.845 169.995 123.185 170.965 ;
        RECT 119.675 169.575 120.025 169.825 ;
        RECT 120.210 169.365 120.380 169.995 ;
        RECT 120.550 169.575 120.880 169.775 ;
        RECT 121.050 169.575 121.380 169.775 ;
        RECT 121.550 169.575 121.970 169.775 ;
        RECT 122.145 169.745 122.315 169.995 ;
        RECT 122.145 169.575 122.840 169.745 ;
        RECT 116.425 168.585 116.855 169.030 ;
        RECT 117.090 168.755 117.260 169.155 ;
        RECT 117.430 168.585 118.150 168.985 ;
        RECT 118.320 168.755 118.490 169.200 ;
        RECT 119.065 168.585 119.465 169.095 ;
        RECT 119.880 168.755 120.380 169.365 ;
        RECT 121.010 169.235 122.235 169.405 ;
        RECT 123.010 169.385 123.185 169.995 ;
        RECT 123.360 170.745 123.695 170.965 ;
        RECT 124.700 170.755 125.055 171.135 ;
        RECT 123.360 170.125 123.615 170.745 ;
        RECT 123.865 170.585 124.095 170.625 ;
        RECT 125.225 170.585 125.475 170.965 ;
        RECT 123.865 170.385 125.475 170.585 ;
        RECT 123.865 170.295 124.050 170.385 ;
        RECT 124.640 170.375 125.475 170.385 ;
        RECT 125.725 170.355 125.975 171.135 ;
        RECT 126.145 170.285 126.405 170.965 ;
        RECT 124.205 170.185 124.535 170.215 ;
        RECT 124.205 170.125 126.005 170.185 ;
        RECT 123.360 170.015 126.065 170.125 ;
        RECT 123.360 169.955 124.535 170.015 ;
        RECT 125.865 169.980 126.065 170.015 ;
        RECT 123.355 169.575 123.845 169.775 ;
        RECT 124.035 169.575 124.510 169.785 ;
        RECT 121.010 168.755 121.340 169.235 ;
        RECT 121.510 168.585 121.735 169.045 ;
        RECT 121.905 168.755 122.235 169.235 ;
        RECT 122.425 168.585 122.675 169.385 ;
        RECT 122.845 168.755 123.185 169.385 ;
        RECT 123.360 168.585 123.815 169.350 ;
        RECT 124.290 169.175 124.510 169.575 ;
        RECT 124.755 169.575 125.085 169.785 ;
        RECT 124.755 169.175 124.965 169.575 ;
        RECT 125.255 169.540 125.665 169.845 ;
        RECT 125.895 169.405 126.065 169.980 ;
        RECT 125.795 169.285 126.065 169.405 ;
        RECT 125.220 169.240 126.065 169.285 ;
        RECT 125.220 169.115 125.975 169.240 ;
        RECT 125.220 168.965 125.390 169.115 ;
        RECT 126.235 169.085 126.405 170.285 ;
        RECT 126.575 170.045 129.165 171.135 ;
        RECT 124.090 168.755 125.390 168.965 ;
        RECT 125.645 168.585 125.975 168.945 ;
        RECT 126.145 168.755 126.405 169.085 ;
        RECT 126.575 169.355 127.785 169.875 ;
        RECT 127.955 169.525 129.165 170.045 ;
        RECT 129.335 169.970 129.625 171.135 ;
        RECT 129.800 169.995 130.135 170.965 ;
        RECT 130.305 169.995 130.475 171.135 ;
        RECT 130.645 170.795 132.675 170.965 ;
        RECT 126.575 168.585 129.165 169.355 ;
        RECT 129.800 169.325 129.970 169.995 ;
        RECT 130.645 169.825 130.815 170.795 ;
        RECT 130.140 169.495 130.395 169.825 ;
        RECT 130.620 169.495 130.815 169.825 ;
        RECT 130.985 170.455 132.110 170.625 ;
        RECT 130.225 169.325 130.395 169.495 ;
        RECT 130.985 169.325 131.155 170.455 ;
        RECT 129.335 168.585 129.625 169.310 ;
        RECT 129.800 168.755 130.055 169.325 ;
        RECT 130.225 169.155 131.155 169.325 ;
        RECT 131.325 170.115 132.335 170.285 ;
        RECT 131.325 169.315 131.495 170.115 ;
        RECT 131.700 169.435 131.975 169.915 ;
        RECT 131.695 169.265 131.975 169.435 ;
        RECT 130.980 169.120 131.155 169.155 ;
        RECT 130.225 168.585 130.555 168.985 ;
        RECT 130.980 168.755 131.510 169.120 ;
        RECT 131.700 168.755 131.975 169.265 ;
        RECT 132.145 168.755 132.335 170.115 ;
        RECT 132.505 170.130 132.675 170.795 ;
        RECT 132.845 170.375 133.015 171.135 ;
        RECT 133.250 170.375 133.765 170.785 ;
        RECT 132.505 169.940 133.255 170.130 ;
        RECT 133.425 169.565 133.765 170.375 ;
        RECT 132.535 169.395 133.765 169.565 ;
        RECT 133.935 169.995 134.320 170.965 ;
        RECT 134.490 170.675 134.815 171.135 ;
        RECT 135.335 170.505 135.615 170.965 ;
        RECT 134.490 170.285 135.615 170.505 ;
        RECT 132.515 168.585 133.025 169.120 ;
        RECT 133.245 168.790 133.490 169.395 ;
        RECT 133.935 169.325 134.215 169.995 ;
        RECT 134.490 169.825 134.940 170.285 ;
        RECT 135.805 170.115 136.205 170.965 ;
        RECT 136.605 170.675 136.875 171.135 ;
        RECT 137.045 170.505 137.330 170.965 ;
        RECT 134.385 169.495 134.940 169.825 ;
        RECT 135.110 169.555 136.205 170.115 ;
        RECT 134.490 169.385 134.940 169.495 ;
        RECT 133.935 168.755 134.320 169.325 ;
        RECT 134.490 169.215 135.615 169.385 ;
        RECT 134.490 168.585 134.815 169.045 ;
        RECT 135.335 168.755 135.615 169.215 ;
        RECT 135.805 168.755 136.205 169.555 ;
        RECT 136.375 170.285 137.330 170.505 ;
        RECT 136.375 169.385 136.585 170.285 ;
        RECT 136.755 169.555 137.445 170.115 ;
        RECT 137.615 170.045 138.825 171.135 ;
        RECT 137.615 169.505 138.135 170.045 ;
        RECT 136.375 169.215 137.330 169.385 ;
        RECT 138.305 169.335 138.825 169.875 ;
        RECT 136.605 168.585 136.875 169.045 ;
        RECT 137.045 168.755 137.330 169.215 ;
        RECT 137.615 168.585 138.825 169.335 ;
        RECT 13.330 168.415 138.910 168.585 ;
        RECT 13.415 167.665 14.625 168.415 ;
        RECT 13.415 167.125 13.935 167.665 ;
        RECT 14.795 167.645 16.465 168.415 ;
        RECT 17.145 167.760 17.475 168.195 ;
        RECT 17.645 167.805 17.815 168.415 ;
        RECT 17.095 167.675 17.475 167.760 ;
        RECT 17.985 167.675 18.315 168.200 ;
        RECT 18.575 167.885 18.785 168.415 ;
        RECT 19.060 167.965 19.845 168.135 ;
        RECT 20.015 167.965 20.420 168.135 ;
        RECT 14.105 166.955 14.625 167.495 ;
        RECT 14.795 167.125 15.545 167.645 ;
        RECT 17.095 167.635 17.320 167.675 ;
        RECT 15.715 166.955 16.465 167.475 ;
        RECT 13.415 165.865 14.625 166.955 ;
        RECT 14.795 165.865 16.465 166.955 ;
        RECT 17.095 167.055 17.265 167.635 ;
        RECT 17.985 167.505 18.185 167.675 ;
        RECT 19.060 167.505 19.230 167.965 ;
        RECT 17.435 167.175 18.185 167.505 ;
        RECT 18.355 167.175 19.230 167.505 ;
        RECT 17.095 167.005 17.310 167.055 ;
        RECT 17.095 166.925 17.485 167.005 ;
        RECT 17.155 166.080 17.485 166.925 ;
        RECT 17.995 166.970 18.185 167.175 ;
        RECT 17.655 165.865 17.825 166.875 ;
        RECT 17.995 166.595 18.890 166.970 ;
        RECT 17.995 166.035 18.335 166.595 ;
        RECT 18.565 165.865 18.880 166.365 ;
        RECT 19.060 166.335 19.230 167.175 ;
        RECT 19.400 167.465 19.865 167.795 ;
        RECT 20.250 167.735 20.420 167.965 ;
        RECT 20.600 167.915 20.970 168.415 ;
        RECT 21.290 167.965 21.965 168.135 ;
        RECT 22.160 167.965 22.495 168.135 ;
        RECT 19.400 166.505 19.720 167.465 ;
        RECT 20.250 167.435 21.080 167.735 ;
        RECT 19.890 166.535 20.080 167.255 ;
        RECT 20.250 166.365 20.420 167.435 ;
        RECT 20.880 167.405 21.080 167.435 ;
        RECT 20.590 167.185 20.760 167.255 ;
        RECT 21.290 167.185 21.460 167.965 ;
        RECT 22.325 167.825 22.495 167.965 ;
        RECT 22.665 167.955 22.915 168.415 ;
        RECT 20.590 167.015 21.460 167.185 ;
        RECT 21.630 167.545 22.155 167.765 ;
        RECT 22.325 167.695 22.550 167.825 ;
        RECT 20.590 166.925 21.100 167.015 ;
        RECT 19.060 166.165 19.945 166.335 ;
        RECT 20.170 166.035 20.420 166.365 ;
        RECT 20.590 165.865 20.760 166.665 ;
        RECT 20.930 166.310 21.100 166.925 ;
        RECT 21.630 166.845 21.800 167.545 ;
        RECT 21.270 166.480 21.800 166.845 ;
        RECT 21.970 166.780 22.210 167.375 ;
        RECT 22.380 166.590 22.550 167.695 ;
        RECT 22.720 166.835 23.000 167.785 ;
        RECT 22.245 166.460 22.550 166.590 ;
        RECT 20.930 166.140 22.035 166.310 ;
        RECT 22.245 166.035 22.495 166.460 ;
        RECT 22.665 165.865 22.930 166.325 ;
        RECT 23.170 166.035 23.355 168.155 ;
        RECT 23.525 168.035 23.855 168.415 ;
        RECT 24.025 167.865 24.195 168.155 ;
        RECT 23.530 167.695 24.195 167.865 ;
        RECT 23.530 166.705 23.760 167.695 ;
        RECT 24.455 167.645 27.045 168.415 ;
        RECT 27.680 167.765 27.950 167.975 ;
        RECT 28.170 167.955 28.500 168.415 ;
        RECT 29.010 167.955 29.760 168.245 ;
        RECT 23.930 166.875 24.280 167.525 ;
        RECT 24.455 167.125 25.665 167.645 ;
        RECT 27.680 167.595 29.015 167.765 ;
        RECT 25.835 166.955 27.045 167.475 ;
        RECT 28.845 167.425 29.015 167.595 ;
        RECT 27.680 167.185 28.030 167.425 ;
        RECT 28.200 167.185 28.675 167.425 ;
        RECT 28.845 167.175 29.220 167.425 ;
        RECT 28.845 167.005 29.015 167.175 ;
        RECT 23.530 166.535 24.195 166.705 ;
        RECT 23.525 165.865 23.855 166.365 ;
        RECT 24.025 166.035 24.195 166.535 ;
        RECT 24.455 165.865 27.045 166.955 ;
        RECT 27.680 166.835 29.015 167.005 ;
        RECT 27.680 166.675 27.960 166.835 ;
        RECT 29.390 166.665 29.760 167.955 ;
        RECT 29.980 167.650 30.435 168.415 ;
        RECT 30.710 168.035 32.010 168.245 ;
        RECT 32.265 168.055 32.595 168.415 ;
        RECT 31.840 167.885 32.010 168.035 ;
        RECT 32.765 167.915 33.025 168.245 ;
        RECT 32.795 167.905 33.025 167.915 ;
        RECT 30.910 167.425 31.130 167.825 ;
        RECT 29.975 167.225 30.465 167.425 ;
        RECT 30.655 167.215 31.130 167.425 ;
        RECT 31.375 167.425 31.585 167.825 ;
        RECT 31.840 167.760 32.595 167.885 ;
        RECT 31.840 167.715 32.685 167.760 ;
        RECT 32.415 167.595 32.685 167.715 ;
        RECT 31.375 167.215 31.705 167.425 ;
        RECT 31.875 167.155 32.285 167.460 ;
        RECT 28.170 165.865 28.420 166.665 ;
        RECT 28.590 166.495 29.760 166.665 ;
        RECT 29.980 166.985 31.155 167.045 ;
        RECT 32.515 167.020 32.685 167.595 ;
        RECT 32.485 166.985 32.685 167.020 ;
        RECT 29.980 166.875 32.685 166.985 ;
        RECT 28.590 166.035 28.920 166.495 ;
        RECT 29.090 165.865 29.305 166.325 ;
        RECT 29.980 166.255 30.235 166.875 ;
        RECT 30.825 166.815 32.625 166.875 ;
        RECT 30.825 166.785 31.155 166.815 ;
        RECT 32.855 166.715 33.025 167.905 ;
        RECT 33.195 167.665 34.405 168.415 ;
        RECT 34.575 167.675 34.915 168.245 ;
        RECT 35.110 167.750 35.280 168.415 ;
        RECT 35.560 168.075 35.780 168.120 ;
        RECT 35.555 167.905 35.780 168.075 ;
        RECT 35.950 167.935 36.395 168.105 ;
        RECT 35.560 167.765 35.780 167.905 ;
        RECT 33.195 167.125 33.715 167.665 ;
        RECT 33.885 166.955 34.405 167.495 ;
        RECT 30.485 166.615 30.670 166.705 ;
        RECT 31.260 166.615 32.095 166.625 ;
        RECT 30.485 166.415 32.095 166.615 ;
        RECT 30.485 166.375 30.715 166.415 ;
        RECT 29.980 166.035 30.315 166.255 ;
        RECT 31.320 165.865 31.675 166.245 ;
        RECT 31.845 166.035 32.095 166.415 ;
        RECT 32.345 165.865 32.595 166.645 ;
        RECT 32.765 166.035 33.025 166.715 ;
        RECT 33.195 165.865 34.405 166.955 ;
        RECT 34.575 166.705 34.750 167.675 ;
        RECT 35.560 167.595 36.055 167.765 ;
        RECT 34.920 167.055 35.090 167.505 ;
        RECT 35.260 167.225 35.710 167.425 ;
        RECT 35.880 167.400 36.055 167.595 ;
        RECT 36.225 167.145 36.395 167.935 ;
        RECT 36.565 167.810 36.815 168.180 ;
        RECT 36.645 167.425 36.815 167.810 ;
        RECT 36.985 167.775 37.235 168.180 ;
        RECT 37.405 167.945 37.575 168.415 ;
        RECT 37.745 167.775 38.085 168.180 ;
        RECT 36.985 167.595 38.085 167.775 ;
        RECT 39.175 167.690 39.465 168.415 ;
        RECT 39.635 167.645 41.305 168.415 ;
        RECT 41.485 168.055 43.555 168.245 ;
        RECT 43.785 168.055 44.115 168.415 ;
        RECT 44.645 168.055 44.975 168.415 ;
        RECT 45.505 168.055 45.835 168.415 ;
        RECT 42.435 168.035 43.555 168.055 ;
        RECT 36.645 167.255 36.840 167.425 ;
        RECT 34.920 166.885 35.315 167.055 ;
        RECT 36.225 167.005 36.500 167.145 ;
        RECT 34.575 166.035 34.835 166.705 ;
        RECT 35.145 166.615 35.315 166.885 ;
        RECT 35.485 166.785 36.500 167.005 ;
        RECT 36.670 167.005 36.840 167.255 ;
        RECT 37.010 167.175 37.570 167.425 ;
        RECT 36.670 166.615 37.225 167.005 ;
        RECT 35.145 166.445 37.225 166.615 ;
        RECT 35.005 165.865 35.335 166.265 ;
        RECT 36.205 165.865 36.605 166.265 ;
        RECT 36.895 166.210 37.225 166.445 ;
        RECT 37.395 166.075 37.570 167.175 ;
        RECT 37.740 166.855 38.085 167.425 ;
        RECT 39.635 167.125 40.385 167.645 ;
        RECT 37.740 165.865 38.085 166.685 ;
        RECT 39.175 165.865 39.465 167.030 ;
        RECT 40.555 166.955 41.305 167.475 ;
        RECT 39.635 165.865 41.305 166.955 ;
        RECT 41.475 166.530 41.765 167.505 ;
        RECT 41.935 166.960 42.265 167.830 ;
        RECT 42.435 167.610 42.625 168.035 ;
        RECT 45.145 167.865 45.335 167.985 ;
        RECT 42.795 167.655 45.335 167.865 ;
        RECT 45.505 167.425 45.845 167.735 ;
        RECT 46.075 167.615 46.770 168.245 ;
        RECT 46.975 167.615 47.285 168.415 ;
        RECT 47.540 167.845 47.715 168.245 ;
        RECT 47.885 168.035 48.215 168.415 ;
        RECT 48.460 167.915 48.690 168.245 ;
        RECT 47.540 167.675 48.170 167.845 ;
        RECT 42.435 167.135 43.295 167.425 ;
        RECT 43.755 167.145 44.725 167.425 ;
        RECT 44.895 167.255 45.845 167.425 ;
        RECT 44.950 167.205 45.845 167.255 ;
        RECT 46.095 167.175 46.430 167.425 ;
        RECT 46.600 167.015 46.770 167.615 ;
        RECT 48.000 167.505 48.170 167.675 ;
        RECT 46.940 167.175 47.275 167.445 ;
        RECT 41.935 166.790 44.545 166.960 ;
        RECT 41.505 165.865 41.765 166.325 ;
        RECT 41.935 166.035 42.195 166.790 ;
        RECT 42.365 165.865 42.695 166.585 ;
        RECT 42.865 166.035 43.055 166.790 ;
        RECT 43.225 165.865 43.555 166.585 ;
        RECT 43.785 166.205 44.045 166.400 ;
        RECT 44.215 166.375 44.545 166.790 ;
        RECT 44.715 166.805 45.835 166.975 ;
        RECT 44.715 166.205 44.905 166.805 ;
        RECT 43.785 166.035 44.905 166.205 ;
        RECT 45.075 165.865 45.405 166.635 ;
        RECT 45.575 166.035 45.835 166.805 ;
        RECT 46.075 165.865 46.335 167.005 ;
        RECT 46.505 166.035 46.835 167.015 ;
        RECT 47.005 165.865 47.285 167.005 ;
        RECT 47.455 166.825 47.820 167.505 ;
        RECT 48.000 167.175 48.350 167.505 ;
        RECT 48.000 166.655 48.170 167.175 ;
        RECT 47.540 166.485 48.170 166.655 ;
        RECT 48.520 166.625 48.690 167.915 ;
        RECT 48.890 166.805 49.170 168.080 ;
        RECT 49.395 168.075 49.665 168.080 ;
        RECT 49.355 167.905 49.665 168.075 ;
        RECT 50.125 168.035 50.455 168.415 ;
        RECT 50.625 168.160 50.960 168.205 ;
        RECT 49.395 166.805 49.665 167.905 ;
        RECT 49.855 166.805 50.195 167.835 ;
        RECT 50.625 167.695 50.965 168.160 ;
        RECT 51.185 167.760 51.515 168.195 ;
        RECT 51.685 167.805 51.855 168.415 ;
        RECT 50.365 167.175 50.625 167.505 ;
        RECT 50.365 166.625 50.535 167.175 ;
        RECT 50.795 167.005 50.965 167.695 ;
        RECT 47.540 166.035 47.715 166.485 ;
        RECT 48.520 166.455 50.535 166.625 ;
        RECT 47.885 165.865 48.215 166.305 ;
        RECT 48.520 166.035 48.690 166.455 ;
        RECT 48.925 165.865 49.595 166.275 ;
        RECT 49.810 166.035 49.980 166.455 ;
        RECT 50.180 165.865 50.510 166.275 ;
        RECT 50.705 166.035 50.965 167.005 ;
        RECT 51.135 167.675 51.515 167.760 ;
        RECT 52.025 167.675 52.355 168.200 ;
        RECT 52.615 167.885 52.825 168.415 ;
        RECT 53.100 167.965 53.885 168.135 ;
        RECT 54.055 167.965 54.460 168.135 ;
        RECT 51.135 167.635 51.360 167.675 ;
        RECT 51.135 167.055 51.305 167.635 ;
        RECT 52.025 167.505 52.225 167.675 ;
        RECT 53.100 167.505 53.270 167.965 ;
        RECT 51.475 167.175 52.225 167.505 ;
        RECT 52.395 167.175 53.270 167.505 ;
        RECT 51.135 167.005 51.350 167.055 ;
        RECT 51.135 166.925 51.525 167.005 ;
        RECT 51.195 166.080 51.525 166.925 ;
        RECT 52.035 166.970 52.225 167.175 ;
        RECT 51.695 165.865 51.865 166.875 ;
        RECT 52.035 166.595 52.930 166.970 ;
        RECT 52.035 166.035 52.375 166.595 ;
        RECT 52.605 165.865 52.920 166.365 ;
        RECT 53.100 166.335 53.270 167.175 ;
        RECT 53.440 167.465 53.905 167.795 ;
        RECT 54.290 167.735 54.460 167.965 ;
        RECT 54.640 167.915 55.010 168.415 ;
        RECT 55.330 167.965 56.005 168.135 ;
        RECT 56.200 167.965 56.535 168.135 ;
        RECT 53.440 166.505 53.760 167.465 ;
        RECT 54.290 167.435 55.120 167.735 ;
        RECT 53.930 166.535 54.120 167.255 ;
        RECT 54.290 166.365 54.460 167.435 ;
        RECT 54.920 167.405 55.120 167.435 ;
        RECT 54.630 167.185 54.800 167.255 ;
        RECT 55.330 167.185 55.500 167.965 ;
        RECT 56.365 167.825 56.535 167.965 ;
        RECT 56.705 167.955 56.955 168.415 ;
        RECT 54.630 167.015 55.500 167.185 ;
        RECT 55.670 167.545 56.195 167.765 ;
        RECT 56.365 167.695 56.590 167.825 ;
        RECT 54.630 166.925 55.140 167.015 ;
        RECT 53.100 166.165 53.985 166.335 ;
        RECT 54.210 166.035 54.460 166.365 ;
        RECT 54.630 165.865 54.800 166.665 ;
        RECT 54.970 166.310 55.140 166.925 ;
        RECT 55.670 166.845 55.840 167.545 ;
        RECT 55.310 166.480 55.840 166.845 ;
        RECT 56.010 166.780 56.250 167.375 ;
        RECT 56.420 166.590 56.590 167.695 ;
        RECT 56.760 166.835 57.040 167.785 ;
        RECT 56.285 166.460 56.590 166.590 ;
        RECT 54.970 166.140 56.075 166.310 ;
        RECT 56.285 166.035 56.535 166.460 ;
        RECT 56.705 165.865 56.970 166.325 ;
        RECT 57.210 166.035 57.395 168.155 ;
        RECT 57.565 168.035 57.895 168.415 ;
        RECT 58.500 168.160 58.835 168.205 ;
        RECT 58.065 167.865 58.235 168.155 ;
        RECT 57.570 167.695 58.235 167.865 ;
        RECT 58.495 167.695 58.835 168.160 ;
        RECT 59.005 168.035 59.335 168.415 ;
        RECT 57.570 166.705 57.800 167.695 ;
        RECT 57.970 166.875 58.320 167.525 ;
        RECT 58.495 167.005 58.665 167.695 ;
        RECT 58.835 167.175 59.095 167.505 ;
        RECT 57.570 166.535 58.235 166.705 ;
        RECT 57.565 165.865 57.895 166.365 ;
        RECT 58.065 166.035 58.235 166.535 ;
        RECT 58.495 166.035 58.755 167.005 ;
        RECT 58.925 166.625 59.095 167.175 ;
        RECT 59.265 166.805 59.605 167.835 ;
        RECT 59.795 167.735 60.065 168.080 ;
        RECT 59.795 167.565 60.105 167.735 ;
        RECT 59.795 166.805 60.065 167.565 ;
        RECT 60.290 166.805 60.570 168.080 ;
        RECT 60.770 167.915 61.000 168.245 ;
        RECT 61.245 168.035 61.575 168.415 ;
        RECT 60.770 166.625 60.940 167.915 ;
        RECT 61.745 167.845 61.920 168.245 ;
        RECT 61.290 167.675 61.920 167.845 ;
        RECT 61.290 167.505 61.460 167.675 ;
        RECT 62.175 167.645 64.765 168.415 ;
        RECT 64.935 167.690 65.225 168.415 ;
        RECT 65.395 167.645 67.065 168.415 ;
        RECT 67.240 167.910 67.575 168.415 ;
        RECT 67.745 167.845 67.985 168.220 ;
        RECT 68.265 168.085 68.435 168.230 ;
        RECT 68.265 167.890 68.640 168.085 ;
        RECT 69.000 167.920 69.395 168.415 ;
        RECT 61.110 167.175 61.460 167.505 ;
        RECT 58.925 166.455 60.940 166.625 ;
        RECT 61.290 166.655 61.460 167.175 ;
        RECT 61.640 166.825 62.005 167.505 ;
        RECT 62.175 167.125 63.385 167.645 ;
        RECT 63.555 166.955 64.765 167.475 ;
        RECT 65.395 167.125 66.145 167.645 ;
        RECT 61.290 166.485 61.920 166.655 ;
        RECT 58.950 165.865 59.280 166.275 ;
        RECT 59.480 166.035 59.650 166.455 ;
        RECT 59.865 165.865 60.535 166.275 ;
        RECT 60.770 166.035 60.940 166.455 ;
        RECT 61.245 165.865 61.575 166.305 ;
        RECT 61.745 166.035 61.920 166.485 ;
        RECT 62.175 165.865 64.765 166.955 ;
        RECT 64.935 165.865 65.225 167.030 ;
        RECT 66.315 166.955 67.065 167.475 ;
        RECT 65.395 165.865 67.065 166.955 ;
        RECT 67.295 166.885 67.595 167.735 ;
        RECT 67.765 167.695 67.985 167.845 ;
        RECT 67.765 167.365 68.300 167.695 ;
        RECT 68.470 167.555 68.640 167.890 ;
        RECT 69.565 167.725 69.805 168.245 ;
        RECT 70.005 167.915 70.335 168.415 ;
        RECT 70.535 167.845 70.705 168.195 ;
        RECT 70.905 168.015 71.235 168.415 ;
        RECT 71.405 167.845 71.575 168.195 ;
        RECT 71.745 168.015 72.125 168.415 ;
        RECT 67.765 166.715 68.000 167.365 ;
        RECT 68.470 167.195 69.455 167.555 ;
        RECT 67.325 166.485 68.000 166.715 ;
        RECT 68.170 167.175 69.455 167.195 ;
        RECT 68.170 167.025 69.030 167.175 ;
        RECT 67.325 166.055 67.495 166.485 ;
        RECT 67.665 165.865 67.995 166.315 ;
        RECT 68.170 166.080 68.455 167.025 ;
        RECT 69.630 166.920 69.805 167.725 ;
        RECT 70.000 167.175 70.350 167.745 ;
        RECT 70.535 167.675 72.145 167.845 ;
        RECT 72.315 167.740 72.585 168.085 ;
        RECT 71.975 167.505 72.145 167.675 ;
        RECT 68.630 166.545 69.325 166.855 ;
        RECT 68.635 165.865 69.320 166.335 ;
        RECT 69.500 166.135 69.805 166.920 ;
        RECT 70.000 166.715 70.320 167.005 ;
        RECT 70.520 166.885 71.230 167.505 ;
        RECT 71.400 167.175 71.805 167.505 ;
        RECT 71.975 167.175 72.245 167.505 ;
        RECT 71.975 167.005 72.145 167.175 ;
        RECT 72.415 167.005 72.585 167.740 ;
        RECT 72.805 167.875 73.030 168.235 ;
        RECT 73.210 168.045 73.540 168.415 ;
        RECT 73.720 167.875 73.975 168.235 ;
        RECT 74.540 168.045 75.285 168.415 ;
        RECT 72.805 167.685 75.290 167.875 ;
        RECT 72.765 167.175 73.035 167.505 ;
        RECT 73.215 167.175 73.650 167.505 ;
        RECT 73.830 167.175 74.405 167.505 ;
        RECT 74.585 167.175 74.865 167.505 ;
        RECT 71.420 166.835 72.145 167.005 ;
        RECT 71.420 166.715 71.590 166.835 ;
        RECT 70.000 166.545 71.590 166.715 ;
        RECT 70.000 166.085 71.655 166.375 ;
        RECT 71.825 165.865 72.105 166.665 ;
        RECT 72.315 166.035 72.585 167.005 ;
        RECT 75.065 166.995 75.290 167.685 ;
        RECT 72.795 166.815 75.290 166.995 ;
        RECT 75.465 166.815 75.800 168.235 ;
        RECT 72.795 166.045 73.085 166.815 ;
        RECT 73.655 166.405 74.845 166.635 ;
        RECT 73.655 166.045 73.915 166.405 ;
        RECT 74.085 165.865 74.415 166.235 ;
        RECT 74.585 166.045 74.845 166.405 ;
        RECT 75.035 165.865 75.365 166.585 ;
        RECT 75.535 166.045 75.800 166.815 ;
        RECT 76.895 167.765 77.155 168.245 ;
        RECT 77.325 167.955 77.655 168.415 ;
        RECT 77.845 167.775 78.045 168.195 ;
        RECT 76.895 166.735 77.065 167.765 ;
        RECT 77.235 167.075 77.465 167.505 ;
        RECT 77.635 167.255 78.045 167.775 ;
        RECT 78.215 167.930 79.005 168.195 ;
        RECT 78.215 167.075 78.470 167.930 ;
        RECT 79.185 167.595 79.515 168.015 ;
        RECT 79.685 167.595 79.945 168.415 ;
        RECT 80.165 167.760 80.495 168.195 ;
        RECT 80.665 167.805 80.835 168.415 ;
        RECT 80.115 167.675 80.495 167.760 ;
        RECT 81.005 167.675 81.335 168.200 ;
        RECT 81.595 167.885 81.805 168.415 ;
        RECT 82.080 167.965 82.865 168.135 ;
        RECT 83.035 167.965 83.440 168.135 ;
        RECT 80.115 167.635 80.340 167.675 ;
        RECT 79.185 167.505 79.435 167.595 ;
        RECT 78.640 167.255 79.435 167.505 ;
        RECT 77.235 166.905 79.025 167.075 ;
        RECT 76.895 166.035 77.170 166.735 ;
        RECT 77.340 166.610 78.055 166.905 ;
        RECT 78.275 166.545 78.605 166.735 ;
        RECT 77.380 165.865 77.595 166.410 ;
        RECT 77.765 166.035 78.240 166.375 ;
        RECT 78.410 166.370 78.605 166.545 ;
        RECT 78.775 166.540 79.025 166.905 ;
        RECT 78.410 165.865 79.025 166.370 ;
        RECT 79.265 166.035 79.435 167.255 ;
        RECT 79.605 166.545 79.945 167.425 ;
        RECT 80.115 167.055 80.285 167.635 ;
        RECT 81.005 167.505 81.205 167.675 ;
        RECT 82.080 167.505 82.250 167.965 ;
        RECT 80.455 167.175 81.205 167.505 ;
        RECT 81.375 167.175 82.250 167.505 ;
        RECT 80.115 167.005 80.330 167.055 ;
        RECT 80.115 166.925 80.505 167.005 ;
        RECT 79.685 165.865 79.945 166.375 ;
        RECT 80.175 166.080 80.505 166.925 ;
        RECT 81.015 166.970 81.205 167.175 ;
        RECT 80.675 165.865 80.845 166.875 ;
        RECT 81.015 166.595 81.910 166.970 ;
        RECT 81.015 166.035 81.355 166.595 ;
        RECT 81.585 165.865 81.900 166.365 ;
        RECT 82.080 166.335 82.250 167.175 ;
        RECT 82.420 167.465 82.885 167.795 ;
        RECT 83.270 167.735 83.440 167.965 ;
        RECT 83.620 167.915 83.990 168.415 ;
        RECT 84.310 167.965 84.985 168.135 ;
        RECT 85.180 167.965 85.515 168.135 ;
        RECT 82.420 166.505 82.740 167.465 ;
        RECT 83.270 167.435 84.100 167.735 ;
        RECT 82.910 166.535 83.100 167.255 ;
        RECT 83.270 166.365 83.440 167.435 ;
        RECT 83.900 167.405 84.100 167.435 ;
        RECT 83.610 167.185 83.780 167.255 ;
        RECT 84.310 167.185 84.480 167.965 ;
        RECT 85.345 167.825 85.515 167.965 ;
        RECT 85.685 167.955 85.935 168.415 ;
        RECT 83.610 167.015 84.480 167.185 ;
        RECT 84.650 167.545 85.175 167.765 ;
        RECT 85.345 167.695 85.570 167.825 ;
        RECT 83.610 166.925 84.120 167.015 ;
        RECT 82.080 166.165 82.965 166.335 ;
        RECT 83.190 166.035 83.440 166.365 ;
        RECT 83.610 165.865 83.780 166.665 ;
        RECT 83.950 166.310 84.120 166.925 ;
        RECT 84.650 166.845 84.820 167.545 ;
        RECT 84.290 166.480 84.820 166.845 ;
        RECT 84.990 166.780 85.230 167.375 ;
        RECT 85.400 166.590 85.570 167.695 ;
        RECT 85.740 166.835 86.020 167.785 ;
        RECT 85.265 166.460 85.570 166.590 ;
        RECT 83.950 166.140 85.055 166.310 ;
        RECT 85.265 166.035 85.515 166.460 ;
        RECT 85.685 165.865 85.950 166.325 ;
        RECT 86.190 166.035 86.375 168.155 ;
        RECT 86.545 168.035 86.875 168.415 ;
        RECT 87.045 167.865 87.215 168.155 ;
        RECT 86.550 167.695 87.215 167.865 ;
        RECT 86.550 166.705 86.780 167.695 ;
        RECT 87.475 167.645 90.065 168.415 ;
        RECT 90.695 167.690 90.985 168.415 ;
        RECT 92.125 167.760 92.455 168.195 ;
        RECT 92.625 167.805 92.795 168.415 ;
        RECT 92.075 167.675 92.455 167.760 ;
        RECT 92.965 167.675 93.295 168.200 ;
        RECT 93.555 167.885 93.765 168.415 ;
        RECT 94.040 167.965 94.825 168.135 ;
        RECT 94.995 167.965 95.400 168.135 ;
        RECT 86.950 166.875 87.300 167.525 ;
        RECT 87.475 167.125 88.685 167.645 ;
        RECT 92.075 167.635 92.300 167.675 ;
        RECT 88.855 166.955 90.065 167.475 ;
        RECT 92.075 167.055 92.245 167.635 ;
        RECT 92.965 167.505 93.165 167.675 ;
        RECT 94.040 167.505 94.210 167.965 ;
        RECT 92.415 167.175 93.165 167.505 ;
        RECT 93.335 167.175 94.210 167.505 ;
        RECT 86.550 166.535 87.215 166.705 ;
        RECT 86.545 165.865 86.875 166.365 ;
        RECT 87.045 166.035 87.215 166.535 ;
        RECT 87.475 165.865 90.065 166.955 ;
        RECT 90.695 165.865 90.985 167.030 ;
        RECT 92.075 167.005 92.290 167.055 ;
        RECT 92.075 166.925 92.465 167.005 ;
        RECT 92.135 166.080 92.465 166.925 ;
        RECT 92.975 166.970 93.165 167.175 ;
        RECT 92.635 165.865 92.805 166.875 ;
        RECT 92.975 166.595 93.870 166.970 ;
        RECT 92.975 166.035 93.315 166.595 ;
        RECT 93.545 165.865 93.860 166.365 ;
        RECT 94.040 166.335 94.210 167.175 ;
        RECT 94.380 167.465 94.845 167.795 ;
        RECT 95.230 167.735 95.400 167.965 ;
        RECT 95.580 167.915 95.950 168.415 ;
        RECT 96.270 167.965 96.945 168.135 ;
        RECT 97.140 167.965 97.475 168.135 ;
        RECT 94.380 166.505 94.700 167.465 ;
        RECT 95.230 167.435 96.060 167.735 ;
        RECT 94.870 166.535 95.060 167.255 ;
        RECT 95.230 166.365 95.400 167.435 ;
        RECT 95.860 167.405 96.060 167.435 ;
        RECT 95.570 167.185 95.740 167.255 ;
        RECT 96.270 167.185 96.440 167.965 ;
        RECT 97.305 167.825 97.475 167.965 ;
        RECT 97.645 167.955 97.895 168.415 ;
        RECT 95.570 167.015 96.440 167.185 ;
        RECT 96.610 167.545 97.135 167.765 ;
        RECT 97.305 167.695 97.530 167.825 ;
        RECT 95.570 166.925 96.080 167.015 ;
        RECT 94.040 166.165 94.925 166.335 ;
        RECT 95.150 166.035 95.400 166.365 ;
        RECT 95.570 165.865 95.740 166.665 ;
        RECT 95.910 166.310 96.080 166.925 ;
        RECT 96.610 166.845 96.780 167.545 ;
        RECT 96.250 166.480 96.780 166.845 ;
        RECT 96.950 166.780 97.190 167.375 ;
        RECT 97.360 166.590 97.530 167.695 ;
        RECT 97.700 166.835 97.980 167.785 ;
        RECT 97.225 166.460 97.530 166.590 ;
        RECT 95.910 166.140 97.015 166.310 ;
        RECT 97.225 166.035 97.475 166.460 ;
        RECT 97.645 165.865 97.910 166.325 ;
        RECT 98.150 166.035 98.335 168.155 ;
        RECT 98.505 168.035 98.835 168.415 ;
        RECT 99.005 167.865 99.175 168.155 ;
        RECT 98.510 167.695 99.175 167.865 ;
        RECT 98.510 166.705 98.740 167.695 ;
        RECT 98.910 166.875 99.260 167.525 ;
        RECT 98.510 166.535 99.175 166.705 ;
        RECT 98.505 165.865 98.835 166.365 ;
        RECT 99.005 166.035 99.175 166.535 ;
        RECT 99.435 166.035 99.715 168.135 ;
        RECT 99.945 167.955 100.115 168.415 ;
        RECT 100.385 168.025 101.635 168.205 ;
        RECT 100.770 167.785 101.135 167.855 ;
        RECT 99.885 167.605 101.135 167.785 ;
        RECT 101.305 167.805 101.635 168.025 ;
        RECT 101.805 167.975 101.975 168.415 ;
        RECT 102.145 167.805 102.485 168.220 ;
        RECT 101.305 167.635 102.485 167.805 ;
        RECT 102.655 167.645 104.325 168.415 ;
        RECT 105.155 167.785 105.485 168.145 ;
        RECT 106.105 167.955 106.355 168.415 ;
        RECT 106.525 167.955 107.085 168.245 ;
        RECT 99.885 167.005 100.160 167.605 ;
        RECT 100.330 167.175 100.685 167.425 ;
        RECT 100.880 167.395 101.345 167.425 ;
        RECT 100.875 167.225 101.345 167.395 ;
        RECT 100.880 167.175 101.345 167.225 ;
        RECT 101.515 167.175 101.845 167.425 ;
        RECT 102.020 167.225 102.485 167.425 ;
        RECT 101.665 167.055 101.845 167.175 ;
        RECT 102.655 167.125 103.405 167.645 ;
        RECT 105.155 167.595 106.545 167.785 ;
        RECT 106.375 167.505 106.545 167.595 ;
        RECT 99.885 166.795 101.495 167.005 ;
        RECT 101.665 166.885 101.995 167.055 ;
        RECT 101.085 166.695 101.495 166.795 ;
        RECT 99.905 165.865 100.690 166.625 ;
        RECT 101.085 166.035 101.470 166.695 ;
        RECT 101.795 166.095 101.995 166.885 ;
        RECT 102.165 165.865 102.485 167.045 ;
        RECT 103.575 166.955 104.325 167.475 ;
        RECT 102.655 165.865 104.325 166.955 ;
        RECT 104.970 167.175 105.645 167.425 ;
        RECT 105.865 167.175 106.205 167.425 ;
        RECT 106.375 167.175 106.665 167.505 ;
        RECT 104.970 166.815 105.235 167.175 ;
        RECT 106.375 166.925 106.545 167.175 ;
        RECT 105.605 166.755 106.545 166.925 ;
        RECT 105.155 165.865 105.435 166.535 ;
        RECT 105.605 166.205 105.905 166.755 ;
        RECT 106.835 166.585 107.085 167.955 ;
        RECT 107.315 167.595 107.525 168.415 ;
        RECT 107.695 167.615 108.025 168.245 ;
        RECT 107.695 167.015 107.945 167.615 ;
        RECT 108.195 167.595 108.425 168.415 ;
        RECT 108.635 167.615 109.330 168.245 ;
        RECT 109.535 167.615 109.845 168.415 ;
        RECT 109.155 167.565 109.330 167.615 ;
        RECT 110.025 167.605 110.295 168.415 ;
        RECT 110.465 167.605 110.795 168.245 ;
        RECT 110.965 167.605 111.205 168.415 ;
        RECT 111.395 167.615 112.090 168.245 ;
        RECT 112.295 167.615 112.605 168.415 ;
        RECT 113.975 167.785 114.355 168.235 ;
        RECT 108.115 167.175 108.445 167.425 ;
        RECT 108.655 167.175 108.990 167.425 ;
        RECT 109.160 167.015 109.330 167.565 ;
        RECT 109.500 167.175 109.835 167.445 ;
        RECT 110.015 167.175 110.365 167.425 ;
        RECT 106.105 165.865 106.435 166.585 ;
        RECT 106.625 166.035 107.085 166.585 ;
        RECT 107.315 165.865 107.525 167.005 ;
        RECT 107.695 166.035 108.025 167.015 ;
        RECT 108.195 165.865 108.425 167.005 ;
        RECT 108.635 165.865 108.895 167.005 ;
        RECT 109.065 166.035 109.395 167.015 ;
        RECT 110.535 167.005 110.705 167.605 ;
        RECT 110.875 167.175 111.225 167.425 ;
        RECT 111.415 167.175 111.750 167.425 ;
        RECT 111.920 167.055 112.090 167.615 ;
        RECT 112.260 167.175 112.595 167.445 ;
        RECT 111.915 167.015 112.090 167.055 ;
        RECT 109.565 165.865 109.845 167.005 ;
        RECT 110.025 165.865 110.355 167.005 ;
        RECT 110.535 166.835 111.215 167.005 ;
        RECT 110.885 166.050 111.215 166.835 ;
        RECT 111.395 165.865 111.655 167.005 ;
        RECT 111.825 166.035 112.155 167.015 ;
        RECT 112.325 165.865 112.605 167.005 ;
        RECT 113.715 166.835 113.945 167.525 ;
        RECT 114.125 167.335 114.355 167.785 ;
        RECT 114.535 167.635 114.765 168.415 ;
        RECT 114.945 167.705 115.375 168.235 ;
        RECT 114.945 167.455 115.190 167.705 ;
        RECT 115.555 167.505 115.765 168.125 ;
        RECT 115.935 167.685 116.265 168.415 ;
        RECT 116.455 167.690 116.745 168.415 ;
        RECT 116.930 167.845 117.185 168.195 ;
        RECT 117.355 168.015 117.685 168.415 ;
        RECT 117.855 167.845 118.025 168.195 ;
        RECT 118.195 168.015 118.575 168.415 ;
        RECT 116.930 167.675 118.595 167.845 ;
        RECT 118.765 167.740 119.040 168.085 ;
        RECT 119.275 167.955 119.520 168.415 ;
        RECT 118.425 167.505 118.595 167.675 ;
        RECT 114.125 166.655 114.465 167.335 ;
        RECT 113.705 166.455 114.465 166.655 ;
        RECT 114.655 167.155 115.190 167.455 ;
        RECT 115.370 167.155 115.765 167.505 ;
        RECT 115.960 167.155 116.250 167.505 ;
        RECT 116.915 167.175 117.260 167.505 ;
        RECT 117.430 167.175 118.255 167.505 ;
        RECT 118.425 167.175 118.700 167.505 ;
        RECT 113.705 166.065 113.965 166.455 ;
        RECT 114.135 165.865 114.465 166.275 ;
        RECT 114.655 166.045 114.985 167.155 ;
        RECT 115.155 166.775 116.195 166.975 ;
        RECT 115.155 166.045 115.345 166.775 ;
        RECT 115.515 165.865 115.845 166.595 ;
        RECT 116.025 166.045 116.195 166.775 ;
        RECT 116.455 165.865 116.745 167.030 ;
        RECT 116.935 166.715 117.260 167.005 ;
        RECT 117.430 166.885 117.625 167.175 ;
        RECT 118.425 167.005 118.595 167.175 ;
        RECT 118.870 167.005 119.040 167.740 ;
        RECT 119.215 167.175 119.530 167.785 ;
        RECT 119.700 167.425 119.950 168.235 ;
        RECT 120.120 167.890 120.380 168.415 ;
        RECT 120.550 167.765 120.810 168.220 ;
        RECT 120.980 167.935 121.240 168.415 ;
        RECT 121.410 167.765 121.670 168.220 ;
        RECT 121.840 167.935 122.100 168.415 ;
        RECT 122.270 167.765 122.530 168.220 ;
        RECT 122.700 167.935 122.960 168.415 ;
        RECT 123.130 167.765 123.390 168.220 ;
        RECT 123.560 167.935 123.860 168.415 ;
        RECT 120.550 167.595 123.860 167.765 ;
        RECT 124.275 167.615 124.970 168.245 ;
        RECT 125.175 167.615 125.485 168.415 ;
        RECT 126.665 167.865 126.835 168.155 ;
        RECT 127.005 168.035 127.335 168.415 ;
        RECT 126.665 167.695 127.330 167.865 ;
        RECT 119.700 167.175 122.720 167.425 ;
        RECT 117.935 166.835 118.595 167.005 ;
        RECT 117.935 166.715 118.105 166.835 ;
        RECT 116.935 166.545 118.105 166.715 ;
        RECT 116.915 166.085 118.105 166.375 ;
        RECT 118.275 165.865 118.555 166.665 ;
        RECT 118.765 166.035 119.040 167.005 ;
        RECT 119.225 165.865 119.520 166.975 ;
        RECT 119.700 166.040 119.950 167.175 ;
        RECT 122.890 167.005 123.860 167.595 ;
        RECT 124.295 167.175 124.630 167.425 ;
        RECT 124.800 167.015 124.970 167.615 ;
        RECT 125.140 167.175 125.475 167.445 ;
        RECT 120.120 165.865 120.380 166.975 ;
        RECT 120.550 166.765 123.860 167.005 ;
        RECT 120.550 166.040 120.810 166.765 ;
        RECT 120.980 165.865 121.240 166.595 ;
        RECT 121.410 166.040 121.670 166.765 ;
        RECT 121.840 165.865 122.100 166.595 ;
        RECT 122.270 166.040 122.530 166.765 ;
        RECT 122.700 165.865 122.960 166.595 ;
        RECT 123.130 166.040 123.390 166.765 ;
        RECT 123.560 165.865 123.855 166.595 ;
        RECT 124.275 165.865 124.535 167.005 ;
        RECT 124.705 166.035 125.035 167.015 ;
        RECT 125.205 165.865 125.485 167.005 ;
        RECT 126.580 166.875 126.930 167.525 ;
        RECT 127.100 166.705 127.330 167.695 ;
        RECT 126.665 166.535 127.330 166.705 ;
        RECT 126.665 166.035 126.835 166.535 ;
        RECT 127.005 165.865 127.335 166.365 ;
        RECT 127.505 166.035 127.690 168.155 ;
        RECT 127.945 167.955 128.195 168.415 ;
        RECT 128.365 167.965 128.700 168.135 ;
        RECT 128.895 167.965 129.570 168.135 ;
        RECT 128.365 167.825 128.535 167.965 ;
        RECT 127.860 166.835 128.140 167.785 ;
        RECT 128.310 167.695 128.535 167.825 ;
        RECT 128.310 166.590 128.480 167.695 ;
        RECT 128.705 167.545 129.230 167.765 ;
        RECT 128.650 166.780 128.890 167.375 ;
        RECT 129.060 166.845 129.230 167.545 ;
        RECT 129.400 167.185 129.570 167.965 ;
        RECT 129.890 167.915 130.260 168.415 ;
        RECT 130.440 167.965 130.845 168.135 ;
        RECT 131.015 167.965 131.800 168.135 ;
        RECT 130.440 167.735 130.610 167.965 ;
        RECT 129.780 167.435 130.610 167.735 ;
        RECT 130.995 167.465 131.460 167.795 ;
        RECT 129.780 167.405 129.980 167.435 ;
        RECT 130.100 167.185 130.270 167.255 ;
        RECT 129.400 167.015 130.270 167.185 ;
        RECT 129.760 166.925 130.270 167.015 ;
        RECT 128.310 166.460 128.615 166.590 ;
        RECT 129.060 166.480 129.590 166.845 ;
        RECT 127.930 165.865 128.195 166.325 ;
        RECT 128.365 166.035 128.615 166.460 ;
        RECT 129.760 166.310 129.930 166.925 ;
        RECT 128.825 166.140 129.930 166.310 ;
        RECT 130.100 165.865 130.270 166.665 ;
        RECT 130.440 166.365 130.610 167.435 ;
        RECT 130.780 166.535 130.970 167.255 ;
        RECT 131.140 166.505 131.460 167.465 ;
        RECT 131.630 167.505 131.800 167.965 ;
        RECT 132.075 167.885 132.285 168.415 ;
        RECT 132.545 167.675 132.875 168.200 ;
        RECT 133.045 167.805 133.215 168.415 ;
        RECT 133.385 167.760 133.715 168.195 ;
        RECT 134.025 167.865 134.195 168.245 ;
        RECT 134.410 168.035 134.740 168.415 ;
        RECT 133.385 167.675 133.765 167.760 ;
        RECT 134.025 167.695 134.740 167.865 ;
        RECT 132.675 167.505 132.875 167.675 ;
        RECT 133.540 167.635 133.765 167.675 ;
        RECT 131.630 167.175 132.505 167.505 ;
        RECT 132.675 167.175 133.425 167.505 ;
        RECT 130.440 166.035 130.690 166.365 ;
        RECT 131.630 166.335 131.800 167.175 ;
        RECT 132.675 166.970 132.865 167.175 ;
        RECT 133.595 167.055 133.765 167.635 ;
        RECT 133.935 167.145 134.290 167.515 ;
        RECT 134.570 167.505 134.740 167.695 ;
        RECT 134.910 167.670 135.165 168.245 ;
        RECT 134.570 167.175 134.825 167.505 ;
        RECT 133.550 167.005 133.765 167.055 ;
        RECT 131.970 166.595 132.865 166.970 ;
        RECT 133.375 166.925 133.765 167.005 ;
        RECT 134.570 166.965 134.740 167.175 ;
        RECT 130.915 166.165 131.800 166.335 ;
        RECT 131.980 165.865 132.295 166.365 ;
        RECT 132.525 166.035 132.865 166.595 ;
        RECT 133.035 165.865 133.205 166.875 ;
        RECT 133.375 166.080 133.705 166.925 ;
        RECT 134.025 166.795 134.740 166.965 ;
        RECT 134.995 166.940 135.165 167.670 ;
        RECT 135.340 167.575 135.600 168.415 ;
        RECT 135.865 167.865 136.035 168.245 ;
        RECT 136.250 168.035 136.580 168.415 ;
        RECT 135.865 167.695 136.580 167.865 ;
        RECT 135.775 167.145 136.130 167.515 ;
        RECT 136.410 167.505 136.580 167.695 ;
        RECT 136.750 167.670 137.005 168.245 ;
        RECT 136.410 167.175 136.665 167.505 ;
        RECT 134.025 166.035 134.195 166.795 ;
        RECT 134.410 165.865 134.740 166.625 ;
        RECT 134.910 166.035 135.165 166.940 ;
        RECT 135.340 165.865 135.600 167.015 ;
        RECT 136.410 166.965 136.580 167.175 ;
        RECT 135.865 166.795 136.580 166.965 ;
        RECT 136.835 166.940 137.005 167.670 ;
        RECT 137.180 167.575 137.440 168.415 ;
        RECT 137.615 167.665 138.825 168.415 ;
        RECT 135.865 166.035 136.035 166.795 ;
        RECT 136.250 165.865 136.580 166.625 ;
        RECT 136.750 166.035 137.005 166.940 ;
        RECT 137.180 165.865 137.440 167.015 ;
        RECT 137.615 166.955 138.135 167.495 ;
        RECT 138.305 167.125 138.825 167.665 ;
        RECT 137.615 165.865 138.825 166.955 ;
        RECT 13.330 165.695 138.910 165.865 ;
        RECT 13.415 164.605 14.625 165.695 ;
        RECT 15.805 165.025 15.975 165.525 ;
        RECT 16.145 165.195 16.475 165.695 ;
        RECT 15.805 164.855 16.470 165.025 ;
        RECT 13.415 163.895 13.935 164.435 ;
        RECT 14.105 164.065 14.625 164.605 ;
        RECT 15.720 164.035 16.070 164.685 ;
        RECT 13.415 163.145 14.625 163.895 ;
        RECT 16.240 163.865 16.470 164.855 ;
        RECT 15.805 163.695 16.470 163.865 ;
        RECT 15.805 163.405 15.975 163.695 ;
        RECT 16.145 163.145 16.475 163.525 ;
        RECT 16.645 163.405 16.830 165.525 ;
        RECT 17.070 165.235 17.335 165.695 ;
        RECT 17.505 165.100 17.755 165.525 ;
        RECT 17.965 165.250 19.070 165.420 ;
        RECT 17.450 164.970 17.755 165.100 ;
        RECT 17.000 163.775 17.280 164.725 ;
        RECT 17.450 163.865 17.620 164.970 ;
        RECT 17.790 164.185 18.030 164.780 ;
        RECT 18.200 164.715 18.730 165.080 ;
        RECT 18.200 164.015 18.370 164.715 ;
        RECT 18.900 164.635 19.070 165.250 ;
        RECT 19.240 164.895 19.410 165.695 ;
        RECT 19.580 165.195 19.830 165.525 ;
        RECT 20.055 165.225 20.940 165.395 ;
        RECT 18.900 164.545 19.410 164.635 ;
        RECT 17.450 163.735 17.675 163.865 ;
        RECT 17.845 163.795 18.370 164.015 ;
        RECT 18.540 164.375 19.410 164.545 ;
        RECT 17.085 163.145 17.335 163.605 ;
        RECT 17.505 163.595 17.675 163.735 ;
        RECT 18.540 163.595 18.710 164.375 ;
        RECT 19.240 164.305 19.410 164.375 ;
        RECT 18.920 164.125 19.120 164.155 ;
        RECT 19.580 164.125 19.750 165.195 ;
        RECT 19.920 164.305 20.110 165.025 ;
        RECT 18.920 163.825 19.750 164.125 ;
        RECT 20.280 164.095 20.600 165.055 ;
        RECT 17.505 163.425 17.840 163.595 ;
        RECT 18.035 163.425 18.710 163.595 ;
        RECT 19.030 163.145 19.400 163.645 ;
        RECT 19.580 163.595 19.750 163.825 ;
        RECT 20.135 163.765 20.600 164.095 ;
        RECT 20.770 164.385 20.940 165.225 ;
        RECT 21.120 165.195 21.435 165.695 ;
        RECT 21.665 164.965 22.005 165.525 ;
        RECT 21.110 164.590 22.005 164.965 ;
        RECT 22.175 164.685 22.345 165.695 ;
        RECT 21.815 164.385 22.005 164.590 ;
        RECT 22.515 164.635 22.845 165.480 ;
        RECT 22.515 164.555 22.905 164.635 ;
        RECT 23.075 164.605 25.665 165.695 ;
        RECT 22.690 164.505 22.905 164.555 ;
        RECT 20.770 164.055 21.645 164.385 ;
        RECT 21.815 164.055 22.565 164.385 ;
        RECT 20.770 163.595 20.940 164.055 ;
        RECT 21.815 163.885 22.015 164.055 ;
        RECT 22.735 163.925 22.905 164.505 ;
        RECT 22.680 163.885 22.905 163.925 ;
        RECT 19.580 163.425 19.985 163.595 ;
        RECT 20.155 163.425 20.940 163.595 ;
        RECT 21.215 163.145 21.425 163.675 ;
        RECT 21.685 163.360 22.015 163.885 ;
        RECT 22.525 163.800 22.905 163.885 ;
        RECT 23.075 163.915 24.285 164.435 ;
        RECT 24.455 164.085 25.665 164.605 ;
        RECT 26.295 164.530 26.585 165.695 ;
        RECT 26.810 164.825 27.095 165.695 ;
        RECT 27.265 165.065 27.525 165.525 ;
        RECT 27.700 165.235 27.955 165.695 ;
        RECT 28.125 165.065 28.385 165.525 ;
        RECT 27.265 164.895 28.385 165.065 ;
        RECT 28.555 164.895 28.865 165.695 ;
        RECT 27.265 164.645 27.525 164.895 ;
        RECT 29.035 164.725 29.345 165.525 ;
        RECT 29.515 165.260 34.860 165.695 ;
        RECT 26.770 164.475 27.525 164.645 ;
        RECT 28.315 164.555 29.345 164.725 ;
        RECT 26.770 163.965 27.175 164.475 ;
        RECT 28.315 164.305 28.485 164.555 ;
        RECT 27.345 164.135 28.485 164.305 ;
        RECT 22.185 163.145 22.355 163.755 ;
        RECT 22.525 163.365 22.855 163.800 ;
        RECT 23.075 163.145 25.665 163.915 ;
        RECT 26.295 163.145 26.585 163.870 ;
        RECT 26.770 163.795 28.420 163.965 ;
        RECT 28.655 163.815 29.005 164.385 ;
        RECT 26.815 163.145 27.095 163.625 ;
        RECT 27.265 163.405 27.525 163.795 ;
        RECT 27.700 163.145 27.955 163.625 ;
        RECT 28.125 163.405 28.420 163.795 ;
        RECT 29.175 163.645 29.345 164.555 ;
        RECT 31.100 163.690 31.440 164.520 ;
        RECT 32.920 164.010 33.270 165.260 ;
        RECT 35.035 164.090 35.315 165.525 ;
        RECT 35.485 164.920 36.195 165.695 ;
        RECT 36.365 164.750 36.695 165.525 ;
        RECT 35.545 164.535 36.695 164.750 ;
        RECT 28.600 163.145 28.875 163.625 ;
        RECT 29.045 163.315 29.345 163.645 ;
        RECT 29.515 163.145 34.860 163.690 ;
        RECT 35.035 163.315 35.375 164.090 ;
        RECT 35.545 163.965 35.830 164.535 ;
        RECT 36.015 164.135 36.485 164.365 ;
        RECT 36.890 164.335 37.105 165.450 ;
        RECT 37.285 164.975 37.615 165.695 ;
        RECT 37.395 164.335 37.625 164.675 ;
        RECT 37.795 164.605 39.465 165.695 ;
        RECT 36.655 164.155 37.105 164.335 ;
        RECT 36.655 164.135 36.985 164.155 ;
        RECT 37.295 164.135 37.625 164.335 ;
        RECT 35.545 163.775 36.255 163.965 ;
        RECT 35.955 163.635 36.255 163.775 ;
        RECT 36.445 163.775 37.625 163.965 ;
        RECT 36.445 163.695 36.775 163.775 ;
        RECT 35.955 163.625 36.270 163.635 ;
        RECT 35.955 163.615 36.280 163.625 ;
        RECT 35.955 163.610 36.290 163.615 ;
        RECT 35.545 163.145 35.715 163.605 ;
        RECT 35.955 163.600 36.295 163.610 ;
        RECT 35.955 163.595 36.300 163.600 ;
        RECT 35.955 163.585 36.305 163.595 ;
        RECT 35.955 163.580 36.310 163.585 ;
        RECT 35.955 163.315 36.315 163.580 ;
        RECT 36.945 163.145 37.115 163.605 ;
        RECT 37.285 163.315 37.625 163.775 ;
        RECT 37.795 163.915 38.545 164.435 ;
        RECT 38.715 164.085 39.465 164.605 ;
        RECT 39.635 164.555 39.905 165.525 ;
        RECT 40.115 164.895 40.395 165.695 ;
        RECT 40.565 165.185 42.220 165.475 ;
        RECT 40.630 164.845 42.220 165.015 ;
        RECT 42.405 164.895 42.735 165.695 ;
        RECT 42.915 165.355 44.345 165.525 ;
        RECT 40.630 164.725 40.800 164.845 ;
        RECT 40.075 164.555 40.800 164.725 ;
        RECT 37.795 163.145 39.465 163.915 ;
        RECT 39.635 163.820 39.805 164.555 ;
        RECT 40.075 164.385 40.245 164.555 ;
        RECT 39.975 164.055 40.245 164.385 ;
        RECT 40.415 164.055 40.820 164.385 ;
        RECT 40.990 164.055 41.700 164.675 ;
        RECT 41.900 164.555 42.220 164.845 ;
        RECT 42.915 164.725 43.165 165.355 ;
        RECT 42.395 164.555 43.165 164.725 ;
        RECT 40.075 163.885 40.245 164.055 ;
        RECT 39.635 163.475 39.905 163.820 ;
        RECT 40.075 163.715 41.685 163.885 ;
        RECT 41.870 163.815 42.220 164.385 ;
        RECT 42.395 163.885 42.565 164.555 ;
        RECT 42.735 164.055 43.140 164.385 ;
        RECT 43.355 164.055 43.605 165.185 ;
        RECT 43.805 164.385 44.005 165.185 ;
        RECT 44.175 164.675 44.345 165.355 ;
        RECT 44.515 164.845 44.830 165.695 ;
        RECT 45.005 164.895 45.445 165.525 ;
        RECT 44.175 164.505 44.965 164.675 ;
        RECT 43.805 164.055 44.050 164.385 ;
        RECT 44.235 164.055 44.625 164.335 ;
        RECT 44.795 164.055 44.965 164.505 ;
        RECT 45.135 163.885 45.445 164.895 ;
        RECT 45.625 164.725 45.955 165.510 ;
        RECT 45.625 164.555 46.305 164.725 ;
        RECT 46.485 164.555 46.815 165.695 ;
        RECT 48.000 165.075 48.175 165.525 ;
        RECT 48.345 165.255 48.675 165.695 ;
        RECT 48.980 165.105 49.150 165.525 ;
        RECT 49.385 165.285 50.055 165.695 ;
        RECT 50.270 165.105 50.440 165.525 ;
        RECT 50.640 165.285 50.970 165.695 ;
        RECT 48.000 164.905 48.630 165.075 ;
        RECT 45.615 164.135 45.965 164.385 ;
        RECT 46.135 163.955 46.305 164.555 ;
        RECT 46.475 164.135 46.825 164.385 ;
        RECT 47.915 164.055 48.280 164.735 ;
        RECT 48.460 164.385 48.630 164.905 ;
        RECT 48.980 164.935 50.995 165.105 ;
        RECT 48.460 164.055 48.810 164.385 ;
        RECT 40.095 163.145 40.475 163.545 ;
        RECT 40.645 163.365 40.815 163.715 ;
        RECT 40.985 163.145 41.315 163.545 ;
        RECT 41.515 163.365 41.685 163.715 ;
        RECT 41.885 163.145 42.215 163.645 ;
        RECT 42.395 163.315 42.885 163.885 ;
        RECT 43.055 163.715 44.215 163.885 ;
        RECT 43.055 163.315 43.285 163.715 ;
        RECT 43.455 163.145 43.875 163.545 ;
        RECT 44.045 163.315 44.215 163.715 ;
        RECT 44.385 163.145 44.835 163.885 ;
        RECT 45.005 163.325 45.445 163.885 ;
        RECT 45.635 163.145 45.875 163.955 ;
        RECT 46.045 163.315 46.375 163.955 ;
        RECT 46.545 163.145 46.815 163.955 ;
        RECT 48.460 163.885 48.630 164.055 ;
        RECT 48.000 163.715 48.630 163.885 ;
        RECT 48.000 163.315 48.175 163.715 ;
        RECT 48.980 163.645 49.150 164.935 ;
        RECT 48.345 163.145 48.675 163.525 ;
        RECT 48.920 163.315 49.150 163.645 ;
        RECT 49.350 163.480 49.630 164.755 ;
        RECT 49.855 164.675 50.125 164.755 ;
        RECT 49.815 164.505 50.125 164.675 ;
        RECT 49.855 163.480 50.125 164.505 ;
        RECT 50.315 163.725 50.655 164.755 ;
        RECT 50.825 164.385 50.995 164.935 ;
        RECT 51.165 164.555 51.425 165.525 ;
        RECT 50.825 164.055 51.085 164.385 ;
        RECT 51.255 163.865 51.425 164.555 ;
        RECT 52.055 164.530 52.345 165.695 ;
        RECT 52.575 164.635 52.905 165.480 ;
        RECT 53.075 164.685 53.245 165.695 ;
        RECT 53.415 164.965 53.755 165.525 ;
        RECT 53.985 165.195 54.300 165.695 ;
        RECT 54.480 165.225 55.365 165.395 ;
        RECT 52.515 164.555 52.905 164.635 ;
        RECT 53.415 164.590 54.310 164.965 ;
        RECT 52.515 164.505 52.730 164.555 ;
        RECT 52.515 163.925 52.685 164.505 ;
        RECT 53.415 164.385 53.605 164.590 ;
        RECT 54.480 164.385 54.650 165.225 ;
        RECT 55.590 165.195 55.840 165.525 ;
        RECT 52.855 164.055 53.605 164.385 ;
        RECT 53.775 164.055 54.650 164.385 ;
        RECT 52.515 163.885 52.740 163.925 ;
        RECT 53.405 163.885 53.605 164.055 ;
        RECT 50.585 163.145 50.915 163.525 ;
        RECT 51.085 163.400 51.425 163.865 ;
        RECT 51.085 163.355 51.420 163.400 ;
        RECT 52.055 163.145 52.345 163.870 ;
        RECT 52.515 163.800 52.895 163.885 ;
        RECT 52.565 163.365 52.895 163.800 ;
        RECT 53.065 163.145 53.235 163.755 ;
        RECT 53.405 163.360 53.735 163.885 ;
        RECT 53.995 163.145 54.205 163.675 ;
        RECT 54.480 163.595 54.650 164.055 ;
        RECT 54.820 164.095 55.140 165.055 ;
        RECT 55.310 164.305 55.500 165.025 ;
        RECT 55.670 164.125 55.840 165.195 ;
        RECT 56.010 164.895 56.180 165.695 ;
        RECT 56.350 165.250 57.455 165.420 ;
        RECT 56.350 164.635 56.520 165.250 ;
        RECT 57.665 165.100 57.915 165.525 ;
        RECT 58.085 165.235 58.350 165.695 ;
        RECT 56.690 164.715 57.220 165.080 ;
        RECT 57.665 164.970 57.970 165.100 ;
        RECT 56.010 164.545 56.520 164.635 ;
        RECT 56.010 164.375 56.880 164.545 ;
        RECT 56.010 164.305 56.180 164.375 ;
        RECT 56.300 164.125 56.500 164.155 ;
        RECT 54.820 163.765 55.285 164.095 ;
        RECT 55.670 163.825 56.500 164.125 ;
        RECT 55.670 163.595 55.840 163.825 ;
        RECT 54.480 163.425 55.265 163.595 ;
        RECT 55.435 163.425 55.840 163.595 ;
        RECT 56.020 163.145 56.390 163.645 ;
        RECT 56.710 163.595 56.880 164.375 ;
        RECT 57.050 164.015 57.220 164.715 ;
        RECT 57.390 164.185 57.630 164.780 ;
        RECT 57.050 163.795 57.575 164.015 ;
        RECT 57.800 163.865 57.970 164.970 ;
        RECT 57.745 163.735 57.970 163.865 ;
        RECT 58.140 163.775 58.420 164.725 ;
        RECT 57.745 163.595 57.915 163.735 ;
        RECT 56.710 163.425 57.385 163.595 ;
        RECT 57.580 163.425 57.915 163.595 ;
        RECT 58.085 163.145 58.335 163.605 ;
        RECT 58.590 163.405 58.775 165.525 ;
        RECT 58.945 165.195 59.275 165.695 ;
        RECT 59.445 165.025 59.615 165.525 ;
        RECT 58.950 164.855 59.615 165.025 ;
        RECT 58.950 163.865 59.180 164.855 ;
        RECT 60.335 164.725 60.645 165.525 ;
        RECT 60.815 164.895 61.125 165.695 ;
        RECT 61.295 165.065 61.555 165.525 ;
        RECT 61.725 165.235 61.980 165.695 ;
        RECT 62.155 165.065 62.415 165.525 ;
        RECT 61.295 164.895 62.415 165.065 ;
        RECT 59.350 164.035 59.700 164.685 ;
        RECT 60.335 164.555 61.365 164.725 ;
        RECT 58.950 163.695 59.615 163.865 ;
        RECT 58.945 163.145 59.275 163.525 ;
        RECT 59.445 163.405 59.615 163.695 ;
        RECT 60.335 163.645 60.505 164.555 ;
        RECT 60.675 163.815 61.025 164.385 ;
        RECT 61.195 164.305 61.365 164.555 ;
        RECT 62.155 164.645 62.415 164.895 ;
        RECT 62.585 164.825 62.870 165.695 ;
        RECT 62.155 164.475 62.910 164.645 ;
        RECT 63.105 164.585 63.400 165.695 ;
        RECT 61.195 164.135 62.335 164.305 ;
        RECT 62.505 163.965 62.910 164.475 ;
        RECT 63.580 164.385 63.830 165.520 ;
        RECT 64.000 164.585 64.260 165.695 ;
        RECT 64.430 164.795 64.690 165.520 ;
        RECT 64.860 164.965 65.120 165.695 ;
        RECT 65.290 164.795 65.550 165.520 ;
        RECT 65.720 164.965 65.980 165.695 ;
        RECT 66.150 164.795 66.410 165.520 ;
        RECT 66.580 164.965 66.840 165.695 ;
        RECT 67.010 164.795 67.270 165.520 ;
        RECT 67.440 164.965 67.735 165.695 ;
        RECT 68.155 165.185 68.415 165.695 ;
        RECT 64.430 164.555 67.740 164.795 ;
        RECT 61.260 163.795 62.910 163.965 ;
        RECT 60.335 163.315 60.635 163.645 ;
        RECT 60.805 163.145 61.080 163.625 ;
        RECT 61.260 163.405 61.555 163.795 ;
        RECT 61.725 163.145 61.980 163.625 ;
        RECT 62.155 163.405 62.415 163.795 ;
        RECT 63.095 163.775 63.410 164.385 ;
        RECT 63.580 164.135 66.600 164.385 ;
        RECT 62.585 163.145 62.865 163.625 ;
        RECT 63.155 163.145 63.400 163.605 ;
        RECT 63.580 163.325 63.830 164.135 ;
        RECT 66.770 163.965 67.740 164.555 ;
        RECT 68.155 164.135 68.495 165.015 ;
        RECT 68.665 164.305 68.835 165.525 ;
        RECT 69.075 165.190 69.690 165.695 ;
        RECT 69.075 164.655 69.325 165.020 ;
        RECT 69.495 165.015 69.690 165.190 ;
        RECT 69.860 165.185 70.335 165.525 ;
        RECT 70.505 165.150 70.720 165.695 ;
        RECT 69.495 164.825 69.825 165.015 ;
        RECT 70.045 164.655 70.760 164.950 ;
        RECT 70.930 164.825 71.205 165.525 ;
        RECT 71.465 165.075 71.635 165.505 ;
        RECT 71.805 165.245 72.135 165.695 ;
        RECT 71.465 164.845 72.140 165.075 ;
        RECT 69.075 164.485 70.865 164.655 ;
        RECT 68.665 164.055 69.460 164.305 ;
        RECT 68.665 163.965 68.915 164.055 ;
        RECT 64.430 163.795 67.740 163.965 ;
        RECT 64.000 163.145 64.260 163.670 ;
        RECT 64.430 163.340 64.690 163.795 ;
        RECT 64.860 163.145 65.120 163.625 ;
        RECT 65.290 163.340 65.550 163.795 ;
        RECT 65.720 163.145 65.980 163.625 ;
        RECT 66.150 163.340 66.410 163.795 ;
        RECT 66.580 163.145 66.840 163.625 ;
        RECT 67.010 163.340 67.270 163.795 ;
        RECT 67.440 163.145 67.740 163.625 ;
        RECT 68.155 163.145 68.415 163.965 ;
        RECT 68.585 163.545 68.915 163.965 ;
        RECT 69.630 163.630 69.885 164.485 ;
        RECT 69.095 163.365 69.885 163.630 ;
        RECT 70.055 163.785 70.465 164.305 ;
        RECT 70.635 164.055 70.865 164.485 ;
        RECT 71.035 163.795 71.205 164.825 ;
        RECT 71.435 163.825 71.735 164.675 ;
        RECT 71.905 164.195 72.140 164.845 ;
        RECT 72.310 164.535 72.595 165.480 ;
        RECT 72.775 165.225 73.460 165.695 ;
        RECT 72.770 164.705 73.465 165.015 ;
        RECT 73.640 164.640 73.945 165.425 ;
        RECT 74.250 165.065 74.535 165.525 ;
        RECT 74.705 165.235 74.975 165.695 ;
        RECT 74.250 164.845 75.205 165.065 ;
        RECT 72.310 164.385 73.170 164.535 ;
        RECT 72.310 164.365 73.595 164.385 ;
        RECT 71.905 163.865 72.440 164.195 ;
        RECT 72.610 164.005 73.595 164.365 ;
        RECT 70.055 163.365 70.255 163.785 ;
        RECT 70.445 163.145 70.775 163.605 ;
        RECT 70.945 163.315 71.205 163.795 ;
        RECT 71.905 163.715 72.125 163.865 ;
        RECT 71.380 163.145 71.715 163.650 ;
        RECT 71.885 163.340 72.125 163.715 ;
        RECT 72.610 163.670 72.780 164.005 ;
        RECT 73.770 163.835 73.945 164.640 ;
        RECT 74.135 164.115 74.825 164.675 ;
        RECT 74.995 163.945 75.205 164.845 ;
        RECT 72.405 163.475 72.780 163.670 ;
        RECT 72.405 163.330 72.575 163.475 ;
        RECT 73.140 163.145 73.535 163.640 ;
        RECT 73.705 163.315 73.945 163.835 ;
        RECT 74.250 163.775 75.205 163.945 ;
        RECT 75.375 164.675 75.775 165.525 ;
        RECT 75.965 165.065 76.245 165.525 ;
        RECT 76.765 165.235 77.090 165.695 ;
        RECT 75.965 164.845 77.090 165.065 ;
        RECT 75.375 164.115 76.470 164.675 ;
        RECT 76.640 164.385 77.090 164.845 ;
        RECT 77.260 164.555 77.645 165.525 ;
        RECT 74.250 163.315 74.535 163.775 ;
        RECT 74.705 163.145 74.975 163.605 ;
        RECT 75.375 163.315 75.775 164.115 ;
        RECT 76.640 164.055 77.195 164.385 ;
        RECT 76.640 163.945 77.090 164.055 ;
        RECT 75.965 163.775 77.090 163.945 ;
        RECT 77.365 163.885 77.645 164.555 ;
        RECT 77.815 164.530 78.105 165.695 ;
        RECT 78.335 164.635 78.665 165.480 ;
        RECT 78.835 164.685 79.005 165.695 ;
        RECT 79.175 164.965 79.515 165.525 ;
        RECT 79.745 165.195 80.060 165.695 ;
        RECT 80.240 165.225 81.125 165.395 ;
        RECT 78.275 164.555 78.665 164.635 ;
        RECT 79.175 164.590 80.070 164.965 ;
        RECT 75.965 163.315 76.245 163.775 ;
        RECT 76.765 163.145 77.090 163.605 ;
        RECT 77.260 163.315 77.645 163.885 ;
        RECT 78.275 164.505 78.490 164.555 ;
        RECT 78.275 163.925 78.445 164.505 ;
        RECT 79.175 164.385 79.365 164.590 ;
        RECT 80.240 164.385 80.410 165.225 ;
        RECT 81.350 165.195 81.600 165.525 ;
        RECT 78.615 164.055 79.365 164.385 ;
        RECT 79.535 164.055 80.410 164.385 ;
        RECT 78.275 163.885 78.500 163.925 ;
        RECT 79.165 163.885 79.365 164.055 ;
        RECT 77.815 163.145 78.105 163.870 ;
        RECT 78.275 163.800 78.655 163.885 ;
        RECT 78.325 163.365 78.655 163.800 ;
        RECT 78.825 163.145 78.995 163.755 ;
        RECT 79.165 163.360 79.495 163.885 ;
        RECT 79.755 163.145 79.965 163.675 ;
        RECT 80.240 163.595 80.410 164.055 ;
        RECT 80.580 164.095 80.900 165.055 ;
        RECT 81.070 164.305 81.260 165.025 ;
        RECT 81.430 164.125 81.600 165.195 ;
        RECT 81.770 164.895 81.940 165.695 ;
        RECT 82.110 165.250 83.215 165.420 ;
        RECT 82.110 164.635 82.280 165.250 ;
        RECT 83.425 165.100 83.675 165.525 ;
        RECT 83.845 165.235 84.110 165.695 ;
        RECT 82.450 164.715 82.980 165.080 ;
        RECT 83.425 164.970 83.730 165.100 ;
        RECT 81.770 164.545 82.280 164.635 ;
        RECT 81.770 164.375 82.640 164.545 ;
        RECT 81.770 164.305 81.940 164.375 ;
        RECT 82.060 164.125 82.260 164.155 ;
        RECT 80.580 163.765 81.045 164.095 ;
        RECT 81.430 163.825 82.260 164.125 ;
        RECT 81.430 163.595 81.600 163.825 ;
        RECT 80.240 163.425 81.025 163.595 ;
        RECT 81.195 163.425 81.600 163.595 ;
        RECT 81.780 163.145 82.150 163.645 ;
        RECT 82.470 163.595 82.640 164.375 ;
        RECT 82.810 164.015 82.980 164.715 ;
        RECT 83.150 164.185 83.390 164.780 ;
        RECT 82.810 163.795 83.335 164.015 ;
        RECT 83.560 163.865 83.730 164.970 ;
        RECT 83.505 163.735 83.730 163.865 ;
        RECT 83.900 163.775 84.180 164.725 ;
        RECT 83.505 163.595 83.675 163.735 ;
        RECT 82.470 163.425 83.145 163.595 ;
        RECT 83.340 163.425 83.675 163.595 ;
        RECT 83.845 163.145 84.095 163.605 ;
        RECT 84.350 163.405 84.535 165.525 ;
        RECT 84.705 165.195 85.035 165.695 ;
        RECT 85.205 165.025 85.375 165.525 ;
        RECT 84.710 164.855 85.375 165.025 ;
        RECT 84.710 163.865 84.940 164.855 ;
        RECT 85.110 164.035 85.460 164.685 ;
        RECT 85.640 164.555 85.975 165.525 ;
        RECT 86.145 164.555 86.315 165.695 ;
        RECT 86.485 165.355 88.515 165.525 ;
        RECT 85.640 163.885 85.810 164.555 ;
        RECT 86.485 164.385 86.655 165.355 ;
        RECT 85.980 164.055 86.235 164.385 ;
        RECT 86.460 164.055 86.655 164.385 ;
        RECT 86.825 165.015 87.950 165.185 ;
        RECT 86.065 163.885 86.235 164.055 ;
        RECT 86.825 163.885 86.995 165.015 ;
        RECT 84.710 163.695 85.375 163.865 ;
        RECT 84.705 163.145 85.035 163.525 ;
        RECT 85.205 163.405 85.375 163.695 ;
        RECT 85.640 163.315 85.895 163.885 ;
        RECT 86.065 163.715 86.995 163.885 ;
        RECT 87.165 164.675 88.175 164.845 ;
        RECT 87.165 163.875 87.335 164.675 ;
        RECT 86.820 163.680 86.995 163.715 ;
        RECT 86.065 163.145 86.395 163.545 ;
        RECT 86.820 163.315 87.350 163.680 ;
        RECT 87.540 163.655 87.815 164.475 ;
        RECT 87.535 163.485 87.815 163.655 ;
        RECT 87.540 163.315 87.815 163.485 ;
        RECT 87.985 163.315 88.175 164.675 ;
        RECT 88.345 164.690 88.515 165.355 ;
        RECT 88.685 164.935 88.855 165.695 ;
        RECT 89.090 164.935 89.605 165.345 ;
        RECT 88.345 164.500 89.095 164.690 ;
        RECT 89.265 164.125 89.605 164.935 ;
        RECT 89.775 164.605 91.445 165.695 ;
        RECT 88.375 163.955 89.605 164.125 ;
        RECT 88.355 163.145 88.865 163.680 ;
        RECT 89.085 163.350 89.330 163.955 ;
        RECT 89.775 163.915 90.525 164.435 ;
        RECT 90.695 164.085 91.445 164.605 ;
        RECT 92.085 164.585 92.380 165.695 ;
        RECT 92.560 164.385 92.810 165.520 ;
        RECT 92.980 164.585 93.240 165.695 ;
        RECT 93.410 164.795 93.670 165.520 ;
        RECT 93.840 164.965 94.100 165.695 ;
        RECT 94.270 164.795 94.530 165.520 ;
        RECT 94.700 164.965 94.960 165.695 ;
        RECT 95.130 164.795 95.390 165.520 ;
        RECT 95.560 164.965 95.820 165.695 ;
        RECT 95.990 164.795 96.250 165.520 ;
        RECT 96.420 164.965 96.715 165.695 ;
        RECT 93.410 164.555 96.720 164.795 ;
        RECT 89.775 163.145 91.445 163.915 ;
        RECT 92.075 163.775 92.390 164.385 ;
        RECT 92.560 164.135 95.580 164.385 ;
        RECT 92.135 163.145 92.380 163.605 ;
        RECT 92.560 163.325 92.810 164.135 ;
        RECT 95.750 163.965 96.720 164.555 ;
        RECT 93.410 163.795 96.720 163.965 ;
        RECT 97.140 164.555 97.475 165.525 ;
        RECT 97.645 164.555 97.815 165.695 ;
        RECT 97.985 165.355 100.015 165.525 ;
        RECT 97.140 163.885 97.310 164.555 ;
        RECT 97.985 164.385 98.155 165.355 ;
        RECT 97.480 164.055 97.735 164.385 ;
        RECT 97.960 164.055 98.155 164.385 ;
        RECT 98.325 165.015 99.450 165.185 ;
        RECT 97.565 163.885 97.735 164.055 ;
        RECT 98.325 163.885 98.495 165.015 ;
        RECT 92.980 163.145 93.240 163.670 ;
        RECT 93.410 163.340 93.670 163.795 ;
        RECT 93.840 163.145 94.100 163.625 ;
        RECT 94.270 163.340 94.530 163.795 ;
        RECT 94.700 163.145 94.960 163.625 ;
        RECT 95.130 163.340 95.390 163.795 ;
        RECT 95.560 163.145 95.820 163.625 ;
        RECT 95.990 163.340 96.250 163.795 ;
        RECT 96.420 163.145 96.720 163.625 ;
        RECT 97.140 163.315 97.395 163.885 ;
        RECT 97.565 163.715 98.495 163.885 ;
        RECT 98.665 164.675 99.675 164.845 ;
        RECT 98.665 163.875 98.835 164.675 ;
        RECT 98.320 163.680 98.495 163.715 ;
        RECT 97.565 163.145 97.895 163.545 ;
        RECT 98.320 163.315 98.850 163.680 ;
        RECT 99.040 163.655 99.315 164.475 ;
        RECT 99.035 163.485 99.315 163.655 ;
        RECT 99.040 163.315 99.315 163.485 ;
        RECT 99.485 163.315 99.675 164.675 ;
        RECT 99.845 164.690 100.015 165.355 ;
        RECT 100.185 164.935 100.355 165.695 ;
        RECT 100.590 164.935 101.105 165.345 ;
        RECT 99.845 164.500 100.595 164.690 ;
        RECT 100.765 164.125 101.105 164.935 ;
        RECT 101.275 164.605 102.945 165.695 ;
        RECT 99.875 163.955 101.105 164.125 ;
        RECT 99.855 163.145 100.365 163.680 ;
        RECT 100.585 163.350 100.830 163.955 ;
        RECT 101.275 163.915 102.025 164.435 ;
        RECT 102.195 164.085 102.945 164.605 ;
        RECT 103.575 164.530 103.865 165.695 ;
        RECT 104.040 164.555 104.360 165.695 ;
        RECT 104.540 164.385 104.735 165.435 ;
        RECT 104.915 164.845 105.245 165.525 ;
        RECT 105.445 164.895 105.700 165.695 ;
        RECT 104.915 164.565 105.265 164.845 ;
        RECT 104.100 164.335 104.360 164.385 ;
        RECT 104.095 164.165 104.360 164.335 ;
        RECT 104.100 164.055 104.360 164.165 ;
        RECT 104.540 164.055 104.925 164.385 ;
        RECT 105.095 164.185 105.265 164.565 ;
        RECT 105.455 164.355 105.700 164.715 ;
        RECT 106.375 164.555 106.605 165.695 ;
        RECT 106.775 164.545 107.105 165.525 ;
        RECT 107.275 164.555 107.485 165.695 ;
        RECT 107.715 164.605 111.225 165.695 ;
        RECT 105.095 164.015 105.615 164.185 ;
        RECT 106.355 164.135 106.685 164.385 ;
        RECT 101.275 163.145 102.945 163.915 ;
        RECT 103.575 163.145 103.865 163.870 ;
        RECT 104.040 163.675 105.255 163.845 ;
        RECT 104.040 163.325 104.330 163.675 ;
        RECT 104.525 163.145 104.855 163.505 ;
        RECT 105.025 163.370 105.255 163.675 ;
        RECT 105.445 163.655 105.615 164.015 ;
        RECT 105.445 163.485 105.645 163.655 ;
        RECT 105.445 163.450 105.615 163.485 ;
        RECT 106.375 163.145 106.605 163.965 ;
        RECT 106.855 163.945 107.105 164.545 ;
        RECT 106.775 163.315 107.105 163.945 ;
        RECT 107.275 163.145 107.485 163.965 ;
        RECT 107.715 163.915 109.365 164.435 ;
        RECT 109.535 164.085 111.225 164.605 ;
        RECT 112.010 164.685 112.310 165.525 ;
        RECT 112.505 164.855 112.755 165.695 ;
        RECT 113.345 165.105 114.150 165.525 ;
        RECT 112.925 164.935 114.490 165.105 ;
        RECT 112.925 164.685 113.095 164.935 ;
        RECT 112.010 164.515 113.095 164.685 ;
        RECT 111.855 164.055 112.185 164.345 ;
        RECT 107.715 163.145 111.225 163.915 ;
        RECT 112.355 163.885 112.525 164.515 ;
        RECT 113.265 164.385 113.585 164.765 ;
        RECT 113.775 164.675 114.150 164.765 ;
        RECT 113.755 164.505 114.150 164.675 ;
        RECT 114.320 164.685 114.490 164.935 ;
        RECT 114.660 164.855 114.990 165.695 ;
        RECT 115.160 164.935 115.825 165.525 ;
        RECT 114.320 164.515 115.240 164.685 ;
        RECT 112.695 164.135 113.025 164.345 ;
        RECT 113.205 164.135 113.585 164.385 ;
        RECT 113.775 164.345 114.150 164.505 ;
        RECT 115.070 164.345 115.240 164.515 ;
        RECT 113.775 164.135 114.260 164.345 ;
        RECT 114.450 164.135 114.900 164.345 ;
        RECT 115.070 164.135 115.405 164.345 ;
        RECT 115.575 163.965 115.825 164.935 ;
        RECT 116.000 164.555 116.255 165.695 ;
        RECT 116.425 164.725 116.755 165.525 ;
        RECT 116.925 164.895 117.155 165.695 ;
        RECT 117.325 164.725 117.655 165.525 ;
        RECT 116.425 164.555 117.655 164.725 ;
        RECT 118.305 164.675 118.635 165.525 ;
        RECT 118.805 164.845 118.975 165.695 ;
        RECT 119.145 164.675 119.475 165.525 ;
        RECT 119.645 164.845 119.815 165.695 ;
        RECT 119.985 164.675 120.315 165.525 ;
        RECT 120.485 164.895 120.655 165.695 ;
        RECT 120.825 164.675 121.155 165.525 ;
        RECT 121.325 164.895 121.495 165.695 ;
        RECT 121.665 164.675 121.995 165.525 ;
        RECT 122.165 164.895 122.335 165.695 ;
        RECT 122.505 164.675 122.835 165.525 ;
        RECT 123.005 164.895 123.175 165.695 ;
        RECT 123.345 164.675 123.675 165.525 ;
        RECT 123.845 164.895 124.015 165.695 ;
        RECT 124.185 164.675 124.515 165.525 ;
        RECT 124.685 164.895 124.855 165.695 ;
        RECT 125.025 164.675 125.355 165.525 ;
        RECT 125.525 164.895 125.695 165.695 ;
        RECT 125.865 164.675 126.195 165.525 ;
        RECT 126.365 164.895 126.535 165.695 ;
        RECT 126.705 164.675 127.035 165.525 ;
        RECT 127.205 164.895 127.375 165.695 ;
        RECT 127.545 164.675 127.875 165.525 ;
        RECT 128.045 164.895 128.215 165.695 ;
        RECT 128.385 164.675 128.715 165.525 ;
        RECT 128.885 164.895 129.055 165.695 ;
        RECT 112.015 163.705 112.525 163.885 ;
        RECT 112.930 163.795 114.630 163.965 ;
        RECT 112.930 163.705 113.315 163.795 ;
        RECT 112.015 163.315 112.345 163.705 ;
        RECT 112.515 163.365 113.700 163.535 ;
        RECT 113.960 163.145 114.130 163.615 ;
        RECT 114.300 163.330 114.630 163.795 ;
        RECT 114.800 163.145 114.970 163.965 ;
        RECT 115.140 163.325 115.825 163.965 ;
        RECT 116.020 163.805 116.240 164.385 ;
        RECT 116.425 163.655 116.605 164.555 ;
        RECT 118.305 164.505 119.815 164.675 ;
        RECT 119.985 164.505 122.335 164.675 ;
        RECT 122.505 164.505 129.165 164.675 ;
        RECT 129.335 164.530 129.625 165.695 ;
        RECT 129.800 164.555 130.135 165.525 ;
        RECT 130.305 164.555 130.475 165.695 ;
        RECT 130.645 165.355 132.675 165.525 ;
        RECT 116.775 163.825 117.150 164.385 ;
        RECT 117.355 164.055 117.665 164.385 ;
        RECT 119.645 164.335 119.815 164.505 ;
        RECT 122.160 164.335 122.335 164.505 ;
        RECT 118.300 164.135 119.475 164.335 ;
        RECT 119.645 164.135 121.955 164.335 ;
        RECT 122.160 164.135 128.720 164.335 ;
        RECT 119.645 163.965 119.815 164.135 ;
        RECT 122.160 163.965 122.335 164.135 ;
        RECT 128.890 163.965 129.165 164.505 ;
        RECT 117.325 163.655 117.655 163.885 ;
        RECT 116.000 163.145 116.255 163.635 ;
        RECT 116.425 163.315 117.655 163.655 ;
        RECT 118.305 163.795 119.815 163.965 ;
        RECT 119.985 163.795 122.335 163.965 ;
        RECT 122.505 163.795 129.165 163.965 ;
        RECT 129.800 163.885 129.970 164.555 ;
        RECT 130.645 164.385 130.815 165.355 ;
        RECT 130.140 164.055 130.395 164.385 ;
        RECT 130.620 164.055 130.815 164.385 ;
        RECT 130.985 165.015 132.110 165.185 ;
        RECT 130.225 163.885 130.395 164.055 ;
        RECT 130.985 163.885 131.155 165.015 ;
        RECT 118.305 163.320 118.635 163.795 ;
        RECT 118.805 163.145 118.975 163.625 ;
        RECT 119.145 163.320 119.475 163.795 ;
        RECT 119.645 163.145 119.815 163.625 ;
        RECT 119.985 163.320 120.315 163.795 ;
        RECT 120.485 163.145 120.655 163.625 ;
        RECT 120.825 163.320 121.155 163.795 ;
        RECT 121.325 163.145 121.495 163.625 ;
        RECT 121.665 163.320 121.995 163.795 ;
        RECT 122.165 163.145 122.335 163.625 ;
        RECT 122.505 163.320 122.835 163.795 ;
        RECT 122.505 163.315 122.755 163.320 ;
        RECT 123.005 163.145 123.175 163.625 ;
        RECT 123.345 163.320 123.675 163.795 ;
        RECT 123.425 163.315 123.595 163.320 ;
        RECT 123.845 163.145 124.015 163.625 ;
        RECT 124.185 163.320 124.515 163.795 ;
        RECT 124.265 163.315 124.435 163.320 ;
        RECT 124.685 163.145 124.855 163.625 ;
        RECT 125.025 163.320 125.355 163.795 ;
        RECT 125.525 163.145 125.695 163.625 ;
        RECT 125.865 163.320 126.195 163.795 ;
        RECT 126.365 163.145 126.535 163.625 ;
        RECT 126.705 163.320 127.035 163.795 ;
        RECT 127.205 163.145 127.375 163.625 ;
        RECT 127.545 163.320 127.875 163.795 ;
        RECT 128.045 163.145 128.215 163.625 ;
        RECT 128.385 163.320 128.715 163.795 ;
        RECT 128.885 163.145 129.055 163.625 ;
        RECT 129.335 163.145 129.625 163.870 ;
        RECT 129.800 163.315 130.055 163.885 ;
        RECT 130.225 163.715 131.155 163.885 ;
        RECT 131.325 164.675 132.335 164.845 ;
        RECT 131.325 163.875 131.495 164.675 ;
        RECT 131.700 163.995 131.975 164.475 ;
        RECT 131.695 163.825 131.975 163.995 ;
        RECT 130.980 163.680 131.155 163.715 ;
        RECT 130.225 163.145 130.555 163.545 ;
        RECT 130.980 163.315 131.510 163.680 ;
        RECT 131.700 163.315 131.975 163.825 ;
        RECT 132.145 163.315 132.335 164.675 ;
        RECT 132.505 164.690 132.675 165.355 ;
        RECT 132.845 164.935 133.015 165.695 ;
        RECT 133.250 164.935 133.765 165.345 ;
        RECT 132.505 164.500 133.255 164.690 ;
        RECT 133.425 164.125 133.765 164.935 ;
        RECT 132.535 163.955 133.765 164.125 ;
        RECT 133.935 164.555 134.320 165.525 ;
        RECT 134.490 165.235 134.815 165.695 ;
        RECT 135.335 165.065 135.615 165.525 ;
        RECT 134.490 164.845 135.615 165.065 ;
        RECT 132.515 163.145 133.025 163.680 ;
        RECT 133.245 163.350 133.490 163.955 ;
        RECT 133.935 163.885 134.215 164.555 ;
        RECT 134.490 164.385 134.940 164.845 ;
        RECT 135.805 164.675 136.205 165.525 ;
        RECT 136.605 165.235 136.875 165.695 ;
        RECT 137.045 165.065 137.330 165.525 ;
        RECT 134.385 164.055 134.940 164.385 ;
        RECT 135.110 164.115 136.205 164.675 ;
        RECT 134.490 163.945 134.940 164.055 ;
        RECT 133.935 163.315 134.320 163.885 ;
        RECT 134.490 163.775 135.615 163.945 ;
        RECT 134.490 163.145 134.815 163.605 ;
        RECT 135.335 163.315 135.615 163.775 ;
        RECT 135.805 163.315 136.205 164.115 ;
        RECT 136.375 164.845 137.330 165.065 ;
        RECT 136.375 163.945 136.585 164.845 ;
        RECT 136.755 164.115 137.445 164.675 ;
        RECT 137.615 164.605 138.825 165.695 ;
        RECT 137.615 164.065 138.135 164.605 ;
        RECT 136.375 163.775 137.330 163.945 ;
        RECT 138.305 163.895 138.825 164.435 ;
        RECT 136.605 163.145 136.875 163.605 ;
        RECT 137.045 163.315 137.330 163.775 ;
        RECT 137.615 163.145 138.825 163.895 ;
        RECT 13.330 162.975 138.910 163.145 ;
        RECT 13.415 162.225 14.625 162.975 ;
        RECT 14.795 162.430 20.140 162.975 ;
        RECT 13.415 161.685 13.935 162.225 ;
        RECT 14.105 161.515 14.625 162.055 ;
        RECT 16.380 161.600 16.720 162.430 ;
        RECT 20.315 162.205 21.985 162.975 ;
        RECT 22.665 162.585 22.995 162.975 ;
        RECT 23.165 162.405 23.335 162.725 ;
        RECT 23.505 162.585 23.835 162.975 ;
        RECT 24.250 162.575 25.205 162.745 ;
        RECT 22.615 162.235 24.865 162.405 ;
        RECT 13.415 160.425 14.625 161.515 ;
        RECT 18.200 160.860 18.550 162.110 ;
        RECT 20.315 161.685 21.065 162.205 ;
        RECT 21.235 161.515 21.985 162.035 ;
        RECT 14.795 160.425 20.140 160.860 ;
        RECT 20.315 160.425 21.985 161.515 ;
        RECT 22.615 161.275 22.785 162.235 ;
        RECT 22.955 161.615 23.200 162.065 ;
        RECT 23.370 161.785 23.920 161.985 ;
        RECT 24.090 161.815 24.465 161.985 ;
        RECT 24.090 161.615 24.260 161.815 ;
        RECT 24.635 161.735 24.865 162.235 ;
        RECT 22.955 161.445 24.260 161.615 ;
        RECT 25.035 161.695 25.205 162.575 ;
        RECT 25.375 162.140 25.665 162.975 ;
        RECT 25.835 162.205 28.425 162.975 ;
        RECT 29.060 162.325 29.330 162.535 ;
        RECT 29.550 162.515 29.880 162.975 ;
        RECT 30.390 162.515 31.140 162.805 ;
        RECT 25.035 161.525 25.665 161.695 ;
        RECT 25.835 161.685 27.045 162.205 ;
        RECT 29.060 162.155 30.395 162.325 ;
        RECT 22.615 160.595 22.995 161.275 ;
        RECT 23.585 160.425 23.755 161.275 ;
        RECT 23.925 161.105 25.165 161.275 ;
        RECT 23.925 160.595 24.255 161.105 ;
        RECT 24.425 160.425 24.595 160.935 ;
        RECT 24.765 160.595 25.165 161.105 ;
        RECT 25.345 160.595 25.665 161.525 ;
        RECT 27.215 161.515 28.425 162.035 ;
        RECT 30.225 161.985 30.395 162.155 ;
        RECT 29.060 161.745 29.410 161.985 ;
        RECT 29.580 161.745 30.055 161.985 ;
        RECT 30.225 161.735 30.600 161.985 ;
        RECT 30.225 161.565 30.395 161.735 ;
        RECT 25.835 160.425 28.425 161.515 ;
        RECT 29.060 161.395 30.395 161.565 ;
        RECT 29.060 161.235 29.340 161.395 ;
        RECT 30.770 161.225 31.140 162.515 ;
        RECT 31.355 162.430 36.700 162.975 ;
        RECT 32.940 161.600 33.280 162.430 ;
        RECT 36.875 162.205 38.545 162.975 ;
        RECT 39.175 162.250 39.465 162.975 ;
        RECT 29.550 160.425 29.800 161.225 ;
        RECT 29.970 161.055 31.140 161.225 ;
        RECT 29.970 160.595 30.300 161.055 ;
        RECT 30.470 160.425 30.685 160.885 ;
        RECT 34.760 160.860 35.110 162.110 ;
        RECT 36.875 161.685 37.625 162.205 ;
        RECT 39.675 162.155 39.905 162.975 ;
        RECT 40.075 162.175 40.405 162.805 ;
        RECT 37.795 161.515 38.545 162.035 ;
        RECT 39.655 161.735 39.985 161.985 ;
        RECT 31.355 160.425 36.700 160.860 ;
        RECT 36.875 160.425 38.545 161.515 ;
        RECT 39.175 160.425 39.465 161.590 ;
        RECT 40.155 161.575 40.405 162.175 ;
        RECT 40.575 162.155 40.785 162.975 ;
        RECT 41.475 162.235 41.940 162.780 ;
        RECT 39.675 160.425 39.905 161.565 ;
        RECT 40.075 160.595 40.405 161.575 ;
        RECT 40.575 160.425 40.785 161.565 ;
        RECT 41.475 161.275 41.645 162.235 ;
        RECT 42.445 162.155 42.615 162.975 ;
        RECT 42.785 162.325 43.115 162.805 ;
        RECT 43.285 162.585 43.635 162.975 ;
        RECT 43.805 162.405 44.035 162.805 ;
        RECT 43.525 162.325 44.035 162.405 ;
        RECT 42.785 162.235 44.035 162.325 ;
        RECT 44.205 162.235 44.525 162.715 ;
        RECT 44.705 162.475 45.035 162.975 ;
        RECT 45.235 162.405 45.405 162.755 ;
        RECT 45.605 162.575 45.935 162.975 ;
        RECT 46.105 162.405 46.275 162.755 ;
        RECT 46.445 162.575 46.825 162.975 ;
        RECT 42.785 162.155 43.695 162.235 ;
        RECT 41.815 161.615 42.060 162.065 ;
        RECT 42.320 161.785 43.015 161.985 ;
        RECT 43.185 161.815 43.785 161.985 ;
        RECT 43.185 161.615 43.355 161.815 ;
        RECT 44.015 161.645 44.185 162.065 ;
        RECT 41.815 161.445 43.355 161.615 ;
        RECT 43.525 161.475 44.185 161.645 ;
        RECT 43.525 161.275 43.695 161.475 ;
        RECT 44.355 161.305 44.525 162.235 ;
        RECT 44.700 161.735 45.050 162.305 ;
        RECT 45.235 162.235 46.845 162.405 ;
        RECT 47.015 162.300 47.285 162.645 ;
        RECT 46.675 162.065 46.845 162.235 ;
        RECT 41.475 161.105 43.695 161.275 ;
        RECT 43.865 161.105 44.525 161.305 ;
        RECT 44.700 161.275 45.020 161.565 ;
        RECT 45.220 161.445 45.930 162.065 ;
        RECT 46.100 161.735 46.505 162.065 ;
        RECT 46.675 161.735 46.945 162.065 ;
        RECT 46.675 161.565 46.845 161.735 ;
        RECT 47.115 161.565 47.285 162.300 ;
        RECT 47.455 162.205 49.125 162.975 ;
        RECT 49.295 162.235 49.615 162.715 ;
        RECT 49.785 162.405 50.015 162.805 ;
        RECT 50.185 162.585 50.535 162.975 ;
        RECT 49.785 162.325 50.295 162.405 ;
        RECT 50.705 162.325 51.035 162.805 ;
        RECT 49.785 162.235 51.035 162.325 ;
        RECT 47.455 161.685 48.205 162.205 ;
        RECT 46.120 161.395 46.845 161.565 ;
        RECT 46.120 161.275 46.290 161.395 ;
        RECT 44.700 161.105 46.290 161.275 ;
        RECT 41.475 160.425 41.775 160.935 ;
        RECT 41.945 160.595 42.275 161.105 ;
        RECT 43.865 160.935 44.035 161.105 ;
        RECT 42.445 160.425 43.075 160.935 ;
        RECT 43.655 160.765 44.035 160.935 ;
        RECT 44.205 160.425 44.505 160.935 ;
        RECT 44.700 160.645 46.355 160.935 ;
        RECT 46.525 160.425 46.805 161.225 ;
        RECT 47.015 160.595 47.285 161.565 ;
        RECT 48.375 161.515 49.125 162.035 ;
        RECT 47.455 160.425 49.125 161.515 ;
        RECT 49.295 161.305 49.465 162.235 ;
        RECT 50.125 162.155 51.035 162.235 ;
        RECT 51.205 162.155 51.375 162.975 ;
        RECT 51.880 162.235 52.345 162.780 ;
        RECT 52.515 162.430 57.860 162.975 ;
        RECT 58.035 162.430 63.380 162.975 ;
        RECT 49.635 161.645 49.805 162.065 ;
        RECT 50.035 161.815 50.635 161.985 ;
        RECT 49.635 161.475 50.295 161.645 ;
        RECT 49.295 161.105 49.955 161.305 ;
        RECT 50.125 161.275 50.295 161.475 ;
        RECT 50.465 161.615 50.635 161.815 ;
        RECT 50.805 161.785 51.500 161.985 ;
        RECT 51.760 161.615 52.005 162.065 ;
        RECT 50.465 161.445 52.005 161.615 ;
        RECT 52.175 161.275 52.345 162.235 ;
        RECT 54.100 161.600 54.440 162.430 ;
        RECT 50.125 161.105 52.345 161.275 ;
        RECT 49.785 160.935 49.955 161.105 ;
        RECT 49.315 160.425 49.615 160.935 ;
        RECT 49.785 160.765 50.165 160.935 ;
        RECT 50.745 160.425 51.375 160.935 ;
        RECT 51.545 160.595 51.875 161.105 ;
        RECT 52.045 160.425 52.345 160.935 ;
        RECT 55.920 160.860 56.270 162.110 ;
        RECT 59.620 161.600 59.960 162.430 ;
        RECT 63.555 162.225 64.765 162.975 ;
        RECT 64.935 162.250 65.225 162.975 ;
        RECT 65.485 162.425 65.655 162.715 ;
        RECT 65.825 162.595 66.155 162.975 ;
        RECT 65.485 162.255 66.150 162.425 ;
        RECT 61.440 160.860 61.790 162.110 ;
        RECT 63.555 161.685 64.075 162.225 ;
        RECT 64.245 161.515 64.765 162.055 ;
        RECT 52.515 160.425 57.860 160.860 ;
        RECT 58.035 160.425 63.380 160.860 ;
        RECT 63.555 160.425 64.765 161.515 ;
        RECT 64.935 160.425 65.225 161.590 ;
        RECT 65.400 161.435 65.750 162.085 ;
        RECT 65.920 161.265 66.150 162.255 ;
        RECT 65.485 161.095 66.150 161.265 ;
        RECT 65.485 160.595 65.655 161.095 ;
        RECT 65.825 160.425 66.155 160.925 ;
        RECT 66.325 160.595 66.510 162.715 ;
        RECT 66.765 162.515 67.015 162.975 ;
        RECT 67.185 162.525 67.520 162.695 ;
        RECT 67.715 162.525 68.390 162.695 ;
        RECT 67.185 162.385 67.355 162.525 ;
        RECT 66.680 161.395 66.960 162.345 ;
        RECT 67.130 162.255 67.355 162.385 ;
        RECT 67.130 161.150 67.300 162.255 ;
        RECT 67.525 162.105 68.050 162.325 ;
        RECT 67.470 161.340 67.710 161.935 ;
        RECT 67.880 161.405 68.050 162.105 ;
        RECT 68.220 161.745 68.390 162.525 ;
        RECT 68.710 162.475 69.080 162.975 ;
        RECT 69.260 162.525 69.665 162.695 ;
        RECT 69.835 162.525 70.620 162.695 ;
        RECT 69.260 162.295 69.430 162.525 ;
        RECT 68.600 161.995 69.430 162.295 ;
        RECT 69.815 162.025 70.280 162.355 ;
        RECT 68.600 161.965 68.800 161.995 ;
        RECT 68.920 161.745 69.090 161.815 ;
        RECT 68.220 161.575 69.090 161.745 ;
        RECT 68.580 161.485 69.090 161.575 ;
        RECT 67.130 161.020 67.435 161.150 ;
        RECT 67.880 161.040 68.410 161.405 ;
        RECT 66.750 160.425 67.015 160.885 ;
        RECT 67.185 160.595 67.435 161.020 ;
        RECT 68.580 160.870 68.750 161.485 ;
        RECT 67.645 160.700 68.750 160.870 ;
        RECT 68.920 160.425 69.090 161.225 ;
        RECT 69.260 160.925 69.430 161.995 ;
        RECT 69.600 161.095 69.790 161.815 ;
        RECT 69.960 161.065 70.280 162.025 ;
        RECT 70.450 162.065 70.620 162.525 ;
        RECT 70.895 162.445 71.105 162.975 ;
        RECT 71.365 162.235 71.695 162.760 ;
        RECT 71.865 162.365 72.035 162.975 ;
        RECT 72.205 162.320 72.535 162.755 ;
        RECT 72.205 162.235 72.585 162.320 ;
        RECT 71.495 162.065 71.695 162.235 ;
        RECT 72.360 162.195 72.585 162.235 ;
        RECT 70.450 161.735 71.325 162.065 ;
        RECT 71.495 161.735 72.245 162.065 ;
        RECT 69.260 160.595 69.510 160.925 ;
        RECT 70.450 160.895 70.620 161.735 ;
        RECT 71.495 161.530 71.685 161.735 ;
        RECT 72.415 161.615 72.585 162.195 ;
        RECT 72.370 161.565 72.585 161.615 ;
        RECT 70.790 161.155 71.685 161.530 ;
        RECT 72.195 161.485 72.585 161.565 ;
        RECT 72.755 162.235 73.140 162.805 ;
        RECT 73.310 162.515 73.635 162.975 ;
        RECT 74.155 162.345 74.435 162.805 ;
        RECT 72.755 161.565 73.035 162.235 ;
        RECT 73.310 162.175 74.435 162.345 ;
        RECT 73.310 162.065 73.760 162.175 ;
        RECT 73.205 161.735 73.760 162.065 ;
        RECT 74.625 162.005 75.025 162.805 ;
        RECT 75.425 162.515 75.695 162.975 ;
        RECT 75.865 162.345 76.150 162.805 ;
        RECT 69.735 160.725 70.620 160.895 ;
        RECT 70.800 160.425 71.115 160.925 ;
        RECT 71.345 160.595 71.685 161.155 ;
        RECT 71.855 160.425 72.025 161.435 ;
        RECT 72.195 160.640 72.525 161.485 ;
        RECT 72.755 160.595 73.140 161.565 ;
        RECT 73.310 161.275 73.760 161.735 ;
        RECT 73.930 161.445 75.025 162.005 ;
        RECT 73.310 161.055 74.435 161.275 ;
        RECT 73.310 160.425 73.635 160.885 ;
        RECT 74.155 160.595 74.435 161.055 ;
        RECT 74.625 160.595 75.025 161.445 ;
        RECT 75.195 162.175 76.150 162.345 ;
        RECT 76.435 162.205 78.105 162.975 ;
        RECT 78.325 162.320 78.655 162.755 ;
        RECT 78.825 162.365 78.995 162.975 ;
        RECT 78.275 162.235 78.655 162.320 ;
        RECT 79.165 162.235 79.495 162.760 ;
        RECT 79.755 162.445 79.965 162.975 ;
        RECT 80.240 162.525 81.025 162.695 ;
        RECT 81.195 162.525 81.600 162.695 ;
        RECT 75.195 161.275 75.405 162.175 ;
        RECT 75.575 161.445 76.265 162.005 ;
        RECT 76.435 161.685 77.185 162.205 ;
        RECT 78.275 162.195 78.500 162.235 ;
        RECT 77.355 161.515 78.105 162.035 ;
        RECT 75.195 161.055 76.150 161.275 ;
        RECT 75.425 160.425 75.695 160.885 ;
        RECT 75.865 160.595 76.150 161.055 ;
        RECT 76.435 160.425 78.105 161.515 ;
        RECT 78.275 161.615 78.445 162.195 ;
        RECT 79.165 162.065 79.365 162.235 ;
        RECT 80.240 162.065 80.410 162.525 ;
        RECT 78.615 161.735 79.365 162.065 ;
        RECT 79.535 161.735 80.410 162.065 ;
        RECT 78.275 161.565 78.490 161.615 ;
        RECT 78.275 161.485 78.665 161.565 ;
        RECT 78.335 160.640 78.665 161.485 ;
        RECT 79.175 161.530 79.365 161.735 ;
        RECT 78.835 160.425 79.005 161.435 ;
        RECT 79.175 161.155 80.070 161.530 ;
        RECT 79.175 160.595 79.515 161.155 ;
        RECT 79.745 160.425 80.060 160.925 ;
        RECT 80.240 160.895 80.410 161.735 ;
        RECT 80.580 162.025 81.045 162.355 ;
        RECT 81.430 162.295 81.600 162.525 ;
        RECT 81.780 162.475 82.150 162.975 ;
        RECT 82.470 162.525 83.145 162.695 ;
        RECT 83.340 162.525 83.675 162.695 ;
        RECT 80.580 161.065 80.900 162.025 ;
        RECT 81.430 161.995 82.260 162.295 ;
        RECT 81.070 161.095 81.260 161.815 ;
        RECT 81.430 160.925 81.600 161.995 ;
        RECT 82.060 161.965 82.260 161.995 ;
        RECT 81.770 161.745 81.940 161.815 ;
        RECT 82.470 161.745 82.640 162.525 ;
        RECT 83.505 162.385 83.675 162.525 ;
        RECT 83.845 162.515 84.095 162.975 ;
        RECT 81.770 161.575 82.640 161.745 ;
        RECT 82.810 162.105 83.335 162.325 ;
        RECT 83.505 162.255 83.730 162.385 ;
        RECT 81.770 161.485 82.280 161.575 ;
        RECT 80.240 160.725 81.125 160.895 ;
        RECT 81.350 160.595 81.600 160.925 ;
        RECT 81.770 160.425 81.940 161.225 ;
        RECT 82.110 160.870 82.280 161.485 ;
        RECT 82.810 161.405 82.980 162.105 ;
        RECT 82.450 161.040 82.980 161.405 ;
        RECT 83.150 161.340 83.390 161.935 ;
        RECT 83.560 161.150 83.730 162.255 ;
        RECT 83.900 161.395 84.180 162.345 ;
        RECT 83.425 161.020 83.730 161.150 ;
        RECT 82.110 160.700 83.215 160.870 ;
        RECT 83.425 160.595 83.675 161.020 ;
        RECT 83.845 160.425 84.110 160.885 ;
        RECT 84.350 160.595 84.535 162.715 ;
        RECT 84.705 162.595 85.035 162.975 ;
        RECT 85.205 162.425 85.375 162.715 ;
        RECT 84.710 162.255 85.375 162.425 ;
        RECT 84.710 161.265 84.940 162.255 ;
        RECT 85.640 162.235 85.895 162.805 ;
        RECT 86.065 162.575 86.395 162.975 ;
        RECT 86.820 162.440 87.350 162.805 ;
        RECT 86.820 162.405 86.995 162.440 ;
        RECT 86.065 162.235 86.995 162.405 ;
        RECT 85.110 161.435 85.460 162.085 ;
        RECT 85.640 161.565 85.810 162.235 ;
        RECT 86.065 162.065 86.235 162.235 ;
        RECT 85.980 161.735 86.235 162.065 ;
        RECT 86.460 161.735 86.655 162.065 ;
        RECT 84.710 161.095 85.375 161.265 ;
        RECT 84.705 160.425 85.035 160.925 ;
        RECT 85.205 160.595 85.375 161.095 ;
        RECT 85.640 160.595 85.975 161.565 ;
        RECT 86.145 160.425 86.315 161.565 ;
        RECT 86.485 160.765 86.655 161.735 ;
        RECT 86.825 161.105 86.995 162.235 ;
        RECT 87.165 161.445 87.335 162.245 ;
        RECT 87.540 161.955 87.815 162.805 ;
        RECT 87.535 161.785 87.815 161.955 ;
        RECT 87.540 161.645 87.815 161.785 ;
        RECT 87.985 161.445 88.175 162.805 ;
        RECT 88.355 162.440 88.865 162.975 ;
        RECT 89.085 162.165 89.330 162.770 ;
        RECT 90.695 162.250 90.985 162.975 ;
        RECT 92.135 162.515 92.380 162.975 ;
        RECT 88.375 161.995 89.605 162.165 ;
        RECT 87.165 161.275 88.175 161.445 ;
        RECT 88.345 161.430 89.095 161.620 ;
        RECT 86.825 160.935 87.950 161.105 ;
        RECT 88.345 160.765 88.515 161.430 ;
        RECT 89.265 161.185 89.605 161.995 ;
        RECT 92.075 161.735 92.390 162.345 ;
        RECT 92.560 161.985 92.810 162.795 ;
        RECT 92.980 162.450 93.240 162.975 ;
        RECT 93.410 162.325 93.670 162.780 ;
        RECT 93.840 162.495 94.100 162.975 ;
        RECT 94.270 162.325 94.530 162.780 ;
        RECT 94.700 162.495 94.960 162.975 ;
        RECT 95.130 162.325 95.390 162.780 ;
        RECT 95.560 162.495 95.820 162.975 ;
        RECT 95.990 162.325 96.250 162.780 ;
        RECT 96.420 162.495 96.720 162.975 ;
        RECT 93.410 162.155 96.720 162.325 ;
        RECT 92.560 161.735 95.580 161.985 ;
        RECT 86.485 160.595 88.515 160.765 ;
        RECT 88.685 160.425 88.855 161.185 ;
        RECT 89.090 160.775 89.605 161.185 ;
        RECT 90.695 160.425 90.985 161.590 ;
        RECT 92.085 160.425 92.380 161.535 ;
        RECT 92.560 160.600 92.810 161.735 ;
        RECT 95.750 161.565 96.720 162.155 ;
        RECT 92.980 160.425 93.240 161.535 ;
        RECT 93.410 161.325 96.720 161.565 ;
        RECT 97.140 162.235 97.395 162.805 ;
        RECT 97.565 162.575 97.895 162.975 ;
        RECT 98.320 162.440 98.850 162.805 ;
        RECT 98.320 162.405 98.495 162.440 ;
        RECT 97.565 162.235 98.495 162.405 ;
        RECT 99.040 162.295 99.315 162.805 ;
        RECT 97.140 161.565 97.310 162.235 ;
        RECT 97.565 162.065 97.735 162.235 ;
        RECT 97.480 161.735 97.735 162.065 ;
        RECT 97.960 161.735 98.155 162.065 ;
        RECT 93.410 160.600 93.670 161.325 ;
        RECT 93.840 160.425 94.100 161.155 ;
        RECT 94.270 160.600 94.530 161.325 ;
        RECT 94.700 160.425 94.960 161.155 ;
        RECT 95.130 160.600 95.390 161.325 ;
        RECT 95.560 160.425 95.820 161.155 ;
        RECT 95.990 160.600 96.250 161.325 ;
        RECT 96.420 160.425 96.715 161.155 ;
        RECT 97.140 160.595 97.475 161.565 ;
        RECT 97.645 160.425 97.815 161.565 ;
        RECT 97.985 160.765 98.155 161.735 ;
        RECT 98.325 161.105 98.495 162.235 ;
        RECT 98.665 161.445 98.835 162.245 ;
        RECT 99.035 162.125 99.315 162.295 ;
        RECT 99.040 161.645 99.315 162.125 ;
        RECT 99.485 161.445 99.675 162.805 ;
        RECT 99.855 162.440 100.365 162.975 ;
        RECT 100.585 162.165 100.830 162.770 ;
        RECT 101.280 162.235 101.535 162.805 ;
        RECT 101.705 162.575 102.035 162.975 ;
        RECT 102.460 162.440 102.990 162.805 ;
        RECT 102.460 162.405 102.635 162.440 ;
        RECT 101.705 162.235 102.635 162.405 ;
        RECT 99.875 161.995 101.105 162.165 ;
        RECT 98.665 161.275 99.675 161.445 ;
        RECT 99.845 161.430 100.595 161.620 ;
        RECT 98.325 160.935 99.450 161.105 ;
        RECT 99.845 160.765 100.015 161.430 ;
        RECT 100.765 161.185 101.105 161.995 ;
        RECT 97.985 160.595 100.015 160.765 ;
        RECT 100.185 160.425 100.355 161.185 ;
        RECT 100.590 160.775 101.105 161.185 ;
        RECT 101.280 161.565 101.450 162.235 ;
        RECT 101.705 162.065 101.875 162.235 ;
        RECT 101.620 161.735 101.875 162.065 ;
        RECT 102.100 161.735 102.295 162.065 ;
        RECT 101.280 160.595 101.615 161.565 ;
        RECT 101.785 160.425 101.955 161.565 ;
        RECT 102.125 160.765 102.295 161.735 ;
        RECT 102.465 161.105 102.635 162.235 ;
        RECT 102.805 161.445 102.975 162.245 ;
        RECT 103.180 161.955 103.455 162.805 ;
        RECT 103.175 161.785 103.455 161.955 ;
        RECT 103.180 161.645 103.455 161.785 ;
        RECT 103.625 161.445 103.815 162.805 ;
        RECT 103.995 162.440 104.505 162.975 ;
        RECT 104.725 162.165 104.970 162.770 ;
        RECT 105.415 162.235 105.800 162.805 ;
        RECT 105.970 162.515 106.295 162.975 ;
        RECT 106.815 162.345 107.095 162.805 ;
        RECT 104.015 161.995 105.245 162.165 ;
        RECT 102.805 161.275 103.815 161.445 ;
        RECT 103.985 161.430 104.735 161.620 ;
        RECT 102.465 160.935 103.590 161.105 ;
        RECT 103.985 160.765 104.155 161.430 ;
        RECT 104.905 161.185 105.245 161.995 ;
        RECT 102.125 160.595 104.155 160.765 ;
        RECT 104.325 160.425 104.495 161.185 ;
        RECT 104.730 160.775 105.245 161.185 ;
        RECT 105.415 161.565 105.695 162.235 ;
        RECT 105.970 162.175 107.095 162.345 ;
        RECT 105.970 162.065 106.420 162.175 ;
        RECT 105.865 161.735 106.420 162.065 ;
        RECT 107.285 162.005 107.685 162.805 ;
        RECT 108.085 162.515 108.355 162.975 ;
        RECT 108.525 162.345 108.810 162.805 ;
        RECT 105.415 160.595 105.800 161.565 ;
        RECT 105.970 161.275 106.420 161.735 ;
        RECT 106.590 161.445 107.685 162.005 ;
        RECT 105.970 161.055 107.095 161.275 ;
        RECT 105.970 160.425 106.295 160.885 ;
        RECT 106.815 160.595 107.095 161.055 ;
        RECT 107.285 160.595 107.685 161.445 ;
        RECT 107.855 162.175 108.810 162.345 ;
        RECT 109.100 162.210 109.555 162.975 ;
        RECT 109.830 162.595 111.130 162.805 ;
        RECT 111.385 162.615 111.715 162.975 ;
        RECT 110.960 162.445 111.130 162.595 ;
        RECT 111.885 162.475 112.145 162.805 ;
        RECT 107.855 161.275 108.065 162.175 ;
        RECT 108.235 161.445 108.925 162.005 ;
        RECT 110.030 161.985 110.250 162.385 ;
        RECT 109.095 161.785 109.585 161.985 ;
        RECT 109.775 161.775 110.250 161.985 ;
        RECT 110.495 161.985 110.705 162.385 ;
        RECT 110.960 162.320 111.715 162.445 ;
        RECT 110.960 162.275 111.805 162.320 ;
        RECT 111.535 162.155 111.805 162.275 ;
        RECT 110.495 161.775 110.825 161.985 ;
        RECT 110.995 161.715 111.405 162.020 ;
        RECT 109.100 161.545 110.275 161.605 ;
        RECT 111.635 161.580 111.805 162.155 ;
        RECT 111.605 161.545 111.805 161.580 ;
        RECT 109.100 161.435 111.805 161.545 ;
        RECT 107.855 161.055 108.810 161.275 ;
        RECT 108.085 160.425 108.355 160.885 ;
        RECT 108.525 160.595 108.810 161.055 ;
        RECT 109.100 160.815 109.355 161.435 ;
        RECT 109.945 161.375 111.745 161.435 ;
        RECT 109.945 161.345 110.275 161.375 ;
        RECT 111.975 161.275 112.145 162.475 ;
        RECT 109.605 161.175 109.790 161.265 ;
        RECT 110.380 161.175 111.215 161.185 ;
        RECT 109.605 160.975 111.215 161.175 ;
        RECT 109.605 160.935 109.835 160.975 ;
        RECT 109.100 160.595 109.435 160.815 ;
        RECT 110.440 160.425 110.795 160.805 ;
        RECT 110.965 160.595 111.215 160.975 ;
        RECT 111.465 160.425 111.715 161.205 ;
        RECT 111.885 160.595 112.145 161.275 ;
        RECT 112.325 162.250 112.655 162.760 ;
        RECT 112.825 162.575 113.155 162.975 ;
        RECT 114.205 162.405 114.535 162.745 ;
        RECT 114.705 162.575 115.035 162.975 ;
        RECT 112.325 161.485 112.515 162.250 ;
        RECT 112.825 162.235 115.190 162.405 ;
        RECT 116.455 162.250 116.745 162.975 ;
        RECT 116.930 162.405 117.185 162.755 ;
        RECT 117.355 162.575 117.685 162.975 ;
        RECT 117.855 162.405 118.025 162.755 ;
        RECT 118.195 162.575 118.575 162.975 ;
        RECT 116.930 162.235 118.595 162.405 ;
        RECT 118.765 162.300 119.040 162.645 ;
        RECT 119.275 162.515 119.520 162.975 ;
        RECT 112.825 162.065 112.995 162.235 ;
        RECT 112.685 161.735 112.995 162.065 ;
        RECT 113.165 161.735 113.470 162.065 ;
        RECT 112.325 160.635 112.655 161.485 ;
        RECT 112.825 160.425 113.075 161.565 ;
        RECT 113.255 161.405 113.470 161.735 ;
        RECT 113.645 161.405 113.930 162.065 ;
        RECT 114.125 161.405 114.390 162.065 ;
        RECT 114.605 161.405 114.850 162.065 ;
        RECT 115.020 161.235 115.190 162.235 ;
        RECT 118.425 162.065 118.595 162.235 ;
        RECT 116.915 161.735 117.260 162.065 ;
        RECT 117.430 161.735 118.255 162.065 ;
        RECT 118.425 161.735 118.700 162.065 ;
        RECT 113.265 161.065 114.555 161.235 ;
        RECT 113.265 160.645 113.515 161.065 ;
        RECT 113.745 160.425 114.075 160.895 ;
        RECT 114.305 160.645 114.555 161.065 ;
        RECT 114.735 161.065 115.190 161.235 ;
        RECT 114.735 160.635 115.065 161.065 ;
        RECT 116.455 160.425 116.745 161.590 ;
        RECT 116.935 161.275 117.260 161.565 ;
        RECT 117.430 161.445 117.625 161.735 ;
        RECT 118.425 161.565 118.595 161.735 ;
        RECT 118.870 161.565 119.040 162.300 ;
        RECT 119.215 161.735 119.530 162.345 ;
        RECT 119.700 161.985 119.950 162.795 ;
        RECT 120.120 162.450 120.380 162.975 ;
        RECT 120.550 162.325 120.810 162.780 ;
        RECT 120.980 162.495 121.240 162.975 ;
        RECT 121.410 162.325 121.670 162.780 ;
        RECT 121.840 162.495 122.100 162.975 ;
        RECT 122.270 162.325 122.530 162.780 ;
        RECT 122.700 162.495 122.960 162.975 ;
        RECT 123.130 162.325 123.390 162.780 ;
        RECT 123.560 162.495 123.860 162.975 ;
        RECT 124.440 162.465 124.680 162.975 ;
        RECT 124.860 162.465 125.140 162.795 ;
        RECT 125.370 162.465 125.585 162.975 ;
        RECT 120.550 162.155 123.860 162.325 ;
        RECT 119.700 161.735 122.720 161.985 ;
        RECT 117.935 161.395 118.595 161.565 ;
        RECT 117.935 161.275 118.105 161.395 ;
        RECT 116.935 161.105 118.105 161.275 ;
        RECT 116.915 160.645 118.105 160.935 ;
        RECT 118.275 160.425 118.555 161.225 ;
        RECT 118.765 160.595 119.040 161.565 ;
        RECT 119.225 160.425 119.520 161.535 ;
        RECT 119.700 160.600 119.950 161.735 ;
        RECT 122.890 161.565 123.860 162.155 ;
        RECT 124.335 161.735 124.690 162.295 ;
        RECT 124.860 161.565 125.030 162.465 ;
        RECT 125.200 161.735 125.465 162.295 ;
        RECT 125.755 162.235 126.370 162.805 ;
        RECT 126.665 162.425 126.835 162.715 ;
        RECT 127.005 162.595 127.335 162.975 ;
        RECT 126.665 162.255 127.330 162.425 ;
        RECT 125.715 161.565 125.885 162.065 ;
        RECT 120.120 160.425 120.380 161.535 ;
        RECT 120.550 161.325 123.860 161.565 ;
        RECT 124.460 161.395 125.885 161.565 ;
        RECT 120.550 160.600 120.810 161.325 ;
        RECT 120.980 160.425 121.240 161.155 ;
        RECT 121.410 160.600 121.670 161.325 ;
        RECT 121.840 160.425 122.100 161.155 ;
        RECT 122.270 160.600 122.530 161.325 ;
        RECT 122.700 160.425 122.960 161.155 ;
        RECT 123.130 160.600 123.390 161.325 ;
        RECT 124.460 161.220 124.850 161.395 ;
        RECT 123.560 160.425 123.855 161.155 ;
        RECT 125.335 160.425 125.665 161.225 ;
        RECT 126.055 161.215 126.370 162.235 ;
        RECT 126.580 161.435 126.930 162.085 ;
        RECT 127.100 161.265 127.330 162.255 ;
        RECT 125.835 160.595 126.370 161.215 ;
        RECT 126.665 161.095 127.330 161.265 ;
        RECT 126.665 160.595 126.835 161.095 ;
        RECT 127.005 160.425 127.335 160.925 ;
        RECT 127.505 160.595 127.690 162.715 ;
        RECT 127.945 162.515 128.195 162.975 ;
        RECT 128.365 162.525 128.700 162.695 ;
        RECT 128.895 162.525 129.570 162.695 ;
        RECT 128.365 162.385 128.535 162.525 ;
        RECT 127.860 161.395 128.140 162.345 ;
        RECT 128.310 162.255 128.535 162.385 ;
        RECT 128.310 161.150 128.480 162.255 ;
        RECT 128.705 162.105 129.230 162.325 ;
        RECT 128.650 161.340 128.890 161.935 ;
        RECT 129.060 161.405 129.230 162.105 ;
        RECT 129.400 161.745 129.570 162.525 ;
        RECT 129.890 162.475 130.260 162.975 ;
        RECT 130.440 162.525 130.845 162.695 ;
        RECT 131.015 162.525 131.800 162.695 ;
        RECT 130.440 162.295 130.610 162.525 ;
        RECT 129.780 161.995 130.610 162.295 ;
        RECT 130.995 162.025 131.460 162.355 ;
        RECT 129.780 161.965 129.980 161.995 ;
        RECT 130.100 161.745 130.270 161.815 ;
        RECT 129.400 161.575 130.270 161.745 ;
        RECT 129.760 161.485 130.270 161.575 ;
        RECT 128.310 161.020 128.615 161.150 ;
        RECT 129.060 161.040 129.590 161.405 ;
        RECT 127.930 160.425 128.195 160.885 ;
        RECT 128.365 160.595 128.615 161.020 ;
        RECT 129.760 160.870 129.930 161.485 ;
        RECT 128.825 160.700 129.930 160.870 ;
        RECT 130.100 160.425 130.270 161.225 ;
        RECT 130.440 160.925 130.610 161.995 ;
        RECT 130.780 161.095 130.970 161.815 ;
        RECT 131.140 161.065 131.460 162.025 ;
        RECT 131.630 162.065 131.800 162.525 ;
        RECT 132.075 162.445 132.285 162.975 ;
        RECT 132.545 162.235 132.875 162.760 ;
        RECT 133.045 162.365 133.215 162.975 ;
        RECT 133.385 162.320 133.715 162.755 ;
        RECT 134.025 162.425 134.195 162.805 ;
        RECT 134.375 162.595 134.705 162.975 ;
        RECT 133.385 162.235 133.765 162.320 ;
        RECT 134.025 162.255 134.690 162.425 ;
        RECT 134.885 162.300 135.145 162.805 ;
        RECT 132.675 162.065 132.875 162.235 ;
        RECT 133.540 162.195 133.765 162.235 ;
        RECT 131.630 161.735 132.505 162.065 ;
        RECT 132.675 161.735 133.425 162.065 ;
        RECT 130.440 160.595 130.690 160.925 ;
        RECT 131.630 160.895 131.800 161.735 ;
        RECT 132.675 161.530 132.865 161.735 ;
        RECT 133.595 161.615 133.765 162.195 ;
        RECT 133.955 161.705 134.285 162.075 ;
        RECT 134.520 162.000 134.690 162.255 ;
        RECT 133.550 161.565 133.765 161.615 ;
        RECT 131.970 161.155 132.865 161.530 ;
        RECT 133.375 161.485 133.765 161.565 ;
        RECT 134.520 161.670 134.805 162.000 ;
        RECT 134.520 161.525 134.690 161.670 ;
        RECT 130.915 160.725 131.800 160.895 ;
        RECT 131.980 160.425 132.295 160.925 ;
        RECT 132.525 160.595 132.865 161.155 ;
        RECT 133.035 160.425 133.205 161.435 ;
        RECT 133.375 160.640 133.705 161.485 ;
        RECT 134.025 161.355 134.690 161.525 ;
        RECT 134.975 161.500 135.145 162.300 ;
        RECT 135.865 162.425 136.035 162.805 ;
        RECT 136.250 162.595 136.580 162.975 ;
        RECT 135.865 162.255 136.580 162.425 ;
        RECT 135.775 161.705 136.130 162.075 ;
        RECT 136.410 162.065 136.580 162.255 ;
        RECT 136.750 162.230 137.005 162.805 ;
        RECT 136.410 161.735 136.665 162.065 ;
        RECT 136.410 161.525 136.580 161.735 ;
        RECT 134.025 160.595 134.195 161.355 ;
        RECT 134.375 160.425 134.705 161.185 ;
        RECT 134.875 160.595 135.145 161.500 ;
        RECT 135.865 161.355 136.580 161.525 ;
        RECT 136.835 161.500 137.005 162.230 ;
        RECT 137.180 162.135 137.440 162.975 ;
        RECT 137.615 162.225 138.825 162.975 ;
        RECT 135.865 160.595 136.035 161.355 ;
        RECT 136.250 160.425 136.580 161.185 ;
        RECT 136.750 160.595 137.005 161.500 ;
        RECT 137.180 160.425 137.440 161.575 ;
        RECT 137.615 161.515 138.135 162.055 ;
        RECT 138.305 161.685 138.825 162.225 ;
        RECT 137.615 160.425 138.825 161.515 ;
        RECT 13.330 160.255 138.910 160.425 ;
        RECT 13.415 159.165 14.625 160.255 ;
        RECT 14.795 159.820 20.140 160.255 ;
        RECT 20.315 159.820 25.660 160.255 ;
        RECT 13.415 158.455 13.935 158.995 ;
        RECT 14.105 158.625 14.625 159.165 ;
        RECT 13.415 157.705 14.625 158.455 ;
        RECT 16.380 158.250 16.720 159.080 ;
        RECT 18.200 158.570 18.550 159.820 ;
        RECT 21.900 158.250 22.240 159.080 ;
        RECT 23.720 158.570 24.070 159.820 ;
        RECT 26.295 159.090 26.585 160.255 ;
        RECT 26.755 159.820 32.100 160.255 ;
        RECT 14.795 157.705 20.140 158.250 ;
        RECT 20.315 157.705 25.660 158.250 ;
        RECT 26.295 157.705 26.585 158.430 ;
        RECT 28.340 158.250 28.680 159.080 ;
        RECT 30.160 158.570 30.510 159.820 ;
        RECT 32.275 159.165 33.945 160.255 ;
        RECT 32.275 158.475 33.025 158.995 ;
        RECT 33.195 158.645 33.945 159.165 ;
        RECT 34.115 159.235 34.490 160.085 ;
        RECT 34.660 159.455 34.910 160.255 ;
        RECT 35.080 159.625 35.330 160.085 ;
        RECT 35.500 159.795 35.750 160.255 ;
        RECT 35.920 159.625 36.170 160.085 ;
        RECT 36.340 159.795 36.590 160.255 ;
        RECT 36.760 159.625 37.010 160.085 ;
        RECT 37.180 159.795 37.430 160.255 ;
        RECT 37.600 159.625 37.850 160.085 ;
        RECT 35.080 159.405 37.850 159.625 ;
        RECT 38.065 159.625 38.380 160.085 ;
        RECT 38.550 159.795 38.800 160.255 ;
        RECT 38.970 159.625 39.220 160.085 ;
        RECT 39.390 159.795 39.640 160.255 ;
        RECT 39.810 159.835 41.780 160.085 ;
        RECT 39.810 159.625 40.020 159.835 ;
        RECT 41.990 159.665 42.280 160.085 ;
        RECT 38.065 159.405 40.020 159.625 ;
        RECT 40.190 159.405 42.280 159.665 ;
        RECT 42.450 159.455 42.700 160.255 ;
        RECT 35.080 159.235 35.330 159.405 ;
        RECT 41.990 159.285 42.280 159.405 ;
        RECT 42.870 159.285 43.120 160.085 ;
        RECT 43.290 159.455 43.540 160.255 ;
        RECT 43.710 159.285 44.065 160.085 ;
        RECT 44.235 159.820 49.580 160.255 ;
        RECT 34.115 159.065 35.330 159.235 ;
        RECT 35.715 159.065 39.760 159.235 ;
        RECT 39.930 159.065 41.800 159.235 ;
        RECT 41.990 159.065 44.065 159.285 ;
        RECT 34.115 158.525 34.350 159.065 ;
        RECT 35.715 158.895 35.885 159.065 ;
        RECT 39.590 158.895 39.760 159.065 ;
        RECT 41.630 158.895 41.800 159.065 ;
        RECT 34.520 158.695 35.885 158.895 ;
        RECT 36.205 158.695 39.420 158.895 ;
        RECT 39.590 158.695 41.460 158.895 ;
        RECT 41.630 158.695 43.675 158.895 ;
        RECT 43.845 158.525 44.065 159.065 ;
        RECT 26.755 157.705 32.100 158.250 ;
        RECT 32.275 157.705 33.945 158.475 ;
        RECT 34.115 158.265 35.790 158.525 ;
        RECT 35.960 158.345 37.890 158.525 ;
        RECT 35.960 158.095 36.210 158.345 ;
        RECT 34.200 157.875 36.210 158.095 ;
        RECT 36.380 157.705 36.550 158.175 ;
        RECT 36.720 157.875 37.050 158.345 ;
        RECT 37.220 157.705 37.390 158.175 ;
        RECT 37.560 157.875 37.890 158.345 ;
        RECT 38.065 157.705 38.340 158.525 ;
        RECT 38.510 158.355 42.240 158.525 ;
        RECT 38.510 158.345 41.460 158.355 ;
        RECT 38.510 157.875 38.840 158.345 ;
        RECT 39.010 157.705 39.180 158.175 ;
        RECT 39.350 157.875 39.680 158.345 ;
        RECT 39.850 157.705 40.020 158.175 ;
        RECT 40.190 157.875 40.520 158.345 ;
        RECT 40.690 157.705 40.860 158.175 ;
        RECT 41.030 157.875 41.360 158.345 ;
        RECT 41.530 157.705 41.800 158.175 ;
        RECT 41.990 158.095 42.240 158.355 ;
        RECT 42.410 158.265 44.065 158.525 ;
        RECT 45.820 158.250 46.160 159.080 ;
        RECT 47.640 158.570 47.990 159.820 ;
        RECT 49.755 159.165 51.425 160.255 ;
        RECT 49.755 158.475 50.505 158.995 ;
        RECT 50.675 158.645 51.425 159.165 ;
        RECT 52.055 159.090 52.345 160.255 ;
        RECT 52.515 159.820 57.860 160.255 ;
        RECT 58.035 159.820 63.380 160.255 ;
        RECT 41.990 157.925 44.000 158.095 ;
        RECT 44.235 157.705 49.580 158.250 ;
        RECT 49.755 157.705 51.425 158.475 ;
        RECT 52.055 157.705 52.345 158.430 ;
        RECT 54.100 158.250 54.440 159.080 ;
        RECT 55.920 158.570 56.270 159.820 ;
        RECT 59.620 158.250 59.960 159.080 ;
        RECT 61.440 158.570 61.790 159.820 ;
        RECT 63.555 159.165 66.145 160.255 ;
        RECT 63.555 158.475 64.765 158.995 ;
        RECT 64.935 158.645 66.145 159.165 ;
        RECT 66.780 159.115 67.115 160.085 ;
        RECT 67.285 159.115 67.455 160.255 ;
        RECT 67.625 159.915 69.655 160.085 ;
        RECT 52.515 157.705 57.860 158.250 ;
        RECT 58.035 157.705 63.380 158.250 ;
        RECT 63.555 157.705 66.145 158.475 ;
        RECT 66.780 158.445 66.950 159.115 ;
        RECT 67.625 158.945 67.795 159.915 ;
        RECT 67.120 158.615 67.375 158.945 ;
        RECT 67.600 158.615 67.795 158.945 ;
        RECT 67.965 159.575 69.090 159.745 ;
        RECT 67.205 158.445 67.375 158.615 ;
        RECT 67.965 158.445 68.135 159.575 ;
        RECT 66.780 157.875 67.035 158.445 ;
        RECT 67.205 158.275 68.135 158.445 ;
        RECT 68.305 159.235 69.315 159.405 ;
        RECT 68.305 158.435 68.475 159.235 ;
        RECT 68.680 158.555 68.955 159.035 ;
        RECT 68.675 158.385 68.955 158.555 ;
        RECT 67.960 158.240 68.135 158.275 ;
        RECT 67.205 157.705 67.535 158.105 ;
        RECT 67.960 157.875 68.490 158.240 ;
        RECT 68.680 157.875 68.955 158.385 ;
        RECT 69.125 157.875 69.315 159.235 ;
        RECT 69.485 159.250 69.655 159.915 ;
        RECT 69.825 159.495 69.995 160.255 ;
        RECT 70.230 159.495 70.745 159.905 ;
        RECT 69.485 159.060 70.235 159.250 ;
        RECT 70.405 158.685 70.745 159.495 ;
        RECT 70.915 159.165 72.125 160.255 ;
        RECT 69.515 158.515 70.745 158.685 ;
        RECT 69.495 157.705 70.005 158.240 ;
        RECT 70.225 157.910 70.470 158.515 ;
        RECT 70.915 158.455 71.435 158.995 ;
        RECT 71.605 158.625 72.125 159.165 ;
        RECT 72.295 159.115 72.680 160.085 ;
        RECT 72.850 159.795 73.175 160.255 ;
        RECT 73.695 159.625 73.975 160.085 ;
        RECT 72.850 159.405 73.975 159.625 ;
        RECT 70.915 157.705 72.125 158.455 ;
        RECT 72.295 158.445 72.575 159.115 ;
        RECT 72.850 158.945 73.300 159.405 ;
        RECT 74.165 159.235 74.565 160.085 ;
        RECT 74.965 159.795 75.235 160.255 ;
        RECT 75.405 159.625 75.690 160.085 ;
        RECT 72.745 158.615 73.300 158.945 ;
        RECT 73.470 158.675 74.565 159.235 ;
        RECT 72.850 158.505 73.300 158.615 ;
        RECT 72.295 157.875 72.680 158.445 ;
        RECT 72.850 158.335 73.975 158.505 ;
        RECT 72.850 157.705 73.175 158.165 ;
        RECT 73.695 157.875 73.975 158.335 ;
        RECT 74.165 157.875 74.565 158.675 ;
        RECT 74.735 159.405 75.690 159.625 ;
        RECT 74.735 158.505 74.945 159.405 ;
        RECT 75.115 158.675 75.805 159.235 ;
        RECT 75.975 159.165 77.645 160.255 ;
        RECT 74.735 158.335 75.690 158.505 ;
        RECT 74.965 157.705 75.235 158.165 ;
        RECT 75.405 157.875 75.690 158.335 ;
        RECT 75.975 158.475 76.725 158.995 ;
        RECT 76.895 158.645 77.645 159.165 ;
        RECT 77.815 159.090 78.105 160.255 ;
        RECT 78.275 159.820 83.620 160.255 ;
        RECT 75.975 157.705 77.645 158.475 ;
        RECT 77.815 157.705 78.105 158.430 ;
        RECT 79.860 158.250 80.200 159.080 ;
        RECT 81.680 158.570 82.030 159.820 ;
        RECT 83.795 159.165 85.005 160.255 ;
        RECT 83.795 158.455 84.315 158.995 ;
        RECT 84.485 158.625 85.005 159.165 ;
        RECT 85.175 159.495 85.690 159.905 ;
        RECT 85.925 159.495 86.095 160.255 ;
        RECT 86.265 159.915 88.295 160.085 ;
        RECT 85.175 158.685 85.515 159.495 ;
        RECT 86.265 159.250 86.435 159.915 ;
        RECT 86.830 159.575 87.955 159.745 ;
        RECT 85.685 159.060 86.435 159.250 ;
        RECT 86.605 159.235 87.615 159.405 ;
        RECT 85.175 158.515 86.405 158.685 ;
        RECT 78.275 157.705 83.620 158.250 ;
        RECT 83.795 157.705 85.005 158.455 ;
        RECT 85.450 157.910 85.695 158.515 ;
        RECT 85.915 157.705 86.425 158.240 ;
        RECT 86.605 157.875 86.795 159.235 ;
        RECT 86.965 158.215 87.240 159.035 ;
        RECT 87.445 158.435 87.615 159.235 ;
        RECT 87.785 158.445 87.955 159.575 ;
        RECT 88.125 158.945 88.295 159.915 ;
        RECT 88.465 159.115 88.635 160.255 ;
        RECT 88.805 159.115 89.140 160.085 ;
        RECT 89.315 159.165 91.905 160.255 ;
        RECT 92.625 159.585 92.795 160.085 ;
        RECT 92.965 159.755 93.295 160.255 ;
        RECT 92.625 159.415 93.290 159.585 ;
        RECT 88.125 158.615 88.320 158.945 ;
        RECT 88.545 158.615 88.800 158.945 ;
        RECT 88.545 158.445 88.715 158.615 ;
        RECT 88.970 158.445 89.140 159.115 ;
        RECT 87.785 158.275 88.715 158.445 ;
        RECT 87.785 158.240 87.960 158.275 ;
        RECT 86.965 158.045 87.245 158.215 ;
        RECT 86.965 157.875 87.240 158.045 ;
        RECT 87.430 157.875 87.960 158.240 ;
        RECT 88.385 157.705 88.715 158.105 ;
        RECT 88.885 157.875 89.140 158.445 ;
        RECT 89.315 158.475 90.525 158.995 ;
        RECT 90.695 158.645 91.905 159.165 ;
        RECT 92.540 158.595 92.890 159.245 ;
        RECT 89.315 157.705 91.905 158.475 ;
        RECT 93.060 158.425 93.290 159.415 ;
        RECT 92.625 158.255 93.290 158.425 ;
        RECT 92.625 157.965 92.795 158.255 ;
        RECT 92.965 157.705 93.295 158.085 ;
        RECT 93.465 157.965 93.650 160.085 ;
        RECT 93.890 159.795 94.155 160.255 ;
        RECT 94.325 159.660 94.575 160.085 ;
        RECT 94.785 159.810 95.890 159.980 ;
        RECT 94.270 159.530 94.575 159.660 ;
        RECT 93.820 158.335 94.100 159.285 ;
        RECT 94.270 158.425 94.440 159.530 ;
        RECT 94.610 158.745 94.850 159.340 ;
        RECT 95.020 159.275 95.550 159.640 ;
        RECT 95.020 158.575 95.190 159.275 ;
        RECT 95.720 159.195 95.890 159.810 ;
        RECT 96.060 159.455 96.230 160.255 ;
        RECT 96.400 159.755 96.650 160.085 ;
        RECT 96.875 159.785 97.760 159.955 ;
        RECT 95.720 159.105 96.230 159.195 ;
        RECT 94.270 158.295 94.495 158.425 ;
        RECT 94.665 158.355 95.190 158.575 ;
        RECT 95.360 158.935 96.230 159.105 ;
        RECT 93.905 157.705 94.155 158.165 ;
        RECT 94.325 158.155 94.495 158.295 ;
        RECT 95.360 158.155 95.530 158.935 ;
        RECT 96.060 158.865 96.230 158.935 ;
        RECT 95.740 158.685 95.940 158.715 ;
        RECT 96.400 158.685 96.570 159.755 ;
        RECT 96.740 158.865 96.930 159.585 ;
        RECT 95.740 158.385 96.570 158.685 ;
        RECT 97.100 158.655 97.420 159.615 ;
        RECT 94.325 157.985 94.660 158.155 ;
        RECT 94.855 157.985 95.530 158.155 ;
        RECT 95.850 157.705 96.220 158.205 ;
        RECT 96.400 158.155 96.570 158.385 ;
        RECT 96.955 158.325 97.420 158.655 ;
        RECT 97.590 158.945 97.760 159.785 ;
        RECT 97.940 159.755 98.255 160.255 ;
        RECT 98.485 159.525 98.825 160.085 ;
        RECT 97.930 159.150 98.825 159.525 ;
        RECT 98.995 159.245 99.165 160.255 ;
        RECT 98.635 158.945 98.825 159.150 ;
        RECT 99.335 159.195 99.665 160.040 ;
        RECT 99.335 159.115 99.725 159.195 ;
        RECT 99.895 159.165 103.405 160.255 ;
        RECT 99.510 159.065 99.725 159.115 ;
        RECT 97.590 158.615 98.465 158.945 ;
        RECT 98.635 158.615 99.385 158.945 ;
        RECT 97.590 158.155 97.760 158.615 ;
        RECT 98.635 158.445 98.835 158.615 ;
        RECT 99.555 158.485 99.725 159.065 ;
        RECT 99.500 158.445 99.725 158.485 ;
        RECT 96.400 157.985 96.805 158.155 ;
        RECT 96.975 157.985 97.760 158.155 ;
        RECT 98.035 157.705 98.245 158.235 ;
        RECT 98.505 157.920 98.835 158.445 ;
        RECT 99.345 158.360 99.725 158.445 ;
        RECT 99.895 158.475 101.545 158.995 ;
        RECT 101.715 158.645 103.405 159.165 ;
        RECT 103.575 159.090 103.865 160.255 ;
        RECT 104.150 159.625 104.435 160.085 ;
        RECT 104.605 159.795 104.875 160.255 ;
        RECT 104.150 159.405 105.105 159.625 ;
        RECT 104.035 158.675 104.725 159.235 ;
        RECT 104.895 158.505 105.105 159.405 ;
        RECT 99.005 157.705 99.175 158.315 ;
        RECT 99.345 157.925 99.675 158.360 ;
        RECT 99.895 157.705 103.405 158.475 ;
        RECT 103.575 157.705 103.865 158.430 ;
        RECT 104.150 158.335 105.105 158.505 ;
        RECT 105.275 159.235 105.675 160.085 ;
        RECT 105.865 159.625 106.145 160.085 ;
        RECT 106.665 159.795 106.990 160.255 ;
        RECT 105.865 159.405 106.990 159.625 ;
        RECT 105.275 158.675 106.370 159.235 ;
        RECT 106.540 158.945 106.990 159.405 ;
        RECT 107.160 159.115 107.545 160.085 ;
        RECT 107.720 159.115 108.040 160.255 ;
        RECT 104.150 157.875 104.435 158.335 ;
        RECT 104.605 157.705 104.875 158.165 ;
        RECT 105.275 157.875 105.675 158.675 ;
        RECT 106.540 158.615 107.095 158.945 ;
        RECT 106.540 158.505 106.990 158.615 ;
        RECT 105.865 158.335 106.990 158.505 ;
        RECT 107.265 158.445 107.545 159.115 ;
        RECT 108.220 158.945 108.415 159.995 ;
        RECT 108.595 159.405 108.925 160.085 ;
        RECT 109.125 159.455 109.380 160.255 ;
        RECT 108.595 159.125 108.945 159.405 ;
        RECT 107.780 158.895 108.040 158.945 ;
        RECT 107.775 158.725 108.040 158.895 ;
        RECT 107.780 158.615 108.040 158.725 ;
        RECT 108.220 158.615 108.605 158.945 ;
        RECT 108.775 158.745 108.945 159.125 ;
        RECT 109.135 158.915 109.380 159.275 ;
        RECT 109.555 159.115 109.835 160.255 ;
        RECT 110.005 159.105 110.335 160.085 ;
        RECT 110.505 159.115 110.765 160.255 ;
        RECT 111.970 159.625 112.255 160.085 ;
        RECT 112.425 159.795 112.695 160.255 ;
        RECT 111.970 159.405 112.925 159.625 ;
        RECT 108.775 158.575 109.295 158.745 ;
        RECT 109.565 158.675 109.900 158.945 ;
        RECT 105.865 157.875 106.145 158.335 ;
        RECT 106.665 157.705 106.990 158.165 ;
        RECT 107.160 157.875 107.545 158.445 ;
        RECT 109.125 158.555 109.295 158.575 ;
        RECT 107.720 158.235 108.935 158.405 ;
        RECT 107.720 157.885 108.010 158.235 ;
        RECT 108.205 157.705 108.535 158.065 ;
        RECT 108.705 157.930 108.935 158.235 ;
        RECT 109.125 158.385 109.325 158.555 ;
        RECT 110.070 158.505 110.240 159.105 ;
        RECT 110.410 158.695 110.745 158.945 ;
        RECT 111.855 158.675 112.545 159.235 ;
        RECT 112.715 158.505 112.925 159.405 ;
        RECT 109.125 158.010 109.295 158.385 ;
        RECT 109.555 157.705 109.865 158.505 ;
        RECT 110.070 157.875 110.765 158.505 ;
        RECT 111.970 158.335 112.925 158.505 ;
        RECT 113.095 159.235 113.495 160.085 ;
        RECT 113.685 159.625 113.965 160.085 ;
        RECT 114.485 159.795 114.810 160.255 ;
        RECT 113.685 159.405 114.810 159.625 ;
        RECT 113.095 158.675 114.190 159.235 ;
        RECT 114.360 158.945 114.810 159.405 ;
        RECT 114.980 159.115 115.365 160.085 ;
        RECT 111.970 157.875 112.255 158.335 ;
        RECT 112.425 157.705 112.695 158.165 ;
        RECT 113.095 157.875 113.495 158.675 ;
        RECT 114.360 158.615 114.915 158.945 ;
        RECT 114.360 158.505 114.810 158.615 ;
        RECT 113.685 158.335 114.810 158.505 ;
        RECT 115.085 158.445 115.365 159.115 ;
        RECT 113.685 157.875 113.965 158.335 ;
        RECT 114.485 157.705 114.810 158.165 ;
        RECT 114.980 157.875 115.365 158.445 ;
        RECT 115.535 159.405 115.795 160.085 ;
        RECT 115.965 159.475 116.215 160.255 ;
        RECT 116.465 159.705 116.715 160.085 ;
        RECT 116.885 159.875 117.240 160.255 ;
        RECT 118.245 159.865 118.580 160.085 ;
        RECT 117.845 159.705 118.075 159.745 ;
        RECT 116.465 159.505 118.075 159.705 ;
        RECT 116.465 159.495 117.300 159.505 ;
        RECT 117.890 159.415 118.075 159.505 ;
        RECT 115.535 158.215 115.705 159.405 ;
        RECT 117.405 159.305 117.735 159.335 ;
        RECT 115.935 159.245 117.735 159.305 ;
        RECT 118.325 159.245 118.580 159.865 ;
        RECT 115.875 159.135 118.580 159.245 ;
        RECT 119.225 159.145 119.520 160.255 ;
        RECT 115.875 159.100 116.075 159.135 ;
        RECT 115.875 158.525 116.045 159.100 ;
        RECT 117.405 159.075 118.580 159.135 ;
        RECT 116.275 158.660 116.685 158.965 ;
        RECT 119.700 158.945 119.950 160.080 ;
        RECT 120.120 159.145 120.380 160.255 ;
        RECT 120.550 159.355 120.810 160.080 ;
        RECT 120.980 159.525 121.240 160.255 ;
        RECT 121.410 159.355 121.670 160.080 ;
        RECT 121.840 159.525 122.100 160.255 ;
        RECT 122.270 159.355 122.530 160.080 ;
        RECT 122.700 159.525 122.960 160.255 ;
        RECT 123.130 159.355 123.390 160.080 ;
        RECT 123.560 159.525 123.855 160.255 ;
        RECT 125.195 159.495 125.710 159.905 ;
        RECT 125.945 159.495 126.115 160.255 ;
        RECT 126.285 159.915 128.315 160.085 ;
        RECT 120.550 159.115 123.860 159.355 ;
        RECT 116.855 158.695 117.185 158.905 ;
        RECT 115.875 158.405 116.145 158.525 ;
        RECT 115.875 158.360 116.720 158.405 ;
        RECT 115.965 158.235 116.720 158.360 ;
        RECT 116.975 158.295 117.185 158.695 ;
        RECT 117.430 158.695 117.905 158.905 ;
        RECT 118.095 158.695 118.585 158.895 ;
        RECT 117.430 158.295 117.650 158.695 ;
        RECT 115.535 158.205 115.765 158.215 ;
        RECT 115.535 157.875 115.795 158.205 ;
        RECT 116.550 158.085 116.720 158.235 ;
        RECT 115.965 157.705 116.295 158.065 ;
        RECT 116.550 157.875 117.850 158.085 ;
        RECT 118.125 157.705 118.580 158.470 ;
        RECT 119.215 158.335 119.530 158.945 ;
        RECT 119.700 158.695 122.720 158.945 ;
        RECT 119.275 157.705 119.520 158.165 ;
        RECT 119.700 157.885 119.950 158.695 ;
        RECT 122.890 158.525 123.860 159.115 ;
        RECT 120.550 158.355 123.860 158.525 ;
        RECT 125.195 158.685 125.535 159.495 ;
        RECT 126.285 159.250 126.455 159.915 ;
        RECT 126.850 159.575 127.975 159.745 ;
        RECT 125.705 159.060 126.455 159.250 ;
        RECT 126.625 159.235 127.635 159.405 ;
        RECT 125.195 158.515 126.425 158.685 ;
        RECT 120.120 157.705 120.380 158.230 ;
        RECT 120.550 157.900 120.810 158.355 ;
        RECT 120.980 157.705 121.240 158.185 ;
        RECT 121.410 157.900 121.670 158.355 ;
        RECT 121.840 157.705 122.100 158.185 ;
        RECT 122.270 157.900 122.530 158.355 ;
        RECT 122.700 157.705 122.960 158.185 ;
        RECT 123.130 157.900 123.390 158.355 ;
        RECT 123.560 157.705 123.860 158.185 ;
        RECT 125.470 157.910 125.715 158.515 ;
        RECT 125.935 157.705 126.445 158.240 ;
        RECT 126.625 157.875 126.815 159.235 ;
        RECT 126.985 158.215 127.260 159.035 ;
        RECT 127.465 158.435 127.635 159.235 ;
        RECT 127.805 158.445 127.975 159.575 ;
        RECT 128.145 158.945 128.315 159.915 ;
        RECT 128.485 159.115 128.655 160.255 ;
        RECT 128.825 159.115 129.160 160.085 ;
        RECT 128.145 158.615 128.340 158.945 ;
        RECT 128.565 158.615 128.820 158.945 ;
        RECT 128.565 158.445 128.735 158.615 ;
        RECT 128.990 158.445 129.160 159.115 ;
        RECT 129.335 159.090 129.625 160.255 ;
        RECT 129.885 159.585 130.055 160.085 ;
        RECT 130.225 159.755 130.555 160.255 ;
        RECT 129.885 159.415 130.550 159.585 ;
        RECT 129.800 158.595 130.150 159.245 ;
        RECT 127.805 158.275 128.735 158.445 ;
        RECT 127.805 158.240 127.980 158.275 ;
        RECT 126.985 158.045 127.265 158.215 ;
        RECT 126.985 157.875 127.260 158.045 ;
        RECT 127.450 157.875 127.980 158.240 ;
        RECT 128.405 157.705 128.735 158.105 ;
        RECT 128.905 157.875 129.160 158.445 ;
        RECT 129.335 157.705 129.625 158.430 ;
        RECT 130.320 158.425 130.550 159.415 ;
        RECT 129.885 158.255 130.550 158.425 ;
        RECT 129.885 157.965 130.055 158.255 ;
        RECT 130.225 157.705 130.555 158.085 ;
        RECT 130.725 157.965 130.910 160.085 ;
        RECT 131.150 159.795 131.415 160.255 ;
        RECT 131.585 159.660 131.835 160.085 ;
        RECT 132.045 159.810 133.150 159.980 ;
        RECT 131.530 159.530 131.835 159.660 ;
        RECT 131.080 158.335 131.360 159.285 ;
        RECT 131.530 158.425 131.700 159.530 ;
        RECT 131.870 158.745 132.110 159.340 ;
        RECT 132.280 159.275 132.810 159.640 ;
        RECT 132.280 158.575 132.450 159.275 ;
        RECT 132.980 159.195 133.150 159.810 ;
        RECT 133.320 159.455 133.490 160.255 ;
        RECT 133.660 159.755 133.910 160.085 ;
        RECT 134.135 159.785 135.020 159.955 ;
        RECT 132.980 159.105 133.490 159.195 ;
        RECT 131.530 158.295 131.755 158.425 ;
        RECT 131.925 158.355 132.450 158.575 ;
        RECT 132.620 158.935 133.490 159.105 ;
        RECT 131.165 157.705 131.415 158.165 ;
        RECT 131.585 158.155 131.755 158.295 ;
        RECT 132.620 158.155 132.790 158.935 ;
        RECT 133.320 158.865 133.490 158.935 ;
        RECT 133.000 158.685 133.200 158.715 ;
        RECT 133.660 158.685 133.830 159.755 ;
        RECT 134.000 158.865 134.190 159.585 ;
        RECT 133.000 158.385 133.830 158.685 ;
        RECT 134.360 158.655 134.680 159.615 ;
        RECT 131.585 157.985 131.920 158.155 ;
        RECT 132.115 157.985 132.790 158.155 ;
        RECT 133.110 157.705 133.480 158.205 ;
        RECT 133.660 158.155 133.830 158.385 ;
        RECT 134.215 158.325 134.680 158.655 ;
        RECT 134.850 158.945 135.020 159.785 ;
        RECT 135.200 159.755 135.515 160.255 ;
        RECT 135.745 159.525 136.085 160.085 ;
        RECT 135.190 159.150 136.085 159.525 ;
        RECT 136.255 159.245 136.425 160.255 ;
        RECT 135.895 158.945 136.085 159.150 ;
        RECT 136.595 159.195 136.925 160.040 ;
        RECT 136.595 159.115 136.985 159.195 ;
        RECT 136.770 159.065 136.985 159.115 ;
        RECT 134.850 158.615 135.725 158.945 ;
        RECT 135.895 158.615 136.645 158.945 ;
        RECT 134.850 158.155 135.020 158.615 ;
        RECT 135.895 158.445 136.095 158.615 ;
        RECT 136.815 158.485 136.985 159.065 ;
        RECT 137.615 159.165 138.825 160.255 ;
        RECT 137.615 158.625 138.135 159.165 ;
        RECT 136.760 158.445 136.985 158.485 ;
        RECT 138.305 158.455 138.825 158.995 ;
        RECT 133.660 157.985 134.065 158.155 ;
        RECT 134.235 157.985 135.020 158.155 ;
        RECT 135.295 157.705 135.505 158.235 ;
        RECT 135.765 157.920 136.095 158.445 ;
        RECT 136.605 158.360 136.985 158.445 ;
        RECT 136.265 157.705 136.435 158.315 ;
        RECT 136.605 157.925 136.935 158.360 ;
        RECT 137.615 157.705 138.825 158.455 ;
        RECT 13.330 157.535 138.910 157.705 ;
        RECT 13.415 156.785 14.625 157.535 ;
        RECT 14.885 156.985 15.055 157.365 ;
        RECT 15.270 157.155 15.600 157.535 ;
        RECT 14.885 156.815 15.600 156.985 ;
        RECT 13.415 156.245 13.935 156.785 ;
        RECT 14.105 156.075 14.625 156.615 ;
        RECT 14.795 156.265 15.150 156.635 ;
        RECT 15.430 156.625 15.600 156.815 ;
        RECT 15.770 156.790 16.025 157.365 ;
        RECT 15.430 156.295 15.685 156.625 ;
        RECT 15.430 156.085 15.600 156.295 ;
        RECT 13.415 154.985 14.625 156.075 ;
        RECT 14.885 155.915 15.600 156.085 ;
        RECT 15.855 156.060 16.025 156.790 ;
        RECT 16.200 156.695 16.460 157.535 ;
        RECT 16.635 156.765 19.225 157.535 ;
        RECT 19.485 156.985 19.655 157.275 ;
        RECT 19.825 157.155 20.155 157.535 ;
        RECT 19.485 156.815 20.150 156.985 ;
        RECT 16.635 156.245 17.845 156.765 ;
        RECT 14.885 155.155 15.055 155.915 ;
        RECT 15.270 154.985 15.600 155.745 ;
        RECT 15.770 155.155 16.025 156.060 ;
        RECT 16.200 154.985 16.460 156.135 ;
        RECT 18.015 156.075 19.225 156.595 ;
        RECT 16.635 154.985 19.225 156.075 ;
        RECT 19.400 155.995 19.750 156.645 ;
        RECT 19.920 155.825 20.150 156.815 ;
        RECT 19.485 155.655 20.150 155.825 ;
        RECT 19.485 155.155 19.655 155.655 ;
        RECT 19.825 154.985 20.155 155.485 ;
        RECT 20.325 155.155 20.510 157.275 ;
        RECT 20.765 157.075 21.015 157.535 ;
        RECT 21.185 157.085 21.520 157.255 ;
        RECT 21.715 157.085 22.390 157.255 ;
        RECT 21.185 156.945 21.355 157.085 ;
        RECT 20.680 155.955 20.960 156.905 ;
        RECT 21.130 156.815 21.355 156.945 ;
        RECT 21.130 155.710 21.300 156.815 ;
        RECT 21.525 156.665 22.050 156.885 ;
        RECT 21.470 155.900 21.710 156.495 ;
        RECT 21.880 155.965 22.050 156.665 ;
        RECT 22.220 156.305 22.390 157.085 ;
        RECT 22.710 157.035 23.080 157.535 ;
        RECT 23.260 157.085 23.665 157.255 ;
        RECT 23.835 157.085 24.620 157.255 ;
        RECT 23.260 156.855 23.430 157.085 ;
        RECT 22.600 156.555 23.430 156.855 ;
        RECT 23.815 156.585 24.280 156.915 ;
        RECT 22.600 156.525 22.800 156.555 ;
        RECT 22.920 156.305 23.090 156.375 ;
        RECT 22.220 156.135 23.090 156.305 ;
        RECT 22.580 156.045 23.090 156.135 ;
        RECT 21.130 155.580 21.435 155.710 ;
        RECT 21.880 155.600 22.410 155.965 ;
        RECT 20.750 154.985 21.015 155.445 ;
        RECT 21.185 155.155 21.435 155.580 ;
        RECT 22.580 155.430 22.750 156.045 ;
        RECT 21.645 155.260 22.750 155.430 ;
        RECT 22.920 154.985 23.090 155.785 ;
        RECT 23.260 155.485 23.430 156.555 ;
        RECT 23.600 155.655 23.790 156.375 ;
        RECT 23.960 155.625 24.280 156.585 ;
        RECT 24.450 156.625 24.620 157.085 ;
        RECT 24.895 157.005 25.105 157.535 ;
        RECT 25.365 156.795 25.695 157.320 ;
        RECT 25.865 156.925 26.035 157.535 ;
        RECT 26.205 156.880 26.535 157.315 ;
        RECT 27.675 156.895 28.015 157.300 ;
        RECT 28.185 157.065 28.355 157.535 ;
        RECT 28.525 156.895 28.775 157.300 ;
        RECT 26.205 156.795 26.585 156.880 ;
        RECT 25.495 156.625 25.695 156.795 ;
        RECT 26.360 156.755 26.585 156.795 ;
        RECT 24.450 156.295 25.325 156.625 ;
        RECT 25.495 156.295 26.245 156.625 ;
        RECT 23.260 155.155 23.510 155.485 ;
        RECT 24.450 155.455 24.620 156.295 ;
        RECT 25.495 156.090 25.685 156.295 ;
        RECT 26.415 156.175 26.585 156.755 ;
        RECT 27.675 156.715 28.775 156.895 ;
        RECT 28.945 156.930 29.195 157.300 ;
        RECT 29.365 157.055 29.810 157.225 ;
        RECT 29.980 157.195 30.200 157.240 ;
        RECT 28.945 156.545 29.115 156.930 ;
        RECT 26.370 156.125 26.585 156.175 ;
        RECT 24.790 155.715 25.685 156.090 ;
        RECT 26.195 156.045 26.585 156.125 ;
        RECT 23.735 155.285 24.620 155.455 ;
        RECT 24.800 154.985 25.115 155.485 ;
        RECT 25.345 155.155 25.685 155.715 ;
        RECT 25.855 154.985 26.025 155.995 ;
        RECT 26.195 155.200 26.525 156.045 ;
        RECT 27.675 155.975 28.020 156.545 ;
        RECT 28.190 156.295 28.750 156.545 ;
        RECT 28.920 156.375 29.115 156.545 ;
        RECT 27.675 154.985 28.020 155.805 ;
        RECT 28.190 155.195 28.365 156.295 ;
        RECT 28.920 156.125 29.090 156.375 ;
        RECT 29.365 156.265 29.535 157.055 ;
        RECT 29.980 157.025 30.205 157.195 ;
        RECT 29.980 156.885 30.200 157.025 ;
        RECT 29.705 156.715 30.200 156.885 ;
        RECT 30.480 156.870 30.650 157.535 ;
        RECT 30.845 156.795 31.185 157.365 ;
        RECT 29.705 156.520 29.880 156.715 ;
        RECT 30.050 156.345 30.500 156.545 ;
        RECT 28.535 155.735 29.090 156.125 ;
        RECT 29.260 156.125 29.535 156.265 ;
        RECT 30.670 156.175 30.840 156.625 ;
        RECT 29.260 155.905 30.275 156.125 ;
        RECT 30.445 156.005 30.840 156.175 ;
        RECT 30.445 155.735 30.615 156.005 ;
        RECT 31.010 155.825 31.185 156.795 ;
        RECT 31.355 156.765 34.865 157.535 ;
        RECT 35.960 157.030 36.295 157.535 ;
        RECT 36.465 156.965 36.705 157.340 ;
        RECT 36.985 157.205 37.155 157.350 ;
        RECT 36.985 157.010 37.360 157.205 ;
        RECT 37.720 157.040 38.115 157.535 ;
        RECT 31.355 156.245 33.005 156.765 ;
        RECT 33.175 156.075 34.865 156.595 ;
        RECT 28.535 155.565 30.615 155.735 ;
        RECT 28.535 155.330 28.865 155.565 ;
        RECT 29.155 154.985 29.555 155.385 ;
        RECT 30.425 154.985 30.755 155.385 ;
        RECT 30.925 155.155 31.185 155.825 ;
        RECT 31.355 154.985 34.865 156.075 ;
        RECT 36.015 156.005 36.315 156.855 ;
        RECT 36.485 156.815 36.705 156.965 ;
        RECT 36.485 156.485 37.020 156.815 ;
        RECT 37.190 156.675 37.360 157.010 ;
        RECT 38.285 156.845 38.525 157.365 ;
        RECT 36.485 155.835 36.720 156.485 ;
        RECT 37.190 156.315 38.175 156.675 ;
        RECT 36.045 155.605 36.720 155.835 ;
        RECT 36.890 156.295 38.175 156.315 ;
        RECT 36.890 156.145 37.750 156.295 ;
        RECT 36.045 155.175 36.215 155.605 ;
        RECT 36.385 154.985 36.715 155.435 ;
        RECT 36.890 155.200 37.175 156.145 ;
        RECT 38.350 156.040 38.525 156.845 ;
        RECT 39.175 156.810 39.465 157.535 ;
        RECT 39.800 157.025 40.040 157.535 ;
        RECT 40.220 157.025 40.500 157.355 ;
        RECT 40.730 157.025 40.945 157.535 ;
        RECT 39.695 156.295 40.050 156.855 ;
        RECT 37.350 155.665 38.045 155.975 ;
        RECT 37.355 154.985 38.040 155.455 ;
        RECT 38.220 155.255 38.525 156.040 ;
        RECT 39.175 154.985 39.465 156.150 ;
        RECT 40.220 156.125 40.390 157.025 ;
        RECT 40.560 156.295 40.825 156.855 ;
        RECT 41.115 156.795 41.730 157.365 ;
        RECT 41.935 156.990 47.280 157.535 ;
        RECT 47.455 156.990 52.800 157.535 ;
        RECT 52.975 156.990 58.320 157.535 ;
        RECT 58.495 156.990 63.840 157.535 ;
        RECT 41.075 156.125 41.245 156.625 ;
        RECT 39.820 155.955 41.245 156.125 ;
        RECT 39.820 155.780 40.210 155.955 ;
        RECT 40.695 154.985 41.025 155.785 ;
        RECT 41.415 155.775 41.730 156.795 ;
        RECT 43.520 156.160 43.860 156.990 ;
        RECT 41.195 155.155 41.730 155.775 ;
        RECT 45.340 155.420 45.690 156.670 ;
        RECT 49.040 156.160 49.380 156.990 ;
        RECT 50.860 155.420 51.210 156.670 ;
        RECT 54.560 156.160 54.900 156.990 ;
        RECT 56.380 155.420 56.730 156.670 ;
        RECT 60.080 156.160 60.420 156.990 ;
        RECT 64.935 156.810 65.225 157.535 ;
        RECT 65.485 156.985 65.655 157.275 ;
        RECT 65.825 157.155 66.155 157.535 ;
        RECT 65.485 156.815 66.150 156.985 ;
        RECT 61.900 155.420 62.250 156.670 ;
        RECT 41.935 154.985 47.280 155.420 ;
        RECT 47.455 154.985 52.800 155.420 ;
        RECT 52.975 154.985 58.320 155.420 ;
        RECT 58.495 154.985 63.840 155.420 ;
        RECT 64.935 154.985 65.225 156.150 ;
        RECT 65.400 155.995 65.750 156.645 ;
        RECT 65.920 155.825 66.150 156.815 ;
        RECT 65.485 155.655 66.150 155.825 ;
        RECT 65.485 155.155 65.655 155.655 ;
        RECT 65.825 154.985 66.155 155.485 ;
        RECT 66.325 155.155 66.510 157.275 ;
        RECT 66.765 157.075 67.015 157.535 ;
        RECT 67.185 157.085 67.520 157.255 ;
        RECT 67.715 157.085 68.390 157.255 ;
        RECT 67.185 156.945 67.355 157.085 ;
        RECT 66.680 155.955 66.960 156.905 ;
        RECT 67.130 156.815 67.355 156.945 ;
        RECT 67.130 155.710 67.300 156.815 ;
        RECT 67.525 156.665 68.050 156.885 ;
        RECT 67.470 155.900 67.710 156.495 ;
        RECT 67.880 155.965 68.050 156.665 ;
        RECT 68.220 156.305 68.390 157.085 ;
        RECT 68.710 157.035 69.080 157.535 ;
        RECT 69.260 157.085 69.665 157.255 ;
        RECT 69.835 157.085 70.620 157.255 ;
        RECT 69.260 156.855 69.430 157.085 ;
        RECT 68.600 156.555 69.430 156.855 ;
        RECT 69.815 156.585 70.280 156.915 ;
        RECT 68.600 156.525 68.800 156.555 ;
        RECT 68.920 156.305 69.090 156.375 ;
        RECT 68.220 156.135 69.090 156.305 ;
        RECT 68.580 156.045 69.090 156.135 ;
        RECT 67.130 155.580 67.435 155.710 ;
        RECT 67.880 155.600 68.410 155.965 ;
        RECT 66.750 154.985 67.015 155.445 ;
        RECT 67.185 155.155 67.435 155.580 ;
        RECT 68.580 155.430 68.750 156.045 ;
        RECT 67.645 155.260 68.750 155.430 ;
        RECT 68.920 154.985 69.090 155.785 ;
        RECT 69.260 155.485 69.430 156.555 ;
        RECT 69.600 155.655 69.790 156.375 ;
        RECT 69.960 155.625 70.280 156.585 ;
        RECT 70.450 156.625 70.620 157.085 ;
        RECT 70.895 157.005 71.105 157.535 ;
        RECT 71.365 156.795 71.695 157.320 ;
        RECT 71.865 156.925 72.035 157.535 ;
        RECT 72.205 156.880 72.535 157.315 ;
        RECT 72.205 156.795 72.585 156.880 ;
        RECT 71.495 156.625 71.695 156.795 ;
        RECT 72.360 156.755 72.585 156.795 ;
        RECT 70.450 156.295 71.325 156.625 ;
        RECT 71.495 156.295 72.245 156.625 ;
        RECT 69.260 155.155 69.510 155.485 ;
        RECT 70.450 155.455 70.620 156.295 ;
        RECT 71.495 156.090 71.685 156.295 ;
        RECT 72.415 156.175 72.585 156.755 ;
        RECT 72.370 156.125 72.585 156.175 ;
        RECT 70.790 155.715 71.685 156.090 ;
        RECT 72.195 156.045 72.585 156.125 ;
        RECT 72.760 156.795 73.015 157.365 ;
        RECT 73.185 157.135 73.515 157.535 ;
        RECT 73.940 157.000 74.470 157.365 ;
        RECT 73.940 156.965 74.115 157.000 ;
        RECT 73.185 156.795 74.115 156.965 ;
        RECT 72.760 156.125 72.930 156.795 ;
        RECT 73.185 156.625 73.355 156.795 ;
        RECT 73.100 156.295 73.355 156.625 ;
        RECT 73.580 156.295 73.775 156.625 ;
        RECT 69.735 155.285 70.620 155.455 ;
        RECT 70.800 154.985 71.115 155.485 ;
        RECT 71.345 155.155 71.685 155.715 ;
        RECT 71.855 154.985 72.025 155.995 ;
        RECT 72.195 155.200 72.525 156.045 ;
        RECT 72.760 155.155 73.095 156.125 ;
        RECT 73.265 154.985 73.435 156.125 ;
        RECT 73.605 155.325 73.775 156.295 ;
        RECT 73.945 155.665 74.115 156.795 ;
        RECT 74.285 156.005 74.455 156.805 ;
        RECT 74.660 156.515 74.935 157.365 ;
        RECT 74.655 156.345 74.935 156.515 ;
        RECT 74.660 156.205 74.935 156.345 ;
        RECT 75.105 156.005 75.295 157.365 ;
        RECT 75.475 157.000 75.985 157.535 ;
        RECT 76.205 156.725 76.450 157.330 ;
        RECT 76.895 156.795 77.280 157.365 ;
        RECT 77.450 157.075 77.775 157.535 ;
        RECT 78.295 156.905 78.575 157.365 ;
        RECT 75.495 156.555 76.725 156.725 ;
        RECT 74.285 155.835 75.295 156.005 ;
        RECT 75.465 155.990 76.215 156.180 ;
        RECT 73.945 155.495 75.070 155.665 ;
        RECT 75.465 155.325 75.635 155.990 ;
        RECT 76.385 155.745 76.725 156.555 ;
        RECT 73.605 155.155 75.635 155.325 ;
        RECT 75.805 154.985 75.975 155.745 ;
        RECT 76.210 155.335 76.725 155.745 ;
        RECT 76.895 156.125 77.175 156.795 ;
        RECT 77.450 156.735 78.575 156.905 ;
        RECT 77.450 156.625 77.900 156.735 ;
        RECT 77.345 156.295 77.900 156.625 ;
        RECT 78.765 156.565 79.165 157.365 ;
        RECT 79.565 157.075 79.835 157.535 ;
        RECT 80.005 156.905 80.290 157.365 ;
        RECT 80.575 156.990 85.920 157.535 ;
        RECT 76.895 155.155 77.280 156.125 ;
        RECT 77.450 155.835 77.900 156.295 ;
        RECT 78.070 156.005 79.165 156.565 ;
        RECT 77.450 155.615 78.575 155.835 ;
        RECT 77.450 154.985 77.775 155.445 ;
        RECT 78.295 155.155 78.575 155.615 ;
        RECT 78.765 155.155 79.165 156.005 ;
        RECT 79.335 156.735 80.290 156.905 ;
        RECT 79.335 155.835 79.545 156.735 ;
        RECT 79.715 156.005 80.405 156.565 ;
        RECT 82.160 156.160 82.500 156.990 ;
        RECT 86.095 156.765 89.605 157.535 ;
        RECT 90.695 156.810 90.985 157.535 ;
        RECT 91.155 156.785 92.365 157.535 ;
        RECT 92.625 156.985 92.795 157.275 ;
        RECT 92.965 157.155 93.295 157.535 ;
        RECT 92.625 156.815 93.290 156.985 ;
        RECT 79.335 155.615 80.290 155.835 ;
        RECT 79.565 154.985 79.835 155.445 ;
        RECT 80.005 155.155 80.290 155.615 ;
        RECT 83.980 155.420 84.330 156.670 ;
        RECT 86.095 156.245 87.745 156.765 ;
        RECT 87.915 156.075 89.605 156.595 ;
        RECT 91.155 156.245 91.675 156.785 ;
        RECT 80.575 154.985 85.920 155.420 ;
        RECT 86.095 154.985 89.605 156.075 ;
        RECT 90.695 154.985 90.985 156.150 ;
        RECT 91.845 156.075 92.365 156.615 ;
        RECT 91.155 154.985 92.365 156.075 ;
        RECT 92.540 155.995 92.890 156.645 ;
        RECT 93.060 155.825 93.290 156.815 ;
        RECT 92.625 155.655 93.290 155.825 ;
        RECT 92.625 155.155 92.795 155.655 ;
        RECT 92.965 154.985 93.295 155.485 ;
        RECT 93.465 155.155 93.650 157.275 ;
        RECT 93.905 157.075 94.155 157.535 ;
        RECT 94.325 157.085 94.660 157.255 ;
        RECT 94.855 157.085 95.530 157.255 ;
        RECT 94.325 156.945 94.495 157.085 ;
        RECT 93.820 155.955 94.100 156.905 ;
        RECT 94.270 156.815 94.495 156.945 ;
        RECT 94.270 155.710 94.440 156.815 ;
        RECT 94.665 156.665 95.190 156.885 ;
        RECT 94.610 155.900 94.850 156.495 ;
        RECT 95.020 155.965 95.190 156.665 ;
        RECT 95.360 156.305 95.530 157.085 ;
        RECT 95.850 157.035 96.220 157.535 ;
        RECT 96.400 157.085 96.805 157.255 ;
        RECT 96.975 157.085 97.760 157.255 ;
        RECT 96.400 156.855 96.570 157.085 ;
        RECT 95.740 156.555 96.570 156.855 ;
        RECT 96.955 156.585 97.420 156.915 ;
        RECT 95.740 156.525 95.940 156.555 ;
        RECT 96.060 156.305 96.230 156.375 ;
        RECT 95.360 156.135 96.230 156.305 ;
        RECT 95.720 156.045 96.230 156.135 ;
        RECT 94.270 155.580 94.575 155.710 ;
        RECT 95.020 155.600 95.550 155.965 ;
        RECT 93.890 154.985 94.155 155.445 ;
        RECT 94.325 155.155 94.575 155.580 ;
        RECT 95.720 155.430 95.890 156.045 ;
        RECT 94.785 155.260 95.890 155.430 ;
        RECT 96.060 154.985 96.230 155.785 ;
        RECT 96.400 155.485 96.570 156.555 ;
        RECT 96.740 155.655 96.930 156.375 ;
        RECT 97.100 155.625 97.420 156.585 ;
        RECT 97.590 156.625 97.760 157.085 ;
        RECT 98.035 157.005 98.245 157.535 ;
        RECT 98.505 156.795 98.835 157.320 ;
        RECT 99.005 156.925 99.175 157.535 ;
        RECT 99.345 156.880 99.675 157.315 ;
        RECT 100.865 156.880 101.195 157.315 ;
        RECT 101.365 156.925 101.535 157.535 ;
        RECT 99.345 156.795 99.725 156.880 ;
        RECT 98.635 156.625 98.835 156.795 ;
        RECT 99.500 156.755 99.725 156.795 ;
        RECT 97.590 156.295 98.465 156.625 ;
        RECT 98.635 156.295 99.385 156.625 ;
        RECT 96.400 155.155 96.650 155.485 ;
        RECT 97.590 155.455 97.760 156.295 ;
        RECT 98.635 156.090 98.825 156.295 ;
        RECT 99.555 156.175 99.725 156.755 ;
        RECT 99.510 156.125 99.725 156.175 ;
        RECT 97.930 155.715 98.825 156.090 ;
        RECT 99.335 156.045 99.725 156.125 ;
        RECT 100.815 156.795 101.195 156.880 ;
        RECT 101.705 156.795 102.035 157.320 ;
        RECT 102.295 157.005 102.505 157.535 ;
        RECT 102.780 157.085 103.565 157.255 ;
        RECT 103.735 157.085 104.140 157.255 ;
        RECT 100.815 156.755 101.040 156.795 ;
        RECT 100.815 156.175 100.985 156.755 ;
        RECT 101.705 156.625 101.905 156.795 ;
        RECT 102.780 156.625 102.950 157.085 ;
        RECT 101.155 156.295 101.905 156.625 ;
        RECT 102.075 156.295 102.950 156.625 ;
        RECT 100.815 156.125 101.030 156.175 ;
        RECT 100.815 156.045 101.205 156.125 ;
        RECT 96.875 155.285 97.760 155.455 ;
        RECT 97.940 154.985 98.255 155.485 ;
        RECT 98.485 155.155 98.825 155.715 ;
        RECT 98.995 154.985 99.165 155.995 ;
        RECT 99.335 155.200 99.665 156.045 ;
        RECT 100.875 155.200 101.205 156.045 ;
        RECT 101.715 156.090 101.905 156.295 ;
        RECT 101.375 154.985 101.545 155.995 ;
        RECT 101.715 155.715 102.610 156.090 ;
        RECT 101.715 155.155 102.055 155.715 ;
        RECT 102.285 154.985 102.600 155.485 ;
        RECT 102.780 155.455 102.950 156.295 ;
        RECT 103.120 156.585 103.585 156.915 ;
        RECT 103.970 156.855 104.140 157.085 ;
        RECT 104.320 157.035 104.690 157.535 ;
        RECT 105.010 157.085 105.685 157.255 ;
        RECT 105.880 157.085 106.215 157.255 ;
        RECT 103.120 155.625 103.440 156.585 ;
        RECT 103.970 156.555 104.800 156.855 ;
        RECT 103.610 155.655 103.800 156.375 ;
        RECT 103.970 155.485 104.140 156.555 ;
        RECT 104.600 156.525 104.800 156.555 ;
        RECT 104.310 156.305 104.480 156.375 ;
        RECT 105.010 156.305 105.180 157.085 ;
        RECT 106.045 156.945 106.215 157.085 ;
        RECT 106.385 157.075 106.635 157.535 ;
        RECT 104.310 156.135 105.180 156.305 ;
        RECT 105.350 156.665 105.875 156.885 ;
        RECT 106.045 156.815 106.270 156.945 ;
        RECT 104.310 156.045 104.820 156.135 ;
        RECT 102.780 155.285 103.665 155.455 ;
        RECT 103.890 155.155 104.140 155.485 ;
        RECT 104.310 154.985 104.480 155.785 ;
        RECT 104.650 155.430 104.820 156.045 ;
        RECT 105.350 155.965 105.520 156.665 ;
        RECT 104.990 155.600 105.520 155.965 ;
        RECT 105.690 155.900 105.930 156.495 ;
        RECT 106.100 155.710 106.270 156.815 ;
        RECT 106.440 155.955 106.720 156.905 ;
        RECT 105.965 155.580 106.270 155.710 ;
        RECT 104.650 155.260 105.755 155.430 ;
        RECT 105.965 155.155 106.215 155.580 ;
        RECT 106.385 154.985 106.650 155.445 ;
        RECT 106.890 155.155 107.075 157.275 ;
        RECT 107.245 157.155 107.575 157.535 ;
        RECT 107.745 156.985 107.915 157.275 ;
        RECT 107.250 156.815 107.915 156.985 ;
        RECT 109.145 156.880 109.475 157.315 ;
        RECT 109.645 156.925 109.815 157.535 ;
        RECT 107.250 155.825 107.480 156.815 ;
        RECT 109.095 156.795 109.475 156.880 ;
        RECT 109.985 156.795 110.315 157.320 ;
        RECT 110.575 157.005 110.785 157.535 ;
        RECT 111.060 157.085 111.845 157.255 ;
        RECT 112.015 157.085 112.420 157.255 ;
        RECT 109.095 156.755 109.320 156.795 ;
        RECT 107.650 155.995 108.000 156.645 ;
        RECT 109.095 156.175 109.265 156.755 ;
        RECT 109.985 156.625 110.185 156.795 ;
        RECT 111.060 156.625 111.230 157.085 ;
        RECT 109.435 156.295 110.185 156.625 ;
        RECT 110.355 156.295 111.230 156.625 ;
        RECT 109.095 156.125 109.310 156.175 ;
        RECT 109.095 156.045 109.485 156.125 ;
        RECT 107.250 155.655 107.915 155.825 ;
        RECT 107.245 154.985 107.575 155.485 ;
        RECT 107.745 155.155 107.915 155.655 ;
        RECT 109.155 155.200 109.485 156.045 ;
        RECT 109.995 156.090 110.185 156.295 ;
        RECT 109.655 154.985 109.825 155.995 ;
        RECT 109.995 155.715 110.890 156.090 ;
        RECT 109.995 155.155 110.335 155.715 ;
        RECT 110.565 154.985 110.880 155.485 ;
        RECT 111.060 155.455 111.230 156.295 ;
        RECT 111.400 156.585 111.865 156.915 ;
        RECT 112.250 156.855 112.420 157.085 ;
        RECT 112.600 157.035 112.970 157.535 ;
        RECT 113.290 157.085 113.965 157.255 ;
        RECT 114.160 157.085 114.495 157.255 ;
        RECT 111.400 155.625 111.720 156.585 ;
        RECT 112.250 156.555 113.080 156.855 ;
        RECT 111.890 155.655 112.080 156.375 ;
        RECT 112.250 155.485 112.420 156.555 ;
        RECT 112.880 156.525 113.080 156.555 ;
        RECT 112.590 156.305 112.760 156.375 ;
        RECT 113.290 156.305 113.460 157.085 ;
        RECT 114.325 156.945 114.495 157.085 ;
        RECT 114.665 157.075 114.915 157.535 ;
        RECT 112.590 156.135 113.460 156.305 ;
        RECT 113.630 156.665 114.155 156.885 ;
        RECT 114.325 156.815 114.550 156.945 ;
        RECT 112.590 156.045 113.100 156.135 ;
        RECT 111.060 155.285 111.945 155.455 ;
        RECT 112.170 155.155 112.420 155.485 ;
        RECT 112.590 154.985 112.760 155.785 ;
        RECT 112.930 155.430 113.100 156.045 ;
        RECT 113.630 155.965 113.800 156.665 ;
        RECT 113.270 155.600 113.800 155.965 ;
        RECT 113.970 155.900 114.210 156.495 ;
        RECT 114.380 155.710 114.550 156.815 ;
        RECT 114.720 155.955 115.000 156.905 ;
        RECT 114.245 155.580 114.550 155.710 ;
        RECT 112.930 155.260 114.035 155.430 ;
        RECT 114.245 155.155 114.495 155.580 ;
        RECT 114.665 154.985 114.930 155.445 ;
        RECT 115.170 155.155 115.355 157.275 ;
        RECT 115.525 157.155 115.855 157.535 ;
        RECT 116.025 156.985 116.195 157.275 ;
        RECT 115.530 156.815 116.195 156.985 ;
        RECT 115.530 155.825 115.760 156.815 ;
        RECT 116.455 156.810 116.745 157.535 ;
        RECT 116.915 156.735 117.225 157.535 ;
        RECT 117.430 156.735 118.125 157.365 ;
        RECT 119.220 156.770 119.675 157.535 ;
        RECT 119.950 157.155 121.250 157.365 ;
        RECT 121.505 157.175 121.835 157.535 ;
        RECT 121.080 157.005 121.250 157.155 ;
        RECT 122.005 157.035 122.265 157.365 ;
        RECT 122.035 157.025 122.265 157.035 ;
        RECT 115.930 155.995 116.280 156.645 ;
        RECT 116.925 156.295 117.260 156.565 ;
        RECT 117.430 156.175 117.600 156.735 ;
        RECT 120.150 156.545 120.370 156.945 ;
        RECT 117.770 156.295 118.105 156.545 ;
        RECT 119.215 156.345 119.705 156.545 ;
        RECT 119.895 156.335 120.370 156.545 ;
        RECT 120.615 156.545 120.825 156.945 ;
        RECT 121.080 156.880 121.835 157.005 ;
        RECT 121.080 156.835 121.925 156.880 ;
        RECT 121.655 156.715 121.925 156.835 ;
        RECT 120.615 156.335 120.945 156.545 ;
        RECT 121.115 156.275 121.525 156.580 ;
        RECT 115.530 155.655 116.195 155.825 ;
        RECT 115.525 154.985 115.855 155.485 ;
        RECT 116.025 155.155 116.195 155.655 ;
        RECT 116.455 154.985 116.745 156.150 ;
        RECT 117.430 156.135 117.605 156.175 ;
        RECT 116.915 154.985 117.195 156.125 ;
        RECT 117.365 155.155 117.695 156.135 ;
        RECT 117.865 154.985 118.125 156.125 ;
        RECT 119.220 156.105 120.395 156.165 ;
        RECT 121.755 156.140 121.925 156.715 ;
        RECT 121.725 156.105 121.925 156.140 ;
        RECT 119.220 155.995 121.925 156.105 ;
        RECT 119.220 155.375 119.475 155.995 ;
        RECT 120.065 155.935 121.865 155.995 ;
        RECT 120.065 155.905 120.395 155.935 ;
        RECT 122.095 155.835 122.265 157.025 ;
        RECT 122.440 156.770 122.895 157.535 ;
        RECT 123.170 157.155 124.470 157.365 ;
        RECT 124.725 157.175 125.055 157.535 ;
        RECT 124.300 157.005 124.470 157.155 ;
        RECT 125.225 157.035 125.485 157.365 ;
        RECT 123.370 156.545 123.590 156.945 ;
        RECT 122.435 156.345 122.925 156.545 ;
        RECT 123.115 156.335 123.590 156.545 ;
        RECT 123.835 156.545 124.045 156.945 ;
        RECT 124.300 156.880 125.055 157.005 ;
        RECT 124.300 156.835 125.145 156.880 ;
        RECT 124.875 156.715 125.145 156.835 ;
        RECT 123.835 156.335 124.165 156.545 ;
        RECT 124.335 156.275 124.745 156.580 ;
        RECT 119.725 155.735 119.910 155.825 ;
        RECT 120.500 155.735 121.335 155.745 ;
        RECT 119.725 155.535 121.335 155.735 ;
        RECT 119.725 155.495 119.955 155.535 ;
        RECT 119.220 155.155 119.555 155.375 ;
        RECT 120.560 154.985 120.915 155.365 ;
        RECT 121.085 155.155 121.335 155.535 ;
        RECT 121.585 154.985 121.835 155.765 ;
        RECT 122.005 155.155 122.265 155.835 ;
        RECT 122.440 156.105 123.615 156.165 ;
        RECT 124.975 156.140 125.145 156.715 ;
        RECT 124.945 156.105 125.145 156.140 ;
        RECT 122.440 155.995 125.145 156.105 ;
        RECT 122.440 155.375 122.695 155.995 ;
        RECT 123.285 155.935 125.085 155.995 ;
        RECT 123.285 155.905 123.615 155.935 ;
        RECT 125.315 155.835 125.485 157.035 ;
        RECT 125.660 156.770 126.115 157.535 ;
        RECT 126.390 157.155 127.690 157.365 ;
        RECT 127.945 157.175 128.275 157.535 ;
        RECT 127.520 157.005 127.690 157.155 ;
        RECT 128.445 157.035 128.705 157.365 ;
        RECT 126.590 156.545 126.810 156.945 ;
        RECT 125.655 156.345 126.145 156.545 ;
        RECT 126.335 156.335 126.810 156.545 ;
        RECT 127.055 156.545 127.265 156.945 ;
        RECT 127.520 156.880 128.275 157.005 ;
        RECT 127.520 156.835 128.365 156.880 ;
        RECT 128.095 156.715 128.365 156.835 ;
        RECT 127.055 156.335 127.385 156.545 ;
        RECT 127.555 156.275 127.965 156.580 ;
        RECT 122.945 155.735 123.130 155.825 ;
        RECT 123.720 155.735 124.555 155.745 ;
        RECT 122.945 155.535 124.555 155.735 ;
        RECT 122.945 155.495 123.175 155.535 ;
        RECT 122.440 155.155 122.775 155.375 ;
        RECT 123.780 154.985 124.135 155.365 ;
        RECT 124.305 155.155 124.555 155.535 ;
        RECT 124.805 154.985 125.055 155.765 ;
        RECT 125.225 155.155 125.485 155.835 ;
        RECT 125.660 156.105 126.835 156.165 ;
        RECT 128.195 156.140 128.365 156.715 ;
        RECT 128.165 156.105 128.365 156.140 ;
        RECT 125.660 155.995 128.365 156.105 ;
        RECT 125.660 155.375 125.915 155.995 ;
        RECT 126.505 155.935 128.305 155.995 ;
        RECT 126.505 155.905 126.835 155.935 ;
        RECT 128.535 155.835 128.705 157.035 ;
        RECT 128.875 156.765 130.545 157.535 ;
        RECT 130.805 156.985 130.975 157.365 ;
        RECT 131.155 157.155 131.485 157.535 ;
        RECT 130.805 156.815 131.470 156.985 ;
        RECT 131.665 156.860 131.925 157.365 ;
        RECT 128.875 156.245 129.625 156.765 ;
        RECT 129.795 156.075 130.545 156.595 ;
        RECT 130.735 156.265 131.065 156.635 ;
        RECT 131.300 156.560 131.470 156.815 ;
        RECT 131.300 156.230 131.585 156.560 ;
        RECT 131.300 156.085 131.470 156.230 ;
        RECT 126.165 155.735 126.350 155.825 ;
        RECT 126.940 155.735 127.775 155.745 ;
        RECT 126.165 155.535 127.775 155.735 ;
        RECT 126.165 155.495 126.395 155.535 ;
        RECT 125.660 155.155 125.995 155.375 ;
        RECT 127.000 154.985 127.355 155.365 ;
        RECT 127.525 155.155 127.775 155.535 ;
        RECT 128.025 154.985 128.275 155.765 ;
        RECT 128.445 155.155 128.705 155.835 ;
        RECT 128.875 154.985 130.545 156.075 ;
        RECT 130.805 155.915 131.470 156.085 ;
        RECT 131.755 156.060 131.925 156.860 ;
        RECT 130.805 155.155 130.975 155.915 ;
        RECT 131.155 154.985 131.485 155.745 ;
        RECT 131.655 155.155 131.925 156.060 ;
        RECT 132.095 156.795 132.480 157.365 ;
        RECT 132.650 157.075 132.975 157.535 ;
        RECT 133.495 156.905 133.775 157.365 ;
        RECT 132.095 156.125 132.375 156.795 ;
        RECT 132.650 156.735 133.775 156.905 ;
        RECT 132.650 156.625 133.100 156.735 ;
        RECT 132.545 156.295 133.100 156.625 ;
        RECT 133.965 156.565 134.365 157.365 ;
        RECT 134.765 157.075 135.035 157.535 ;
        RECT 135.205 156.905 135.490 157.365 ;
        RECT 132.095 155.155 132.480 156.125 ;
        RECT 132.650 155.835 133.100 156.295 ;
        RECT 133.270 156.005 134.365 156.565 ;
        RECT 132.650 155.615 133.775 155.835 ;
        RECT 132.650 154.985 132.975 155.445 ;
        RECT 133.495 155.155 133.775 155.615 ;
        RECT 133.965 155.155 134.365 156.005 ;
        RECT 134.535 156.735 135.490 156.905 ;
        RECT 135.865 156.985 136.035 157.365 ;
        RECT 136.250 157.155 136.580 157.535 ;
        RECT 135.865 156.815 136.580 156.985 ;
        RECT 134.535 155.835 134.745 156.735 ;
        RECT 134.915 156.005 135.605 156.565 ;
        RECT 135.775 156.265 136.130 156.635 ;
        RECT 136.410 156.625 136.580 156.815 ;
        RECT 136.750 156.790 137.005 157.365 ;
        RECT 136.410 156.295 136.665 156.625 ;
        RECT 136.410 156.085 136.580 156.295 ;
        RECT 135.865 155.915 136.580 156.085 ;
        RECT 136.835 156.060 137.005 156.790 ;
        RECT 137.180 156.695 137.440 157.535 ;
        RECT 137.615 156.785 138.825 157.535 ;
        RECT 134.535 155.615 135.490 155.835 ;
        RECT 134.765 154.985 135.035 155.445 ;
        RECT 135.205 155.155 135.490 155.615 ;
        RECT 135.865 155.155 136.035 155.915 ;
        RECT 136.250 154.985 136.580 155.745 ;
        RECT 136.750 155.155 137.005 156.060 ;
        RECT 137.180 154.985 137.440 156.135 ;
        RECT 137.615 156.075 138.135 156.615 ;
        RECT 138.305 156.245 138.825 156.785 ;
        RECT 137.615 154.985 138.825 156.075 ;
        RECT 13.330 154.815 138.910 154.985 ;
        RECT 13.415 153.725 14.625 154.815 ;
        RECT 13.415 153.015 13.935 153.555 ;
        RECT 14.105 153.185 14.625 153.725 ;
        RECT 14.795 153.845 15.065 154.615 ;
        RECT 15.235 154.035 15.565 154.815 ;
        RECT 15.770 154.210 15.955 154.615 ;
        RECT 16.125 154.390 16.460 154.815 ;
        RECT 15.770 154.035 16.435 154.210 ;
        RECT 14.795 153.675 15.925 153.845 ;
        RECT 13.415 152.265 14.625 153.015 ;
        RECT 14.795 152.765 14.965 153.675 ;
        RECT 15.135 152.925 15.495 153.505 ;
        RECT 15.675 153.175 15.925 153.675 ;
        RECT 16.095 153.005 16.435 154.035 ;
        RECT 16.635 153.725 18.305 154.815 ;
        RECT 15.750 152.835 16.435 153.005 ;
        RECT 16.635 153.035 17.385 153.555 ;
        RECT 17.555 153.205 18.305 153.725 ;
        RECT 18.485 153.675 18.815 154.815 ;
        RECT 19.345 153.845 19.675 154.630 ;
        RECT 18.995 153.675 19.675 153.845 ;
        RECT 19.855 153.945 20.130 154.645 ;
        RECT 20.300 154.270 20.555 154.815 ;
        RECT 20.725 154.305 21.205 154.645 ;
        RECT 21.380 154.260 21.985 154.815 ;
        RECT 21.370 154.160 21.985 154.260 ;
        RECT 21.370 154.135 21.555 154.160 ;
        RECT 18.475 153.255 18.825 153.505 ;
        RECT 18.995 153.075 19.165 153.675 ;
        RECT 19.335 153.255 19.685 153.505 ;
        RECT 14.795 152.435 15.055 152.765 ;
        RECT 15.265 152.265 15.540 152.745 ;
        RECT 15.750 152.435 15.955 152.835 ;
        RECT 16.125 152.265 16.460 152.665 ;
        RECT 16.635 152.265 18.305 153.035 ;
        RECT 18.485 152.265 18.755 153.075 ;
        RECT 18.925 152.435 19.255 153.075 ;
        RECT 19.425 152.265 19.665 153.075 ;
        RECT 19.855 152.915 20.025 153.945 ;
        RECT 20.300 153.815 21.055 154.065 ;
        RECT 21.225 153.890 21.555 154.135 ;
        RECT 20.300 153.780 21.070 153.815 ;
        RECT 20.300 153.770 21.085 153.780 ;
        RECT 20.195 153.755 21.090 153.770 ;
        RECT 20.195 153.740 21.110 153.755 ;
        RECT 20.195 153.730 21.130 153.740 ;
        RECT 20.195 153.720 21.155 153.730 ;
        RECT 20.195 153.690 21.225 153.720 ;
        RECT 20.195 153.660 21.245 153.690 ;
        RECT 20.195 153.630 21.265 153.660 ;
        RECT 20.195 153.605 21.295 153.630 ;
        RECT 20.195 153.570 21.330 153.605 ;
        RECT 20.195 153.565 21.360 153.570 ;
        RECT 20.195 153.170 20.425 153.565 ;
        RECT 20.970 153.560 21.360 153.565 ;
        RECT 20.995 153.550 21.360 153.560 ;
        RECT 21.010 153.545 21.360 153.550 ;
        RECT 21.025 153.540 21.360 153.545 ;
        RECT 21.725 153.540 21.985 153.990 ;
        RECT 22.165 153.845 22.495 154.630 ;
        RECT 22.165 153.675 22.845 153.845 ;
        RECT 23.025 153.675 23.355 154.815 ;
        RECT 23.570 154.025 24.105 154.645 ;
        RECT 21.025 153.535 21.985 153.540 ;
        RECT 21.035 153.525 21.985 153.535 ;
        RECT 21.045 153.520 21.985 153.525 ;
        RECT 21.055 153.510 21.985 153.520 ;
        RECT 21.060 153.500 21.985 153.510 ;
        RECT 21.065 153.495 21.985 153.500 ;
        RECT 21.075 153.480 21.985 153.495 ;
        RECT 21.080 153.465 21.985 153.480 ;
        RECT 21.090 153.440 21.985 153.465 ;
        RECT 20.595 152.970 20.925 153.395 ;
        RECT 20.675 152.945 20.925 152.970 ;
        RECT 19.855 152.435 20.115 152.915 ;
        RECT 20.285 152.265 20.535 152.805 ;
        RECT 20.705 152.485 20.925 152.945 ;
        RECT 21.095 153.370 21.985 153.440 ;
        RECT 21.095 152.645 21.265 153.370 ;
        RECT 22.155 153.255 22.505 153.505 ;
        RECT 21.435 152.815 21.985 153.200 ;
        RECT 22.675 153.075 22.845 153.675 ;
        RECT 23.015 153.255 23.365 153.505 ;
        RECT 21.095 152.475 21.985 152.645 ;
        RECT 22.175 152.265 22.415 153.075 ;
        RECT 22.585 152.435 22.915 153.075 ;
        RECT 23.085 152.265 23.355 153.075 ;
        RECT 23.570 153.005 23.885 154.025 ;
        RECT 24.275 154.015 24.605 154.815 ;
        RECT 25.090 153.845 25.480 154.020 ;
        RECT 24.055 153.675 25.480 153.845 ;
        RECT 24.055 153.175 24.225 153.675 ;
        RECT 23.570 152.435 24.185 153.005 ;
        RECT 24.475 152.945 24.740 153.505 ;
        RECT 24.910 152.775 25.080 153.675 ;
        RECT 26.295 153.650 26.585 154.815 ;
        RECT 26.755 154.385 27.095 154.645 ;
        RECT 25.250 152.945 25.605 153.505 ;
        RECT 24.355 152.265 24.570 152.775 ;
        RECT 24.800 152.445 25.080 152.775 ;
        RECT 25.260 152.265 25.500 152.775 ;
        RECT 26.295 152.265 26.585 152.990 ;
        RECT 26.755 152.985 27.015 154.385 ;
        RECT 27.265 154.015 27.595 154.815 ;
        RECT 28.060 153.845 28.310 154.645 ;
        RECT 28.495 154.095 28.825 154.815 ;
        RECT 29.045 153.845 29.295 154.645 ;
        RECT 29.465 154.435 29.800 154.815 ;
        RECT 27.205 153.675 29.395 153.845 ;
        RECT 27.205 153.505 27.520 153.675 ;
        RECT 27.190 153.255 27.520 153.505 ;
        RECT 26.755 152.475 27.095 152.985 ;
        RECT 27.265 152.265 27.535 153.065 ;
        RECT 27.715 152.535 27.995 153.505 ;
        RECT 28.175 152.535 28.475 153.505 ;
        RECT 28.655 152.540 29.005 153.505 ;
        RECT 29.225 152.765 29.395 153.675 ;
        RECT 29.565 152.945 29.805 154.255 ;
        RECT 29.975 153.725 33.485 154.815 ;
        RECT 35.075 154.355 35.290 154.815 ;
        RECT 35.460 154.185 35.790 154.645 ;
        RECT 29.975 153.035 31.625 153.555 ;
        RECT 31.795 153.205 33.485 153.725 ;
        RECT 34.620 154.015 35.790 154.185 ;
        RECT 35.960 154.015 36.210 154.815 ;
        RECT 29.225 152.435 29.720 152.765 ;
        RECT 29.975 152.265 33.485 153.035 ;
        RECT 34.620 152.725 34.990 154.015 ;
        RECT 36.420 153.845 36.700 154.005 ;
        RECT 35.365 153.675 36.700 153.845 ;
        RECT 36.875 153.725 39.465 154.815 ;
        RECT 39.640 154.390 39.975 154.815 ;
        RECT 40.145 154.210 40.330 154.615 ;
        RECT 35.365 153.505 35.535 153.675 ;
        RECT 35.160 153.255 35.535 153.505 ;
        RECT 35.705 153.255 36.180 153.495 ;
        RECT 36.350 153.255 36.700 153.495 ;
        RECT 35.365 153.085 35.535 153.255 ;
        RECT 35.365 152.915 36.700 153.085 ;
        RECT 34.620 152.435 35.370 152.725 ;
        RECT 35.880 152.265 36.210 152.725 ;
        RECT 36.430 152.705 36.700 152.915 ;
        RECT 36.875 153.035 38.085 153.555 ;
        RECT 38.255 153.205 39.465 153.725 ;
        RECT 39.665 154.035 40.330 154.210 ;
        RECT 40.535 154.035 40.865 154.815 ;
        RECT 36.875 152.265 39.465 153.035 ;
        RECT 39.665 153.005 40.005 154.035 ;
        RECT 41.035 153.845 41.305 154.615 ;
        RECT 40.175 153.675 41.305 153.845 ;
        RECT 41.565 153.885 41.735 154.645 ;
        RECT 41.950 154.055 42.280 154.815 ;
        RECT 41.565 153.715 42.280 153.885 ;
        RECT 42.450 153.740 42.705 154.645 ;
        RECT 40.175 153.175 40.425 153.675 ;
        RECT 39.665 152.835 40.350 153.005 ;
        RECT 40.605 152.925 40.965 153.505 ;
        RECT 39.640 152.265 39.975 152.665 ;
        RECT 40.145 152.435 40.350 152.835 ;
        RECT 41.135 152.765 41.305 153.675 ;
        RECT 41.475 153.165 41.830 153.535 ;
        RECT 42.110 153.505 42.280 153.715 ;
        RECT 42.110 153.175 42.365 153.505 ;
        RECT 42.110 152.985 42.280 153.175 ;
        RECT 42.535 153.010 42.705 153.740 ;
        RECT 42.880 153.665 43.140 154.815 ;
        RECT 43.315 154.380 48.660 154.815 ;
        RECT 40.560 152.265 40.835 152.745 ;
        RECT 41.045 152.435 41.305 152.765 ;
        RECT 41.565 152.815 42.280 152.985 ;
        RECT 41.565 152.435 41.735 152.815 ;
        RECT 41.950 152.265 42.280 152.645 ;
        RECT 42.450 152.435 42.705 153.010 ;
        RECT 42.880 152.265 43.140 153.105 ;
        RECT 44.900 152.810 45.240 153.640 ;
        RECT 46.720 153.130 47.070 154.380 ;
        RECT 48.835 153.725 51.425 154.815 ;
        RECT 48.835 153.035 50.045 153.555 ;
        RECT 50.215 153.205 51.425 153.725 ;
        RECT 52.055 153.650 52.345 154.815 ;
        RECT 52.515 153.725 54.185 154.815 ;
        RECT 54.360 154.390 54.695 154.815 ;
        RECT 54.865 154.210 55.050 154.615 ;
        RECT 52.515 153.035 53.265 153.555 ;
        RECT 53.435 153.205 54.185 153.725 ;
        RECT 54.385 154.035 55.050 154.210 ;
        RECT 55.255 154.035 55.585 154.815 ;
        RECT 43.315 152.265 48.660 152.810 ;
        RECT 48.835 152.265 51.425 153.035 ;
        RECT 52.055 152.265 52.345 152.990 ;
        RECT 52.515 152.265 54.185 153.035 ;
        RECT 54.385 153.005 54.725 154.035 ;
        RECT 55.755 153.845 56.025 154.615 ;
        RECT 56.200 154.390 56.535 154.815 ;
        RECT 56.705 154.210 56.890 154.615 ;
        RECT 54.895 153.675 56.025 153.845 ;
        RECT 54.895 153.175 55.145 153.675 ;
        RECT 54.385 152.835 55.070 153.005 ;
        RECT 55.325 152.925 55.685 153.505 ;
        RECT 54.360 152.265 54.695 152.665 ;
        RECT 54.865 152.435 55.070 152.835 ;
        RECT 55.855 152.765 56.025 153.675 ;
        RECT 56.225 154.035 56.890 154.210 ;
        RECT 57.095 154.035 57.425 154.815 ;
        RECT 56.225 153.005 56.565 154.035 ;
        RECT 57.595 153.845 57.865 154.615 ;
        RECT 56.735 153.675 57.865 153.845 ;
        RECT 58.035 153.675 58.315 154.815 ;
        RECT 56.735 153.175 56.985 153.675 ;
        RECT 56.225 152.835 56.910 153.005 ;
        RECT 57.165 152.925 57.525 153.505 ;
        RECT 55.280 152.265 55.555 152.745 ;
        RECT 55.765 152.435 56.025 152.765 ;
        RECT 56.200 152.265 56.535 152.665 ;
        RECT 56.705 152.435 56.910 152.835 ;
        RECT 57.695 152.765 57.865 153.675 ;
        RECT 58.485 153.665 58.815 154.645 ;
        RECT 58.985 153.675 59.245 154.815 ;
        RECT 59.415 153.725 62.005 154.815 ;
        RECT 62.695 153.755 63.025 154.600 ;
        RECT 63.195 153.805 63.365 154.815 ;
        RECT 63.535 154.085 63.875 154.645 ;
        RECT 64.105 154.315 64.420 154.815 ;
        RECT 64.600 154.345 65.485 154.515 ;
        RECT 58.045 153.235 58.380 153.505 ;
        RECT 58.550 153.065 58.720 153.665 ;
        RECT 58.890 153.255 59.225 153.505 ;
        RECT 57.120 152.265 57.395 152.745 ;
        RECT 57.605 152.435 57.865 152.765 ;
        RECT 58.035 152.265 58.345 153.065 ;
        RECT 58.550 152.435 59.245 153.065 ;
        RECT 59.415 153.035 60.625 153.555 ;
        RECT 60.795 153.205 62.005 153.725 ;
        RECT 62.635 153.675 63.025 153.755 ;
        RECT 63.535 153.710 64.430 154.085 ;
        RECT 62.635 153.625 62.850 153.675 ;
        RECT 62.635 153.045 62.805 153.625 ;
        RECT 63.535 153.505 63.725 153.710 ;
        RECT 64.600 153.505 64.770 154.345 ;
        RECT 65.710 154.315 65.960 154.645 ;
        RECT 62.975 153.175 63.725 153.505 ;
        RECT 63.895 153.175 64.770 153.505 ;
        RECT 59.415 152.265 62.005 153.035 ;
        RECT 62.635 153.005 62.860 153.045 ;
        RECT 63.525 153.005 63.725 153.175 ;
        RECT 62.635 152.920 63.015 153.005 ;
        RECT 62.685 152.485 63.015 152.920 ;
        RECT 63.185 152.265 63.355 152.875 ;
        RECT 63.525 152.480 63.855 153.005 ;
        RECT 64.115 152.265 64.325 152.795 ;
        RECT 64.600 152.715 64.770 153.175 ;
        RECT 64.940 153.215 65.260 154.175 ;
        RECT 65.430 153.425 65.620 154.145 ;
        RECT 65.790 153.245 65.960 154.315 ;
        RECT 66.130 154.015 66.300 154.815 ;
        RECT 66.470 154.370 67.575 154.540 ;
        RECT 66.470 153.755 66.640 154.370 ;
        RECT 67.785 154.220 68.035 154.645 ;
        RECT 68.205 154.355 68.470 154.815 ;
        RECT 66.810 153.835 67.340 154.200 ;
        RECT 67.785 154.090 68.090 154.220 ;
        RECT 66.130 153.665 66.640 153.755 ;
        RECT 66.130 153.495 67.000 153.665 ;
        RECT 66.130 153.425 66.300 153.495 ;
        RECT 66.420 153.245 66.620 153.275 ;
        RECT 64.940 152.885 65.405 153.215 ;
        RECT 65.790 152.945 66.620 153.245 ;
        RECT 65.790 152.715 65.960 152.945 ;
        RECT 64.600 152.545 65.385 152.715 ;
        RECT 65.555 152.545 65.960 152.715 ;
        RECT 66.140 152.265 66.510 152.765 ;
        RECT 66.830 152.715 67.000 153.495 ;
        RECT 67.170 153.135 67.340 153.835 ;
        RECT 67.510 153.305 67.750 153.900 ;
        RECT 67.170 152.915 67.695 153.135 ;
        RECT 67.920 152.985 68.090 154.090 ;
        RECT 67.865 152.855 68.090 152.985 ;
        RECT 68.260 152.895 68.540 153.845 ;
        RECT 67.865 152.715 68.035 152.855 ;
        RECT 66.830 152.545 67.505 152.715 ;
        RECT 67.700 152.545 68.035 152.715 ;
        RECT 68.205 152.265 68.455 152.725 ;
        RECT 68.710 152.525 68.895 154.645 ;
        RECT 69.065 154.315 69.395 154.815 ;
        RECT 69.565 154.145 69.735 154.645 ;
        RECT 69.070 153.975 69.735 154.145 ;
        RECT 69.070 152.985 69.300 153.975 ;
        RECT 69.470 153.155 69.820 153.805 ;
        RECT 70.000 153.675 70.335 154.645 ;
        RECT 70.505 153.675 70.675 154.815 ;
        RECT 70.845 154.475 72.875 154.645 ;
        RECT 70.000 153.005 70.170 153.675 ;
        RECT 70.845 153.505 71.015 154.475 ;
        RECT 70.340 153.175 70.595 153.505 ;
        RECT 70.820 153.175 71.015 153.505 ;
        RECT 71.185 154.135 72.310 154.305 ;
        RECT 70.425 153.005 70.595 153.175 ;
        RECT 71.185 153.005 71.355 154.135 ;
        RECT 69.070 152.815 69.735 152.985 ;
        RECT 69.065 152.265 69.395 152.645 ;
        RECT 69.565 152.525 69.735 152.815 ;
        RECT 70.000 152.435 70.255 153.005 ;
        RECT 70.425 152.835 71.355 153.005 ;
        RECT 71.525 153.795 72.535 153.965 ;
        RECT 71.525 152.995 71.695 153.795 ;
        RECT 71.900 153.115 72.175 153.595 ;
        RECT 71.895 152.945 72.175 153.115 ;
        RECT 71.180 152.800 71.355 152.835 ;
        RECT 70.425 152.265 70.755 152.665 ;
        RECT 71.180 152.435 71.710 152.800 ;
        RECT 71.900 152.435 72.175 152.945 ;
        RECT 72.345 152.435 72.535 153.795 ;
        RECT 72.705 153.810 72.875 154.475 ;
        RECT 73.045 154.055 73.215 154.815 ;
        RECT 73.450 154.055 73.965 154.465 ;
        RECT 72.705 153.620 73.455 153.810 ;
        RECT 73.625 153.245 73.965 154.055 ;
        RECT 74.190 153.945 74.475 154.815 ;
        RECT 74.645 154.185 74.905 154.645 ;
        RECT 75.080 154.355 75.335 154.815 ;
        RECT 75.505 154.185 75.765 154.645 ;
        RECT 74.645 154.015 75.765 154.185 ;
        RECT 75.935 154.015 76.245 154.815 ;
        RECT 74.645 153.765 74.905 154.015 ;
        RECT 76.415 153.845 76.725 154.645 ;
        RECT 72.735 153.075 73.965 153.245 ;
        RECT 74.150 153.595 74.905 153.765 ;
        RECT 75.695 153.675 76.725 153.845 ;
        RECT 74.150 153.085 74.555 153.595 ;
        RECT 75.695 153.425 75.865 153.675 ;
        RECT 74.725 153.255 75.865 153.425 ;
        RECT 72.715 152.265 73.225 152.800 ;
        RECT 73.445 152.470 73.690 153.075 ;
        RECT 74.150 152.915 75.800 153.085 ;
        RECT 76.035 152.935 76.385 153.505 ;
        RECT 74.195 152.265 74.475 152.745 ;
        RECT 74.645 152.525 74.905 152.915 ;
        RECT 75.080 152.265 75.335 152.745 ;
        RECT 75.505 152.525 75.800 152.915 ;
        RECT 76.555 152.765 76.725 153.675 ;
        RECT 77.815 153.650 78.105 154.815 ;
        RECT 78.275 153.725 79.945 154.815 ;
        RECT 78.275 153.035 79.025 153.555 ;
        RECT 79.195 153.205 79.945 153.725 ;
        RECT 80.120 153.675 80.455 154.645 ;
        RECT 80.625 153.675 80.795 154.815 ;
        RECT 80.965 154.475 82.995 154.645 ;
        RECT 75.980 152.265 76.255 152.745 ;
        RECT 76.425 152.435 76.725 152.765 ;
        RECT 77.815 152.265 78.105 152.990 ;
        RECT 78.275 152.265 79.945 153.035 ;
        RECT 80.120 153.005 80.290 153.675 ;
        RECT 80.965 153.505 81.135 154.475 ;
        RECT 80.460 153.175 80.715 153.505 ;
        RECT 80.940 153.175 81.135 153.505 ;
        RECT 81.305 154.135 82.430 154.305 ;
        RECT 80.545 153.005 80.715 153.175 ;
        RECT 81.305 153.005 81.475 154.135 ;
        RECT 80.120 152.435 80.375 153.005 ;
        RECT 80.545 152.835 81.475 153.005 ;
        RECT 81.645 153.795 82.655 153.965 ;
        RECT 81.645 152.995 81.815 153.795 ;
        RECT 81.300 152.800 81.475 152.835 ;
        RECT 80.545 152.265 80.875 152.665 ;
        RECT 81.300 152.435 81.830 152.800 ;
        RECT 82.020 152.775 82.295 153.595 ;
        RECT 82.015 152.605 82.295 152.775 ;
        RECT 82.020 152.435 82.295 152.605 ;
        RECT 82.465 152.435 82.655 153.795 ;
        RECT 82.825 153.810 82.995 154.475 ;
        RECT 83.165 154.055 83.335 154.815 ;
        RECT 83.570 154.055 84.085 154.465 ;
        RECT 82.825 153.620 83.575 153.810 ;
        RECT 83.745 153.245 84.085 154.055 ;
        RECT 84.370 154.185 84.655 154.645 ;
        RECT 84.825 154.355 85.095 154.815 ;
        RECT 84.370 153.965 85.325 154.185 ;
        RECT 82.855 153.075 84.085 153.245 ;
        RECT 84.255 153.235 84.945 153.795 ;
        RECT 82.835 152.265 83.345 152.800 ;
        RECT 83.565 152.470 83.810 153.075 ;
        RECT 85.115 153.065 85.325 153.965 ;
        RECT 84.370 152.895 85.325 153.065 ;
        RECT 85.495 153.795 85.895 154.645 ;
        RECT 86.085 154.185 86.365 154.645 ;
        RECT 86.885 154.355 87.210 154.815 ;
        RECT 86.085 153.965 87.210 154.185 ;
        RECT 85.495 153.235 86.590 153.795 ;
        RECT 86.760 153.505 87.210 153.965 ;
        RECT 87.380 153.675 87.765 154.645 ;
        RECT 87.935 154.380 93.280 154.815 ;
        RECT 84.370 152.435 84.655 152.895 ;
        RECT 84.825 152.265 85.095 152.725 ;
        RECT 85.495 152.435 85.895 153.235 ;
        RECT 86.760 153.175 87.315 153.505 ;
        RECT 86.760 153.065 87.210 153.175 ;
        RECT 86.085 152.895 87.210 153.065 ;
        RECT 87.485 153.005 87.765 153.675 ;
        RECT 86.085 152.435 86.365 152.895 ;
        RECT 86.885 152.265 87.210 152.725 ;
        RECT 87.380 152.435 87.765 153.005 ;
        RECT 89.520 152.810 89.860 153.640 ;
        RECT 91.340 153.130 91.690 154.380 ;
        RECT 93.455 153.725 94.665 154.815 ;
        RECT 93.455 153.015 93.975 153.555 ;
        RECT 94.145 153.185 94.665 153.725 ;
        RECT 94.840 153.675 95.175 154.645 ;
        RECT 95.345 153.675 95.515 154.815 ;
        RECT 95.685 154.475 97.715 154.645 ;
        RECT 87.935 152.265 93.280 152.810 ;
        RECT 93.455 152.265 94.665 153.015 ;
        RECT 94.840 153.005 95.010 153.675 ;
        RECT 95.685 153.505 95.855 154.475 ;
        RECT 95.180 153.175 95.435 153.505 ;
        RECT 95.660 153.175 95.855 153.505 ;
        RECT 96.025 154.135 97.150 154.305 ;
        RECT 95.265 153.005 95.435 153.175 ;
        RECT 96.025 153.005 96.195 154.135 ;
        RECT 94.840 152.435 95.095 153.005 ;
        RECT 95.265 152.835 96.195 153.005 ;
        RECT 96.365 153.795 97.375 153.965 ;
        RECT 96.365 152.995 96.535 153.795 ;
        RECT 96.740 153.115 97.015 153.595 ;
        RECT 96.735 152.945 97.015 153.115 ;
        RECT 96.020 152.800 96.195 152.835 ;
        RECT 95.265 152.265 95.595 152.665 ;
        RECT 96.020 152.435 96.550 152.800 ;
        RECT 96.740 152.435 97.015 152.945 ;
        RECT 97.185 152.435 97.375 153.795 ;
        RECT 97.545 153.810 97.715 154.475 ;
        RECT 97.885 154.055 98.055 154.815 ;
        RECT 98.290 154.055 98.805 154.465 ;
        RECT 97.545 153.620 98.295 153.810 ;
        RECT 98.465 153.245 98.805 154.055 ;
        RECT 97.575 153.075 98.805 153.245 ;
        RECT 98.980 153.675 99.315 154.645 ;
        RECT 99.485 153.675 99.655 154.815 ;
        RECT 99.825 154.475 101.855 154.645 ;
        RECT 97.555 152.265 98.065 152.800 ;
        RECT 98.285 152.470 98.530 153.075 ;
        RECT 98.980 153.005 99.150 153.675 ;
        RECT 99.825 153.505 99.995 154.475 ;
        RECT 99.320 153.175 99.575 153.505 ;
        RECT 99.800 153.175 99.995 153.505 ;
        RECT 100.165 154.135 101.290 154.305 ;
        RECT 99.405 153.005 99.575 153.175 ;
        RECT 100.165 153.005 100.335 154.135 ;
        RECT 98.980 152.435 99.235 153.005 ;
        RECT 99.405 152.835 100.335 153.005 ;
        RECT 100.505 153.795 101.515 153.965 ;
        RECT 100.505 152.995 100.675 153.795 ;
        RECT 100.160 152.800 100.335 152.835 ;
        RECT 99.405 152.265 99.735 152.665 ;
        RECT 100.160 152.435 100.690 152.800 ;
        RECT 100.880 152.775 101.155 153.595 ;
        RECT 100.875 152.605 101.155 152.775 ;
        RECT 100.880 152.435 101.155 152.605 ;
        RECT 101.325 152.435 101.515 153.795 ;
        RECT 101.685 153.810 101.855 154.475 ;
        RECT 102.025 154.055 102.195 154.815 ;
        RECT 102.430 154.055 102.945 154.465 ;
        RECT 101.685 153.620 102.435 153.810 ;
        RECT 102.605 153.245 102.945 154.055 ;
        RECT 103.575 153.650 103.865 154.815 ;
        RECT 104.610 154.185 104.895 154.645 ;
        RECT 105.065 154.355 105.335 154.815 ;
        RECT 104.610 153.965 105.565 154.185 ;
        RECT 101.715 153.075 102.945 153.245 ;
        RECT 104.495 153.235 105.185 153.795 ;
        RECT 101.695 152.265 102.205 152.800 ;
        RECT 102.425 152.470 102.670 153.075 ;
        RECT 105.355 153.065 105.565 153.965 ;
        RECT 103.575 152.265 103.865 152.990 ;
        RECT 104.610 152.895 105.565 153.065 ;
        RECT 105.735 153.795 106.135 154.645 ;
        RECT 106.325 154.185 106.605 154.645 ;
        RECT 107.125 154.355 107.450 154.815 ;
        RECT 106.325 153.965 107.450 154.185 ;
        RECT 105.735 153.235 106.830 153.795 ;
        RECT 107.000 153.505 107.450 153.965 ;
        RECT 107.620 153.675 108.005 154.645 ;
        RECT 108.215 153.675 108.445 154.815 ;
        RECT 104.610 152.435 104.895 152.895 ;
        RECT 105.065 152.265 105.335 152.725 ;
        RECT 105.735 152.435 106.135 153.235 ;
        RECT 107.000 153.175 107.555 153.505 ;
        RECT 107.000 153.065 107.450 153.175 ;
        RECT 106.325 152.895 107.450 153.065 ;
        RECT 107.725 153.005 108.005 153.675 ;
        RECT 108.615 153.665 108.945 154.645 ;
        RECT 109.115 153.675 109.325 154.815 ;
        RECT 110.475 153.675 110.735 154.815 ;
        RECT 110.905 153.665 111.235 154.645 ;
        RECT 111.405 153.675 111.685 154.815 ;
        RECT 111.855 153.725 115.365 154.815 ;
        RECT 108.195 153.255 108.525 153.505 ;
        RECT 106.325 152.435 106.605 152.895 ;
        RECT 107.125 152.265 107.450 152.725 ;
        RECT 107.620 152.435 108.005 153.005 ;
        RECT 108.215 152.265 108.445 153.085 ;
        RECT 108.695 153.065 108.945 153.665 ;
        RECT 110.495 153.255 110.830 153.505 ;
        RECT 108.615 152.435 108.945 153.065 ;
        RECT 109.115 152.265 109.325 153.085 ;
        RECT 111.000 153.065 111.170 153.665 ;
        RECT 111.340 153.235 111.675 153.505 ;
        RECT 110.475 152.435 111.170 153.065 ;
        RECT 111.375 152.265 111.685 153.065 ;
        RECT 111.855 153.035 113.505 153.555 ;
        RECT 113.675 153.205 115.365 153.725 ;
        RECT 115.535 154.055 116.050 154.465 ;
        RECT 116.285 154.055 116.455 154.815 ;
        RECT 116.625 154.475 118.655 154.645 ;
        RECT 115.535 153.245 115.875 154.055 ;
        RECT 116.625 153.810 116.795 154.475 ;
        RECT 117.190 154.135 118.315 154.305 ;
        RECT 116.045 153.620 116.795 153.810 ;
        RECT 116.965 153.795 117.975 153.965 ;
        RECT 115.535 153.075 116.765 153.245 ;
        RECT 111.855 152.265 115.365 153.035 ;
        RECT 115.810 152.470 116.055 153.075 ;
        RECT 116.275 152.265 116.785 152.800 ;
        RECT 116.965 152.435 117.155 153.795 ;
        RECT 117.325 153.455 117.600 153.595 ;
        RECT 117.325 153.285 117.605 153.455 ;
        RECT 117.325 152.435 117.600 153.285 ;
        RECT 117.805 152.995 117.975 153.795 ;
        RECT 118.145 153.005 118.315 154.135 ;
        RECT 118.485 153.505 118.655 154.475 ;
        RECT 118.825 153.675 118.995 154.815 ;
        RECT 119.165 153.675 119.500 154.645 ;
        RECT 118.485 153.175 118.680 153.505 ;
        RECT 118.905 153.175 119.160 153.505 ;
        RECT 118.905 153.005 119.075 153.175 ;
        RECT 119.330 153.005 119.500 153.675 ;
        RECT 119.680 153.665 119.940 154.815 ;
        RECT 120.115 153.740 120.370 154.645 ;
        RECT 120.540 154.055 120.870 154.815 ;
        RECT 121.085 153.885 121.255 154.645 ;
        RECT 122.065 154.145 122.235 154.645 ;
        RECT 122.405 154.315 122.735 154.815 ;
        RECT 122.065 153.975 122.730 154.145 ;
        RECT 118.145 152.835 119.075 153.005 ;
        RECT 118.145 152.800 118.320 152.835 ;
        RECT 117.790 152.435 118.320 152.800 ;
        RECT 118.745 152.265 119.075 152.665 ;
        RECT 119.245 152.435 119.500 153.005 ;
        RECT 119.680 152.265 119.940 153.105 ;
        RECT 120.115 153.010 120.285 153.740 ;
        RECT 120.540 153.715 121.255 153.885 ;
        RECT 120.540 153.505 120.710 153.715 ;
        RECT 120.455 153.175 120.710 153.505 ;
        RECT 120.115 152.435 120.370 153.010 ;
        RECT 120.540 152.985 120.710 153.175 ;
        RECT 120.990 153.165 121.345 153.535 ;
        RECT 121.980 153.155 122.330 153.805 ;
        RECT 122.500 152.985 122.730 153.975 ;
        RECT 120.540 152.815 121.255 152.985 ;
        RECT 120.540 152.265 120.870 152.645 ;
        RECT 121.085 152.435 121.255 152.815 ;
        RECT 122.065 152.815 122.730 152.985 ;
        RECT 122.065 152.525 122.235 152.815 ;
        RECT 122.405 152.265 122.735 152.645 ;
        RECT 122.905 152.525 123.090 154.645 ;
        RECT 123.330 154.355 123.595 154.815 ;
        RECT 123.765 154.220 124.015 154.645 ;
        RECT 124.225 154.370 125.330 154.540 ;
        RECT 123.710 154.090 124.015 154.220 ;
        RECT 123.260 152.895 123.540 153.845 ;
        RECT 123.710 152.985 123.880 154.090 ;
        RECT 124.050 153.305 124.290 153.900 ;
        RECT 124.460 153.835 124.990 154.200 ;
        RECT 124.460 153.135 124.630 153.835 ;
        RECT 125.160 153.755 125.330 154.370 ;
        RECT 125.500 154.015 125.670 154.815 ;
        RECT 125.840 154.315 126.090 154.645 ;
        RECT 126.315 154.345 127.200 154.515 ;
        RECT 125.160 153.665 125.670 153.755 ;
        RECT 123.710 152.855 123.935 152.985 ;
        RECT 124.105 152.915 124.630 153.135 ;
        RECT 124.800 153.495 125.670 153.665 ;
        RECT 123.345 152.265 123.595 152.725 ;
        RECT 123.765 152.715 123.935 152.855 ;
        RECT 124.800 152.715 124.970 153.495 ;
        RECT 125.500 153.425 125.670 153.495 ;
        RECT 125.180 153.245 125.380 153.275 ;
        RECT 125.840 153.245 126.010 154.315 ;
        RECT 126.180 153.425 126.370 154.145 ;
        RECT 125.180 152.945 126.010 153.245 ;
        RECT 126.540 153.215 126.860 154.175 ;
        RECT 123.765 152.545 124.100 152.715 ;
        RECT 124.295 152.545 124.970 152.715 ;
        RECT 125.290 152.265 125.660 152.765 ;
        RECT 125.840 152.715 126.010 152.945 ;
        RECT 126.395 152.885 126.860 153.215 ;
        RECT 127.030 153.505 127.200 154.345 ;
        RECT 127.380 154.315 127.695 154.815 ;
        RECT 127.925 154.085 128.265 154.645 ;
        RECT 127.370 153.710 128.265 154.085 ;
        RECT 128.435 153.805 128.605 154.815 ;
        RECT 128.075 153.505 128.265 153.710 ;
        RECT 128.775 153.755 129.105 154.600 ;
        RECT 128.775 153.675 129.165 153.755 ;
        RECT 128.950 153.625 129.165 153.675 ;
        RECT 129.335 153.650 129.625 154.815 ;
        RECT 129.795 153.675 130.180 154.645 ;
        RECT 130.350 154.355 130.675 154.815 ;
        RECT 131.195 154.185 131.475 154.645 ;
        RECT 130.350 153.965 131.475 154.185 ;
        RECT 127.030 153.175 127.905 153.505 ;
        RECT 128.075 153.175 128.825 153.505 ;
        RECT 127.030 152.715 127.200 153.175 ;
        RECT 128.075 153.005 128.275 153.175 ;
        RECT 128.995 153.045 129.165 153.625 ;
        RECT 128.940 153.005 129.165 153.045 ;
        RECT 125.840 152.545 126.245 152.715 ;
        RECT 126.415 152.545 127.200 152.715 ;
        RECT 127.475 152.265 127.685 152.795 ;
        RECT 127.945 152.480 128.275 153.005 ;
        RECT 128.785 152.920 129.165 153.005 ;
        RECT 129.795 153.005 130.075 153.675 ;
        RECT 130.350 153.505 130.800 153.965 ;
        RECT 131.665 153.795 132.065 154.645 ;
        RECT 132.465 154.355 132.735 154.815 ;
        RECT 132.905 154.185 133.190 154.645 ;
        RECT 130.245 153.175 130.800 153.505 ;
        RECT 130.970 153.235 132.065 153.795 ;
        RECT 130.350 153.065 130.800 153.175 ;
        RECT 128.445 152.265 128.615 152.875 ;
        RECT 128.785 152.485 129.115 152.920 ;
        RECT 129.335 152.265 129.625 152.990 ;
        RECT 129.795 152.435 130.180 153.005 ;
        RECT 130.350 152.895 131.475 153.065 ;
        RECT 130.350 152.265 130.675 152.725 ;
        RECT 131.195 152.435 131.475 152.895 ;
        RECT 131.665 152.435 132.065 153.235 ;
        RECT 132.235 153.965 133.190 154.185 ;
        RECT 132.235 153.065 132.445 153.965 ;
        RECT 134.025 153.885 134.195 154.645 ;
        RECT 134.410 154.055 134.740 154.815 ;
        RECT 132.615 153.235 133.305 153.795 ;
        RECT 134.025 153.715 134.740 153.885 ;
        RECT 134.910 153.740 135.165 154.645 ;
        RECT 133.935 153.165 134.290 153.535 ;
        RECT 134.570 153.505 134.740 153.715 ;
        RECT 134.570 153.175 134.825 153.505 ;
        RECT 132.235 152.895 133.190 153.065 ;
        RECT 134.570 152.985 134.740 153.175 ;
        RECT 134.995 153.010 135.165 153.740 ;
        RECT 135.340 153.665 135.600 154.815 ;
        RECT 135.865 153.885 136.035 154.645 ;
        RECT 136.250 154.055 136.580 154.815 ;
        RECT 135.865 153.715 136.580 153.885 ;
        RECT 136.750 153.740 137.005 154.645 ;
        RECT 135.775 153.165 136.130 153.535 ;
        RECT 136.410 153.505 136.580 153.715 ;
        RECT 136.410 153.175 136.665 153.505 ;
        RECT 132.465 152.265 132.735 152.725 ;
        RECT 132.905 152.435 133.190 152.895 ;
        RECT 134.025 152.815 134.740 152.985 ;
        RECT 134.025 152.435 134.195 152.815 ;
        RECT 134.410 152.265 134.740 152.645 ;
        RECT 134.910 152.435 135.165 153.010 ;
        RECT 135.340 152.265 135.600 153.105 ;
        RECT 136.410 152.985 136.580 153.175 ;
        RECT 136.835 153.010 137.005 153.740 ;
        RECT 137.180 153.665 137.440 154.815 ;
        RECT 137.615 153.725 138.825 154.815 ;
        RECT 137.615 153.185 138.135 153.725 ;
        RECT 135.865 152.815 136.580 152.985 ;
        RECT 135.865 152.435 136.035 152.815 ;
        RECT 136.250 152.265 136.580 152.645 ;
        RECT 136.750 152.435 137.005 153.010 ;
        RECT 137.180 152.265 137.440 153.105 ;
        RECT 138.305 153.015 138.825 153.555 ;
        RECT 137.615 152.265 138.825 153.015 ;
        RECT 13.330 152.095 138.910 152.265 ;
        RECT 13.415 151.345 14.625 152.095 ;
        RECT 13.415 150.805 13.935 151.345 ;
        RECT 14.795 151.325 16.465 152.095 ;
        RECT 16.635 151.445 16.895 151.925 ;
        RECT 17.065 151.635 17.395 152.095 ;
        RECT 17.585 151.455 17.785 151.875 ;
        RECT 14.105 150.635 14.625 151.175 ;
        RECT 14.795 150.805 15.545 151.325 ;
        RECT 15.715 150.635 16.465 151.155 ;
        RECT 13.415 149.545 14.625 150.635 ;
        RECT 14.795 149.545 16.465 150.635 ;
        RECT 16.635 150.415 16.805 151.445 ;
        RECT 16.975 150.755 17.205 151.185 ;
        RECT 17.375 150.935 17.785 151.455 ;
        RECT 17.955 151.610 18.745 151.875 ;
        RECT 17.955 150.755 18.210 151.610 ;
        RECT 18.925 151.275 19.255 151.695 ;
        RECT 19.425 151.275 19.685 152.095 ;
        RECT 19.940 151.595 20.435 151.925 ;
        RECT 18.925 151.185 19.175 151.275 ;
        RECT 18.380 150.935 19.175 151.185 ;
        RECT 16.975 150.585 18.765 150.755 ;
        RECT 16.635 149.715 16.910 150.415 ;
        RECT 17.080 150.290 17.795 150.585 ;
        RECT 18.015 150.225 18.345 150.415 ;
        RECT 17.120 149.545 17.335 150.090 ;
        RECT 17.505 149.715 17.980 150.055 ;
        RECT 18.150 150.050 18.345 150.225 ;
        RECT 18.515 150.220 18.765 150.585 ;
        RECT 18.150 149.545 18.765 150.050 ;
        RECT 19.005 149.715 19.175 150.935 ;
        RECT 19.345 150.225 19.685 151.105 ;
        RECT 19.855 150.105 20.095 151.415 ;
        RECT 20.265 150.685 20.435 151.595 ;
        RECT 20.655 150.855 21.005 151.820 ;
        RECT 21.185 150.855 21.485 151.825 ;
        RECT 21.665 150.855 21.945 151.825 ;
        RECT 22.125 151.295 22.395 152.095 ;
        RECT 22.565 151.375 22.905 151.885 ;
        RECT 23.165 151.545 23.335 151.835 ;
        RECT 23.505 151.715 23.835 152.095 ;
        RECT 23.165 151.375 23.830 151.545 ;
        RECT 22.140 150.855 22.470 151.105 ;
        RECT 22.140 150.685 22.455 150.855 ;
        RECT 20.265 150.515 22.455 150.685 ;
        RECT 19.425 149.545 19.685 150.055 ;
        RECT 19.860 149.545 20.195 149.925 ;
        RECT 20.365 149.715 20.615 150.515 ;
        RECT 20.835 149.545 21.165 150.265 ;
        RECT 21.350 149.715 21.600 150.515 ;
        RECT 22.065 149.545 22.395 150.345 ;
        RECT 22.645 149.975 22.905 151.375 ;
        RECT 23.080 150.555 23.430 151.205 ;
        RECT 23.600 150.385 23.830 151.375 ;
        RECT 22.565 149.715 22.905 149.975 ;
        RECT 23.165 150.215 23.830 150.385 ;
        RECT 23.165 149.715 23.335 150.215 ;
        RECT 23.505 149.545 23.835 150.045 ;
        RECT 24.005 149.715 24.190 151.835 ;
        RECT 24.445 151.635 24.695 152.095 ;
        RECT 24.865 151.645 25.200 151.815 ;
        RECT 25.395 151.645 26.070 151.815 ;
        RECT 24.865 151.505 25.035 151.645 ;
        RECT 24.360 150.515 24.640 151.465 ;
        RECT 24.810 151.375 25.035 151.505 ;
        RECT 24.810 150.270 24.980 151.375 ;
        RECT 25.205 151.225 25.730 151.445 ;
        RECT 25.150 150.460 25.390 151.055 ;
        RECT 25.560 150.525 25.730 151.225 ;
        RECT 25.900 150.865 26.070 151.645 ;
        RECT 26.390 151.595 26.760 152.095 ;
        RECT 26.940 151.645 27.345 151.815 ;
        RECT 27.515 151.645 28.300 151.815 ;
        RECT 26.940 151.415 27.110 151.645 ;
        RECT 26.280 151.115 27.110 151.415 ;
        RECT 27.495 151.145 27.960 151.475 ;
        RECT 26.280 151.085 26.480 151.115 ;
        RECT 26.600 150.865 26.770 150.935 ;
        RECT 25.900 150.695 26.770 150.865 ;
        RECT 26.260 150.605 26.770 150.695 ;
        RECT 24.810 150.140 25.115 150.270 ;
        RECT 25.560 150.160 26.090 150.525 ;
        RECT 24.430 149.545 24.695 150.005 ;
        RECT 24.865 149.715 25.115 150.140 ;
        RECT 26.260 149.990 26.430 150.605 ;
        RECT 25.325 149.820 26.430 149.990 ;
        RECT 26.600 149.545 26.770 150.345 ;
        RECT 26.940 150.045 27.110 151.115 ;
        RECT 27.280 150.215 27.470 150.935 ;
        RECT 27.640 150.185 27.960 151.145 ;
        RECT 28.130 151.185 28.300 151.645 ;
        RECT 28.575 151.565 28.785 152.095 ;
        RECT 29.045 151.355 29.375 151.880 ;
        RECT 29.545 151.485 29.715 152.095 ;
        RECT 29.885 151.440 30.215 151.875 ;
        RECT 29.885 151.355 30.265 151.440 ;
        RECT 29.175 151.185 29.375 151.355 ;
        RECT 30.040 151.315 30.265 151.355 ;
        RECT 28.130 150.855 29.005 151.185 ;
        RECT 29.175 150.855 29.925 151.185 ;
        RECT 26.940 149.715 27.190 150.045 ;
        RECT 28.130 150.015 28.300 150.855 ;
        RECT 29.175 150.650 29.365 150.855 ;
        RECT 30.095 150.735 30.265 151.315 ;
        RECT 30.475 151.275 30.705 152.095 ;
        RECT 30.875 151.295 31.205 151.925 ;
        RECT 30.455 150.855 30.785 151.105 ;
        RECT 30.050 150.685 30.265 150.735 ;
        RECT 30.955 150.695 31.205 151.295 ;
        RECT 31.375 151.275 31.585 152.095 ;
        RECT 32.745 151.285 33.015 152.095 ;
        RECT 33.185 151.285 33.515 151.925 ;
        RECT 33.685 151.285 33.925 152.095 ;
        RECT 34.120 151.330 34.575 152.095 ;
        RECT 34.850 151.715 36.150 151.925 ;
        RECT 36.405 151.735 36.735 152.095 ;
        RECT 35.980 151.565 36.150 151.715 ;
        RECT 36.905 151.595 37.165 151.925 ;
        RECT 32.735 150.855 33.085 151.105 ;
        RECT 28.470 150.275 29.365 150.650 ;
        RECT 29.875 150.605 30.265 150.685 ;
        RECT 27.415 149.845 28.300 150.015 ;
        RECT 28.480 149.545 28.795 150.045 ;
        RECT 29.025 149.715 29.365 150.275 ;
        RECT 29.535 149.545 29.705 150.555 ;
        RECT 29.875 149.760 30.205 150.605 ;
        RECT 30.475 149.545 30.705 150.685 ;
        RECT 30.875 149.715 31.205 150.695 ;
        RECT 33.255 150.685 33.425 151.285 ;
        RECT 35.050 151.105 35.270 151.505 ;
        RECT 33.595 150.855 33.945 151.105 ;
        RECT 34.115 150.905 34.605 151.105 ;
        RECT 34.795 150.895 35.270 151.105 ;
        RECT 35.515 151.105 35.725 151.505 ;
        RECT 35.980 151.440 36.735 151.565 ;
        RECT 35.980 151.395 36.825 151.440 ;
        RECT 36.555 151.275 36.825 151.395 ;
        RECT 35.515 150.895 35.845 151.105 ;
        RECT 36.015 150.835 36.425 151.140 ;
        RECT 31.375 149.545 31.585 150.685 ;
        RECT 32.745 149.545 33.075 150.685 ;
        RECT 33.255 150.515 33.935 150.685 ;
        RECT 33.605 149.730 33.935 150.515 ;
        RECT 34.120 150.665 35.295 150.725 ;
        RECT 36.655 150.700 36.825 151.275 ;
        RECT 36.625 150.665 36.825 150.700 ;
        RECT 34.120 150.555 36.825 150.665 ;
        RECT 34.120 149.935 34.375 150.555 ;
        RECT 34.965 150.495 36.765 150.555 ;
        RECT 34.965 150.465 35.295 150.495 ;
        RECT 36.995 150.395 37.165 151.595 ;
        RECT 37.335 151.325 39.005 152.095 ;
        RECT 39.175 151.370 39.465 152.095 ;
        RECT 39.635 151.705 40.895 151.885 ;
        RECT 37.335 150.805 38.085 151.325 ;
        RECT 38.255 150.635 39.005 151.155 ;
        RECT 34.625 150.295 34.810 150.385 ;
        RECT 35.400 150.295 36.235 150.305 ;
        RECT 34.625 150.095 36.235 150.295 ;
        RECT 34.625 150.055 34.855 150.095 ;
        RECT 34.120 149.715 34.455 149.935 ;
        RECT 35.460 149.545 35.815 149.925 ;
        RECT 35.985 149.715 36.235 150.095 ;
        RECT 36.485 149.545 36.735 150.325 ;
        RECT 36.905 149.715 37.165 150.395 ;
        RECT 37.335 149.545 39.005 150.635 ;
        RECT 39.175 149.545 39.465 150.710 ;
        RECT 39.635 150.190 39.875 151.515 ;
        RECT 40.045 151.355 40.395 151.535 ;
        RECT 40.565 151.485 40.895 151.705 ;
        RECT 41.085 151.655 41.255 152.095 ;
        RECT 41.425 151.485 41.765 151.900 ;
        RECT 41.935 151.550 47.280 152.095 ;
        RECT 40.565 151.355 41.765 151.485 ;
        RECT 40.045 150.345 40.215 151.355 ;
        RECT 40.735 151.315 41.765 151.355 ;
        RECT 40.385 150.765 40.555 151.185 ;
        RECT 40.770 150.935 41.135 151.105 ;
        RECT 40.385 150.515 40.785 150.765 ;
        RECT 40.955 150.735 41.135 150.935 ;
        RECT 41.305 150.905 41.765 151.105 ;
        RECT 40.955 150.565 41.275 150.735 ;
        RECT 40.045 150.135 40.885 150.345 ;
        RECT 39.685 149.545 39.895 150.005 ;
        RECT 40.385 149.715 40.885 150.135 ;
        RECT 41.075 149.775 41.275 150.565 ;
        RECT 41.445 149.545 41.765 150.725 ;
        RECT 43.520 150.720 43.860 151.550 ;
        RECT 47.455 151.325 50.045 152.095 ;
        RECT 50.265 151.440 50.595 151.875 ;
        RECT 50.765 151.485 50.935 152.095 ;
        RECT 50.215 151.355 50.595 151.440 ;
        RECT 51.105 151.355 51.435 151.880 ;
        RECT 51.695 151.565 51.905 152.095 ;
        RECT 52.180 151.645 52.965 151.815 ;
        RECT 53.135 151.645 53.540 151.815 ;
        RECT 45.340 149.980 45.690 151.230 ;
        RECT 47.455 150.805 48.665 151.325 ;
        RECT 50.215 151.315 50.440 151.355 ;
        RECT 48.835 150.635 50.045 151.155 ;
        RECT 41.935 149.545 47.280 149.980 ;
        RECT 47.455 149.545 50.045 150.635 ;
        RECT 50.215 150.735 50.385 151.315 ;
        RECT 51.105 151.185 51.305 151.355 ;
        RECT 52.180 151.185 52.350 151.645 ;
        RECT 50.555 150.855 51.305 151.185 ;
        RECT 51.475 150.855 52.350 151.185 ;
        RECT 50.215 150.685 50.430 150.735 ;
        RECT 50.215 150.605 50.605 150.685 ;
        RECT 50.275 149.760 50.605 150.605 ;
        RECT 51.115 150.650 51.305 150.855 ;
        RECT 50.775 149.545 50.945 150.555 ;
        RECT 51.115 150.275 52.010 150.650 ;
        RECT 51.115 149.715 51.455 150.275 ;
        RECT 51.685 149.545 52.000 150.045 ;
        RECT 52.180 150.015 52.350 150.855 ;
        RECT 52.520 151.145 52.985 151.475 ;
        RECT 53.370 151.415 53.540 151.645 ;
        RECT 53.720 151.595 54.090 152.095 ;
        RECT 54.410 151.645 55.085 151.815 ;
        RECT 55.280 151.645 55.615 151.815 ;
        RECT 52.520 150.185 52.840 151.145 ;
        RECT 53.370 151.115 54.200 151.415 ;
        RECT 53.010 150.215 53.200 150.935 ;
        RECT 53.370 150.045 53.540 151.115 ;
        RECT 54.000 151.085 54.200 151.115 ;
        RECT 53.710 150.865 53.880 150.935 ;
        RECT 54.410 150.865 54.580 151.645 ;
        RECT 55.445 151.505 55.615 151.645 ;
        RECT 55.785 151.635 56.035 152.095 ;
        RECT 53.710 150.695 54.580 150.865 ;
        RECT 54.750 151.225 55.275 151.445 ;
        RECT 55.445 151.375 55.670 151.505 ;
        RECT 53.710 150.605 54.220 150.695 ;
        RECT 52.180 149.845 53.065 150.015 ;
        RECT 53.290 149.715 53.540 150.045 ;
        RECT 53.710 149.545 53.880 150.345 ;
        RECT 54.050 149.990 54.220 150.605 ;
        RECT 54.750 150.525 54.920 151.225 ;
        RECT 54.390 150.160 54.920 150.525 ;
        RECT 55.090 150.460 55.330 151.055 ;
        RECT 55.500 150.270 55.670 151.375 ;
        RECT 55.840 150.515 56.120 151.465 ;
        RECT 55.365 150.140 55.670 150.270 ;
        RECT 54.050 149.820 55.155 149.990 ;
        RECT 55.365 149.715 55.615 150.140 ;
        RECT 55.785 149.545 56.050 150.005 ;
        RECT 56.290 149.715 56.475 151.835 ;
        RECT 56.645 151.715 56.975 152.095 ;
        RECT 57.145 151.545 57.315 151.835 ;
        RECT 56.650 151.375 57.315 151.545 ;
        RECT 57.665 151.545 57.835 151.835 ;
        RECT 58.005 151.715 58.335 152.095 ;
        RECT 57.665 151.375 58.330 151.545 ;
        RECT 56.650 150.385 56.880 151.375 ;
        RECT 57.050 150.555 57.400 151.205 ;
        RECT 57.580 150.555 57.930 151.205 ;
        RECT 58.100 150.385 58.330 151.375 ;
        RECT 56.650 150.215 57.315 150.385 ;
        RECT 56.645 149.545 56.975 150.045 ;
        RECT 57.145 149.715 57.315 150.215 ;
        RECT 57.665 150.215 58.330 150.385 ;
        RECT 57.665 149.715 57.835 150.215 ;
        RECT 58.005 149.545 58.335 150.045 ;
        RECT 58.505 149.715 58.690 151.835 ;
        RECT 58.945 151.635 59.195 152.095 ;
        RECT 59.365 151.645 59.700 151.815 ;
        RECT 59.895 151.645 60.570 151.815 ;
        RECT 59.365 151.505 59.535 151.645 ;
        RECT 58.860 150.515 59.140 151.465 ;
        RECT 59.310 151.375 59.535 151.505 ;
        RECT 59.310 150.270 59.480 151.375 ;
        RECT 59.705 151.225 60.230 151.445 ;
        RECT 59.650 150.460 59.890 151.055 ;
        RECT 60.060 150.525 60.230 151.225 ;
        RECT 60.400 150.865 60.570 151.645 ;
        RECT 60.890 151.595 61.260 152.095 ;
        RECT 61.440 151.645 61.845 151.815 ;
        RECT 62.015 151.645 62.800 151.815 ;
        RECT 61.440 151.415 61.610 151.645 ;
        RECT 60.780 151.115 61.610 151.415 ;
        RECT 61.995 151.145 62.460 151.475 ;
        RECT 60.780 151.085 60.980 151.115 ;
        RECT 61.100 150.865 61.270 150.935 ;
        RECT 60.400 150.695 61.270 150.865 ;
        RECT 60.760 150.605 61.270 150.695 ;
        RECT 59.310 150.140 59.615 150.270 ;
        RECT 60.060 150.160 60.590 150.525 ;
        RECT 58.930 149.545 59.195 150.005 ;
        RECT 59.365 149.715 59.615 150.140 ;
        RECT 60.760 149.990 60.930 150.605 ;
        RECT 59.825 149.820 60.930 149.990 ;
        RECT 61.100 149.545 61.270 150.345 ;
        RECT 61.440 150.045 61.610 151.115 ;
        RECT 61.780 150.215 61.970 150.935 ;
        RECT 62.140 150.185 62.460 151.145 ;
        RECT 62.630 151.185 62.800 151.645 ;
        RECT 63.075 151.565 63.285 152.095 ;
        RECT 63.545 151.355 63.875 151.880 ;
        RECT 64.045 151.485 64.215 152.095 ;
        RECT 64.385 151.440 64.715 151.875 ;
        RECT 64.385 151.355 64.765 151.440 ;
        RECT 64.935 151.370 65.225 152.095 ;
        RECT 65.875 151.585 66.115 152.095 ;
        RECT 63.675 151.185 63.875 151.355 ;
        RECT 64.540 151.315 64.765 151.355 ;
        RECT 62.630 150.855 63.505 151.185 ;
        RECT 63.675 150.855 64.425 151.185 ;
        RECT 61.440 149.715 61.690 150.045 ;
        RECT 62.630 150.015 62.800 150.855 ;
        RECT 63.675 150.650 63.865 150.855 ;
        RECT 64.595 150.735 64.765 151.315 ;
        RECT 65.860 150.855 66.115 151.415 ;
        RECT 66.285 151.355 66.615 151.890 ;
        RECT 66.830 151.355 67.000 152.095 ;
        RECT 67.210 151.445 67.540 151.915 ;
        RECT 67.710 151.615 67.880 152.095 ;
        RECT 68.050 151.445 68.380 151.915 ;
        RECT 68.550 151.615 68.720 152.095 ;
        RECT 64.550 150.685 64.765 150.735 ;
        RECT 62.970 150.275 63.865 150.650 ;
        RECT 64.375 150.605 64.765 150.685 ;
        RECT 61.915 149.845 62.800 150.015 ;
        RECT 62.980 149.545 63.295 150.045 ;
        RECT 63.525 149.715 63.865 150.275 ;
        RECT 64.035 149.545 64.205 150.555 ;
        RECT 64.375 149.760 64.705 150.605 ;
        RECT 64.935 149.545 65.225 150.710 ;
        RECT 66.285 150.685 66.465 151.355 ;
        RECT 67.210 151.275 68.905 151.445 ;
        RECT 69.125 151.440 69.455 151.875 ;
        RECT 69.625 151.485 69.795 152.095 ;
        RECT 66.635 150.855 67.010 151.185 ;
        RECT 67.180 150.935 68.390 151.105 ;
        RECT 67.180 150.685 67.385 150.935 ;
        RECT 68.560 150.685 68.905 151.275 ;
        RECT 65.925 150.515 67.385 150.685 ;
        RECT 68.050 150.515 68.905 150.685 ;
        RECT 69.075 151.355 69.455 151.440 ;
        RECT 69.965 151.355 70.295 151.880 ;
        RECT 70.555 151.565 70.765 152.095 ;
        RECT 71.040 151.645 71.825 151.815 ;
        RECT 71.995 151.645 72.400 151.815 ;
        RECT 69.075 151.315 69.300 151.355 ;
        RECT 69.075 150.735 69.245 151.315 ;
        RECT 69.965 151.185 70.165 151.355 ;
        RECT 71.040 151.185 71.210 151.645 ;
        RECT 69.415 150.855 70.165 151.185 ;
        RECT 70.335 150.855 71.210 151.185 ;
        RECT 69.075 150.685 69.290 150.735 ;
        RECT 69.075 150.605 69.465 150.685 ;
        RECT 65.925 149.715 66.285 150.515 ;
        RECT 68.050 150.345 68.380 150.515 ;
        RECT 66.830 149.545 67.000 150.345 ;
        RECT 67.210 150.175 68.380 150.345 ;
        RECT 67.210 149.715 67.540 150.175 ;
        RECT 67.710 149.545 67.880 150.005 ;
        RECT 68.050 149.715 68.380 150.175 ;
        RECT 68.550 149.545 68.720 150.345 ;
        RECT 69.135 149.760 69.465 150.605 ;
        RECT 69.975 150.650 70.165 150.855 ;
        RECT 69.635 149.545 69.805 150.555 ;
        RECT 69.975 150.275 70.870 150.650 ;
        RECT 69.975 149.715 70.315 150.275 ;
        RECT 70.545 149.545 70.860 150.045 ;
        RECT 71.040 150.015 71.210 150.855 ;
        RECT 71.380 151.145 71.845 151.475 ;
        RECT 72.230 151.415 72.400 151.645 ;
        RECT 72.580 151.595 72.950 152.095 ;
        RECT 73.270 151.645 73.945 151.815 ;
        RECT 74.140 151.645 74.475 151.815 ;
        RECT 71.380 150.185 71.700 151.145 ;
        RECT 72.230 151.115 73.060 151.415 ;
        RECT 71.870 150.215 72.060 150.935 ;
        RECT 72.230 150.045 72.400 151.115 ;
        RECT 72.860 151.085 73.060 151.115 ;
        RECT 72.570 150.865 72.740 150.935 ;
        RECT 73.270 150.865 73.440 151.645 ;
        RECT 74.305 151.505 74.475 151.645 ;
        RECT 74.645 151.635 74.895 152.095 ;
        RECT 72.570 150.695 73.440 150.865 ;
        RECT 73.610 151.225 74.135 151.445 ;
        RECT 74.305 151.375 74.530 151.505 ;
        RECT 72.570 150.605 73.080 150.695 ;
        RECT 71.040 149.845 71.925 150.015 ;
        RECT 72.150 149.715 72.400 150.045 ;
        RECT 72.570 149.545 72.740 150.345 ;
        RECT 72.910 149.990 73.080 150.605 ;
        RECT 73.610 150.525 73.780 151.225 ;
        RECT 73.250 150.160 73.780 150.525 ;
        RECT 73.950 150.460 74.190 151.055 ;
        RECT 74.360 150.270 74.530 151.375 ;
        RECT 74.700 150.515 74.980 151.465 ;
        RECT 74.225 150.140 74.530 150.270 ;
        RECT 72.910 149.820 74.015 149.990 ;
        RECT 74.225 149.715 74.475 150.140 ;
        RECT 74.645 149.545 74.910 150.005 ;
        RECT 75.150 149.715 75.335 151.835 ;
        RECT 75.505 151.715 75.835 152.095 ;
        RECT 76.005 151.545 76.175 151.835 ;
        RECT 75.510 151.375 76.175 151.545 ;
        RECT 76.525 151.545 76.695 151.835 ;
        RECT 76.865 151.715 77.195 152.095 ;
        RECT 76.525 151.375 77.190 151.545 ;
        RECT 75.510 150.385 75.740 151.375 ;
        RECT 75.910 150.555 76.260 151.205 ;
        RECT 76.440 150.555 76.790 151.205 ;
        RECT 76.960 150.385 77.190 151.375 ;
        RECT 75.510 150.215 76.175 150.385 ;
        RECT 75.505 149.545 75.835 150.045 ;
        RECT 76.005 149.715 76.175 150.215 ;
        RECT 76.525 150.215 77.190 150.385 ;
        RECT 76.525 149.715 76.695 150.215 ;
        RECT 76.865 149.545 77.195 150.045 ;
        RECT 77.365 149.715 77.550 151.835 ;
        RECT 77.805 151.635 78.055 152.095 ;
        RECT 78.225 151.645 78.560 151.815 ;
        RECT 78.755 151.645 79.430 151.815 ;
        RECT 78.225 151.505 78.395 151.645 ;
        RECT 77.720 150.515 78.000 151.465 ;
        RECT 78.170 151.375 78.395 151.505 ;
        RECT 78.170 150.270 78.340 151.375 ;
        RECT 78.565 151.225 79.090 151.445 ;
        RECT 78.510 150.460 78.750 151.055 ;
        RECT 78.920 150.525 79.090 151.225 ;
        RECT 79.260 150.865 79.430 151.645 ;
        RECT 79.750 151.595 80.120 152.095 ;
        RECT 80.300 151.645 80.705 151.815 ;
        RECT 80.875 151.645 81.660 151.815 ;
        RECT 80.300 151.415 80.470 151.645 ;
        RECT 79.640 151.115 80.470 151.415 ;
        RECT 80.855 151.145 81.320 151.475 ;
        RECT 79.640 151.085 79.840 151.115 ;
        RECT 79.960 150.865 80.130 150.935 ;
        RECT 79.260 150.695 80.130 150.865 ;
        RECT 79.620 150.605 80.130 150.695 ;
        RECT 78.170 150.140 78.475 150.270 ;
        RECT 78.920 150.160 79.450 150.525 ;
        RECT 77.790 149.545 78.055 150.005 ;
        RECT 78.225 149.715 78.475 150.140 ;
        RECT 79.620 149.990 79.790 150.605 ;
        RECT 78.685 149.820 79.790 149.990 ;
        RECT 79.960 149.545 80.130 150.345 ;
        RECT 80.300 150.045 80.470 151.115 ;
        RECT 80.640 150.215 80.830 150.935 ;
        RECT 81.000 150.185 81.320 151.145 ;
        RECT 81.490 151.185 81.660 151.645 ;
        RECT 81.935 151.565 82.145 152.095 ;
        RECT 82.405 151.355 82.735 151.880 ;
        RECT 82.905 151.485 83.075 152.095 ;
        RECT 83.245 151.440 83.575 151.875 ;
        RECT 83.245 151.355 83.625 151.440 ;
        RECT 82.535 151.185 82.735 151.355 ;
        RECT 83.400 151.315 83.625 151.355 ;
        RECT 81.490 150.855 82.365 151.185 ;
        RECT 82.535 150.855 83.285 151.185 ;
        RECT 80.300 149.715 80.550 150.045 ;
        RECT 81.490 150.015 81.660 150.855 ;
        RECT 82.535 150.650 82.725 150.855 ;
        RECT 83.455 150.735 83.625 151.315 ;
        RECT 83.410 150.685 83.625 150.735 ;
        RECT 81.830 150.275 82.725 150.650 ;
        RECT 83.235 150.605 83.625 150.685 ;
        RECT 83.800 151.355 84.055 151.925 ;
        RECT 84.225 151.695 84.555 152.095 ;
        RECT 84.980 151.560 85.510 151.925 ;
        RECT 85.700 151.755 85.975 151.925 ;
        RECT 85.695 151.585 85.975 151.755 ;
        RECT 84.980 151.525 85.155 151.560 ;
        RECT 84.225 151.355 85.155 151.525 ;
        RECT 83.800 150.685 83.970 151.355 ;
        RECT 84.225 151.185 84.395 151.355 ;
        RECT 84.140 150.855 84.395 151.185 ;
        RECT 84.620 150.855 84.815 151.185 ;
        RECT 80.775 149.845 81.660 150.015 ;
        RECT 81.840 149.545 82.155 150.045 ;
        RECT 82.385 149.715 82.725 150.275 ;
        RECT 82.895 149.545 83.065 150.555 ;
        RECT 83.235 149.760 83.565 150.605 ;
        RECT 83.800 149.715 84.135 150.685 ;
        RECT 84.305 149.545 84.475 150.685 ;
        RECT 84.645 149.885 84.815 150.855 ;
        RECT 84.985 150.225 85.155 151.355 ;
        RECT 85.325 150.565 85.495 151.365 ;
        RECT 85.700 150.765 85.975 151.585 ;
        RECT 86.145 150.565 86.335 151.925 ;
        RECT 86.515 151.560 87.025 152.095 ;
        RECT 87.245 151.285 87.490 151.890 ;
        RECT 87.935 151.325 90.525 152.095 ;
        RECT 90.695 151.370 90.985 152.095 ;
        RECT 91.160 151.355 91.415 151.925 ;
        RECT 91.585 151.695 91.915 152.095 ;
        RECT 92.340 151.560 92.870 151.925 ;
        RECT 92.340 151.525 92.515 151.560 ;
        RECT 91.585 151.355 92.515 151.525 ;
        RECT 86.535 151.115 87.765 151.285 ;
        RECT 85.325 150.395 86.335 150.565 ;
        RECT 86.505 150.550 87.255 150.740 ;
        RECT 84.985 150.055 86.110 150.225 ;
        RECT 86.505 149.885 86.675 150.550 ;
        RECT 87.425 150.305 87.765 151.115 ;
        RECT 87.935 150.805 89.145 151.325 ;
        RECT 89.315 150.635 90.525 151.155 ;
        RECT 84.645 149.715 86.675 149.885 ;
        RECT 86.845 149.545 87.015 150.305 ;
        RECT 87.250 149.895 87.765 150.305 ;
        RECT 87.935 149.545 90.525 150.635 ;
        RECT 90.695 149.545 90.985 150.710 ;
        RECT 91.160 150.685 91.330 151.355 ;
        RECT 91.585 151.185 91.755 151.355 ;
        RECT 91.500 150.855 91.755 151.185 ;
        RECT 91.980 150.855 92.175 151.185 ;
        RECT 91.160 149.715 91.495 150.685 ;
        RECT 91.665 149.545 91.835 150.685 ;
        RECT 92.005 149.885 92.175 150.855 ;
        RECT 92.345 150.225 92.515 151.355 ;
        RECT 92.685 150.565 92.855 151.365 ;
        RECT 93.060 151.075 93.335 151.925 ;
        RECT 93.055 150.905 93.335 151.075 ;
        RECT 93.060 150.765 93.335 150.905 ;
        RECT 93.505 150.565 93.695 151.925 ;
        RECT 93.875 151.560 94.385 152.095 ;
        RECT 94.605 151.285 94.850 151.890 ;
        RECT 95.295 151.355 95.680 151.925 ;
        RECT 95.850 151.635 96.175 152.095 ;
        RECT 96.695 151.465 96.975 151.925 ;
        RECT 93.895 151.115 95.125 151.285 ;
        RECT 92.685 150.395 93.695 150.565 ;
        RECT 93.865 150.550 94.615 150.740 ;
        RECT 92.345 150.055 93.470 150.225 ;
        RECT 93.865 149.885 94.035 150.550 ;
        RECT 94.785 150.305 95.125 151.115 ;
        RECT 92.005 149.715 94.035 149.885 ;
        RECT 94.205 149.545 94.375 150.305 ;
        RECT 94.610 149.895 95.125 150.305 ;
        RECT 95.295 150.685 95.575 151.355 ;
        RECT 95.850 151.295 96.975 151.465 ;
        RECT 95.850 151.185 96.300 151.295 ;
        RECT 95.745 150.855 96.300 151.185 ;
        RECT 97.165 151.125 97.565 151.925 ;
        RECT 97.965 151.635 98.235 152.095 ;
        RECT 98.405 151.465 98.690 151.925 ;
        RECT 98.975 151.550 104.320 152.095 ;
        RECT 104.495 151.550 109.840 152.095 ;
        RECT 110.015 151.550 115.360 152.095 ;
        RECT 95.295 149.715 95.680 150.685 ;
        RECT 95.850 150.395 96.300 150.855 ;
        RECT 96.470 150.565 97.565 151.125 ;
        RECT 95.850 150.175 96.975 150.395 ;
        RECT 95.850 149.545 96.175 150.005 ;
        RECT 96.695 149.715 96.975 150.175 ;
        RECT 97.165 149.715 97.565 150.565 ;
        RECT 97.735 151.295 98.690 151.465 ;
        RECT 97.735 150.395 97.945 151.295 ;
        RECT 98.115 150.565 98.805 151.125 ;
        RECT 100.560 150.720 100.900 151.550 ;
        RECT 97.735 150.175 98.690 150.395 ;
        RECT 97.965 149.545 98.235 150.005 ;
        RECT 98.405 149.715 98.690 150.175 ;
        RECT 102.380 149.980 102.730 151.230 ;
        RECT 106.080 150.720 106.420 151.550 ;
        RECT 107.900 149.980 108.250 151.230 ;
        RECT 111.600 150.720 111.940 151.550 ;
        RECT 116.455 151.370 116.745 152.095 ;
        RECT 117.835 151.295 118.145 152.095 ;
        RECT 118.350 151.295 119.045 151.925 ;
        RECT 119.215 151.325 122.725 152.095 ;
        RECT 122.895 151.345 124.105 152.095 ;
        RECT 124.280 151.355 124.535 151.925 ;
        RECT 124.705 151.695 125.035 152.095 ;
        RECT 125.460 151.560 125.990 151.925 ;
        RECT 126.180 151.755 126.455 151.925 ;
        RECT 126.175 151.585 126.455 151.755 ;
        RECT 125.460 151.525 125.635 151.560 ;
        RECT 124.705 151.355 125.635 151.525 ;
        RECT 118.350 151.245 118.525 151.295 ;
        RECT 113.420 149.980 113.770 151.230 ;
        RECT 117.845 150.855 118.180 151.125 ;
        RECT 98.975 149.545 104.320 149.980 ;
        RECT 104.495 149.545 109.840 149.980 ;
        RECT 110.015 149.545 115.360 149.980 ;
        RECT 116.455 149.545 116.745 150.710 ;
        RECT 118.350 150.695 118.520 151.245 ;
        RECT 118.690 150.855 119.025 151.105 ;
        RECT 119.215 150.805 120.865 151.325 ;
        RECT 117.835 149.545 118.115 150.685 ;
        RECT 118.285 149.715 118.615 150.695 ;
        RECT 118.785 149.545 119.045 150.685 ;
        RECT 121.035 150.635 122.725 151.155 ;
        RECT 122.895 150.805 123.415 151.345 ;
        RECT 123.585 150.635 124.105 151.175 ;
        RECT 119.215 149.545 122.725 150.635 ;
        RECT 122.895 149.545 124.105 150.635 ;
        RECT 124.280 150.685 124.450 151.355 ;
        RECT 124.705 151.185 124.875 151.355 ;
        RECT 124.620 150.855 124.875 151.185 ;
        RECT 125.100 150.855 125.295 151.185 ;
        RECT 124.280 149.715 124.615 150.685 ;
        RECT 124.785 149.545 124.955 150.685 ;
        RECT 125.125 149.885 125.295 150.855 ;
        RECT 125.465 150.225 125.635 151.355 ;
        RECT 125.805 150.565 125.975 151.365 ;
        RECT 126.180 150.765 126.455 151.585 ;
        RECT 126.625 150.565 126.815 151.925 ;
        RECT 126.995 151.560 127.505 152.095 ;
        RECT 127.725 151.285 127.970 151.890 ;
        RECT 128.415 151.325 131.925 152.095 ;
        RECT 132.645 151.545 132.815 151.925 ;
        RECT 132.995 151.715 133.325 152.095 ;
        RECT 132.645 151.375 133.310 151.545 ;
        RECT 133.505 151.420 133.765 151.925 ;
        RECT 127.015 151.115 128.245 151.285 ;
        RECT 125.805 150.395 126.815 150.565 ;
        RECT 126.985 150.550 127.735 150.740 ;
        RECT 125.465 150.055 126.590 150.225 ;
        RECT 126.985 149.885 127.155 150.550 ;
        RECT 127.905 150.305 128.245 151.115 ;
        RECT 128.415 150.805 130.065 151.325 ;
        RECT 130.235 150.635 131.925 151.155 ;
        RECT 132.575 150.825 132.905 151.195 ;
        RECT 133.140 151.120 133.310 151.375 ;
        RECT 133.140 150.790 133.425 151.120 ;
        RECT 133.140 150.645 133.310 150.790 ;
        RECT 125.125 149.715 127.155 149.885 ;
        RECT 127.325 149.545 127.495 150.305 ;
        RECT 127.730 149.895 128.245 150.305 ;
        RECT 128.415 149.545 131.925 150.635 ;
        RECT 132.645 150.475 133.310 150.645 ;
        RECT 133.595 150.620 133.765 151.420 ;
        RECT 133.935 151.325 137.445 152.095 ;
        RECT 137.615 151.345 138.825 152.095 ;
        RECT 133.935 150.805 135.585 151.325 ;
        RECT 135.755 150.635 137.445 151.155 ;
        RECT 132.645 149.715 132.815 150.475 ;
        RECT 132.995 149.545 133.325 150.305 ;
        RECT 133.495 149.715 133.765 150.620 ;
        RECT 133.935 149.545 137.445 150.635 ;
        RECT 137.615 150.635 138.135 151.175 ;
        RECT 138.305 150.805 138.825 151.345 ;
        RECT 137.615 149.545 138.825 150.635 ;
        RECT 13.330 149.375 138.910 149.545 ;
        RECT 13.415 148.285 14.625 149.375 ;
        RECT 14.795 148.285 16.465 149.375 ;
        RECT 16.725 148.705 16.895 149.205 ;
        RECT 17.065 148.875 17.395 149.375 ;
        RECT 16.725 148.535 17.390 148.705 ;
        RECT 13.415 147.575 13.935 148.115 ;
        RECT 14.105 147.745 14.625 148.285 ;
        RECT 14.795 147.595 15.545 148.115 ;
        RECT 15.715 147.765 16.465 148.285 ;
        RECT 16.640 147.715 16.990 148.365 ;
        RECT 13.415 146.825 14.625 147.575 ;
        RECT 14.795 146.825 16.465 147.595 ;
        RECT 17.160 147.545 17.390 148.535 ;
        RECT 16.725 147.375 17.390 147.545 ;
        RECT 16.725 147.085 16.895 147.375 ;
        RECT 17.065 146.825 17.395 147.205 ;
        RECT 17.565 147.085 17.750 149.205 ;
        RECT 17.990 148.915 18.255 149.375 ;
        RECT 18.425 148.780 18.675 149.205 ;
        RECT 18.885 148.930 19.990 149.100 ;
        RECT 18.370 148.650 18.675 148.780 ;
        RECT 17.920 147.455 18.200 148.405 ;
        RECT 18.370 147.545 18.540 148.650 ;
        RECT 18.710 147.865 18.950 148.460 ;
        RECT 19.120 148.395 19.650 148.760 ;
        RECT 19.120 147.695 19.290 148.395 ;
        RECT 19.820 148.315 19.990 148.930 ;
        RECT 20.160 148.575 20.330 149.375 ;
        RECT 20.500 148.875 20.750 149.205 ;
        RECT 20.975 148.905 21.860 149.075 ;
        RECT 19.820 148.225 20.330 148.315 ;
        RECT 18.370 147.415 18.595 147.545 ;
        RECT 18.765 147.475 19.290 147.695 ;
        RECT 19.460 148.055 20.330 148.225 ;
        RECT 18.005 146.825 18.255 147.285 ;
        RECT 18.425 147.275 18.595 147.415 ;
        RECT 19.460 147.275 19.630 148.055 ;
        RECT 20.160 147.985 20.330 148.055 ;
        RECT 19.840 147.805 20.040 147.835 ;
        RECT 20.500 147.805 20.670 148.875 ;
        RECT 20.840 147.985 21.030 148.705 ;
        RECT 19.840 147.505 20.670 147.805 ;
        RECT 21.200 147.775 21.520 148.735 ;
        RECT 18.425 147.105 18.760 147.275 ;
        RECT 18.955 147.105 19.630 147.275 ;
        RECT 19.950 146.825 20.320 147.325 ;
        RECT 20.500 147.275 20.670 147.505 ;
        RECT 21.055 147.445 21.520 147.775 ;
        RECT 21.690 148.065 21.860 148.905 ;
        RECT 22.040 148.875 22.355 149.375 ;
        RECT 22.585 148.645 22.925 149.205 ;
        RECT 22.030 148.270 22.925 148.645 ;
        RECT 23.095 148.365 23.265 149.375 ;
        RECT 22.735 148.065 22.925 148.270 ;
        RECT 23.435 148.315 23.765 149.160 ;
        RECT 23.995 148.655 24.455 149.205 ;
        RECT 24.645 148.655 24.975 149.375 ;
        RECT 23.435 148.235 23.825 148.315 ;
        RECT 23.610 148.185 23.825 148.235 ;
        RECT 21.690 147.735 22.565 148.065 ;
        RECT 22.735 147.735 23.485 148.065 ;
        RECT 21.690 147.275 21.860 147.735 ;
        RECT 22.735 147.565 22.935 147.735 ;
        RECT 23.655 147.605 23.825 148.185 ;
        RECT 23.600 147.565 23.825 147.605 ;
        RECT 20.500 147.105 20.905 147.275 ;
        RECT 21.075 147.105 21.860 147.275 ;
        RECT 22.135 146.825 22.345 147.355 ;
        RECT 22.605 147.040 22.935 147.565 ;
        RECT 23.445 147.480 23.825 147.565 ;
        RECT 23.105 146.825 23.275 147.435 ;
        RECT 23.445 147.045 23.775 147.480 ;
        RECT 23.995 147.285 24.245 148.655 ;
        RECT 25.175 148.485 25.475 149.035 ;
        RECT 25.645 148.705 25.925 149.375 ;
        RECT 24.535 148.315 25.475 148.485 ;
        RECT 24.535 148.065 24.705 148.315 ;
        RECT 25.845 148.065 26.110 148.425 ;
        RECT 26.295 148.210 26.585 149.375 ;
        RECT 26.755 148.235 27.015 149.375 ;
        RECT 27.185 148.225 27.515 149.205 ;
        RECT 27.685 148.235 27.965 149.375 ;
        RECT 28.135 148.235 28.395 149.375 ;
        RECT 28.635 148.865 30.250 149.195 ;
        RECT 27.275 148.185 27.450 148.225 ;
        RECT 24.415 147.735 24.705 148.065 ;
        RECT 24.875 147.815 25.215 148.065 ;
        RECT 25.435 147.815 26.110 148.065 ;
        RECT 26.775 147.815 27.110 148.065 ;
        RECT 24.535 147.645 24.705 147.735 ;
        RECT 24.535 147.455 25.925 147.645 ;
        RECT 27.280 147.625 27.450 148.185 ;
        RECT 28.645 148.065 28.815 148.625 ;
        RECT 29.075 148.525 30.250 148.695 ;
        RECT 30.420 148.575 30.700 149.375 ;
        RECT 29.075 148.235 29.405 148.525 ;
        RECT 30.080 148.405 30.250 148.525 ;
        RECT 29.575 148.065 29.820 148.355 ;
        RECT 30.080 148.235 30.740 148.405 ;
        RECT 30.910 148.235 31.185 149.205 ;
        RECT 31.560 148.405 31.890 149.205 ;
        RECT 32.060 148.575 32.390 149.375 ;
        RECT 32.690 148.405 33.020 149.205 ;
        RECT 33.665 148.575 33.915 149.375 ;
        RECT 31.560 148.235 33.995 148.405 ;
        RECT 34.185 148.235 34.355 149.375 ;
        RECT 34.525 148.235 34.865 149.205 ;
        RECT 30.570 148.065 30.740 148.235 ;
        RECT 27.620 147.795 27.955 148.065 ;
        RECT 28.140 147.815 28.475 148.065 ;
        RECT 28.645 147.735 29.360 148.065 ;
        RECT 29.575 147.735 30.400 148.065 ;
        RECT 30.570 147.735 30.845 148.065 ;
        RECT 28.645 147.645 28.895 147.735 ;
        RECT 23.995 146.995 24.555 147.285 ;
        RECT 24.725 146.825 24.975 147.285 ;
        RECT 25.595 147.095 25.925 147.455 ;
        RECT 26.295 146.825 26.585 147.550 ;
        RECT 26.755 146.995 27.450 147.625 ;
        RECT 27.655 146.825 27.965 147.625 ;
        RECT 28.135 146.825 28.395 147.645 ;
        RECT 28.565 147.225 28.895 147.645 ;
        RECT 30.570 147.565 30.740 147.735 ;
        RECT 29.075 147.395 30.740 147.565 ;
        RECT 31.015 147.500 31.185 148.235 ;
        RECT 31.355 147.815 31.705 148.065 ;
        RECT 31.890 147.605 32.060 148.235 ;
        RECT 32.230 147.815 32.560 148.015 ;
        RECT 32.730 147.815 33.060 148.015 ;
        RECT 33.230 147.815 33.650 148.015 ;
        RECT 33.825 147.985 33.995 148.235 ;
        RECT 33.825 147.815 34.520 147.985 ;
        RECT 34.690 147.675 34.865 148.235 ;
        RECT 29.075 146.995 29.335 147.395 ;
        RECT 29.505 146.825 29.835 147.225 ;
        RECT 30.005 147.045 30.175 147.395 ;
        RECT 30.345 146.825 30.720 147.225 ;
        RECT 30.910 147.155 31.185 147.500 ;
        RECT 31.560 146.995 32.060 147.605 ;
        RECT 32.690 147.475 33.915 147.645 ;
        RECT 34.635 147.625 34.865 147.675 ;
        RECT 32.690 146.995 33.020 147.475 ;
        RECT 33.190 146.825 33.415 147.285 ;
        RECT 33.585 146.995 33.915 147.475 ;
        RECT 34.105 146.825 34.355 147.625 ;
        RECT 34.525 146.995 34.865 147.625 ;
        RECT 35.035 148.505 35.310 149.205 ;
        RECT 35.520 148.830 35.735 149.375 ;
        RECT 35.905 148.865 36.380 149.205 ;
        RECT 36.550 148.870 37.165 149.375 ;
        RECT 36.550 148.695 36.745 148.870 ;
        RECT 35.035 147.475 35.205 148.505 ;
        RECT 35.480 148.335 36.195 148.630 ;
        RECT 36.415 148.505 36.745 148.695 ;
        RECT 36.915 148.335 37.165 148.700 ;
        RECT 35.375 148.165 37.165 148.335 ;
        RECT 35.375 147.735 35.605 148.165 ;
        RECT 35.035 146.995 35.295 147.475 ;
        RECT 35.775 147.465 36.185 147.985 ;
        RECT 35.465 146.825 35.795 147.285 ;
        RECT 35.985 147.045 36.185 147.465 ;
        RECT 36.355 147.310 36.610 148.165 ;
        RECT 37.405 147.985 37.575 149.205 ;
        RECT 37.825 148.865 38.085 149.375 ;
        RECT 36.780 147.735 37.575 147.985 ;
        RECT 37.745 147.815 38.085 148.695 ;
        RECT 38.260 148.575 38.575 149.375 ;
        RECT 38.840 149.020 39.920 149.190 ;
        RECT 38.840 148.405 39.010 149.020 ;
        RECT 37.325 147.645 37.575 147.735 ;
        RECT 36.355 147.045 37.145 147.310 ;
        RECT 37.325 147.225 37.655 147.645 ;
        RECT 37.825 146.825 38.085 147.645 ;
        RECT 38.255 147.395 38.525 148.405 ;
        RECT 38.695 148.235 39.010 148.405 ;
        RECT 38.695 147.565 38.865 148.235 ;
        RECT 39.180 148.065 39.415 148.745 ;
        RECT 39.585 148.235 39.920 149.020 ;
        RECT 40.095 148.285 42.685 149.375 ;
        RECT 39.035 147.735 39.415 148.065 ;
        RECT 39.585 147.735 39.920 148.065 ;
        RECT 40.095 147.595 41.305 148.115 ;
        RECT 41.475 147.765 42.685 148.285 ;
        RECT 43.335 148.485 43.595 149.195 ;
        RECT 43.765 148.665 44.095 149.375 ;
        RECT 44.265 148.485 44.495 149.195 ;
        RECT 43.335 148.245 44.495 148.485 ;
        RECT 44.675 148.465 44.945 149.195 ;
        RECT 45.125 148.645 45.465 149.375 ;
        RECT 44.675 148.245 45.445 148.465 ;
        RECT 43.325 147.735 43.625 148.065 ;
        RECT 43.805 147.755 44.330 148.065 ;
        RECT 44.510 147.755 44.975 148.065 ;
        RECT 38.695 147.395 39.920 147.565 ;
        RECT 38.325 146.825 38.655 147.225 ;
        RECT 38.825 147.125 38.995 147.395 ;
        RECT 39.165 146.825 39.495 147.225 ;
        RECT 39.665 147.125 39.920 147.395 ;
        RECT 40.095 146.825 42.685 147.595 ;
        RECT 43.335 146.825 43.625 147.555 ;
        RECT 43.805 147.115 44.035 147.755 ;
        RECT 45.155 147.575 45.445 148.245 ;
        RECT 44.215 147.375 45.445 147.575 ;
        RECT 44.215 147.005 44.525 147.375 ;
        RECT 44.705 146.825 45.375 147.195 ;
        RECT 45.635 147.005 45.895 149.195 ;
        RECT 46.075 148.285 49.585 149.375 ;
        RECT 49.755 148.820 50.360 149.375 ;
        RECT 50.535 148.865 51.015 149.205 ;
        RECT 51.185 148.830 51.440 149.375 ;
        RECT 49.755 148.720 50.370 148.820 ;
        RECT 50.185 148.695 50.370 148.720 ;
        RECT 46.075 147.595 47.725 148.115 ;
        RECT 47.895 147.765 49.585 148.285 ;
        RECT 49.755 148.100 50.015 148.550 ;
        RECT 50.185 148.450 50.515 148.695 ;
        RECT 50.685 148.375 51.440 148.625 ;
        RECT 51.610 148.505 51.885 149.205 ;
        RECT 50.670 148.340 51.440 148.375 ;
        RECT 50.655 148.330 51.440 148.340 ;
        RECT 50.650 148.315 51.545 148.330 ;
        RECT 50.630 148.300 51.545 148.315 ;
        RECT 50.610 148.290 51.545 148.300 ;
        RECT 50.585 148.280 51.545 148.290 ;
        RECT 50.515 148.250 51.545 148.280 ;
        RECT 50.495 148.220 51.545 148.250 ;
        RECT 50.475 148.190 51.545 148.220 ;
        RECT 50.445 148.165 51.545 148.190 ;
        RECT 50.410 148.130 51.545 148.165 ;
        RECT 50.380 148.125 51.545 148.130 ;
        RECT 50.380 148.120 50.770 148.125 ;
        RECT 50.380 148.110 50.745 148.120 ;
        RECT 50.380 148.105 50.730 148.110 ;
        RECT 50.380 148.100 50.715 148.105 ;
        RECT 49.755 148.095 50.715 148.100 ;
        RECT 49.755 148.085 50.705 148.095 ;
        RECT 49.755 148.080 50.695 148.085 ;
        RECT 49.755 148.070 50.685 148.080 ;
        RECT 49.755 148.060 50.680 148.070 ;
        RECT 49.755 148.055 50.675 148.060 ;
        RECT 49.755 148.040 50.665 148.055 ;
        RECT 49.755 148.025 50.660 148.040 ;
        RECT 49.755 148.000 50.650 148.025 ;
        RECT 49.755 147.930 50.645 148.000 ;
        RECT 46.075 146.825 49.585 147.595 ;
        RECT 49.755 147.375 50.305 147.760 ;
        RECT 50.475 147.205 50.645 147.930 ;
        RECT 49.755 147.035 50.645 147.205 ;
        RECT 50.815 147.530 51.145 147.955 ;
        RECT 51.315 147.730 51.545 148.125 ;
        RECT 50.815 147.045 51.035 147.530 ;
        RECT 51.715 147.475 51.885 148.505 ;
        RECT 52.055 148.210 52.345 149.375 ;
        RECT 52.605 148.705 52.775 149.205 ;
        RECT 52.945 148.875 53.275 149.375 ;
        RECT 52.605 148.535 53.270 148.705 ;
        RECT 52.520 147.715 52.870 148.365 ;
        RECT 51.205 146.825 51.455 147.365 ;
        RECT 51.625 146.995 51.885 147.475 ;
        RECT 52.055 146.825 52.345 147.550 ;
        RECT 53.040 147.545 53.270 148.535 ;
        RECT 52.605 147.375 53.270 147.545 ;
        RECT 52.605 147.085 52.775 147.375 ;
        RECT 52.945 146.825 53.275 147.205 ;
        RECT 53.445 147.085 53.630 149.205 ;
        RECT 53.870 148.915 54.135 149.375 ;
        RECT 54.305 148.780 54.555 149.205 ;
        RECT 54.765 148.930 55.870 149.100 ;
        RECT 54.250 148.650 54.555 148.780 ;
        RECT 53.800 147.455 54.080 148.405 ;
        RECT 54.250 147.545 54.420 148.650 ;
        RECT 54.590 147.865 54.830 148.460 ;
        RECT 55.000 148.395 55.530 148.760 ;
        RECT 55.000 147.695 55.170 148.395 ;
        RECT 55.700 148.315 55.870 148.930 ;
        RECT 56.040 148.575 56.210 149.375 ;
        RECT 56.380 148.875 56.630 149.205 ;
        RECT 56.855 148.905 57.740 149.075 ;
        RECT 55.700 148.225 56.210 148.315 ;
        RECT 54.250 147.415 54.475 147.545 ;
        RECT 54.645 147.475 55.170 147.695 ;
        RECT 55.340 148.055 56.210 148.225 ;
        RECT 53.885 146.825 54.135 147.285 ;
        RECT 54.305 147.275 54.475 147.415 ;
        RECT 55.340 147.275 55.510 148.055 ;
        RECT 56.040 147.985 56.210 148.055 ;
        RECT 55.720 147.805 55.920 147.835 ;
        RECT 56.380 147.805 56.550 148.875 ;
        RECT 56.720 147.985 56.910 148.705 ;
        RECT 55.720 147.505 56.550 147.805 ;
        RECT 57.080 147.775 57.400 148.735 ;
        RECT 54.305 147.105 54.640 147.275 ;
        RECT 54.835 147.105 55.510 147.275 ;
        RECT 55.830 146.825 56.200 147.325 ;
        RECT 56.380 147.275 56.550 147.505 ;
        RECT 56.935 147.445 57.400 147.775 ;
        RECT 57.570 148.065 57.740 148.905 ;
        RECT 57.920 148.875 58.235 149.375 ;
        RECT 58.465 148.645 58.805 149.205 ;
        RECT 57.910 148.270 58.805 148.645 ;
        RECT 58.975 148.365 59.145 149.375 ;
        RECT 58.615 148.065 58.805 148.270 ;
        RECT 59.315 148.315 59.645 149.160 ;
        RECT 59.315 148.235 59.705 148.315 ;
        RECT 59.875 148.285 63.385 149.375 ;
        RECT 64.475 148.820 65.080 149.375 ;
        RECT 65.255 148.865 65.735 149.205 ;
        RECT 65.905 148.830 66.160 149.375 ;
        RECT 64.475 148.720 65.090 148.820 ;
        RECT 64.905 148.695 65.090 148.720 ;
        RECT 59.490 148.185 59.705 148.235 ;
        RECT 57.570 147.735 58.445 148.065 ;
        RECT 58.615 147.735 59.365 148.065 ;
        RECT 57.570 147.275 57.740 147.735 ;
        RECT 58.615 147.565 58.815 147.735 ;
        RECT 59.535 147.605 59.705 148.185 ;
        RECT 59.480 147.565 59.705 147.605 ;
        RECT 56.380 147.105 56.785 147.275 ;
        RECT 56.955 147.105 57.740 147.275 ;
        RECT 58.015 146.825 58.225 147.355 ;
        RECT 58.485 147.040 58.815 147.565 ;
        RECT 59.325 147.480 59.705 147.565 ;
        RECT 59.875 147.595 61.525 148.115 ;
        RECT 61.695 147.765 63.385 148.285 ;
        RECT 64.475 148.100 64.735 148.550 ;
        RECT 64.905 148.450 65.235 148.695 ;
        RECT 65.405 148.375 66.160 148.625 ;
        RECT 66.330 148.505 66.605 149.205 ;
        RECT 65.390 148.340 66.160 148.375 ;
        RECT 65.375 148.330 66.160 148.340 ;
        RECT 65.370 148.315 66.265 148.330 ;
        RECT 65.350 148.300 66.265 148.315 ;
        RECT 65.330 148.290 66.265 148.300 ;
        RECT 65.305 148.280 66.265 148.290 ;
        RECT 65.235 148.250 66.265 148.280 ;
        RECT 65.215 148.220 66.265 148.250 ;
        RECT 65.195 148.190 66.265 148.220 ;
        RECT 65.165 148.165 66.265 148.190 ;
        RECT 65.130 148.130 66.265 148.165 ;
        RECT 65.100 148.125 66.265 148.130 ;
        RECT 65.100 148.120 65.490 148.125 ;
        RECT 65.100 148.110 65.465 148.120 ;
        RECT 65.100 148.105 65.450 148.110 ;
        RECT 65.100 148.100 65.435 148.105 ;
        RECT 64.475 148.095 65.435 148.100 ;
        RECT 64.475 148.085 65.425 148.095 ;
        RECT 64.475 148.080 65.415 148.085 ;
        RECT 64.475 148.070 65.405 148.080 ;
        RECT 64.475 148.060 65.400 148.070 ;
        RECT 64.475 148.055 65.395 148.060 ;
        RECT 64.475 148.040 65.385 148.055 ;
        RECT 64.475 148.025 65.380 148.040 ;
        RECT 64.475 148.000 65.370 148.025 ;
        RECT 64.475 147.930 65.365 148.000 ;
        RECT 58.985 146.825 59.155 147.435 ;
        RECT 59.325 147.045 59.655 147.480 ;
        RECT 59.875 146.825 63.385 147.595 ;
        RECT 64.475 147.375 65.025 147.760 ;
        RECT 65.195 147.205 65.365 147.930 ;
        RECT 64.475 147.035 65.365 147.205 ;
        RECT 65.535 147.530 65.865 147.955 ;
        RECT 66.035 147.730 66.265 148.125 ;
        RECT 65.535 147.045 65.755 147.530 ;
        RECT 66.435 147.475 66.605 148.505 ;
        RECT 65.925 146.825 66.175 147.365 ;
        RECT 66.345 146.995 66.605 147.475 ;
        RECT 66.775 148.185 67.115 149.205 ;
        RECT 67.285 148.185 67.975 149.375 ;
        RECT 68.145 148.405 68.475 149.205 ;
        RECT 68.645 148.575 68.815 149.375 ;
        RECT 68.985 148.745 69.315 149.205 ;
        RECT 69.485 148.915 69.655 149.375 ;
        RECT 69.825 148.745 70.155 149.205 ;
        RECT 68.985 148.405 70.155 148.745 ;
        RECT 70.325 148.575 70.495 149.375 ;
        RECT 70.665 148.405 70.995 149.205 ;
        RECT 71.165 148.575 71.855 149.375 ;
        RECT 72.025 148.405 72.355 149.205 ;
        RECT 72.525 148.575 72.695 149.375 ;
        RECT 72.865 148.405 73.195 149.205 ;
        RECT 68.145 148.185 73.195 148.405 ;
        RECT 73.365 148.185 73.695 149.375 ;
        RECT 74.135 148.235 74.520 149.205 ;
        RECT 74.690 148.915 75.015 149.375 ;
        RECT 75.535 148.745 75.815 149.205 ;
        RECT 74.690 148.525 75.815 148.745 ;
        RECT 66.775 147.645 66.950 148.185 ;
        RECT 67.120 147.815 67.470 148.015 ;
        RECT 67.695 147.815 69.315 148.015 ;
        RECT 69.485 147.815 69.790 148.185 ;
        RECT 69.960 147.815 71.170 148.015 ;
        RECT 71.435 147.845 73.190 148.015 ;
        RECT 71.480 147.815 73.190 147.845 ;
        RECT 67.695 147.645 67.975 147.815 ;
        RECT 69.485 147.645 69.655 147.815 ;
        RECT 66.775 147.455 67.975 147.645 ;
        RECT 66.775 146.995 67.115 147.455 ;
        RECT 68.145 147.375 69.655 147.645 ;
        RECT 69.825 147.455 73.195 147.645 ;
        RECT 69.825 147.375 71.415 147.455 ;
        RECT 67.285 146.825 67.535 147.285 ;
        RECT 67.725 146.995 71.415 147.205 ;
        RECT 71.605 146.825 71.855 147.285 ;
        RECT 72.025 146.995 72.355 147.455 ;
        RECT 72.525 146.825 72.695 147.285 ;
        RECT 72.865 146.995 73.195 147.455 ;
        RECT 73.365 146.825 73.695 147.645 ;
        RECT 74.135 147.565 74.415 148.235 ;
        RECT 74.690 148.065 75.140 148.525 ;
        RECT 76.005 148.355 76.405 149.205 ;
        RECT 76.805 148.915 77.075 149.375 ;
        RECT 77.245 148.745 77.530 149.205 ;
        RECT 74.585 147.735 75.140 148.065 ;
        RECT 75.310 147.795 76.405 148.355 ;
        RECT 74.690 147.625 75.140 147.735 ;
        RECT 74.135 146.995 74.520 147.565 ;
        RECT 74.690 147.455 75.815 147.625 ;
        RECT 74.690 146.825 75.015 147.285 ;
        RECT 75.535 146.995 75.815 147.455 ;
        RECT 76.005 146.995 76.405 147.795 ;
        RECT 76.575 148.525 77.530 148.745 ;
        RECT 76.575 147.625 76.785 148.525 ;
        RECT 76.955 147.795 77.645 148.355 ;
        RECT 77.815 148.210 78.105 149.375 ;
        RECT 79.255 148.315 79.585 149.160 ;
        RECT 79.755 148.365 79.925 149.375 ;
        RECT 80.095 148.645 80.435 149.205 ;
        RECT 80.665 148.875 80.980 149.375 ;
        RECT 81.160 148.905 82.045 149.075 ;
        RECT 79.195 148.235 79.585 148.315 ;
        RECT 80.095 148.270 80.990 148.645 ;
        RECT 79.195 148.185 79.410 148.235 ;
        RECT 76.575 147.455 77.530 147.625 ;
        RECT 79.195 147.605 79.365 148.185 ;
        RECT 80.095 148.065 80.285 148.270 ;
        RECT 81.160 148.065 81.330 148.905 ;
        RECT 82.270 148.875 82.520 149.205 ;
        RECT 79.535 147.735 80.285 148.065 ;
        RECT 80.455 147.735 81.330 148.065 ;
        RECT 79.195 147.565 79.420 147.605 ;
        RECT 80.085 147.565 80.285 147.735 ;
        RECT 76.805 146.825 77.075 147.285 ;
        RECT 77.245 146.995 77.530 147.455 ;
        RECT 77.815 146.825 78.105 147.550 ;
        RECT 79.195 147.480 79.575 147.565 ;
        RECT 79.245 147.045 79.575 147.480 ;
        RECT 79.745 146.825 79.915 147.435 ;
        RECT 80.085 147.040 80.415 147.565 ;
        RECT 80.675 146.825 80.885 147.355 ;
        RECT 81.160 147.275 81.330 147.735 ;
        RECT 81.500 147.775 81.820 148.735 ;
        RECT 81.990 147.985 82.180 148.705 ;
        RECT 82.350 147.805 82.520 148.875 ;
        RECT 82.690 148.575 82.860 149.375 ;
        RECT 83.030 148.930 84.135 149.100 ;
        RECT 83.030 148.315 83.200 148.930 ;
        RECT 84.345 148.780 84.595 149.205 ;
        RECT 84.765 148.915 85.030 149.375 ;
        RECT 83.370 148.395 83.900 148.760 ;
        RECT 84.345 148.650 84.650 148.780 ;
        RECT 82.690 148.225 83.200 148.315 ;
        RECT 82.690 148.055 83.560 148.225 ;
        RECT 82.690 147.985 82.860 148.055 ;
        RECT 82.980 147.805 83.180 147.835 ;
        RECT 81.500 147.445 81.965 147.775 ;
        RECT 82.350 147.505 83.180 147.805 ;
        RECT 82.350 147.275 82.520 147.505 ;
        RECT 81.160 147.105 81.945 147.275 ;
        RECT 82.115 147.105 82.520 147.275 ;
        RECT 82.700 146.825 83.070 147.325 ;
        RECT 83.390 147.275 83.560 148.055 ;
        RECT 83.730 147.695 83.900 148.395 ;
        RECT 84.070 147.865 84.310 148.460 ;
        RECT 83.730 147.475 84.255 147.695 ;
        RECT 84.480 147.545 84.650 148.650 ;
        RECT 84.425 147.415 84.650 147.545 ;
        RECT 84.820 147.455 85.100 148.405 ;
        RECT 84.425 147.275 84.595 147.415 ;
        RECT 83.390 147.105 84.065 147.275 ;
        RECT 84.260 147.105 84.595 147.275 ;
        RECT 84.765 146.825 85.015 147.285 ;
        RECT 85.270 147.085 85.455 149.205 ;
        RECT 85.625 148.875 85.955 149.375 ;
        RECT 86.125 148.705 86.295 149.205 ;
        RECT 85.630 148.535 86.295 148.705 ;
        RECT 86.645 148.705 86.815 149.205 ;
        RECT 86.985 148.875 87.315 149.375 ;
        RECT 86.645 148.535 87.310 148.705 ;
        RECT 85.630 147.545 85.860 148.535 ;
        RECT 86.030 147.715 86.380 148.365 ;
        RECT 86.560 147.715 86.910 148.365 ;
        RECT 87.080 147.545 87.310 148.535 ;
        RECT 85.630 147.375 86.295 147.545 ;
        RECT 85.625 146.825 85.955 147.205 ;
        RECT 86.125 147.085 86.295 147.375 ;
        RECT 86.645 147.375 87.310 147.545 ;
        RECT 86.645 147.085 86.815 147.375 ;
        RECT 86.985 146.825 87.315 147.205 ;
        RECT 87.485 147.085 87.670 149.205 ;
        RECT 87.910 148.915 88.175 149.375 ;
        RECT 88.345 148.780 88.595 149.205 ;
        RECT 88.805 148.930 89.910 149.100 ;
        RECT 88.290 148.650 88.595 148.780 ;
        RECT 87.840 147.455 88.120 148.405 ;
        RECT 88.290 147.545 88.460 148.650 ;
        RECT 88.630 147.865 88.870 148.460 ;
        RECT 89.040 148.395 89.570 148.760 ;
        RECT 89.040 147.695 89.210 148.395 ;
        RECT 89.740 148.315 89.910 148.930 ;
        RECT 90.080 148.575 90.250 149.375 ;
        RECT 90.420 148.875 90.670 149.205 ;
        RECT 90.895 148.905 91.780 149.075 ;
        RECT 89.740 148.225 90.250 148.315 ;
        RECT 88.290 147.415 88.515 147.545 ;
        RECT 88.685 147.475 89.210 147.695 ;
        RECT 89.380 148.055 90.250 148.225 ;
        RECT 87.925 146.825 88.175 147.285 ;
        RECT 88.345 147.275 88.515 147.415 ;
        RECT 89.380 147.275 89.550 148.055 ;
        RECT 90.080 147.985 90.250 148.055 ;
        RECT 89.760 147.805 89.960 147.835 ;
        RECT 90.420 147.805 90.590 148.875 ;
        RECT 90.760 147.985 90.950 148.705 ;
        RECT 89.760 147.505 90.590 147.805 ;
        RECT 91.120 147.775 91.440 148.735 ;
        RECT 88.345 147.105 88.680 147.275 ;
        RECT 88.875 147.105 89.550 147.275 ;
        RECT 89.870 146.825 90.240 147.325 ;
        RECT 90.420 147.275 90.590 147.505 ;
        RECT 90.975 147.445 91.440 147.775 ;
        RECT 91.610 148.065 91.780 148.905 ;
        RECT 91.960 148.875 92.275 149.375 ;
        RECT 92.505 148.645 92.845 149.205 ;
        RECT 91.950 148.270 92.845 148.645 ;
        RECT 93.015 148.365 93.185 149.375 ;
        RECT 92.655 148.065 92.845 148.270 ;
        RECT 93.355 148.315 93.685 149.160 ;
        RECT 94.925 148.705 95.095 149.205 ;
        RECT 95.265 148.875 95.595 149.375 ;
        RECT 94.925 148.535 95.590 148.705 ;
        RECT 93.355 148.235 93.745 148.315 ;
        RECT 93.530 148.185 93.745 148.235 ;
        RECT 91.610 147.735 92.485 148.065 ;
        RECT 92.655 147.735 93.405 148.065 ;
        RECT 91.610 147.275 91.780 147.735 ;
        RECT 92.655 147.565 92.855 147.735 ;
        RECT 93.575 147.605 93.745 148.185 ;
        RECT 94.840 147.715 95.190 148.365 ;
        RECT 93.520 147.565 93.745 147.605 ;
        RECT 90.420 147.105 90.825 147.275 ;
        RECT 90.995 147.105 91.780 147.275 ;
        RECT 92.055 146.825 92.265 147.355 ;
        RECT 92.525 147.040 92.855 147.565 ;
        RECT 93.365 147.480 93.745 147.565 ;
        RECT 95.360 147.545 95.590 148.535 ;
        RECT 93.025 146.825 93.195 147.435 ;
        RECT 93.365 147.045 93.695 147.480 ;
        RECT 94.925 147.375 95.590 147.545 ;
        RECT 94.925 147.085 95.095 147.375 ;
        RECT 95.265 146.825 95.595 147.205 ;
        RECT 95.765 147.085 95.950 149.205 ;
        RECT 96.190 148.915 96.455 149.375 ;
        RECT 96.625 148.780 96.875 149.205 ;
        RECT 97.085 148.930 98.190 149.100 ;
        RECT 96.570 148.650 96.875 148.780 ;
        RECT 96.120 147.455 96.400 148.405 ;
        RECT 96.570 147.545 96.740 148.650 ;
        RECT 96.910 147.865 97.150 148.460 ;
        RECT 97.320 148.395 97.850 148.760 ;
        RECT 97.320 147.695 97.490 148.395 ;
        RECT 98.020 148.315 98.190 148.930 ;
        RECT 98.360 148.575 98.530 149.375 ;
        RECT 98.700 148.875 98.950 149.205 ;
        RECT 99.175 148.905 100.060 149.075 ;
        RECT 98.020 148.225 98.530 148.315 ;
        RECT 96.570 147.415 96.795 147.545 ;
        RECT 96.965 147.475 97.490 147.695 ;
        RECT 97.660 148.055 98.530 148.225 ;
        RECT 96.205 146.825 96.455 147.285 ;
        RECT 96.625 147.275 96.795 147.415 ;
        RECT 97.660 147.275 97.830 148.055 ;
        RECT 98.360 147.985 98.530 148.055 ;
        RECT 98.040 147.805 98.240 147.835 ;
        RECT 98.700 147.805 98.870 148.875 ;
        RECT 99.040 147.985 99.230 148.705 ;
        RECT 98.040 147.505 98.870 147.805 ;
        RECT 99.400 147.775 99.720 148.735 ;
        RECT 96.625 147.105 96.960 147.275 ;
        RECT 97.155 147.105 97.830 147.275 ;
        RECT 98.150 146.825 98.520 147.325 ;
        RECT 98.700 147.275 98.870 147.505 ;
        RECT 99.255 147.445 99.720 147.775 ;
        RECT 99.890 148.065 100.060 148.905 ;
        RECT 100.240 148.875 100.555 149.375 ;
        RECT 100.785 148.645 101.125 149.205 ;
        RECT 100.230 148.270 101.125 148.645 ;
        RECT 101.295 148.365 101.465 149.375 ;
        RECT 100.935 148.065 101.125 148.270 ;
        RECT 101.635 148.315 101.965 149.160 ;
        RECT 101.635 148.235 102.025 148.315 ;
        RECT 102.195 148.285 103.405 149.375 ;
        RECT 101.810 148.185 102.025 148.235 ;
        RECT 99.890 147.735 100.765 148.065 ;
        RECT 100.935 147.735 101.685 148.065 ;
        RECT 99.890 147.275 100.060 147.735 ;
        RECT 100.935 147.565 101.135 147.735 ;
        RECT 101.855 147.605 102.025 148.185 ;
        RECT 101.800 147.565 102.025 147.605 ;
        RECT 98.700 147.105 99.105 147.275 ;
        RECT 99.275 147.105 100.060 147.275 ;
        RECT 100.335 146.825 100.545 147.355 ;
        RECT 100.805 147.040 101.135 147.565 ;
        RECT 101.645 147.480 102.025 147.565 ;
        RECT 102.195 147.575 102.715 148.115 ;
        RECT 102.885 147.745 103.405 148.285 ;
        RECT 103.575 148.210 103.865 149.375 ;
        RECT 104.035 148.235 104.420 149.205 ;
        RECT 104.590 148.915 104.915 149.375 ;
        RECT 105.435 148.745 105.715 149.205 ;
        RECT 104.590 148.525 105.715 148.745 ;
        RECT 101.305 146.825 101.475 147.435 ;
        RECT 101.645 147.045 101.975 147.480 ;
        RECT 102.195 146.825 103.405 147.575 ;
        RECT 104.035 147.565 104.315 148.235 ;
        RECT 104.590 148.065 105.040 148.525 ;
        RECT 105.905 148.355 106.305 149.205 ;
        RECT 106.705 148.915 106.975 149.375 ;
        RECT 107.145 148.745 107.430 149.205 ;
        RECT 104.485 147.735 105.040 148.065 ;
        RECT 105.210 147.795 106.305 148.355 ;
        RECT 104.590 147.625 105.040 147.735 ;
        RECT 103.575 146.825 103.865 147.550 ;
        RECT 104.035 146.995 104.420 147.565 ;
        RECT 104.590 147.455 105.715 147.625 ;
        RECT 104.590 146.825 104.915 147.285 ;
        RECT 105.435 146.995 105.715 147.455 ;
        RECT 105.905 146.995 106.305 147.795 ;
        RECT 106.475 148.525 107.430 148.745 ;
        RECT 106.475 147.625 106.685 148.525 ;
        RECT 106.855 147.795 107.545 148.355 ;
        RECT 107.715 148.235 108.100 149.205 ;
        RECT 108.270 148.915 108.595 149.375 ;
        RECT 109.115 148.745 109.395 149.205 ;
        RECT 108.270 148.525 109.395 148.745 ;
        RECT 106.475 147.455 107.430 147.625 ;
        RECT 106.705 146.825 106.975 147.285 ;
        RECT 107.145 146.995 107.430 147.455 ;
        RECT 107.715 147.565 107.995 148.235 ;
        RECT 108.270 148.065 108.720 148.525 ;
        RECT 109.585 148.355 109.985 149.205 ;
        RECT 110.385 148.915 110.655 149.375 ;
        RECT 110.825 148.745 111.110 149.205 ;
        RECT 108.165 147.735 108.720 148.065 ;
        RECT 108.890 147.795 109.985 148.355 ;
        RECT 108.270 147.625 108.720 147.735 ;
        RECT 107.715 146.995 108.100 147.565 ;
        RECT 108.270 147.455 109.395 147.625 ;
        RECT 108.270 146.825 108.595 147.285 ;
        RECT 109.115 146.995 109.395 147.455 ;
        RECT 109.585 146.995 109.985 147.795 ;
        RECT 110.155 148.525 111.110 148.745 ;
        RECT 110.155 147.625 110.365 148.525 ;
        RECT 111.600 148.405 111.930 149.205 ;
        RECT 112.100 148.575 112.430 149.375 ;
        RECT 112.730 148.405 113.060 149.205 ;
        RECT 113.705 148.575 113.955 149.375 ;
        RECT 110.535 147.795 111.225 148.355 ;
        RECT 111.600 148.235 114.035 148.405 ;
        RECT 114.225 148.235 114.395 149.375 ;
        RECT 114.565 148.235 114.905 149.205 ;
        RECT 111.395 147.815 111.745 148.065 ;
        RECT 110.155 147.455 111.110 147.625 ;
        RECT 111.930 147.605 112.100 148.235 ;
        RECT 112.270 147.815 112.600 148.015 ;
        RECT 112.770 147.815 113.100 148.015 ;
        RECT 113.270 147.815 113.690 148.015 ;
        RECT 113.865 147.985 114.035 148.235 ;
        RECT 113.865 147.815 114.560 147.985 ;
        RECT 110.385 146.825 110.655 147.285 ;
        RECT 110.825 146.995 111.110 147.455 ;
        RECT 111.600 146.995 112.100 147.605 ;
        RECT 112.730 147.475 113.955 147.645 ;
        RECT 114.730 147.625 114.905 148.235 ;
        RECT 112.730 146.995 113.060 147.475 ;
        RECT 113.230 146.825 113.455 147.285 ;
        RECT 113.625 146.995 113.955 147.475 ;
        RECT 114.145 146.825 114.395 147.625 ;
        RECT 114.565 146.995 114.905 147.625 ;
        RECT 115.110 148.585 115.645 149.205 ;
        RECT 115.110 147.565 115.425 148.585 ;
        RECT 115.815 148.575 116.145 149.375 ;
        RECT 117.375 148.940 122.720 149.375 ;
        RECT 122.895 148.940 128.240 149.375 ;
        RECT 116.630 148.405 117.020 148.580 ;
        RECT 115.595 148.235 117.020 148.405 ;
        RECT 115.595 147.735 115.765 148.235 ;
        RECT 115.110 146.995 115.725 147.565 ;
        RECT 116.015 147.505 116.280 148.065 ;
        RECT 116.450 147.335 116.620 148.235 ;
        RECT 116.790 147.505 117.145 148.065 ;
        RECT 118.960 147.370 119.300 148.200 ;
        RECT 120.780 147.690 121.130 148.940 ;
        RECT 124.480 147.370 124.820 148.200 ;
        RECT 126.300 147.690 126.650 148.940 ;
        RECT 129.335 148.210 129.625 149.375 ;
        RECT 129.885 148.705 130.055 149.205 ;
        RECT 130.225 148.875 130.555 149.375 ;
        RECT 129.885 148.535 130.550 148.705 ;
        RECT 129.800 147.715 130.150 148.365 ;
        RECT 115.895 146.825 116.110 147.335 ;
        RECT 116.340 147.005 116.620 147.335 ;
        RECT 116.800 146.825 117.040 147.335 ;
        RECT 117.375 146.825 122.720 147.370 ;
        RECT 122.895 146.825 128.240 147.370 ;
        RECT 129.335 146.825 129.625 147.550 ;
        RECT 130.320 147.545 130.550 148.535 ;
        RECT 129.885 147.375 130.550 147.545 ;
        RECT 129.885 147.085 130.055 147.375 ;
        RECT 130.225 146.825 130.555 147.205 ;
        RECT 130.725 147.085 130.910 149.205 ;
        RECT 131.150 148.915 131.415 149.375 ;
        RECT 131.585 148.780 131.835 149.205 ;
        RECT 132.045 148.930 133.150 149.100 ;
        RECT 131.530 148.650 131.835 148.780 ;
        RECT 131.080 147.455 131.360 148.405 ;
        RECT 131.530 147.545 131.700 148.650 ;
        RECT 131.870 147.865 132.110 148.460 ;
        RECT 132.280 148.395 132.810 148.760 ;
        RECT 132.280 147.695 132.450 148.395 ;
        RECT 132.980 148.315 133.150 148.930 ;
        RECT 133.320 148.575 133.490 149.375 ;
        RECT 133.660 148.875 133.910 149.205 ;
        RECT 134.135 148.905 135.020 149.075 ;
        RECT 132.980 148.225 133.490 148.315 ;
        RECT 131.530 147.415 131.755 147.545 ;
        RECT 131.925 147.475 132.450 147.695 ;
        RECT 132.620 148.055 133.490 148.225 ;
        RECT 131.165 146.825 131.415 147.285 ;
        RECT 131.585 147.275 131.755 147.415 ;
        RECT 132.620 147.275 132.790 148.055 ;
        RECT 133.320 147.985 133.490 148.055 ;
        RECT 133.000 147.805 133.200 147.835 ;
        RECT 133.660 147.805 133.830 148.875 ;
        RECT 134.000 147.985 134.190 148.705 ;
        RECT 133.000 147.505 133.830 147.805 ;
        RECT 134.360 147.775 134.680 148.735 ;
        RECT 131.585 147.105 131.920 147.275 ;
        RECT 132.115 147.105 132.790 147.275 ;
        RECT 133.110 146.825 133.480 147.325 ;
        RECT 133.660 147.275 133.830 147.505 ;
        RECT 134.215 147.445 134.680 147.775 ;
        RECT 134.850 148.065 135.020 148.905 ;
        RECT 135.200 148.875 135.515 149.375 ;
        RECT 135.745 148.645 136.085 149.205 ;
        RECT 135.190 148.270 136.085 148.645 ;
        RECT 136.255 148.365 136.425 149.375 ;
        RECT 135.895 148.065 136.085 148.270 ;
        RECT 136.595 148.315 136.925 149.160 ;
        RECT 136.595 148.235 136.985 148.315 ;
        RECT 136.770 148.185 136.985 148.235 ;
        RECT 134.850 147.735 135.725 148.065 ;
        RECT 135.895 147.735 136.645 148.065 ;
        RECT 134.850 147.275 135.020 147.735 ;
        RECT 135.895 147.565 136.095 147.735 ;
        RECT 136.815 147.605 136.985 148.185 ;
        RECT 137.615 148.285 138.825 149.375 ;
        RECT 137.615 147.745 138.135 148.285 ;
        RECT 136.760 147.565 136.985 147.605 ;
        RECT 138.305 147.575 138.825 148.115 ;
        RECT 133.660 147.105 134.065 147.275 ;
        RECT 134.235 147.105 135.020 147.275 ;
        RECT 135.295 146.825 135.505 147.355 ;
        RECT 135.765 147.040 136.095 147.565 ;
        RECT 136.605 147.480 136.985 147.565 ;
        RECT 136.265 146.825 136.435 147.435 ;
        RECT 136.605 147.045 136.935 147.480 ;
        RECT 137.615 146.825 138.825 147.575 ;
        RECT 13.330 146.655 138.910 146.825 ;
        RECT 13.415 145.905 14.625 146.655 ;
        RECT 15.805 146.105 15.975 146.395 ;
        RECT 16.145 146.275 16.475 146.655 ;
        RECT 15.805 145.935 16.470 146.105 ;
        RECT 13.415 145.365 13.935 145.905 ;
        RECT 14.105 145.195 14.625 145.735 ;
        RECT 13.415 144.105 14.625 145.195 ;
        RECT 15.720 145.115 16.070 145.765 ;
        RECT 16.240 144.945 16.470 145.935 ;
        RECT 15.805 144.775 16.470 144.945 ;
        RECT 15.805 144.275 15.975 144.775 ;
        RECT 16.145 144.105 16.475 144.605 ;
        RECT 16.645 144.275 16.830 146.395 ;
        RECT 17.085 146.195 17.335 146.655 ;
        RECT 17.505 146.205 17.840 146.375 ;
        RECT 18.035 146.205 18.710 146.375 ;
        RECT 17.505 146.065 17.675 146.205 ;
        RECT 17.000 145.075 17.280 146.025 ;
        RECT 17.450 145.935 17.675 146.065 ;
        RECT 17.450 144.830 17.620 145.935 ;
        RECT 17.845 145.785 18.370 146.005 ;
        RECT 17.790 145.020 18.030 145.615 ;
        RECT 18.200 145.085 18.370 145.785 ;
        RECT 18.540 145.425 18.710 146.205 ;
        RECT 19.030 146.155 19.400 146.655 ;
        RECT 19.580 146.205 19.985 146.375 ;
        RECT 20.155 146.205 20.940 146.375 ;
        RECT 19.580 145.975 19.750 146.205 ;
        RECT 18.920 145.675 19.750 145.975 ;
        RECT 20.135 145.705 20.600 146.035 ;
        RECT 18.920 145.645 19.120 145.675 ;
        RECT 19.240 145.425 19.410 145.495 ;
        RECT 18.540 145.255 19.410 145.425 ;
        RECT 18.900 145.165 19.410 145.255 ;
        RECT 17.450 144.700 17.755 144.830 ;
        RECT 18.200 144.720 18.730 145.085 ;
        RECT 17.070 144.105 17.335 144.565 ;
        RECT 17.505 144.275 17.755 144.700 ;
        RECT 18.900 144.550 19.070 145.165 ;
        RECT 17.965 144.380 19.070 144.550 ;
        RECT 19.240 144.105 19.410 144.905 ;
        RECT 19.580 144.605 19.750 145.675 ;
        RECT 19.920 144.775 20.110 145.495 ;
        RECT 20.280 144.745 20.600 145.705 ;
        RECT 20.770 145.745 20.940 146.205 ;
        RECT 21.215 146.125 21.425 146.655 ;
        RECT 21.685 145.915 22.015 146.440 ;
        RECT 22.185 146.045 22.355 146.655 ;
        RECT 22.525 146.000 22.855 146.435 ;
        RECT 22.525 145.915 22.905 146.000 ;
        RECT 21.815 145.745 22.015 145.915 ;
        RECT 22.680 145.875 22.905 145.915 ;
        RECT 20.770 145.415 21.645 145.745 ;
        RECT 21.815 145.415 22.565 145.745 ;
        RECT 19.580 144.275 19.830 144.605 ;
        RECT 20.770 144.575 20.940 145.415 ;
        RECT 21.815 145.210 22.005 145.415 ;
        RECT 22.735 145.295 22.905 145.875 ;
        RECT 23.095 145.845 23.335 146.655 ;
        RECT 23.505 145.845 23.835 146.485 ;
        RECT 24.005 145.845 24.275 146.655 ;
        RECT 24.475 145.845 24.715 146.655 ;
        RECT 24.885 145.845 25.215 146.485 ;
        RECT 25.385 145.845 25.655 146.655 ;
        RECT 25.835 146.110 31.180 146.655 ;
        RECT 23.075 145.415 23.425 145.665 ;
        RECT 22.690 145.245 22.905 145.295 ;
        RECT 23.595 145.245 23.765 145.845 ;
        RECT 23.935 145.415 24.285 145.665 ;
        RECT 24.455 145.415 24.805 145.665 ;
        RECT 24.975 145.245 25.145 145.845 ;
        RECT 25.315 145.415 25.665 145.665 ;
        RECT 27.420 145.280 27.760 146.110 ;
        RECT 32.315 145.835 32.545 146.655 ;
        RECT 32.715 145.855 33.045 146.485 ;
        RECT 21.110 144.835 22.005 145.210 ;
        RECT 22.515 145.165 22.905 145.245 ;
        RECT 20.055 144.405 20.940 144.575 ;
        RECT 21.120 144.105 21.435 144.605 ;
        RECT 21.665 144.275 22.005 144.835 ;
        RECT 22.175 144.105 22.345 145.115 ;
        RECT 22.515 144.320 22.845 145.165 ;
        RECT 23.085 145.075 23.765 145.245 ;
        RECT 23.085 144.290 23.415 145.075 ;
        RECT 23.945 144.105 24.275 145.245 ;
        RECT 24.465 145.075 25.145 145.245 ;
        RECT 24.465 144.290 24.795 145.075 ;
        RECT 25.325 144.105 25.655 145.245 ;
        RECT 29.240 144.540 29.590 145.790 ;
        RECT 32.295 145.415 32.625 145.665 ;
        RECT 32.795 145.255 33.045 145.855 ;
        RECT 33.215 145.835 33.425 146.655 ;
        RECT 33.655 145.855 34.350 146.485 ;
        RECT 34.555 145.855 34.865 146.655 ;
        RECT 35.125 146.085 35.295 146.485 ;
        RECT 35.535 146.255 35.865 146.655 ;
        RECT 36.135 146.315 37.540 146.485 ;
        RECT 36.135 146.085 36.305 146.315 ;
        RECT 35.125 145.915 36.305 146.085 ;
        RECT 37.370 146.085 37.540 146.315 ;
        RECT 37.710 146.275 38.040 146.655 ;
        RECT 33.675 145.415 34.010 145.665 ;
        RECT 34.180 145.295 34.350 145.855 ;
        RECT 36.475 145.745 36.665 145.975 ;
        RECT 34.520 145.415 34.855 145.685 ;
        RECT 35.095 145.415 35.280 145.745 ;
        RECT 35.535 145.415 36.010 145.745 ;
        RECT 36.320 145.415 36.665 145.745 ;
        RECT 36.925 145.415 37.120 145.990 ;
        RECT 37.370 145.915 38.065 146.085 ;
        RECT 38.235 146.070 38.545 146.485 ;
        RECT 37.895 145.745 38.065 145.915 ;
        RECT 37.390 145.415 37.725 145.745 ;
        RECT 37.895 145.415 38.205 145.745 ;
        RECT 34.175 145.255 34.350 145.295 ;
        RECT 25.835 144.105 31.180 144.540 ;
        RECT 32.315 144.105 32.545 145.245 ;
        RECT 32.715 144.275 33.045 145.255 ;
        RECT 33.215 144.105 33.425 145.245 ;
        RECT 33.655 144.105 33.915 145.245 ;
        RECT 34.085 144.275 34.415 145.255 ;
        RECT 37.895 145.245 38.065 145.415 ;
        RECT 34.585 144.105 34.865 145.245 ;
        RECT 35.125 145.075 38.065 145.245 ;
        RECT 35.125 144.275 35.295 145.075 ;
        RECT 38.375 144.955 38.545 146.070 ;
        RECT 39.175 145.930 39.465 146.655 ;
        RECT 39.635 146.275 40.525 146.445 ;
        RECT 39.635 145.720 40.185 146.105 ;
        RECT 40.355 145.550 40.525 146.275 ;
        RECT 39.635 145.480 40.525 145.550 ;
        RECT 40.695 145.950 40.915 146.435 ;
        RECT 41.085 146.115 41.335 146.655 ;
        RECT 41.505 146.005 41.765 146.485 ;
        RECT 40.695 145.525 41.025 145.950 ;
        RECT 39.635 145.455 40.530 145.480 ;
        RECT 39.635 145.440 40.540 145.455 ;
        RECT 39.635 145.425 40.545 145.440 ;
        RECT 39.635 145.420 40.555 145.425 ;
        RECT 39.635 145.410 40.560 145.420 ;
        RECT 39.635 145.400 40.565 145.410 ;
        RECT 39.635 145.395 40.575 145.400 ;
        RECT 39.635 145.385 40.585 145.395 ;
        RECT 39.635 145.380 40.595 145.385 ;
        RECT 36.055 144.735 37.615 144.905 ;
        RECT 36.055 144.275 36.305 144.735 ;
        RECT 36.505 144.105 37.175 144.485 ;
        RECT 37.365 144.275 37.615 144.735 ;
        RECT 37.790 144.105 38.035 144.565 ;
        RECT 38.205 144.315 38.545 144.955 ;
        RECT 39.175 144.105 39.465 145.270 ;
        RECT 39.635 144.930 39.895 145.380 ;
        RECT 40.260 145.375 40.595 145.380 ;
        RECT 40.260 145.370 40.610 145.375 ;
        RECT 40.260 145.360 40.625 145.370 ;
        RECT 40.260 145.355 40.650 145.360 ;
        RECT 41.195 145.355 41.425 145.750 ;
        RECT 40.260 145.350 41.425 145.355 ;
        RECT 40.290 145.315 41.425 145.350 ;
        RECT 40.325 145.290 41.425 145.315 ;
        RECT 40.355 145.260 41.425 145.290 ;
        RECT 40.375 145.230 41.425 145.260 ;
        RECT 40.395 145.200 41.425 145.230 ;
        RECT 40.465 145.190 41.425 145.200 ;
        RECT 40.490 145.180 41.425 145.190 ;
        RECT 40.510 145.165 41.425 145.180 ;
        RECT 40.530 145.150 41.425 145.165 ;
        RECT 40.535 145.140 41.320 145.150 ;
        RECT 40.550 145.105 41.320 145.140 ;
        RECT 40.065 144.785 40.395 145.030 ;
        RECT 40.565 144.855 41.320 145.105 ;
        RECT 41.595 144.975 41.765 146.005 ;
        RECT 41.935 145.905 43.145 146.655 ;
        RECT 43.325 146.060 43.575 146.485 ;
        RECT 43.745 146.230 44.075 146.655 ;
        RECT 44.245 146.235 45.335 146.485 ;
        RECT 45.525 146.235 46.615 146.485 ;
        RECT 44.245 146.060 44.415 146.235 ;
        RECT 41.935 145.365 42.455 145.905 ;
        RECT 43.325 145.890 44.415 146.060 ;
        RECT 44.585 145.895 46.275 146.065 ;
        RECT 46.445 146.060 46.615 146.235 ;
        RECT 46.785 146.230 47.115 146.655 ;
        RECT 47.285 146.060 47.605 146.485 ;
        RECT 42.625 145.195 43.145 145.735 ;
        RECT 43.380 145.635 44.010 145.665 ;
        RECT 43.375 145.465 44.010 145.635 ;
        RECT 44.300 145.465 44.930 145.665 ;
        RECT 45.100 145.255 45.390 145.895 ;
        RECT 46.445 145.890 47.605 146.060 ;
        RECT 48.005 145.975 48.175 146.350 ;
        RECT 47.975 145.805 48.175 145.975 ;
        RECT 48.365 146.125 48.595 146.430 ;
        RECT 48.765 146.295 49.095 146.655 ;
        RECT 49.290 146.125 49.580 146.475 ;
        RECT 48.365 145.955 49.580 146.125 ;
        RECT 49.755 145.855 50.450 146.485 ;
        RECT 50.655 145.855 50.965 146.655 ;
        RECT 51.340 145.875 51.840 146.485 ;
        RECT 48.005 145.785 48.175 145.805 ;
        RECT 45.675 145.465 46.330 145.665 ;
        RECT 46.620 145.635 47.730 145.665 ;
        RECT 46.595 145.465 47.730 145.635 ;
        RECT 48.005 145.615 48.525 145.785 ;
        RECT 40.065 144.760 40.250 144.785 ;
        RECT 39.635 144.660 40.250 144.760 ;
        RECT 39.635 144.105 40.240 144.660 ;
        RECT 40.415 144.275 40.895 144.615 ;
        RECT 41.065 144.105 41.320 144.650 ;
        RECT 41.490 144.275 41.765 144.975 ;
        RECT 41.935 144.105 43.145 145.195 ;
        RECT 43.325 145.085 45.390 145.255 ;
        RECT 43.325 144.275 43.575 145.085 ;
        RECT 43.745 144.445 43.995 144.915 ;
        RECT 44.165 144.615 44.495 145.085 ;
        RECT 44.665 144.445 44.835 144.915 ;
        RECT 45.005 144.615 45.390 145.085 ;
        RECT 45.605 145.085 47.535 145.255 ;
        RECT 47.920 145.085 48.165 145.445 ;
        RECT 48.355 145.235 48.525 145.615 ;
        RECT 48.695 145.415 49.080 145.745 ;
        RECT 49.260 145.415 49.520 145.745 ;
        RECT 49.775 145.415 50.110 145.665 ;
        RECT 45.605 144.445 45.855 145.085 ;
        RECT 43.745 144.275 45.855 144.445 ;
        RECT 46.025 144.105 46.195 144.915 ;
        RECT 46.365 144.275 46.695 145.085 ;
        RECT 46.865 144.105 47.035 144.915 ;
        RECT 47.205 144.275 47.535 145.085 ;
        RECT 48.355 144.955 48.705 145.235 ;
        RECT 47.920 144.105 48.175 144.905 ;
        RECT 48.375 144.275 48.705 144.955 ;
        RECT 48.885 144.365 49.080 145.415 ;
        RECT 50.280 145.255 50.450 145.855 ;
        RECT 50.620 145.415 50.955 145.685 ;
        RECT 51.135 145.415 51.485 145.665 ;
        RECT 49.260 144.105 49.580 145.245 ;
        RECT 49.755 144.105 50.015 145.245 ;
        RECT 50.185 144.275 50.515 145.255 ;
        RECT 51.670 145.245 51.840 145.875 ;
        RECT 52.470 146.005 52.800 146.485 ;
        RECT 52.970 146.195 53.195 146.655 ;
        RECT 53.365 146.005 53.695 146.485 ;
        RECT 52.470 145.835 53.695 146.005 ;
        RECT 53.885 145.855 54.135 146.655 ;
        RECT 54.305 145.855 54.645 146.485 ;
        RECT 54.815 146.275 55.705 146.445 ;
        RECT 52.010 145.465 52.340 145.665 ;
        RECT 52.510 145.465 52.840 145.665 ;
        RECT 53.010 145.465 53.430 145.665 ;
        RECT 53.605 145.495 54.300 145.665 ;
        RECT 53.605 145.245 53.775 145.495 ;
        RECT 54.470 145.245 54.645 145.855 ;
        RECT 54.815 145.720 55.365 146.105 ;
        RECT 55.535 145.550 55.705 146.275 ;
        RECT 50.685 144.105 50.965 145.245 ;
        RECT 51.340 145.075 53.775 145.245 ;
        RECT 51.340 144.275 51.670 145.075 ;
        RECT 51.840 144.105 52.170 144.905 ;
        RECT 52.470 144.275 52.800 145.075 ;
        RECT 53.445 144.105 53.695 144.905 ;
        RECT 53.965 144.105 54.135 145.245 ;
        RECT 54.305 144.275 54.645 145.245 ;
        RECT 54.815 145.480 55.705 145.550 ;
        RECT 55.875 145.950 56.095 146.435 ;
        RECT 56.265 146.115 56.515 146.655 ;
        RECT 56.685 146.005 56.945 146.485 ;
        RECT 55.875 145.525 56.205 145.950 ;
        RECT 54.815 145.455 55.710 145.480 ;
        RECT 54.815 145.440 55.720 145.455 ;
        RECT 54.815 145.425 55.725 145.440 ;
        RECT 54.815 145.420 55.735 145.425 ;
        RECT 54.815 145.410 55.740 145.420 ;
        RECT 54.815 145.400 55.745 145.410 ;
        RECT 54.815 145.395 55.755 145.400 ;
        RECT 54.815 145.385 55.765 145.395 ;
        RECT 54.815 145.380 55.775 145.385 ;
        RECT 54.815 144.930 55.075 145.380 ;
        RECT 55.440 145.375 55.775 145.380 ;
        RECT 55.440 145.370 55.790 145.375 ;
        RECT 55.440 145.360 55.805 145.370 ;
        RECT 55.440 145.355 55.830 145.360 ;
        RECT 56.375 145.355 56.605 145.750 ;
        RECT 55.440 145.350 56.605 145.355 ;
        RECT 55.470 145.315 56.605 145.350 ;
        RECT 55.505 145.290 56.605 145.315 ;
        RECT 55.535 145.260 56.605 145.290 ;
        RECT 55.555 145.230 56.605 145.260 ;
        RECT 55.575 145.200 56.605 145.230 ;
        RECT 55.645 145.190 56.605 145.200 ;
        RECT 55.670 145.180 56.605 145.190 ;
        RECT 55.690 145.165 56.605 145.180 ;
        RECT 55.710 145.150 56.605 145.165 ;
        RECT 55.715 145.140 56.500 145.150 ;
        RECT 55.730 145.105 56.500 145.140 ;
        RECT 55.245 144.785 55.575 145.030 ;
        RECT 55.745 144.855 56.500 145.105 ;
        RECT 56.775 144.975 56.945 146.005 ;
        RECT 57.135 145.845 57.375 146.655 ;
        RECT 57.545 145.845 57.875 146.485 ;
        RECT 58.045 145.845 58.315 146.655 ;
        RECT 58.495 146.110 63.840 146.655 ;
        RECT 57.115 145.415 57.465 145.665 ;
        RECT 57.635 145.245 57.805 145.845 ;
        RECT 57.975 145.415 58.325 145.665 ;
        RECT 60.080 145.280 60.420 146.110 ;
        RECT 64.935 145.930 65.225 146.655 ;
        RECT 65.395 145.905 66.605 146.655 ;
        RECT 55.245 144.760 55.430 144.785 ;
        RECT 54.815 144.660 55.430 144.760 ;
        RECT 54.815 144.105 55.420 144.660 ;
        RECT 55.595 144.275 56.075 144.615 ;
        RECT 56.245 144.105 56.500 144.650 ;
        RECT 56.670 144.275 56.945 144.975 ;
        RECT 57.125 145.075 57.805 145.245 ;
        RECT 57.125 144.290 57.455 145.075 ;
        RECT 57.985 144.105 58.315 145.245 ;
        RECT 61.900 144.540 62.250 145.790 ;
        RECT 65.395 145.365 65.915 145.905 ;
        RECT 66.775 145.835 67.035 146.655 ;
        RECT 67.205 145.835 67.535 146.255 ;
        RECT 67.715 146.170 68.505 146.435 ;
        RECT 67.285 145.745 67.535 145.835 ;
        RECT 58.495 144.105 63.840 144.540 ;
        RECT 64.935 144.105 65.225 145.270 ;
        RECT 66.085 145.195 66.605 145.735 ;
        RECT 65.395 144.105 66.605 145.195 ;
        RECT 66.775 144.785 67.115 145.665 ;
        RECT 67.285 145.495 68.080 145.745 ;
        RECT 66.775 144.105 67.035 144.615 ;
        RECT 67.285 144.275 67.455 145.495 ;
        RECT 68.250 145.315 68.505 146.170 ;
        RECT 68.675 146.015 68.875 146.435 ;
        RECT 69.065 146.195 69.395 146.655 ;
        RECT 68.675 145.495 69.085 146.015 ;
        RECT 69.565 146.005 69.825 146.485 ;
        RECT 69.995 146.275 70.885 146.445 ;
        RECT 69.255 145.315 69.485 145.745 ;
        RECT 67.695 145.145 69.485 145.315 ;
        RECT 67.695 144.780 67.945 145.145 ;
        RECT 68.115 144.785 68.445 144.975 ;
        RECT 68.665 144.850 69.380 145.145 ;
        RECT 69.655 144.975 69.825 146.005 ;
        RECT 69.995 145.720 70.545 146.105 ;
        RECT 70.715 145.550 70.885 146.275 ;
        RECT 68.115 144.610 68.310 144.785 ;
        RECT 67.695 144.105 68.310 144.610 ;
        RECT 68.480 144.275 68.955 144.615 ;
        RECT 69.125 144.105 69.340 144.650 ;
        RECT 69.550 144.275 69.825 144.975 ;
        RECT 69.995 145.480 70.885 145.550 ;
        RECT 71.055 145.975 71.275 146.435 ;
        RECT 71.445 146.115 71.695 146.655 ;
        RECT 71.865 146.005 72.125 146.485 ;
        RECT 71.055 145.950 71.305 145.975 ;
        RECT 71.055 145.525 71.385 145.950 ;
        RECT 69.995 145.455 70.890 145.480 ;
        RECT 69.995 145.440 70.900 145.455 ;
        RECT 69.995 145.425 70.905 145.440 ;
        RECT 69.995 145.420 70.915 145.425 ;
        RECT 69.995 145.410 70.920 145.420 ;
        RECT 69.995 145.400 70.925 145.410 ;
        RECT 69.995 145.395 70.935 145.400 ;
        RECT 69.995 145.385 70.945 145.395 ;
        RECT 69.995 145.380 70.955 145.385 ;
        RECT 69.995 144.930 70.255 145.380 ;
        RECT 70.620 145.375 70.955 145.380 ;
        RECT 70.620 145.370 70.970 145.375 ;
        RECT 70.620 145.360 70.985 145.370 ;
        RECT 70.620 145.355 71.010 145.360 ;
        RECT 71.555 145.355 71.785 145.750 ;
        RECT 70.620 145.350 71.785 145.355 ;
        RECT 70.650 145.315 71.785 145.350 ;
        RECT 70.685 145.290 71.785 145.315 ;
        RECT 70.715 145.260 71.785 145.290 ;
        RECT 70.735 145.230 71.785 145.260 ;
        RECT 70.755 145.200 71.785 145.230 ;
        RECT 70.825 145.190 71.785 145.200 ;
        RECT 70.850 145.180 71.785 145.190 ;
        RECT 70.870 145.165 71.785 145.180 ;
        RECT 70.890 145.150 71.785 145.165 ;
        RECT 70.895 145.140 71.680 145.150 ;
        RECT 70.910 145.105 71.680 145.140 ;
        RECT 70.425 144.785 70.755 145.030 ;
        RECT 70.925 144.855 71.680 145.105 ;
        RECT 71.955 144.975 72.125 146.005 ;
        RECT 72.355 145.835 72.565 146.655 ;
        RECT 72.735 145.855 73.065 146.485 ;
        RECT 72.735 145.255 72.985 145.855 ;
        RECT 73.235 145.835 73.465 146.655 ;
        RECT 74.135 146.145 74.440 146.655 ;
        RECT 73.155 145.415 73.485 145.665 ;
        RECT 74.135 145.415 74.450 145.975 ;
        RECT 74.620 145.665 74.870 146.475 ;
        RECT 75.040 146.130 75.300 146.655 ;
        RECT 75.480 145.665 75.730 146.475 ;
        RECT 75.900 146.095 76.160 146.655 ;
        RECT 76.330 146.005 76.590 146.460 ;
        RECT 76.760 146.175 77.020 146.655 ;
        RECT 77.190 146.005 77.450 146.460 ;
        RECT 77.620 146.175 77.880 146.655 ;
        RECT 78.050 146.005 78.310 146.460 ;
        RECT 78.480 146.175 78.725 146.655 ;
        RECT 78.895 146.005 79.170 146.460 ;
        RECT 79.340 146.175 79.585 146.655 ;
        RECT 79.755 146.005 80.015 146.460 ;
        RECT 80.195 146.175 80.445 146.655 ;
        RECT 80.615 146.005 80.875 146.460 ;
        RECT 81.055 146.175 81.305 146.655 ;
        RECT 81.475 146.005 81.735 146.460 ;
        RECT 81.915 146.175 82.175 146.655 ;
        RECT 82.345 146.005 82.605 146.460 ;
        RECT 82.775 146.175 83.075 146.655 ;
        RECT 83.425 146.105 83.595 146.395 ;
        RECT 83.765 146.275 84.095 146.655 ;
        RECT 76.330 145.835 83.075 146.005 ;
        RECT 83.425 145.935 84.090 146.105 ;
        RECT 74.620 145.415 81.740 145.665 ;
        RECT 70.425 144.760 70.610 144.785 ;
        RECT 69.995 144.660 70.610 144.760 ;
        RECT 69.995 144.105 70.600 144.660 ;
        RECT 70.775 144.275 71.255 144.615 ;
        RECT 71.425 144.105 71.680 144.650 ;
        RECT 71.850 144.275 72.125 144.975 ;
        RECT 72.355 144.105 72.565 145.245 ;
        RECT 72.735 144.275 73.065 145.255 ;
        RECT 73.235 144.105 73.465 145.245 ;
        RECT 74.145 144.105 74.440 144.915 ;
        RECT 74.620 144.275 74.865 145.415 ;
        RECT 75.040 144.105 75.300 144.915 ;
        RECT 75.480 144.280 75.730 145.415 ;
        RECT 81.910 145.245 83.075 145.835 ;
        RECT 76.330 145.020 83.075 145.245 ;
        RECT 83.340 145.115 83.690 145.765 ;
        RECT 76.330 145.005 81.735 145.020 ;
        RECT 75.900 144.110 76.160 144.905 ;
        RECT 76.330 144.280 76.590 145.005 ;
        RECT 76.760 144.110 77.020 144.835 ;
        RECT 77.190 144.280 77.450 145.005 ;
        RECT 77.620 144.110 77.880 144.835 ;
        RECT 78.050 144.280 78.310 145.005 ;
        RECT 78.480 144.110 78.740 144.835 ;
        RECT 78.910 144.280 79.170 145.005 ;
        RECT 79.340 144.110 79.585 144.835 ;
        RECT 79.755 144.280 80.015 145.005 ;
        RECT 80.200 144.110 80.445 144.835 ;
        RECT 80.615 144.280 80.875 145.005 ;
        RECT 81.060 144.110 81.305 144.835 ;
        RECT 81.475 144.280 81.735 145.005 ;
        RECT 81.920 144.110 82.175 144.835 ;
        RECT 82.345 144.280 82.635 145.020 ;
        RECT 83.860 144.945 84.090 145.935 ;
        RECT 75.900 144.105 82.175 144.110 ;
        RECT 82.805 144.105 83.075 144.850 ;
        RECT 83.425 144.775 84.090 144.945 ;
        RECT 83.425 144.275 83.595 144.775 ;
        RECT 83.765 144.105 84.095 144.605 ;
        RECT 84.265 144.275 84.450 146.395 ;
        RECT 84.705 146.195 84.955 146.655 ;
        RECT 85.125 146.205 85.460 146.375 ;
        RECT 85.655 146.205 86.330 146.375 ;
        RECT 85.125 146.065 85.295 146.205 ;
        RECT 84.620 145.075 84.900 146.025 ;
        RECT 85.070 145.935 85.295 146.065 ;
        RECT 85.070 144.830 85.240 145.935 ;
        RECT 85.465 145.785 85.990 146.005 ;
        RECT 85.410 145.020 85.650 145.615 ;
        RECT 85.820 145.085 85.990 145.785 ;
        RECT 86.160 145.425 86.330 146.205 ;
        RECT 86.650 146.155 87.020 146.655 ;
        RECT 87.200 146.205 87.605 146.375 ;
        RECT 87.775 146.205 88.560 146.375 ;
        RECT 87.200 145.975 87.370 146.205 ;
        RECT 86.540 145.675 87.370 145.975 ;
        RECT 87.755 145.705 88.220 146.035 ;
        RECT 86.540 145.645 86.740 145.675 ;
        RECT 86.860 145.425 87.030 145.495 ;
        RECT 86.160 145.255 87.030 145.425 ;
        RECT 86.520 145.165 87.030 145.255 ;
        RECT 85.070 144.700 85.375 144.830 ;
        RECT 85.820 144.720 86.350 145.085 ;
        RECT 84.690 144.105 84.955 144.565 ;
        RECT 85.125 144.275 85.375 144.700 ;
        RECT 86.520 144.550 86.690 145.165 ;
        RECT 85.585 144.380 86.690 144.550 ;
        RECT 86.860 144.105 87.030 144.905 ;
        RECT 87.200 144.605 87.370 145.675 ;
        RECT 87.540 144.775 87.730 145.495 ;
        RECT 87.900 144.745 88.220 145.705 ;
        RECT 88.390 145.745 88.560 146.205 ;
        RECT 88.835 146.125 89.045 146.655 ;
        RECT 89.305 145.915 89.635 146.440 ;
        RECT 89.805 146.045 89.975 146.655 ;
        RECT 90.145 146.000 90.475 146.435 ;
        RECT 90.145 145.915 90.525 146.000 ;
        RECT 90.695 145.930 90.985 146.655 ;
        RECT 89.435 145.745 89.635 145.915 ;
        RECT 90.300 145.875 90.525 145.915 ;
        RECT 88.390 145.415 89.265 145.745 ;
        RECT 89.435 145.415 90.185 145.745 ;
        RECT 87.200 144.275 87.450 144.605 ;
        RECT 88.390 144.575 88.560 145.415 ;
        RECT 89.435 145.210 89.625 145.415 ;
        RECT 90.355 145.295 90.525 145.875 ;
        RECT 91.155 145.885 92.825 146.655 ;
        RECT 93.545 146.105 93.715 146.395 ;
        RECT 93.885 146.275 94.215 146.655 ;
        RECT 93.545 145.935 94.210 146.105 ;
        RECT 91.155 145.365 91.905 145.885 ;
        RECT 90.310 145.245 90.525 145.295 ;
        RECT 88.730 144.835 89.625 145.210 ;
        RECT 90.135 145.165 90.525 145.245 ;
        RECT 87.675 144.405 88.560 144.575 ;
        RECT 88.740 144.105 89.055 144.605 ;
        RECT 89.285 144.275 89.625 144.835 ;
        RECT 89.795 144.105 89.965 145.115 ;
        RECT 90.135 144.320 90.465 145.165 ;
        RECT 90.695 144.105 90.985 145.270 ;
        RECT 92.075 145.195 92.825 145.715 ;
        RECT 91.155 144.105 92.825 145.195 ;
        RECT 93.460 145.115 93.810 145.765 ;
        RECT 93.980 144.945 94.210 145.935 ;
        RECT 93.545 144.775 94.210 144.945 ;
        RECT 93.545 144.275 93.715 144.775 ;
        RECT 93.885 144.105 94.215 144.605 ;
        RECT 94.385 144.275 94.570 146.395 ;
        RECT 94.825 146.195 95.075 146.655 ;
        RECT 95.245 146.205 95.580 146.375 ;
        RECT 95.775 146.205 96.450 146.375 ;
        RECT 95.245 146.065 95.415 146.205 ;
        RECT 94.740 145.075 95.020 146.025 ;
        RECT 95.190 145.935 95.415 146.065 ;
        RECT 95.190 144.830 95.360 145.935 ;
        RECT 95.585 145.785 96.110 146.005 ;
        RECT 95.530 145.020 95.770 145.615 ;
        RECT 95.940 145.085 96.110 145.785 ;
        RECT 96.280 145.425 96.450 146.205 ;
        RECT 96.770 146.155 97.140 146.655 ;
        RECT 97.320 146.205 97.725 146.375 ;
        RECT 97.895 146.205 98.680 146.375 ;
        RECT 97.320 145.975 97.490 146.205 ;
        RECT 96.660 145.675 97.490 145.975 ;
        RECT 97.875 145.705 98.340 146.035 ;
        RECT 96.660 145.645 96.860 145.675 ;
        RECT 96.980 145.425 97.150 145.495 ;
        RECT 96.280 145.255 97.150 145.425 ;
        RECT 96.640 145.165 97.150 145.255 ;
        RECT 95.190 144.700 95.495 144.830 ;
        RECT 95.940 144.720 96.470 145.085 ;
        RECT 94.810 144.105 95.075 144.565 ;
        RECT 95.245 144.275 95.495 144.700 ;
        RECT 96.640 144.550 96.810 145.165 ;
        RECT 95.705 144.380 96.810 144.550 ;
        RECT 96.980 144.105 97.150 144.905 ;
        RECT 97.320 144.605 97.490 145.675 ;
        RECT 97.660 144.775 97.850 145.495 ;
        RECT 98.020 144.745 98.340 145.705 ;
        RECT 98.510 145.745 98.680 146.205 ;
        RECT 98.955 146.125 99.165 146.655 ;
        RECT 99.425 145.915 99.755 146.440 ;
        RECT 99.925 146.045 100.095 146.655 ;
        RECT 100.265 146.000 100.595 146.435 ;
        RECT 100.265 145.915 100.645 146.000 ;
        RECT 99.555 145.745 99.755 145.915 ;
        RECT 100.420 145.875 100.645 145.915 ;
        RECT 98.510 145.415 99.385 145.745 ;
        RECT 99.555 145.415 100.305 145.745 ;
        RECT 97.320 144.275 97.570 144.605 ;
        RECT 98.510 144.575 98.680 145.415 ;
        RECT 99.555 145.210 99.745 145.415 ;
        RECT 100.475 145.295 100.645 145.875 ;
        RECT 100.430 145.245 100.645 145.295 ;
        RECT 98.850 144.835 99.745 145.210 ;
        RECT 100.255 145.165 100.645 145.245 ;
        RECT 100.820 145.915 101.075 146.485 ;
        RECT 101.245 146.255 101.575 146.655 ;
        RECT 102.000 146.120 102.530 146.485 ;
        RECT 102.720 146.315 102.995 146.485 ;
        RECT 102.715 146.145 102.995 146.315 ;
        RECT 102.000 146.085 102.175 146.120 ;
        RECT 101.245 145.915 102.175 146.085 ;
        RECT 100.820 145.245 100.990 145.915 ;
        RECT 101.245 145.745 101.415 145.915 ;
        RECT 101.160 145.415 101.415 145.745 ;
        RECT 101.640 145.415 101.835 145.745 ;
        RECT 97.795 144.405 98.680 144.575 ;
        RECT 98.860 144.105 99.175 144.605 ;
        RECT 99.405 144.275 99.745 144.835 ;
        RECT 99.915 144.105 100.085 145.115 ;
        RECT 100.255 144.320 100.585 145.165 ;
        RECT 100.820 144.275 101.155 145.245 ;
        RECT 101.325 144.105 101.495 145.245 ;
        RECT 101.665 144.445 101.835 145.415 ;
        RECT 102.005 144.785 102.175 145.915 ;
        RECT 102.345 145.125 102.515 145.925 ;
        RECT 102.720 145.325 102.995 146.145 ;
        RECT 103.165 145.125 103.355 146.485 ;
        RECT 103.535 146.120 104.045 146.655 ;
        RECT 104.265 145.845 104.510 146.450 ;
        RECT 104.960 145.915 105.215 146.485 ;
        RECT 105.385 146.255 105.715 146.655 ;
        RECT 106.140 146.120 106.670 146.485 ;
        RECT 106.860 146.315 107.135 146.485 ;
        RECT 106.855 146.145 107.135 146.315 ;
        RECT 106.140 146.085 106.315 146.120 ;
        RECT 105.385 145.915 106.315 146.085 ;
        RECT 103.555 145.675 104.785 145.845 ;
        RECT 102.345 144.955 103.355 145.125 ;
        RECT 103.525 145.110 104.275 145.300 ;
        RECT 102.005 144.615 103.130 144.785 ;
        RECT 103.525 144.445 103.695 145.110 ;
        RECT 104.445 144.865 104.785 145.675 ;
        RECT 101.665 144.275 103.695 144.445 ;
        RECT 103.865 144.105 104.035 144.865 ;
        RECT 104.270 144.455 104.785 144.865 ;
        RECT 104.960 145.245 105.130 145.915 ;
        RECT 105.385 145.745 105.555 145.915 ;
        RECT 105.300 145.415 105.555 145.745 ;
        RECT 105.780 145.415 105.975 145.745 ;
        RECT 104.960 144.275 105.295 145.245 ;
        RECT 105.465 144.105 105.635 145.245 ;
        RECT 105.805 144.445 105.975 145.415 ;
        RECT 106.145 144.785 106.315 145.915 ;
        RECT 106.485 145.125 106.655 145.925 ;
        RECT 106.860 145.325 107.135 146.145 ;
        RECT 107.305 145.125 107.495 146.485 ;
        RECT 107.675 146.120 108.185 146.655 ;
        RECT 108.405 145.845 108.650 146.450 ;
        RECT 109.185 146.105 109.355 146.395 ;
        RECT 109.525 146.275 109.855 146.655 ;
        RECT 109.185 145.935 109.850 146.105 ;
        RECT 107.695 145.675 108.925 145.845 ;
        RECT 106.485 144.955 107.495 145.125 ;
        RECT 107.665 145.110 108.415 145.300 ;
        RECT 106.145 144.615 107.270 144.785 ;
        RECT 107.665 144.445 107.835 145.110 ;
        RECT 108.585 144.865 108.925 145.675 ;
        RECT 109.100 145.115 109.450 145.765 ;
        RECT 109.620 144.945 109.850 145.935 ;
        RECT 105.805 144.275 107.835 144.445 ;
        RECT 108.005 144.105 108.175 144.865 ;
        RECT 108.410 144.455 108.925 144.865 ;
        RECT 109.185 144.775 109.850 144.945 ;
        RECT 109.185 144.275 109.355 144.775 ;
        RECT 109.525 144.105 109.855 144.605 ;
        RECT 110.025 144.275 110.210 146.395 ;
        RECT 110.465 146.195 110.715 146.655 ;
        RECT 110.885 146.205 111.220 146.375 ;
        RECT 111.415 146.205 112.090 146.375 ;
        RECT 110.885 146.065 111.055 146.205 ;
        RECT 110.380 145.075 110.660 146.025 ;
        RECT 110.830 145.935 111.055 146.065 ;
        RECT 110.830 144.830 111.000 145.935 ;
        RECT 111.225 145.785 111.750 146.005 ;
        RECT 111.170 145.020 111.410 145.615 ;
        RECT 111.580 145.085 111.750 145.785 ;
        RECT 111.920 145.425 112.090 146.205 ;
        RECT 112.410 146.155 112.780 146.655 ;
        RECT 112.960 146.205 113.365 146.375 ;
        RECT 113.535 146.205 114.320 146.375 ;
        RECT 112.960 145.975 113.130 146.205 ;
        RECT 112.300 145.675 113.130 145.975 ;
        RECT 113.515 145.705 113.980 146.035 ;
        RECT 112.300 145.645 112.500 145.675 ;
        RECT 112.620 145.425 112.790 145.495 ;
        RECT 111.920 145.255 112.790 145.425 ;
        RECT 112.280 145.165 112.790 145.255 ;
        RECT 110.830 144.700 111.135 144.830 ;
        RECT 111.580 144.720 112.110 145.085 ;
        RECT 110.450 144.105 110.715 144.565 ;
        RECT 110.885 144.275 111.135 144.700 ;
        RECT 112.280 144.550 112.450 145.165 ;
        RECT 111.345 144.380 112.450 144.550 ;
        RECT 112.620 144.105 112.790 144.905 ;
        RECT 112.960 144.605 113.130 145.675 ;
        RECT 113.300 144.775 113.490 145.495 ;
        RECT 113.660 144.745 113.980 145.705 ;
        RECT 114.150 145.745 114.320 146.205 ;
        RECT 114.595 146.125 114.805 146.655 ;
        RECT 115.065 145.915 115.395 146.440 ;
        RECT 115.565 146.045 115.735 146.655 ;
        RECT 115.905 146.000 116.235 146.435 ;
        RECT 115.905 145.915 116.285 146.000 ;
        RECT 116.455 145.930 116.745 146.655 ;
        RECT 117.005 146.105 117.175 146.395 ;
        RECT 117.345 146.275 117.675 146.655 ;
        RECT 117.005 145.935 117.670 146.105 ;
        RECT 115.195 145.745 115.395 145.915 ;
        RECT 116.060 145.875 116.285 145.915 ;
        RECT 114.150 145.415 115.025 145.745 ;
        RECT 115.195 145.415 115.945 145.745 ;
        RECT 112.960 144.275 113.210 144.605 ;
        RECT 114.150 144.575 114.320 145.415 ;
        RECT 115.195 145.210 115.385 145.415 ;
        RECT 116.115 145.295 116.285 145.875 ;
        RECT 116.070 145.245 116.285 145.295 ;
        RECT 114.490 144.835 115.385 145.210 ;
        RECT 115.895 145.165 116.285 145.245 ;
        RECT 113.435 144.405 114.320 144.575 ;
        RECT 114.500 144.105 114.815 144.605 ;
        RECT 115.045 144.275 115.385 144.835 ;
        RECT 115.555 144.105 115.725 145.115 ;
        RECT 115.895 144.320 116.225 145.165 ;
        RECT 116.455 144.105 116.745 145.270 ;
        RECT 116.920 145.115 117.270 145.765 ;
        RECT 117.440 144.945 117.670 145.935 ;
        RECT 117.005 144.775 117.670 144.945 ;
        RECT 117.005 144.275 117.175 144.775 ;
        RECT 117.345 144.105 117.675 144.605 ;
        RECT 117.845 144.275 118.030 146.395 ;
        RECT 118.285 146.195 118.535 146.655 ;
        RECT 118.705 146.205 119.040 146.375 ;
        RECT 119.235 146.205 119.910 146.375 ;
        RECT 118.705 146.065 118.875 146.205 ;
        RECT 118.200 145.075 118.480 146.025 ;
        RECT 118.650 145.935 118.875 146.065 ;
        RECT 118.650 144.830 118.820 145.935 ;
        RECT 119.045 145.785 119.570 146.005 ;
        RECT 118.990 145.020 119.230 145.615 ;
        RECT 119.400 145.085 119.570 145.785 ;
        RECT 119.740 145.425 119.910 146.205 ;
        RECT 120.230 146.155 120.600 146.655 ;
        RECT 120.780 146.205 121.185 146.375 ;
        RECT 121.355 146.205 122.140 146.375 ;
        RECT 120.780 145.975 120.950 146.205 ;
        RECT 120.120 145.675 120.950 145.975 ;
        RECT 121.335 145.705 121.800 146.035 ;
        RECT 120.120 145.645 120.320 145.675 ;
        RECT 120.440 145.425 120.610 145.495 ;
        RECT 119.740 145.255 120.610 145.425 ;
        RECT 120.100 145.165 120.610 145.255 ;
        RECT 118.650 144.700 118.955 144.830 ;
        RECT 119.400 144.720 119.930 145.085 ;
        RECT 118.270 144.105 118.535 144.565 ;
        RECT 118.705 144.275 118.955 144.700 ;
        RECT 120.100 144.550 120.270 145.165 ;
        RECT 119.165 144.380 120.270 144.550 ;
        RECT 120.440 144.105 120.610 144.905 ;
        RECT 120.780 144.605 120.950 145.675 ;
        RECT 121.120 144.775 121.310 145.495 ;
        RECT 121.480 144.745 121.800 145.705 ;
        RECT 121.970 145.745 122.140 146.205 ;
        RECT 122.415 146.125 122.625 146.655 ;
        RECT 122.885 145.915 123.215 146.440 ;
        RECT 123.385 146.045 123.555 146.655 ;
        RECT 123.725 146.000 124.055 146.435 ;
        RECT 123.725 145.915 124.105 146.000 ;
        RECT 123.015 145.745 123.215 145.915 ;
        RECT 123.880 145.875 124.105 145.915 ;
        RECT 121.970 145.415 122.845 145.745 ;
        RECT 123.015 145.415 123.765 145.745 ;
        RECT 120.780 144.275 121.030 144.605 ;
        RECT 121.970 144.575 122.140 145.415 ;
        RECT 123.015 145.210 123.205 145.415 ;
        RECT 123.935 145.295 124.105 145.875 ;
        RECT 124.275 145.885 125.945 146.655 ;
        RECT 124.275 145.365 125.025 145.885 ;
        RECT 126.320 145.875 126.820 146.485 ;
        RECT 123.890 145.245 124.105 145.295 ;
        RECT 122.310 144.835 123.205 145.210 ;
        RECT 123.715 145.165 124.105 145.245 ;
        RECT 125.195 145.195 125.945 145.715 ;
        RECT 126.115 145.415 126.465 145.665 ;
        RECT 126.650 145.245 126.820 145.875 ;
        RECT 127.450 146.005 127.780 146.485 ;
        RECT 127.950 146.195 128.175 146.655 ;
        RECT 128.345 146.005 128.675 146.485 ;
        RECT 127.450 145.835 128.675 146.005 ;
        RECT 128.865 145.855 129.115 146.655 ;
        RECT 129.285 145.855 129.625 146.485 ;
        RECT 129.960 146.145 130.200 146.655 ;
        RECT 130.380 146.145 130.660 146.475 ;
        RECT 130.890 146.145 131.105 146.655 ;
        RECT 126.990 145.465 127.320 145.665 ;
        RECT 127.490 145.465 127.820 145.665 ;
        RECT 127.990 145.465 128.410 145.665 ;
        RECT 128.585 145.495 129.280 145.665 ;
        RECT 128.585 145.245 128.755 145.495 ;
        RECT 129.450 145.245 129.625 145.855 ;
        RECT 129.855 145.415 130.210 145.975 ;
        RECT 130.380 145.245 130.550 146.145 ;
        RECT 130.720 145.415 130.985 145.975 ;
        RECT 131.275 145.915 131.890 146.485 ;
        RECT 131.235 145.245 131.405 145.745 ;
        RECT 121.255 144.405 122.140 144.575 ;
        RECT 122.320 144.105 122.635 144.605 ;
        RECT 122.865 144.275 123.205 144.835 ;
        RECT 123.375 144.105 123.545 145.115 ;
        RECT 123.715 144.320 124.045 145.165 ;
        RECT 124.275 144.105 125.945 145.195 ;
        RECT 126.320 145.075 128.755 145.245 ;
        RECT 126.320 144.275 126.650 145.075 ;
        RECT 126.820 144.105 127.150 144.905 ;
        RECT 127.450 144.275 127.780 145.075 ;
        RECT 128.425 144.105 128.675 144.905 ;
        RECT 128.945 144.105 129.115 145.245 ;
        RECT 129.285 144.275 129.625 145.245 ;
        RECT 129.980 145.075 131.405 145.245 ;
        RECT 129.980 144.900 130.370 145.075 ;
        RECT 130.855 144.105 131.185 144.905 ;
        RECT 131.575 144.895 131.890 145.915 ;
        RECT 132.095 145.885 133.765 146.655 ;
        RECT 134.025 146.105 134.195 146.485 ;
        RECT 134.410 146.275 134.740 146.655 ;
        RECT 134.025 145.935 134.740 146.105 ;
        RECT 132.095 145.365 132.845 145.885 ;
        RECT 133.015 145.195 133.765 145.715 ;
        RECT 133.935 145.385 134.290 145.755 ;
        RECT 134.570 145.745 134.740 145.935 ;
        RECT 134.910 145.910 135.165 146.485 ;
        RECT 134.570 145.415 134.825 145.745 ;
        RECT 134.570 145.205 134.740 145.415 ;
        RECT 131.355 144.275 131.890 144.895 ;
        RECT 132.095 144.105 133.765 145.195 ;
        RECT 134.025 145.035 134.740 145.205 ;
        RECT 134.995 145.180 135.165 145.910 ;
        RECT 135.340 145.815 135.600 146.655 ;
        RECT 135.865 146.105 136.035 146.485 ;
        RECT 136.250 146.275 136.580 146.655 ;
        RECT 135.865 145.935 136.580 146.105 ;
        RECT 135.775 145.385 136.130 145.755 ;
        RECT 136.410 145.745 136.580 145.935 ;
        RECT 136.750 145.910 137.005 146.485 ;
        RECT 136.410 145.415 136.665 145.745 ;
        RECT 134.025 144.275 134.195 145.035 ;
        RECT 134.410 144.105 134.740 144.865 ;
        RECT 134.910 144.275 135.165 145.180 ;
        RECT 135.340 144.105 135.600 145.255 ;
        RECT 136.410 145.205 136.580 145.415 ;
        RECT 135.865 145.035 136.580 145.205 ;
        RECT 136.835 145.180 137.005 145.910 ;
        RECT 137.180 145.815 137.440 146.655 ;
        RECT 137.615 145.905 138.825 146.655 ;
        RECT 135.865 144.275 136.035 145.035 ;
        RECT 136.250 144.105 136.580 144.865 ;
        RECT 136.750 144.275 137.005 145.180 ;
        RECT 137.180 144.105 137.440 145.255 ;
        RECT 137.615 145.195 138.135 145.735 ;
        RECT 138.305 145.365 138.825 145.905 ;
        RECT 137.615 144.105 138.825 145.195 ;
        RECT 13.330 143.935 138.910 144.105 ;
        RECT 13.415 142.845 14.625 143.935 ;
        RECT 14.795 142.845 18.305 143.935 ;
        RECT 13.415 142.135 13.935 142.675 ;
        RECT 14.105 142.305 14.625 142.845 ;
        RECT 14.795 142.155 16.445 142.675 ;
        RECT 16.615 142.325 18.305 142.845 ;
        RECT 18.475 143.065 18.750 143.765 ;
        RECT 18.920 143.390 19.175 143.935 ;
        RECT 19.345 143.425 19.825 143.765 ;
        RECT 20.000 143.380 20.605 143.935 ;
        RECT 20.775 143.500 26.120 143.935 ;
        RECT 19.990 143.280 20.605 143.380 ;
        RECT 19.990 143.255 20.175 143.280 ;
        RECT 13.415 141.385 14.625 142.135 ;
        RECT 14.795 141.385 18.305 142.155 ;
        RECT 18.475 142.035 18.645 143.065 ;
        RECT 18.920 142.935 19.675 143.185 ;
        RECT 19.845 143.010 20.175 143.255 ;
        RECT 18.920 142.900 19.690 142.935 ;
        RECT 18.920 142.890 19.705 142.900 ;
        RECT 18.815 142.875 19.710 142.890 ;
        RECT 18.815 142.860 19.730 142.875 ;
        RECT 18.815 142.850 19.750 142.860 ;
        RECT 18.815 142.840 19.775 142.850 ;
        RECT 18.815 142.810 19.845 142.840 ;
        RECT 18.815 142.780 19.865 142.810 ;
        RECT 18.815 142.750 19.885 142.780 ;
        RECT 18.815 142.725 19.915 142.750 ;
        RECT 18.815 142.690 19.950 142.725 ;
        RECT 18.815 142.685 19.980 142.690 ;
        RECT 18.815 142.290 19.045 142.685 ;
        RECT 19.590 142.680 19.980 142.685 ;
        RECT 19.615 142.670 19.980 142.680 ;
        RECT 19.630 142.665 19.980 142.670 ;
        RECT 19.645 142.660 19.980 142.665 ;
        RECT 20.345 142.660 20.605 143.110 ;
        RECT 19.645 142.655 20.605 142.660 ;
        RECT 19.655 142.645 20.605 142.655 ;
        RECT 19.665 142.640 20.605 142.645 ;
        RECT 19.675 142.630 20.605 142.640 ;
        RECT 19.680 142.620 20.605 142.630 ;
        RECT 19.685 142.615 20.605 142.620 ;
        RECT 19.695 142.600 20.605 142.615 ;
        RECT 19.700 142.585 20.605 142.600 ;
        RECT 19.710 142.560 20.605 142.585 ;
        RECT 19.215 142.090 19.545 142.515 ;
        RECT 18.475 141.555 18.735 142.035 ;
        RECT 18.905 141.385 19.155 141.925 ;
        RECT 19.325 141.605 19.545 142.090 ;
        RECT 19.715 142.490 20.605 142.560 ;
        RECT 19.715 141.765 19.885 142.490 ;
        RECT 20.055 141.935 20.605 142.320 ;
        RECT 22.360 141.930 22.700 142.760 ;
        RECT 24.180 142.250 24.530 143.500 ;
        RECT 26.295 142.770 26.585 143.935 ;
        RECT 26.755 143.500 32.100 143.935 ;
        RECT 19.715 141.595 20.605 141.765 ;
        RECT 20.775 141.385 26.120 141.930 ;
        RECT 26.295 141.385 26.585 142.110 ;
        RECT 28.340 141.930 28.680 142.760 ;
        RECT 30.160 142.250 30.510 143.500 ;
        RECT 32.275 142.845 33.485 143.935 ;
        RECT 32.275 142.135 32.795 142.675 ;
        RECT 32.965 142.305 33.485 142.845 ;
        RECT 33.655 142.370 34.005 143.765 ;
        RECT 34.175 143.135 34.580 143.935 ;
        RECT 34.750 143.595 36.285 143.765 ;
        RECT 34.750 142.965 34.920 143.595 ;
        RECT 34.175 142.795 34.920 142.965 ;
        RECT 26.755 141.385 32.100 141.930 ;
        RECT 32.275 141.385 33.485 142.135 ;
        RECT 33.655 141.555 33.925 142.370 ;
        RECT 34.175 142.295 34.345 142.795 ;
        RECT 35.090 142.625 35.360 143.370 ;
        RECT 34.515 142.295 34.850 142.625 ;
        RECT 35.020 142.295 35.360 142.625 ;
        RECT 35.550 142.625 35.785 143.370 ;
        RECT 35.955 142.965 36.285 143.595 ;
        RECT 36.470 143.135 36.705 143.935 ;
        RECT 36.875 142.965 37.165 143.765 ;
        RECT 37.535 143.265 37.815 143.935 ;
        RECT 37.985 143.045 38.285 143.595 ;
        RECT 38.485 143.215 38.815 143.935 ;
        RECT 39.005 143.215 39.465 143.765 ;
        RECT 35.955 142.795 37.165 142.965 ;
        RECT 35.550 142.295 35.840 142.625 ;
        RECT 36.010 142.295 36.410 142.625 ;
        RECT 36.580 142.125 36.750 142.795 ;
        RECT 37.350 142.625 37.615 142.985 ;
        RECT 37.985 142.875 38.925 143.045 ;
        RECT 38.755 142.625 38.925 142.875 ;
        RECT 36.920 142.295 37.165 142.625 ;
        RECT 37.350 142.375 38.025 142.625 ;
        RECT 38.245 142.375 38.585 142.625 ;
        RECT 38.755 142.295 39.045 142.625 ;
        RECT 38.755 142.205 38.925 142.295 ;
        RECT 34.095 141.385 34.765 142.125 ;
        RECT 34.935 141.955 36.330 142.125 ;
        RECT 34.935 141.610 35.230 141.955 ;
        RECT 35.410 141.385 35.785 141.785 ;
        RECT 36.000 141.610 36.330 141.955 ;
        RECT 36.580 141.555 37.165 142.125 ;
        RECT 37.535 142.015 38.925 142.205 ;
        RECT 37.535 141.655 37.865 142.015 ;
        RECT 39.215 141.845 39.465 143.215 ;
        RECT 39.635 142.845 42.225 143.935 ;
        RECT 38.485 141.385 38.735 141.845 ;
        RECT 38.905 141.555 39.465 141.845 ;
        RECT 39.635 142.155 40.845 142.675 ;
        RECT 41.015 142.325 42.225 142.845 ;
        RECT 42.395 142.795 42.665 143.765 ;
        RECT 42.875 143.135 43.155 143.935 ;
        RECT 43.325 143.425 44.980 143.715 ;
        RECT 43.390 143.085 44.980 143.255 ;
        RECT 43.390 142.965 43.560 143.085 ;
        RECT 42.835 142.795 43.560 142.965 ;
        RECT 39.635 141.385 42.225 142.155 ;
        RECT 42.395 142.060 42.565 142.795 ;
        RECT 42.835 142.625 43.005 142.795 ;
        RECT 42.735 142.295 43.005 142.625 ;
        RECT 43.175 142.295 43.580 142.625 ;
        RECT 43.750 142.295 44.460 142.915 ;
        RECT 44.660 142.795 44.980 143.085 ;
        RECT 45.155 142.795 45.415 143.765 ;
        RECT 45.610 143.525 45.940 143.935 ;
        RECT 46.140 143.345 46.310 143.765 ;
        RECT 46.525 143.525 47.195 143.935 ;
        RECT 47.430 143.345 47.600 143.765 ;
        RECT 47.905 143.495 48.235 143.935 ;
        RECT 45.585 143.175 47.600 143.345 ;
        RECT 48.405 143.315 48.580 143.765 ;
        RECT 42.835 142.125 43.005 142.295 ;
        RECT 42.395 141.715 42.665 142.060 ;
        RECT 42.835 141.955 44.445 142.125 ;
        RECT 44.630 142.055 44.980 142.625 ;
        RECT 45.155 142.105 45.325 142.795 ;
        RECT 45.585 142.625 45.755 143.175 ;
        RECT 45.495 142.295 45.755 142.625 ;
        RECT 42.855 141.385 43.235 141.785 ;
        RECT 43.405 141.605 43.575 141.955 ;
        RECT 43.745 141.385 44.075 141.785 ;
        RECT 44.275 141.605 44.445 141.955 ;
        RECT 44.645 141.385 44.975 141.885 ;
        RECT 45.155 141.640 45.495 142.105 ;
        RECT 45.925 141.965 46.265 142.995 ;
        RECT 46.455 142.575 46.725 142.995 ;
        RECT 46.455 142.405 46.765 142.575 ;
        RECT 45.160 141.595 45.495 141.640 ;
        RECT 45.665 141.385 45.995 141.765 ;
        RECT 46.455 141.720 46.725 142.405 ;
        RECT 46.950 141.720 47.230 142.995 ;
        RECT 47.430 141.885 47.600 143.175 ;
        RECT 47.950 143.145 48.580 143.315 ;
        RECT 47.950 142.625 48.120 143.145 ;
        RECT 47.770 142.295 48.120 142.625 ;
        RECT 48.300 142.295 48.665 142.975 ;
        RECT 47.950 142.125 48.120 142.295 ;
        RECT 47.950 141.955 48.580 142.125 ;
        RECT 47.430 141.555 47.660 141.885 ;
        RECT 47.905 141.385 48.235 141.765 ;
        RECT 48.405 141.555 48.580 141.955 ;
        RECT 48.835 141.665 49.115 143.765 ;
        RECT 49.305 143.175 50.090 143.935 ;
        RECT 50.485 143.105 50.870 143.765 ;
        RECT 50.485 143.005 50.895 143.105 ;
        RECT 49.285 142.795 50.895 143.005 ;
        RECT 51.195 142.915 51.395 143.705 ;
        RECT 49.285 142.195 49.560 142.795 ;
        RECT 51.065 142.745 51.395 142.915 ;
        RECT 51.565 142.755 51.885 143.935 ;
        RECT 52.055 142.770 52.345 143.935 ;
        RECT 52.525 143.325 52.855 143.755 ;
        RECT 53.035 143.495 53.230 143.935 ;
        RECT 53.400 143.325 53.730 143.755 ;
        RECT 52.525 143.155 53.730 143.325 ;
        RECT 52.525 142.825 53.420 143.155 ;
        RECT 53.900 142.985 54.175 143.755 ;
        RECT 54.355 143.500 59.700 143.935 ;
        RECT 59.875 143.500 65.220 143.935 ;
        RECT 53.590 142.795 54.175 142.985 ;
        RECT 51.065 142.625 51.245 142.745 ;
        RECT 49.730 142.375 50.085 142.625 ;
        RECT 50.280 142.575 50.745 142.625 ;
        RECT 50.275 142.405 50.745 142.575 ;
        RECT 50.280 142.375 50.745 142.405 ;
        RECT 50.915 142.375 51.245 142.625 ;
        RECT 51.420 142.375 51.885 142.575 ;
        RECT 52.530 142.295 52.825 142.625 ;
        RECT 53.005 142.295 53.420 142.625 ;
        RECT 49.285 142.015 50.535 142.195 ;
        RECT 50.170 141.945 50.535 142.015 ;
        RECT 50.705 141.995 51.885 142.165 ;
        RECT 49.345 141.385 49.515 141.845 ;
        RECT 50.705 141.775 51.035 141.995 ;
        RECT 49.785 141.595 51.035 141.775 ;
        RECT 51.205 141.385 51.375 141.825 ;
        RECT 51.545 141.580 51.885 141.995 ;
        RECT 52.055 141.385 52.345 142.110 ;
        RECT 52.525 141.385 52.825 142.115 ;
        RECT 53.005 141.675 53.235 142.295 ;
        RECT 53.590 142.125 53.765 142.795 ;
        RECT 53.435 141.945 53.765 142.125 ;
        RECT 53.935 141.975 54.175 142.625 ;
        RECT 53.435 141.565 53.660 141.945 ;
        RECT 55.940 141.930 56.280 142.760 ;
        RECT 57.760 142.250 58.110 143.500 ;
        RECT 61.460 141.930 61.800 142.760 ;
        RECT 63.280 142.250 63.630 143.500 ;
        RECT 65.395 142.845 67.985 143.935 ;
        RECT 65.395 142.155 66.605 142.675 ;
        RECT 66.775 142.325 67.985 142.845 ;
        RECT 68.155 143.215 68.615 143.765 ;
        RECT 68.805 143.215 69.135 143.935 ;
        RECT 53.830 141.385 54.160 141.775 ;
        RECT 54.355 141.385 59.700 141.930 ;
        RECT 59.875 141.385 65.220 141.930 ;
        RECT 65.395 141.385 67.985 142.155 ;
        RECT 68.155 141.845 68.405 143.215 ;
        RECT 69.335 143.045 69.635 143.595 ;
        RECT 69.805 143.265 70.085 143.935 ;
        RECT 68.695 142.875 69.635 143.045 ;
        RECT 68.695 142.625 68.865 142.875 ;
        RECT 70.005 142.625 70.270 142.985 ;
        RECT 70.455 142.845 73.045 143.935 ;
        RECT 68.575 142.295 68.865 142.625 ;
        RECT 69.035 142.375 69.375 142.625 ;
        RECT 69.595 142.375 70.270 142.625 ;
        RECT 68.695 142.205 68.865 142.295 ;
        RECT 68.695 142.015 70.085 142.205 ;
        RECT 68.155 141.555 68.715 141.845 ;
        RECT 68.885 141.385 69.135 141.845 ;
        RECT 69.755 141.655 70.085 142.015 ;
        RECT 70.455 142.155 71.665 142.675 ;
        RECT 71.835 142.325 73.045 142.845 ;
        RECT 73.675 143.175 74.190 143.585 ;
        RECT 74.425 143.175 74.595 143.935 ;
        RECT 74.765 143.595 76.795 143.765 ;
        RECT 73.675 142.365 74.015 143.175 ;
        RECT 74.765 142.930 74.935 143.595 ;
        RECT 75.330 143.255 76.455 143.425 ;
        RECT 74.185 142.740 74.935 142.930 ;
        RECT 75.105 142.915 76.115 143.085 ;
        RECT 73.675 142.195 74.905 142.365 ;
        RECT 70.455 141.385 73.045 142.155 ;
        RECT 73.950 141.590 74.195 142.195 ;
        RECT 74.415 141.385 74.925 141.920 ;
        RECT 75.105 141.555 75.295 142.915 ;
        RECT 75.465 142.575 75.740 142.715 ;
        RECT 75.465 142.405 75.745 142.575 ;
        RECT 75.465 141.555 75.740 142.405 ;
        RECT 75.945 142.115 76.115 142.915 ;
        RECT 76.285 142.125 76.455 143.255 ;
        RECT 76.625 142.625 76.795 143.595 ;
        RECT 76.965 142.795 77.135 143.935 ;
        RECT 77.305 142.795 77.640 143.765 ;
        RECT 76.625 142.295 76.820 142.625 ;
        RECT 77.045 142.295 77.300 142.625 ;
        RECT 77.045 142.125 77.215 142.295 ;
        RECT 77.470 142.125 77.640 142.795 ;
        RECT 77.815 142.770 78.105 143.935 ;
        RECT 78.275 142.845 81.785 143.935 ;
        RECT 76.285 141.955 77.215 142.125 ;
        RECT 76.285 141.920 76.460 141.955 ;
        RECT 75.930 141.555 76.460 141.920 ;
        RECT 76.885 141.385 77.215 141.785 ;
        RECT 77.385 141.555 77.640 142.125 ;
        RECT 78.275 142.155 79.925 142.675 ;
        RECT 80.095 142.325 81.785 142.845 ;
        RECT 81.955 143.175 82.470 143.585 ;
        RECT 82.705 143.175 82.875 143.935 ;
        RECT 83.045 143.595 85.075 143.765 ;
        RECT 81.955 142.365 82.295 143.175 ;
        RECT 83.045 142.930 83.215 143.595 ;
        RECT 83.610 143.255 84.735 143.425 ;
        RECT 82.465 142.740 83.215 142.930 ;
        RECT 83.385 142.915 84.395 143.085 ;
        RECT 81.955 142.195 83.185 142.365 ;
        RECT 77.815 141.385 78.105 142.110 ;
        RECT 78.275 141.385 81.785 142.155 ;
        RECT 82.230 141.590 82.475 142.195 ;
        RECT 82.695 141.385 83.205 141.920 ;
        RECT 83.385 141.555 83.575 142.915 ;
        RECT 83.745 141.895 84.020 142.715 ;
        RECT 84.225 142.115 84.395 142.915 ;
        RECT 84.565 142.125 84.735 143.255 ;
        RECT 84.905 142.625 85.075 143.595 ;
        RECT 85.245 142.795 85.415 143.935 ;
        RECT 85.585 142.795 85.920 143.765 ;
        RECT 84.905 142.295 85.100 142.625 ;
        RECT 85.325 142.295 85.580 142.625 ;
        RECT 85.325 142.125 85.495 142.295 ;
        RECT 85.750 142.125 85.920 142.795 ;
        RECT 84.565 141.955 85.495 142.125 ;
        RECT 84.565 141.920 84.740 141.955 ;
        RECT 83.745 141.725 84.025 141.895 ;
        RECT 83.745 141.555 84.020 141.725 ;
        RECT 84.210 141.555 84.740 141.920 ;
        RECT 85.165 141.385 85.495 141.785 ;
        RECT 85.665 141.555 85.920 142.125 ;
        RECT 86.095 142.795 86.480 143.765 ;
        RECT 86.650 143.475 86.975 143.935 ;
        RECT 87.495 143.305 87.775 143.765 ;
        RECT 86.650 143.085 87.775 143.305 ;
        RECT 86.095 142.125 86.375 142.795 ;
        RECT 86.650 142.625 87.100 143.085 ;
        RECT 87.965 142.915 88.365 143.765 ;
        RECT 88.765 143.475 89.035 143.935 ;
        RECT 89.205 143.305 89.490 143.765 ;
        RECT 86.545 142.295 87.100 142.625 ;
        RECT 87.270 142.355 88.365 142.915 ;
        RECT 86.650 142.185 87.100 142.295 ;
        RECT 86.095 141.555 86.480 142.125 ;
        RECT 86.650 142.015 87.775 142.185 ;
        RECT 86.650 141.385 86.975 141.845 ;
        RECT 87.495 141.555 87.775 142.015 ;
        RECT 87.965 141.555 88.365 142.355 ;
        RECT 88.535 143.085 89.490 143.305 ;
        RECT 88.535 142.185 88.745 143.085 ;
        RECT 88.915 142.355 89.605 142.915 ;
        RECT 89.775 142.845 93.285 143.935 ;
        RECT 93.545 143.265 93.715 143.765 ;
        RECT 93.885 143.435 94.215 143.935 ;
        RECT 93.545 143.095 94.210 143.265 ;
        RECT 88.535 142.015 89.490 142.185 ;
        RECT 88.765 141.385 89.035 141.845 ;
        RECT 89.205 141.555 89.490 142.015 ;
        RECT 89.775 142.155 91.425 142.675 ;
        RECT 91.595 142.325 93.285 142.845 ;
        RECT 93.460 142.275 93.810 142.925 ;
        RECT 89.775 141.385 93.285 142.155 ;
        RECT 93.980 142.105 94.210 143.095 ;
        RECT 93.545 141.935 94.210 142.105 ;
        RECT 93.545 141.645 93.715 141.935 ;
        RECT 93.885 141.385 94.215 141.765 ;
        RECT 94.385 141.645 94.570 143.765 ;
        RECT 94.810 143.475 95.075 143.935 ;
        RECT 95.245 143.340 95.495 143.765 ;
        RECT 95.705 143.490 96.810 143.660 ;
        RECT 95.190 143.210 95.495 143.340 ;
        RECT 94.740 142.015 95.020 142.965 ;
        RECT 95.190 142.105 95.360 143.210 ;
        RECT 95.530 142.425 95.770 143.020 ;
        RECT 95.940 142.955 96.470 143.320 ;
        RECT 95.940 142.255 96.110 142.955 ;
        RECT 96.640 142.875 96.810 143.490 ;
        RECT 96.980 143.135 97.150 143.935 ;
        RECT 97.320 143.435 97.570 143.765 ;
        RECT 97.795 143.465 98.680 143.635 ;
        RECT 96.640 142.785 97.150 142.875 ;
        RECT 95.190 141.975 95.415 142.105 ;
        RECT 95.585 142.035 96.110 142.255 ;
        RECT 96.280 142.615 97.150 142.785 ;
        RECT 94.825 141.385 95.075 141.845 ;
        RECT 95.245 141.835 95.415 141.975 ;
        RECT 96.280 141.835 96.450 142.615 ;
        RECT 96.980 142.545 97.150 142.615 ;
        RECT 96.660 142.365 96.860 142.395 ;
        RECT 97.320 142.365 97.490 143.435 ;
        RECT 97.660 142.545 97.850 143.265 ;
        RECT 96.660 142.065 97.490 142.365 ;
        RECT 98.020 142.335 98.340 143.295 ;
        RECT 95.245 141.665 95.580 141.835 ;
        RECT 95.775 141.665 96.450 141.835 ;
        RECT 96.770 141.385 97.140 141.885 ;
        RECT 97.320 141.835 97.490 142.065 ;
        RECT 97.875 142.005 98.340 142.335 ;
        RECT 98.510 142.625 98.680 143.465 ;
        RECT 98.860 143.435 99.175 143.935 ;
        RECT 99.405 143.205 99.745 143.765 ;
        RECT 98.850 142.830 99.745 143.205 ;
        RECT 99.915 142.925 100.085 143.935 ;
        RECT 99.555 142.625 99.745 142.830 ;
        RECT 100.255 142.875 100.585 143.720 ;
        RECT 100.255 142.795 100.645 142.875 ;
        RECT 100.815 142.845 103.405 143.935 ;
        RECT 100.430 142.745 100.645 142.795 ;
        RECT 98.510 142.295 99.385 142.625 ;
        RECT 99.555 142.295 100.305 142.625 ;
        RECT 98.510 141.835 98.680 142.295 ;
        RECT 99.555 142.125 99.755 142.295 ;
        RECT 100.475 142.165 100.645 142.745 ;
        RECT 100.420 142.125 100.645 142.165 ;
        RECT 97.320 141.665 97.725 141.835 ;
        RECT 97.895 141.665 98.680 141.835 ;
        RECT 98.955 141.385 99.165 141.915 ;
        RECT 99.425 141.600 99.755 142.125 ;
        RECT 100.265 142.040 100.645 142.125 ;
        RECT 100.815 142.155 102.025 142.675 ;
        RECT 102.195 142.325 103.405 142.845 ;
        RECT 103.575 142.770 103.865 143.935 ;
        RECT 104.035 142.795 104.420 143.765 ;
        RECT 104.590 143.475 104.915 143.935 ;
        RECT 105.435 143.305 105.715 143.765 ;
        RECT 104.590 143.085 105.715 143.305 ;
        RECT 99.925 141.385 100.095 141.995 ;
        RECT 100.265 141.605 100.595 142.040 ;
        RECT 100.815 141.385 103.405 142.155 ;
        RECT 104.035 142.125 104.315 142.795 ;
        RECT 104.590 142.625 105.040 143.085 ;
        RECT 105.905 142.915 106.305 143.765 ;
        RECT 106.705 143.475 106.975 143.935 ;
        RECT 107.145 143.305 107.430 143.765 ;
        RECT 104.485 142.295 105.040 142.625 ;
        RECT 105.210 142.355 106.305 142.915 ;
        RECT 104.590 142.185 105.040 142.295 ;
        RECT 103.575 141.385 103.865 142.110 ;
        RECT 104.035 141.555 104.420 142.125 ;
        RECT 104.590 142.015 105.715 142.185 ;
        RECT 104.590 141.385 104.915 141.845 ;
        RECT 105.435 141.555 105.715 142.015 ;
        RECT 105.905 141.555 106.305 142.355 ;
        RECT 106.475 143.085 107.430 143.305 ;
        RECT 106.475 142.185 106.685 143.085 ;
        RECT 106.855 142.355 107.545 142.915 ;
        RECT 108.635 142.795 108.975 143.765 ;
        RECT 109.145 142.795 109.315 143.935 ;
        RECT 109.585 143.135 109.835 143.935 ;
        RECT 110.480 142.965 110.810 143.765 ;
        RECT 111.110 143.135 111.440 143.935 ;
        RECT 111.610 142.965 111.940 143.765 ;
        RECT 112.405 143.265 112.575 143.765 ;
        RECT 112.745 143.435 113.075 143.935 ;
        RECT 112.405 143.095 113.070 143.265 ;
        RECT 109.505 142.795 111.940 142.965 ;
        RECT 108.635 142.185 108.810 142.795 ;
        RECT 109.505 142.545 109.675 142.795 ;
        RECT 108.980 142.375 109.675 142.545 ;
        RECT 109.850 142.375 110.270 142.575 ;
        RECT 110.440 142.375 110.770 142.575 ;
        RECT 110.940 142.375 111.270 142.575 ;
        RECT 106.475 142.015 107.430 142.185 ;
        RECT 106.705 141.385 106.975 141.845 ;
        RECT 107.145 141.555 107.430 142.015 ;
        RECT 108.635 141.555 108.975 142.185 ;
        RECT 109.145 141.385 109.395 142.185 ;
        RECT 109.585 142.035 110.810 142.205 ;
        RECT 109.585 141.555 109.915 142.035 ;
        RECT 110.085 141.385 110.310 141.845 ;
        RECT 110.480 141.555 110.810 142.035 ;
        RECT 111.440 142.165 111.610 142.795 ;
        RECT 111.795 142.375 112.145 142.625 ;
        RECT 112.320 142.275 112.670 142.925 ;
        RECT 111.440 141.555 111.940 142.165 ;
        RECT 112.840 142.105 113.070 143.095 ;
        RECT 112.405 141.935 113.070 142.105 ;
        RECT 112.405 141.645 112.575 141.935 ;
        RECT 112.745 141.385 113.075 141.765 ;
        RECT 113.245 141.645 113.430 143.765 ;
        RECT 113.670 143.475 113.935 143.935 ;
        RECT 114.105 143.340 114.355 143.765 ;
        RECT 114.565 143.490 115.670 143.660 ;
        RECT 114.050 143.210 114.355 143.340 ;
        RECT 113.600 142.015 113.880 142.965 ;
        RECT 114.050 142.105 114.220 143.210 ;
        RECT 114.390 142.425 114.630 143.020 ;
        RECT 114.800 142.955 115.330 143.320 ;
        RECT 114.800 142.255 114.970 142.955 ;
        RECT 115.500 142.875 115.670 143.490 ;
        RECT 115.840 143.135 116.010 143.935 ;
        RECT 116.180 143.435 116.430 143.765 ;
        RECT 116.655 143.465 117.540 143.635 ;
        RECT 115.500 142.785 116.010 142.875 ;
        RECT 114.050 141.975 114.275 142.105 ;
        RECT 114.445 142.035 114.970 142.255 ;
        RECT 115.140 142.615 116.010 142.785 ;
        RECT 113.685 141.385 113.935 141.845 ;
        RECT 114.105 141.835 114.275 141.975 ;
        RECT 115.140 141.835 115.310 142.615 ;
        RECT 115.840 142.545 116.010 142.615 ;
        RECT 115.520 142.365 115.720 142.395 ;
        RECT 116.180 142.365 116.350 143.435 ;
        RECT 116.520 142.545 116.710 143.265 ;
        RECT 115.520 142.065 116.350 142.365 ;
        RECT 116.880 142.335 117.200 143.295 ;
        RECT 114.105 141.665 114.440 141.835 ;
        RECT 114.635 141.665 115.310 141.835 ;
        RECT 115.630 141.385 116.000 141.885 ;
        RECT 116.180 141.835 116.350 142.065 ;
        RECT 116.735 142.005 117.200 142.335 ;
        RECT 117.370 142.625 117.540 143.465 ;
        RECT 117.720 143.435 118.035 143.935 ;
        RECT 118.265 143.205 118.605 143.765 ;
        RECT 117.710 142.830 118.605 143.205 ;
        RECT 118.775 142.925 118.945 143.935 ;
        RECT 118.415 142.625 118.605 142.830 ;
        RECT 119.115 142.875 119.445 143.720 ;
        RECT 119.860 142.965 120.250 143.140 ;
        RECT 120.735 143.135 121.065 143.935 ;
        RECT 121.235 143.145 121.770 143.765 ;
        RECT 119.115 142.795 119.505 142.875 ;
        RECT 119.860 142.795 121.285 142.965 ;
        RECT 119.290 142.745 119.505 142.795 ;
        RECT 117.370 142.295 118.245 142.625 ;
        RECT 118.415 142.295 119.165 142.625 ;
        RECT 117.370 141.835 117.540 142.295 ;
        RECT 118.415 142.125 118.615 142.295 ;
        RECT 119.335 142.165 119.505 142.745 ;
        RECT 119.280 142.125 119.505 142.165 ;
        RECT 116.180 141.665 116.585 141.835 ;
        RECT 116.755 141.665 117.540 141.835 ;
        RECT 117.815 141.385 118.025 141.915 ;
        RECT 118.285 141.600 118.615 142.125 ;
        RECT 119.125 142.040 119.505 142.125 ;
        RECT 119.735 142.065 120.090 142.625 ;
        RECT 118.785 141.385 118.955 141.995 ;
        RECT 119.125 141.605 119.455 142.040 ;
        RECT 120.260 141.895 120.430 142.795 ;
        RECT 120.600 142.065 120.865 142.625 ;
        RECT 121.115 142.295 121.285 142.795 ;
        RECT 121.455 142.125 121.770 143.145 ;
        RECT 121.975 142.845 123.185 143.935 ;
        RECT 119.840 141.385 120.080 141.895 ;
        RECT 120.260 141.565 120.540 141.895 ;
        RECT 120.770 141.385 120.985 141.895 ;
        RECT 121.155 141.555 121.770 142.125 ;
        RECT 121.975 142.135 122.495 142.675 ;
        RECT 122.665 142.305 123.185 142.845 ;
        RECT 123.540 142.965 123.930 143.140 ;
        RECT 124.415 143.135 124.745 143.935 ;
        RECT 124.915 143.145 125.450 143.765 ;
        RECT 123.540 142.795 124.965 142.965 ;
        RECT 121.975 141.385 123.185 142.135 ;
        RECT 123.415 142.065 123.770 142.625 ;
        RECT 123.940 141.895 124.110 142.795 ;
        RECT 124.280 142.065 124.545 142.625 ;
        RECT 124.795 142.295 124.965 142.795 ;
        RECT 125.135 142.125 125.450 143.145 ;
        RECT 125.860 142.965 126.190 143.765 ;
        RECT 126.360 143.135 126.690 143.935 ;
        RECT 126.990 142.965 127.320 143.765 ;
        RECT 127.965 143.135 128.215 143.935 ;
        RECT 125.860 142.795 128.295 142.965 ;
        RECT 128.485 142.795 128.655 143.935 ;
        RECT 128.825 142.795 129.165 143.765 ;
        RECT 125.655 142.375 126.005 142.625 ;
        RECT 126.190 142.165 126.360 142.795 ;
        RECT 126.530 142.375 126.860 142.575 ;
        RECT 127.030 142.375 127.360 142.575 ;
        RECT 127.530 142.375 127.950 142.575 ;
        RECT 128.125 142.545 128.295 142.795 ;
        RECT 128.125 142.375 128.820 142.545 ;
        RECT 128.990 142.235 129.165 142.795 ;
        RECT 129.335 142.770 129.625 143.935 ;
        RECT 129.885 143.265 130.055 143.765 ;
        RECT 130.225 143.435 130.555 143.935 ;
        RECT 129.885 143.095 130.550 143.265 ;
        RECT 129.800 142.275 130.150 142.925 ;
        RECT 123.520 141.385 123.760 141.895 ;
        RECT 123.940 141.565 124.220 141.895 ;
        RECT 124.450 141.385 124.665 141.895 ;
        RECT 124.835 141.555 125.450 142.125 ;
        RECT 125.860 141.555 126.360 142.165 ;
        RECT 126.990 142.035 128.215 142.205 ;
        RECT 128.935 142.185 129.165 142.235 ;
        RECT 126.990 141.555 127.320 142.035 ;
        RECT 127.490 141.385 127.715 141.845 ;
        RECT 127.885 141.555 128.215 142.035 ;
        RECT 128.405 141.385 128.655 142.185 ;
        RECT 128.825 141.555 129.165 142.185 ;
        RECT 129.335 141.385 129.625 142.110 ;
        RECT 130.320 142.105 130.550 143.095 ;
        RECT 129.885 141.935 130.550 142.105 ;
        RECT 129.885 141.645 130.055 141.935 ;
        RECT 130.225 141.385 130.555 141.765 ;
        RECT 130.725 141.645 130.910 143.765 ;
        RECT 131.150 143.475 131.415 143.935 ;
        RECT 131.585 143.340 131.835 143.765 ;
        RECT 132.045 143.490 133.150 143.660 ;
        RECT 131.530 143.210 131.835 143.340 ;
        RECT 131.080 142.015 131.360 142.965 ;
        RECT 131.530 142.105 131.700 143.210 ;
        RECT 131.870 142.425 132.110 143.020 ;
        RECT 132.280 142.955 132.810 143.320 ;
        RECT 132.280 142.255 132.450 142.955 ;
        RECT 132.980 142.875 133.150 143.490 ;
        RECT 133.320 143.135 133.490 143.935 ;
        RECT 133.660 143.435 133.910 143.765 ;
        RECT 134.135 143.465 135.020 143.635 ;
        RECT 132.980 142.785 133.490 142.875 ;
        RECT 131.530 141.975 131.755 142.105 ;
        RECT 131.925 142.035 132.450 142.255 ;
        RECT 132.620 142.615 133.490 142.785 ;
        RECT 131.165 141.385 131.415 141.845 ;
        RECT 131.585 141.835 131.755 141.975 ;
        RECT 132.620 141.835 132.790 142.615 ;
        RECT 133.320 142.545 133.490 142.615 ;
        RECT 133.000 142.365 133.200 142.395 ;
        RECT 133.660 142.365 133.830 143.435 ;
        RECT 134.000 142.545 134.190 143.265 ;
        RECT 133.000 142.065 133.830 142.365 ;
        RECT 134.360 142.335 134.680 143.295 ;
        RECT 131.585 141.665 131.920 141.835 ;
        RECT 132.115 141.665 132.790 141.835 ;
        RECT 133.110 141.385 133.480 141.885 ;
        RECT 133.660 141.835 133.830 142.065 ;
        RECT 134.215 142.005 134.680 142.335 ;
        RECT 134.850 142.625 135.020 143.465 ;
        RECT 135.200 143.435 135.515 143.935 ;
        RECT 135.745 143.205 136.085 143.765 ;
        RECT 135.190 142.830 136.085 143.205 ;
        RECT 136.255 142.925 136.425 143.935 ;
        RECT 135.895 142.625 136.085 142.830 ;
        RECT 136.595 142.875 136.925 143.720 ;
        RECT 136.595 142.795 136.985 142.875 ;
        RECT 136.770 142.745 136.985 142.795 ;
        RECT 134.850 142.295 135.725 142.625 ;
        RECT 135.895 142.295 136.645 142.625 ;
        RECT 134.850 141.835 135.020 142.295 ;
        RECT 135.895 142.125 136.095 142.295 ;
        RECT 136.815 142.165 136.985 142.745 ;
        RECT 137.615 142.845 138.825 143.935 ;
        RECT 137.615 142.305 138.135 142.845 ;
        RECT 136.760 142.125 136.985 142.165 ;
        RECT 138.305 142.135 138.825 142.675 ;
        RECT 133.660 141.665 134.065 141.835 ;
        RECT 134.235 141.665 135.020 141.835 ;
        RECT 135.295 141.385 135.505 141.915 ;
        RECT 135.765 141.600 136.095 142.125 ;
        RECT 136.605 142.040 136.985 142.125 ;
        RECT 136.265 141.385 136.435 141.995 ;
        RECT 136.605 141.605 136.935 142.040 ;
        RECT 137.615 141.385 138.825 142.135 ;
        RECT 13.330 141.215 138.910 141.385 ;
        RECT 13.415 140.465 14.625 141.215 ;
        RECT 14.795 140.670 20.140 141.215 ;
        RECT 13.415 139.925 13.935 140.465 ;
        RECT 14.105 139.755 14.625 140.295 ;
        RECT 16.380 139.840 16.720 140.670 ;
        RECT 20.315 140.445 21.985 141.215 ;
        RECT 13.415 138.665 14.625 139.755 ;
        RECT 18.200 139.100 18.550 140.350 ;
        RECT 20.315 139.925 21.065 140.445 ;
        RECT 22.165 140.405 22.435 141.215 ;
        RECT 22.605 140.405 22.935 141.045 ;
        RECT 23.105 140.405 23.345 141.215 ;
        RECT 23.535 140.670 28.880 141.215 ;
        RECT 21.235 139.755 21.985 140.275 ;
        RECT 22.155 139.975 22.505 140.225 ;
        RECT 22.675 139.805 22.845 140.405 ;
        RECT 23.015 139.975 23.365 140.225 ;
        RECT 25.120 139.840 25.460 140.670 ;
        RECT 29.055 140.445 32.565 141.215 ;
        RECT 33.285 140.875 33.455 140.910 ;
        RECT 33.255 140.705 33.455 140.875 ;
        RECT 14.795 138.665 20.140 139.100 ;
        RECT 20.315 138.665 21.985 139.755 ;
        RECT 22.165 138.665 22.495 139.805 ;
        RECT 22.675 139.635 23.355 139.805 ;
        RECT 23.025 138.850 23.355 139.635 ;
        RECT 26.940 139.100 27.290 140.350 ;
        RECT 29.055 139.925 30.705 140.445 ;
        RECT 33.285 140.345 33.455 140.705 ;
        RECT 33.645 140.685 33.875 140.990 ;
        RECT 34.045 140.855 34.375 141.215 ;
        RECT 34.570 140.685 34.860 141.035 ;
        RECT 33.645 140.515 34.860 140.685 ;
        RECT 35.045 140.485 35.345 141.215 ;
        RECT 30.875 139.755 32.565 140.275 ;
        RECT 33.285 140.175 33.805 140.345 ;
        RECT 35.525 140.305 35.755 140.925 ;
        RECT 35.955 140.655 36.180 141.035 ;
        RECT 36.350 140.825 36.680 141.215 ;
        RECT 35.955 140.475 36.285 140.655 ;
        RECT 23.535 138.665 28.880 139.100 ;
        RECT 29.055 138.665 32.565 139.755 ;
        RECT 33.200 139.645 33.445 140.005 ;
        RECT 33.635 139.795 33.805 140.175 ;
        RECT 33.975 139.975 34.360 140.305 ;
        RECT 34.540 140.195 34.800 140.305 ;
        RECT 34.540 140.025 34.805 140.195 ;
        RECT 34.540 139.975 34.800 140.025 ;
        RECT 35.050 139.975 35.345 140.305 ;
        RECT 35.525 139.975 35.940 140.305 ;
        RECT 33.635 139.515 33.985 139.795 ;
        RECT 33.200 138.665 33.455 139.465 ;
        RECT 33.655 138.835 33.985 139.515 ;
        RECT 34.165 138.925 34.360 139.975 ;
        RECT 36.110 139.805 36.285 140.475 ;
        RECT 36.455 139.975 36.695 140.625 ;
        RECT 36.875 140.445 38.545 141.215 ;
        RECT 39.175 140.490 39.465 141.215 ;
        RECT 39.635 140.670 44.980 141.215 ;
        RECT 46.240 140.705 46.480 141.215 ;
        RECT 46.660 140.705 46.940 141.035 ;
        RECT 47.170 140.705 47.385 141.215 ;
        RECT 36.875 139.925 37.625 140.445 ;
        RECT 34.540 138.665 34.860 139.805 ;
        RECT 35.045 139.445 35.940 139.775 ;
        RECT 36.110 139.615 36.695 139.805 ;
        RECT 37.795 139.755 38.545 140.275 ;
        RECT 41.220 139.840 41.560 140.670 ;
        RECT 35.045 139.275 36.250 139.445 ;
        RECT 35.045 138.845 35.375 139.275 ;
        RECT 35.555 138.665 35.750 139.105 ;
        RECT 35.920 138.845 36.250 139.275 ;
        RECT 36.420 138.845 36.695 139.615 ;
        RECT 36.875 138.665 38.545 139.755 ;
        RECT 39.175 138.665 39.465 139.830 ;
        RECT 43.040 139.100 43.390 140.350 ;
        RECT 46.135 139.975 46.490 140.535 ;
        RECT 46.660 139.805 46.830 140.705 ;
        RECT 47.000 139.975 47.265 140.535 ;
        RECT 47.555 140.475 48.170 141.045 ;
        RECT 47.515 139.805 47.685 140.305 ;
        RECT 46.260 139.635 47.685 139.805 ;
        RECT 46.260 139.460 46.650 139.635 ;
        RECT 39.635 138.665 44.980 139.100 ;
        RECT 47.135 138.665 47.465 139.465 ;
        RECT 47.855 139.455 48.170 140.475 ;
        RECT 47.635 138.835 48.170 139.455 ;
        RECT 48.410 140.475 49.025 141.045 ;
        RECT 49.195 140.705 49.410 141.215 ;
        RECT 49.640 140.705 49.920 141.035 ;
        RECT 50.100 140.705 50.340 141.215 ;
        RECT 51.595 140.835 52.485 141.005 ;
        RECT 48.410 139.455 48.725 140.475 ;
        RECT 48.895 139.805 49.065 140.305 ;
        RECT 49.315 139.975 49.580 140.535 ;
        RECT 49.750 139.805 49.920 140.705 ;
        RECT 50.090 139.975 50.445 140.535 ;
        RECT 51.595 140.280 52.145 140.665 ;
        RECT 52.315 140.110 52.485 140.835 ;
        RECT 51.595 140.040 52.485 140.110 ;
        RECT 52.655 140.510 52.875 140.995 ;
        RECT 53.045 140.675 53.295 141.215 ;
        RECT 53.465 140.565 53.725 141.045 ;
        RECT 52.655 140.085 52.985 140.510 ;
        RECT 51.595 140.015 52.490 140.040 ;
        RECT 51.595 140.000 52.500 140.015 ;
        RECT 51.595 139.985 52.505 140.000 ;
        RECT 51.595 139.980 52.515 139.985 ;
        RECT 51.595 139.970 52.520 139.980 ;
        RECT 51.595 139.960 52.525 139.970 ;
        RECT 51.595 139.955 52.535 139.960 ;
        RECT 51.595 139.945 52.545 139.955 ;
        RECT 51.595 139.940 52.555 139.945 ;
        RECT 48.895 139.635 50.320 139.805 ;
        RECT 48.410 138.835 48.945 139.455 ;
        RECT 49.115 138.665 49.445 139.465 ;
        RECT 49.930 139.460 50.320 139.635 ;
        RECT 51.595 139.490 51.855 139.940 ;
        RECT 52.220 139.935 52.555 139.940 ;
        RECT 52.220 139.930 52.570 139.935 ;
        RECT 52.220 139.920 52.585 139.930 ;
        RECT 52.220 139.915 52.610 139.920 ;
        RECT 53.155 139.915 53.385 140.310 ;
        RECT 52.220 139.910 53.385 139.915 ;
        RECT 52.250 139.875 53.385 139.910 ;
        RECT 52.285 139.850 53.385 139.875 ;
        RECT 52.315 139.820 53.385 139.850 ;
        RECT 52.335 139.790 53.385 139.820 ;
        RECT 52.355 139.760 53.385 139.790 ;
        RECT 52.425 139.750 53.385 139.760 ;
        RECT 52.450 139.740 53.385 139.750 ;
        RECT 52.470 139.725 53.385 139.740 ;
        RECT 52.490 139.710 53.385 139.725 ;
        RECT 52.495 139.700 53.280 139.710 ;
        RECT 52.510 139.665 53.280 139.700 ;
        RECT 52.025 139.345 52.355 139.590 ;
        RECT 52.525 139.415 53.280 139.665 ;
        RECT 53.555 139.535 53.725 140.565 ;
        RECT 53.945 140.560 54.275 140.995 ;
        RECT 54.445 140.605 54.615 141.215 ;
        RECT 53.895 140.475 54.275 140.560 ;
        RECT 54.785 140.475 55.115 141.000 ;
        RECT 55.375 140.685 55.585 141.215 ;
        RECT 55.860 140.765 56.645 140.935 ;
        RECT 56.815 140.765 57.220 140.935 ;
        RECT 53.895 140.435 54.120 140.475 ;
        RECT 53.895 139.855 54.065 140.435 ;
        RECT 54.785 140.305 54.985 140.475 ;
        RECT 55.860 140.305 56.030 140.765 ;
        RECT 54.235 139.975 54.985 140.305 ;
        RECT 55.155 139.975 56.030 140.305 ;
        RECT 53.895 139.805 54.110 139.855 ;
        RECT 53.895 139.725 54.285 139.805 ;
        RECT 52.025 139.320 52.210 139.345 ;
        RECT 51.595 139.220 52.210 139.320 ;
        RECT 51.595 138.665 52.200 139.220 ;
        RECT 52.375 138.835 52.855 139.175 ;
        RECT 53.025 138.665 53.280 139.210 ;
        RECT 53.450 138.835 53.725 139.535 ;
        RECT 53.955 138.880 54.285 139.725 ;
        RECT 54.795 139.770 54.985 139.975 ;
        RECT 54.455 138.665 54.625 139.675 ;
        RECT 54.795 139.395 55.690 139.770 ;
        RECT 54.795 138.835 55.135 139.395 ;
        RECT 55.365 138.665 55.680 139.165 ;
        RECT 55.860 139.135 56.030 139.975 ;
        RECT 56.200 140.265 56.665 140.595 ;
        RECT 57.050 140.535 57.220 140.765 ;
        RECT 57.400 140.715 57.770 141.215 ;
        RECT 58.090 140.765 58.765 140.935 ;
        RECT 58.960 140.765 59.295 140.935 ;
        RECT 56.200 139.305 56.520 140.265 ;
        RECT 57.050 140.235 57.880 140.535 ;
        RECT 56.690 139.335 56.880 140.055 ;
        RECT 57.050 139.165 57.220 140.235 ;
        RECT 57.680 140.205 57.880 140.235 ;
        RECT 57.390 139.985 57.560 140.055 ;
        RECT 58.090 139.985 58.260 140.765 ;
        RECT 59.125 140.625 59.295 140.765 ;
        RECT 59.465 140.755 59.715 141.215 ;
        RECT 57.390 139.815 58.260 139.985 ;
        RECT 58.430 140.345 58.955 140.565 ;
        RECT 59.125 140.495 59.350 140.625 ;
        RECT 57.390 139.725 57.900 139.815 ;
        RECT 55.860 138.965 56.745 139.135 ;
        RECT 56.970 138.835 57.220 139.165 ;
        RECT 57.390 138.665 57.560 139.465 ;
        RECT 57.730 139.110 57.900 139.725 ;
        RECT 58.430 139.645 58.600 140.345 ;
        RECT 58.070 139.280 58.600 139.645 ;
        RECT 58.770 139.580 59.010 140.175 ;
        RECT 59.180 139.390 59.350 140.495 ;
        RECT 59.520 139.635 59.800 140.585 ;
        RECT 59.045 139.260 59.350 139.390 ;
        RECT 57.730 138.940 58.835 139.110 ;
        RECT 59.045 138.835 59.295 139.260 ;
        RECT 59.465 138.665 59.730 139.125 ;
        RECT 59.970 138.835 60.155 140.955 ;
        RECT 60.325 140.835 60.655 141.215 ;
        RECT 60.825 140.665 60.995 140.955 ;
        RECT 60.330 140.495 60.995 140.665 ;
        RECT 60.330 139.505 60.560 140.495 ;
        RECT 61.255 140.445 64.765 141.215 ;
        RECT 64.935 140.490 65.225 141.215 ;
        RECT 66.405 140.665 66.575 140.955 ;
        RECT 66.745 140.835 67.075 141.215 ;
        RECT 66.405 140.495 67.070 140.665 ;
        RECT 60.730 139.675 61.080 140.325 ;
        RECT 61.255 139.925 62.905 140.445 ;
        RECT 63.075 139.755 64.765 140.275 ;
        RECT 60.330 139.335 60.995 139.505 ;
        RECT 60.325 138.665 60.655 139.165 ;
        RECT 60.825 138.835 60.995 139.335 ;
        RECT 61.255 138.665 64.765 139.755 ;
        RECT 64.935 138.665 65.225 139.830 ;
        RECT 66.320 139.675 66.670 140.325 ;
        RECT 66.840 139.505 67.070 140.495 ;
        RECT 66.405 139.335 67.070 139.505 ;
        RECT 66.405 138.835 66.575 139.335 ;
        RECT 66.745 138.665 67.075 139.165 ;
        RECT 67.245 138.835 67.430 140.955 ;
        RECT 67.685 140.755 67.935 141.215 ;
        RECT 68.105 140.765 68.440 140.935 ;
        RECT 68.635 140.765 69.310 140.935 ;
        RECT 68.105 140.625 68.275 140.765 ;
        RECT 67.600 139.635 67.880 140.585 ;
        RECT 68.050 140.495 68.275 140.625 ;
        RECT 68.050 139.390 68.220 140.495 ;
        RECT 68.445 140.345 68.970 140.565 ;
        RECT 68.390 139.580 68.630 140.175 ;
        RECT 68.800 139.645 68.970 140.345 ;
        RECT 69.140 139.985 69.310 140.765 ;
        RECT 69.630 140.715 70.000 141.215 ;
        RECT 70.180 140.765 70.585 140.935 ;
        RECT 70.755 140.765 71.540 140.935 ;
        RECT 70.180 140.535 70.350 140.765 ;
        RECT 69.520 140.235 70.350 140.535 ;
        RECT 70.735 140.265 71.200 140.595 ;
        RECT 69.520 140.205 69.720 140.235 ;
        RECT 69.840 139.985 70.010 140.055 ;
        RECT 69.140 139.815 70.010 139.985 ;
        RECT 69.500 139.725 70.010 139.815 ;
        RECT 68.050 139.260 68.355 139.390 ;
        RECT 68.800 139.280 69.330 139.645 ;
        RECT 67.670 138.665 67.935 139.125 ;
        RECT 68.105 138.835 68.355 139.260 ;
        RECT 69.500 139.110 69.670 139.725 ;
        RECT 68.565 138.940 69.670 139.110 ;
        RECT 69.840 138.665 70.010 139.465 ;
        RECT 70.180 139.165 70.350 140.235 ;
        RECT 70.520 139.335 70.710 140.055 ;
        RECT 70.880 139.305 71.200 140.265 ;
        RECT 71.370 140.305 71.540 140.765 ;
        RECT 71.815 140.685 72.025 141.215 ;
        RECT 72.285 140.475 72.615 141.000 ;
        RECT 72.785 140.605 72.955 141.215 ;
        RECT 73.125 140.560 73.455 140.995 ;
        RECT 73.675 140.670 79.020 141.215 ;
        RECT 79.195 140.670 84.540 141.215 ;
        RECT 84.715 140.670 90.060 141.215 ;
        RECT 73.125 140.475 73.505 140.560 ;
        RECT 72.415 140.305 72.615 140.475 ;
        RECT 73.280 140.435 73.505 140.475 ;
        RECT 71.370 139.975 72.245 140.305 ;
        RECT 72.415 139.975 73.165 140.305 ;
        RECT 70.180 138.835 70.430 139.165 ;
        RECT 71.370 139.135 71.540 139.975 ;
        RECT 72.415 139.770 72.605 139.975 ;
        RECT 73.335 139.855 73.505 140.435 ;
        RECT 73.290 139.805 73.505 139.855 ;
        RECT 75.260 139.840 75.600 140.670 ;
        RECT 71.710 139.395 72.605 139.770 ;
        RECT 73.115 139.725 73.505 139.805 ;
        RECT 70.655 138.965 71.540 139.135 ;
        RECT 71.720 138.665 72.035 139.165 ;
        RECT 72.265 138.835 72.605 139.395 ;
        RECT 72.775 138.665 72.945 139.675 ;
        RECT 73.115 138.880 73.445 139.725 ;
        RECT 77.080 139.100 77.430 140.350 ;
        RECT 80.780 139.840 81.120 140.670 ;
        RECT 82.600 139.100 82.950 140.350 ;
        RECT 86.300 139.840 86.640 140.670 ;
        RECT 90.695 140.490 90.985 141.215 ;
        RECT 91.155 140.670 96.500 141.215 ;
        RECT 88.120 139.100 88.470 140.350 ;
        RECT 92.740 139.840 93.080 140.670 ;
        RECT 97.140 140.475 97.395 141.045 ;
        RECT 97.565 140.815 97.895 141.215 ;
        RECT 98.320 140.680 98.850 141.045 ;
        RECT 99.040 140.875 99.315 141.045 ;
        RECT 99.035 140.705 99.315 140.875 ;
        RECT 98.320 140.645 98.495 140.680 ;
        RECT 97.565 140.475 98.495 140.645 ;
        RECT 73.675 138.665 79.020 139.100 ;
        RECT 79.195 138.665 84.540 139.100 ;
        RECT 84.715 138.665 90.060 139.100 ;
        RECT 90.695 138.665 90.985 139.830 ;
        RECT 94.560 139.100 94.910 140.350 ;
        RECT 97.140 139.805 97.310 140.475 ;
        RECT 97.565 140.305 97.735 140.475 ;
        RECT 97.480 139.975 97.735 140.305 ;
        RECT 97.960 139.975 98.155 140.305 ;
        RECT 91.155 138.665 96.500 139.100 ;
        RECT 97.140 138.835 97.475 139.805 ;
        RECT 97.645 138.665 97.815 139.805 ;
        RECT 97.985 139.005 98.155 139.975 ;
        RECT 98.325 139.345 98.495 140.475 ;
        RECT 98.665 139.685 98.835 140.485 ;
        RECT 99.040 139.885 99.315 140.705 ;
        RECT 99.485 139.685 99.675 141.045 ;
        RECT 99.855 140.680 100.365 141.215 ;
        RECT 100.585 140.405 100.830 141.010 ;
        RECT 101.275 140.445 104.785 141.215 ;
        RECT 99.875 140.235 101.105 140.405 ;
        RECT 98.665 139.515 99.675 139.685 ;
        RECT 99.845 139.670 100.595 139.860 ;
        RECT 98.325 139.175 99.450 139.345 ;
        RECT 99.845 139.005 100.015 139.670 ;
        RECT 100.765 139.425 101.105 140.235 ;
        RECT 101.275 139.925 102.925 140.445 ;
        RECT 103.095 139.755 104.785 140.275 ;
        RECT 97.985 138.835 100.015 139.005 ;
        RECT 100.185 138.665 100.355 139.425 ;
        RECT 100.590 139.015 101.105 139.425 ;
        RECT 101.275 138.665 104.785 139.755 ;
        RECT 105.420 139.615 105.755 141.035 ;
        RECT 105.935 140.845 106.680 141.215 ;
        RECT 107.245 140.675 107.500 141.035 ;
        RECT 107.680 140.845 108.010 141.215 ;
        RECT 108.190 140.675 108.415 141.035 ;
        RECT 105.930 140.485 108.415 140.675 ;
        RECT 105.930 139.795 106.155 140.485 ;
        RECT 108.635 140.445 110.305 141.215 ;
        RECT 106.355 139.975 106.635 140.305 ;
        RECT 106.815 139.975 107.390 140.305 ;
        RECT 107.570 139.975 108.005 140.305 ;
        RECT 108.185 139.975 108.455 140.305 ;
        RECT 108.635 139.925 109.385 140.445 ;
        RECT 110.680 140.435 111.180 141.045 ;
        RECT 105.930 139.615 108.425 139.795 ;
        RECT 109.555 139.755 110.305 140.275 ;
        RECT 110.475 139.975 110.825 140.225 ;
        RECT 111.010 139.805 111.180 140.435 ;
        RECT 111.810 140.565 112.140 141.045 ;
        RECT 112.310 140.755 112.535 141.215 ;
        RECT 112.705 140.565 113.035 141.045 ;
        RECT 111.810 140.395 113.035 140.565 ;
        RECT 113.225 140.415 113.475 141.215 ;
        RECT 113.645 140.415 113.985 141.045 ;
        RECT 111.350 140.025 111.680 140.225 ;
        RECT 111.850 140.025 112.180 140.225 ;
        RECT 112.350 140.025 112.770 140.225 ;
        RECT 112.945 140.055 113.640 140.225 ;
        RECT 112.945 139.805 113.115 140.055 ;
        RECT 113.810 139.805 113.985 140.415 ;
        RECT 105.420 138.845 105.685 139.615 ;
        RECT 105.855 138.665 106.185 139.385 ;
        RECT 106.375 139.205 107.565 139.435 ;
        RECT 106.375 138.845 106.635 139.205 ;
        RECT 106.805 138.665 107.135 139.035 ;
        RECT 107.305 138.845 107.565 139.205 ;
        RECT 108.135 138.845 108.425 139.615 ;
        RECT 108.635 138.665 110.305 139.755 ;
        RECT 110.680 139.635 113.115 139.805 ;
        RECT 110.680 138.835 111.010 139.635 ;
        RECT 111.180 138.665 111.510 139.465 ;
        RECT 111.810 138.835 112.140 139.635 ;
        RECT 112.785 138.665 113.035 139.465 ;
        RECT 113.305 138.665 113.475 139.805 ;
        RECT 113.645 138.835 113.985 139.805 ;
        RECT 114.190 140.475 114.805 141.045 ;
        RECT 114.975 140.705 115.190 141.215 ;
        RECT 115.420 140.705 115.700 141.035 ;
        RECT 115.880 140.705 116.120 141.215 ;
        RECT 114.190 139.455 114.505 140.475 ;
        RECT 114.675 139.805 114.845 140.305 ;
        RECT 115.095 139.975 115.360 140.535 ;
        RECT 115.530 139.805 115.700 140.705 ;
        RECT 115.870 139.975 116.225 140.535 ;
        RECT 116.455 140.490 116.745 141.215 ;
        RECT 116.915 140.670 122.260 141.215 ;
        RECT 118.500 139.840 118.840 140.670 ;
        RECT 122.435 140.445 124.105 141.215 ;
        RECT 124.735 140.715 124.995 141.045 ;
        RECT 125.165 140.855 125.495 141.215 ;
        RECT 125.750 140.835 127.050 141.045 ;
        RECT 114.675 139.635 116.100 139.805 ;
        RECT 114.190 138.835 114.725 139.455 ;
        RECT 114.895 138.665 115.225 139.465 ;
        RECT 115.710 139.460 116.100 139.635 ;
        RECT 116.455 138.665 116.745 139.830 ;
        RECT 120.320 139.100 120.670 140.350 ;
        RECT 122.435 139.925 123.185 140.445 ;
        RECT 123.355 139.755 124.105 140.275 ;
        RECT 116.915 138.665 122.260 139.100 ;
        RECT 122.435 138.665 124.105 139.755 ;
        RECT 124.735 139.515 124.905 140.715 ;
        RECT 125.750 140.685 125.920 140.835 ;
        RECT 125.165 140.560 125.920 140.685 ;
        RECT 125.075 140.515 125.920 140.560 ;
        RECT 125.075 140.395 125.345 140.515 ;
        RECT 125.075 139.820 125.245 140.395 ;
        RECT 125.475 139.955 125.885 140.260 ;
        RECT 126.175 140.225 126.385 140.625 ;
        RECT 126.055 140.015 126.385 140.225 ;
        RECT 126.630 140.225 126.850 140.625 ;
        RECT 127.325 140.450 127.780 141.215 ;
        RECT 128.045 140.665 128.215 140.955 ;
        RECT 128.385 140.835 128.715 141.215 ;
        RECT 128.045 140.495 128.710 140.665 ;
        RECT 126.630 140.015 127.105 140.225 ;
        RECT 127.295 140.025 127.785 140.225 ;
        RECT 125.075 139.785 125.275 139.820 ;
        RECT 126.605 139.785 127.780 139.845 ;
        RECT 125.075 139.675 127.780 139.785 ;
        RECT 127.960 139.675 128.310 140.325 ;
        RECT 125.135 139.615 126.935 139.675 ;
        RECT 126.605 139.585 126.935 139.615 ;
        RECT 124.735 138.835 124.995 139.515 ;
        RECT 125.165 138.665 125.415 139.445 ;
        RECT 125.665 139.415 126.500 139.425 ;
        RECT 127.090 139.415 127.275 139.505 ;
        RECT 125.665 139.215 127.275 139.415 ;
        RECT 125.665 138.835 125.915 139.215 ;
        RECT 127.045 139.175 127.275 139.215 ;
        RECT 127.525 139.055 127.780 139.675 ;
        RECT 128.480 139.505 128.710 140.495 ;
        RECT 126.085 138.665 126.440 139.045 ;
        RECT 127.445 138.835 127.780 139.055 ;
        RECT 128.045 139.335 128.710 139.505 ;
        RECT 128.045 138.835 128.215 139.335 ;
        RECT 128.385 138.665 128.715 139.165 ;
        RECT 128.885 138.835 129.070 140.955 ;
        RECT 129.325 140.755 129.575 141.215 ;
        RECT 129.745 140.765 130.080 140.935 ;
        RECT 130.275 140.765 130.950 140.935 ;
        RECT 129.745 140.625 129.915 140.765 ;
        RECT 129.240 139.635 129.520 140.585 ;
        RECT 129.690 140.495 129.915 140.625 ;
        RECT 129.690 139.390 129.860 140.495 ;
        RECT 130.085 140.345 130.610 140.565 ;
        RECT 130.030 139.580 130.270 140.175 ;
        RECT 130.440 139.645 130.610 140.345 ;
        RECT 130.780 139.985 130.950 140.765 ;
        RECT 131.270 140.715 131.640 141.215 ;
        RECT 131.820 140.765 132.225 140.935 ;
        RECT 132.395 140.765 133.180 140.935 ;
        RECT 131.820 140.535 131.990 140.765 ;
        RECT 131.160 140.235 131.990 140.535 ;
        RECT 132.375 140.265 132.840 140.595 ;
        RECT 131.160 140.205 131.360 140.235 ;
        RECT 131.480 139.985 131.650 140.055 ;
        RECT 130.780 139.815 131.650 139.985 ;
        RECT 131.140 139.725 131.650 139.815 ;
        RECT 129.690 139.260 129.995 139.390 ;
        RECT 130.440 139.280 130.970 139.645 ;
        RECT 129.310 138.665 129.575 139.125 ;
        RECT 129.745 138.835 129.995 139.260 ;
        RECT 131.140 139.110 131.310 139.725 ;
        RECT 130.205 138.940 131.310 139.110 ;
        RECT 131.480 138.665 131.650 139.465 ;
        RECT 131.820 139.165 131.990 140.235 ;
        RECT 132.160 139.335 132.350 140.055 ;
        RECT 132.520 139.305 132.840 140.265 ;
        RECT 133.010 140.305 133.180 140.765 ;
        RECT 133.455 140.685 133.665 141.215 ;
        RECT 133.925 140.475 134.255 141.000 ;
        RECT 134.425 140.605 134.595 141.215 ;
        RECT 134.765 140.560 135.095 140.995 ;
        RECT 135.865 140.665 136.035 141.045 ;
        RECT 136.250 140.835 136.580 141.215 ;
        RECT 134.765 140.475 135.145 140.560 ;
        RECT 135.865 140.495 136.580 140.665 ;
        RECT 134.055 140.305 134.255 140.475 ;
        RECT 134.920 140.435 135.145 140.475 ;
        RECT 133.010 139.975 133.885 140.305 ;
        RECT 134.055 139.975 134.805 140.305 ;
        RECT 131.820 138.835 132.070 139.165 ;
        RECT 133.010 139.135 133.180 139.975 ;
        RECT 134.055 139.770 134.245 139.975 ;
        RECT 134.975 139.855 135.145 140.435 ;
        RECT 135.775 139.945 136.130 140.315 ;
        RECT 136.410 140.305 136.580 140.495 ;
        RECT 136.750 140.470 137.005 141.045 ;
        RECT 136.410 139.975 136.665 140.305 ;
        RECT 134.930 139.805 135.145 139.855 ;
        RECT 133.350 139.395 134.245 139.770 ;
        RECT 134.755 139.725 135.145 139.805 ;
        RECT 136.410 139.765 136.580 139.975 ;
        RECT 132.295 138.965 133.180 139.135 ;
        RECT 133.360 138.665 133.675 139.165 ;
        RECT 133.905 138.835 134.245 139.395 ;
        RECT 134.415 138.665 134.585 139.675 ;
        RECT 134.755 138.880 135.085 139.725 ;
        RECT 135.865 139.595 136.580 139.765 ;
        RECT 136.835 139.740 137.005 140.470 ;
        RECT 137.180 140.375 137.440 141.215 ;
        RECT 137.615 140.465 138.825 141.215 ;
        RECT 135.865 138.835 136.035 139.595 ;
        RECT 136.250 138.665 136.580 139.425 ;
        RECT 136.750 138.835 137.005 139.740 ;
        RECT 137.180 138.665 137.440 139.815 ;
        RECT 137.615 139.755 138.135 140.295 ;
        RECT 138.305 139.925 138.825 140.465 ;
        RECT 137.615 138.665 138.825 139.755 ;
        RECT 13.330 138.495 138.910 138.665 ;
        RECT 13.415 137.405 14.625 138.495 ;
        RECT 14.795 137.405 18.305 138.495 ;
        RECT 13.415 136.695 13.935 137.235 ;
        RECT 14.105 136.865 14.625 137.405 ;
        RECT 14.795 136.715 16.445 137.235 ;
        RECT 16.615 136.885 18.305 137.405 ;
        RECT 18.475 138.065 18.815 138.325 ;
        RECT 13.415 135.945 14.625 136.695 ;
        RECT 14.795 135.945 18.305 136.715 ;
        RECT 18.475 136.665 18.735 138.065 ;
        RECT 18.985 137.695 19.315 138.495 ;
        RECT 19.780 137.525 20.030 138.325 ;
        RECT 20.215 137.775 20.545 138.495 ;
        RECT 20.765 137.525 21.015 138.325 ;
        RECT 21.185 138.115 21.520 138.495 ;
        RECT 18.925 137.355 21.115 137.525 ;
        RECT 18.925 137.185 19.240 137.355 ;
        RECT 18.910 136.935 19.240 137.185 ;
        RECT 18.475 136.155 18.815 136.665 ;
        RECT 18.985 135.945 19.255 136.745 ;
        RECT 19.435 136.215 19.715 137.185 ;
        RECT 19.895 136.215 20.195 137.185 ;
        RECT 20.375 136.220 20.725 137.185 ;
        RECT 20.945 136.445 21.115 137.355 ;
        RECT 21.285 136.625 21.525 137.935 ;
        RECT 21.730 137.705 22.265 138.325 ;
        RECT 21.730 136.685 22.045 137.705 ;
        RECT 22.435 137.695 22.765 138.495 ;
        RECT 23.250 137.525 23.640 137.700 ;
        RECT 22.215 137.355 23.640 137.525 ;
        RECT 23.995 137.625 24.270 138.325 ;
        RECT 24.440 137.950 24.695 138.495 ;
        RECT 24.865 137.985 25.345 138.325 ;
        RECT 25.520 137.940 26.125 138.495 ;
        RECT 25.510 137.840 26.125 137.940 ;
        RECT 25.510 137.815 25.695 137.840 ;
        RECT 22.215 136.855 22.385 137.355 ;
        RECT 20.945 136.115 21.440 136.445 ;
        RECT 21.730 136.115 22.345 136.685 ;
        RECT 22.635 136.625 22.900 137.185 ;
        RECT 23.070 136.455 23.240 137.355 ;
        RECT 23.410 136.625 23.765 137.185 ;
        RECT 23.995 136.595 24.165 137.625 ;
        RECT 24.440 137.495 25.195 137.745 ;
        RECT 25.365 137.570 25.695 137.815 ;
        RECT 24.440 137.460 25.210 137.495 ;
        RECT 24.440 137.450 25.225 137.460 ;
        RECT 24.335 137.435 25.230 137.450 ;
        RECT 24.335 137.420 25.250 137.435 ;
        RECT 24.335 137.410 25.270 137.420 ;
        RECT 24.335 137.400 25.295 137.410 ;
        RECT 24.335 137.370 25.365 137.400 ;
        RECT 24.335 137.340 25.385 137.370 ;
        RECT 24.335 137.310 25.405 137.340 ;
        RECT 24.335 137.285 25.435 137.310 ;
        RECT 24.335 137.250 25.470 137.285 ;
        RECT 24.335 137.245 25.500 137.250 ;
        RECT 24.335 136.850 24.565 137.245 ;
        RECT 25.110 137.240 25.500 137.245 ;
        RECT 25.135 137.230 25.500 137.240 ;
        RECT 25.150 137.225 25.500 137.230 ;
        RECT 25.165 137.220 25.500 137.225 ;
        RECT 25.865 137.220 26.125 137.670 ;
        RECT 26.295 137.330 26.585 138.495 ;
        RECT 26.765 137.525 27.095 138.310 ;
        RECT 26.765 137.355 27.445 137.525 ;
        RECT 27.625 137.355 27.955 138.495 ;
        RECT 28.135 138.060 33.480 138.495 ;
        RECT 25.165 137.215 26.125 137.220 ;
        RECT 25.175 137.205 26.125 137.215 ;
        RECT 25.185 137.200 26.125 137.205 ;
        RECT 25.195 137.190 26.125 137.200 ;
        RECT 25.200 137.180 26.125 137.190 ;
        RECT 25.205 137.175 26.125 137.180 ;
        RECT 25.215 137.160 26.125 137.175 ;
        RECT 25.220 137.145 26.125 137.160 ;
        RECT 25.230 137.120 26.125 137.145 ;
        RECT 24.735 136.650 25.065 137.075 ;
        RECT 22.515 135.945 22.730 136.455 ;
        RECT 22.960 136.125 23.240 136.455 ;
        RECT 23.420 135.945 23.660 136.455 ;
        RECT 23.995 136.115 24.255 136.595 ;
        RECT 24.425 135.945 24.675 136.485 ;
        RECT 24.845 136.165 25.065 136.650 ;
        RECT 25.235 137.050 26.125 137.120 ;
        RECT 25.235 136.325 25.405 137.050 ;
        RECT 26.755 136.935 27.105 137.185 ;
        RECT 25.575 136.495 26.125 136.880 ;
        RECT 27.275 136.755 27.445 137.355 ;
        RECT 27.615 136.935 27.965 137.185 ;
        RECT 25.235 136.155 26.125 136.325 ;
        RECT 26.295 135.945 26.585 136.670 ;
        RECT 26.775 135.945 27.015 136.755 ;
        RECT 27.185 136.115 27.515 136.755 ;
        RECT 27.685 135.945 27.955 136.755 ;
        RECT 29.720 136.490 30.060 137.320 ;
        RECT 31.540 136.810 31.890 138.060 ;
        RECT 33.665 137.545 33.940 138.315 ;
        RECT 34.110 137.885 34.440 138.315 ;
        RECT 34.610 138.055 34.805 138.495 ;
        RECT 34.985 137.885 35.315 138.315 ;
        RECT 35.495 138.060 40.840 138.495 ;
        RECT 41.015 138.060 46.360 138.495 ;
        RECT 34.110 137.715 35.315 137.885 ;
        RECT 33.665 137.355 34.250 137.545 ;
        RECT 34.420 137.385 35.315 137.715 ;
        RECT 33.665 136.535 33.905 137.185 ;
        RECT 34.075 136.685 34.250 137.355 ;
        RECT 34.420 136.855 34.835 137.185 ;
        RECT 35.015 136.855 35.310 137.185 ;
        RECT 34.075 136.505 34.405 136.685 ;
        RECT 28.135 135.945 33.480 136.490 ;
        RECT 33.680 135.945 34.010 136.335 ;
        RECT 34.180 136.125 34.405 136.505 ;
        RECT 34.605 136.235 34.835 136.855 ;
        RECT 35.015 135.945 35.315 136.675 ;
        RECT 37.080 136.490 37.420 137.320 ;
        RECT 38.900 136.810 39.250 138.060 ;
        RECT 42.600 136.490 42.940 137.320 ;
        RECT 44.420 136.810 44.770 138.060 ;
        RECT 46.535 137.405 49.125 138.495 ;
        RECT 46.535 136.715 47.745 137.235 ;
        RECT 47.915 136.885 49.125 137.405 ;
        RECT 49.305 137.525 49.635 138.310 ;
        RECT 49.305 137.355 49.985 137.525 ;
        RECT 50.165 137.355 50.495 138.495 ;
        RECT 50.685 137.525 51.015 138.310 ;
        RECT 50.685 137.355 51.365 137.525 ;
        RECT 51.545 137.355 51.875 138.495 ;
        RECT 49.295 136.935 49.645 137.185 ;
        RECT 49.815 136.755 49.985 137.355 ;
        RECT 50.155 136.935 50.505 137.185 ;
        RECT 50.675 136.935 51.025 137.185 ;
        RECT 51.195 136.755 51.365 137.355 ;
        RECT 52.055 137.330 52.345 138.495 ;
        RECT 52.515 137.395 52.835 138.325 ;
        RECT 53.015 137.815 53.415 138.325 ;
        RECT 53.585 137.985 53.755 138.495 ;
        RECT 53.925 137.815 54.255 138.325 ;
        RECT 53.015 137.645 54.255 137.815 ;
        RECT 54.425 137.645 54.595 138.495 ;
        RECT 55.185 137.645 55.565 138.325 ;
        RECT 55.735 138.060 61.080 138.495 ;
        RECT 52.515 137.225 53.145 137.395 ;
        RECT 51.535 136.935 51.885 137.185 ;
        RECT 35.495 135.945 40.840 136.490 ;
        RECT 41.015 135.945 46.360 136.490 ;
        RECT 46.535 135.945 49.125 136.715 ;
        RECT 49.315 135.945 49.555 136.755 ;
        RECT 49.725 136.115 50.055 136.755 ;
        RECT 50.225 135.945 50.495 136.755 ;
        RECT 50.695 135.945 50.935 136.755 ;
        RECT 51.105 136.115 51.435 136.755 ;
        RECT 51.605 135.945 51.875 136.755 ;
        RECT 52.055 135.945 52.345 136.670 ;
        RECT 52.515 135.945 52.805 136.780 ;
        RECT 52.975 136.345 53.145 137.225 ;
        RECT 53.920 137.305 55.225 137.475 ;
        RECT 53.315 136.685 53.545 137.185 ;
        RECT 53.920 137.105 54.090 137.305 ;
        RECT 53.715 136.935 54.090 137.105 ;
        RECT 54.260 136.935 54.810 137.135 ;
        RECT 54.980 136.855 55.225 137.305 ;
        RECT 55.395 136.685 55.565 137.645 ;
        RECT 53.315 136.515 55.565 136.685 ;
        RECT 52.975 136.175 53.930 136.345 ;
        RECT 54.345 135.945 54.675 136.335 ;
        RECT 54.845 136.195 55.015 136.515 ;
        RECT 57.320 136.490 57.660 137.320 ;
        RECT 59.140 136.810 59.490 138.060 ;
        RECT 61.255 137.405 63.845 138.495 ;
        RECT 64.565 137.825 64.735 138.325 ;
        RECT 64.905 137.995 65.235 138.495 ;
        RECT 64.565 137.655 65.230 137.825 ;
        RECT 61.255 136.715 62.465 137.235 ;
        RECT 62.635 136.885 63.845 137.405 ;
        RECT 64.480 136.835 64.830 137.485 ;
        RECT 55.185 135.945 55.515 136.335 ;
        RECT 55.735 135.945 61.080 136.490 ;
        RECT 61.255 135.945 63.845 136.715 ;
        RECT 65.000 136.665 65.230 137.655 ;
        RECT 64.565 136.495 65.230 136.665 ;
        RECT 64.565 136.205 64.735 136.495 ;
        RECT 64.905 135.945 65.235 136.325 ;
        RECT 65.405 136.205 65.590 138.325 ;
        RECT 65.830 138.035 66.095 138.495 ;
        RECT 66.265 137.900 66.515 138.325 ;
        RECT 66.725 138.050 67.830 138.220 ;
        RECT 66.210 137.770 66.515 137.900 ;
        RECT 65.760 136.575 66.040 137.525 ;
        RECT 66.210 136.665 66.380 137.770 ;
        RECT 66.550 136.985 66.790 137.580 ;
        RECT 66.960 137.515 67.490 137.880 ;
        RECT 66.960 136.815 67.130 137.515 ;
        RECT 67.660 137.435 67.830 138.050 ;
        RECT 68.000 137.695 68.170 138.495 ;
        RECT 68.340 137.995 68.590 138.325 ;
        RECT 68.815 138.025 69.700 138.195 ;
        RECT 67.660 137.345 68.170 137.435 ;
        RECT 66.210 136.535 66.435 136.665 ;
        RECT 66.605 136.595 67.130 136.815 ;
        RECT 67.300 137.175 68.170 137.345 ;
        RECT 65.845 135.945 66.095 136.405 ;
        RECT 66.265 136.395 66.435 136.535 ;
        RECT 67.300 136.395 67.470 137.175 ;
        RECT 68.000 137.105 68.170 137.175 ;
        RECT 67.680 136.925 67.880 136.955 ;
        RECT 68.340 136.925 68.510 137.995 ;
        RECT 68.680 137.105 68.870 137.825 ;
        RECT 67.680 136.625 68.510 136.925 ;
        RECT 69.040 136.895 69.360 137.855 ;
        RECT 66.265 136.225 66.600 136.395 ;
        RECT 66.795 136.225 67.470 136.395 ;
        RECT 67.790 135.945 68.160 136.445 ;
        RECT 68.340 136.395 68.510 136.625 ;
        RECT 68.895 136.565 69.360 136.895 ;
        RECT 69.530 137.185 69.700 138.025 ;
        RECT 69.880 137.995 70.195 138.495 ;
        RECT 70.425 137.765 70.765 138.325 ;
        RECT 69.870 137.390 70.765 137.765 ;
        RECT 70.935 137.485 71.105 138.495 ;
        RECT 70.575 137.185 70.765 137.390 ;
        RECT 71.275 137.435 71.605 138.280 ;
        RECT 71.775 137.580 71.945 138.495 ;
        RECT 71.275 137.355 71.665 137.435 ;
        RECT 71.450 137.305 71.665 137.355 ;
        RECT 69.530 136.855 70.405 137.185 ;
        RECT 70.575 136.855 71.325 137.185 ;
        RECT 69.530 136.395 69.700 136.855 ;
        RECT 70.575 136.685 70.775 136.855 ;
        RECT 71.495 136.725 71.665 137.305 ;
        RECT 71.440 136.685 71.665 136.725 ;
        RECT 68.340 136.225 68.745 136.395 ;
        RECT 68.915 136.225 69.700 136.395 ;
        RECT 69.975 135.945 70.185 136.475 ;
        RECT 70.445 136.160 70.775 136.685 ;
        RECT 71.285 136.600 71.665 136.685 ;
        RECT 72.300 137.355 72.635 138.325 ;
        RECT 72.805 137.355 72.975 138.495 ;
        RECT 73.145 138.155 75.175 138.325 ;
        RECT 72.300 136.685 72.470 137.355 ;
        RECT 73.145 137.185 73.315 138.155 ;
        RECT 72.640 136.855 72.895 137.185 ;
        RECT 73.120 136.855 73.315 137.185 ;
        RECT 73.485 137.815 74.610 137.985 ;
        RECT 72.725 136.685 72.895 136.855 ;
        RECT 73.485 136.685 73.655 137.815 ;
        RECT 70.945 135.945 71.115 136.555 ;
        RECT 71.285 136.165 71.615 136.600 ;
        RECT 71.785 135.945 71.955 136.460 ;
        RECT 72.300 136.115 72.555 136.685 ;
        RECT 72.725 136.515 73.655 136.685 ;
        RECT 73.825 137.475 74.835 137.645 ;
        RECT 73.825 136.675 73.995 137.475 ;
        RECT 74.200 137.135 74.475 137.275 ;
        RECT 74.195 136.965 74.475 137.135 ;
        RECT 73.480 136.480 73.655 136.515 ;
        RECT 72.725 135.945 73.055 136.345 ;
        RECT 73.480 136.115 74.010 136.480 ;
        RECT 74.200 136.115 74.475 136.965 ;
        RECT 74.645 136.115 74.835 137.475 ;
        RECT 75.005 137.490 75.175 138.155 ;
        RECT 75.345 137.735 75.515 138.495 ;
        RECT 75.750 137.735 76.265 138.145 ;
        RECT 75.005 137.300 75.755 137.490 ;
        RECT 75.925 136.925 76.265 137.735 ;
        RECT 76.435 137.405 77.645 138.495 ;
        RECT 75.035 136.755 76.265 136.925 ;
        RECT 75.015 135.945 75.525 136.480 ;
        RECT 75.745 136.150 75.990 136.755 ;
        RECT 76.435 136.695 76.955 137.235 ;
        RECT 77.125 136.865 77.645 137.405 ;
        RECT 77.815 137.330 78.105 138.495 ;
        RECT 78.365 137.825 78.535 138.325 ;
        RECT 78.705 137.995 79.035 138.495 ;
        RECT 78.365 137.655 79.030 137.825 ;
        RECT 78.280 136.835 78.630 137.485 ;
        RECT 76.435 135.945 77.645 136.695 ;
        RECT 77.815 135.945 78.105 136.670 ;
        RECT 78.800 136.665 79.030 137.655 ;
        RECT 78.365 136.495 79.030 136.665 ;
        RECT 78.365 136.205 78.535 136.495 ;
        RECT 78.705 135.945 79.035 136.325 ;
        RECT 79.205 136.205 79.390 138.325 ;
        RECT 79.630 138.035 79.895 138.495 ;
        RECT 80.065 137.900 80.315 138.325 ;
        RECT 80.525 138.050 81.630 138.220 ;
        RECT 80.010 137.770 80.315 137.900 ;
        RECT 79.560 136.575 79.840 137.525 ;
        RECT 80.010 136.665 80.180 137.770 ;
        RECT 80.350 136.985 80.590 137.580 ;
        RECT 80.760 137.515 81.290 137.880 ;
        RECT 80.760 136.815 80.930 137.515 ;
        RECT 81.460 137.435 81.630 138.050 ;
        RECT 81.800 137.695 81.970 138.495 ;
        RECT 82.140 137.995 82.390 138.325 ;
        RECT 82.615 138.025 83.500 138.195 ;
        RECT 81.460 137.345 81.970 137.435 ;
        RECT 80.010 136.535 80.235 136.665 ;
        RECT 80.405 136.595 80.930 136.815 ;
        RECT 81.100 137.175 81.970 137.345 ;
        RECT 79.645 135.945 79.895 136.405 ;
        RECT 80.065 136.395 80.235 136.535 ;
        RECT 81.100 136.395 81.270 137.175 ;
        RECT 81.800 137.105 81.970 137.175 ;
        RECT 81.480 136.925 81.680 136.955 ;
        RECT 82.140 136.925 82.310 137.995 ;
        RECT 82.480 137.105 82.670 137.825 ;
        RECT 81.480 136.625 82.310 136.925 ;
        RECT 82.840 136.895 83.160 137.855 ;
        RECT 80.065 136.225 80.400 136.395 ;
        RECT 80.595 136.225 81.270 136.395 ;
        RECT 81.590 135.945 81.960 136.445 ;
        RECT 82.140 136.395 82.310 136.625 ;
        RECT 82.695 136.565 83.160 136.895 ;
        RECT 83.330 137.185 83.500 138.025 ;
        RECT 83.680 137.995 83.995 138.495 ;
        RECT 84.225 137.765 84.565 138.325 ;
        RECT 83.670 137.390 84.565 137.765 ;
        RECT 84.735 137.485 84.905 138.495 ;
        RECT 84.375 137.185 84.565 137.390 ;
        RECT 85.075 137.435 85.405 138.280 ;
        RECT 85.575 137.580 85.745 138.495 ;
        RECT 85.075 137.355 85.465 137.435 ;
        RECT 85.250 137.305 85.465 137.355 ;
        RECT 83.330 136.855 84.205 137.185 ;
        RECT 84.375 136.855 85.125 137.185 ;
        RECT 83.330 136.395 83.500 136.855 ;
        RECT 84.375 136.685 84.575 136.855 ;
        RECT 85.295 136.725 85.465 137.305 ;
        RECT 85.240 136.685 85.465 136.725 ;
        RECT 82.140 136.225 82.545 136.395 ;
        RECT 82.715 136.225 83.500 136.395 ;
        RECT 83.775 135.945 83.985 136.475 ;
        RECT 84.245 136.160 84.575 136.685 ;
        RECT 85.085 136.600 85.465 136.685 ;
        RECT 86.100 137.355 86.435 138.325 ;
        RECT 86.605 137.355 86.775 138.495 ;
        RECT 86.945 138.155 88.975 138.325 ;
        RECT 86.100 136.685 86.270 137.355 ;
        RECT 86.945 137.185 87.115 138.155 ;
        RECT 86.440 136.855 86.695 137.185 ;
        RECT 86.920 136.855 87.115 137.185 ;
        RECT 87.285 137.815 88.410 137.985 ;
        RECT 86.525 136.685 86.695 136.855 ;
        RECT 87.285 136.685 87.455 137.815 ;
        RECT 84.745 135.945 84.915 136.555 ;
        RECT 85.085 136.165 85.415 136.600 ;
        RECT 85.585 135.945 85.755 136.460 ;
        RECT 86.100 136.115 86.355 136.685 ;
        RECT 86.525 136.515 87.455 136.685 ;
        RECT 87.625 137.475 88.635 137.645 ;
        RECT 87.625 136.675 87.795 137.475 ;
        RECT 87.280 136.480 87.455 136.515 ;
        RECT 86.525 135.945 86.855 136.345 ;
        RECT 87.280 136.115 87.810 136.480 ;
        RECT 88.000 136.455 88.275 137.275 ;
        RECT 87.995 136.285 88.275 136.455 ;
        RECT 88.000 136.115 88.275 136.285 ;
        RECT 88.445 136.115 88.635 137.475 ;
        RECT 88.805 137.490 88.975 138.155 ;
        RECT 89.145 137.735 89.315 138.495 ;
        RECT 89.550 137.735 90.065 138.145 ;
        RECT 88.805 137.300 89.555 137.490 ;
        RECT 89.725 136.925 90.065 137.735 ;
        RECT 90.235 137.405 93.745 138.495 ;
        RECT 88.835 136.755 90.065 136.925 ;
        RECT 88.815 135.945 89.325 136.480 ;
        RECT 89.545 136.150 89.790 136.755 ;
        RECT 90.235 136.715 91.885 137.235 ;
        RECT 92.055 136.885 93.745 137.405 ;
        RECT 94.380 137.355 94.715 138.325 ;
        RECT 94.885 137.355 95.055 138.495 ;
        RECT 95.225 138.155 97.255 138.325 ;
        RECT 90.235 135.945 93.745 136.715 ;
        RECT 94.380 136.685 94.550 137.355 ;
        RECT 95.225 137.185 95.395 138.155 ;
        RECT 94.720 136.855 94.975 137.185 ;
        RECT 95.200 136.855 95.395 137.185 ;
        RECT 95.565 137.815 96.690 137.985 ;
        RECT 94.805 136.685 94.975 136.855 ;
        RECT 95.565 136.685 95.735 137.815 ;
        RECT 94.380 136.115 94.635 136.685 ;
        RECT 94.805 136.515 95.735 136.685 ;
        RECT 95.905 137.475 96.915 137.645 ;
        RECT 95.905 136.675 96.075 137.475 ;
        RECT 96.280 136.795 96.555 137.275 ;
        RECT 96.275 136.625 96.555 136.795 ;
        RECT 95.560 136.480 95.735 136.515 ;
        RECT 94.805 135.945 95.135 136.345 ;
        RECT 95.560 136.115 96.090 136.480 ;
        RECT 96.280 136.115 96.555 136.625 ;
        RECT 96.725 136.115 96.915 137.475 ;
        RECT 97.085 137.490 97.255 138.155 ;
        RECT 97.425 137.735 97.595 138.495 ;
        RECT 97.830 137.735 98.345 138.145 ;
        RECT 97.085 137.300 97.835 137.490 ;
        RECT 98.005 136.925 98.345 137.735 ;
        RECT 97.115 136.755 98.345 136.925 ;
        RECT 98.515 137.355 98.900 138.325 ;
        RECT 99.070 138.035 99.395 138.495 ;
        RECT 99.915 137.865 100.195 138.325 ;
        RECT 99.070 137.645 100.195 137.865 ;
        RECT 97.095 135.945 97.605 136.480 ;
        RECT 97.825 136.150 98.070 136.755 ;
        RECT 98.515 136.685 98.795 137.355 ;
        RECT 99.070 137.185 99.520 137.645 ;
        RECT 100.385 137.475 100.785 138.325 ;
        RECT 101.185 138.035 101.455 138.495 ;
        RECT 101.625 137.865 101.910 138.325 ;
        RECT 98.965 136.855 99.520 137.185 ;
        RECT 99.690 136.915 100.785 137.475 ;
        RECT 99.070 136.745 99.520 136.855 ;
        RECT 98.515 136.115 98.900 136.685 ;
        RECT 99.070 136.575 100.195 136.745 ;
        RECT 99.070 135.945 99.395 136.405 ;
        RECT 99.915 136.115 100.195 136.575 ;
        RECT 100.385 136.115 100.785 136.915 ;
        RECT 100.955 137.645 101.910 137.865 ;
        RECT 100.955 136.745 101.165 137.645 ;
        RECT 101.335 136.915 102.025 137.475 ;
        RECT 102.195 137.405 103.405 138.495 ;
        RECT 100.955 136.575 101.910 136.745 ;
        RECT 101.185 135.945 101.455 136.405 ;
        RECT 101.625 136.115 101.910 136.575 ;
        RECT 102.195 136.695 102.715 137.235 ;
        RECT 102.885 136.865 103.405 137.405 ;
        RECT 103.575 137.330 103.865 138.495 ;
        RECT 104.035 137.405 106.625 138.495 ;
        RECT 104.035 136.715 105.245 137.235 ;
        RECT 105.415 136.885 106.625 137.405 ;
        RECT 107.260 137.545 107.525 138.315 ;
        RECT 107.695 137.775 108.025 138.495 ;
        RECT 108.215 137.955 108.475 138.315 ;
        RECT 108.645 138.125 108.975 138.495 ;
        RECT 109.145 137.955 109.405 138.315 ;
        RECT 108.215 137.725 109.405 137.955 ;
        RECT 109.975 137.545 110.265 138.315 ;
        RECT 102.195 135.945 103.405 136.695 ;
        RECT 103.575 135.945 103.865 136.670 ;
        RECT 104.035 135.945 106.625 136.715 ;
        RECT 107.260 136.125 107.595 137.545 ;
        RECT 107.770 137.365 110.265 137.545 ;
        RECT 110.480 137.545 110.745 138.315 ;
        RECT 110.915 137.775 111.245 138.495 ;
        RECT 111.435 137.955 111.695 138.315 ;
        RECT 111.865 138.125 112.195 138.495 ;
        RECT 112.365 137.955 112.625 138.315 ;
        RECT 111.435 137.725 112.625 137.955 ;
        RECT 113.195 137.545 113.485 138.315 ;
        RECT 107.770 136.675 107.995 137.365 ;
        RECT 108.195 136.855 108.475 137.185 ;
        RECT 108.655 136.855 109.230 137.185 ;
        RECT 109.410 136.855 109.845 137.185 ;
        RECT 110.025 136.855 110.295 137.185 ;
        RECT 107.770 136.485 110.255 136.675 ;
        RECT 107.775 135.945 108.520 136.315 ;
        RECT 109.085 136.125 109.340 136.485 ;
        RECT 109.520 135.945 109.850 136.315 ;
        RECT 110.030 136.125 110.255 136.485 ;
        RECT 110.480 136.125 110.815 137.545 ;
        RECT 110.990 137.365 113.485 137.545 ;
        RECT 113.730 137.705 114.265 138.325 ;
        RECT 110.990 136.675 111.215 137.365 ;
        RECT 111.415 136.855 111.695 137.185 ;
        RECT 111.875 136.855 112.450 137.185 ;
        RECT 112.630 136.855 113.065 137.185 ;
        RECT 113.245 136.855 113.515 137.185 ;
        RECT 113.730 136.685 114.045 137.705 ;
        RECT 114.435 137.695 114.765 138.495 ;
        RECT 115.250 137.525 115.640 137.700 ;
        RECT 114.215 137.355 115.640 137.525 ;
        RECT 115.995 137.405 117.665 138.495 ;
        RECT 114.215 136.855 114.385 137.355 ;
        RECT 110.990 136.485 113.475 136.675 ;
        RECT 110.995 135.945 111.740 136.315 ;
        RECT 112.305 136.125 112.560 136.485 ;
        RECT 112.740 135.945 113.070 136.315 ;
        RECT 113.250 136.125 113.475 136.485 ;
        RECT 113.730 136.115 114.345 136.685 ;
        RECT 114.635 136.625 114.900 137.185 ;
        RECT 115.070 136.455 115.240 137.355 ;
        RECT 115.410 136.625 115.765 137.185 ;
        RECT 115.995 136.715 116.745 137.235 ;
        RECT 116.915 136.885 117.665 137.405 ;
        RECT 117.835 137.645 118.095 138.325 ;
        RECT 118.265 137.715 118.515 138.495 ;
        RECT 118.765 137.945 119.015 138.325 ;
        RECT 119.185 138.115 119.540 138.495 ;
        RECT 120.545 138.105 120.880 138.325 ;
        RECT 120.145 137.945 120.375 137.985 ;
        RECT 118.765 137.745 120.375 137.945 ;
        RECT 118.765 137.735 119.600 137.745 ;
        RECT 120.190 137.655 120.375 137.745 ;
        RECT 114.515 135.945 114.730 136.455 ;
        RECT 114.960 136.125 115.240 136.455 ;
        RECT 115.420 135.945 115.660 136.455 ;
        RECT 115.995 135.945 117.665 136.715 ;
        RECT 117.835 136.445 118.005 137.645 ;
        RECT 119.705 137.545 120.035 137.575 ;
        RECT 118.235 137.485 120.035 137.545 ;
        RECT 120.625 137.485 120.880 138.105 ;
        RECT 121.055 138.060 126.400 138.495 ;
        RECT 118.175 137.375 120.880 137.485 ;
        RECT 118.175 137.340 118.375 137.375 ;
        RECT 118.175 136.765 118.345 137.340 ;
        RECT 119.705 137.315 120.880 137.375 ;
        RECT 118.575 136.900 118.985 137.205 ;
        RECT 119.155 136.935 119.485 137.145 ;
        RECT 118.175 136.645 118.445 136.765 ;
        RECT 118.175 136.600 119.020 136.645 ;
        RECT 118.265 136.475 119.020 136.600 ;
        RECT 119.275 136.535 119.485 136.935 ;
        RECT 119.730 136.935 120.205 137.145 ;
        RECT 120.395 136.935 120.885 137.135 ;
        RECT 119.730 136.535 119.950 136.935 ;
        RECT 117.835 136.115 118.095 136.445 ;
        RECT 118.850 136.325 119.020 136.475 ;
        RECT 118.265 135.945 118.595 136.305 ;
        RECT 118.850 136.115 120.150 136.325 ;
        RECT 120.425 135.945 120.880 136.710 ;
        RECT 122.640 136.490 122.980 137.320 ;
        RECT 124.460 136.810 124.810 138.060 ;
        RECT 127.220 137.525 127.610 137.700 ;
        RECT 128.095 137.695 128.425 138.495 ;
        RECT 128.595 137.705 129.130 138.325 ;
        RECT 127.220 137.355 128.645 137.525 ;
        RECT 127.095 136.625 127.450 137.185 ;
        RECT 121.055 135.945 126.400 136.490 ;
        RECT 127.620 136.455 127.790 137.355 ;
        RECT 127.960 136.625 128.225 137.185 ;
        RECT 128.475 136.855 128.645 137.355 ;
        RECT 128.815 136.685 129.130 137.705 ;
        RECT 129.335 137.330 129.625 138.495 ;
        RECT 130.000 137.525 130.330 138.325 ;
        RECT 130.500 137.695 130.830 138.495 ;
        RECT 131.130 137.525 131.460 138.325 ;
        RECT 132.105 137.695 132.355 138.495 ;
        RECT 130.000 137.355 132.435 137.525 ;
        RECT 132.625 137.355 132.795 138.495 ;
        RECT 132.965 137.355 133.305 138.325 ;
        RECT 129.795 136.935 130.145 137.185 ;
        RECT 130.330 136.725 130.500 137.355 ;
        RECT 130.670 136.935 131.000 137.135 ;
        RECT 131.170 136.935 131.500 137.135 ;
        RECT 131.670 136.935 132.090 137.135 ;
        RECT 132.265 137.105 132.435 137.355 ;
        RECT 132.265 136.935 132.960 137.105 ;
        RECT 127.200 135.945 127.440 136.455 ;
        RECT 127.620 136.125 127.900 136.455 ;
        RECT 128.130 135.945 128.345 136.455 ;
        RECT 128.515 136.115 129.130 136.685 ;
        RECT 129.335 135.945 129.625 136.670 ;
        RECT 130.000 136.115 130.500 136.725 ;
        RECT 131.130 136.595 132.355 136.765 ;
        RECT 133.130 136.745 133.305 137.355 ;
        RECT 131.130 136.115 131.460 136.595 ;
        RECT 131.630 135.945 131.855 136.405 ;
        RECT 132.025 136.115 132.355 136.595 ;
        RECT 132.545 135.945 132.795 136.745 ;
        RECT 132.965 136.115 133.305 136.745 ;
        RECT 133.475 137.645 133.735 138.325 ;
        RECT 133.905 137.715 134.155 138.495 ;
        RECT 134.405 137.945 134.655 138.325 ;
        RECT 134.825 138.115 135.180 138.495 ;
        RECT 136.185 138.105 136.520 138.325 ;
        RECT 135.785 137.945 136.015 137.985 ;
        RECT 134.405 137.745 136.015 137.945 ;
        RECT 134.405 137.735 135.240 137.745 ;
        RECT 135.830 137.655 136.015 137.745 ;
        RECT 133.475 136.445 133.645 137.645 ;
        RECT 135.345 137.545 135.675 137.575 ;
        RECT 133.875 137.485 135.675 137.545 ;
        RECT 136.265 137.485 136.520 138.105 ;
        RECT 133.815 137.375 136.520 137.485 ;
        RECT 133.815 137.340 134.015 137.375 ;
        RECT 133.815 136.765 133.985 137.340 ;
        RECT 135.345 137.315 136.520 137.375 ;
        RECT 137.615 137.405 138.825 138.495 ;
        RECT 134.215 136.900 134.625 137.205 ;
        RECT 134.795 136.935 135.125 137.145 ;
        RECT 133.815 136.645 134.085 136.765 ;
        RECT 133.815 136.600 134.660 136.645 ;
        RECT 133.905 136.475 134.660 136.600 ;
        RECT 134.915 136.535 135.125 136.935 ;
        RECT 135.370 136.935 135.845 137.145 ;
        RECT 136.035 136.935 136.525 137.135 ;
        RECT 135.370 136.535 135.590 136.935 ;
        RECT 137.615 136.865 138.135 137.405 ;
        RECT 133.475 136.115 133.735 136.445 ;
        RECT 134.490 136.325 134.660 136.475 ;
        RECT 133.905 135.945 134.235 136.305 ;
        RECT 134.490 136.115 135.790 136.325 ;
        RECT 136.065 135.945 136.520 136.710 ;
        RECT 138.305 136.695 138.825 137.235 ;
        RECT 137.615 135.945 138.825 136.695 ;
        RECT 13.330 135.775 138.910 135.945 ;
        RECT 13.415 135.025 14.625 135.775 ;
        RECT 13.415 134.485 13.935 135.025 ;
        RECT 14.795 134.975 15.105 135.775 ;
        RECT 15.310 134.975 16.005 135.605 ;
        RECT 16.265 135.225 16.435 135.515 ;
        RECT 16.605 135.395 16.935 135.775 ;
        RECT 16.265 135.055 16.930 135.225 ;
        RECT 14.105 134.315 14.625 134.855 ;
        RECT 14.805 134.535 15.140 134.805 ;
        RECT 15.310 134.375 15.480 134.975 ;
        RECT 15.650 134.535 15.985 134.785 ;
        RECT 13.415 133.225 14.625 134.315 ;
        RECT 14.795 133.225 15.075 134.365 ;
        RECT 15.245 133.395 15.575 134.375 ;
        RECT 15.745 133.225 16.005 134.365 ;
        RECT 16.180 134.235 16.530 134.885 ;
        RECT 16.700 134.065 16.930 135.055 ;
        RECT 16.265 133.895 16.930 134.065 ;
        RECT 16.265 133.395 16.435 133.895 ;
        RECT 16.605 133.225 16.935 133.725 ;
        RECT 17.105 133.395 17.290 135.515 ;
        RECT 17.545 135.315 17.795 135.775 ;
        RECT 17.965 135.325 18.300 135.495 ;
        RECT 18.495 135.325 19.170 135.495 ;
        RECT 17.965 135.185 18.135 135.325 ;
        RECT 17.460 134.195 17.740 135.145 ;
        RECT 17.910 135.055 18.135 135.185 ;
        RECT 17.910 133.950 18.080 135.055 ;
        RECT 18.305 134.905 18.830 135.125 ;
        RECT 18.250 134.140 18.490 134.735 ;
        RECT 18.660 134.205 18.830 134.905 ;
        RECT 19.000 134.545 19.170 135.325 ;
        RECT 19.490 135.275 19.860 135.775 ;
        RECT 20.040 135.325 20.445 135.495 ;
        RECT 20.615 135.325 21.400 135.495 ;
        RECT 20.040 135.095 20.210 135.325 ;
        RECT 19.380 134.795 20.210 135.095 ;
        RECT 20.595 134.825 21.060 135.155 ;
        RECT 19.380 134.765 19.580 134.795 ;
        RECT 19.700 134.545 19.870 134.615 ;
        RECT 19.000 134.375 19.870 134.545 ;
        RECT 19.360 134.285 19.870 134.375 ;
        RECT 17.910 133.820 18.215 133.950 ;
        RECT 18.660 133.840 19.190 134.205 ;
        RECT 17.530 133.225 17.795 133.685 ;
        RECT 17.965 133.395 18.215 133.820 ;
        RECT 19.360 133.670 19.530 134.285 ;
        RECT 18.425 133.500 19.530 133.670 ;
        RECT 19.700 133.225 19.870 134.025 ;
        RECT 20.040 133.725 20.210 134.795 ;
        RECT 20.380 133.895 20.570 134.615 ;
        RECT 20.740 133.865 21.060 134.825 ;
        RECT 21.230 134.865 21.400 135.325 ;
        RECT 21.675 135.245 21.885 135.775 ;
        RECT 22.145 135.035 22.475 135.560 ;
        RECT 22.645 135.165 22.815 135.775 ;
        RECT 22.985 135.120 23.315 135.555 ;
        RECT 23.535 135.125 23.795 135.605 ;
        RECT 23.965 135.235 24.215 135.775 ;
        RECT 22.985 135.035 23.365 135.120 ;
        RECT 22.275 134.865 22.475 135.035 ;
        RECT 23.140 134.995 23.365 135.035 ;
        RECT 21.230 134.535 22.105 134.865 ;
        RECT 22.275 134.535 23.025 134.865 ;
        RECT 20.040 133.395 20.290 133.725 ;
        RECT 21.230 133.695 21.400 134.535 ;
        RECT 22.275 134.330 22.465 134.535 ;
        RECT 23.195 134.415 23.365 134.995 ;
        RECT 23.150 134.365 23.365 134.415 ;
        RECT 21.570 133.955 22.465 134.330 ;
        RECT 22.975 134.285 23.365 134.365 ;
        RECT 20.515 133.525 21.400 133.695 ;
        RECT 21.580 133.225 21.895 133.725 ;
        RECT 22.125 133.395 22.465 133.955 ;
        RECT 22.635 133.225 22.805 134.235 ;
        RECT 22.975 133.440 23.305 134.285 ;
        RECT 23.535 134.095 23.705 135.125 ;
        RECT 24.385 135.070 24.605 135.555 ;
        RECT 23.875 134.475 24.105 134.870 ;
        RECT 24.275 134.645 24.605 135.070 ;
        RECT 24.775 135.395 25.665 135.565 ;
        RECT 24.775 134.670 24.945 135.395 ;
        RECT 25.920 135.275 26.415 135.605 ;
        RECT 25.115 134.840 25.665 135.225 ;
        RECT 24.775 134.600 25.665 134.670 ;
        RECT 24.770 134.575 25.665 134.600 ;
        RECT 24.760 134.560 25.665 134.575 ;
        RECT 24.755 134.545 25.665 134.560 ;
        RECT 24.745 134.540 25.665 134.545 ;
        RECT 24.740 134.530 25.665 134.540 ;
        RECT 24.735 134.520 25.665 134.530 ;
        RECT 24.725 134.515 25.665 134.520 ;
        RECT 24.715 134.505 25.665 134.515 ;
        RECT 24.705 134.500 25.665 134.505 ;
        RECT 24.705 134.495 25.040 134.500 ;
        RECT 24.690 134.490 25.040 134.495 ;
        RECT 24.675 134.480 25.040 134.490 ;
        RECT 24.650 134.475 25.040 134.480 ;
        RECT 23.875 134.470 25.040 134.475 ;
        RECT 23.875 134.435 25.010 134.470 ;
        RECT 23.875 134.410 24.975 134.435 ;
        RECT 23.875 134.380 24.945 134.410 ;
        RECT 23.875 134.350 24.925 134.380 ;
        RECT 23.875 134.320 24.905 134.350 ;
        RECT 23.875 134.310 24.835 134.320 ;
        RECT 23.875 134.300 24.810 134.310 ;
        RECT 23.875 134.285 24.790 134.300 ;
        RECT 23.875 134.270 24.770 134.285 ;
        RECT 23.980 134.260 24.765 134.270 ;
        RECT 23.980 134.225 24.750 134.260 ;
        RECT 23.535 133.395 23.810 134.095 ;
        RECT 23.980 133.975 24.735 134.225 ;
        RECT 24.905 133.905 25.235 134.150 ;
        RECT 25.405 134.050 25.665 134.500 ;
        RECT 25.050 133.880 25.235 133.905 ;
        RECT 25.050 133.780 25.665 133.880 ;
        RECT 25.835 133.785 26.075 135.095 ;
        RECT 26.245 134.365 26.415 135.275 ;
        RECT 26.635 134.535 26.985 135.500 ;
        RECT 27.165 134.535 27.465 135.505 ;
        RECT 27.645 134.535 27.925 135.505 ;
        RECT 28.105 134.975 28.375 135.775 ;
        RECT 28.545 135.055 28.885 135.565 ;
        RECT 28.120 134.535 28.450 134.785 ;
        RECT 28.120 134.365 28.435 134.535 ;
        RECT 26.245 134.195 28.435 134.365 ;
        RECT 23.980 133.225 24.235 133.770 ;
        RECT 24.405 133.395 24.885 133.735 ;
        RECT 25.060 133.225 25.665 133.780 ;
        RECT 25.840 133.225 26.175 133.605 ;
        RECT 26.345 133.395 26.595 134.195 ;
        RECT 26.815 133.225 27.145 133.945 ;
        RECT 27.330 133.395 27.580 134.195 ;
        RECT 28.045 133.225 28.375 134.025 ;
        RECT 28.625 133.655 28.885 135.055 ;
        RECT 29.065 135.045 29.365 135.775 ;
        RECT 29.545 134.865 29.775 135.485 ;
        RECT 29.975 135.215 30.200 135.595 ;
        RECT 30.370 135.385 30.700 135.775 ;
        RECT 29.975 135.035 30.305 135.215 ;
        RECT 29.070 134.535 29.365 134.865 ;
        RECT 29.545 134.535 29.960 134.865 ;
        RECT 30.130 134.365 30.305 135.035 ;
        RECT 30.475 134.535 30.715 135.185 ;
        RECT 30.895 135.145 31.235 135.605 ;
        RECT 31.405 135.315 31.575 135.775 ;
        RECT 32.205 135.340 32.565 135.605 ;
        RECT 32.210 135.335 32.565 135.340 ;
        RECT 32.215 135.325 32.565 135.335 ;
        RECT 32.220 135.320 32.565 135.325 ;
        RECT 32.225 135.310 32.565 135.320 ;
        RECT 32.805 135.315 32.975 135.775 ;
        RECT 32.230 135.305 32.565 135.310 ;
        RECT 32.240 135.295 32.565 135.305 ;
        RECT 32.250 135.285 32.565 135.295 ;
        RECT 31.745 135.145 32.075 135.225 ;
        RECT 30.895 134.955 32.075 135.145 ;
        RECT 32.265 135.145 32.565 135.285 ;
        RECT 32.265 134.955 32.975 135.145 ;
        RECT 30.895 134.585 31.225 134.785 ;
        RECT 31.535 134.765 31.865 134.785 ;
        RECT 31.415 134.585 31.865 134.765 ;
        RECT 28.545 133.395 28.885 133.655 ;
        RECT 29.065 134.005 29.960 134.335 ;
        RECT 30.130 134.175 30.715 134.365 ;
        RECT 30.895 134.245 31.125 134.585 ;
        RECT 29.065 133.835 30.270 134.005 ;
        RECT 29.065 133.405 29.395 133.835 ;
        RECT 29.575 133.225 29.770 133.665 ;
        RECT 29.940 133.405 30.270 133.835 ;
        RECT 30.440 133.405 30.715 134.175 ;
        RECT 30.905 133.225 31.235 133.945 ;
        RECT 31.415 133.470 31.630 134.585 ;
        RECT 32.035 134.555 32.505 134.785 ;
        RECT 32.690 134.385 32.975 134.955 ;
        RECT 33.145 134.830 33.485 135.605 ;
        RECT 33.655 135.165 33.995 135.580 ;
        RECT 34.165 135.335 34.335 135.775 ;
        RECT 34.505 135.385 35.755 135.565 ;
        RECT 34.505 135.165 34.835 135.385 ;
        RECT 36.025 135.315 36.195 135.775 ;
        RECT 33.655 134.995 34.835 135.165 ;
        RECT 35.005 135.145 35.370 135.215 ;
        RECT 35.005 134.965 36.255 135.145 ;
        RECT 31.825 134.170 32.975 134.385 ;
        RECT 31.825 133.395 32.155 134.170 ;
        RECT 32.325 133.225 33.035 134.000 ;
        RECT 33.205 133.395 33.485 134.830 ;
        RECT 33.655 134.585 34.120 134.785 ;
        RECT 34.295 134.535 34.625 134.785 ;
        RECT 34.795 134.755 35.260 134.785 ;
        RECT 34.795 134.585 35.265 134.755 ;
        RECT 34.795 134.535 35.260 134.585 ;
        RECT 35.455 134.535 35.810 134.785 ;
        RECT 34.295 134.415 34.475 134.535 ;
        RECT 33.655 133.225 33.975 134.405 ;
        RECT 34.145 134.245 34.475 134.415 ;
        RECT 35.980 134.365 36.255 134.965 ;
        RECT 34.145 133.455 34.345 134.245 ;
        RECT 34.645 134.155 36.255 134.365 ;
        RECT 34.645 134.055 35.055 134.155 ;
        RECT 34.670 133.395 35.055 134.055 ;
        RECT 35.450 133.225 36.235 133.985 ;
        RECT 36.425 133.395 36.705 135.495 ;
        RECT 36.875 135.005 38.545 135.775 ;
        RECT 39.175 135.050 39.465 135.775 ;
        RECT 39.635 135.230 44.980 135.775 ;
        RECT 46.160 135.275 46.655 135.605 ;
        RECT 36.875 134.485 37.625 135.005 ;
        RECT 37.795 134.315 38.545 134.835 ;
        RECT 41.220 134.400 41.560 135.230 ;
        RECT 36.875 133.225 38.545 134.315 ;
        RECT 39.175 133.225 39.465 134.390 ;
        RECT 43.040 133.660 43.390 134.910 ;
        RECT 46.075 133.785 46.315 135.095 ;
        RECT 46.485 134.365 46.655 135.275 ;
        RECT 46.875 134.535 47.225 135.500 ;
        RECT 47.405 134.535 47.705 135.505 ;
        RECT 47.885 134.535 48.165 135.505 ;
        RECT 48.345 134.975 48.615 135.775 ;
        RECT 48.785 135.055 49.125 135.565 ;
        RECT 49.345 135.120 49.675 135.555 ;
        RECT 49.845 135.165 50.015 135.775 ;
        RECT 48.360 134.535 48.690 134.785 ;
        RECT 48.360 134.365 48.675 134.535 ;
        RECT 46.485 134.195 48.675 134.365 ;
        RECT 39.635 133.225 44.980 133.660 ;
        RECT 46.080 133.225 46.415 133.605 ;
        RECT 46.585 133.395 46.835 134.195 ;
        RECT 47.055 133.225 47.385 133.945 ;
        RECT 47.570 133.395 47.820 134.195 ;
        RECT 48.285 133.225 48.615 134.025 ;
        RECT 48.865 133.655 49.125 135.055 ;
        RECT 49.295 135.035 49.675 135.120 ;
        RECT 50.185 135.035 50.515 135.560 ;
        RECT 50.775 135.245 50.985 135.775 ;
        RECT 51.260 135.325 52.045 135.495 ;
        RECT 52.215 135.325 52.620 135.495 ;
        RECT 49.295 134.995 49.520 135.035 ;
        RECT 49.295 134.415 49.465 134.995 ;
        RECT 50.185 134.865 50.385 135.035 ;
        RECT 51.260 134.865 51.430 135.325 ;
        RECT 49.635 134.535 50.385 134.865 ;
        RECT 50.555 134.535 51.430 134.865 ;
        RECT 49.295 134.365 49.510 134.415 ;
        RECT 49.295 134.285 49.685 134.365 ;
        RECT 48.785 133.395 49.125 133.655 ;
        RECT 49.355 133.440 49.685 134.285 ;
        RECT 50.195 134.330 50.385 134.535 ;
        RECT 49.855 133.225 50.025 134.235 ;
        RECT 50.195 133.955 51.090 134.330 ;
        RECT 50.195 133.395 50.535 133.955 ;
        RECT 50.765 133.225 51.080 133.725 ;
        RECT 51.260 133.695 51.430 134.535 ;
        RECT 51.600 134.825 52.065 135.155 ;
        RECT 52.450 135.095 52.620 135.325 ;
        RECT 52.800 135.275 53.170 135.775 ;
        RECT 53.490 135.325 54.165 135.495 ;
        RECT 54.360 135.325 54.695 135.495 ;
        RECT 51.600 133.865 51.920 134.825 ;
        RECT 52.450 134.795 53.280 135.095 ;
        RECT 52.090 133.895 52.280 134.615 ;
        RECT 52.450 133.725 52.620 134.795 ;
        RECT 53.080 134.765 53.280 134.795 ;
        RECT 52.790 134.545 52.960 134.615 ;
        RECT 53.490 134.545 53.660 135.325 ;
        RECT 54.525 135.185 54.695 135.325 ;
        RECT 54.865 135.315 55.115 135.775 ;
        RECT 52.790 134.375 53.660 134.545 ;
        RECT 53.830 134.905 54.355 135.125 ;
        RECT 54.525 135.055 54.750 135.185 ;
        RECT 52.790 134.285 53.300 134.375 ;
        RECT 51.260 133.525 52.145 133.695 ;
        RECT 52.370 133.395 52.620 133.725 ;
        RECT 52.790 133.225 52.960 134.025 ;
        RECT 53.130 133.670 53.300 134.285 ;
        RECT 53.830 134.205 54.000 134.905 ;
        RECT 53.470 133.840 54.000 134.205 ;
        RECT 54.170 134.140 54.410 134.735 ;
        RECT 54.580 133.950 54.750 135.055 ;
        RECT 54.920 134.195 55.200 135.145 ;
        RECT 54.445 133.820 54.750 133.950 ;
        RECT 53.130 133.500 54.235 133.670 ;
        RECT 54.445 133.395 54.695 133.820 ;
        RECT 54.865 133.225 55.130 133.685 ;
        RECT 55.370 133.395 55.555 135.515 ;
        RECT 55.725 135.395 56.055 135.775 ;
        RECT 56.225 135.225 56.395 135.515 ;
        RECT 56.655 135.230 62.000 135.775 ;
        RECT 55.730 135.055 56.395 135.225 ;
        RECT 55.730 134.065 55.960 135.055 ;
        RECT 56.130 134.235 56.480 134.885 ;
        RECT 58.240 134.400 58.580 135.230 ;
        RECT 62.175 135.005 64.765 135.775 ;
        RECT 64.935 135.050 65.225 135.775 ;
        RECT 65.485 135.225 65.655 135.515 ;
        RECT 65.825 135.395 66.155 135.775 ;
        RECT 65.485 135.055 66.150 135.225 ;
        RECT 55.730 133.895 56.395 134.065 ;
        RECT 55.725 133.225 56.055 133.725 ;
        RECT 56.225 133.395 56.395 133.895 ;
        RECT 60.060 133.660 60.410 134.910 ;
        RECT 62.175 134.485 63.385 135.005 ;
        RECT 63.555 134.315 64.765 134.835 ;
        RECT 56.655 133.225 62.000 133.660 ;
        RECT 62.175 133.225 64.765 134.315 ;
        RECT 64.935 133.225 65.225 134.390 ;
        RECT 65.400 134.235 65.750 134.885 ;
        RECT 65.920 134.065 66.150 135.055 ;
        RECT 65.485 133.895 66.150 134.065 ;
        RECT 65.485 133.395 65.655 133.895 ;
        RECT 65.825 133.225 66.155 133.725 ;
        RECT 66.325 133.395 66.510 135.515 ;
        RECT 66.765 135.315 67.015 135.775 ;
        RECT 67.185 135.325 67.520 135.495 ;
        RECT 67.715 135.325 68.390 135.495 ;
        RECT 67.185 135.185 67.355 135.325 ;
        RECT 66.680 134.195 66.960 135.145 ;
        RECT 67.130 135.055 67.355 135.185 ;
        RECT 67.130 133.950 67.300 135.055 ;
        RECT 67.525 134.905 68.050 135.125 ;
        RECT 67.470 134.140 67.710 134.735 ;
        RECT 67.880 134.205 68.050 134.905 ;
        RECT 68.220 134.545 68.390 135.325 ;
        RECT 68.710 135.275 69.080 135.775 ;
        RECT 69.260 135.325 69.665 135.495 ;
        RECT 69.835 135.325 70.620 135.495 ;
        RECT 69.260 135.095 69.430 135.325 ;
        RECT 68.600 134.795 69.430 135.095 ;
        RECT 69.815 134.825 70.280 135.155 ;
        RECT 68.600 134.765 68.800 134.795 ;
        RECT 68.920 134.545 69.090 134.615 ;
        RECT 68.220 134.375 69.090 134.545 ;
        RECT 68.580 134.285 69.090 134.375 ;
        RECT 67.130 133.820 67.435 133.950 ;
        RECT 67.880 133.840 68.410 134.205 ;
        RECT 66.750 133.225 67.015 133.685 ;
        RECT 67.185 133.395 67.435 133.820 ;
        RECT 68.580 133.670 68.750 134.285 ;
        RECT 67.645 133.500 68.750 133.670 ;
        RECT 68.920 133.225 69.090 134.025 ;
        RECT 69.260 133.725 69.430 134.795 ;
        RECT 69.600 133.895 69.790 134.615 ;
        RECT 69.960 133.865 70.280 134.825 ;
        RECT 70.450 134.865 70.620 135.325 ;
        RECT 70.895 135.245 71.105 135.775 ;
        RECT 71.365 135.035 71.695 135.560 ;
        RECT 71.865 135.165 72.035 135.775 ;
        RECT 72.205 135.120 72.535 135.555 ;
        RECT 72.205 135.035 72.585 135.120 ;
        RECT 71.495 134.865 71.695 135.035 ;
        RECT 72.360 134.995 72.585 135.035 ;
        RECT 70.450 134.535 71.325 134.865 ;
        RECT 71.495 134.535 72.245 134.865 ;
        RECT 69.260 133.395 69.510 133.725 ;
        RECT 70.450 133.695 70.620 134.535 ;
        RECT 71.495 134.330 71.685 134.535 ;
        RECT 72.415 134.415 72.585 134.995 ;
        RECT 72.775 134.965 73.015 135.775 ;
        RECT 73.185 134.965 73.515 135.605 ;
        RECT 73.685 134.965 73.955 135.775 ;
        RECT 72.755 134.535 73.105 134.785 ;
        RECT 72.370 134.365 72.585 134.415 ;
        RECT 73.275 134.365 73.445 134.965 ;
        RECT 74.135 134.955 74.395 135.775 ;
        RECT 74.565 134.955 74.895 135.375 ;
        RECT 75.075 135.290 75.865 135.555 ;
        RECT 74.645 134.865 74.895 134.955 ;
        RECT 73.615 134.535 73.965 134.785 ;
        RECT 70.790 133.955 71.685 134.330 ;
        RECT 72.195 134.285 72.585 134.365 ;
        RECT 69.735 133.525 70.620 133.695 ;
        RECT 70.800 133.225 71.115 133.725 ;
        RECT 71.345 133.395 71.685 133.955 ;
        RECT 71.855 133.225 72.025 134.235 ;
        RECT 72.195 133.440 72.525 134.285 ;
        RECT 72.765 134.195 73.445 134.365 ;
        RECT 72.765 133.410 73.095 134.195 ;
        RECT 73.625 133.225 73.955 134.365 ;
        RECT 74.135 133.905 74.475 134.785 ;
        RECT 74.645 134.615 75.440 134.865 ;
        RECT 74.135 133.225 74.395 133.735 ;
        RECT 74.645 133.395 74.815 134.615 ;
        RECT 75.610 134.435 75.865 135.290 ;
        RECT 76.035 135.135 76.235 135.555 ;
        RECT 76.425 135.315 76.755 135.775 ;
        RECT 76.035 134.615 76.445 135.135 ;
        RECT 76.925 135.125 77.185 135.605 ;
        RECT 76.615 134.435 76.845 134.865 ;
        RECT 75.055 134.265 76.845 134.435 ;
        RECT 75.055 133.900 75.305 134.265 ;
        RECT 75.475 133.905 75.805 134.095 ;
        RECT 76.025 133.970 76.740 134.265 ;
        RECT 77.015 134.095 77.185 135.125 ;
        RECT 77.630 134.965 77.875 135.570 ;
        RECT 78.095 135.240 78.605 135.775 ;
        RECT 75.475 133.730 75.670 133.905 ;
        RECT 75.055 133.225 75.670 133.730 ;
        RECT 75.840 133.395 76.315 133.735 ;
        RECT 76.485 133.225 76.700 133.770 ;
        RECT 76.910 133.395 77.185 134.095 ;
        RECT 77.355 134.795 78.585 134.965 ;
        RECT 77.355 133.985 77.695 134.795 ;
        RECT 77.865 134.230 78.615 134.420 ;
        RECT 77.355 133.575 77.870 133.985 ;
        RECT 78.105 133.225 78.275 133.985 ;
        RECT 78.445 133.565 78.615 134.230 ;
        RECT 78.785 134.245 78.975 135.605 ;
        RECT 79.145 134.755 79.420 135.605 ;
        RECT 79.610 135.240 80.140 135.605 ;
        RECT 80.565 135.375 80.895 135.775 ;
        RECT 79.965 135.205 80.140 135.240 ;
        RECT 79.145 134.585 79.425 134.755 ;
        RECT 79.145 134.445 79.420 134.585 ;
        RECT 79.625 134.245 79.795 135.045 ;
        RECT 78.785 134.075 79.795 134.245 ;
        RECT 79.965 135.035 80.895 135.205 ;
        RECT 81.065 135.035 81.320 135.605 ;
        RECT 81.585 135.225 81.755 135.515 ;
        RECT 81.925 135.395 82.255 135.775 ;
        RECT 81.585 135.055 82.250 135.225 ;
        RECT 79.965 133.905 80.135 135.035 ;
        RECT 80.725 134.865 80.895 135.035 ;
        RECT 79.010 133.735 80.135 133.905 ;
        RECT 80.305 134.535 80.500 134.865 ;
        RECT 80.725 134.535 80.980 134.865 ;
        RECT 80.305 133.565 80.475 134.535 ;
        RECT 81.150 134.365 81.320 135.035 ;
        RECT 78.445 133.395 80.475 133.565 ;
        RECT 80.645 133.225 80.815 134.365 ;
        RECT 80.985 133.395 81.320 134.365 ;
        RECT 81.500 134.235 81.850 134.885 ;
        RECT 82.020 134.065 82.250 135.055 ;
        RECT 81.585 133.895 82.250 134.065 ;
        RECT 81.585 133.395 81.755 133.895 ;
        RECT 81.925 133.225 82.255 133.725 ;
        RECT 82.425 133.395 82.610 135.515 ;
        RECT 82.865 135.315 83.115 135.775 ;
        RECT 83.285 135.325 83.620 135.495 ;
        RECT 83.815 135.325 84.490 135.495 ;
        RECT 83.285 135.185 83.455 135.325 ;
        RECT 82.780 134.195 83.060 135.145 ;
        RECT 83.230 135.055 83.455 135.185 ;
        RECT 83.230 133.950 83.400 135.055 ;
        RECT 83.625 134.905 84.150 135.125 ;
        RECT 83.570 134.140 83.810 134.735 ;
        RECT 83.980 134.205 84.150 134.905 ;
        RECT 84.320 134.545 84.490 135.325 ;
        RECT 84.810 135.275 85.180 135.775 ;
        RECT 85.360 135.325 85.765 135.495 ;
        RECT 85.935 135.325 86.720 135.495 ;
        RECT 85.360 135.095 85.530 135.325 ;
        RECT 84.700 134.795 85.530 135.095 ;
        RECT 85.915 134.825 86.380 135.155 ;
        RECT 84.700 134.765 84.900 134.795 ;
        RECT 85.020 134.545 85.190 134.615 ;
        RECT 84.320 134.375 85.190 134.545 ;
        RECT 84.680 134.285 85.190 134.375 ;
        RECT 83.230 133.820 83.535 133.950 ;
        RECT 83.980 133.840 84.510 134.205 ;
        RECT 82.850 133.225 83.115 133.685 ;
        RECT 83.285 133.395 83.535 133.820 ;
        RECT 84.680 133.670 84.850 134.285 ;
        RECT 83.745 133.500 84.850 133.670 ;
        RECT 85.020 133.225 85.190 134.025 ;
        RECT 85.360 133.725 85.530 134.795 ;
        RECT 85.700 133.895 85.890 134.615 ;
        RECT 86.060 133.865 86.380 134.825 ;
        RECT 86.550 134.865 86.720 135.325 ;
        RECT 86.995 135.245 87.205 135.775 ;
        RECT 87.465 135.035 87.795 135.560 ;
        RECT 87.965 135.165 88.135 135.775 ;
        RECT 88.305 135.120 88.635 135.555 ;
        RECT 88.805 135.260 88.975 135.775 ;
        RECT 88.305 135.035 88.685 135.120 ;
        RECT 87.595 134.865 87.795 135.035 ;
        RECT 88.460 134.995 88.685 135.035 ;
        RECT 86.550 134.535 87.425 134.865 ;
        RECT 87.595 134.535 88.345 134.865 ;
        RECT 85.360 133.395 85.610 133.725 ;
        RECT 86.550 133.695 86.720 134.535 ;
        RECT 87.595 134.330 87.785 134.535 ;
        RECT 88.515 134.415 88.685 134.995 ;
        RECT 89.315 135.025 90.525 135.775 ;
        RECT 90.695 135.050 90.985 135.775 ;
        RECT 89.315 134.485 89.835 135.025 ;
        RECT 91.155 135.005 92.825 135.775 ;
        RECT 93.085 135.225 93.255 135.515 ;
        RECT 93.425 135.395 93.755 135.775 ;
        RECT 93.085 135.055 93.750 135.225 ;
        RECT 88.470 134.365 88.685 134.415 ;
        RECT 86.890 133.955 87.785 134.330 ;
        RECT 88.295 134.285 88.685 134.365 ;
        RECT 90.005 134.315 90.525 134.855 ;
        RECT 91.155 134.485 91.905 135.005 ;
        RECT 85.835 133.525 86.720 133.695 ;
        RECT 86.900 133.225 87.215 133.725 ;
        RECT 87.445 133.395 87.785 133.955 ;
        RECT 87.955 133.225 88.125 134.235 ;
        RECT 88.295 133.440 88.625 134.285 ;
        RECT 88.795 133.225 88.965 134.140 ;
        RECT 89.315 133.225 90.525 134.315 ;
        RECT 90.695 133.225 90.985 134.390 ;
        RECT 92.075 134.315 92.825 134.835 ;
        RECT 91.155 133.225 92.825 134.315 ;
        RECT 93.000 134.235 93.350 134.885 ;
        RECT 93.520 134.065 93.750 135.055 ;
        RECT 93.085 133.895 93.750 134.065 ;
        RECT 93.085 133.395 93.255 133.895 ;
        RECT 93.425 133.225 93.755 133.725 ;
        RECT 93.925 133.395 94.110 135.515 ;
        RECT 94.365 135.315 94.615 135.775 ;
        RECT 94.785 135.325 95.120 135.495 ;
        RECT 95.315 135.325 95.990 135.495 ;
        RECT 94.785 135.185 94.955 135.325 ;
        RECT 94.280 134.195 94.560 135.145 ;
        RECT 94.730 135.055 94.955 135.185 ;
        RECT 94.730 133.950 94.900 135.055 ;
        RECT 95.125 134.905 95.650 135.125 ;
        RECT 95.070 134.140 95.310 134.735 ;
        RECT 95.480 134.205 95.650 134.905 ;
        RECT 95.820 134.545 95.990 135.325 ;
        RECT 96.310 135.275 96.680 135.775 ;
        RECT 96.860 135.325 97.265 135.495 ;
        RECT 97.435 135.325 98.220 135.495 ;
        RECT 96.860 135.095 97.030 135.325 ;
        RECT 96.200 134.795 97.030 135.095 ;
        RECT 97.415 134.825 97.880 135.155 ;
        RECT 96.200 134.765 96.400 134.795 ;
        RECT 96.520 134.545 96.690 134.615 ;
        RECT 95.820 134.375 96.690 134.545 ;
        RECT 96.180 134.285 96.690 134.375 ;
        RECT 94.730 133.820 95.035 133.950 ;
        RECT 95.480 133.840 96.010 134.205 ;
        RECT 94.350 133.225 94.615 133.685 ;
        RECT 94.785 133.395 95.035 133.820 ;
        RECT 96.180 133.670 96.350 134.285 ;
        RECT 95.245 133.500 96.350 133.670 ;
        RECT 96.520 133.225 96.690 134.025 ;
        RECT 96.860 133.725 97.030 134.795 ;
        RECT 97.200 133.895 97.390 134.615 ;
        RECT 97.560 133.865 97.880 134.825 ;
        RECT 98.050 134.865 98.220 135.325 ;
        RECT 98.495 135.245 98.705 135.775 ;
        RECT 98.965 135.035 99.295 135.560 ;
        RECT 99.465 135.165 99.635 135.775 ;
        RECT 99.805 135.120 100.135 135.555 ;
        RECT 99.805 135.035 100.185 135.120 ;
        RECT 99.095 134.865 99.295 135.035 ;
        RECT 99.960 134.995 100.185 135.035 ;
        RECT 98.050 134.535 98.925 134.865 ;
        RECT 99.095 134.535 99.845 134.865 ;
        RECT 96.860 133.395 97.110 133.725 ;
        RECT 98.050 133.695 98.220 134.535 ;
        RECT 99.095 134.330 99.285 134.535 ;
        RECT 100.015 134.415 100.185 134.995 ;
        RECT 99.970 134.365 100.185 134.415 ;
        RECT 98.390 133.955 99.285 134.330 ;
        RECT 99.795 134.285 100.185 134.365 ;
        RECT 100.360 135.035 100.615 135.605 ;
        RECT 100.785 135.375 101.115 135.775 ;
        RECT 101.540 135.240 102.070 135.605 ;
        RECT 101.540 135.205 101.715 135.240 ;
        RECT 100.785 135.035 101.715 135.205 ;
        RECT 100.360 134.365 100.530 135.035 ;
        RECT 100.785 134.865 100.955 135.035 ;
        RECT 100.700 134.535 100.955 134.865 ;
        RECT 101.180 134.535 101.375 134.865 ;
        RECT 97.335 133.525 98.220 133.695 ;
        RECT 98.400 133.225 98.715 133.725 ;
        RECT 98.945 133.395 99.285 133.955 ;
        RECT 99.455 133.225 99.625 134.235 ;
        RECT 99.795 133.440 100.125 134.285 ;
        RECT 100.360 133.395 100.695 134.365 ;
        RECT 100.865 133.225 101.035 134.365 ;
        RECT 101.205 133.565 101.375 134.535 ;
        RECT 101.545 133.905 101.715 135.035 ;
        RECT 101.885 134.245 102.055 135.045 ;
        RECT 102.260 134.755 102.535 135.605 ;
        RECT 102.255 134.585 102.535 134.755 ;
        RECT 102.260 134.445 102.535 134.585 ;
        RECT 102.705 134.245 102.895 135.605 ;
        RECT 103.075 135.240 103.585 135.775 ;
        RECT 103.805 134.965 104.050 135.570 ;
        RECT 104.495 135.025 105.705 135.775 ;
        RECT 105.965 135.225 106.135 135.515 ;
        RECT 106.305 135.395 106.635 135.775 ;
        RECT 105.965 135.055 106.630 135.225 ;
        RECT 103.095 134.795 104.325 134.965 ;
        RECT 101.885 134.075 102.895 134.245 ;
        RECT 103.065 134.230 103.815 134.420 ;
        RECT 101.545 133.735 102.670 133.905 ;
        RECT 103.065 133.565 103.235 134.230 ;
        RECT 103.985 133.985 104.325 134.795 ;
        RECT 104.495 134.485 105.015 135.025 ;
        RECT 105.185 134.315 105.705 134.855 ;
        RECT 101.205 133.395 103.235 133.565 ;
        RECT 103.405 133.225 103.575 133.985 ;
        RECT 103.810 133.575 104.325 133.985 ;
        RECT 104.495 133.225 105.705 134.315 ;
        RECT 105.880 134.235 106.230 134.885 ;
        RECT 106.400 134.065 106.630 135.055 ;
        RECT 105.965 133.895 106.630 134.065 ;
        RECT 105.965 133.395 106.135 133.895 ;
        RECT 106.305 133.225 106.635 133.725 ;
        RECT 106.805 133.395 106.990 135.515 ;
        RECT 107.245 135.315 107.495 135.775 ;
        RECT 107.665 135.325 108.000 135.495 ;
        RECT 108.195 135.325 108.870 135.495 ;
        RECT 107.665 135.185 107.835 135.325 ;
        RECT 107.160 134.195 107.440 135.145 ;
        RECT 107.610 135.055 107.835 135.185 ;
        RECT 107.610 133.950 107.780 135.055 ;
        RECT 108.005 134.905 108.530 135.125 ;
        RECT 107.950 134.140 108.190 134.735 ;
        RECT 108.360 134.205 108.530 134.905 ;
        RECT 108.700 134.545 108.870 135.325 ;
        RECT 109.190 135.275 109.560 135.775 ;
        RECT 109.740 135.325 110.145 135.495 ;
        RECT 110.315 135.325 111.100 135.495 ;
        RECT 109.740 135.095 109.910 135.325 ;
        RECT 109.080 134.795 109.910 135.095 ;
        RECT 110.295 134.825 110.760 135.155 ;
        RECT 109.080 134.765 109.280 134.795 ;
        RECT 109.400 134.545 109.570 134.615 ;
        RECT 108.700 134.375 109.570 134.545 ;
        RECT 109.060 134.285 109.570 134.375 ;
        RECT 107.610 133.820 107.915 133.950 ;
        RECT 108.360 133.840 108.890 134.205 ;
        RECT 107.230 133.225 107.495 133.685 ;
        RECT 107.665 133.395 107.915 133.820 ;
        RECT 109.060 133.670 109.230 134.285 ;
        RECT 108.125 133.500 109.230 133.670 ;
        RECT 109.400 133.225 109.570 134.025 ;
        RECT 109.740 133.725 109.910 134.795 ;
        RECT 110.080 133.895 110.270 134.615 ;
        RECT 110.440 133.865 110.760 134.825 ;
        RECT 110.930 134.865 111.100 135.325 ;
        RECT 111.375 135.245 111.585 135.775 ;
        RECT 111.845 135.035 112.175 135.560 ;
        RECT 112.345 135.165 112.515 135.775 ;
        RECT 112.685 135.120 113.015 135.555 ;
        RECT 113.235 135.275 113.535 135.605 ;
        RECT 113.705 135.295 113.980 135.775 ;
        RECT 112.685 135.035 113.065 135.120 ;
        RECT 111.975 134.865 112.175 135.035 ;
        RECT 112.840 134.995 113.065 135.035 ;
        RECT 110.930 134.535 111.805 134.865 ;
        RECT 111.975 134.535 112.725 134.865 ;
        RECT 109.740 133.395 109.990 133.725 ;
        RECT 110.930 133.695 111.100 134.535 ;
        RECT 111.975 134.330 112.165 134.535 ;
        RECT 112.895 134.415 113.065 134.995 ;
        RECT 112.850 134.365 113.065 134.415 ;
        RECT 111.270 133.955 112.165 134.330 ;
        RECT 112.675 134.285 113.065 134.365 ;
        RECT 113.235 134.365 113.405 135.275 ;
        RECT 114.160 135.125 114.455 135.515 ;
        RECT 114.625 135.295 114.880 135.775 ;
        RECT 115.055 135.125 115.315 135.515 ;
        RECT 115.485 135.295 115.765 135.775 ;
        RECT 113.575 134.535 113.925 135.105 ;
        RECT 114.160 134.955 115.810 135.125 ;
        RECT 116.455 135.050 116.745 135.775 ;
        RECT 117.005 135.225 117.175 135.515 ;
        RECT 117.345 135.395 117.675 135.775 ;
        RECT 117.005 135.055 117.670 135.225 ;
        RECT 114.095 134.615 115.235 134.785 ;
        RECT 114.095 134.365 114.265 134.615 ;
        RECT 115.405 134.445 115.810 134.955 ;
        RECT 110.215 133.525 111.100 133.695 ;
        RECT 111.280 133.225 111.595 133.725 ;
        RECT 111.825 133.395 112.165 133.955 ;
        RECT 112.335 133.225 112.505 134.235 ;
        RECT 112.675 133.440 113.005 134.285 ;
        RECT 113.235 134.195 114.265 134.365 ;
        RECT 115.055 134.275 115.810 134.445 ;
        RECT 113.235 133.395 113.545 134.195 ;
        RECT 115.055 134.025 115.315 134.275 ;
        RECT 113.715 133.225 114.025 134.025 ;
        RECT 114.195 133.855 115.315 134.025 ;
        RECT 114.195 133.395 114.455 133.855 ;
        RECT 114.625 133.225 114.880 133.685 ;
        RECT 115.055 133.395 115.315 133.855 ;
        RECT 115.485 133.225 115.770 134.095 ;
        RECT 116.455 133.225 116.745 134.390 ;
        RECT 116.920 134.235 117.270 134.885 ;
        RECT 117.440 134.065 117.670 135.055 ;
        RECT 117.005 133.895 117.670 134.065 ;
        RECT 117.005 133.395 117.175 133.895 ;
        RECT 117.345 133.225 117.675 133.725 ;
        RECT 117.845 133.395 118.030 135.515 ;
        RECT 118.285 135.315 118.535 135.775 ;
        RECT 118.705 135.325 119.040 135.495 ;
        RECT 119.235 135.325 119.910 135.495 ;
        RECT 118.705 135.185 118.875 135.325 ;
        RECT 118.200 134.195 118.480 135.145 ;
        RECT 118.650 135.055 118.875 135.185 ;
        RECT 118.650 133.950 118.820 135.055 ;
        RECT 119.045 134.905 119.570 135.125 ;
        RECT 118.990 134.140 119.230 134.735 ;
        RECT 119.400 134.205 119.570 134.905 ;
        RECT 119.740 134.545 119.910 135.325 ;
        RECT 120.230 135.275 120.600 135.775 ;
        RECT 120.780 135.325 121.185 135.495 ;
        RECT 121.355 135.325 122.140 135.495 ;
        RECT 120.780 135.095 120.950 135.325 ;
        RECT 120.120 134.795 120.950 135.095 ;
        RECT 121.335 134.825 121.800 135.155 ;
        RECT 120.120 134.765 120.320 134.795 ;
        RECT 120.440 134.545 120.610 134.615 ;
        RECT 119.740 134.375 120.610 134.545 ;
        RECT 120.100 134.285 120.610 134.375 ;
        RECT 118.650 133.820 118.955 133.950 ;
        RECT 119.400 133.840 119.930 134.205 ;
        RECT 118.270 133.225 118.535 133.685 ;
        RECT 118.705 133.395 118.955 133.820 ;
        RECT 120.100 133.670 120.270 134.285 ;
        RECT 119.165 133.500 120.270 133.670 ;
        RECT 120.440 133.225 120.610 134.025 ;
        RECT 120.780 133.725 120.950 134.795 ;
        RECT 121.120 133.895 121.310 134.615 ;
        RECT 121.480 133.865 121.800 134.825 ;
        RECT 121.970 134.865 122.140 135.325 ;
        RECT 122.415 135.245 122.625 135.775 ;
        RECT 122.885 135.035 123.215 135.560 ;
        RECT 123.385 135.165 123.555 135.775 ;
        RECT 123.725 135.120 124.055 135.555 ;
        RECT 123.725 135.035 124.105 135.120 ;
        RECT 123.015 134.865 123.215 135.035 ;
        RECT 123.880 134.995 124.105 135.035 ;
        RECT 121.970 134.535 122.845 134.865 ;
        RECT 123.015 134.535 123.765 134.865 ;
        RECT 120.780 133.395 121.030 133.725 ;
        RECT 121.970 133.695 122.140 134.535 ;
        RECT 123.015 134.330 123.205 134.535 ;
        RECT 123.935 134.415 124.105 134.995 ;
        RECT 124.275 135.005 126.865 135.775 ;
        RECT 127.125 135.225 127.295 135.515 ;
        RECT 127.465 135.395 127.795 135.775 ;
        RECT 127.125 135.055 127.790 135.225 ;
        RECT 124.275 134.485 125.485 135.005 ;
        RECT 123.890 134.365 124.105 134.415 ;
        RECT 122.310 133.955 123.205 134.330 ;
        RECT 123.715 134.285 124.105 134.365 ;
        RECT 125.655 134.315 126.865 134.835 ;
        RECT 121.255 133.525 122.140 133.695 ;
        RECT 122.320 133.225 122.635 133.725 ;
        RECT 122.865 133.395 123.205 133.955 ;
        RECT 123.375 133.225 123.545 134.235 ;
        RECT 123.715 133.440 124.045 134.285 ;
        RECT 124.275 133.225 126.865 134.315 ;
        RECT 127.040 134.235 127.390 134.885 ;
        RECT 127.560 134.065 127.790 135.055 ;
        RECT 127.125 133.895 127.790 134.065 ;
        RECT 127.125 133.395 127.295 133.895 ;
        RECT 127.465 133.225 127.795 133.725 ;
        RECT 127.965 133.395 128.150 135.515 ;
        RECT 128.405 135.315 128.655 135.775 ;
        RECT 128.825 135.325 129.160 135.495 ;
        RECT 129.355 135.325 130.030 135.495 ;
        RECT 128.825 135.185 128.995 135.325 ;
        RECT 128.320 134.195 128.600 135.145 ;
        RECT 128.770 135.055 128.995 135.185 ;
        RECT 128.770 133.950 128.940 135.055 ;
        RECT 129.165 134.905 129.690 135.125 ;
        RECT 129.110 134.140 129.350 134.735 ;
        RECT 129.520 134.205 129.690 134.905 ;
        RECT 129.860 134.545 130.030 135.325 ;
        RECT 130.350 135.275 130.720 135.775 ;
        RECT 130.900 135.325 131.305 135.495 ;
        RECT 131.475 135.325 132.260 135.495 ;
        RECT 130.900 135.095 131.070 135.325 ;
        RECT 130.240 134.795 131.070 135.095 ;
        RECT 131.455 134.825 131.920 135.155 ;
        RECT 130.240 134.765 130.440 134.795 ;
        RECT 130.560 134.545 130.730 134.615 ;
        RECT 129.860 134.375 130.730 134.545 ;
        RECT 130.220 134.285 130.730 134.375 ;
        RECT 128.770 133.820 129.075 133.950 ;
        RECT 129.520 133.840 130.050 134.205 ;
        RECT 128.390 133.225 128.655 133.685 ;
        RECT 128.825 133.395 129.075 133.820 ;
        RECT 130.220 133.670 130.390 134.285 ;
        RECT 129.285 133.500 130.390 133.670 ;
        RECT 130.560 133.225 130.730 134.025 ;
        RECT 130.900 133.725 131.070 134.795 ;
        RECT 131.240 133.895 131.430 134.615 ;
        RECT 131.600 133.865 131.920 134.825 ;
        RECT 132.090 134.865 132.260 135.325 ;
        RECT 132.535 135.245 132.745 135.775 ;
        RECT 133.005 135.035 133.335 135.560 ;
        RECT 133.505 135.165 133.675 135.775 ;
        RECT 133.845 135.120 134.175 135.555 ;
        RECT 133.845 135.035 134.225 135.120 ;
        RECT 133.135 134.865 133.335 135.035 ;
        RECT 134.000 134.995 134.225 135.035 ;
        RECT 132.090 134.535 132.965 134.865 ;
        RECT 133.135 134.535 133.885 134.865 ;
        RECT 130.900 133.395 131.150 133.725 ;
        RECT 132.090 133.695 132.260 134.535 ;
        RECT 133.135 134.330 133.325 134.535 ;
        RECT 134.055 134.415 134.225 134.995 ;
        RECT 134.395 135.025 135.605 135.775 ;
        RECT 135.865 135.225 136.035 135.605 ;
        RECT 136.250 135.395 136.580 135.775 ;
        RECT 135.865 135.055 136.580 135.225 ;
        RECT 134.395 134.485 134.915 135.025 ;
        RECT 134.010 134.365 134.225 134.415 ;
        RECT 132.430 133.955 133.325 134.330 ;
        RECT 133.835 134.285 134.225 134.365 ;
        RECT 135.085 134.315 135.605 134.855 ;
        RECT 135.775 134.505 136.130 134.875 ;
        RECT 136.410 134.865 136.580 135.055 ;
        RECT 136.750 135.030 137.005 135.605 ;
        RECT 136.410 134.535 136.665 134.865 ;
        RECT 136.410 134.325 136.580 134.535 ;
        RECT 131.375 133.525 132.260 133.695 ;
        RECT 132.440 133.225 132.755 133.725 ;
        RECT 132.985 133.395 133.325 133.955 ;
        RECT 133.495 133.225 133.665 134.235 ;
        RECT 133.835 133.440 134.165 134.285 ;
        RECT 134.395 133.225 135.605 134.315 ;
        RECT 135.865 134.155 136.580 134.325 ;
        RECT 136.835 134.300 137.005 135.030 ;
        RECT 137.180 134.935 137.440 135.775 ;
        RECT 137.615 135.025 138.825 135.775 ;
        RECT 135.865 133.395 136.035 134.155 ;
        RECT 136.250 133.225 136.580 133.985 ;
        RECT 136.750 133.395 137.005 134.300 ;
        RECT 137.180 133.225 137.440 134.375 ;
        RECT 137.615 134.315 138.135 134.855 ;
        RECT 138.305 134.485 138.825 135.025 ;
        RECT 137.615 133.225 138.825 134.315 ;
        RECT 13.330 133.055 138.910 133.225 ;
        RECT 13.415 131.965 14.625 133.055 ;
        RECT 14.795 131.965 17.385 133.055 ;
        RECT 18.105 132.385 18.275 132.885 ;
        RECT 18.445 132.555 18.775 133.055 ;
        RECT 18.105 132.215 18.770 132.385 ;
        RECT 13.415 131.255 13.935 131.795 ;
        RECT 14.105 131.425 14.625 131.965 ;
        RECT 14.795 131.275 16.005 131.795 ;
        RECT 16.175 131.445 17.385 131.965 ;
        RECT 18.020 131.395 18.370 132.045 ;
        RECT 13.415 130.505 14.625 131.255 ;
        RECT 14.795 130.505 17.385 131.275 ;
        RECT 18.540 131.225 18.770 132.215 ;
        RECT 18.105 131.055 18.770 131.225 ;
        RECT 18.105 130.765 18.275 131.055 ;
        RECT 18.445 130.505 18.775 130.885 ;
        RECT 18.945 130.765 19.130 132.885 ;
        RECT 19.370 132.595 19.635 133.055 ;
        RECT 19.805 132.460 20.055 132.885 ;
        RECT 20.265 132.610 21.370 132.780 ;
        RECT 19.750 132.330 20.055 132.460 ;
        RECT 19.300 131.135 19.580 132.085 ;
        RECT 19.750 131.225 19.920 132.330 ;
        RECT 20.090 131.545 20.330 132.140 ;
        RECT 20.500 132.075 21.030 132.440 ;
        RECT 20.500 131.375 20.670 132.075 ;
        RECT 21.200 131.995 21.370 132.610 ;
        RECT 21.540 132.255 21.710 133.055 ;
        RECT 21.880 132.555 22.130 132.885 ;
        RECT 22.355 132.585 23.240 132.755 ;
        RECT 21.200 131.905 21.710 131.995 ;
        RECT 19.750 131.095 19.975 131.225 ;
        RECT 20.145 131.155 20.670 131.375 ;
        RECT 20.840 131.735 21.710 131.905 ;
        RECT 19.385 130.505 19.635 130.965 ;
        RECT 19.805 130.955 19.975 131.095 ;
        RECT 20.840 130.955 21.010 131.735 ;
        RECT 21.540 131.665 21.710 131.735 ;
        RECT 21.220 131.485 21.420 131.515 ;
        RECT 21.880 131.485 22.050 132.555 ;
        RECT 22.220 131.665 22.410 132.385 ;
        RECT 21.220 131.185 22.050 131.485 ;
        RECT 22.580 131.455 22.900 132.415 ;
        RECT 19.805 130.785 20.140 130.955 ;
        RECT 20.335 130.785 21.010 130.955 ;
        RECT 21.330 130.505 21.700 131.005 ;
        RECT 21.880 130.955 22.050 131.185 ;
        RECT 22.435 131.125 22.900 131.455 ;
        RECT 23.070 131.745 23.240 132.585 ;
        RECT 23.420 132.555 23.735 133.055 ;
        RECT 23.965 132.325 24.305 132.885 ;
        RECT 23.410 131.950 24.305 132.325 ;
        RECT 24.475 132.045 24.645 133.055 ;
        RECT 24.115 131.745 24.305 131.950 ;
        RECT 24.815 131.995 25.145 132.840 ;
        RECT 24.815 131.915 25.205 131.995 ;
        RECT 24.990 131.865 25.205 131.915 ;
        RECT 26.295 131.890 26.585 133.055 ;
        RECT 26.755 132.500 27.360 133.055 ;
        RECT 27.535 132.545 28.015 132.885 ;
        RECT 28.185 132.510 28.440 133.055 ;
        RECT 26.755 132.400 27.370 132.500 ;
        RECT 27.185 132.375 27.370 132.400 ;
        RECT 23.070 131.415 23.945 131.745 ;
        RECT 24.115 131.415 24.865 131.745 ;
        RECT 23.070 130.955 23.240 131.415 ;
        RECT 24.115 131.245 24.315 131.415 ;
        RECT 25.035 131.285 25.205 131.865 ;
        RECT 26.755 131.780 27.015 132.230 ;
        RECT 27.185 132.130 27.515 132.375 ;
        RECT 27.685 132.055 28.440 132.305 ;
        RECT 28.610 132.185 28.885 132.885 ;
        RECT 27.670 132.020 28.440 132.055 ;
        RECT 27.655 132.010 28.440 132.020 ;
        RECT 27.650 131.995 28.545 132.010 ;
        RECT 27.630 131.980 28.545 131.995 ;
        RECT 27.610 131.970 28.545 131.980 ;
        RECT 27.585 131.960 28.545 131.970 ;
        RECT 27.515 131.930 28.545 131.960 ;
        RECT 27.495 131.900 28.545 131.930 ;
        RECT 27.475 131.870 28.545 131.900 ;
        RECT 27.445 131.845 28.545 131.870 ;
        RECT 27.410 131.810 28.545 131.845 ;
        RECT 27.380 131.805 28.545 131.810 ;
        RECT 27.380 131.800 27.770 131.805 ;
        RECT 27.380 131.790 27.745 131.800 ;
        RECT 27.380 131.785 27.730 131.790 ;
        RECT 27.380 131.780 27.715 131.785 ;
        RECT 26.755 131.775 27.715 131.780 ;
        RECT 26.755 131.765 27.705 131.775 ;
        RECT 26.755 131.760 27.695 131.765 ;
        RECT 26.755 131.750 27.685 131.760 ;
        RECT 26.755 131.740 27.680 131.750 ;
        RECT 26.755 131.735 27.675 131.740 ;
        RECT 26.755 131.720 27.665 131.735 ;
        RECT 26.755 131.705 27.660 131.720 ;
        RECT 26.755 131.680 27.650 131.705 ;
        RECT 26.755 131.610 27.645 131.680 ;
        RECT 24.980 131.245 25.205 131.285 ;
        RECT 21.880 130.785 22.285 130.955 ;
        RECT 22.455 130.785 23.240 130.955 ;
        RECT 23.515 130.505 23.725 131.035 ;
        RECT 23.985 130.720 24.315 131.245 ;
        RECT 24.825 131.160 25.205 131.245 ;
        RECT 24.485 130.505 24.655 131.115 ;
        RECT 24.825 130.725 25.155 131.160 ;
        RECT 26.295 130.505 26.585 131.230 ;
        RECT 26.755 131.055 27.305 131.440 ;
        RECT 27.475 130.885 27.645 131.610 ;
        RECT 26.755 130.715 27.645 130.885 ;
        RECT 27.815 131.210 28.145 131.635 ;
        RECT 28.315 131.410 28.545 131.805 ;
        RECT 27.815 130.725 28.035 131.210 ;
        RECT 28.715 131.155 28.885 132.185 ;
        RECT 29.065 132.085 29.395 132.870 ;
        RECT 29.065 131.915 29.745 132.085 ;
        RECT 29.925 131.915 30.255 133.055 ;
        RECT 31.355 132.205 31.735 132.885 ;
        RECT 32.325 132.205 32.495 133.055 ;
        RECT 32.665 132.375 32.995 132.885 ;
        RECT 33.165 132.545 33.335 133.055 ;
        RECT 33.505 132.375 33.905 132.885 ;
        RECT 32.665 132.205 33.905 132.375 ;
        RECT 29.055 131.495 29.405 131.745 ;
        RECT 29.575 131.315 29.745 131.915 ;
        RECT 29.915 131.495 30.265 131.745 ;
        RECT 28.205 130.505 28.455 131.045 ;
        RECT 28.625 130.675 28.885 131.155 ;
        RECT 29.075 130.505 29.315 131.315 ;
        RECT 29.485 130.675 29.815 131.315 ;
        RECT 29.985 130.505 30.255 131.315 ;
        RECT 31.355 131.245 31.525 132.205 ;
        RECT 31.695 131.865 33.000 132.035 ;
        RECT 34.085 131.955 34.405 132.885 ;
        RECT 34.665 132.385 34.835 132.885 ;
        RECT 35.005 132.555 35.335 133.055 ;
        RECT 34.665 132.215 35.330 132.385 ;
        RECT 31.695 131.415 31.940 131.865 ;
        RECT 32.110 131.495 32.660 131.695 ;
        RECT 32.830 131.665 33.000 131.865 ;
        RECT 33.775 131.785 34.405 131.955 ;
        RECT 32.830 131.495 33.205 131.665 ;
        RECT 33.375 131.245 33.605 131.745 ;
        RECT 31.355 131.075 33.605 131.245 ;
        RECT 31.405 130.505 31.735 130.895 ;
        RECT 31.905 130.755 32.075 131.075 ;
        RECT 33.775 130.905 33.945 131.785 ;
        RECT 34.580 131.395 34.930 132.045 ;
        RECT 32.245 130.505 32.575 130.895 ;
        RECT 32.990 130.735 33.945 130.905 ;
        RECT 34.115 130.505 34.405 131.340 ;
        RECT 35.100 131.225 35.330 132.215 ;
        RECT 34.665 131.055 35.330 131.225 ;
        RECT 34.665 130.765 34.835 131.055 ;
        RECT 35.005 130.505 35.335 130.885 ;
        RECT 35.505 130.765 35.690 132.885 ;
        RECT 35.930 132.595 36.195 133.055 ;
        RECT 36.365 132.460 36.615 132.885 ;
        RECT 36.825 132.610 37.930 132.780 ;
        RECT 36.310 132.330 36.615 132.460 ;
        RECT 35.860 131.135 36.140 132.085 ;
        RECT 36.310 131.225 36.480 132.330 ;
        RECT 36.650 131.545 36.890 132.140 ;
        RECT 37.060 132.075 37.590 132.440 ;
        RECT 37.060 131.375 37.230 132.075 ;
        RECT 37.760 131.995 37.930 132.610 ;
        RECT 38.100 132.255 38.270 133.055 ;
        RECT 38.440 132.555 38.690 132.885 ;
        RECT 38.915 132.585 39.800 132.755 ;
        RECT 37.760 131.905 38.270 131.995 ;
        RECT 36.310 131.095 36.535 131.225 ;
        RECT 36.705 131.155 37.230 131.375 ;
        RECT 37.400 131.735 38.270 131.905 ;
        RECT 35.945 130.505 36.195 130.965 ;
        RECT 36.365 130.955 36.535 131.095 ;
        RECT 37.400 130.955 37.570 131.735 ;
        RECT 38.100 131.665 38.270 131.735 ;
        RECT 37.780 131.485 37.980 131.515 ;
        RECT 38.440 131.485 38.610 132.555 ;
        RECT 38.780 131.665 38.970 132.385 ;
        RECT 37.780 131.185 38.610 131.485 ;
        RECT 39.140 131.455 39.460 132.415 ;
        RECT 36.365 130.785 36.700 130.955 ;
        RECT 36.895 130.785 37.570 130.955 ;
        RECT 37.890 130.505 38.260 131.005 ;
        RECT 38.440 130.955 38.610 131.185 ;
        RECT 38.995 131.125 39.460 131.455 ;
        RECT 39.630 131.745 39.800 132.585 ;
        RECT 39.980 132.555 40.295 133.055 ;
        RECT 40.525 132.325 40.865 132.885 ;
        RECT 39.970 131.950 40.865 132.325 ;
        RECT 41.035 132.045 41.205 133.055 ;
        RECT 40.675 131.745 40.865 131.950 ;
        RECT 41.375 131.995 41.705 132.840 ;
        RECT 41.945 132.445 42.275 132.875 ;
        RECT 42.455 132.615 42.650 133.055 ;
        RECT 42.820 132.445 43.150 132.875 ;
        RECT 41.945 132.275 43.150 132.445 ;
        RECT 41.375 131.915 41.765 131.995 ;
        RECT 41.945 131.945 42.840 132.275 ;
        RECT 43.320 132.105 43.595 132.875 ;
        RECT 43.775 132.500 44.380 133.055 ;
        RECT 44.555 132.545 45.035 132.885 ;
        RECT 45.205 132.510 45.460 133.055 ;
        RECT 43.775 132.400 44.390 132.500 ;
        RECT 44.205 132.375 44.390 132.400 ;
        RECT 41.550 131.865 41.765 131.915 ;
        RECT 39.630 131.415 40.505 131.745 ;
        RECT 40.675 131.415 41.425 131.745 ;
        RECT 39.630 130.955 39.800 131.415 ;
        RECT 40.675 131.245 40.875 131.415 ;
        RECT 41.595 131.285 41.765 131.865 ;
        RECT 43.010 131.915 43.595 132.105 ;
        RECT 41.950 131.415 42.245 131.745 ;
        RECT 42.425 131.415 42.840 131.745 ;
        RECT 41.540 131.245 41.765 131.285 ;
        RECT 38.440 130.785 38.845 130.955 ;
        RECT 39.015 130.785 39.800 130.955 ;
        RECT 40.075 130.505 40.285 131.035 ;
        RECT 40.545 130.720 40.875 131.245 ;
        RECT 41.385 131.160 41.765 131.245 ;
        RECT 41.045 130.505 41.215 131.115 ;
        RECT 41.385 130.725 41.715 131.160 ;
        RECT 41.945 130.505 42.245 131.235 ;
        RECT 42.425 130.795 42.655 131.415 ;
        RECT 43.010 131.245 43.185 131.915 ;
        RECT 43.775 131.780 44.035 132.230 ;
        RECT 44.205 132.130 44.535 132.375 ;
        RECT 44.705 132.055 45.460 132.305 ;
        RECT 45.630 132.185 45.905 132.885 ;
        RECT 46.075 132.500 46.680 133.055 ;
        RECT 46.855 132.545 47.335 132.885 ;
        RECT 47.505 132.510 47.760 133.055 ;
        RECT 46.075 132.400 46.690 132.500 ;
        RECT 46.505 132.375 46.690 132.400 ;
        RECT 44.690 132.020 45.460 132.055 ;
        RECT 44.675 132.010 45.460 132.020 ;
        RECT 44.670 131.995 45.565 132.010 ;
        RECT 44.650 131.980 45.565 131.995 ;
        RECT 44.630 131.970 45.565 131.980 ;
        RECT 44.605 131.960 45.565 131.970 ;
        RECT 44.535 131.930 45.565 131.960 ;
        RECT 44.515 131.900 45.565 131.930 ;
        RECT 44.495 131.870 45.565 131.900 ;
        RECT 44.465 131.845 45.565 131.870 ;
        RECT 44.430 131.810 45.565 131.845 ;
        RECT 44.400 131.805 45.565 131.810 ;
        RECT 44.400 131.800 44.790 131.805 ;
        RECT 44.400 131.790 44.765 131.800 ;
        RECT 44.400 131.785 44.750 131.790 ;
        RECT 44.400 131.780 44.735 131.785 ;
        RECT 43.775 131.775 44.735 131.780 ;
        RECT 43.775 131.765 44.725 131.775 ;
        RECT 43.775 131.760 44.715 131.765 ;
        RECT 43.775 131.750 44.705 131.760 ;
        RECT 42.855 131.065 43.185 131.245 ;
        RECT 43.355 131.095 43.595 131.745 ;
        RECT 43.775 131.740 44.700 131.750 ;
        RECT 43.775 131.735 44.695 131.740 ;
        RECT 43.775 131.720 44.685 131.735 ;
        RECT 43.775 131.705 44.680 131.720 ;
        RECT 43.775 131.680 44.670 131.705 ;
        RECT 43.775 131.610 44.665 131.680 ;
        RECT 42.855 130.685 43.080 131.065 ;
        RECT 43.775 131.055 44.325 131.440 ;
        RECT 43.250 130.505 43.580 130.895 ;
        RECT 44.495 130.885 44.665 131.610 ;
        RECT 43.775 130.715 44.665 130.885 ;
        RECT 44.835 131.210 45.165 131.635 ;
        RECT 45.335 131.410 45.565 131.805 ;
        RECT 44.835 130.725 45.055 131.210 ;
        RECT 45.735 131.155 45.905 132.185 ;
        RECT 46.075 131.780 46.335 132.230 ;
        RECT 46.505 132.130 46.835 132.375 ;
        RECT 47.005 132.055 47.760 132.305 ;
        RECT 47.930 132.185 48.205 132.885 ;
        RECT 46.990 132.020 47.760 132.055 ;
        RECT 46.975 132.010 47.760 132.020 ;
        RECT 46.970 131.995 47.865 132.010 ;
        RECT 46.950 131.980 47.865 131.995 ;
        RECT 46.930 131.970 47.865 131.980 ;
        RECT 46.905 131.960 47.865 131.970 ;
        RECT 46.835 131.930 47.865 131.960 ;
        RECT 46.815 131.900 47.865 131.930 ;
        RECT 46.795 131.870 47.865 131.900 ;
        RECT 46.765 131.845 47.865 131.870 ;
        RECT 46.730 131.810 47.865 131.845 ;
        RECT 46.700 131.805 47.865 131.810 ;
        RECT 46.700 131.800 47.090 131.805 ;
        RECT 46.700 131.790 47.065 131.800 ;
        RECT 46.700 131.785 47.050 131.790 ;
        RECT 46.700 131.780 47.035 131.785 ;
        RECT 46.075 131.775 47.035 131.780 ;
        RECT 46.075 131.765 47.025 131.775 ;
        RECT 46.075 131.760 47.015 131.765 ;
        RECT 46.075 131.750 47.005 131.760 ;
        RECT 46.075 131.740 47.000 131.750 ;
        RECT 46.075 131.735 46.995 131.740 ;
        RECT 46.075 131.720 46.985 131.735 ;
        RECT 46.075 131.705 46.980 131.720 ;
        RECT 46.075 131.680 46.970 131.705 ;
        RECT 46.075 131.610 46.965 131.680 ;
        RECT 45.225 130.505 45.475 131.045 ;
        RECT 45.645 130.675 45.905 131.155 ;
        RECT 46.075 131.055 46.625 131.440 ;
        RECT 46.795 130.885 46.965 131.610 ;
        RECT 46.075 130.715 46.965 130.885 ;
        RECT 47.135 131.210 47.465 131.635 ;
        RECT 47.635 131.410 47.865 131.805 ;
        RECT 47.135 130.725 47.355 131.210 ;
        RECT 48.035 131.155 48.205 132.185 ;
        RECT 48.385 132.085 48.715 132.870 ;
        RECT 48.385 131.915 49.065 132.085 ;
        RECT 49.245 131.915 49.575 133.055 ;
        RECT 49.755 132.500 50.360 133.055 ;
        RECT 50.535 132.545 51.015 132.885 ;
        RECT 51.185 132.510 51.440 133.055 ;
        RECT 49.755 132.400 50.370 132.500 ;
        RECT 50.185 132.375 50.370 132.400 ;
        RECT 48.375 131.495 48.725 131.745 ;
        RECT 48.895 131.315 49.065 131.915 ;
        RECT 49.755 131.780 50.015 132.230 ;
        RECT 50.185 132.130 50.515 132.375 ;
        RECT 50.685 132.055 51.440 132.305 ;
        RECT 51.610 132.185 51.885 132.885 ;
        RECT 50.670 132.020 51.440 132.055 ;
        RECT 50.655 132.010 51.440 132.020 ;
        RECT 50.650 131.995 51.545 132.010 ;
        RECT 50.630 131.980 51.545 131.995 ;
        RECT 50.610 131.970 51.545 131.980 ;
        RECT 50.585 131.960 51.545 131.970 ;
        RECT 50.515 131.930 51.545 131.960 ;
        RECT 50.495 131.900 51.545 131.930 ;
        RECT 50.475 131.870 51.545 131.900 ;
        RECT 50.445 131.845 51.545 131.870 ;
        RECT 50.410 131.810 51.545 131.845 ;
        RECT 50.380 131.805 51.545 131.810 ;
        RECT 50.380 131.800 50.770 131.805 ;
        RECT 50.380 131.790 50.745 131.800 ;
        RECT 50.380 131.785 50.730 131.790 ;
        RECT 50.380 131.780 50.715 131.785 ;
        RECT 49.755 131.775 50.715 131.780 ;
        RECT 49.755 131.765 50.705 131.775 ;
        RECT 49.755 131.760 50.695 131.765 ;
        RECT 49.755 131.750 50.685 131.760 ;
        RECT 49.235 131.495 49.585 131.745 ;
        RECT 49.755 131.740 50.680 131.750 ;
        RECT 49.755 131.735 50.675 131.740 ;
        RECT 49.755 131.720 50.665 131.735 ;
        RECT 49.755 131.705 50.660 131.720 ;
        RECT 49.755 131.680 50.650 131.705 ;
        RECT 49.755 131.610 50.645 131.680 ;
        RECT 47.525 130.505 47.775 131.045 ;
        RECT 47.945 130.675 48.205 131.155 ;
        RECT 48.395 130.505 48.635 131.315 ;
        RECT 48.805 130.675 49.135 131.315 ;
        RECT 49.305 130.505 49.575 131.315 ;
        RECT 49.755 131.055 50.305 131.440 ;
        RECT 50.475 130.885 50.645 131.610 ;
        RECT 49.755 130.715 50.645 130.885 ;
        RECT 50.815 131.210 51.145 131.635 ;
        RECT 51.315 131.410 51.545 131.805 ;
        RECT 50.815 131.185 51.065 131.210 ;
        RECT 50.815 130.725 51.035 131.185 ;
        RECT 51.715 131.155 51.885 132.185 ;
        RECT 52.055 131.890 52.345 133.055 ;
        RECT 52.515 132.620 57.860 133.055 ;
        RECT 58.035 132.620 63.380 133.055 ;
        RECT 51.205 130.505 51.455 131.045 ;
        RECT 51.625 130.675 51.885 131.155 ;
        RECT 52.055 130.505 52.345 131.230 ;
        RECT 54.100 131.050 54.440 131.880 ;
        RECT 55.920 131.370 56.270 132.620 ;
        RECT 59.620 131.050 59.960 131.880 ;
        RECT 61.440 131.370 61.790 132.620 ;
        RECT 63.555 131.965 67.065 133.055 ;
        RECT 63.555 131.275 65.205 131.795 ;
        RECT 65.375 131.445 67.065 131.965 ;
        RECT 67.730 132.265 68.265 132.885 ;
        RECT 52.515 130.505 57.860 131.050 ;
        RECT 58.035 130.505 63.380 131.050 ;
        RECT 63.555 130.505 67.065 131.275 ;
        RECT 67.730 131.245 68.045 132.265 ;
        RECT 68.435 132.255 68.765 133.055 ;
        RECT 69.250 132.085 69.640 132.260 ;
        RECT 68.215 131.915 69.640 132.085 ;
        RECT 70.180 132.085 70.570 132.260 ;
        RECT 71.055 132.255 71.385 133.055 ;
        RECT 71.555 132.265 72.090 132.885 ;
        RECT 70.180 131.915 71.605 132.085 ;
        RECT 68.215 131.415 68.385 131.915 ;
        RECT 67.730 130.675 68.345 131.245 ;
        RECT 68.635 131.185 68.900 131.745 ;
        RECT 69.070 131.015 69.240 131.915 ;
        RECT 69.410 131.185 69.765 131.745 ;
        RECT 70.055 131.185 70.410 131.745 ;
        RECT 70.580 131.015 70.750 131.915 ;
        RECT 70.920 131.185 71.185 131.745 ;
        RECT 71.435 131.415 71.605 131.915 ;
        RECT 71.775 131.245 72.090 132.265 ;
        RECT 68.515 130.505 68.730 131.015 ;
        RECT 68.960 130.685 69.240 131.015 ;
        RECT 69.420 130.505 69.660 131.015 ;
        RECT 70.160 130.505 70.400 131.015 ;
        RECT 70.580 130.685 70.860 131.015 ;
        RECT 71.090 130.505 71.305 131.015 ;
        RECT 71.475 130.675 72.090 131.245 ;
        RECT 72.295 132.335 72.755 132.885 ;
        RECT 72.945 132.335 73.275 133.055 ;
        RECT 72.295 130.965 72.545 132.335 ;
        RECT 73.475 132.165 73.775 132.715 ;
        RECT 73.945 132.385 74.225 133.055 ;
        RECT 72.835 131.995 73.775 132.165 ;
        RECT 72.835 131.745 73.005 131.995 ;
        RECT 74.145 131.745 74.410 132.105 ;
        RECT 74.595 131.965 77.185 133.055 ;
        RECT 72.715 131.415 73.005 131.745 ;
        RECT 73.175 131.495 73.515 131.745 ;
        RECT 73.735 131.495 74.410 131.745 ;
        RECT 72.835 131.325 73.005 131.415 ;
        RECT 72.835 131.135 74.225 131.325 ;
        RECT 72.295 130.675 72.855 130.965 ;
        RECT 73.025 130.505 73.275 130.965 ;
        RECT 73.895 130.775 74.225 131.135 ;
        RECT 74.595 131.275 75.805 131.795 ;
        RECT 75.975 131.445 77.185 131.965 ;
        RECT 77.815 131.890 78.105 133.055 ;
        RECT 78.735 131.915 78.995 133.055 ;
        RECT 79.235 132.545 80.850 132.875 ;
        RECT 79.245 131.745 79.415 132.305 ;
        RECT 79.675 132.205 80.850 132.375 ;
        RECT 81.020 132.255 81.300 133.055 ;
        RECT 79.675 131.915 80.005 132.205 ;
        RECT 80.680 132.085 80.850 132.205 ;
        RECT 80.175 131.745 80.420 132.035 ;
        RECT 80.680 131.915 81.340 132.085 ;
        RECT 81.510 131.915 81.785 132.885 ;
        RECT 81.955 132.500 82.560 133.055 ;
        RECT 82.735 132.545 83.215 132.885 ;
        RECT 83.385 132.510 83.640 133.055 ;
        RECT 81.955 132.400 82.570 132.500 ;
        RECT 82.385 132.375 82.570 132.400 ;
        RECT 81.170 131.745 81.340 131.915 ;
        RECT 78.740 131.495 79.075 131.745 ;
        RECT 79.245 131.415 79.960 131.745 ;
        RECT 80.175 131.415 81.000 131.745 ;
        RECT 81.170 131.415 81.445 131.745 ;
        RECT 79.245 131.325 79.495 131.415 ;
        RECT 74.595 130.505 77.185 131.275 ;
        RECT 77.815 130.505 78.105 131.230 ;
        RECT 78.735 130.505 78.995 131.325 ;
        RECT 79.165 130.905 79.495 131.325 ;
        RECT 81.170 131.245 81.340 131.415 ;
        RECT 79.675 131.075 81.340 131.245 ;
        RECT 81.615 131.180 81.785 131.915 ;
        RECT 81.955 131.780 82.215 132.230 ;
        RECT 82.385 132.130 82.715 132.375 ;
        RECT 82.885 132.055 83.640 132.305 ;
        RECT 83.810 132.185 84.085 132.885 ;
        RECT 84.345 132.385 84.515 132.885 ;
        RECT 84.685 132.555 85.015 133.055 ;
        RECT 84.345 132.215 85.010 132.385 ;
        RECT 82.870 132.020 83.640 132.055 ;
        RECT 82.855 132.010 83.640 132.020 ;
        RECT 82.850 131.995 83.745 132.010 ;
        RECT 82.830 131.980 83.745 131.995 ;
        RECT 82.810 131.970 83.745 131.980 ;
        RECT 82.785 131.960 83.745 131.970 ;
        RECT 82.715 131.930 83.745 131.960 ;
        RECT 82.695 131.900 83.745 131.930 ;
        RECT 82.675 131.870 83.745 131.900 ;
        RECT 82.645 131.845 83.745 131.870 ;
        RECT 82.610 131.810 83.745 131.845 ;
        RECT 82.580 131.805 83.745 131.810 ;
        RECT 82.580 131.800 82.970 131.805 ;
        RECT 82.580 131.790 82.945 131.800 ;
        RECT 82.580 131.785 82.930 131.790 ;
        RECT 82.580 131.780 82.915 131.785 ;
        RECT 81.955 131.775 82.915 131.780 ;
        RECT 81.955 131.765 82.905 131.775 ;
        RECT 81.955 131.760 82.895 131.765 ;
        RECT 81.955 131.750 82.885 131.760 ;
        RECT 81.955 131.740 82.880 131.750 ;
        RECT 81.955 131.735 82.875 131.740 ;
        RECT 81.955 131.720 82.865 131.735 ;
        RECT 81.955 131.705 82.860 131.720 ;
        RECT 81.955 131.680 82.850 131.705 ;
        RECT 81.955 131.610 82.845 131.680 ;
        RECT 79.675 130.675 79.935 131.075 ;
        RECT 80.105 130.505 80.435 130.905 ;
        RECT 80.605 130.725 80.775 131.075 ;
        RECT 80.945 130.505 81.320 130.905 ;
        RECT 81.510 130.835 81.785 131.180 ;
        RECT 81.955 131.055 82.505 131.440 ;
        RECT 82.675 130.885 82.845 131.610 ;
        RECT 81.955 130.715 82.845 130.885 ;
        RECT 83.015 131.210 83.345 131.635 ;
        RECT 83.515 131.410 83.745 131.805 ;
        RECT 83.015 130.725 83.235 131.210 ;
        RECT 83.915 131.155 84.085 132.185 ;
        RECT 84.260 131.395 84.610 132.045 ;
        RECT 84.780 131.225 85.010 132.215 ;
        RECT 83.405 130.505 83.655 131.045 ;
        RECT 83.825 130.675 84.085 131.155 ;
        RECT 84.345 131.055 85.010 131.225 ;
        RECT 84.345 130.765 84.515 131.055 ;
        RECT 84.685 130.505 85.015 130.885 ;
        RECT 85.185 130.765 85.370 132.885 ;
        RECT 85.610 132.595 85.875 133.055 ;
        RECT 86.045 132.460 86.295 132.885 ;
        RECT 86.505 132.610 87.610 132.780 ;
        RECT 85.990 132.330 86.295 132.460 ;
        RECT 85.540 131.135 85.820 132.085 ;
        RECT 85.990 131.225 86.160 132.330 ;
        RECT 86.330 131.545 86.570 132.140 ;
        RECT 86.740 132.075 87.270 132.440 ;
        RECT 86.740 131.375 86.910 132.075 ;
        RECT 87.440 131.995 87.610 132.610 ;
        RECT 87.780 132.255 87.950 133.055 ;
        RECT 88.120 132.555 88.370 132.885 ;
        RECT 88.595 132.585 89.480 132.755 ;
        RECT 87.440 131.905 87.950 131.995 ;
        RECT 85.990 131.095 86.215 131.225 ;
        RECT 86.385 131.155 86.910 131.375 ;
        RECT 87.080 131.735 87.950 131.905 ;
        RECT 85.625 130.505 85.875 130.965 ;
        RECT 86.045 130.955 86.215 131.095 ;
        RECT 87.080 130.955 87.250 131.735 ;
        RECT 87.780 131.665 87.950 131.735 ;
        RECT 87.460 131.485 87.660 131.515 ;
        RECT 88.120 131.485 88.290 132.555 ;
        RECT 88.460 131.665 88.650 132.385 ;
        RECT 87.460 131.185 88.290 131.485 ;
        RECT 88.820 131.455 89.140 132.415 ;
        RECT 86.045 130.785 86.380 130.955 ;
        RECT 86.575 130.785 87.250 130.955 ;
        RECT 87.570 130.505 87.940 131.005 ;
        RECT 88.120 130.955 88.290 131.185 ;
        RECT 88.675 131.125 89.140 131.455 ;
        RECT 89.310 131.745 89.480 132.585 ;
        RECT 89.660 132.555 89.975 133.055 ;
        RECT 90.205 132.325 90.545 132.885 ;
        RECT 89.650 131.950 90.545 132.325 ;
        RECT 90.715 132.045 90.885 133.055 ;
        RECT 90.355 131.745 90.545 131.950 ;
        RECT 91.055 131.995 91.385 132.840 ;
        RECT 91.555 132.140 91.725 133.055 ;
        RECT 91.055 131.915 91.445 131.995 ;
        RECT 92.075 131.965 93.745 133.055 ;
        RECT 94.465 132.385 94.635 132.885 ;
        RECT 94.805 132.555 95.135 133.055 ;
        RECT 94.465 132.215 95.130 132.385 ;
        RECT 91.230 131.865 91.445 131.915 ;
        RECT 89.310 131.415 90.185 131.745 ;
        RECT 90.355 131.415 91.105 131.745 ;
        RECT 89.310 130.955 89.480 131.415 ;
        RECT 90.355 131.245 90.555 131.415 ;
        RECT 91.275 131.285 91.445 131.865 ;
        RECT 91.220 131.245 91.445 131.285 ;
        RECT 88.120 130.785 88.525 130.955 ;
        RECT 88.695 130.785 89.480 130.955 ;
        RECT 89.755 130.505 89.965 131.035 ;
        RECT 90.225 130.720 90.555 131.245 ;
        RECT 91.065 131.160 91.445 131.245 ;
        RECT 92.075 131.275 92.825 131.795 ;
        RECT 92.995 131.445 93.745 131.965 ;
        RECT 94.380 131.395 94.730 132.045 ;
        RECT 90.725 130.505 90.895 131.115 ;
        RECT 91.065 130.725 91.395 131.160 ;
        RECT 91.565 130.505 91.735 131.020 ;
        RECT 92.075 130.505 93.745 131.275 ;
        RECT 94.900 131.225 95.130 132.215 ;
        RECT 94.465 131.055 95.130 131.225 ;
        RECT 94.465 130.765 94.635 131.055 ;
        RECT 94.805 130.505 95.135 130.885 ;
        RECT 95.305 130.765 95.490 132.885 ;
        RECT 95.730 132.595 95.995 133.055 ;
        RECT 96.165 132.460 96.415 132.885 ;
        RECT 96.625 132.610 97.730 132.780 ;
        RECT 96.110 132.330 96.415 132.460 ;
        RECT 95.660 131.135 95.940 132.085 ;
        RECT 96.110 131.225 96.280 132.330 ;
        RECT 96.450 131.545 96.690 132.140 ;
        RECT 96.860 132.075 97.390 132.440 ;
        RECT 96.860 131.375 97.030 132.075 ;
        RECT 97.560 131.995 97.730 132.610 ;
        RECT 97.900 132.255 98.070 133.055 ;
        RECT 98.240 132.555 98.490 132.885 ;
        RECT 98.715 132.585 99.600 132.755 ;
        RECT 97.560 131.905 98.070 131.995 ;
        RECT 96.110 131.095 96.335 131.225 ;
        RECT 96.505 131.155 97.030 131.375 ;
        RECT 97.200 131.735 98.070 131.905 ;
        RECT 95.745 130.505 95.995 130.965 ;
        RECT 96.165 130.955 96.335 131.095 ;
        RECT 97.200 130.955 97.370 131.735 ;
        RECT 97.900 131.665 98.070 131.735 ;
        RECT 97.580 131.485 97.780 131.515 ;
        RECT 98.240 131.485 98.410 132.555 ;
        RECT 98.580 131.665 98.770 132.385 ;
        RECT 97.580 131.185 98.410 131.485 ;
        RECT 98.940 131.455 99.260 132.415 ;
        RECT 96.165 130.785 96.500 130.955 ;
        RECT 96.695 130.785 97.370 130.955 ;
        RECT 97.690 130.505 98.060 131.005 ;
        RECT 98.240 130.955 98.410 131.185 ;
        RECT 98.795 131.125 99.260 131.455 ;
        RECT 99.430 131.745 99.600 132.585 ;
        RECT 99.780 132.555 100.095 133.055 ;
        RECT 100.325 132.325 100.665 132.885 ;
        RECT 99.770 131.950 100.665 132.325 ;
        RECT 100.835 132.045 101.005 133.055 ;
        RECT 100.475 131.745 100.665 131.950 ;
        RECT 101.175 131.995 101.505 132.840 ;
        RECT 101.175 131.915 101.565 131.995 ;
        RECT 101.735 131.965 103.405 133.055 ;
        RECT 101.350 131.865 101.565 131.915 ;
        RECT 99.430 131.415 100.305 131.745 ;
        RECT 100.475 131.415 101.225 131.745 ;
        RECT 99.430 130.955 99.600 131.415 ;
        RECT 100.475 131.245 100.675 131.415 ;
        RECT 101.395 131.285 101.565 131.865 ;
        RECT 101.340 131.245 101.565 131.285 ;
        RECT 98.240 130.785 98.645 130.955 ;
        RECT 98.815 130.785 99.600 130.955 ;
        RECT 99.875 130.505 100.085 131.035 ;
        RECT 100.345 130.720 100.675 131.245 ;
        RECT 101.185 131.160 101.565 131.245 ;
        RECT 101.735 131.275 102.485 131.795 ;
        RECT 102.655 131.445 103.405 131.965 ;
        RECT 103.575 131.890 103.865 133.055 ;
        RECT 104.035 131.915 104.420 132.885 ;
        RECT 104.590 132.595 104.915 133.055 ;
        RECT 105.435 132.425 105.715 132.885 ;
        RECT 104.590 132.205 105.715 132.425 ;
        RECT 100.845 130.505 101.015 131.115 ;
        RECT 101.185 130.725 101.515 131.160 ;
        RECT 101.735 130.505 103.405 131.275 ;
        RECT 104.035 131.245 104.315 131.915 ;
        RECT 104.590 131.745 105.040 132.205 ;
        RECT 105.905 132.035 106.305 132.885 ;
        RECT 106.705 132.595 106.975 133.055 ;
        RECT 107.145 132.425 107.430 132.885 ;
        RECT 104.485 131.415 105.040 131.745 ;
        RECT 105.210 131.475 106.305 132.035 ;
        RECT 104.590 131.305 105.040 131.415 ;
        RECT 103.575 130.505 103.865 131.230 ;
        RECT 104.035 130.675 104.420 131.245 ;
        RECT 104.590 131.135 105.715 131.305 ;
        RECT 104.590 130.505 104.915 130.965 ;
        RECT 105.435 130.675 105.715 131.135 ;
        RECT 105.905 130.675 106.305 131.475 ;
        RECT 106.475 132.205 107.430 132.425 ;
        RECT 106.475 131.305 106.685 132.205 ;
        RECT 106.855 131.475 107.545 132.035 ;
        RECT 107.715 131.915 108.055 132.885 ;
        RECT 108.225 131.915 108.395 133.055 ;
        RECT 108.665 132.255 108.915 133.055 ;
        RECT 109.560 132.085 109.890 132.885 ;
        RECT 110.190 132.255 110.520 133.055 ;
        RECT 110.690 132.085 111.020 132.885 ;
        RECT 108.585 131.915 111.020 132.085 ;
        RECT 111.400 132.105 111.665 132.875 ;
        RECT 111.835 132.335 112.165 133.055 ;
        RECT 112.355 132.515 112.615 132.875 ;
        RECT 112.785 132.685 113.115 133.055 ;
        RECT 113.285 132.515 113.545 132.875 ;
        RECT 112.355 132.285 113.545 132.515 ;
        RECT 114.115 132.105 114.405 132.875 ;
        RECT 107.715 131.305 107.890 131.915 ;
        RECT 108.585 131.665 108.755 131.915 ;
        RECT 108.060 131.495 108.755 131.665 ;
        RECT 108.930 131.495 109.350 131.695 ;
        RECT 109.520 131.495 109.850 131.695 ;
        RECT 110.020 131.495 110.350 131.695 ;
        RECT 106.475 131.135 107.430 131.305 ;
        RECT 106.705 130.505 106.975 130.965 ;
        RECT 107.145 130.675 107.430 131.135 ;
        RECT 107.715 130.675 108.055 131.305 ;
        RECT 108.225 130.505 108.475 131.305 ;
        RECT 108.665 131.155 109.890 131.325 ;
        RECT 108.665 130.675 108.995 131.155 ;
        RECT 109.165 130.505 109.390 130.965 ;
        RECT 109.560 130.675 109.890 131.155 ;
        RECT 110.520 131.285 110.690 131.915 ;
        RECT 110.875 131.495 111.225 131.745 ;
        RECT 110.520 130.675 111.020 131.285 ;
        RECT 111.400 130.685 111.735 132.105 ;
        RECT 111.910 131.925 114.405 132.105 ;
        RECT 114.615 131.965 116.285 133.055 ;
        RECT 111.910 131.235 112.135 131.925 ;
        RECT 112.335 131.415 112.615 131.745 ;
        RECT 112.795 131.415 113.370 131.745 ;
        RECT 113.550 131.415 113.985 131.745 ;
        RECT 114.165 131.415 114.435 131.745 ;
        RECT 114.615 131.275 115.365 131.795 ;
        RECT 115.535 131.445 116.285 131.965 ;
        RECT 116.455 131.915 116.795 132.885 ;
        RECT 116.965 131.915 117.135 133.055 ;
        RECT 117.405 132.255 117.655 133.055 ;
        RECT 118.300 132.085 118.630 132.885 ;
        RECT 118.930 132.255 119.260 133.055 ;
        RECT 119.430 132.085 119.760 132.885 ;
        RECT 117.325 131.915 119.760 132.085 ;
        RECT 120.170 132.265 120.705 132.885 ;
        RECT 116.455 131.305 116.630 131.915 ;
        RECT 117.325 131.665 117.495 131.915 ;
        RECT 116.800 131.495 117.495 131.665 ;
        RECT 117.670 131.495 118.090 131.695 ;
        RECT 118.260 131.495 118.590 131.695 ;
        RECT 118.760 131.495 119.090 131.695 ;
        RECT 111.910 131.045 114.395 131.235 ;
        RECT 111.915 130.505 112.660 130.875 ;
        RECT 113.225 130.685 113.480 131.045 ;
        RECT 113.660 130.505 113.990 130.875 ;
        RECT 114.170 130.685 114.395 131.045 ;
        RECT 114.615 130.505 116.285 131.275 ;
        RECT 116.455 130.675 116.795 131.305 ;
        RECT 116.965 130.505 117.215 131.305 ;
        RECT 117.405 131.155 118.630 131.325 ;
        RECT 117.405 130.675 117.735 131.155 ;
        RECT 117.905 130.505 118.130 130.965 ;
        RECT 118.300 130.675 118.630 131.155 ;
        RECT 119.260 131.285 119.430 131.915 ;
        RECT 119.615 131.495 119.965 131.745 ;
        RECT 119.260 130.675 119.760 131.285 ;
        RECT 120.170 131.245 120.485 132.265 ;
        RECT 120.875 132.255 121.205 133.055 ;
        RECT 121.690 132.085 122.080 132.260 ;
        RECT 120.655 131.915 122.080 132.085 ;
        RECT 122.435 131.965 125.025 133.055 ;
        RECT 120.655 131.415 120.825 131.915 ;
        RECT 120.170 130.675 120.785 131.245 ;
        RECT 121.075 131.185 121.340 131.745 ;
        RECT 121.510 131.015 121.680 131.915 ;
        RECT 121.850 131.185 122.205 131.745 ;
        RECT 122.435 131.275 123.645 131.795 ;
        RECT 123.815 131.445 125.025 131.965 ;
        RECT 125.860 132.085 126.190 132.885 ;
        RECT 126.360 132.255 126.690 133.055 ;
        RECT 126.990 132.085 127.320 132.885 ;
        RECT 127.965 132.255 128.215 133.055 ;
        RECT 125.860 131.915 128.295 132.085 ;
        RECT 128.485 131.915 128.655 133.055 ;
        RECT 128.825 131.915 129.165 132.885 ;
        RECT 125.655 131.495 126.005 131.745 ;
        RECT 126.190 131.285 126.360 131.915 ;
        RECT 126.530 131.495 126.860 131.695 ;
        RECT 127.030 131.495 127.360 131.695 ;
        RECT 127.530 131.495 127.950 131.695 ;
        RECT 128.125 131.665 128.295 131.915 ;
        RECT 128.935 131.865 129.165 131.915 ;
        RECT 129.335 131.890 129.625 133.055 ;
        RECT 129.830 132.265 130.365 132.885 ;
        RECT 128.125 131.495 128.820 131.665 ;
        RECT 120.955 130.505 121.170 131.015 ;
        RECT 121.400 130.685 121.680 131.015 ;
        RECT 121.860 130.505 122.100 131.015 ;
        RECT 122.435 130.505 125.025 131.275 ;
        RECT 125.860 130.675 126.360 131.285 ;
        RECT 126.990 131.155 128.215 131.325 ;
        RECT 128.990 131.305 129.165 131.865 ;
        RECT 126.990 130.675 127.320 131.155 ;
        RECT 127.490 130.505 127.715 130.965 ;
        RECT 127.885 130.675 128.215 131.155 ;
        RECT 128.405 130.505 128.655 131.305 ;
        RECT 128.825 130.675 129.165 131.305 ;
        RECT 129.830 131.245 130.145 132.265 ;
        RECT 130.535 132.255 130.865 133.055 ;
        RECT 132.130 132.265 132.665 132.885 ;
        RECT 131.350 132.085 131.740 132.260 ;
        RECT 130.315 131.915 131.740 132.085 ;
        RECT 130.315 131.415 130.485 131.915 ;
        RECT 129.335 130.505 129.625 131.230 ;
        RECT 129.830 130.675 130.445 131.245 ;
        RECT 130.735 131.185 131.000 131.745 ;
        RECT 131.170 131.015 131.340 131.915 ;
        RECT 131.510 131.185 131.865 131.745 ;
        RECT 132.130 131.245 132.445 132.265 ;
        RECT 132.835 132.255 133.165 133.055 ;
        RECT 133.650 132.085 134.040 132.260 ;
        RECT 132.615 131.915 134.040 132.085 ;
        RECT 134.395 131.965 135.605 133.055 ;
        RECT 132.615 131.415 132.785 131.915 ;
        RECT 130.615 130.505 130.830 131.015 ;
        RECT 131.060 130.685 131.340 131.015 ;
        RECT 131.520 130.505 131.760 131.015 ;
        RECT 132.130 130.675 132.745 131.245 ;
        RECT 133.035 131.185 133.300 131.745 ;
        RECT 133.470 131.015 133.640 131.915 ;
        RECT 133.810 131.185 134.165 131.745 ;
        RECT 134.395 131.255 134.915 131.795 ;
        RECT 135.085 131.425 135.605 131.965 ;
        RECT 135.865 132.125 136.035 132.885 ;
        RECT 136.250 132.295 136.580 133.055 ;
        RECT 135.865 131.955 136.580 132.125 ;
        RECT 136.750 131.980 137.005 132.885 ;
        RECT 135.775 131.405 136.130 131.775 ;
        RECT 136.410 131.745 136.580 131.955 ;
        RECT 136.410 131.415 136.665 131.745 ;
        RECT 132.915 130.505 133.130 131.015 ;
        RECT 133.360 130.685 133.640 131.015 ;
        RECT 133.820 130.505 134.060 131.015 ;
        RECT 134.395 130.505 135.605 131.255 ;
        RECT 136.410 131.225 136.580 131.415 ;
        RECT 136.835 131.250 137.005 131.980 ;
        RECT 137.180 131.905 137.440 133.055 ;
        RECT 137.615 131.965 138.825 133.055 ;
        RECT 137.615 131.425 138.135 131.965 ;
        RECT 135.865 131.055 136.580 131.225 ;
        RECT 135.865 130.675 136.035 131.055 ;
        RECT 136.250 130.505 136.580 130.885 ;
        RECT 136.750 130.675 137.005 131.250 ;
        RECT 137.180 130.505 137.440 131.345 ;
        RECT 138.305 131.255 138.825 131.795 ;
        RECT 137.615 130.505 138.825 131.255 ;
        RECT 13.330 130.335 138.910 130.505 ;
        RECT 13.415 129.585 14.625 130.335 ;
        RECT 14.795 129.790 20.140 130.335 ;
        RECT 13.415 129.045 13.935 129.585 ;
        RECT 14.105 128.875 14.625 129.415 ;
        RECT 16.380 128.960 16.720 129.790 ;
        RECT 20.315 129.565 21.985 130.335 ;
        RECT 22.205 129.680 22.535 130.115 ;
        RECT 22.705 129.725 22.875 130.335 ;
        RECT 22.155 129.595 22.535 129.680 ;
        RECT 23.045 129.595 23.375 130.120 ;
        RECT 23.635 129.805 23.845 130.335 ;
        RECT 24.120 129.885 24.905 130.055 ;
        RECT 25.075 129.885 25.480 130.055 ;
        RECT 13.415 127.785 14.625 128.875 ;
        RECT 18.200 128.220 18.550 129.470 ;
        RECT 20.315 129.045 21.065 129.565 ;
        RECT 22.155 129.555 22.380 129.595 ;
        RECT 21.235 128.875 21.985 129.395 ;
        RECT 14.795 127.785 20.140 128.220 ;
        RECT 20.315 127.785 21.985 128.875 ;
        RECT 22.155 128.975 22.325 129.555 ;
        RECT 23.045 129.425 23.245 129.595 ;
        RECT 24.120 129.425 24.290 129.885 ;
        RECT 22.495 129.095 23.245 129.425 ;
        RECT 23.415 129.095 24.290 129.425 ;
        RECT 22.155 128.925 22.370 128.975 ;
        RECT 22.155 128.845 22.545 128.925 ;
        RECT 22.215 128.000 22.545 128.845 ;
        RECT 23.055 128.890 23.245 129.095 ;
        RECT 22.715 127.785 22.885 128.795 ;
        RECT 23.055 128.515 23.950 128.890 ;
        RECT 23.055 127.955 23.395 128.515 ;
        RECT 23.625 127.785 23.940 128.285 ;
        RECT 24.120 128.255 24.290 129.095 ;
        RECT 24.460 129.385 24.925 129.715 ;
        RECT 25.310 129.655 25.480 129.885 ;
        RECT 25.660 129.835 26.030 130.335 ;
        RECT 26.350 129.885 27.025 130.055 ;
        RECT 27.220 129.885 27.555 130.055 ;
        RECT 24.460 128.425 24.780 129.385 ;
        RECT 25.310 129.355 26.140 129.655 ;
        RECT 24.950 128.455 25.140 129.175 ;
        RECT 25.310 128.285 25.480 129.355 ;
        RECT 25.940 129.325 26.140 129.355 ;
        RECT 25.650 129.105 25.820 129.175 ;
        RECT 26.350 129.105 26.520 129.885 ;
        RECT 27.385 129.745 27.555 129.885 ;
        RECT 27.725 129.875 27.975 130.335 ;
        RECT 25.650 128.935 26.520 129.105 ;
        RECT 26.690 129.465 27.215 129.685 ;
        RECT 27.385 129.615 27.610 129.745 ;
        RECT 25.650 128.845 26.160 128.935 ;
        RECT 24.120 128.085 25.005 128.255 ;
        RECT 25.230 127.955 25.480 128.285 ;
        RECT 25.650 127.785 25.820 128.585 ;
        RECT 25.990 128.230 26.160 128.845 ;
        RECT 26.690 128.765 26.860 129.465 ;
        RECT 26.330 128.400 26.860 128.765 ;
        RECT 27.030 128.700 27.270 129.295 ;
        RECT 27.440 128.510 27.610 129.615 ;
        RECT 27.780 128.755 28.060 129.705 ;
        RECT 27.305 128.380 27.610 128.510 ;
        RECT 25.990 128.060 27.095 128.230 ;
        RECT 27.305 127.955 27.555 128.380 ;
        RECT 27.725 127.785 27.990 128.245 ;
        RECT 28.230 127.955 28.415 130.075 ;
        RECT 28.585 129.955 28.915 130.335 ;
        RECT 29.085 129.785 29.255 130.075 ;
        RECT 29.515 129.790 34.860 130.335 ;
        RECT 28.590 129.615 29.255 129.785 ;
        RECT 28.590 128.625 28.820 129.615 ;
        RECT 28.990 128.795 29.340 129.445 ;
        RECT 31.100 128.960 31.440 129.790 ;
        RECT 35.035 129.685 35.295 130.165 ;
        RECT 35.465 129.795 35.715 130.335 ;
        RECT 28.590 128.455 29.255 128.625 ;
        RECT 28.585 127.785 28.915 128.285 ;
        RECT 29.085 127.955 29.255 128.455 ;
        RECT 32.920 128.220 33.270 129.470 ;
        RECT 35.035 128.655 35.205 129.685 ;
        RECT 35.885 129.655 36.105 130.115 ;
        RECT 35.855 129.630 36.105 129.655 ;
        RECT 35.375 129.035 35.605 129.430 ;
        RECT 35.775 129.205 36.105 129.630 ;
        RECT 36.275 129.955 37.165 130.125 ;
        RECT 36.275 129.230 36.445 129.955 ;
        RECT 36.615 129.400 37.165 129.785 ;
        RECT 37.335 129.565 39.005 130.335 ;
        RECT 39.175 129.610 39.465 130.335 ;
        RECT 39.635 129.585 40.845 130.335 ;
        RECT 41.015 129.595 41.480 130.140 ;
        RECT 36.275 129.160 37.165 129.230 ;
        RECT 36.270 129.135 37.165 129.160 ;
        RECT 36.260 129.120 37.165 129.135 ;
        RECT 36.255 129.105 37.165 129.120 ;
        RECT 36.245 129.100 37.165 129.105 ;
        RECT 36.240 129.090 37.165 129.100 ;
        RECT 36.235 129.080 37.165 129.090 ;
        RECT 36.225 129.075 37.165 129.080 ;
        RECT 36.215 129.065 37.165 129.075 ;
        RECT 36.205 129.060 37.165 129.065 ;
        RECT 36.205 129.055 36.540 129.060 ;
        RECT 36.190 129.050 36.540 129.055 ;
        RECT 36.175 129.040 36.540 129.050 ;
        RECT 36.150 129.035 36.540 129.040 ;
        RECT 35.375 129.030 36.540 129.035 ;
        RECT 35.375 128.995 36.510 129.030 ;
        RECT 35.375 128.970 36.475 128.995 ;
        RECT 35.375 128.940 36.445 128.970 ;
        RECT 35.375 128.910 36.425 128.940 ;
        RECT 35.375 128.880 36.405 128.910 ;
        RECT 35.375 128.870 36.335 128.880 ;
        RECT 35.375 128.860 36.310 128.870 ;
        RECT 35.375 128.845 36.290 128.860 ;
        RECT 35.375 128.830 36.270 128.845 ;
        RECT 35.480 128.820 36.265 128.830 ;
        RECT 35.480 128.785 36.250 128.820 ;
        RECT 29.515 127.785 34.860 128.220 ;
        RECT 35.035 127.955 35.310 128.655 ;
        RECT 35.480 128.535 36.235 128.785 ;
        RECT 36.405 128.465 36.735 128.710 ;
        RECT 36.905 128.610 37.165 129.060 ;
        RECT 37.335 129.045 38.085 129.565 ;
        RECT 38.255 128.875 39.005 129.395 ;
        RECT 39.635 129.045 40.155 129.585 ;
        RECT 36.550 128.440 36.735 128.465 ;
        RECT 36.550 128.340 37.165 128.440 ;
        RECT 35.480 127.785 35.735 128.330 ;
        RECT 35.905 127.955 36.385 128.295 ;
        RECT 36.560 127.785 37.165 128.340 ;
        RECT 37.335 127.785 39.005 128.875 ;
        RECT 39.175 127.785 39.465 128.950 ;
        RECT 40.325 128.875 40.845 129.415 ;
        RECT 39.635 127.785 40.845 128.875 ;
        RECT 41.015 128.635 41.185 129.595 ;
        RECT 41.985 129.515 42.155 130.335 ;
        RECT 42.325 129.685 42.655 130.165 ;
        RECT 42.825 129.945 43.175 130.335 ;
        RECT 43.345 129.765 43.575 130.165 ;
        RECT 43.065 129.685 43.575 129.765 ;
        RECT 42.325 129.595 43.575 129.685 ;
        RECT 43.745 129.595 44.065 130.075 ;
        RECT 42.325 129.515 43.235 129.595 ;
        RECT 41.355 128.975 41.600 129.425 ;
        RECT 41.860 129.145 42.555 129.345 ;
        RECT 42.725 129.175 43.325 129.345 ;
        RECT 42.725 128.975 42.895 129.175 ;
        RECT 43.555 129.005 43.725 129.425 ;
        RECT 41.355 128.805 42.895 128.975 ;
        RECT 43.065 128.835 43.725 129.005 ;
        RECT 43.065 128.635 43.235 128.835 ;
        RECT 43.895 128.665 44.065 129.595 ;
        RECT 44.235 129.585 45.445 130.335 ;
        RECT 45.665 129.680 45.995 130.115 ;
        RECT 46.165 129.725 46.335 130.335 ;
        RECT 45.615 129.595 45.995 129.680 ;
        RECT 46.505 129.595 46.835 130.120 ;
        RECT 47.095 129.805 47.305 130.335 ;
        RECT 47.580 129.885 48.365 130.055 ;
        RECT 48.535 129.885 48.940 130.055 ;
        RECT 44.235 129.045 44.755 129.585 ;
        RECT 45.615 129.555 45.840 129.595 ;
        RECT 44.925 128.875 45.445 129.415 ;
        RECT 41.015 128.465 43.235 128.635 ;
        RECT 43.405 128.465 44.065 128.665 ;
        RECT 41.015 127.785 41.315 128.295 ;
        RECT 41.485 127.955 41.815 128.465 ;
        RECT 43.405 128.295 43.575 128.465 ;
        RECT 41.985 127.785 42.615 128.295 ;
        RECT 43.195 128.125 43.575 128.295 ;
        RECT 43.745 127.785 44.045 128.295 ;
        RECT 44.235 127.785 45.445 128.875 ;
        RECT 45.615 128.975 45.785 129.555 ;
        RECT 46.505 129.425 46.705 129.595 ;
        RECT 47.580 129.425 47.750 129.885 ;
        RECT 45.955 129.095 46.705 129.425 ;
        RECT 46.875 129.095 47.750 129.425 ;
        RECT 45.615 128.925 45.830 128.975 ;
        RECT 45.615 128.845 46.005 128.925 ;
        RECT 45.675 128.000 46.005 128.845 ;
        RECT 46.515 128.890 46.705 129.095 ;
        RECT 46.175 127.785 46.345 128.795 ;
        RECT 46.515 128.515 47.410 128.890 ;
        RECT 46.515 127.955 46.855 128.515 ;
        RECT 47.085 127.785 47.400 128.285 ;
        RECT 47.580 128.255 47.750 129.095 ;
        RECT 47.920 129.385 48.385 129.715 ;
        RECT 48.770 129.655 48.940 129.885 ;
        RECT 49.120 129.835 49.490 130.335 ;
        RECT 49.810 129.885 50.485 130.055 ;
        RECT 50.680 129.885 51.015 130.055 ;
        RECT 47.920 128.425 48.240 129.385 ;
        RECT 48.770 129.355 49.600 129.655 ;
        RECT 48.410 128.455 48.600 129.175 ;
        RECT 48.770 128.285 48.940 129.355 ;
        RECT 49.400 129.325 49.600 129.355 ;
        RECT 49.110 129.105 49.280 129.175 ;
        RECT 49.810 129.105 49.980 129.885 ;
        RECT 50.845 129.745 51.015 129.885 ;
        RECT 51.185 129.875 51.435 130.335 ;
        RECT 49.110 128.935 49.980 129.105 ;
        RECT 50.150 129.465 50.675 129.685 ;
        RECT 50.845 129.615 51.070 129.745 ;
        RECT 49.110 128.845 49.620 128.935 ;
        RECT 47.580 128.085 48.465 128.255 ;
        RECT 48.690 127.955 48.940 128.285 ;
        RECT 49.110 127.785 49.280 128.585 ;
        RECT 49.450 128.230 49.620 128.845 ;
        RECT 50.150 128.765 50.320 129.465 ;
        RECT 49.790 128.400 50.320 128.765 ;
        RECT 50.490 128.700 50.730 129.295 ;
        RECT 50.900 128.510 51.070 129.615 ;
        RECT 51.240 128.755 51.520 129.705 ;
        RECT 50.765 128.380 51.070 128.510 ;
        RECT 49.450 128.060 50.555 128.230 ;
        RECT 50.765 127.955 51.015 128.380 ;
        RECT 51.185 127.785 51.450 128.245 ;
        RECT 51.690 127.955 51.875 130.075 ;
        RECT 52.045 129.955 52.375 130.335 ;
        RECT 52.545 129.785 52.715 130.075 ;
        RECT 52.975 129.790 58.320 130.335 ;
        RECT 59.015 129.875 59.260 130.335 ;
        RECT 52.050 129.615 52.715 129.785 ;
        RECT 52.050 128.625 52.280 129.615 ;
        RECT 52.450 128.795 52.800 129.445 ;
        RECT 54.560 128.960 54.900 129.790 ;
        RECT 52.050 128.455 52.715 128.625 ;
        RECT 52.045 127.785 52.375 128.285 ;
        RECT 52.545 127.955 52.715 128.455 ;
        RECT 56.380 128.220 56.730 129.470 ;
        RECT 58.955 129.095 59.270 129.705 ;
        RECT 59.440 129.345 59.690 130.155 ;
        RECT 59.860 129.810 60.120 130.335 ;
        RECT 60.290 129.685 60.550 130.140 ;
        RECT 60.720 129.855 60.980 130.335 ;
        RECT 61.150 129.685 61.410 130.140 ;
        RECT 61.580 129.855 61.840 130.335 ;
        RECT 62.010 129.685 62.270 130.140 ;
        RECT 62.440 129.855 62.700 130.335 ;
        RECT 62.870 129.685 63.130 130.140 ;
        RECT 63.300 129.855 63.600 130.335 ;
        RECT 60.290 129.515 63.600 129.685 ;
        RECT 64.935 129.610 65.225 130.335 ;
        RECT 65.405 129.525 65.675 130.335 ;
        RECT 65.845 129.525 66.175 130.165 ;
        RECT 66.345 129.525 66.585 130.335 ;
        RECT 66.775 129.585 67.985 130.335 ;
        RECT 59.440 129.095 62.460 129.345 ;
        RECT 52.975 127.785 58.320 128.220 ;
        RECT 58.965 127.785 59.260 128.895 ;
        RECT 59.440 127.960 59.690 129.095 ;
        RECT 62.630 128.925 63.600 129.515 ;
        RECT 65.395 129.095 65.745 129.345 ;
        RECT 59.860 127.785 60.120 128.895 ;
        RECT 60.290 128.685 63.600 128.925 ;
        RECT 60.290 127.960 60.550 128.685 ;
        RECT 60.720 127.785 60.980 128.515 ;
        RECT 61.150 127.960 61.410 128.685 ;
        RECT 61.580 127.785 61.840 128.515 ;
        RECT 62.010 127.960 62.270 128.685 ;
        RECT 62.440 127.785 62.700 128.515 ;
        RECT 62.870 127.960 63.130 128.685 ;
        RECT 63.300 127.785 63.595 128.515 ;
        RECT 64.935 127.785 65.225 128.950 ;
        RECT 65.915 128.925 66.085 129.525 ;
        RECT 66.255 129.095 66.605 129.345 ;
        RECT 66.775 129.045 67.295 129.585 ;
        RECT 68.155 129.535 68.850 130.165 ;
        RECT 69.055 129.535 69.365 130.335 ;
        RECT 69.995 129.535 70.305 130.335 ;
        RECT 70.510 129.535 71.205 130.165 ;
        RECT 71.375 129.790 76.720 130.335 ;
        RECT 65.405 127.785 65.735 128.925 ;
        RECT 65.915 128.755 66.595 128.925 ;
        RECT 67.465 128.875 67.985 129.415 ;
        RECT 68.175 129.095 68.510 129.345 ;
        RECT 68.680 128.935 68.850 129.535 ;
        RECT 69.020 129.095 69.355 129.365 ;
        RECT 70.005 129.095 70.340 129.365 ;
        RECT 70.510 128.935 70.680 129.535 ;
        RECT 70.850 129.095 71.185 129.345 ;
        RECT 72.960 128.960 73.300 129.790 ;
        RECT 76.895 129.565 78.565 130.335 ;
        RECT 66.265 127.970 66.595 128.755 ;
        RECT 66.775 127.785 67.985 128.875 ;
        RECT 68.155 127.785 68.415 128.925 ;
        RECT 68.585 127.955 68.915 128.935 ;
        RECT 69.085 127.785 69.365 128.925 ;
        RECT 69.995 127.785 70.275 128.925 ;
        RECT 70.445 127.955 70.775 128.935 ;
        RECT 70.945 127.785 71.205 128.925 ;
        RECT 74.780 128.220 75.130 129.470 ;
        RECT 76.895 129.045 77.645 129.565 ;
        RECT 79.235 129.515 79.465 130.335 ;
        RECT 79.635 129.535 79.965 130.165 ;
        RECT 77.815 128.875 78.565 129.395 ;
        RECT 79.215 129.095 79.545 129.345 ;
        RECT 79.715 128.935 79.965 129.535 ;
        RECT 80.135 129.515 80.345 130.335 ;
        RECT 80.575 129.515 80.835 130.335 ;
        RECT 81.005 129.515 81.335 129.935 ;
        RECT 81.515 129.765 81.775 130.165 ;
        RECT 81.945 129.935 82.275 130.335 ;
        RECT 82.445 129.765 82.615 130.115 ;
        RECT 82.785 129.935 83.160 130.335 ;
        RECT 81.515 129.595 83.180 129.765 ;
        RECT 83.350 129.660 83.625 130.005 ;
        RECT 81.085 129.425 81.335 129.515 ;
        RECT 83.010 129.425 83.180 129.595 ;
        RECT 80.580 129.095 80.915 129.345 ;
        RECT 81.085 129.095 81.800 129.425 ;
        RECT 82.015 129.095 82.840 129.425 ;
        RECT 83.010 129.095 83.285 129.425 ;
        RECT 71.375 127.785 76.720 128.220 ;
        RECT 76.895 127.785 78.565 128.875 ;
        RECT 79.235 127.785 79.465 128.925 ;
        RECT 79.635 127.955 79.965 128.935 ;
        RECT 80.135 127.785 80.345 128.925 ;
        RECT 80.575 127.785 80.835 128.925 ;
        RECT 81.085 128.535 81.255 129.095 ;
        RECT 81.515 128.635 81.845 128.925 ;
        RECT 82.015 128.805 82.260 129.095 ;
        RECT 83.010 128.925 83.180 129.095 ;
        RECT 83.455 128.925 83.625 129.660 ;
        RECT 82.520 128.755 83.180 128.925 ;
        RECT 82.520 128.635 82.690 128.755 ;
        RECT 81.515 128.465 82.690 128.635 ;
        RECT 81.075 127.965 82.690 128.295 ;
        RECT 82.860 127.785 83.140 128.585 ;
        RECT 83.350 127.955 83.625 128.925 ;
        RECT 84.720 129.595 84.975 130.165 ;
        RECT 85.145 129.935 85.475 130.335 ;
        RECT 85.900 129.800 86.430 130.165 ;
        RECT 85.900 129.765 86.075 129.800 ;
        RECT 85.145 129.595 86.075 129.765 ;
        RECT 84.720 128.925 84.890 129.595 ;
        RECT 85.145 129.425 85.315 129.595 ;
        RECT 85.060 129.095 85.315 129.425 ;
        RECT 85.540 129.095 85.735 129.425 ;
        RECT 84.720 127.955 85.055 128.925 ;
        RECT 85.225 127.785 85.395 128.925 ;
        RECT 85.565 128.125 85.735 129.095 ;
        RECT 85.905 128.465 86.075 129.595 ;
        RECT 86.245 128.805 86.415 129.605 ;
        RECT 86.620 129.315 86.895 130.165 ;
        RECT 86.615 129.145 86.895 129.315 ;
        RECT 86.620 129.005 86.895 129.145 ;
        RECT 87.065 128.805 87.255 130.165 ;
        RECT 87.435 129.800 87.945 130.335 ;
        RECT 88.165 129.525 88.410 130.130 ;
        RECT 88.855 129.565 90.525 130.335 ;
        RECT 90.695 129.610 90.985 130.335 ;
        RECT 91.155 129.790 96.500 130.335 ;
        RECT 87.455 129.355 88.685 129.525 ;
        RECT 86.245 128.635 87.255 128.805 ;
        RECT 87.425 128.790 88.175 128.980 ;
        RECT 85.905 128.295 87.030 128.465 ;
        RECT 87.425 128.125 87.595 128.790 ;
        RECT 88.345 128.545 88.685 129.355 ;
        RECT 88.855 129.045 89.605 129.565 ;
        RECT 89.775 128.875 90.525 129.395 ;
        RECT 92.740 128.960 93.080 129.790 ;
        RECT 97.600 129.595 97.855 130.165 ;
        RECT 98.025 129.935 98.355 130.335 ;
        RECT 98.780 129.800 99.310 130.165 ;
        RECT 98.780 129.765 98.955 129.800 ;
        RECT 98.025 129.595 98.955 129.765 ;
        RECT 85.565 127.955 87.595 128.125 ;
        RECT 87.765 127.785 87.935 128.545 ;
        RECT 88.170 128.135 88.685 128.545 ;
        RECT 88.855 127.785 90.525 128.875 ;
        RECT 90.695 127.785 90.985 128.950 ;
        RECT 94.560 128.220 94.910 129.470 ;
        RECT 97.600 128.925 97.770 129.595 ;
        RECT 98.025 129.425 98.195 129.595 ;
        RECT 97.940 129.095 98.195 129.425 ;
        RECT 98.420 129.095 98.615 129.425 ;
        RECT 91.155 127.785 96.500 128.220 ;
        RECT 97.600 127.955 97.935 128.925 ;
        RECT 98.105 127.785 98.275 128.925 ;
        RECT 98.445 128.125 98.615 129.095 ;
        RECT 98.785 128.465 98.955 129.595 ;
        RECT 99.125 128.805 99.295 129.605 ;
        RECT 99.500 129.315 99.775 130.165 ;
        RECT 99.495 129.145 99.775 129.315 ;
        RECT 99.500 129.005 99.775 129.145 ;
        RECT 99.945 128.805 100.135 130.165 ;
        RECT 100.315 129.800 100.825 130.335 ;
        RECT 101.045 129.525 101.290 130.130 ;
        RECT 101.735 129.790 107.080 130.335 ;
        RECT 107.255 129.790 112.600 130.335 ;
        RECT 100.335 129.355 101.565 129.525 ;
        RECT 99.125 128.635 100.135 128.805 ;
        RECT 100.305 128.790 101.055 128.980 ;
        RECT 98.785 128.295 99.910 128.465 ;
        RECT 100.305 128.125 100.475 128.790 ;
        RECT 101.225 128.545 101.565 129.355 ;
        RECT 103.320 128.960 103.660 129.790 ;
        RECT 98.445 127.955 100.475 128.125 ;
        RECT 100.645 127.785 100.815 128.545 ;
        RECT 101.050 128.135 101.565 128.545 ;
        RECT 105.140 128.220 105.490 129.470 ;
        RECT 108.840 128.960 109.180 129.790 ;
        RECT 112.775 129.535 113.115 130.165 ;
        RECT 113.285 129.535 113.535 130.335 ;
        RECT 113.725 129.685 114.055 130.165 ;
        RECT 114.225 129.875 114.450 130.335 ;
        RECT 114.620 129.685 114.950 130.165 ;
        RECT 110.660 128.220 111.010 129.470 ;
        RECT 112.775 128.925 112.950 129.535 ;
        RECT 113.725 129.515 114.950 129.685 ;
        RECT 115.580 129.555 116.080 130.165 ;
        RECT 116.455 129.610 116.745 130.335 ;
        RECT 116.950 129.595 117.565 130.165 ;
        RECT 117.735 129.825 117.950 130.335 ;
        RECT 118.180 129.825 118.460 130.155 ;
        RECT 118.640 129.825 118.880 130.335 ;
        RECT 113.120 129.175 113.815 129.345 ;
        RECT 113.645 128.925 113.815 129.175 ;
        RECT 113.990 129.145 114.410 129.345 ;
        RECT 114.580 129.145 114.910 129.345 ;
        RECT 115.080 129.145 115.410 129.345 ;
        RECT 115.580 128.925 115.750 129.555 ;
        RECT 115.935 129.095 116.285 129.345 ;
        RECT 101.735 127.785 107.080 128.220 ;
        RECT 107.255 127.785 112.600 128.220 ;
        RECT 112.775 127.955 113.115 128.925 ;
        RECT 113.285 127.785 113.455 128.925 ;
        RECT 113.645 128.755 116.080 128.925 ;
        RECT 113.725 127.785 113.975 128.585 ;
        RECT 114.620 127.955 114.950 128.755 ;
        RECT 115.250 127.785 115.580 128.585 ;
        RECT 115.750 127.955 116.080 128.755 ;
        RECT 116.455 127.785 116.745 128.950 ;
        RECT 116.950 128.575 117.265 129.595 ;
        RECT 117.435 128.925 117.605 129.425 ;
        RECT 117.855 129.095 118.120 129.655 ;
        RECT 118.290 128.925 118.460 129.825 ;
        RECT 119.215 129.790 124.560 130.335 ;
        RECT 118.630 129.095 118.985 129.655 ;
        RECT 120.800 128.960 121.140 129.790 ;
        RECT 124.940 129.555 125.440 130.165 ;
        RECT 117.435 128.755 118.860 128.925 ;
        RECT 116.950 127.955 117.485 128.575 ;
        RECT 117.655 127.785 117.985 128.585 ;
        RECT 118.470 128.580 118.860 128.755 ;
        RECT 122.620 128.220 122.970 129.470 ;
        RECT 124.735 129.095 125.085 129.345 ;
        RECT 125.270 128.925 125.440 129.555 ;
        RECT 126.070 129.685 126.400 130.165 ;
        RECT 126.570 129.875 126.795 130.335 ;
        RECT 126.965 129.685 127.295 130.165 ;
        RECT 126.070 129.515 127.295 129.685 ;
        RECT 127.485 129.535 127.735 130.335 ;
        RECT 127.905 129.535 128.245 130.165 ;
        RECT 128.505 129.785 128.675 130.075 ;
        RECT 128.845 129.955 129.175 130.335 ;
        RECT 128.505 129.615 129.170 129.785 ;
        RECT 128.015 129.485 128.245 129.535 ;
        RECT 125.610 129.145 125.940 129.345 ;
        RECT 126.110 129.145 126.440 129.345 ;
        RECT 126.610 129.145 127.030 129.345 ;
        RECT 127.205 129.175 127.900 129.345 ;
        RECT 127.205 128.925 127.375 129.175 ;
        RECT 128.070 128.925 128.245 129.485 ;
        RECT 124.940 128.755 127.375 128.925 ;
        RECT 119.215 127.785 124.560 128.220 ;
        RECT 124.940 127.955 125.270 128.755 ;
        RECT 125.440 127.785 125.770 128.585 ;
        RECT 126.070 127.955 126.400 128.755 ;
        RECT 127.045 127.785 127.295 128.585 ;
        RECT 127.565 127.785 127.735 128.925 ;
        RECT 127.905 127.955 128.245 128.925 ;
        RECT 128.420 128.795 128.770 129.445 ;
        RECT 128.940 128.625 129.170 129.615 ;
        RECT 128.505 128.455 129.170 128.625 ;
        RECT 128.505 127.955 128.675 128.455 ;
        RECT 128.845 127.785 129.175 128.285 ;
        RECT 129.345 127.955 129.530 130.075 ;
        RECT 129.785 129.875 130.035 130.335 ;
        RECT 130.205 129.885 130.540 130.055 ;
        RECT 130.735 129.885 131.410 130.055 ;
        RECT 130.205 129.745 130.375 129.885 ;
        RECT 129.700 128.755 129.980 129.705 ;
        RECT 130.150 129.615 130.375 129.745 ;
        RECT 130.150 128.510 130.320 129.615 ;
        RECT 130.545 129.465 131.070 129.685 ;
        RECT 130.490 128.700 130.730 129.295 ;
        RECT 130.900 128.765 131.070 129.465 ;
        RECT 131.240 129.105 131.410 129.885 ;
        RECT 131.730 129.835 132.100 130.335 ;
        RECT 132.280 129.885 132.685 130.055 ;
        RECT 132.855 129.885 133.640 130.055 ;
        RECT 132.280 129.655 132.450 129.885 ;
        RECT 131.620 129.355 132.450 129.655 ;
        RECT 132.835 129.385 133.300 129.715 ;
        RECT 131.620 129.325 131.820 129.355 ;
        RECT 131.940 129.105 132.110 129.175 ;
        RECT 131.240 128.935 132.110 129.105 ;
        RECT 131.600 128.845 132.110 128.935 ;
        RECT 130.150 128.380 130.455 128.510 ;
        RECT 130.900 128.400 131.430 128.765 ;
        RECT 129.770 127.785 130.035 128.245 ;
        RECT 130.205 127.955 130.455 128.380 ;
        RECT 131.600 128.230 131.770 128.845 ;
        RECT 130.665 128.060 131.770 128.230 ;
        RECT 131.940 127.785 132.110 128.585 ;
        RECT 132.280 128.285 132.450 129.355 ;
        RECT 132.620 128.455 132.810 129.175 ;
        RECT 132.980 128.425 133.300 129.385 ;
        RECT 133.470 129.425 133.640 129.885 ;
        RECT 133.915 129.805 134.125 130.335 ;
        RECT 134.385 129.595 134.715 130.120 ;
        RECT 134.885 129.725 135.055 130.335 ;
        RECT 135.225 129.680 135.555 130.115 ;
        RECT 135.865 129.785 136.035 130.165 ;
        RECT 136.250 129.955 136.580 130.335 ;
        RECT 135.225 129.595 135.605 129.680 ;
        RECT 135.865 129.615 136.580 129.785 ;
        RECT 134.515 129.425 134.715 129.595 ;
        RECT 135.380 129.555 135.605 129.595 ;
        RECT 133.470 129.095 134.345 129.425 ;
        RECT 134.515 129.095 135.265 129.425 ;
        RECT 132.280 127.955 132.530 128.285 ;
        RECT 133.470 128.255 133.640 129.095 ;
        RECT 134.515 128.890 134.705 129.095 ;
        RECT 135.435 128.975 135.605 129.555 ;
        RECT 135.775 129.065 136.130 129.435 ;
        RECT 136.410 129.425 136.580 129.615 ;
        RECT 136.750 129.590 137.005 130.165 ;
        RECT 136.410 129.095 136.665 129.425 ;
        RECT 135.390 128.925 135.605 128.975 ;
        RECT 133.810 128.515 134.705 128.890 ;
        RECT 135.215 128.845 135.605 128.925 ;
        RECT 136.410 128.885 136.580 129.095 ;
        RECT 132.755 128.085 133.640 128.255 ;
        RECT 133.820 127.785 134.135 128.285 ;
        RECT 134.365 127.955 134.705 128.515 ;
        RECT 134.875 127.785 135.045 128.795 ;
        RECT 135.215 128.000 135.545 128.845 ;
        RECT 135.865 128.715 136.580 128.885 ;
        RECT 136.835 128.860 137.005 129.590 ;
        RECT 137.180 129.495 137.440 130.335 ;
        RECT 137.615 129.585 138.825 130.335 ;
        RECT 135.865 127.955 136.035 128.715 ;
        RECT 136.250 127.785 136.580 128.545 ;
        RECT 136.750 127.955 137.005 128.860 ;
        RECT 137.180 127.785 137.440 128.935 ;
        RECT 137.615 128.875 138.135 129.415 ;
        RECT 138.305 129.045 138.825 129.585 ;
        RECT 137.615 127.785 138.825 128.875 ;
        RECT 13.330 127.615 138.910 127.785 ;
        RECT 13.415 126.525 14.625 127.615 ;
        RECT 14.795 127.180 20.140 127.615 ;
        RECT 13.415 125.815 13.935 126.355 ;
        RECT 14.105 125.985 14.625 126.525 ;
        RECT 13.415 125.065 14.625 125.815 ;
        RECT 16.380 125.610 16.720 126.440 ;
        RECT 18.200 125.930 18.550 127.180 ;
        RECT 20.315 126.525 22.905 127.615 ;
        RECT 20.315 125.835 21.525 126.355 ;
        RECT 21.695 126.005 22.905 126.525 ;
        RECT 23.665 126.445 23.995 127.615 ;
        RECT 24.195 126.275 24.525 127.445 ;
        RECT 24.725 126.445 25.055 127.615 ;
        RECT 25.255 126.275 25.615 127.445 ;
        RECT 25.785 126.475 26.115 127.615 ;
        RECT 26.295 126.450 26.585 127.615 ;
        RECT 27.005 126.885 27.300 127.615 ;
        RECT 27.470 126.715 27.730 127.440 ;
        RECT 27.900 126.885 28.160 127.615 ;
        RECT 28.330 126.715 28.590 127.440 ;
        RECT 28.760 126.885 29.020 127.615 ;
        RECT 29.190 126.715 29.450 127.440 ;
        RECT 29.620 126.885 29.880 127.615 ;
        RECT 30.050 126.715 30.310 127.440 ;
        RECT 27.000 126.475 30.310 126.715 ;
        RECT 30.480 126.505 30.740 127.615 ;
        RECT 24.195 125.995 25.615 126.275 ;
        RECT 14.795 125.065 20.140 125.610 ;
        RECT 20.315 125.065 22.905 125.835 ;
        RECT 24.205 125.065 24.535 125.755 ;
        RECT 25.255 125.660 25.615 125.995 ;
        RECT 25.785 125.725 26.125 126.305 ;
        RECT 27.000 125.885 27.970 126.475 ;
        RECT 30.910 126.305 31.160 127.440 ;
        RECT 31.340 126.505 31.635 127.615 ;
        RECT 31.815 127.180 37.160 127.615 ;
        RECT 37.335 127.180 42.680 127.615 ;
        RECT 42.855 127.180 48.200 127.615 ;
        RECT 28.140 126.055 31.160 126.305 ;
        RECT 24.995 125.235 25.615 125.660 ;
        RECT 25.785 125.065 26.115 125.555 ;
        RECT 26.295 125.065 26.585 125.790 ;
        RECT 27.000 125.715 30.310 125.885 ;
        RECT 27.000 125.065 27.300 125.545 ;
        RECT 27.470 125.260 27.730 125.715 ;
        RECT 27.900 125.065 28.160 125.545 ;
        RECT 28.330 125.260 28.590 125.715 ;
        RECT 28.760 125.065 29.020 125.545 ;
        RECT 29.190 125.260 29.450 125.715 ;
        RECT 29.620 125.065 29.880 125.545 ;
        RECT 30.050 125.260 30.310 125.715 ;
        RECT 30.480 125.065 30.740 125.590 ;
        RECT 30.910 125.245 31.160 126.055 ;
        RECT 31.330 125.695 31.645 126.305 ;
        RECT 33.400 125.610 33.740 126.440 ;
        RECT 35.220 125.930 35.570 127.180 ;
        RECT 38.920 125.610 39.260 126.440 ;
        RECT 40.740 125.930 41.090 127.180 ;
        RECT 44.440 125.610 44.780 126.440 ;
        RECT 46.260 125.930 46.610 127.180 ;
        RECT 48.375 126.525 51.885 127.615 ;
        RECT 48.375 125.835 50.025 126.355 ;
        RECT 50.195 126.005 51.885 126.525 ;
        RECT 52.055 126.450 52.345 127.615 ;
        RECT 52.515 126.525 56.025 127.615 ;
        RECT 52.515 125.835 54.165 126.355 ;
        RECT 54.335 126.005 56.025 126.525 ;
        RECT 56.205 126.645 56.535 127.430 ;
        RECT 56.205 126.475 56.885 126.645 ;
        RECT 57.065 126.475 57.395 127.615 ;
        RECT 57.575 126.525 58.785 127.615 ;
        RECT 56.195 126.055 56.545 126.305 ;
        RECT 56.715 125.875 56.885 126.475 ;
        RECT 57.055 126.055 57.405 126.305 ;
        RECT 31.340 125.065 31.585 125.525 ;
        RECT 31.815 125.065 37.160 125.610 ;
        RECT 37.335 125.065 42.680 125.610 ;
        RECT 42.855 125.065 48.200 125.610 ;
        RECT 48.375 125.065 51.885 125.835 ;
        RECT 52.055 125.065 52.345 125.790 ;
        RECT 52.515 125.065 56.025 125.835 ;
        RECT 56.215 125.065 56.455 125.875 ;
        RECT 56.625 125.235 56.955 125.875 ;
        RECT 57.125 125.065 57.395 125.875 ;
        RECT 57.575 125.815 58.095 126.355 ;
        RECT 58.265 125.985 58.785 126.525 ;
        RECT 58.965 126.595 59.295 127.445 ;
        RECT 59.465 126.765 59.635 127.615 ;
        RECT 59.805 126.595 60.135 127.445 ;
        RECT 60.305 126.765 60.475 127.615 ;
        RECT 60.645 126.595 60.975 127.445 ;
        RECT 61.145 126.815 61.315 127.615 ;
        RECT 61.485 126.595 61.815 127.445 ;
        RECT 61.985 126.815 62.155 127.615 ;
        RECT 62.325 126.595 62.655 127.445 ;
        RECT 62.825 126.815 62.995 127.615 ;
        RECT 63.165 126.595 63.495 127.445 ;
        RECT 63.665 126.815 63.835 127.615 ;
        RECT 64.005 126.595 64.335 127.445 ;
        RECT 64.505 126.815 64.675 127.615 ;
        RECT 64.845 126.595 65.175 127.445 ;
        RECT 65.345 126.815 65.515 127.615 ;
        RECT 65.685 126.595 66.015 127.445 ;
        RECT 66.185 126.815 66.355 127.615 ;
        RECT 66.525 126.595 66.855 127.445 ;
        RECT 67.025 126.815 67.195 127.615 ;
        RECT 67.365 126.595 67.695 127.445 ;
        RECT 67.865 126.815 68.035 127.615 ;
        RECT 68.205 126.595 68.535 127.445 ;
        RECT 68.705 126.815 68.875 127.615 ;
        RECT 69.045 126.595 69.375 127.445 ;
        RECT 69.545 126.815 69.715 127.615 ;
        RECT 58.965 126.425 60.475 126.595 ;
        RECT 60.645 126.425 62.995 126.595 ;
        RECT 63.165 126.425 69.825 126.595 ;
        RECT 69.995 126.525 71.205 127.615 ;
        RECT 60.305 126.255 60.475 126.425 ;
        RECT 62.820 126.255 62.995 126.425 ;
        RECT 58.960 126.055 60.135 126.255 ;
        RECT 60.305 126.055 62.615 126.255 ;
        RECT 62.820 126.055 69.380 126.255 ;
        RECT 60.305 125.885 60.475 126.055 ;
        RECT 62.820 125.885 62.995 126.055 ;
        RECT 69.550 125.885 69.825 126.425 ;
        RECT 57.575 125.065 58.785 125.815 ;
        RECT 58.965 125.715 60.475 125.885 ;
        RECT 60.645 125.715 62.995 125.885 ;
        RECT 63.165 125.715 69.825 125.885 ;
        RECT 69.995 125.815 70.515 126.355 ;
        RECT 70.685 125.985 71.205 126.525 ;
        RECT 71.375 126.475 71.760 127.445 ;
        RECT 71.930 127.155 72.255 127.615 ;
        RECT 72.775 126.985 73.055 127.445 ;
        RECT 71.930 126.765 73.055 126.985 ;
        RECT 58.965 125.240 59.295 125.715 ;
        RECT 59.465 125.065 59.635 125.545 ;
        RECT 59.805 125.240 60.135 125.715 ;
        RECT 60.305 125.065 60.475 125.545 ;
        RECT 60.645 125.240 60.975 125.715 ;
        RECT 61.145 125.065 61.315 125.545 ;
        RECT 61.485 125.240 61.815 125.715 ;
        RECT 61.985 125.065 62.155 125.545 ;
        RECT 62.325 125.240 62.655 125.715 ;
        RECT 62.825 125.065 62.995 125.545 ;
        RECT 63.165 125.240 63.495 125.715 ;
        RECT 63.165 125.235 63.415 125.240 ;
        RECT 63.665 125.065 63.835 125.545 ;
        RECT 64.005 125.240 64.335 125.715 ;
        RECT 64.085 125.235 64.255 125.240 ;
        RECT 64.505 125.065 64.675 125.545 ;
        RECT 64.845 125.240 65.175 125.715 ;
        RECT 64.925 125.235 65.095 125.240 ;
        RECT 65.345 125.065 65.515 125.545 ;
        RECT 65.685 125.240 66.015 125.715 ;
        RECT 66.185 125.065 66.355 125.545 ;
        RECT 66.525 125.240 66.855 125.715 ;
        RECT 67.025 125.065 67.195 125.545 ;
        RECT 67.365 125.240 67.695 125.715 ;
        RECT 67.865 125.065 68.035 125.545 ;
        RECT 68.205 125.240 68.535 125.715 ;
        RECT 68.705 125.065 68.875 125.545 ;
        RECT 69.045 125.240 69.375 125.715 ;
        RECT 69.545 125.065 69.715 125.545 ;
        RECT 69.995 125.065 71.205 125.815 ;
        RECT 71.375 125.805 71.655 126.475 ;
        RECT 71.930 126.305 72.380 126.765 ;
        RECT 73.245 126.595 73.645 127.445 ;
        RECT 74.045 127.155 74.315 127.615 ;
        RECT 74.485 126.985 74.770 127.445 ;
        RECT 71.825 125.975 72.380 126.305 ;
        RECT 72.550 126.035 73.645 126.595 ;
        RECT 71.930 125.865 72.380 125.975 ;
        RECT 71.375 125.235 71.760 125.805 ;
        RECT 71.930 125.695 73.055 125.865 ;
        RECT 71.930 125.065 72.255 125.525 ;
        RECT 72.775 125.235 73.055 125.695 ;
        RECT 73.245 125.235 73.645 126.035 ;
        RECT 73.815 126.765 74.770 126.985 ;
        RECT 73.815 125.865 74.025 126.765 ;
        RECT 75.055 126.745 75.330 127.445 ;
        RECT 75.500 127.070 75.755 127.615 ;
        RECT 75.925 127.105 76.405 127.445 ;
        RECT 76.580 127.060 77.185 127.615 ;
        RECT 76.570 126.960 77.185 127.060 ;
        RECT 76.570 126.935 76.755 126.960 ;
        RECT 74.195 126.035 74.885 126.595 ;
        RECT 73.815 125.695 74.770 125.865 ;
        RECT 74.045 125.065 74.315 125.525 ;
        RECT 74.485 125.235 74.770 125.695 ;
        RECT 75.055 125.715 75.225 126.745 ;
        RECT 75.500 126.615 76.255 126.865 ;
        RECT 76.425 126.690 76.755 126.935 ;
        RECT 75.500 126.580 76.270 126.615 ;
        RECT 75.500 126.570 76.285 126.580 ;
        RECT 75.395 126.555 76.290 126.570 ;
        RECT 75.395 126.540 76.310 126.555 ;
        RECT 75.395 126.530 76.330 126.540 ;
        RECT 75.395 126.520 76.355 126.530 ;
        RECT 75.395 126.490 76.425 126.520 ;
        RECT 75.395 126.460 76.445 126.490 ;
        RECT 75.395 126.430 76.465 126.460 ;
        RECT 75.395 126.405 76.495 126.430 ;
        RECT 75.395 126.370 76.530 126.405 ;
        RECT 75.395 126.365 76.560 126.370 ;
        RECT 75.395 125.970 75.625 126.365 ;
        RECT 76.170 126.360 76.560 126.365 ;
        RECT 76.195 126.350 76.560 126.360 ;
        RECT 76.210 126.345 76.560 126.350 ;
        RECT 76.225 126.340 76.560 126.345 ;
        RECT 76.925 126.340 77.185 126.790 ;
        RECT 77.815 126.450 78.105 127.615 ;
        RECT 78.275 127.105 79.465 127.395 ;
        RECT 78.295 126.765 79.465 126.935 ;
        RECT 79.635 126.815 79.915 127.615 ;
        RECT 78.295 126.475 78.620 126.765 ;
        RECT 79.295 126.645 79.465 126.765 ;
        RECT 76.225 126.335 77.185 126.340 ;
        RECT 76.235 126.325 77.185 126.335 ;
        RECT 76.245 126.320 77.185 126.325 ;
        RECT 76.255 126.310 77.185 126.320 ;
        RECT 76.260 126.300 77.185 126.310 ;
        RECT 78.790 126.305 78.985 126.595 ;
        RECT 79.295 126.475 79.955 126.645 ;
        RECT 80.125 126.475 80.400 127.445 ;
        RECT 81.035 126.475 81.295 127.615 ;
        RECT 81.535 127.105 83.150 127.435 ;
        RECT 79.785 126.305 79.955 126.475 ;
        RECT 76.265 126.295 77.185 126.300 ;
        RECT 76.275 126.280 77.185 126.295 ;
        RECT 76.280 126.265 77.185 126.280 ;
        RECT 76.290 126.240 77.185 126.265 ;
        RECT 75.795 125.770 76.125 126.195 ;
        RECT 75.875 125.745 76.125 125.770 ;
        RECT 75.055 125.235 75.315 125.715 ;
        RECT 75.485 125.065 75.735 125.605 ;
        RECT 75.905 125.285 76.125 125.745 ;
        RECT 76.295 126.170 77.185 126.240 ;
        RECT 76.295 125.445 76.465 126.170 ;
        RECT 76.635 125.615 77.185 126.000 ;
        RECT 78.275 125.975 78.620 126.305 ;
        RECT 78.790 125.975 79.615 126.305 ;
        RECT 79.785 125.975 80.060 126.305 ;
        RECT 79.785 125.805 79.955 125.975 ;
        RECT 76.295 125.275 77.185 125.445 ;
        RECT 77.815 125.065 78.105 125.790 ;
        RECT 78.290 125.635 79.955 125.805 ;
        RECT 80.230 125.740 80.400 126.475 ;
        RECT 81.545 126.305 81.715 126.865 ;
        RECT 81.975 126.765 83.150 126.935 ;
        RECT 83.320 126.815 83.600 127.615 ;
        RECT 81.975 126.475 82.305 126.765 ;
        RECT 82.980 126.645 83.150 126.765 ;
        RECT 82.475 126.305 82.720 126.595 ;
        RECT 82.980 126.475 83.640 126.645 ;
        RECT 83.810 126.475 84.085 127.445 ;
        RECT 83.470 126.305 83.640 126.475 ;
        RECT 81.040 126.055 81.375 126.305 ;
        RECT 81.545 125.975 82.260 126.305 ;
        RECT 82.475 125.975 83.300 126.305 ;
        RECT 83.470 125.975 83.745 126.305 ;
        RECT 81.545 125.885 81.795 125.975 ;
        RECT 78.290 125.285 78.545 125.635 ;
        RECT 78.715 125.065 79.045 125.465 ;
        RECT 79.215 125.285 79.385 125.635 ;
        RECT 79.555 125.065 79.935 125.465 ;
        RECT 80.125 125.395 80.400 125.740 ;
        RECT 81.035 125.065 81.295 125.885 ;
        RECT 81.465 125.465 81.795 125.885 ;
        RECT 83.470 125.805 83.640 125.975 ;
        RECT 81.975 125.635 83.640 125.805 ;
        RECT 83.915 125.740 84.085 126.475 ;
        RECT 81.975 125.235 82.235 125.635 ;
        RECT 82.405 125.065 82.735 125.465 ;
        RECT 82.905 125.285 83.075 125.635 ;
        RECT 83.245 125.065 83.620 125.465 ;
        RECT 83.810 125.395 84.085 125.740 ;
        RECT 84.720 126.475 85.055 127.445 ;
        RECT 85.225 126.475 85.395 127.615 ;
        RECT 85.565 127.275 87.595 127.445 ;
        RECT 84.720 125.805 84.890 126.475 ;
        RECT 85.565 126.305 85.735 127.275 ;
        RECT 85.060 125.975 85.315 126.305 ;
        RECT 85.540 125.975 85.735 126.305 ;
        RECT 85.905 126.935 87.030 127.105 ;
        RECT 85.145 125.805 85.315 125.975 ;
        RECT 85.905 125.805 86.075 126.935 ;
        RECT 84.720 125.235 84.975 125.805 ;
        RECT 85.145 125.635 86.075 125.805 ;
        RECT 86.245 126.595 87.255 126.765 ;
        RECT 86.245 125.795 86.415 126.595 ;
        RECT 86.620 125.915 86.895 126.395 ;
        RECT 86.615 125.745 86.895 125.915 ;
        RECT 85.900 125.600 86.075 125.635 ;
        RECT 85.145 125.065 85.475 125.465 ;
        RECT 85.900 125.235 86.430 125.600 ;
        RECT 86.620 125.235 86.895 125.745 ;
        RECT 87.065 125.235 87.255 126.595 ;
        RECT 87.425 126.610 87.595 127.275 ;
        RECT 87.765 126.855 87.935 127.615 ;
        RECT 88.170 126.855 88.685 127.265 ;
        RECT 88.855 127.180 94.200 127.615 ;
        RECT 87.425 126.420 88.175 126.610 ;
        RECT 88.345 126.045 88.685 126.855 ;
        RECT 87.455 125.875 88.685 126.045 ;
        RECT 87.435 125.065 87.945 125.600 ;
        RECT 88.165 125.270 88.410 125.875 ;
        RECT 90.440 125.610 90.780 126.440 ;
        RECT 92.260 125.930 92.610 127.180 ;
        RECT 94.375 126.525 95.585 127.615 ;
        RECT 95.845 126.945 96.015 127.445 ;
        RECT 96.185 127.115 96.515 127.615 ;
        RECT 95.845 126.775 96.510 126.945 ;
        RECT 94.375 125.815 94.895 126.355 ;
        RECT 95.065 125.985 95.585 126.525 ;
        RECT 95.760 125.955 96.110 126.605 ;
        RECT 88.855 125.065 94.200 125.610 ;
        RECT 94.375 125.065 95.585 125.815 ;
        RECT 96.280 125.785 96.510 126.775 ;
        RECT 95.845 125.615 96.510 125.785 ;
        RECT 95.845 125.325 96.015 125.615 ;
        RECT 96.185 125.065 96.515 125.445 ;
        RECT 96.685 125.325 96.870 127.445 ;
        RECT 97.110 127.155 97.375 127.615 ;
        RECT 97.545 127.020 97.795 127.445 ;
        RECT 98.005 127.170 99.110 127.340 ;
        RECT 97.490 126.890 97.795 127.020 ;
        RECT 97.040 125.695 97.320 126.645 ;
        RECT 97.490 125.785 97.660 126.890 ;
        RECT 97.830 126.105 98.070 126.700 ;
        RECT 98.240 126.635 98.770 127.000 ;
        RECT 98.240 125.935 98.410 126.635 ;
        RECT 98.940 126.555 99.110 127.170 ;
        RECT 99.280 126.815 99.450 127.615 ;
        RECT 99.620 127.115 99.870 127.445 ;
        RECT 100.095 127.145 100.980 127.315 ;
        RECT 98.940 126.465 99.450 126.555 ;
        RECT 97.490 125.655 97.715 125.785 ;
        RECT 97.885 125.715 98.410 125.935 ;
        RECT 98.580 126.295 99.450 126.465 ;
        RECT 97.125 125.065 97.375 125.525 ;
        RECT 97.545 125.515 97.715 125.655 ;
        RECT 98.580 125.515 98.750 126.295 ;
        RECT 99.280 126.225 99.450 126.295 ;
        RECT 98.960 126.045 99.160 126.075 ;
        RECT 99.620 126.045 99.790 127.115 ;
        RECT 99.960 126.225 100.150 126.945 ;
        RECT 98.960 125.745 99.790 126.045 ;
        RECT 100.320 126.015 100.640 126.975 ;
        RECT 97.545 125.345 97.880 125.515 ;
        RECT 98.075 125.345 98.750 125.515 ;
        RECT 99.070 125.065 99.440 125.565 ;
        RECT 99.620 125.515 99.790 125.745 ;
        RECT 100.175 125.685 100.640 126.015 ;
        RECT 100.810 126.305 100.980 127.145 ;
        RECT 101.160 127.115 101.475 127.615 ;
        RECT 101.705 126.885 102.045 127.445 ;
        RECT 101.150 126.510 102.045 126.885 ;
        RECT 102.215 126.605 102.385 127.615 ;
        RECT 101.855 126.305 102.045 126.510 ;
        RECT 102.555 126.555 102.885 127.400 ;
        RECT 102.555 126.475 102.945 126.555 ;
        RECT 102.730 126.425 102.945 126.475 ;
        RECT 103.575 126.450 103.865 127.615 ;
        RECT 104.040 126.475 104.375 127.445 ;
        RECT 104.545 126.475 104.715 127.615 ;
        RECT 104.885 127.275 106.915 127.445 ;
        RECT 100.810 125.975 101.685 126.305 ;
        RECT 101.855 125.975 102.605 126.305 ;
        RECT 100.810 125.515 100.980 125.975 ;
        RECT 101.855 125.805 102.055 125.975 ;
        RECT 102.775 125.845 102.945 126.425 ;
        RECT 102.720 125.805 102.945 125.845 ;
        RECT 99.620 125.345 100.025 125.515 ;
        RECT 100.195 125.345 100.980 125.515 ;
        RECT 101.255 125.065 101.465 125.595 ;
        RECT 101.725 125.280 102.055 125.805 ;
        RECT 102.565 125.720 102.945 125.805 ;
        RECT 104.040 125.805 104.210 126.475 ;
        RECT 104.885 126.305 105.055 127.275 ;
        RECT 104.380 125.975 104.635 126.305 ;
        RECT 104.860 125.975 105.055 126.305 ;
        RECT 105.225 126.935 106.350 127.105 ;
        RECT 104.465 125.805 104.635 125.975 ;
        RECT 105.225 125.805 105.395 126.935 ;
        RECT 102.225 125.065 102.395 125.675 ;
        RECT 102.565 125.285 102.895 125.720 ;
        RECT 103.575 125.065 103.865 125.790 ;
        RECT 104.040 125.235 104.295 125.805 ;
        RECT 104.465 125.635 105.395 125.805 ;
        RECT 105.565 126.595 106.575 126.765 ;
        RECT 105.565 125.795 105.735 126.595 ;
        RECT 105.940 125.915 106.215 126.395 ;
        RECT 105.935 125.745 106.215 125.915 ;
        RECT 105.220 125.600 105.395 125.635 ;
        RECT 104.465 125.065 104.795 125.465 ;
        RECT 105.220 125.235 105.750 125.600 ;
        RECT 105.940 125.235 106.215 125.745 ;
        RECT 106.385 125.235 106.575 126.595 ;
        RECT 106.745 126.610 106.915 127.275 ;
        RECT 107.085 126.855 107.255 127.615 ;
        RECT 107.490 126.855 108.005 127.265 ;
        RECT 106.745 126.420 107.495 126.610 ;
        RECT 107.665 126.045 108.005 126.855 ;
        RECT 106.775 125.875 108.005 126.045 ;
        RECT 108.175 126.475 108.560 127.445 ;
        RECT 108.730 127.155 109.055 127.615 ;
        RECT 109.575 126.985 109.855 127.445 ;
        RECT 108.730 126.765 109.855 126.985 ;
        RECT 106.755 125.065 107.265 125.600 ;
        RECT 107.485 125.270 107.730 125.875 ;
        RECT 108.175 125.805 108.455 126.475 ;
        RECT 108.730 126.305 109.180 126.765 ;
        RECT 110.045 126.595 110.445 127.445 ;
        RECT 110.845 127.155 111.115 127.615 ;
        RECT 111.285 126.985 111.570 127.445 ;
        RECT 108.625 125.975 109.180 126.305 ;
        RECT 109.350 126.035 110.445 126.595 ;
        RECT 108.730 125.865 109.180 125.975 ;
        RECT 108.175 125.235 108.560 125.805 ;
        RECT 108.730 125.695 109.855 125.865 ;
        RECT 108.730 125.065 109.055 125.525 ;
        RECT 109.575 125.235 109.855 125.695 ;
        RECT 110.045 125.235 110.445 126.035 ;
        RECT 110.615 126.765 111.570 126.985 ;
        RECT 112.405 126.945 112.575 127.445 ;
        RECT 112.745 127.115 113.075 127.615 ;
        RECT 112.405 126.775 113.070 126.945 ;
        RECT 110.615 125.865 110.825 126.765 ;
        RECT 110.995 126.035 111.685 126.595 ;
        RECT 112.320 125.955 112.670 126.605 ;
        RECT 110.615 125.695 111.570 125.865 ;
        RECT 112.840 125.785 113.070 126.775 ;
        RECT 110.845 125.065 111.115 125.525 ;
        RECT 111.285 125.235 111.570 125.695 ;
        RECT 112.405 125.615 113.070 125.785 ;
        RECT 112.405 125.325 112.575 125.615 ;
        RECT 112.745 125.065 113.075 125.445 ;
        RECT 113.245 125.325 113.430 127.445 ;
        RECT 113.670 127.155 113.935 127.615 ;
        RECT 114.105 127.020 114.355 127.445 ;
        RECT 114.565 127.170 115.670 127.340 ;
        RECT 114.050 126.890 114.355 127.020 ;
        RECT 113.600 125.695 113.880 126.645 ;
        RECT 114.050 125.785 114.220 126.890 ;
        RECT 114.390 126.105 114.630 126.700 ;
        RECT 114.800 126.635 115.330 127.000 ;
        RECT 114.800 125.935 114.970 126.635 ;
        RECT 115.500 126.555 115.670 127.170 ;
        RECT 115.840 126.815 116.010 127.615 ;
        RECT 116.180 127.115 116.430 127.445 ;
        RECT 116.655 127.145 117.540 127.315 ;
        RECT 115.500 126.465 116.010 126.555 ;
        RECT 114.050 125.655 114.275 125.785 ;
        RECT 114.445 125.715 114.970 125.935 ;
        RECT 115.140 126.295 116.010 126.465 ;
        RECT 113.685 125.065 113.935 125.525 ;
        RECT 114.105 125.515 114.275 125.655 ;
        RECT 115.140 125.515 115.310 126.295 ;
        RECT 115.840 126.225 116.010 126.295 ;
        RECT 115.520 126.045 115.720 126.075 ;
        RECT 116.180 126.045 116.350 127.115 ;
        RECT 116.520 126.225 116.710 126.945 ;
        RECT 115.520 125.745 116.350 126.045 ;
        RECT 116.880 126.015 117.200 126.975 ;
        RECT 114.105 125.345 114.440 125.515 ;
        RECT 114.635 125.345 115.310 125.515 ;
        RECT 115.630 125.065 116.000 125.565 ;
        RECT 116.180 125.515 116.350 125.745 ;
        RECT 116.735 125.685 117.200 126.015 ;
        RECT 117.370 126.305 117.540 127.145 ;
        RECT 117.720 127.115 118.035 127.615 ;
        RECT 118.265 126.885 118.605 127.445 ;
        RECT 117.710 126.510 118.605 126.885 ;
        RECT 118.775 126.605 118.945 127.615 ;
        RECT 118.415 126.305 118.605 126.510 ;
        RECT 119.115 126.555 119.445 127.400 ;
        RECT 119.675 127.180 125.020 127.615 ;
        RECT 119.115 126.475 119.505 126.555 ;
        RECT 119.290 126.425 119.505 126.475 ;
        RECT 117.370 125.975 118.245 126.305 ;
        RECT 118.415 125.975 119.165 126.305 ;
        RECT 117.370 125.515 117.540 125.975 ;
        RECT 118.415 125.805 118.615 125.975 ;
        RECT 119.335 125.845 119.505 126.425 ;
        RECT 119.280 125.805 119.505 125.845 ;
        RECT 116.180 125.345 116.585 125.515 ;
        RECT 116.755 125.345 117.540 125.515 ;
        RECT 117.815 125.065 118.025 125.595 ;
        RECT 118.285 125.280 118.615 125.805 ;
        RECT 119.125 125.720 119.505 125.805 ;
        RECT 118.785 125.065 118.955 125.675 ;
        RECT 119.125 125.285 119.455 125.720 ;
        RECT 121.260 125.610 121.600 126.440 ;
        RECT 123.080 125.930 123.430 127.180 ;
        RECT 125.195 126.525 128.705 127.615 ;
        RECT 125.195 125.835 126.845 126.355 ;
        RECT 127.015 126.005 128.705 126.525 ;
        RECT 129.335 126.450 129.625 127.615 ;
        RECT 129.795 126.765 130.055 127.445 ;
        RECT 130.225 126.835 130.475 127.615 ;
        RECT 130.725 127.065 130.975 127.445 ;
        RECT 131.145 127.235 131.500 127.615 ;
        RECT 132.505 127.225 132.840 127.445 ;
        RECT 132.105 127.065 132.335 127.105 ;
        RECT 130.725 126.865 132.335 127.065 ;
        RECT 130.725 126.855 131.560 126.865 ;
        RECT 132.150 126.775 132.335 126.865 ;
        RECT 119.675 125.065 125.020 125.610 ;
        RECT 125.195 125.065 128.705 125.835 ;
        RECT 129.335 125.065 129.625 125.790 ;
        RECT 129.795 125.565 129.965 126.765 ;
        RECT 131.665 126.665 131.995 126.695 ;
        RECT 130.195 126.605 131.995 126.665 ;
        RECT 132.585 126.605 132.840 127.225 ;
        RECT 130.135 126.495 132.840 126.605 ;
        RECT 134.025 126.685 134.195 127.445 ;
        RECT 134.410 126.855 134.740 127.615 ;
        RECT 134.025 126.515 134.740 126.685 ;
        RECT 134.910 126.540 135.165 127.445 ;
        RECT 130.135 126.460 130.335 126.495 ;
        RECT 130.135 125.885 130.305 126.460 ;
        RECT 131.665 126.435 132.840 126.495 ;
        RECT 130.535 126.020 130.945 126.325 ;
        RECT 131.115 126.055 131.445 126.265 ;
        RECT 130.135 125.765 130.405 125.885 ;
        RECT 130.135 125.720 130.980 125.765 ;
        RECT 130.225 125.595 130.980 125.720 ;
        RECT 131.235 125.655 131.445 126.055 ;
        RECT 131.690 126.055 132.165 126.265 ;
        RECT 132.355 126.055 132.845 126.255 ;
        RECT 131.690 125.655 131.910 126.055 ;
        RECT 133.935 125.965 134.290 126.335 ;
        RECT 134.570 126.305 134.740 126.515 ;
        RECT 134.570 125.975 134.825 126.305 ;
        RECT 129.795 125.235 130.055 125.565 ;
        RECT 130.810 125.445 130.980 125.595 ;
        RECT 130.225 125.065 130.555 125.425 ;
        RECT 130.810 125.235 132.110 125.445 ;
        RECT 132.385 125.065 132.840 125.830 ;
        RECT 134.570 125.785 134.740 125.975 ;
        RECT 134.995 125.810 135.165 126.540 ;
        RECT 135.340 126.465 135.600 127.615 ;
        RECT 135.865 126.685 136.035 127.445 ;
        RECT 136.250 126.855 136.580 127.615 ;
        RECT 135.865 126.515 136.580 126.685 ;
        RECT 136.750 126.540 137.005 127.445 ;
        RECT 135.775 125.965 136.130 126.335 ;
        RECT 136.410 126.305 136.580 126.515 ;
        RECT 136.410 125.975 136.665 126.305 ;
        RECT 134.025 125.615 134.740 125.785 ;
        RECT 134.025 125.235 134.195 125.615 ;
        RECT 134.410 125.065 134.740 125.445 ;
        RECT 134.910 125.235 135.165 125.810 ;
        RECT 135.340 125.065 135.600 125.905 ;
        RECT 136.410 125.785 136.580 125.975 ;
        RECT 136.835 125.810 137.005 126.540 ;
        RECT 137.180 126.465 137.440 127.615 ;
        RECT 137.615 126.525 138.825 127.615 ;
        RECT 137.615 125.985 138.135 126.525 ;
        RECT 135.865 125.615 136.580 125.785 ;
        RECT 135.865 125.235 136.035 125.615 ;
        RECT 136.250 125.065 136.580 125.445 ;
        RECT 136.750 125.235 137.005 125.810 ;
        RECT 137.180 125.065 137.440 125.905 ;
        RECT 138.305 125.815 138.825 126.355 ;
        RECT 137.615 125.065 138.825 125.815 ;
        RECT 13.330 124.895 138.910 125.065 ;
        RECT 13.415 124.145 14.625 124.895 ;
        RECT 14.795 124.350 20.140 124.895 ;
        RECT 13.415 123.605 13.935 124.145 ;
        RECT 14.105 123.435 14.625 123.975 ;
        RECT 16.380 123.520 16.720 124.350 ;
        RECT 20.315 124.125 22.905 124.895 ;
        RECT 23.535 124.245 23.795 124.725 ;
        RECT 23.965 124.355 24.215 124.895 ;
        RECT 13.415 122.345 14.625 123.435 ;
        RECT 18.200 122.780 18.550 124.030 ;
        RECT 20.315 123.605 21.525 124.125 ;
        RECT 21.695 123.435 22.905 123.955 ;
        RECT 14.795 122.345 20.140 122.780 ;
        RECT 20.315 122.345 22.905 123.435 ;
        RECT 23.535 123.215 23.705 124.245 ;
        RECT 24.385 124.215 24.605 124.675 ;
        RECT 24.355 124.190 24.605 124.215 ;
        RECT 23.875 123.595 24.105 123.990 ;
        RECT 24.275 123.765 24.605 124.190 ;
        RECT 24.775 124.515 25.665 124.685 ;
        RECT 24.775 123.790 24.945 124.515 ;
        RECT 25.115 123.960 25.665 124.345 ;
        RECT 25.835 124.125 27.505 124.895 ;
        RECT 28.145 124.245 28.475 124.720 ;
        RECT 28.645 124.415 28.815 124.895 ;
        RECT 28.985 124.245 29.315 124.720 ;
        RECT 29.485 124.415 29.655 124.895 ;
        RECT 29.825 124.245 30.155 124.720 ;
        RECT 30.325 124.415 30.495 124.895 ;
        RECT 30.665 124.245 30.995 124.720 ;
        RECT 31.165 124.415 31.335 124.895 ;
        RECT 31.505 124.245 31.835 124.720 ;
        RECT 32.005 124.415 32.175 124.895 ;
        RECT 32.345 124.720 32.595 124.725 ;
        RECT 32.345 124.245 32.675 124.720 ;
        RECT 32.845 124.415 33.015 124.895 ;
        RECT 33.265 124.720 33.435 124.725 ;
        RECT 33.185 124.245 33.515 124.720 ;
        RECT 33.685 124.415 33.855 124.895 ;
        RECT 34.105 124.720 34.275 124.725 ;
        RECT 34.025 124.245 34.355 124.720 ;
        RECT 34.525 124.415 34.695 124.895 ;
        RECT 34.865 124.245 35.195 124.720 ;
        RECT 35.365 124.415 35.535 124.895 ;
        RECT 35.705 124.245 36.035 124.720 ;
        RECT 36.205 124.415 36.375 124.895 ;
        RECT 36.545 124.245 36.875 124.720 ;
        RECT 37.045 124.415 37.215 124.895 ;
        RECT 37.385 124.245 37.715 124.720 ;
        RECT 37.885 124.415 38.055 124.895 ;
        RECT 38.225 124.245 38.555 124.720 ;
        RECT 38.725 124.415 38.895 124.895 ;
        RECT 24.775 123.720 25.665 123.790 ;
        RECT 24.770 123.695 25.665 123.720 ;
        RECT 24.760 123.680 25.665 123.695 ;
        RECT 24.755 123.665 25.665 123.680 ;
        RECT 24.745 123.660 25.665 123.665 ;
        RECT 24.740 123.650 25.665 123.660 ;
        RECT 24.735 123.640 25.665 123.650 ;
        RECT 24.725 123.635 25.665 123.640 ;
        RECT 24.715 123.625 25.665 123.635 ;
        RECT 24.705 123.620 25.665 123.625 ;
        RECT 24.705 123.615 25.040 123.620 ;
        RECT 24.690 123.610 25.040 123.615 ;
        RECT 24.675 123.600 25.040 123.610 ;
        RECT 24.650 123.595 25.040 123.600 ;
        RECT 23.875 123.590 25.040 123.595 ;
        RECT 23.875 123.555 25.010 123.590 ;
        RECT 23.875 123.530 24.975 123.555 ;
        RECT 23.875 123.500 24.945 123.530 ;
        RECT 23.875 123.470 24.925 123.500 ;
        RECT 23.875 123.440 24.905 123.470 ;
        RECT 23.875 123.430 24.835 123.440 ;
        RECT 23.875 123.420 24.810 123.430 ;
        RECT 23.875 123.405 24.790 123.420 ;
        RECT 23.875 123.390 24.770 123.405 ;
        RECT 23.980 123.380 24.765 123.390 ;
        RECT 23.980 123.345 24.750 123.380 ;
        RECT 23.535 122.515 23.810 123.215 ;
        RECT 23.980 123.095 24.735 123.345 ;
        RECT 24.905 123.025 25.235 123.270 ;
        RECT 25.405 123.170 25.665 123.620 ;
        RECT 25.835 123.605 26.585 124.125 ;
        RECT 28.145 124.075 29.655 124.245 ;
        RECT 29.825 124.075 32.175 124.245 ;
        RECT 32.345 124.075 39.005 124.245 ;
        RECT 39.175 124.170 39.465 124.895 ;
        RECT 39.635 124.350 44.980 124.895 ;
        RECT 45.155 124.350 50.500 124.895 ;
        RECT 26.755 123.435 27.505 123.955 ;
        RECT 29.485 123.905 29.655 124.075 ;
        RECT 32.000 123.905 32.175 124.075 ;
        RECT 28.140 123.705 29.315 123.905 ;
        RECT 29.485 123.705 31.795 123.905 ;
        RECT 32.000 123.705 38.560 123.905 ;
        RECT 29.485 123.535 29.655 123.705 ;
        RECT 32.000 123.535 32.175 123.705 ;
        RECT 38.730 123.535 39.005 124.075 ;
        RECT 25.050 123.000 25.235 123.025 ;
        RECT 25.050 122.900 25.665 123.000 ;
        RECT 23.980 122.345 24.235 122.890 ;
        RECT 24.405 122.515 24.885 122.855 ;
        RECT 25.060 122.345 25.665 122.900 ;
        RECT 25.835 122.345 27.505 123.435 ;
        RECT 28.145 123.365 29.655 123.535 ;
        RECT 29.825 123.365 32.175 123.535 ;
        RECT 32.345 123.365 39.005 123.535 ;
        RECT 41.220 123.520 41.560 124.350 ;
        RECT 28.145 122.515 28.475 123.365 ;
        RECT 28.645 122.345 28.815 123.195 ;
        RECT 28.985 122.515 29.315 123.365 ;
        RECT 29.485 122.345 29.655 123.195 ;
        RECT 29.825 122.515 30.155 123.365 ;
        RECT 30.325 122.345 30.495 123.145 ;
        RECT 30.665 122.515 30.995 123.365 ;
        RECT 31.165 122.345 31.335 123.145 ;
        RECT 31.505 122.515 31.835 123.365 ;
        RECT 32.005 122.345 32.175 123.145 ;
        RECT 32.345 122.515 32.675 123.365 ;
        RECT 32.845 122.345 33.015 123.145 ;
        RECT 33.185 122.515 33.515 123.365 ;
        RECT 33.685 122.345 33.855 123.145 ;
        RECT 34.025 122.515 34.355 123.365 ;
        RECT 34.525 122.345 34.695 123.145 ;
        RECT 34.865 122.515 35.195 123.365 ;
        RECT 35.365 122.345 35.535 123.145 ;
        RECT 35.705 122.515 36.035 123.365 ;
        RECT 36.205 122.345 36.375 123.145 ;
        RECT 36.545 122.515 36.875 123.365 ;
        RECT 37.045 122.345 37.215 123.145 ;
        RECT 37.385 122.515 37.715 123.365 ;
        RECT 37.885 122.345 38.055 123.145 ;
        RECT 38.225 122.515 38.555 123.365 ;
        RECT 38.725 122.345 38.895 123.145 ;
        RECT 39.175 122.345 39.465 123.510 ;
        RECT 43.040 122.780 43.390 124.030 ;
        RECT 46.740 123.520 47.080 124.350 ;
        RECT 50.675 124.125 53.265 124.895 ;
        RECT 54.010 124.265 54.295 124.725 ;
        RECT 54.465 124.435 54.735 124.895 ;
        RECT 48.560 122.780 48.910 124.030 ;
        RECT 50.675 123.605 51.885 124.125 ;
        RECT 54.010 124.095 54.965 124.265 ;
        RECT 52.055 123.435 53.265 123.955 ;
        RECT 39.635 122.345 44.980 122.780 ;
        RECT 45.155 122.345 50.500 122.780 ;
        RECT 50.675 122.345 53.265 123.435 ;
        RECT 53.895 123.365 54.585 123.925 ;
        RECT 54.755 123.195 54.965 124.095 ;
        RECT 54.010 122.975 54.965 123.195 ;
        RECT 55.135 123.925 55.535 124.725 ;
        RECT 55.725 124.265 56.005 124.725 ;
        RECT 56.525 124.435 56.850 124.895 ;
        RECT 55.725 124.095 56.850 124.265 ;
        RECT 57.020 124.155 57.405 124.725 ;
        RECT 57.665 124.345 57.835 124.635 ;
        RECT 58.005 124.515 58.335 124.895 ;
        RECT 57.665 124.175 58.330 124.345 ;
        RECT 56.400 123.985 56.850 124.095 ;
        RECT 55.135 123.365 56.230 123.925 ;
        RECT 56.400 123.655 56.955 123.985 ;
        RECT 54.010 122.515 54.295 122.975 ;
        RECT 54.465 122.345 54.735 122.805 ;
        RECT 55.135 122.515 55.535 123.365 ;
        RECT 56.400 123.195 56.850 123.655 ;
        RECT 57.125 123.485 57.405 124.155 ;
        RECT 55.725 122.975 56.850 123.195 ;
        RECT 55.725 122.515 56.005 122.975 ;
        RECT 56.525 122.345 56.850 122.805 ;
        RECT 57.020 122.515 57.405 123.485 ;
        RECT 57.580 123.355 57.930 124.005 ;
        RECT 58.100 123.185 58.330 124.175 ;
        RECT 57.665 123.015 58.330 123.185 ;
        RECT 57.665 122.515 57.835 123.015 ;
        RECT 58.005 122.345 58.335 122.845 ;
        RECT 58.505 122.515 58.690 124.635 ;
        RECT 58.945 124.435 59.195 124.895 ;
        RECT 59.365 124.445 59.700 124.615 ;
        RECT 59.895 124.445 60.570 124.615 ;
        RECT 59.365 124.305 59.535 124.445 ;
        RECT 58.860 123.315 59.140 124.265 ;
        RECT 59.310 124.175 59.535 124.305 ;
        RECT 59.310 123.070 59.480 124.175 ;
        RECT 59.705 124.025 60.230 124.245 ;
        RECT 59.650 123.260 59.890 123.855 ;
        RECT 60.060 123.325 60.230 124.025 ;
        RECT 60.400 123.665 60.570 124.445 ;
        RECT 60.890 124.395 61.260 124.895 ;
        RECT 61.440 124.445 61.845 124.615 ;
        RECT 62.015 124.445 62.800 124.615 ;
        RECT 61.440 124.215 61.610 124.445 ;
        RECT 60.780 123.915 61.610 124.215 ;
        RECT 61.995 123.945 62.460 124.275 ;
        RECT 60.780 123.885 60.980 123.915 ;
        RECT 61.100 123.665 61.270 123.735 ;
        RECT 60.400 123.495 61.270 123.665 ;
        RECT 60.760 123.405 61.270 123.495 ;
        RECT 59.310 122.940 59.615 123.070 ;
        RECT 60.060 122.960 60.590 123.325 ;
        RECT 58.930 122.345 59.195 122.805 ;
        RECT 59.365 122.515 59.615 122.940 ;
        RECT 60.760 122.790 60.930 123.405 ;
        RECT 59.825 122.620 60.930 122.790 ;
        RECT 61.100 122.345 61.270 123.145 ;
        RECT 61.440 122.845 61.610 123.915 ;
        RECT 61.780 123.015 61.970 123.735 ;
        RECT 62.140 122.985 62.460 123.945 ;
        RECT 62.630 123.985 62.800 124.445 ;
        RECT 63.075 124.365 63.285 124.895 ;
        RECT 63.545 124.155 63.875 124.680 ;
        RECT 64.045 124.285 64.215 124.895 ;
        RECT 64.385 124.240 64.715 124.675 ;
        RECT 64.385 124.155 64.765 124.240 ;
        RECT 64.935 124.170 65.225 124.895 ;
        RECT 65.485 124.345 65.655 124.635 ;
        RECT 65.825 124.515 66.155 124.895 ;
        RECT 65.485 124.175 66.150 124.345 ;
        RECT 63.675 123.985 63.875 124.155 ;
        RECT 64.540 124.115 64.765 124.155 ;
        RECT 62.630 123.655 63.505 123.985 ;
        RECT 63.675 123.655 64.425 123.985 ;
        RECT 61.440 122.515 61.690 122.845 ;
        RECT 62.630 122.815 62.800 123.655 ;
        RECT 63.675 123.450 63.865 123.655 ;
        RECT 64.595 123.535 64.765 124.115 ;
        RECT 64.550 123.485 64.765 123.535 ;
        RECT 62.970 123.075 63.865 123.450 ;
        RECT 64.375 123.405 64.765 123.485 ;
        RECT 61.915 122.645 62.800 122.815 ;
        RECT 62.980 122.345 63.295 122.845 ;
        RECT 63.525 122.515 63.865 123.075 ;
        RECT 64.035 122.345 64.205 123.355 ;
        RECT 64.375 122.560 64.705 123.405 ;
        RECT 64.935 122.345 65.225 123.510 ;
        RECT 65.400 123.355 65.750 124.005 ;
        RECT 65.920 123.185 66.150 124.175 ;
        RECT 65.485 123.015 66.150 123.185 ;
        RECT 65.485 122.515 65.655 123.015 ;
        RECT 65.825 122.345 66.155 122.845 ;
        RECT 66.325 122.515 66.510 124.635 ;
        RECT 66.765 124.435 67.015 124.895 ;
        RECT 67.185 124.445 67.520 124.615 ;
        RECT 67.715 124.445 68.390 124.615 ;
        RECT 67.185 124.305 67.355 124.445 ;
        RECT 66.680 123.315 66.960 124.265 ;
        RECT 67.130 124.175 67.355 124.305 ;
        RECT 67.130 123.070 67.300 124.175 ;
        RECT 67.525 124.025 68.050 124.245 ;
        RECT 67.470 123.260 67.710 123.855 ;
        RECT 67.880 123.325 68.050 124.025 ;
        RECT 68.220 123.665 68.390 124.445 ;
        RECT 68.710 124.395 69.080 124.895 ;
        RECT 69.260 124.445 69.665 124.615 ;
        RECT 69.835 124.445 70.620 124.615 ;
        RECT 69.260 124.215 69.430 124.445 ;
        RECT 68.600 123.915 69.430 124.215 ;
        RECT 69.815 123.945 70.280 124.275 ;
        RECT 68.600 123.885 68.800 123.915 ;
        RECT 68.920 123.665 69.090 123.735 ;
        RECT 68.220 123.495 69.090 123.665 ;
        RECT 68.580 123.405 69.090 123.495 ;
        RECT 67.130 122.940 67.435 123.070 ;
        RECT 67.880 122.960 68.410 123.325 ;
        RECT 66.750 122.345 67.015 122.805 ;
        RECT 67.185 122.515 67.435 122.940 ;
        RECT 68.580 122.790 68.750 123.405 ;
        RECT 67.645 122.620 68.750 122.790 ;
        RECT 68.920 122.345 69.090 123.145 ;
        RECT 69.260 122.845 69.430 123.915 ;
        RECT 69.600 123.015 69.790 123.735 ;
        RECT 69.960 122.985 70.280 123.945 ;
        RECT 70.450 123.985 70.620 124.445 ;
        RECT 70.895 124.365 71.105 124.895 ;
        RECT 71.365 124.155 71.695 124.680 ;
        RECT 71.865 124.285 72.035 124.895 ;
        RECT 72.205 124.240 72.535 124.675 ;
        RECT 72.870 124.265 73.155 124.725 ;
        RECT 73.325 124.435 73.595 124.895 ;
        RECT 72.205 124.155 72.585 124.240 ;
        RECT 71.495 123.985 71.695 124.155 ;
        RECT 72.360 124.115 72.585 124.155 ;
        RECT 70.450 123.655 71.325 123.985 ;
        RECT 71.495 123.655 72.245 123.985 ;
        RECT 69.260 122.515 69.510 122.845 ;
        RECT 70.450 122.815 70.620 123.655 ;
        RECT 71.495 123.450 71.685 123.655 ;
        RECT 72.415 123.535 72.585 124.115 ;
        RECT 72.870 124.095 73.825 124.265 ;
        RECT 72.370 123.485 72.585 123.535 ;
        RECT 70.790 123.075 71.685 123.450 ;
        RECT 72.195 123.405 72.585 123.485 ;
        RECT 69.735 122.645 70.620 122.815 ;
        RECT 70.800 122.345 71.115 122.845 ;
        RECT 71.345 122.515 71.685 123.075 ;
        RECT 71.855 122.345 72.025 123.355 ;
        RECT 72.195 122.560 72.525 123.405 ;
        RECT 72.755 123.365 73.445 123.925 ;
        RECT 73.615 123.195 73.825 124.095 ;
        RECT 72.870 122.975 73.825 123.195 ;
        RECT 73.995 123.925 74.395 124.725 ;
        RECT 74.585 124.265 74.865 124.725 ;
        RECT 75.385 124.435 75.710 124.895 ;
        RECT 74.585 124.095 75.710 124.265 ;
        RECT 75.880 124.155 76.265 124.725 ;
        RECT 75.260 123.985 75.710 124.095 ;
        RECT 73.995 123.365 75.090 123.925 ;
        RECT 75.260 123.655 75.815 123.985 ;
        RECT 72.870 122.515 73.155 122.975 ;
        RECT 73.325 122.345 73.595 122.805 ;
        RECT 73.995 122.515 74.395 123.365 ;
        RECT 75.260 123.195 75.710 123.655 ;
        RECT 75.985 123.485 76.265 124.155 ;
        RECT 76.435 124.125 78.105 124.895 ;
        RECT 78.280 124.155 78.535 124.725 ;
        RECT 78.705 124.495 79.035 124.895 ;
        RECT 79.460 124.360 79.990 124.725 ;
        RECT 79.460 124.325 79.635 124.360 ;
        RECT 78.705 124.155 79.635 124.325 ;
        RECT 80.180 124.215 80.455 124.725 ;
        RECT 76.435 123.605 77.185 124.125 ;
        RECT 74.585 122.975 75.710 123.195 ;
        RECT 74.585 122.515 74.865 122.975 ;
        RECT 75.385 122.345 75.710 122.805 ;
        RECT 75.880 122.515 76.265 123.485 ;
        RECT 77.355 123.435 78.105 123.955 ;
        RECT 76.435 122.345 78.105 123.435 ;
        RECT 78.280 123.485 78.450 124.155 ;
        RECT 78.705 123.985 78.875 124.155 ;
        RECT 78.620 123.655 78.875 123.985 ;
        RECT 79.100 123.655 79.295 123.985 ;
        RECT 78.280 122.515 78.615 123.485 ;
        RECT 78.785 122.345 78.955 123.485 ;
        RECT 79.125 122.685 79.295 123.655 ;
        RECT 79.465 123.025 79.635 124.155 ;
        RECT 79.805 123.365 79.975 124.165 ;
        RECT 80.175 124.045 80.455 124.215 ;
        RECT 80.180 123.565 80.455 124.045 ;
        RECT 80.625 123.365 80.815 124.725 ;
        RECT 80.995 124.360 81.505 124.895 ;
        RECT 81.725 124.085 81.970 124.690 ;
        RECT 82.965 124.345 83.135 124.635 ;
        RECT 83.305 124.515 83.635 124.895 ;
        RECT 82.965 124.175 83.630 124.345 ;
        RECT 81.015 123.915 82.245 124.085 ;
        RECT 79.805 123.195 80.815 123.365 ;
        RECT 80.985 123.350 81.735 123.540 ;
        RECT 79.465 122.855 80.590 123.025 ;
        RECT 80.985 122.685 81.155 123.350 ;
        RECT 81.905 123.105 82.245 123.915 ;
        RECT 82.880 123.355 83.230 124.005 ;
        RECT 83.400 123.185 83.630 124.175 ;
        RECT 79.125 122.515 81.155 122.685 ;
        RECT 81.325 122.345 81.495 123.105 ;
        RECT 81.730 122.695 82.245 123.105 ;
        RECT 82.965 123.015 83.630 123.185 ;
        RECT 82.965 122.515 83.135 123.015 ;
        RECT 83.305 122.345 83.635 122.845 ;
        RECT 83.805 122.515 83.990 124.635 ;
        RECT 84.245 124.435 84.495 124.895 ;
        RECT 84.665 124.445 85.000 124.615 ;
        RECT 85.195 124.445 85.870 124.615 ;
        RECT 84.665 124.305 84.835 124.445 ;
        RECT 84.160 123.315 84.440 124.265 ;
        RECT 84.610 124.175 84.835 124.305 ;
        RECT 84.610 123.070 84.780 124.175 ;
        RECT 85.005 124.025 85.530 124.245 ;
        RECT 84.950 123.260 85.190 123.855 ;
        RECT 85.360 123.325 85.530 124.025 ;
        RECT 85.700 123.665 85.870 124.445 ;
        RECT 86.190 124.395 86.560 124.895 ;
        RECT 86.740 124.445 87.145 124.615 ;
        RECT 87.315 124.445 88.100 124.615 ;
        RECT 86.740 124.215 86.910 124.445 ;
        RECT 86.080 123.915 86.910 124.215 ;
        RECT 87.295 123.945 87.760 124.275 ;
        RECT 86.080 123.885 86.280 123.915 ;
        RECT 86.400 123.665 86.570 123.735 ;
        RECT 85.700 123.495 86.570 123.665 ;
        RECT 86.060 123.405 86.570 123.495 ;
        RECT 84.610 122.940 84.915 123.070 ;
        RECT 85.360 122.960 85.890 123.325 ;
        RECT 84.230 122.345 84.495 122.805 ;
        RECT 84.665 122.515 84.915 122.940 ;
        RECT 86.060 122.790 86.230 123.405 ;
        RECT 85.125 122.620 86.230 122.790 ;
        RECT 86.400 122.345 86.570 123.145 ;
        RECT 86.740 122.845 86.910 123.915 ;
        RECT 87.080 123.015 87.270 123.735 ;
        RECT 87.440 122.985 87.760 123.945 ;
        RECT 87.930 123.985 88.100 124.445 ;
        RECT 88.375 124.365 88.585 124.895 ;
        RECT 88.845 124.155 89.175 124.680 ;
        RECT 89.345 124.285 89.515 124.895 ;
        RECT 89.685 124.240 90.015 124.675 ;
        RECT 90.185 124.380 90.355 124.895 ;
        RECT 89.685 124.155 90.065 124.240 ;
        RECT 90.695 124.170 90.985 124.895 ;
        RECT 88.975 123.985 89.175 124.155 ;
        RECT 89.840 124.115 90.065 124.155 ;
        RECT 87.930 123.655 88.805 123.985 ;
        RECT 88.975 123.655 89.725 123.985 ;
        RECT 86.740 122.515 86.990 122.845 ;
        RECT 87.930 122.815 88.100 123.655 ;
        RECT 88.975 123.450 89.165 123.655 ;
        RECT 89.895 123.535 90.065 124.115 ;
        RECT 89.850 123.485 90.065 123.535 ;
        RECT 91.160 124.155 91.415 124.725 ;
        RECT 91.585 124.495 91.915 124.895 ;
        RECT 92.340 124.360 92.870 124.725 ;
        RECT 92.340 124.325 92.515 124.360 ;
        RECT 91.585 124.155 92.515 124.325 ;
        RECT 88.270 123.075 89.165 123.450 ;
        RECT 89.675 123.405 90.065 123.485 ;
        RECT 87.215 122.645 88.100 122.815 ;
        RECT 88.280 122.345 88.595 122.845 ;
        RECT 88.825 122.515 89.165 123.075 ;
        RECT 89.335 122.345 89.505 123.355 ;
        RECT 89.675 122.560 90.005 123.405 ;
        RECT 90.175 122.345 90.345 123.260 ;
        RECT 90.695 122.345 90.985 123.510 ;
        RECT 91.160 123.485 91.330 124.155 ;
        RECT 91.585 123.985 91.755 124.155 ;
        RECT 91.500 123.655 91.755 123.985 ;
        RECT 91.980 123.655 92.175 123.985 ;
        RECT 91.160 122.515 91.495 123.485 ;
        RECT 91.665 122.345 91.835 123.485 ;
        RECT 92.005 122.685 92.175 123.655 ;
        RECT 92.345 123.025 92.515 124.155 ;
        RECT 92.685 123.365 92.855 124.165 ;
        RECT 93.060 123.875 93.335 124.725 ;
        RECT 93.055 123.705 93.335 123.875 ;
        RECT 93.060 123.565 93.335 123.705 ;
        RECT 93.505 123.365 93.695 124.725 ;
        RECT 93.875 124.360 94.385 124.895 ;
        RECT 94.605 124.085 94.850 124.690 ;
        RECT 95.845 124.345 96.015 124.635 ;
        RECT 96.185 124.515 96.515 124.895 ;
        RECT 95.845 124.175 96.510 124.345 ;
        RECT 93.895 123.915 95.125 124.085 ;
        RECT 92.685 123.195 93.695 123.365 ;
        RECT 93.865 123.350 94.615 123.540 ;
        RECT 92.345 122.855 93.470 123.025 ;
        RECT 93.865 122.685 94.035 123.350 ;
        RECT 94.785 123.105 95.125 123.915 ;
        RECT 95.760 123.355 96.110 124.005 ;
        RECT 96.280 123.185 96.510 124.175 ;
        RECT 92.005 122.515 94.035 122.685 ;
        RECT 94.205 122.345 94.375 123.105 ;
        RECT 94.610 122.695 95.125 123.105 ;
        RECT 95.845 123.015 96.510 123.185 ;
        RECT 95.845 122.515 96.015 123.015 ;
        RECT 96.185 122.345 96.515 122.845 ;
        RECT 96.685 122.515 96.870 124.635 ;
        RECT 97.125 124.435 97.375 124.895 ;
        RECT 97.545 124.445 97.880 124.615 ;
        RECT 98.075 124.445 98.750 124.615 ;
        RECT 97.545 124.305 97.715 124.445 ;
        RECT 97.040 123.315 97.320 124.265 ;
        RECT 97.490 124.175 97.715 124.305 ;
        RECT 97.490 123.070 97.660 124.175 ;
        RECT 97.885 124.025 98.410 124.245 ;
        RECT 97.830 123.260 98.070 123.855 ;
        RECT 98.240 123.325 98.410 124.025 ;
        RECT 98.580 123.665 98.750 124.445 ;
        RECT 99.070 124.395 99.440 124.895 ;
        RECT 99.620 124.445 100.025 124.615 ;
        RECT 100.195 124.445 100.980 124.615 ;
        RECT 99.620 124.215 99.790 124.445 ;
        RECT 98.960 123.915 99.790 124.215 ;
        RECT 100.175 123.945 100.640 124.275 ;
        RECT 98.960 123.885 99.160 123.915 ;
        RECT 99.280 123.665 99.450 123.735 ;
        RECT 98.580 123.495 99.450 123.665 ;
        RECT 98.940 123.405 99.450 123.495 ;
        RECT 97.490 122.940 97.795 123.070 ;
        RECT 98.240 122.960 98.770 123.325 ;
        RECT 97.110 122.345 97.375 122.805 ;
        RECT 97.545 122.515 97.795 122.940 ;
        RECT 98.940 122.790 99.110 123.405 ;
        RECT 98.005 122.620 99.110 122.790 ;
        RECT 99.280 122.345 99.450 123.145 ;
        RECT 99.620 122.845 99.790 123.915 ;
        RECT 99.960 123.015 100.150 123.735 ;
        RECT 100.320 122.985 100.640 123.945 ;
        RECT 100.810 123.985 100.980 124.445 ;
        RECT 101.255 124.365 101.465 124.895 ;
        RECT 101.725 124.155 102.055 124.680 ;
        RECT 102.225 124.285 102.395 124.895 ;
        RECT 102.565 124.240 102.895 124.675 ;
        RECT 103.165 124.425 103.455 124.895 ;
        RECT 103.625 124.255 103.955 124.725 ;
        RECT 104.125 124.425 104.835 124.895 ;
        RECT 105.005 124.255 105.335 124.725 ;
        RECT 105.505 124.425 105.675 124.895 ;
        RECT 105.845 124.255 106.175 124.725 ;
        RECT 102.565 124.155 102.945 124.240 ;
        RECT 101.855 123.985 102.055 124.155 ;
        RECT 102.720 124.115 102.945 124.155 ;
        RECT 100.810 123.655 101.685 123.985 ;
        RECT 101.855 123.655 102.605 123.985 ;
        RECT 99.620 122.515 99.870 122.845 ;
        RECT 100.810 122.815 100.980 123.655 ;
        RECT 101.855 123.450 102.045 123.655 ;
        RECT 102.775 123.535 102.945 124.115 ;
        RECT 102.730 123.485 102.945 123.535 ;
        RECT 101.150 123.075 102.045 123.450 ;
        RECT 102.555 123.405 102.945 123.485 ;
        RECT 103.115 124.075 106.175 124.255 ;
        RECT 106.345 124.075 106.620 124.895 ;
        RECT 106.795 124.350 112.140 124.895 ;
        RECT 103.115 123.525 103.575 124.075 ;
        RECT 103.745 123.695 104.335 123.905 ;
        RECT 104.525 123.695 105.575 123.905 ;
        RECT 105.745 123.695 106.575 123.905 ;
        RECT 100.095 122.645 100.980 122.815 ;
        RECT 101.160 122.345 101.475 122.845 ;
        RECT 101.705 122.515 102.045 123.075 ;
        RECT 102.215 122.345 102.385 123.355 ;
        RECT 102.555 122.560 102.885 123.405 ;
        RECT 103.115 123.355 103.875 123.525 ;
        RECT 104.070 123.355 104.335 123.695 ;
        RECT 104.625 123.355 106.560 123.525 ;
        RECT 108.380 123.520 108.720 124.350 ;
        RECT 112.315 124.125 115.825 124.895 ;
        RECT 116.455 124.170 116.745 124.895 ;
        RECT 117.465 124.345 117.635 124.725 ;
        RECT 117.850 124.515 118.180 124.895 ;
        RECT 117.465 124.175 118.180 124.345 ;
        RECT 103.245 122.685 103.495 123.185 ;
        RECT 103.665 122.855 103.875 123.355 ;
        RECT 104.085 122.685 104.295 123.185 ;
        RECT 104.625 122.855 104.875 123.355 ;
        RECT 105.045 122.685 105.295 123.185 ;
        RECT 103.245 122.515 105.295 122.685 ;
        RECT 105.465 122.515 105.715 123.355 ;
        RECT 105.885 122.345 106.135 123.185 ;
        RECT 106.305 122.515 106.560 123.355 ;
        RECT 110.200 122.780 110.550 124.030 ;
        RECT 112.315 123.605 113.965 124.125 ;
        RECT 114.135 123.435 115.825 123.955 ;
        RECT 117.375 123.625 117.730 123.995 ;
        RECT 118.010 123.985 118.180 124.175 ;
        RECT 118.350 124.150 118.605 124.725 ;
        RECT 118.010 123.655 118.265 123.985 ;
        RECT 106.795 122.345 112.140 122.780 ;
        RECT 112.315 122.345 115.825 123.435 ;
        RECT 116.455 122.345 116.745 123.510 ;
        RECT 118.010 123.445 118.180 123.655 ;
        RECT 117.465 123.275 118.180 123.445 ;
        RECT 118.435 123.420 118.605 124.150 ;
        RECT 118.780 124.055 119.040 124.895 ;
        RECT 119.215 124.125 122.725 124.895 ;
        RECT 119.215 123.605 120.865 124.125 ;
        RECT 123.560 124.115 124.060 124.725 ;
        RECT 117.465 122.515 117.635 123.275 ;
        RECT 117.850 122.345 118.180 123.105 ;
        RECT 118.350 122.515 118.605 123.420 ;
        RECT 118.780 122.345 119.040 123.495 ;
        RECT 121.035 123.435 122.725 123.955 ;
        RECT 123.355 123.655 123.705 123.905 ;
        RECT 123.890 123.485 124.060 124.115 ;
        RECT 124.690 124.245 125.020 124.725 ;
        RECT 125.190 124.435 125.415 124.895 ;
        RECT 125.585 124.245 125.915 124.725 ;
        RECT 124.690 124.075 125.915 124.245 ;
        RECT 126.105 124.095 126.355 124.895 ;
        RECT 126.525 124.095 126.865 124.725 ;
        RECT 127.125 124.345 127.295 124.635 ;
        RECT 127.465 124.515 127.795 124.895 ;
        RECT 127.125 124.175 127.790 124.345 ;
        RECT 126.635 124.045 126.865 124.095 ;
        RECT 124.230 123.705 124.560 123.905 ;
        RECT 124.730 123.705 125.060 123.905 ;
        RECT 125.230 123.705 125.650 123.905 ;
        RECT 125.825 123.735 126.520 123.905 ;
        RECT 125.825 123.485 125.995 123.735 ;
        RECT 126.690 123.485 126.865 124.045 ;
        RECT 119.215 122.345 122.725 123.435 ;
        RECT 123.560 123.315 125.995 123.485 ;
        RECT 123.560 122.515 123.890 123.315 ;
        RECT 124.060 122.345 124.390 123.145 ;
        RECT 124.690 122.515 125.020 123.315 ;
        RECT 125.665 122.345 125.915 123.145 ;
        RECT 126.185 122.345 126.355 123.485 ;
        RECT 126.525 122.515 126.865 123.485 ;
        RECT 127.040 123.355 127.390 124.005 ;
        RECT 127.560 123.185 127.790 124.175 ;
        RECT 127.125 123.015 127.790 123.185 ;
        RECT 127.125 122.515 127.295 123.015 ;
        RECT 127.465 122.345 127.795 122.845 ;
        RECT 127.965 122.515 128.150 124.635 ;
        RECT 128.405 124.435 128.655 124.895 ;
        RECT 128.825 124.445 129.160 124.615 ;
        RECT 129.355 124.445 130.030 124.615 ;
        RECT 128.825 124.305 128.995 124.445 ;
        RECT 128.320 123.315 128.600 124.265 ;
        RECT 128.770 124.175 128.995 124.305 ;
        RECT 128.770 123.070 128.940 124.175 ;
        RECT 129.165 124.025 129.690 124.245 ;
        RECT 129.110 123.260 129.350 123.855 ;
        RECT 129.520 123.325 129.690 124.025 ;
        RECT 129.860 123.665 130.030 124.445 ;
        RECT 130.350 124.395 130.720 124.895 ;
        RECT 130.900 124.445 131.305 124.615 ;
        RECT 131.475 124.445 132.260 124.615 ;
        RECT 130.900 124.215 131.070 124.445 ;
        RECT 130.240 123.915 131.070 124.215 ;
        RECT 131.455 123.945 131.920 124.275 ;
        RECT 130.240 123.885 130.440 123.915 ;
        RECT 130.560 123.665 130.730 123.735 ;
        RECT 129.860 123.495 130.730 123.665 ;
        RECT 130.220 123.405 130.730 123.495 ;
        RECT 128.770 122.940 129.075 123.070 ;
        RECT 129.520 122.960 130.050 123.325 ;
        RECT 128.390 122.345 128.655 122.805 ;
        RECT 128.825 122.515 129.075 122.940 ;
        RECT 130.220 122.790 130.390 123.405 ;
        RECT 129.285 122.620 130.390 122.790 ;
        RECT 130.560 122.345 130.730 123.145 ;
        RECT 130.900 122.845 131.070 123.915 ;
        RECT 131.240 123.015 131.430 123.735 ;
        RECT 131.600 122.985 131.920 123.945 ;
        RECT 132.090 123.985 132.260 124.445 ;
        RECT 132.535 124.365 132.745 124.895 ;
        RECT 133.005 124.155 133.335 124.680 ;
        RECT 133.505 124.285 133.675 124.895 ;
        RECT 133.845 124.240 134.175 124.675 ;
        RECT 133.845 124.155 134.225 124.240 ;
        RECT 133.135 123.985 133.335 124.155 ;
        RECT 134.000 124.115 134.225 124.155 ;
        RECT 132.090 123.655 132.965 123.985 ;
        RECT 133.135 123.655 133.885 123.985 ;
        RECT 130.900 122.515 131.150 122.845 ;
        RECT 132.090 122.815 132.260 123.655 ;
        RECT 133.135 123.450 133.325 123.655 ;
        RECT 134.055 123.535 134.225 124.115 ;
        RECT 134.395 124.125 136.985 124.895 ;
        RECT 137.615 124.145 138.825 124.895 ;
        RECT 134.395 123.605 135.605 124.125 ;
        RECT 134.010 123.485 134.225 123.535 ;
        RECT 132.430 123.075 133.325 123.450 ;
        RECT 133.835 123.405 134.225 123.485 ;
        RECT 135.775 123.435 136.985 123.955 ;
        RECT 131.375 122.645 132.260 122.815 ;
        RECT 132.440 122.345 132.755 122.845 ;
        RECT 132.985 122.515 133.325 123.075 ;
        RECT 133.495 122.345 133.665 123.355 ;
        RECT 133.835 122.560 134.165 123.405 ;
        RECT 134.395 122.345 136.985 123.435 ;
        RECT 137.615 123.435 138.135 123.975 ;
        RECT 138.305 123.605 138.825 124.145 ;
        RECT 137.615 122.345 138.825 123.435 ;
        RECT 13.330 122.175 138.910 122.345 ;
        RECT 13.415 121.085 14.625 122.175 ;
        RECT 14.795 121.085 16.005 122.175 ;
        RECT 16.235 121.115 16.565 121.960 ;
        RECT 16.735 121.165 16.905 122.175 ;
        RECT 17.075 121.445 17.415 122.005 ;
        RECT 17.645 121.675 17.960 122.175 ;
        RECT 18.140 121.705 19.025 121.875 ;
        RECT 13.415 120.375 13.935 120.915 ;
        RECT 14.105 120.545 14.625 121.085 ;
        RECT 14.795 120.375 15.315 120.915 ;
        RECT 15.485 120.545 16.005 121.085 ;
        RECT 16.175 121.035 16.565 121.115 ;
        RECT 17.075 121.070 17.970 121.445 ;
        RECT 16.175 120.985 16.390 121.035 ;
        RECT 16.175 120.405 16.345 120.985 ;
        RECT 17.075 120.865 17.265 121.070 ;
        RECT 18.140 120.865 18.310 121.705 ;
        RECT 19.250 121.675 19.500 122.005 ;
        RECT 16.515 120.535 17.265 120.865 ;
        RECT 17.435 120.535 18.310 120.865 ;
        RECT 13.415 119.625 14.625 120.375 ;
        RECT 14.795 119.625 16.005 120.375 ;
        RECT 16.175 120.365 16.400 120.405 ;
        RECT 17.065 120.365 17.265 120.535 ;
        RECT 16.175 120.280 16.555 120.365 ;
        RECT 16.225 119.845 16.555 120.280 ;
        RECT 16.725 119.625 16.895 120.235 ;
        RECT 17.065 119.840 17.395 120.365 ;
        RECT 17.655 119.625 17.865 120.155 ;
        RECT 18.140 120.075 18.310 120.535 ;
        RECT 18.480 120.575 18.800 121.535 ;
        RECT 18.970 120.785 19.160 121.505 ;
        RECT 19.330 120.605 19.500 121.675 ;
        RECT 19.670 121.375 19.840 122.175 ;
        RECT 20.010 121.730 21.115 121.900 ;
        RECT 20.010 121.115 20.180 121.730 ;
        RECT 21.325 121.580 21.575 122.005 ;
        RECT 21.745 121.715 22.010 122.175 ;
        RECT 20.350 121.195 20.880 121.560 ;
        RECT 21.325 121.450 21.630 121.580 ;
        RECT 19.670 121.025 20.180 121.115 ;
        RECT 19.670 120.855 20.540 121.025 ;
        RECT 19.670 120.785 19.840 120.855 ;
        RECT 19.960 120.605 20.160 120.635 ;
        RECT 18.480 120.245 18.945 120.575 ;
        RECT 19.330 120.305 20.160 120.605 ;
        RECT 19.330 120.075 19.500 120.305 ;
        RECT 18.140 119.905 18.925 120.075 ;
        RECT 19.095 119.905 19.500 120.075 ;
        RECT 19.680 119.625 20.050 120.125 ;
        RECT 20.370 120.075 20.540 120.855 ;
        RECT 20.710 120.495 20.880 121.195 ;
        RECT 21.050 120.665 21.290 121.260 ;
        RECT 20.710 120.275 21.235 120.495 ;
        RECT 21.460 120.345 21.630 121.450 ;
        RECT 21.405 120.215 21.630 120.345 ;
        RECT 21.800 120.255 22.080 121.205 ;
        RECT 21.405 120.075 21.575 120.215 ;
        RECT 20.370 119.905 21.045 120.075 ;
        RECT 21.240 119.905 21.575 120.075 ;
        RECT 21.745 119.625 21.995 120.085 ;
        RECT 22.250 119.885 22.435 122.005 ;
        RECT 22.605 121.675 22.935 122.175 ;
        RECT 23.105 121.505 23.275 122.005 ;
        RECT 22.610 121.335 23.275 121.505 ;
        RECT 22.610 120.345 22.840 121.335 ;
        RECT 23.555 121.285 23.815 121.995 ;
        RECT 23.985 121.465 24.315 122.175 ;
        RECT 24.485 121.285 24.715 121.995 ;
        RECT 23.010 120.515 23.360 121.165 ;
        RECT 23.555 121.045 24.715 121.285 ;
        RECT 24.895 121.265 25.165 121.995 ;
        RECT 25.345 121.445 25.685 122.175 ;
        RECT 24.895 121.045 25.665 121.265 ;
        RECT 23.545 120.535 23.845 120.865 ;
        RECT 24.025 120.555 24.550 120.865 ;
        RECT 24.730 120.555 25.195 120.865 ;
        RECT 22.610 120.175 23.275 120.345 ;
        RECT 22.605 119.625 22.935 120.005 ;
        RECT 23.105 119.885 23.275 120.175 ;
        RECT 23.555 119.625 23.845 120.355 ;
        RECT 24.025 119.915 24.255 120.555 ;
        RECT 25.375 120.375 25.665 121.045 ;
        RECT 24.435 120.175 25.665 120.375 ;
        RECT 24.435 119.805 24.745 120.175 ;
        RECT 24.925 119.625 25.595 119.995 ;
        RECT 25.855 119.805 26.115 121.995 ;
        RECT 26.295 121.010 26.585 122.175 ;
        RECT 26.755 121.085 27.965 122.175 ;
        RECT 26.755 120.375 27.275 120.915 ;
        RECT 27.445 120.545 27.965 121.085 ;
        RECT 28.145 121.065 28.440 122.175 ;
        RECT 28.620 120.865 28.870 122.000 ;
        RECT 29.040 121.065 29.300 122.175 ;
        RECT 29.470 121.275 29.730 122.000 ;
        RECT 29.900 121.445 30.160 122.175 ;
        RECT 30.330 121.275 30.590 122.000 ;
        RECT 30.760 121.445 31.020 122.175 ;
        RECT 31.190 121.275 31.450 122.000 ;
        RECT 31.620 121.445 31.880 122.175 ;
        RECT 32.050 121.275 32.310 122.000 ;
        RECT 32.480 121.445 32.775 122.175 ;
        RECT 33.195 121.745 33.535 122.005 ;
        RECT 29.470 121.035 32.780 121.275 ;
        RECT 26.295 119.625 26.585 120.350 ;
        RECT 26.755 119.625 27.965 120.375 ;
        RECT 28.135 120.255 28.450 120.865 ;
        RECT 28.620 120.615 31.640 120.865 ;
        RECT 28.195 119.625 28.440 120.085 ;
        RECT 28.620 119.805 28.870 120.615 ;
        RECT 31.810 120.445 32.780 121.035 ;
        RECT 29.470 120.275 32.780 120.445 ;
        RECT 33.195 120.345 33.455 121.745 ;
        RECT 33.705 121.375 34.035 122.175 ;
        RECT 34.500 121.205 34.750 122.005 ;
        RECT 34.935 121.455 35.265 122.175 ;
        RECT 35.485 121.205 35.735 122.005 ;
        RECT 35.905 121.795 36.240 122.175 ;
        RECT 33.645 121.035 35.835 121.205 ;
        RECT 33.645 120.865 33.960 121.035 ;
        RECT 33.630 120.615 33.960 120.865 ;
        RECT 29.040 119.625 29.300 120.150 ;
        RECT 29.470 119.820 29.730 120.275 ;
        RECT 29.900 119.625 30.160 120.105 ;
        RECT 30.330 119.820 30.590 120.275 ;
        RECT 30.760 119.625 31.020 120.105 ;
        RECT 31.190 119.820 31.450 120.275 ;
        RECT 31.620 119.625 31.880 120.105 ;
        RECT 32.050 119.820 32.310 120.275 ;
        RECT 32.480 119.625 32.780 120.105 ;
        RECT 33.195 119.835 33.535 120.345 ;
        RECT 33.705 119.625 33.975 120.425 ;
        RECT 34.155 119.895 34.435 120.865 ;
        RECT 34.615 119.895 34.915 120.865 ;
        RECT 35.095 119.900 35.445 120.865 ;
        RECT 35.665 120.125 35.835 121.035 ;
        RECT 36.005 120.305 36.245 121.615 ;
        RECT 36.505 121.555 36.675 121.985 ;
        RECT 36.845 121.725 37.175 122.175 ;
        RECT 36.505 121.325 37.180 121.555 ;
        RECT 36.475 120.305 36.775 121.155 ;
        RECT 36.945 120.675 37.180 121.325 ;
        RECT 37.350 121.015 37.635 121.960 ;
        RECT 37.815 121.705 38.500 122.175 ;
        RECT 37.810 121.185 38.505 121.495 ;
        RECT 38.680 121.120 38.985 121.905 ;
        RECT 37.350 120.865 38.210 121.015 ;
        RECT 37.350 120.845 38.635 120.865 ;
        RECT 36.945 120.345 37.480 120.675 ;
        RECT 37.650 120.485 38.635 120.845 ;
        RECT 36.945 120.195 37.165 120.345 ;
        RECT 35.665 119.795 36.160 120.125 ;
        RECT 36.420 119.625 36.755 120.130 ;
        RECT 36.925 119.820 37.165 120.195 ;
        RECT 37.650 120.150 37.820 120.485 ;
        RECT 38.810 120.315 38.985 121.120 ;
        RECT 37.445 119.955 37.820 120.150 ;
        RECT 37.445 119.810 37.615 119.955 ;
        RECT 38.180 119.625 38.575 120.120 ;
        RECT 38.745 119.795 38.985 120.315 ;
        RECT 39.175 120.570 39.455 122.005 ;
        RECT 39.625 121.400 40.335 122.175 ;
        RECT 40.505 121.230 40.835 122.005 ;
        RECT 39.685 121.015 40.835 121.230 ;
        RECT 39.175 119.795 39.515 120.570 ;
        RECT 39.685 120.445 39.970 121.015 ;
        RECT 40.155 120.615 40.625 120.845 ;
        RECT 41.030 120.815 41.245 121.930 ;
        RECT 41.425 121.455 41.755 122.175 ;
        RECT 42.430 121.375 42.680 122.175 ;
        RECT 42.850 121.545 43.180 122.005 ;
        RECT 43.350 121.715 43.565 122.175 ;
        RECT 44.235 121.740 49.580 122.175 ;
        RECT 42.850 121.375 44.020 121.545 ;
        RECT 41.940 121.205 42.220 121.365 ;
        RECT 41.535 120.815 41.765 121.155 ;
        RECT 41.940 121.035 43.275 121.205 ;
        RECT 43.105 120.865 43.275 121.035 ;
        RECT 40.795 120.635 41.245 120.815 ;
        RECT 40.795 120.615 41.125 120.635 ;
        RECT 41.435 120.615 41.765 120.815 ;
        RECT 41.940 120.615 42.290 120.855 ;
        RECT 42.460 120.615 42.935 120.855 ;
        RECT 43.105 120.615 43.480 120.865 ;
        RECT 43.105 120.445 43.275 120.615 ;
        RECT 39.685 120.255 40.395 120.445 ;
        RECT 40.095 120.115 40.395 120.255 ;
        RECT 40.585 120.255 41.765 120.445 ;
        RECT 40.585 120.175 40.915 120.255 ;
        RECT 40.095 120.105 40.410 120.115 ;
        RECT 40.095 120.095 40.420 120.105 ;
        RECT 40.095 120.090 40.430 120.095 ;
        RECT 39.685 119.625 39.855 120.085 ;
        RECT 40.095 120.080 40.435 120.090 ;
        RECT 40.095 120.075 40.440 120.080 ;
        RECT 40.095 120.065 40.445 120.075 ;
        RECT 40.095 120.060 40.450 120.065 ;
        RECT 40.095 119.795 40.455 120.060 ;
        RECT 41.085 119.625 41.255 120.085 ;
        RECT 41.425 119.795 41.765 120.255 ;
        RECT 41.940 120.275 43.275 120.445 ;
        RECT 41.940 120.065 42.210 120.275 ;
        RECT 43.650 120.085 44.020 121.375 ;
        RECT 45.820 120.170 46.160 121.000 ;
        RECT 47.640 120.490 47.990 121.740 ;
        RECT 49.755 121.085 51.425 122.175 ;
        RECT 49.755 120.395 50.505 120.915 ;
        RECT 50.675 120.565 51.425 121.085 ;
        RECT 52.055 121.010 52.345 122.175 ;
        RECT 52.525 121.565 52.855 121.995 ;
        RECT 53.035 121.735 53.230 122.175 ;
        RECT 53.400 121.565 53.730 121.995 ;
        RECT 52.525 121.395 53.730 121.565 ;
        RECT 52.525 121.065 53.420 121.395 ;
        RECT 53.900 121.225 54.175 121.995 ;
        RECT 54.445 121.505 54.615 122.005 ;
        RECT 54.785 121.675 55.115 122.175 ;
        RECT 54.445 121.335 55.110 121.505 ;
        RECT 53.590 121.035 54.175 121.225 ;
        RECT 52.530 120.535 52.825 120.865 ;
        RECT 53.005 120.535 53.420 120.865 ;
        RECT 42.430 119.625 42.760 120.085 ;
        RECT 43.270 119.795 44.020 120.085 ;
        RECT 44.235 119.625 49.580 120.170 ;
        RECT 49.755 119.625 51.425 120.395 ;
        RECT 52.055 119.625 52.345 120.350 ;
        RECT 52.525 119.625 52.825 120.355 ;
        RECT 53.005 119.915 53.235 120.535 ;
        RECT 53.590 120.365 53.765 121.035 ;
        RECT 53.435 120.185 53.765 120.365 ;
        RECT 53.935 120.215 54.175 120.865 ;
        RECT 54.360 120.515 54.710 121.165 ;
        RECT 54.880 120.345 55.110 121.335 ;
        RECT 53.435 119.805 53.660 120.185 ;
        RECT 54.445 120.175 55.110 120.345 ;
        RECT 53.830 119.625 54.160 120.015 ;
        RECT 54.445 119.885 54.615 120.175 ;
        RECT 54.785 119.625 55.115 120.005 ;
        RECT 55.285 119.885 55.470 122.005 ;
        RECT 55.710 121.715 55.975 122.175 ;
        RECT 56.145 121.580 56.395 122.005 ;
        RECT 56.605 121.730 57.710 121.900 ;
        RECT 56.090 121.450 56.395 121.580 ;
        RECT 55.640 120.255 55.920 121.205 ;
        RECT 56.090 120.345 56.260 121.450 ;
        RECT 56.430 120.665 56.670 121.260 ;
        RECT 56.840 121.195 57.370 121.560 ;
        RECT 56.840 120.495 57.010 121.195 ;
        RECT 57.540 121.115 57.710 121.730 ;
        RECT 57.880 121.375 58.050 122.175 ;
        RECT 58.220 121.675 58.470 122.005 ;
        RECT 58.695 121.705 59.580 121.875 ;
        RECT 57.540 121.025 58.050 121.115 ;
        RECT 56.090 120.215 56.315 120.345 ;
        RECT 56.485 120.275 57.010 120.495 ;
        RECT 57.180 120.855 58.050 121.025 ;
        RECT 55.725 119.625 55.975 120.085 ;
        RECT 56.145 120.075 56.315 120.215 ;
        RECT 57.180 120.075 57.350 120.855 ;
        RECT 57.880 120.785 58.050 120.855 ;
        RECT 57.560 120.605 57.760 120.635 ;
        RECT 58.220 120.605 58.390 121.675 ;
        RECT 58.560 120.785 58.750 121.505 ;
        RECT 57.560 120.305 58.390 120.605 ;
        RECT 58.920 120.575 59.240 121.535 ;
        RECT 56.145 119.905 56.480 120.075 ;
        RECT 56.675 119.905 57.350 120.075 ;
        RECT 57.670 119.625 58.040 120.125 ;
        RECT 58.220 120.075 58.390 120.305 ;
        RECT 58.775 120.245 59.240 120.575 ;
        RECT 59.410 120.865 59.580 121.705 ;
        RECT 59.760 121.675 60.075 122.175 ;
        RECT 60.305 121.445 60.645 122.005 ;
        RECT 59.750 121.070 60.645 121.445 ;
        RECT 60.815 121.165 60.985 122.175 ;
        RECT 60.455 120.865 60.645 121.070 ;
        RECT 61.155 121.115 61.485 121.960 ;
        RECT 61.155 121.035 61.545 121.115 ;
        RECT 61.725 121.065 62.020 122.175 ;
        RECT 61.330 120.985 61.545 121.035 ;
        RECT 59.410 120.535 60.285 120.865 ;
        RECT 60.455 120.535 61.205 120.865 ;
        RECT 59.410 120.075 59.580 120.535 ;
        RECT 60.455 120.365 60.655 120.535 ;
        RECT 61.375 120.405 61.545 120.985 ;
        RECT 62.200 120.865 62.450 122.000 ;
        RECT 62.620 121.065 62.880 122.175 ;
        RECT 63.050 121.275 63.310 122.000 ;
        RECT 63.480 121.445 63.740 122.175 ;
        RECT 63.910 121.275 64.170 122.000 ;
        RECT 64.340 121.445 64.600 122.175 ;
        RECT 64.770 121.275 65.030 122.000 ;
        RECT 65.200 121.445 65.460 122.175 ;
        RECT 65.630 121.275 65.890 122.000 ;
        RECT 66.060 121.445 66.355 122.175 ;
        RECT 66.860 121.555 67.035 122.005 ;
        RECT 67.205 121.735 67.535 122.175 ;
        RECT 67.840 121.585 68.010 122.005 ;
        RECT 68.245 121.765 68.915 122.175 ;
        RECT 69.130 121.585 69.300 122.005 ;
        RECT 69.500 121.765 69.830 122.175 ;
        RECT 66.860 121.385 67.490 121.555 ;
        RECT 63.050 121.035 66.360 121.275 ;
        RECT 61.320 120.365 61.545 120.405 ;
        RECT 58.220 119.905 58.625 120.075 ;
        RECT 58.795 119.905 59.580 120.075 ;
        RECT 59.855 119.625 60.065 120.155 ;
        RECT 60.325 119.840 60.655 120.365 ;
        RECT 61.165 120.280 61.545 120.365 ;
        RECT 60.825 119.625 60.995 120.235 ;
        RECT 61.165 119.845 61.495 120.280 ;
        RECT 61.715 120.255 62.030 120.865 ;
        RECT 62.200 120.615 65.220 120.865 ;
        RECT 61.775 119.625 62.020 120.085 ;
        RECT 62.200 119.805 62.450 120.615 ;
        RECT 65.390 120.445 66.360 121.035 ;
        RECT 66.775 120.535 67.140 121.215 ;
        RECT 67.320 120.865 67.490 121.385 ;
        RECT 67.840 121.415 69.855 121.585 ;
        RECT 67.320 120.535 67.670 120.865 ;
        RECT 63.050 120.275 66.360 120.445 ;
        RECT 67.320 120.365 67.490 120.535 ;
        RECT 62.620 119.625 62.880 120.150 ;
        RECT 63.050 119.820 63.310 120.275 ;
        RECT 63.480 119.625 63.740 120.105 ;
        RECT 63.910 119.820 64.170 120.275 ;
        RECT 64.340 119.625 64.600 120.105 ;
        RECT 64.770 119.820 65.030 120.275 ;
        RECT 65.200 119.625 65.460 120.105 ;
        RECT 65.630 119.820 65.890 120.275 ;
        RECT 66.860 120.195 67.490 120.365 ;
        RECT 66.060 119.625 66.360 120.105 ;
        RECT 66.860 119.795 67.035 120.195 ;
        RECT 67.840 120.125 68.010 121.415 ;
        RECT 67.205 119.625 67.535 120.005 ;
        RECT 67.780 119.795 68.010 120.125 ;
        RECT 68.210 119.960 68.490 121.235 ;
        RECT 68.715 121.155 68.985 121.235 ;
        RECT 68.675 120.985 68.985 121.155 ;
        RECT 68.715 119.960 68.985 120.985 ;
        RECT 69.175 120.205 69.515 121.235 ;
        RECT 69.685 120.865 69.855 121.415 ;
        RECT 70.025 121.035 70.285 122.005 ;
        RECT 69.685 120.535 69.945 120.865 ;
        RECT 70.115 120.345 70.285 121.035 ;
        RECT 69.445 119.625 69.775 120.005 ;
        RECT 69.945 119.880 70.285 120.345 ;
        RECT 70.455 121.035 70.840 122.005 ;
        RECT 71.010 121.715 71.335 122.175 ;
        RECT 71.855 121.545 72.135 122.005 ;
        RECT 71.010 121.325 72.135 121.545 ;
        RECT 70.455 120.365 70.735 121.035 ;
        RECT 71.010 120.865 71.460 121.325 ;
        RECT 72.325 121.155 72.725 122.005 ;
        RECT 73.125 121.715 73.395 122.175 ;
        RECT 73.565 121.545 73.850 122.005 ;
        RECT 74.135 121.665 75.330 121.955 ;
        RECT 70.905 120.535 71.460 120.865 ;
        RECT 71.630 120.595 72.725 121.155 ;
        RECT 71.010 120.425 71.460 120.535 ;
        RECT 69.945 119.835 70.280 119.880 ;
        RECT 70.455 119.795 70.840 120.365 ;
        RECT 71.010 120.255 72.135 120.425 ;
        RECT 71.010 119.625 71.335 120.085 ;
        RECT 71.855 119.795 72.135 120.255 ;
        RECT 72.325 119.795 72.725 120.595 ;
        RECT 72.895 121.325 73.850 121.545 ;
        RECT 74.155 121.325 75.320 121.495 ;
        RECT 75.500 121.375 75.780 122.175 ;
        RECT 72.895 120.425 73.105 121.325 ;
        RECT 73.275 120.595 73.965 121.155 ;
        RECT 74.155 121.035 74.485 121.325 ;
        RECT 75.150 121.205 75.320 121.325 ;
        RECT 74.655 120.865 74.880 121.155 ;
        RECT 75.150 121.035 75.820 121.205 ;
        RECT 75.990 121.035 76.265 122.005 ;
        RECT 75.650 120.865 75.820 121.035 ;
        RECT 74.135 120.535 74.485 120.865 ;
        RECT 74.655 120.535 75.480 120.865 ;
        RECT 75.650 120.535 75.925 120.865 ;
        RECT 72.895 120.255 73.850 120.425 ;
        RECT 75.650 120.365 75.820 120.535 ;
        RECT 73.125 119.625 73.395 120.085 ;
        RECT 73.565 119.795 73.850 120.255 ;
        RECT 74.155 120.195 75.820 120.365 ;
        RECT 76.095 120.300 76.265 121.035 ;
        RECT 76.435 120.970 76.725 122.175 ;
        RECT 77.815 121.010 78.105 122.175 ;
        RECT 78.275 121.035 78.535 122.175 ;
        RECT 78.705 121.025 79.035 122.005 ;
        RECT 79.205 121.035 79.485 122.175 ;
        RECT 79.655 121.085 83.165 122.175 ;
        RECT 83.885 121.505 84.055 122.005 ;
        RECT 84.225 121.675 84.555 122.175 ;
        RECT 83.885 121.335 84.550 121.505 ;
        RECT 78.295 120.615 78.630 120.865 ;
        RECT 78.800 120.475 78.970 121.025 ;
        RECT 79.140 120.595 79.475 120.865 ;
        RECT 74.155 119.845 74.410 120.195 ;
        RECT 74.580 119.625 74.910 120.025 ;
        RECT 75.080 119.845 75.250 120.195 ;
        RECT 75.420 119.625 75.800 120.025 ;
        RECT 75.990 119.955 76.265 120.300 ;
        RECT 76.435 119.625 76.725 120.455 ;
        RECT 78.795 120.425 78.970 120.475 ;
        RECT 77.815 119.625 78.105 120.350 ;
        RECT 78.275 119.795 78.970 120.425 ;
        RECT 79.175 119.625 79.485 120.425 ;
        RECT 79.655 120.395 81.305 120.915 ;
        RECT 81.475 120.565 83.165 121.085 ;
        RECT 83.800 120.515 84.150 121.165 ;
        RECT 79.655 119.625 83.165 120.395 ;
        RECT 84.320 120.345 84.550 121.335 ;
        RECT 83.885 120.175 84.550 120.345 ;
        RECT 83.885 119.885 84.055 120.175 ;
        RECT 84.225 119.625 84.555 120.005 ;
        RECT 84.725 119.885 84.910 122.005 ;
        RECT 85.150 121.715 85.415 122.175 ;
        RECT 85.585 121.580 85.835 122.005 ;
        RECT 86.045 121.730 87.150 121.900 ;
        RECT 85.530 121.450 85.835 121.580 ;
        RECT 85.080 120.255 85.360 121.205 ;
        RECT 85.530 120.345 85.700 121.450 ;
        RECT 85.870 120.665 86.110 121.260 ;
        RECT 86.280 121.195 86.810 121.560 ;
        RECT 86.280 120.495 86.450 121.195 ;
        RECT 86.980 121.115 87.150 121.730 ;
        RECT 87.320 121.375 87.490 122.175 ;
        RECT 87.660 121.675 87.910 122.005 ;
        RECT 88.135 121.705 89.020 121.875 ;
        RECT 86.980 121.025 87.490 121.115 ;
        RECT 85.530 120.215 85.755 120.345 ;
        RECT 85.925 120.275 86.450 120.495 ;
        RECT 86.620 120.855 87.490 121.025 ;
        RECT 85.165 119.625 85.415 120.085 ;
        RECT 85.585 120.075 85.755 120.215 ;
        RECT 86.620 120.075 86.790 120.855 ;
        RECT 87.320 120.785 87.490 120.855 ;
        RECT 87.000 120.605 87.200 120.635 ;
        RECT 87.660 120.605 87.830 121.675 ;
        RECT 88.000 120.785 88.190 121.505 ;
        RECT 87.000 120.305 87.830 120.605 ;
        RECT 88.360 120.575 88.680 121.535 ;
        RECT 85.585 119.905 85.920 120.075 ;
        RECT 86.115 119.905 86.790 120.075 ;
        RECT 87.110 119.625 87.480 120.125 ;
        RECT 87.660 120.075 87.830 120.305 ;
        RECT 88.215 120.245 88.680 120.575 ;
        RECT 88.850 120.865 89.020 121.705 ;
        RECT 89.200 121.675 89.515 122.175 ;
        RECT 89.745 121.445 90.085 122.005 ;
        RECT 89.190 121.070 90.085 121.445 ;
        RECT 90.255 121.165 90.425 122.175 ;
        RECT 89.895 120.865 90.085 121.070 ;
        RECT 90.595 121.115 90.925 121.960 ;
        RECT 91.095 121.260 91.265 122.175 ;
        RECT 91.615 121.740 96.960 122.175 ;
        RECT 90.595 121.035 90.985 121.115 ;
        RECT 90.770 120.985 90.985 121.035 ;
        RECT 88.850 120.535 89.725 120.865 ;
        RECT 89.895 120.535 90.645 120.865 ;
        RECT 88.850 120.075 89.020 120.535 ;
        RECT 89.895 120.365 90.095 120.535 ;
        RECT 90.815 120.405 90.985 120.985 ;
        RECT 90.760 120.365 90.985 120.405 ;
        RECT 87.660 119.905 88.065 120.075 ;
        RECT 88.235 119.905 89.020 120.075 ;
        RECT 89.295 119.625 89.505 120.155 ;
        RECT 89.765 119.840 90.095 120.365 ;
        RECT 90.605 120.280 90.985 120.365 ;
        RECT 90.265 119.625 90.435 120.235 ;
        RECT 90.605 119.845 90.935 120.280 ;
        RECT 93.200 120.170 93.540 121.000 ;
        RECT 95.020 120.490 95.370 121.740 ;
        RECT 97.135 121.085 100.645 122.175 ;
        RECT 97.135 120.395 98.785 120.915 ;
        RECT 98.955 120.565 100.645 121.085 ;
        RECT 101.795 121.035 102.005 122.175 ;
        RECT 102.175 121.025 102.505 122.005 ;
        RECT 102.675 121.035 102.905 122.175 ;
        RECT 91.105 119.625 91.275 120.140 ;
        RECT 91.615 119.625 96.960 120.170 ;
        RECT 97.135 119.625 100.645 120.395 ;
        RECT 101.795 119.625 102.005 120.445 ;
        RECT 102.175 120.425 102.425 121.025 ;
        RECT 103.575 121.010 103.865 122.175 ;
        RECT 104.035 121.670 104.665 122.175 ;
        RECT 104.050 121.135 104.305 121.500 ;
        RECT 104.475 121.495 104.665 121.670 ;
        RECT 104.845 121.665 105.320 122.005 ;
        RECT 104.475 121.305 104.805 121.495 ;
        RECT 105.030 121.135 105.280 121.430 ;
        RECT 105.505 121.330 105.720 122.175 ;
        RECT 105.920 121.335 106.195 122.005 ;
        RECT 104.050 120.965 105.840 121.135 ;
        RECT 106.025 120.985 106.195 121.335 ;
        RECT 106.365 121.165 106.625 122.175 ;
        RECT 106.795 121.085 109.385 122.175 ;
        RECT 102.595 120.615 102.925 120.865 ;
        RECT 102.175 119.795 102.505 120.425 ;
        RECT 102.675 119.625 102.905 120.445 ;
        RECT 103.575 119.625 103.865 120.350 ;
        RECT 104.035 120.305 104.420 120.785 ;
        RECT 104.590 120.110 104.845 120.965 ;
        RECT 104.055 119.845 104.845 120.110 ;
        RECT 105.015 120.290 105.425 120.785 ;
        RECT 105.610 120.535 105.840 120.965 ;
        RECT 106.010 120.465 106.625 120.985 ;
        RECT 105.015 119.845 105.245 120.290 ;
        RECT 106.010 120.255 106.180 120.465 ;
        RECT 106.795 120.395 108.005 120.915 ;
        RECT 108.175 120.565 109.385 121.085 ;
        RECT 109.555 121.035 109.895 122.005 ;
        RECT 110.065 121.035 110.235 122.175 ;
        RECT 110.505 121.375 110.755 122.175 ;
        RECT 111.400 121.205 111.730 122.005 ;
        RECT 112.030 121.375 112.360 122.175 ;
        RECT 112.530 121.205 112.860 122.005 ;
        RECT 113.325 121.505 113.495 122.005 ;
        RECT 113.665 121.675 113.995 122.175 ;
        RECT 113.325 121.335 113.990 121.505 ;
        RECT 110.425 121.035 112.860 121.205 ;
        RECT 109.555 120.475 109.730 121.035 ;
        RECT 110.425 120.785 110.595 121.035 ;
        RECT 109.900 120.615 110.595 120.785 ;
        RECT 110.770 120.615 111.190 120.815 ;
        RECT 111.360 120.615 111.690 120.815 ;
        RECT 111.860 120.615 112.190 120.815 ;
        RECT 109.555 120.425 109.785 120.475 ;
        RECT 105.425 119.625 105.755 120.120 ;
        RECT 105.930 119.795 106.180 120.255 ;
        RECT 106.350 119.625 106.625 120.285 ;
        RECT 106.795 119.625 109.385 120.395 ;
        RECT 109.555 119.795 109.895 120.425 ;
        RECT 110.065 119.625 110.315 120.425 ;
        RECT 110.505 120.275 111.730 120.445 ;
        RECT 110.505 119.795 110.835 120.275 ;
        RECT 111.005 119.625 111.230 120.085 ;
        RECT 111.400 119.795 111.730 120.275 ;
        RECT 112.360 120.405 112.530 121.035 ;
        RECT 112.715 120.615 113.065 120.865 ;
        RECT 113.240 120.515 113.590 121.165 ;
        RECT 112.360 119.795 112.860 120.405 ;
        RECT 113.760 120.345 113.990 121.335 ;
        RECT 113.325 120.175 113.990 120.345 ;
        RECT 113.325 119.885 113.495 120.175 ;
        RECT 113.665 119.625 113.995 120.005 ;
        RECT 114.165 119.885 114.350 122.005 ;
        RECT 114.590 121.715 114.855 122.175 ;
        RECT 115.025 121.580 115.275 122.005 ;
        RECT 115.485 121.730 116.590 121.900 ;
        RECT 114.970 121.450 115.275 121.580 ;
        RECT 114.520 120.255 114.800 121.205 ;
        RECT 114.970 120.345 115.140 121.450 ;
        RECT 115.310 120.665 115.550 121.260 ;
        RECT 115.720 121.195 116.250 121.560 ;
        RECT 115.720 120.495 115.890 121.195 ;
        RECT 116.420 121.115 116.590 121.730 ;
        RECT 116.760 121.375 116.930 122.175 ;
        RECT 117.100 121.675 117.350 122.005 ;
        RECT 117.575 121.705 118.460 121.875 ;
        RECT 116.420 121.025 116.930 121.115 ;
        RECT 114.970 120.215 115.195 120.345 ;
        RECT 115.365 120.275 115.890 120.495 ;
        RECT 116.060 120.855 116.930 121.025 ;
        RECT 114.605 119.625 114.855 120.085 ;
        RECT 115.025 120.075 115.195 120.215 ;
        RECT 116.060 120.075 116.230 120.855 ;
        RECT 116.760 120.785 116.930 120.855 ;
        RECT 116.440 120.605 116.640 120.635 ;
        RECT 117.100 120.605 117.270 121.675 ;
        RECT 117.440 120.785 117.630 121.505 ;
        RECT 116.440 120.305 117.270 120.605 ;
        RECT 117.800 120.575 118.120 121.535 ;
        RECT 115.025 119.905 115.360 120.075 ;
        RECT 115.555 119.905 116.230 120.075 ;
        RECT 116.550 119.625 116.920 120.125 ;
        RECT 117.100 120.075 117.270 120.305 ;
        RECT 117.655 120.245 118.120 120.575 ;
        RECT 118.290 120.865 118.460 121.705 ;
        RECT 118.640 121.675 118.955 122.175 ;
        RECT 119.185 121.445 119.525 122.005 ;
        RECT 118.630 121.070 119.525 121.445 ;
        RECT 119.695 121.165 119.865 122.175 ;
        RECT 119.335 120.865 119.525 121.070 ;
        RECT 120.035 121.115 120.365 121.960 ;
        RECT 120.630 121.385 121.165 122.005 ;
        RECT 120.035 121.035 120.425 121.115 ;
        RECT 120.210 120.985 120.425 121.035 ;
        RECT 118.290 120.535 119.165 120.865 ;
        RECT 119.335 120.535 120.085 120.865 ;
        RECT 118.290 120.075 118.460 120.535 ;
        RECT 119.335 120.365 119.535 120.535 ;
        RECT 120.255 120.405 120.425 120.985 ;
        RECT 120.200 120.365 120.425 120.405 ;
        RECT 117.100 119.905 117.505 120.075 ;
        RECT 117.675 119.905 118.460 120.075 ;
        RECT 118.735 119.625 118.945 120.155 ;
        RECT 119.205 119.840 119.535 120.365 ;
        RECT 120.045 120.280 120.425 120.365 ;
        RECT 120.630 120.365 120.945 121.385 ;
        RECT 121.335 121.375 121.665 122.175 ;
        RECT 122.895 121.740 128.240 122.175 ;
        RECT 122.150 121.205 122.540 121.380 ;
        RECT 121.115 121.035 122.540 121.205 ;
        RECT 121.115 120.535 121.285 121.035 ;
        RECT 119.705 119.625 119.875 120.235 ;
        RECT 120.045 119.845 120.375 120.280 ;
        RECT 120.630 119.795 121.245 120.365 ;
        RECT 121.535 120.305 121.800 120.865 ;
        RECT 121.970 120.135 122.140 121.035 ;
        RECT 122.310 120.305 122.665 120.865 ;
        RECT 124.480 120.170 124.820 121.000 ;
        RECT 126.300 120.490 126.650 121.740 ;
        RECT 129.335 121.010 129.625 122.175 ;
        RECT 129.980 121.205 130.370 121.380 ;
        RECT 130.855 121.375 131.185 122.175 ;
        RECT 131.355 121.385 131.890 122.005 ;
        RECT 129.980 121.035 131.405 121.205 ;
        RECT 121.415 119.625 121.630 120.135 ;
        RECT 121.860 119.805 122.140 120.135 ;
        RECT 122.320 119.625 122.560 120.135 ;
        RECT 122.895 119.625 128.240 120.170 ;
        RECT 129.335 119.625 129.625 120.350 ;
        RECT 129.855 120.305 130.210 120.865 ;
        RECT 130.380 120.135 130.550 121.035 ;
        RECT 130.720 120.305 130.985 120.865 ;
        RECT 131.235 120.535 131.405 121.035 ;
        RECT 131.575 120.365 131.890 121.385 ;
        RECT 129.960 119.625 130.200 120.135 ;
        RECT 130.380 119.805 130.660 120.135 ;
        RECT 130.890 119.625 131.105 120.135 ;
        RECT 131.275 119.795 131.890 120.365 ;
        RECT 132.130 121.385 132.665 122.005 ;
        RECT 132.130 120.365 132.445 121.385 ;
        RECT 132.835 121.375 133.165 122.175 ;
        RECT 133.650 121.205 134.040 121.380 ;
        RECT 132.615 121.035 134.040 121.205 ;
        RECT 134.395 121.085 135.605 122.175 ;
        RECT 132.615 120.535 132.785 121.035 ;
        RECT 132.130 119.795 132.745 120.365 ;
        RECT 133.035 120.305 133.300 120.865 ;
        RECT 133.470 120.135 133.640 121.035 ;
        RECT 133.810 120.305 134.165 120.865 ;
        RECT 134.395 120.375 134.915 120.915 ;
        RECT 135.085 120.545 135.605 121.085 ;
        RECT 135.865 121.245 136.035 122.005 ;
        RECT 136.250 121.415 136.580 122.175 ;
        RECT 135.865 121.075 136.580 121.245 ;
        RECT 136.750 121.100 137.005 122.005 ;
        RECT 135.775 120.525 136.130 120.895 ;
        RECT 136.410 120.865 136.580 121.075 ;
        RECT 136.410 120.535 136.665 120.865 ;
        RECT 132.915 119.625 133.130 120.135 ;
        RECT 133.360 119.805 133.640 120.135 ;
        RECT 133.820 119.625 134.060 120.135 ;
        RECT 134.395 119.625 135.605 120.375 ;
        RECT 136.410 120.345 136.580 120.535 ;
        RECT 136.835 120.370 137.005 121.100 ;
        RECT 137.180 121.025 137.440 122.175 ;
        RECT 137.615 121.085 138.825 122.175 ;
        RECT 137.615 120.545 138.135 121.085 ;
        RECT 135.865 120.175 136.580 120.345 ;
        RECT 135.865 119.795 136.035 120.175 ;
        RECT 136.250 119.625 136.580 120.005 ;
        RECT 136.750 119.795 137.005 120.370 ;
        RECT 137.180 119.625 137.440 120.465 ;
        RECT 138.305 120.375 138.825 120.915 ;
        RECT 137.615 119.625 138.825 120.375 ;
        RECT 13.330 119.455 138.910 119.625 ;
        RECT 13.415 118.705 14.625 119.455 ;
        RECT 13.415 118.165 13.935 118.705 ;
        RECT 14.795 118.685 16.465 119.455 ;
        RECT 16.670 118.715 17.285 119.285 ;
        RECT 17.455 118.945 17.670 119.455 ;
        RECT 17.900 118.945 18.180 119.275 ;
        RECT 18.360 118.945 18.600 119.455 ;
        RECT 14.105 117.995 14.625 118.535 ;
        RECT 14.795 118.165 15.545 118.685 ;
        RECT 15.715 117.995 16.465 118.515 ;
        RECT 13.415 116.905 14.625 117.995 ;
        RECT 14.795 116.905 16.465 117.995 ;
        RECT 16.670 117.695 16.985 118.715 ;
        RECT 17.155 118.045 17.325 118.545 ;
        RECT 17.575 118.215 17.840 118.775 ;
        RECT 18.010 118.045 18.180 118.945 ;
        RECT 18.350 118.215 18.705 118.775 ;
        RECT 18.935 118.635 19.195 119.455 ;
        RECT 19.365 118.635 19.695 119.055 ;
        RECT 19.875 118.970 20.665 119.235 ;
        RECT 19.445 118.545 19.695 118.635 ;
        RECT 17.155 117.875 18.580 118.045 ;
        RECT 16.670 117.075 17.205 117.695 ;
        RECT 17.375 116.905 17.705 117.705 ;
        RECT 18.190 117.700 18.580 117.875 ;
        RECT 18.935 117.585 19.275 118.465 ;
        RECT 19.445 118.295 20.240 118.545 ;
        RECT 18.935 116.905 19.195 117.415 ;
        RECT 19.445 117.075 19.615 118.295 ;
        RECT 20.410 118.115 20.665 118.970 ;
        RECT 20.835 118.815 21.035 119.235 ;
        RECT 21.225 118.995 21.555 119.455 ;
        RECT 20.835 118.295 21.245 118.815 ;
        RECT 21.725 118.805 21.985 119.285 ;
        RECT 21.415 118.115 21.645 118.545 ;
        RECT 19.855 117.945 21.645 118.115 ;
        RECT 19.855 117.580 20.105 117.945 ;
        RECT 20.275 117.585 20.605 117.775 ;
        RECT 20.825 117.650 21.540 117.945 ;
        RECT 21.815 117.775 21.985 118.805 ;
        RECT 22.245 118.905 22.415 119.195 ;
        RECT 22.585 119.075 22.915 119.455 ;
        RECT 22.245 118.735 22.910 118.905 ;
        RECT 22.160 117.915 22.510 118.565 ;
        RECT 20.275 117.410 20.470 117.585 ;
        RECT 19.855 116.905 20.470 117.410 ;
        RECT 20.640 117.075 21.115 117.415 ;
        RECT 21.285 116.905 21.500 117.450 ;
        RECT 21.710 117.075 21.985 117.775 ;
        RECT 22.680 117.745 22.910 118.735 ;
        RECT 22.245 117.575 22.910 117.745 ;
        RECT 22.245 117.075 22.415 117.575 ;
        RECT 22.585 116.905 22.915 117.405 ;
        RECT 23.085 117.075 23.270 119.195 ;
        RECT 23.525 118.995 23.775 119.455 ;
        RECT 23.945 119.005 24.280 119.175 ;
        RECT 24.475 119.005 25.150 119.175 ;
        RECT 23.945 118.865 24.115 119.005 ;
        RECT 23.440 117.875 23.720 118.825 ;
        RECT 23.890 118.735 24.115 118.865 ;
        RECT 23.890 117.630 24.060 118.735 ;
        RECT 24.285 118.585 24.810 118.805 ;
        RECT 24.230 117.820 24.470 118.415 ;
        RECT 24.640 117.885 24.810 118.585 ;
        RECT 24.980 118.225 25.150 119.005 ;
        RECT 25.470 118.955 25.840 119.455 ;
        RECT 26.020 119.005 26.425 119.175 ;
        RECT 26.595 119.005 27.380 119.175 ;
        RECT 26.020 118.775 26.190 119.005 ;
        RECT 25.360 118.475 26.190 118.775 ;
        RECT 26.575 118.505 27.040 118.835 ;
        RECT 25.360 118.445 25.560 118.475 ;
        RECT 25.680 118.225 25.850 118.295 ;
        RECT 24.980 118.055 25.850 118.225 ;
        RECT 25.340 117.965 25.850 118.055 ;
        RECT 23.890 117.500 24.195 117.630 ;
        RECT 24.640 117.520 25.170 117.885 ;
        RECT 23.510 116.905 23.775 117.365 ;
        RECT 23.945 117.075 24.195 117.500 ;
        RECT 25.340 117.350 25.510 117.965 ;
        RECT 24.405 117.180 25.510 117.350 ;
        RECT 25.680 116.905 25.850 117.705 ;
        RECT 26.020 117.405 26.190 118.475 ;
        RECT 26.360 117.575 26.550 118.295 ;
        RECT 26.720 117.545 27.040 118.505 ;
        RECT 27.210 118.545 27.380 119.005 ;
        RECT 27.655 118.925 27.865 119.455 ;
        RECT 28.125 118.715 28.455 119.240 ;
        RECT 28.625 118.845 28.795 119.455 ;
        RECT 28.965 118.800 29.295 119.235 ;
        RECT 29.680 118.945 29.920 119.455 ;
        RECT 30.100 118.945 30.380 119.275 ;
        RECT 30.610 118.945 30.825 119.455 ;
        RECT 28.965 118.715 29.345 118.800 ;
        RECT 28.255 118.545 28.455 118.715 ;
        RECT 29.120 118.675 29.345 118.715 ;
        RECT 27.210 118.215 28.085 118.545 ;
        RECT 28.255 118.215 29.005 118.545 ;
        RECT 26.020 117.075 26.270 117.405 ;
        RECT 27.210 117.375 27.380 118.215 ;
        RECT 28.255 118.010 28.445 118.215 ;
        RECT 29.175 118.095 29.345 118.675 ;
        RECT 29.575 118.215 29.930 118.775 ;
        RECT 29.130 118.045 29.345 118.095 ;
        RECT 30.100 118.045 30.270 118.945 ;
        RECT 30.440 118.215 30.705 118.775 ;
        RECT 30.995 118.715 31.610 119.285 ;
        RECT 31.905 118.905 32.075 119.195 ;
        RECT 32.245 119.075 32.575 119.455 ;
        RECT 31.905 118.735 32.570 118.905 ;
        RECT 30.955 118.045 31.125 118.545 ;
        RECT 27.550 117.635 28.445 118.010 ;
        RECT 28.955 117.965 29.345 118.045 ;
        RECT 26.495 117.205 27.380 117.375 ;
        RECT 27.560 116.905 27.875 117.405 ;
        RECT 28.105 117.075 28.445 117.635 ;
        RECT 28.615 116.905 28.785 117.915 ;
        RECT 28.955 117.120 29.285 117.965 ;
        RECT 29.700 117.875 31.125 118.045 ;
        RECT 29.700 117.700 30.090 117.875 ;
        RECT 30.575 116.905 30.905 117.705 ;
        RECT 31.295 117.695 31.610 118.715 ;
        RECT 31.820 117.915 32.170 118.565 ;
        RECT 32.340 117.745 32.570 118.735 ;
        RECT 31.075 117.075 31.610 117.695 ;
        RECT 31.905 117.575 32.570 117.745 ;
        RECT 31.905 117.075 32.075 117.575 ;
        RECT 32.245 116.905 32.575 117.405 ;
        RECT 32.745 117.075 32.930 119.195 ;
        RECT 33.185 118.995 33.435 119.455 ;
        RECT 33.605 119.005 33.940 119.175 ;
        RECT 34.135 119.005 34.810 119.175 ;
        RECT 33.605 118.865 33.775 119.005 ;
        RECT 33.100 117.875 33.380 118.825 ;
        RECT 33.550 118.735 33.775 118.865 ;
        RECT 33.550 117.630 33.720 118.735 ;
        RECT 33.945 118.585 34.470 118.805 ;
        RECT 33.890 117.820 34.130 118.415 ;
        RECT 34.300 117.885 34.470 118.585 ;
        RECT 34.640 118.225 34.810 119.005 ;
        RECT 35.130 118.955 35.500 119.455 ;
        RECT 35.680 119.005 36.085 119.175 ;
        RECT 36.255 119.005 37.040 119.175 ;
        RECT 35.680 118.775 35.850 119.005 ;
        RECT 35.020 118.475 35.850 118.775 ;
        RECT 36.235 118.505 36.700 118.835 ;
        RECT 35.020 118.445 35.220 118.475 ;
        RECT 35.340 118.225 35.510 118.295 ;
        RECT 34.640 118.055 35.510 118.225 ;
        RECT 35.000 117.965 35.510 118.055 ;
        RECT 33.550 117.500 33.855 117.630 ;
        RECT 34.300 117.520 34.830 117.885 ;
        RECT 33.170 116.905 33.435 117.365 ;
        RECT 33.605 117.075 33.855 117.500 ;
        RECT 35.000 117.350 35.170 117.965 ;
        RECT 34.065 117.180 35.170 117.350 ;
        RECT 35.340 116.905 35.510 117.705 ;
        RECT 35.680 117.405 35.850 118.475 ;
        RECT 36.020 117.575 36.210 118.295 ;
        RECT 36.380 117.545 36.700 118.505 ;
        RECT 36.870 118.545 37.040 119.005 ;
        RECT 37.315 118.925 37.525 119.455 ;
        RECT 37.785 118.715 38.115 119.240 ;
        RECT 38.285 118.845 38.455 119.455 ;
        RECT 38.625 118.800 38.955 119.235 ;
        RECT 38.625 118.715 39.005 118.800 ;
        RECT 39.175 118.730 39.465 119.455 ;
        RECT 37.915 118.545 38.115 118.715 ;
        RECT 38.780 118.675 39.005 118.715 ;
        RECT 36.870 118.215 37.745 118.545 ;
        RECT 37.915 118.215 38.665 118.545 ;
        RECT 35.680 117.075 35.930 117.405 ;
        RECT 36.870 117.375 37.040 118.215 ;
        RECT 37.915 118.010 38.105 118.215 ;
        RECT 38.835 118.095 39.005 118.675 ;
        RECT 38.790 118.045 39.005 118.095 ;
        RECT 39.635 118.510 39.975 119.285 ;
        RECT 40.145 118.995 40.315 119.455 ;
        RECT 40.555 119.020 40.915 119.285 ;
        RECT 40.555 119.015 40.910 119.020 ;
        RECT 40.555 119.005 40.905 119.015 ;
        RECT 40.555 119.000 40.900 119.005 ;
        RECT 40.555 118.990 40.895 119.000 ;
        RECT 41.545 118.995 41.715 119.455 ;
        RECT 40.555 118.985 40.890 118.990 ;
        RECT 40.555 118.975 40.880 118.985 ;
        RECT 40.555 118.965 40.870 118.975 ;
        RECT 40.555 118.825 40.855 118.965 ;
        RECT 40.145 118.635 40.855 118.825 ;
        RECT 41.045 118.825 41.375 118.905 ;
        RECT 41.885 118.825 42.225 119.285 ;
        RECT 41.045 118.635 42.225 118.825 ;
        RECT 42.595 118.825 42.925 119.185 ;
        RECT 43.545 118.995 43.795 119.455 ;
        RECT 43.965 118.995 44.525 119.285 ;
        RECT 42.595 118.635 43.985 118.825 ;
        RECT 37.210 117.635 38.105 118.010 ;
        RECT 38.615 117.965 39.005 118.045 ;
        RECT 36.155 117.205 37.040 117.375 ;
        RECT 37.220 116.905 37.535 117.405 ;
        RECT 37.765 117.075 38.105 117.635 ;
        RECT 38.275 116.905 38.445 117.915 ;
        RECT 38.615 117.120 38.945 117.965 ;
        RECT 39.175 116.905 39.465 118.070 ;
        RECT 39.635 117.075 39.915 118.510 ;
        RECT 40.145 118.065 40.430 118.635 ;
        RECT 43.815 118.545 43.985 118.635 ;
        RECT 40.615 118.235 41.085 118.465 ;
        RECT 41.255 118.445 41.585 118.465 ;
        RECT 41.255 118.265 41.705 118.445 ;
        RECT 41.895 118.265 42.225 118.465 ;
        RECT 40.145 117.850 41.295 118.065 ;
        RECT 40.085 116.905 40.795 117.680 ;
        RECT 40.965 117.075 41.295 117.850 ;
        RECT 41.490 117.150 41.705 118.265 ;
        RECT 41.995 117.925 42.225 118.265 ;
        RECT 42.410 118.215 43.085 118.465 ;
        RECT 43.305 118.215 43.645 118.465 ;
        RECT 43.815 118.215 44.105 118.545 ;
        RECT 42.410 117.855 42.675 118.215 ;
        RECT 43.815 117.965 43.985 118.215 ;
        RECT 43.045 117.795 43.985 117.965 ;
        RECT 41.885 116.905 42.215 117.625 ;
        RECT 42.595 116.905 42.875 117.575 ;
        RECT 43.045 117.245 43.345 117.795 ;
        RECT 44.275 117.625 44.525 118.995 ;
        RECT 44.695 118.685 46.365 119.455 ;
        RECT 47.005 118.725 47.305 119.455 ;
        RECT 44.695 118.165 45.445 118.685 ;
        RECT 47.485 118.545 47.715 119.165 ;
        RECT 47.915 118.895 48.140 119.275 ;
        RECT 48.310 119.065 48.640 119.455 ;
        RECT 48.925 118.905 49.095 119.195 ;
        RECT 49.265 119.075 49.595 119.455 ;
        RECT 47.915 118.715 48.245 118.895 ;
        RECT 45.615 117.995 46.365 118.515 ;
        RECT 47.010 118.215 47.305 118.545 ;
        RECT 47.485 118.215 47.900 118.545 ;
        RECT 48.070 118.045 48.245 118.715 ;
        RECT 48.415 118.215 48.655 118.865 ;
        RECT 48.925 118.735 49.590 118.905 ;
        RECT 43.545 116.905 43.875 117.625 ;
        RECT 44.065 117.075 44.525 117.625 ;
        RECT 44.695 116.905 46.365 117.995 ;
        RECT 47.005 117.685 47.900 118.015 ;
        RECT 48.070 117.855 48.655 118.045 ;
        RECT 48.840 117.915 49.190 118.565 ;
        RECT 47.005 117.515 48.210 117.685 ;
        RECT 47.005 117.085 47.335 117.515 ;
        RECT 47.515 116.905 47.710 117.345 ;
        RECT 47.880 117.085 48.210 117.515 ;
        RECT 48.380 117.085 48.655 117.855 ;
        RECT 49.360 117.745 49.590 118.735 ;
        RECT 48.925 117.575 49.590 117.745 ;
        RECT 48.925 117.075 49.095 117.575 ;
        RECT 49.265 116.905 49.595 117.405 ;
        RECT 49.765 117.075 49.950 119.195 ;
        RECT 50.205 118.995 50.455 119.455 ;
        RECT 50.625 119.005 50.960 119.175 ;
        RECT 51.155 119.005 51.830 119.175 ;
        RECT 50.625 118.865 50.795 119.005 ;
        RECT 50.120 117.875 50.400 118.825 ;
        RECT 50.570 118.735 50.795 118.865 ;
        RECT 50.570 117.630 50.740 118.735 ;
        RECT 50.965 118.585 51.490 118.805 ;
        RECT 50.910 117.820 51.150 118.415 ;
        RECT 51.320 117.885 51.490 118.585 ;
        RECT 51.660 118.225 51.830 119.005 ;
        RECT 52.150 118.955 52.520 119.455 ;
        RECT 52.700 119.005 53.105 119.175 ;
        RECT 53.275 119.005 54.060 119.175 ;
        RECT 52.700 118.775 52.870 119.005 ;
        RECT 52.040 118.475 52.870 118.775 ;
        RECT 53.255 118.505 53.720 118.835 ;
        RECT 52.040 118.445 52.240 118.475 ;
        RECT 52.360 118.225 52.530 118.295 ;
        RECT 51.660 118.055 52.530 118.225 ;
        RECT 52.020 117.965 52.530 118.055 ;
        RECT 50.570 117.500 50.875 117.630 ;
        RECT 51.320 117.520 51.850 117.885 ;
        RECT 50.190 116.905 50.455 117.365 ;
        RECT 50.625 117.075 50.875 117.500 ;
        RECT 52.020 117.350 52.190 117.965 ;
        RECT 51.085 117.180 52.190 117.350 ;
        RECT 52.360 116.905 52.530 117.705 ;
        RECT 52.700 117.405 52.870 118.475 ;
        RECT 53.040 117.575 53.230 118.295 ;
        RECT 53.400 117.545 53.720 118.505 ;
        RECT 53.890 118.545 54.060 119.005 ;
        RECT 54.335 118.925 54.545 119.455 ;
        RECT 54.805 118.715 55.135 119.240 ;
        RECT 55.305 118.845 55.475 119.455 ;
        RECT 55.645 118.800 55.975 119.235 ;
        RECT 56.255 118.995 56.500 119.455 ;
        RECT 55.645 118.715 56.025 118.800 ;
        RECT 54.935 118.545 55.135 118.715 ;
        RECT 55.800 118.675 56.025 118.715 ;
        RECT 53.890 118.215 54.765 118.545 ;
        RECT 54.935 118.215 55.685 118.545 ;
        RECT 52.700 117.075 52.950 117.405 ;
        RECT 53.890 117.375 54.060 118.215 ;
        RECT 54.935 118.010 55.125 118.215 ;
        RECT 55.855 118.095 56.025 118.675 ;
        RECT 56.195 118.215 56.510 118.825 ;
        RECT 56.680 118.465 56.930 119.275 ;
        RECT 57.100 118.930 57.360 119.455 ;
        RECT 57.530 118.805 57.790 119.260 ;
        RECT 57.960 118.975 58.220 119.455 ;
        RECT 58.390 118.805 58.650 119.260 ;
        RECT 58.820 118.975 59.080 119.455 ;
        RECT 59.250 118.805 59.510 119.260 ;
        RECT 59.680 118.975 59.940 119.455 ;
        RECT 60.110 118.805 60.370 119.260 ;
        RECT 60.540 118.975 60.840 119.455 ;
        RECT 61.370 118.825 61.655 119.285 ;
        RECT 61.825 118.995 62.095 119.455 ;
        RECT 57.530 118.635 60.840 118.805 ;
        RECT 61.370 118.655 62.325 118.825 ;
        RECT 56.680 118.215 59.700 118.465 ;
        RECT 55.810 118.045 56.025 118.095 ;
        RECT 54.230 117.635 55.125 118.010 ;
        RECT 55.635 117.965 56.025 118.045 ;
        RECT 53.175 117.205 54.060 117.375 ;
        RECT 54.240 116.905 54.555 117.405 ;
        RECT 54.785 117.075 55.125 117.635 ;
        RECT 55.295 116.905 55.465 117.915 ;
        RECT 55.635 117.120 55.965 117.965 ;
        RECT 56.205 116.905 56.500 118.015 ;
        RECT 56.680 117.080 56.930 118.215 ;
        RECT 59.870 118.045 60.840 118.635 ;
        RECT 57.100 116.905 57.360 118.015 ;
        RECT 57.530 117.805 60.840 118.045 ;
        RECT 61.255 117.925 61.945 118.485 ;
        RECT 57.530 117.080 57.790 117.805 ;
        RECT 57.960 116.905 58.220 117.635 ;
        RECT 58.390 117.080 58.650 117.805 ;
        RECT 58.820 116.905 59.080 117.635 ;
        RECT 59.250 117.080 59.510 117.805 ;
        RECT 59.680 116.905 59.940 117.635 ;
        RECT 60.110 117.080 60.370 117.805 ;
        RECT 62.115 117.755 62.325 118.655 ;
        RECT 60.540 116.905 60.835 117.635 ;
        RECT 61.370 117.535 62.325 117.755 ;
        RECT 62.495 118.485 62.895 119.285 ;
        RECT 63.085 118.825 63.365 119.285 ;
        RECT 63.885 118.995 64.210 119.455 ;
        RECT 63.085 118.655 64.210 118.825 ;
        RECT 64.380 118.715 64.765 119.285 ;
        RECT 64.935 118.730 65.225 119.455 ;
        RECT 65.485 118.905 65.655 119.195 ;
        RECT 65.825 119.075 66.155 119.455 ;
        RECT 65.485 118.735 66.150 118.905 ;
        RECT 63.760 118.545 64.210 118.655 ;
        RECT 62.495 117.925 63.590 118.485 ;
        RECT 63.760 118.215 64.315 118.545 ;
        RECT 61.370 117.075 61.655 117.535 ;
        RECT 61.825 116.905 62.095 117.365 ;
        RECT 62.495 117.075 62.895 117.925 ;
        RECT 63.760 117.755 64.210 118.215 ;
        RECT 64.485 118.045 64.765 118.715 ;
        RECT 63.085 117.535 64.210 117.755 ;
        RECT 63.085 117.075 63.365 117.535 ;
        RECT 63.885 116.905 64.210 117.365 ;
        RECT 64.380 117.075 64.765 118.045 ;
        RECT 64.935 116.905 65.225 118.070 ;
        RECT 65.400 117.915 65.750 118.565 ;
        RECT 65.920 117.745 66.150 118.735 ;
        RECT 65.485 117.575 66.150 117.745 ;
        RECT 65.485 117.075 65.655 117.575 ;
        RECT 65.825 116.905 66.155 117.405 ;
        RECT 66.325 117.075 66.510 119.195 ;
        RECT 66.765 118.995 67.015 119.455 ;
        RECT 67.185 119.005 67.520 119.175 ;
        RECT 67.715 119.005 68.390 119.175 ;
        RECT 67.185 118.865 67.355 119.005 ;
        RECT 66.680 117.875 66.960 118.825 ;
        RECT 67.130 118.735 67.355 118.865 ;
        RECT 67.130 117.630 67.300 118.735 ;
        RECT 67.525 118.585 68.050 118.805 ;
        RECT 67.470 117.820 67.710 118.415 ;
        RECT 67.880 117.885 68.050 118.585 ;
        RECT 68.220 118.225 68.390 119.005 ;
        RECT 68.710 118.955 69.080 119.455 ;
        RECT 69.260 119.005 69.665 119.175 ;
        RECT 69.835 119.005 70.620 119.175 ;
        RECT 69.260 118.775 69.430 119.005 ;
        RECT 68.600 118.475 69.430 118.775 ;
        RECT 69.815 118.505 70.280 118.835 ;
        RECT 68.600 118.445 68.800 118.475 ;
        RECT 68.920 118.225 69.090 118.295 ;
        RECT 68.220 118.055 69.090 118.225 ;
        RECT 68.580 117.965 69.090 118.055 ;
        RECT 67.130 117.500 67.435 117.630 ;
        RECT 67.880 117.520 68.410 117.885 ;
        RECT 66.750 116.905 67.015 117.365 ;
        RECT 67.185 117.075 67.435 117.500 ;
        RECT 68.580 117.350 68.750 117.965 ;
        RECT 67.645 117.180 68.750 117.350 ;
        RECT 68.920 116.905 69.090 117.705 ;
        RECT 69.260 117.405 69.430 118.475 ;
        RECT 69.600 117.575 69.790 118.295 ;
        RECT 69.960 117.545 70.280 118.505 ;
        RECT 70.450 118.545 70.620 119.005 ;
        RECT 70.895 118.925 71.105 119.455 ;
        RECT 71.365 118.715 71.695 119.240 ;
        RECT 71.865 118.845 72.035 119.455 ;
        RECT 72.205 118.800 72.535 119.235 ;
        RECT 72.205 118.715 72.585 118.800 ;
        RECT 71.495 118.545 71.695 118.715 ;
        RECT 72.360 118.675 72.585 118.715 ;
        RECT 70.450 118.215 71.325 118.545 ;
        RECT 71.495 118.215 72.245 118.545 ;
        RECT 69.260 117.075 69.510 117.405 ;
        RECT 70.450 117.375 70.620 118.215 ;
        RECT 71.495 118.010 71.685 118.215 ;
        RECT 72.415 118.095 72.585 118.675 ;
        RECT 72.370 118.045 72.585 118.095 ;
        RECT 70.790 117.635 71.685 118.010 ;
        RECT 72.195 117.965 72.585 118.045 ;
        RECT 72.790 118.715 73.405 119.285 ;
        RECT 73.575 118.945 73.790 119.455 ;
        RECT 74.020 118.945 74.300 119.275 ;
        RECT 74.480 118.945 74.720 119.455 ;
        RECT 69.735 117.205 70.620 117.375 ;
        RECT 70.800 116.905 71.115 117.405 ;
        RECT 71.345 117.075 71.685 117.635 ;
        RECT 71.855 116.905 72.025 117.915 ;
        RECT 72.195 117.120 72.525 117.965 ;
        RECT 72.790 117.695 73.105 118.715 ;
        RECT 73.275 118.045 73.445 118.545 ;
        RECT 73.695 118.215 73.960 118.775 ;
        RECT 74.130 118.045 74.300 118.945 ;
        RECT 75.060 118.925 75.350 119.275 ;
        RECT 75.545 119.095 75.875 119.455 ;
        RECT 76.045 118.925 76.275 119.230 ;
        RECT 74.470 118.215 74.825 118.775 ;
        RECT 75.060 118.755 76.275 118.925 ;
        RECT 76.465 118.585 76.635 119.150 ;
        RECT 76.985 118.905 77.155 119.195 ;
        RECT 77.325 119.075 77.655 119.455 ;
        RECT 76.985 118.735 77.650 118.905 ;
        RECT 75.120 118.435 75.380 118.545 ;
        RECT 75.115 118.265 75.380 118.435 ;
        RECT 75.120 118.215 75.380 118.265 ;
        RECT 75.560 118.215 75.945 118.545 ;
        RECT 76.115 118.415 76.635 118.585 ;
        RECT 73.275 117.875 74.700 118.045 ;
        RECT 72.790 117.075 73.325 117.695 ;
        RECT 73.495 116.905 73.825 117.705 ;
        RECT 74.310 117.700 74.700 117.875 ;
        RECT 75.060 116.905 75.380 118.045 ;
        RECT 75.560 117.165 75.755 118.215 ;
        RECT 76.115 118.035 76.285 118.415 ;
        RECT 75.935 117.755 76.285 118.035 ;
        RECT 76.475 117.885 76.720 118.245 ;
        RECT 76.900 117.915 77.250 118.565 ;
        RECT 75.935 117.075 76.265 117.755 ;
        RECT 77.420 117.745 77.650 118.735 ;
        RECT 76.465 116.905 76.720 117.705 ;
        RECT 76.985 117.575 77.650 117.745 ;
        RECT 76.985 117.075 77.155 117.575 ;
        RECT 77.325 116.905 77.655 117.405 ;
        RECT 77.825 117.075 78.010 119.195 ;
        RECT 78.265 118.995 78.515 119.455 ;
        RECT 78.685 119.005 79.020 119.175 ;
        RECT 79.215 119.005 79.890 119.175 ;
        RECT 78.685 118.865 78.855 119.005 ;
        RECT 78.180 117.875 78.460 118.825 ;
        RECT 78.630 118.735 78.855 118.865 ;
        RECT 78.630 117.630 78.800 118.735 ;
        RECT 79.025 118.585 79.550 118.805 ;
        RECT 78.970 117.820 79.210 118.415 ;
        RECT 79.380 117.885 79.550 118.585 ;
        RECT 79.720 118.225 79.890 119.005 ;
        RECT 80.210 118.955 80.580 119.455 ;
        RECT 80.760 119.005 81.165 119.175 ;
        RECT 81.335 119.005 82.120 119.175 ;
        RECT 80.760 118.775 80.930 119.005 ;
        RECT 80.100 118.475 80.930 118.775 ;
        RECT 81.315 118.505 81.780 118.835 ;
        RECT 80.100 118.445 80.300 118.475 ;
        RECT 80.420 118.225 80.590 118.295 ;
        RECT 79.720 118.055 80.590 118.225 ;
        RECT 80.080 117.965 80.590 118.055 ;
        RECT 78.630 117.500 78.935 117.630 ;
        RECT 79.380 117.520 79.910 117.885 ;
        RECT 78.250 116.905 78.515 117.365 ;
        RECT 78.685 117.075 78.935 117.500 ;
        RECT 80.080 117.350 80.250 117.965 ;
        RECT 79.145 117.180 80.250 117.350 ;
        RECT 80.420 116.905 80.590 117.705 ;
        RECT 80.760 117.405 80.930 118.475 ;
        RECT 81.100 117.575 81.290 118.295 ;
        RECT 81.460 117.545 81.780 118.505 ;
        RECT 81.950 118.545 82.120 119.005 ;
        RECT 82.395 118.925 82.605 119.455 ;
        RECT 82.865 118.715 83.195 119.240 ;
        RECT 83.365 118.845 83.535 119.455 ;
        RECT 83.705 118.800 84.035 119.235 ;
        RECT 84.205 118.940 84.375 119.455 ;
        RECT 83.705 118.715 84.085 118.800 ;
        RECT 82.995 118.545 83.195 118.715 ;
        RECT 83.860 118.675 84.085 118.715 ;
        RECT 81.950 118.215 82.825 118.545 ;
        RECT 82.995 118.215 83.745 118.545 ;
        RECT 80.760 117.075 81.010 117.405 ;
        RECT 81.950 117.375 82.120 118.215 ;
        RECT 82.995 118.010 83.185 118.215 ;
        RECT 83.915 118.095 84.085 118.675 ;
        RECT 84.715 118.685 87.305 119.455 ;
        RECT 87.475 118.955 87.775 119.285 ;
        RECT 87.945 118.975 88.220 119.455 ;
        RECT 84.715 118.165 85.925 118.685 ;
        RECT 83.870 118.045 84.085 118.095 ;
        RECT 82.290 117.635 83.185 118.010 ;
        RECT 83.695 117.965 84.085 118.045 ;
        RECT 86.095 117.995 87.305 118.515 ;
        RECT 81.235 117.205 82.120 117.375 ;
        RECT 82.300 116.905 82.615 117.405 ;
        RECT 82.845 117.075 83.185 117.635 ;
        RECT 83.355 116.905 83.525 117.915 ;
        RECT 83.695 117.120 84.025 117.965 ;
        RECT 84.195 116.905 84.365 117.820 ;
        RECT 84.715 116.905 87.305 117.995 ;
        RECT 87.475 118.045 87.645 118.955 ;
        RECT 88.400 118.805 88.695 119.195 ;
        RECT 88.865 118.975 89.120 119.455 ;
        RECT 89.295 118.805 89.555 119.195 ;
        RECT 89.725 118.975 90.005 119.455 ;
        RECT 87.815 118.215 88.165 118.785 ;
        RECT 88.400 118.635 90.050 118.805 ;
        RECT 90.695 118.730 90.985 119.455 ;
        RECT 91.215 118.995 91.460 119.455 ;
        RECT 88.335 118.295 89.475 118.465 ;
        RECT 88.335 118.045 88.505 118.295 ;
        RECT 89.645 118.125 90.050 118.635 ;
        RECT 91.155 118.215 91.470 118.825 ;
        RECT 91.640 118.465 91.890 119.275 ;
        RECT 92.060 118.930 92.320 119.455 ;
        RECT 92.490 118.805 92.750 119.260 ;
        RECT 92.920 118.975 93.180 119.455 ;
        RECT 93.350 118.805 93.610 119.260 ;
        RECT 93.780 118.975 94.040 119.455 ;
        RECT 94.210 118.805 94.470 119.260 ;
        RECT 94.640 118.975 94.900 119.455 ;
        RECT 95.070 118.805 95.330 119.260 ;
        RECT 95.500 118.975 95.800 119.455 ;
        RECT 92.490 118.635 95.800 118.805 ;
        RECT 96.255 118.635 96.485 119.455 ;
        RECT 96.655 118.655 96.985 119.285 ;
        RECT 91.640 118.215 94.660 118.465 ;
        RECT 87.475 117.875 88.505 118.045 ;
        RECT 89.295 117.955 90.050 118.125 ;
        RECT 87.475 117.075 87.785 117.875 ;
        RECT 89.295 117.705 89.555 117.955 ;
        RECT 87.955 116.905 88.265 117.705 ;
        RECT 88.435 117.535 89.555 117.705 ;
        RECT 88.435 117.075 88.695 117.535 ;
        RECT 88.865 116.905 89.120 117.365 ;
        RECT 89.295 117.075 89.555 117.535 ;
        RECT 89.725 116.905 90.010 117.775 ;
        RECT 90.695 116.905 90.985 118.070 ;
        RECT 91.165 116.905 91.460 118.015 ;
        RECT 91.640 117.080 91.890 118.215 ;
        RECT 94.830 118.045 95.800 118.635 ;
        RECT 96.235 118.215 96.565 118.465 ;
        RECT 96.735 118.055 96.985 118.655 ;
        RECT 97.155 118.635 97.365 119.455 ;
        RECT 97.595 118.705 98.805 119.455 ;
        RECT 98.975 118.795 99.250 119.455 ;
        RECT 99.420 118.825 99.670 119.285 ;
        RECT 99.845 118.960 100.175 119.455 ;
        RECT 97.595 118.165 98.115 118.705 ;
        RECT 99.420 118.615 99.590 118.825 ;
        RECT 100.355 118.790 100.585 119.235 ;
        RECT 92.060 116.905 92.320 118.015 ;
        RECT 92.490 117.805 95.800 118.045 ;
        RECT 92.490 117.080 92.750 117.805 ;
        RECT 92.920 116.905 93.180 117.635 ;
        RECT 93.350 117.080 93.610 117.805 ;
        RECT 93.780 116.905 94.040 117.635 ;
        RECT 94.210 117.080 94.470 117.805 ;
        RECT 94.640 116.905 94.900 117.635 ;
        RECT 95.070 117.080 95.330 117.805 ;
        RECT 95.500 116.905 95.795 117.635 ;
        RECT 96.255 116.905 96.485 118.045 ;
        RECT 96.655 117.075 96.985 118.055 ;
        RECT 97.155 116.905 97.365 118.045 ;
        RECT 98.285 117.995 98.805 118.535 ;
        RECT 98.975 118.095 99.590 118.615 ;
        RECT 99.760 118.115 99.990 118.545 ;
        RECT 100.175 118.295 100.585 118.790 ;
        RECT 100.755 118.970 101.545 119.235 ;
        RECT 100.755 118.115 101.010 118.970 ;
        RECT 101.735 118.815 102.025 119.285 ;
        RECT 102.225 118.985 102.395 119.455 ;
        RECT 102.565 118.815 102.895 119.285 ;
        RECT 103.065 118.985 103.235 119.455 ;
        RECT 103.405 118.815 103.735 119.285 ;
        RECT 103.905 118.985 104.075 119.455 ;
        RECT 104.245 118.815 104.575 119.285 ;
        RECT 104.745 118.985 104.915 119.455 ;
        RECT 105.085 118.815 105.415 119.285 ;
        RECT 105.585 118.985 105.755 119.455 ;
        RECT 105.925 118.815 106.255 119.285 ;
        RECT 106.425 118.985 106.595 119.455 ;
        RECT 106.765 118.815 107.095 119.285 ;
        RECT 101.180 118.295 101.565 118.775 ;
        RECT 101.735 118.635 107.095 118.815 ;
        RECT 107.265 118.635 107.540 119.455 ;
        RECT 107.715 118.955 107.975 119.285 ;
        RECT 108.185 118.975 108.460 119.455 ;
        RECT 97.595 116.905 98.805 117.995 ;
        RECT 98.975 116.905 99.235 117.915 ;
        RECT 99.405 117.755 99.575 118.095 ;
        RECT 99.760 117.945 101.550 118.115 ;
        RECT 99.405 117.745 99.665 117.755 ;
        RECT 99.405 117.075 99.680 117.745 ;
        RECT 99.880 116.905 100.095 117.750 ;
        RECT 100.320 117.650 100.570 117.945 ;
        RECT 100.795 117.585 101.125 117.775 ;
        RECT 100.280 117.075 100.755 117.415 ;
        RECT 100.935 117.410 101.125 117.585 ;
        RECT 101.295 117.580 101.550 117.945 ;
        RECT 101.735 117.755 102.025 118.635 ;
        RECT 102.215 118.255 102.635 118.465 ;
        RECT 102.865 118.265 103.775 118.465 ;
        RECT 102.465 118.095 102.635 118.255 ;
        RECT 103.945 118.255 105.535 118.465 ;
        RECT 105.805 118.255 107.540 118.465 ;
        RECT 103.945 118.095 104.115 118.255 ;
        RECT 102.465 117.925 104.115 118.095 ;
        RECT 104.285 117.915 105.375 118.085 ;
        RECT 101.735 117.585 104.115 117.755 ;
        RECT 100.935 116.905 101.565 117.410 ;
        RECT 101.735 117.075 102.015 117.585 ;
        RECT 103.025 117.575 104.115 117.585 ;
        RECT 103.025 117.415 103.275 117.575 ;
        RECT 103.865 117.415 104.115 117.575 ;
        RECT 102.185 117.075 102.435 117.415 ;
        RECT 102.605 117.245 102.855 117.405 ;
        RECT 103.445 117.245 103.695 117.405 ;
        RECT 104.285 117.245 104.535 117.915 ;
        RECT 102.605 117.075 104.535 117.245 ;
        RECT 104.705 117.455 104.955 117.745 ;
        RECT 105.125 117.625 105.375 117.915 ;
        RECT 105.545 117.915 107.480 118.085 ;
        RECT 105.545 117.455 105.795 117.915 ;
        RECT 104.705 117.075 105.795 117.455 ;
        RECT 105.965 116.905 106.215 117.745 ;
        RECT 106.385 117.075 106.635 117.915 ;
        RECT 106.805 116.905 107.055 117.745 ;
        RECT 107.225 117.075 107.480 117.915 ;
        RECT 107.715 118.045 107.885 118.955 ;
        RECT 108.670 118.885 108.875 119.285 ;
        RECT 109.045 119.055 109.380 119.455 ;
        RECT 108.055 118.215 108.415 118.795 ;
        RECT 108.670 118.715 109.355 118.885 ;
        RECT 108.595 118.045 108.845 118.545 ;
        RECT 107.715 117.875 108.845 118.045 ;
        RECT 107.715 117.105 107.985 117.875 ;
        RECT 109.015 117.685 109.355 118.715 ;
        RECT 109.555 118.685 113.065 119.455 ;
        RECT 114.265 119.075 115.435 119.285 ;
        RECT 114.265 119.055 114.595 119.075 ;
        RECT 109.555 118.165 111.205 118.685 ;
        RECT 114.155 118.635 115.015 118.885 ;
        RECT 115.185 118.825 115.435 119.075 ;
        RECT 115.605 118.995 115.775 119.455 ;
        RECT 115.945 118.825 116.285 119.285 ;
        RECT 115.185 118.655 116.285 118.825 ;
        RECT 116.455 118.730 116.745 119.455 ;
        RECT 116.915 118.955 117.175 119.285 ;
        RECT 117.345 119.095 117.675 119.455 ;
        RECT 117.930 119.075 119.230 119.285 ;
        RECT 111.375 117.995 113.065 118.515 ;
        RECT 108.155 116.905 108.485 117.685 ;
        RECT 108.690 117.510 109.355 117.685 ;
        RECT 108.690 117.105 108.875 117.510 ;
        RECT 109.045 116.905 109.380 117.330 ;
        RECT 109.555 116.905 113.065 117.995 ;
        RECT 114.155 118.045 114.435 118.635 ;
        RECT 114.605 118.215 115.355 118.465 ;
        RECT 115.525 118.215 116.285 118.465 ;
        RECT 114.155 117.875 115.855 118.045 ;
        RECT 114.260 116.905 114.515 117.705 ;
        RECT 114.685 117.075 115.015 117.875 ;
        RECT 115.185 116.905 115.355 117.705 ;
        RECT 115.525 117.075 115.855 117.875 ;
        RECT 116.025 116.905 116.285 118.045 ;
        RECT 116.455 116.905 116.745 118.070 ;
        RECT 116.915 117.755 117.085 118.955 ;
        RECT 117.930 118.925 118.100 119.075 ;
        RECT 117.345 118.800 118.100 118.925 ;
        RECT 117.255 118.755 118.100 118.800 ;
        RECT 117.255 118.635 117.525 118.755 ;
        RECT 117.255 118.060 117.425 118.635 ;
        RECT 117.655 118.195 118.065 118.500 ;
        RECT 118.355 118.465 118.565 118.865 ;
        RECT 118.235 118.255 118.565 118.465 ;
        RECT 118.810 118.465 119.030 118.865 ;
        RECT 119.505 118.690 119.960 119.455 ;
        RECT 120.135 118.955 120.435 119.285 ;
        RECT 120.605 118.975 120.880 119.455 ;
        RECT 118.810 118.255 119.285 118.465 ;
        RECT 119.475 118.265 119.965 118.465 ;
        RECT 117.255 118.025 117.455 118.060 ;
        RECT 118.785 118.025 119.960 118.085 ;
        RECT 117.255 117.915 119.960 118.025 ;
        RECT 117.315 117.855 119.115 117.915 ;
        RECT 118.785 117.825 119.115 117.855 ;
        RECT 116.915 117.075 117.175 117.755 ;
        RECT 117.345 116.905 117.595 117.685 ;
        RECT 117.845 117.655 118.680 117.665 ;
        RECT 119.270 117.655 119.455 117.745 ;
        RECT 117.845 117.455 119.455 117.655 ;
        RECT 117.845 117.075 118.095 117.455 ;
        RECT 119.225 117.415 119.455 117.455 ;
        RECT 119.705 117.295 119.960 117.915 ;
        RECT 118.265 116.905 118.620 117.285 ;
        RECT 119.625 117.075 119.960 117.295 ;
        RECT 120.135 118.045 120.305 118.955 ;
        RECT 121.060 118.805 121.355 119.195 ;
        RECT 121.525 118.975 121.780 119.455 ;
        RECT 121.955 118.805 122.215 119.195 ;
        RECT 122.385 118.975 122.665 119.455 ;
        RECT 120.475 118.215 120.825 118.785 ;
        RECT 121.060 118.635 122.710 118.805 ;
        RECT 123.560 118.675 124.060 119.285 ;
        RECT 120.995 118.295 122.135 118.465 ;
        RECT 120.995 118.045 121.165 118.295 ;
        RECT 122.305 118.125 122.710 118.635 ;
        RECT 123.355 118.215 123.705 118.465 ;
        RECT 120.135 117.875 121.165 118.045 ;
        RECT 121.955 117.955 122.710 118.125 ;
        RECT 123.890 118.045 124.060 118.675 ;
        RECT 124.690 118.805 125.020 119.285 ;
        RECT 125.190 118.995 125.415 119.455 ;
        RECT 125.585 118.805 125.915 119.285 ;
        RECT 124.690 118.635 125.915 118.805 ;
        RECT 126.105 118.655 126.355 119.455 ;
        RECT 126.525 118.655 126.865 119.285 ;
        RECT 127.125 118.905 127.295 119.195 ;
        RECT 127.465 119.075 127.795 119.455 ;
        RECT 127.125 118.735 127.790 118.905 ;
        RECT 124.230 118.265 124.560 118.465 ;
        RECT 124.730 118.265 125.060 118.465 ;
        RECT 125.230 118.265 125.650 118.465 ;
        RECT 125.825 118.295 126.520 118.465 ;
        RECT 125.825 118.045 125.995 118.295 ;
        RECT 126.690 118.045 126.865 118.655 ;
        RECT 120.135 117.075 120.445 117.875 ;
        RECT 121.955 117.705 122.215 117.955 ;
        RECT 123.560 117.875 125.995 118.045 ;
        RECT 120.615 116.905 120.925 117.705 ;
        RECT 121.095 117.535 122.215 117.705 ;
        RECT 121.095 117.075 121.355 117.535 ;
        RECT 121.525 116.905 121.780 117.365 ;
        RECT 121.955 117.075 122.215 117.535 ;
        RECT 122.385 116.905 122.670 117.775 ;
        RECT 123.560 117.075 123.890 117.875 ;
        RECT 124.060 116.905 124.390 117.705 ;
        RECT 124.690 117.075 125.020 117.875 ;
        RECT 125.665 116.905 125.915 117.705 ;
        RECT 126.185 116.905 126.355 118.045 ;
        RECT 126.525 117.075 126.865 118.045 ;
        RECT 127.040 117.915 127.390 118.565 ;
        RECT 127.560 117.745 127.790 118.735 ;
        RECT 127.125 117.575 127.790 117.745 ;
        RECT 127.125 117.075 127.295 117.575 ;
        RECT 127.465 116.905 127.795 117.405 ;
        RECT 127.965 117.075 128.150 119.195 ;
        RECT 128.405 118.995 128.655 119.455 ;
        RECT 128.825 119.005 129.160 119.175 ;
        RECT 129.355 119.005 130.030 119.175 ;
        RECT 128.825 118.865 128.995 119.005 ;
        RECT 128.320 117.875 128.600 118.825 ;
        RECT 128.770 118.735 128.995 118.865 ;
        RECT 128.770 117.630 128.940 118.735 ;
        RECT 129.165 118.585 129.690 118.805 ;
        RECT 129.110 117.820 129.350 118.415 ;
        RECT 129.520 117.885 129.690 118.585 ;
        RECT 129.860 118.225 130.030 119.005 ;
        RECT 130.350 118.955 130.720 119.455 ;
        RECT 130.900 119.005 131.305 119.175 ;
        RECT 131.475 119.005 132.260 119.175 ;
        RECT 130.900 118.775 131.070 119.005 ;
        RECT 130.240 118.475 131.070 118.775 ;
        RECT 131.455 118.505 131.920 118.835 ;
        RECT 130.240 118.445 130.440 118.475 ;
        RECT 130.560 118.225 130.730 118.295 ;
        RECT 129.860 118.055 130.730 118.225 ;
        RECT 130.220 117.965 130.730 118.055 ;
        RECT 128.770 117.500 129.075 117.630 ;
        RECT 129.520 117.520 130.050 117.885 ;
        RECT 128.390 116.905 128.655 117.365 ;
        RECT 128.825 117.075 129.075 117.500 ;
        RECT 130.220 117.350 130.390 117.965 ;
        RECT 129.285 117.180 130.390 117.350 ;
        RECT 130.560 116.905 130.730 117.705 ;
        RECT 130.900 117.405 131.070 118.475 ;
        RECT 131.240 117.575 131.430 118.295 ;
        RECT 131.600 117.545 131.920 118.505 ;
        RECT 132.090 118.545 132.260 119.005 ;
        RECT 132.535 118.925 132.745 119.455 ;
        RECT 133.005 118.715 133.335 119.240 ;
        RECT 133.505 118.845 133.675 119.455 ;
        RECT 133.845 118.800 134.175 119.235 ;
        RECT 134.560 118.945 134.800 119.455 ;
        RECT 134.980 118.945 135.260 119.275 ;
        RECT 135.490 118.945 135.705 119.455 ;
        RECT 133.845 118.715 134.225 118.800 ;
        RECT 133.135 118.545 133.335 118.715 ;
        RECT 134.000 118.675 134.225 118.715 ;
        RECT 132.090 118.215 132.965 118.545 ;
        RECT 133.135 118.215 133.885 118.545 ;
        RECT 130.900 117.075 131.150 117.405 ;
        RECT 132.090 117.375 132.260 118.215 ;
        RECT 133.135 118.010 133.325 118.215 ;
        RECT 134.055 118.095 134.225 118.675 ;
        RECT 134.455 118.215 134.810 118.775 ;
        RECT 134.010 118.045 134.225 118.095 ;
        RECT 134.980 118.045 135.150 118.945 ;
        RECT 135.320 118.215 135.585 118.775 ;
        RECT 135.875 118.715 136.490 119.285 ;
        RECT 135.835 118.045 136.005 118.545 ;
        RECT 132.430 117.635 133.325 118.010 ;
        RECT 133.835 117.965 134.225 118.045 ;
        RECT 131.375 117.205 132.260 117.375 ;
        RECT 132.440 116.905 132.755 117.405 ;
        RECT 132.985 117.075 133.325 117.635 ;
        RECT 133.495 116.905 133.665 117.915 ;
        RECT 133.835 117.120 134.165 117.965 ;
        RECT 134.580 117.875 136.005 118.045 ;
        RECT 134.580 117.700 134.970 117.875 ;
        RECT 135.455 116.905 135.785 117.705 ;
        RECT 136.175 117.695 136.490 118.715 ;
        RECT 137.615 118.705 138.825 119.455 ;
        RECT 135.955 117.075 136.490 117.695 ;
        RECT 137.615 117.995 138.135 118.535 ;
        RECT 138.305 118.165 138.825 118.705 ;
        RECT 137.615 116.905 138.825 117.995 ;
        RECT 13.330 116.735 138.910 116.905 ;
        RECT 13.415 115.645 14.625 116.735 ;
        RECT 14.795 115.645 18.305 116.735 ;
        RECT 13.415 114.935 13.935 115.475 ;
        RECT 14.105 115.105 14.625 115.645 ;
        RECT 14.795 114.955 16.445 115.475 ;
        RECT 16.615 115.125 18.305 115.645 ;
        RECT 18.935 115.865 19.210 116.565 ;
        RECT 19.420 116.190 19.635 116.735 ;
        RECT 19.805 116.225 20.280 116.565 ;
        RECT 20.450 116.230 21.065 116.735 ;
        RECT 20.450 116.055 20.645 116.230 ;
        RECT 13.415 114.185 14.625 114.935 ;
        RECT 14.795 114.185 18.305 114.955 ;
        RECT 18.935 114.835 19.105 115.865 ;
        RECT 19.380 115.695 20.095 115.990 ;
        RECT 20.315 115.865 20.645 116.055 ;
        RECT 20.815 115.695 21.065 116.060 ;
        RECT 19.275 115.525 21.065 115.695 ;
        RECT 19.275 115.095 19.505 115.525 ;
        RECT 18.935 114.355 19.195 114.835 ;
        RECT 19.675 114.825 20.085 115.345 ;
        RECT 19.365 114.185 19.695 114.645 ;
        RECT 19.885 114.405 20.085 114.825 ;
        RECT 20.255 114.670 20.510 115.525 ;
        RECT 21.305 115.345 21.475 116.565 ;
        RECT 21.725 116.225 21.985 116.735 ;
        RECT 20.680 115.095 21.475 115.345 ;
        RECT 21.645 115.175 21.985 116.055 ;
        RECT 22.155 115.595 22.435 116.735 ;
        RECT 22.605 115.585 22.935 116.565 ;
        RECT 23.105 115.595 23.365 116.735 ;
        RECT 22.165 115.155 22.500 115.425 ;
        RECT 21.225 115.005 21.475 115.095 ;
        RECT 20.255 114.405 21.045 114.670 ;
        RECT 21.225 114.585 21.555 115.005 ;
        RECT 21.725 114.185 21.985 115.005 ;
        RECT 22.670 114.985 22.840 115.585 ;
        RECT 23.010 115.175 23.345 115.425 ;
        RECT 22.155 114.185 22.465 114.985 ;
        RECT 22.670 114.355 23.365 114.985 ;
        RECT 23.545 114.365 23.805 116.555 ;
        RECT 23.975 116.005 24.315 116.735 ;
        RECT 24.495 115.825 24.765 116.555 ;
        RECT 23.995 115.605 24.765 115.825 ;
        RECT 24.945 115.845 25.175 116.555 ;
        RECT 25.345 116.025 25.675 116.735 ;
        RECT 25.845 115.845 26.105 116.555 ;
        RECT 24.945 115.605 26.105 115.845 ;
        RECT 23.995 114.935 24.285 115.605 ;
        RECT 26.295 115.570 26.585 116.735 ;
        RECT 26.765 115.935 27.095 116.735 ;
        RECT 27.275 116.395 28.705 116.565 ;
        RECT 27.275 115.765 27.525 116.395 ;
        RECT 26.755 115.595 27.525 115.765 ;
        RECT 24.465 115.115 24.930 115.425 ;
        RECT 25.110 115.115 25.635 115.425 ;
        RECT 23.995 114.735 25.225 114.935 ;
        RECT 24.065 114.185 24.735 114.555 ;
        RECT 24.915 114.365 25.225 114.735 ;
        RECT 25.405 114.475 25.635 115.115 ;
        RECT 25.815 115.095 26.115 115.425 ;
        RECT 26.755 114.925 26.925 115.595 ;
        RECT 27.095 115.095 27.500 115.425 ;
        RECT 27.715 115.095 27.965 116.225 ;
        RECT 28.165 115.425 28.365 116.225 ;
        RECT 28.535 115.715 28.705 116.395 ;
        RECT 28.875 115.885 29.190 116.735 ;
        RECT 29.365 115.935 29.805 116.565 ;
        RECT 28.535 115.545 29.325 115.715 ;
        RECT 28.165 115.095 28.410 115.425 ;
        RECT 28.595 115.095 28.985 115.375 ;
        RECT 29.155 115.095 29.325 115.545 ;
        RECT 29.495 114.925 29.805 115.935 ;
        RECT 29.975 115.645 31.645 116.735 ;
        RECT 25.815 114.185 26.105 114.915 ;
        RECT 26.295 114.185 26.585 114.910 ;
        RECT 26.755 114.355 27.245 114.925 ;
        RECT 27.415 114.755 28.575 114.925 ;
        RECT 27.415 114.355 27.645 114.755 ;
        RECT 27.815 114.185 28.235 114.585 ;
        RECT 28.405 114.355 28.575 114.755 ;
        RECT 28.745 114.185 29.195 114.925 ;
        RECT 29.365 114.365 29.805 114.925 ;
        RECT 29.975 114.955 30.725 115.475 ;
        RECT 30.895 115.125 31.645 115.645 ;
        RECT 31.970 115.725 32.270 116.565 ;
        RECT 32.465 115.895 32.715 116.735 ;
        RECT 33.305 116.145 34.110 116.565 ;
        RECT 32.885 115.975 34.450 116.145 ;
        RECT 32.885 115.725 33.055 115.975 ;
        RECT 31.970 115.555 33.055 115.725 ;
        RECT 31.815 115.095 32.145 115.385 ;
        RECT 29.975 114.185 31.645 114.955 ;
        RECT 32.315 114.925 32.485 115.555 ;
        RECT 33.225 115.425 33.545 115.805 ;
        RECT 33.735 115.715 34.110 115.805 ;
        RECT 33.715 115.545 34.110 115.715 ;
        RECT 34.280 115.725 34.450 115.975 ;
        RECT 34.620 115.895 34.950 116.735 ;
        RECT 35.120 115.975 35.785 116.565 ;
        RECT 34.280 115.555 35.200 115.725 ;
        RECT 32.655 115.175 32.985 115.385 ;
        RECT 33.165 115.175 33.545 115.425 ;
        RECT 33.735 115.385 34.110 115.545 ;
        RECT 35.030 115.385 35.200 115.555 ;
        RECT 33.735 115.175 34.220 115.385 ;
        RECT 34.410 115.175 34.860 115.385 ;
        RECT 35.030 115.175 35.365 115.385 ;
        RECT 35.535 115.005 35.785 115.975 ;
        RECT 31.975 114.745 32.485 114.925 ;
        RECT 32.890 114.835 34.590 115.005 ;
        RECT 32.890 114.745 33.275 114.835 ;
        RECT 31.975 114.355 32.305 114.745 ;
        RECT 32.475 114.405 33.660 114.575 ;
        RECT 33.920 114.185 34.090 114.655 ;
        RECT 34.260 114.370 34.590 114.835 ;
        RECT 34.760 114.185 34.930 115.005 ;
        RECT 35.100 114.365 35.785 115.005 ;
        RECT 35.955 115.865 36.230 116.565 ;
        RECT 36.440 116.190 36.655 116.735 ;
        RECT 36.825 116.225 37.300 116.565 ;
        RECT 37.470 116.230 38.085 116.735 ;
        RECT 37.470 116.055 37.665 116.230 ;
        RECT 35.955 114.835 36.125 115.865 ;
        RECT 36.400 115.695 37.115 115.990 ;
        RECT 37.335 115.865 37.665 116.055 ;
        RECT 37.835 115.695 38.085 116.060 ;
        RECT 36.295 115.525 38.085 115.695 ;
        RECT 36.295 115.095 36.525 115.525 ;
        RECT 35.955 114.355 36.215 114.835 ;
        RECT 36.695 114.825 37.105 115.345 ;
        RECT 36.385 114.185 36.715 114.645 ;
        RECT 36.905 114.405 37.105 114.825 ;
        RECT 37.275 114.670 37.530 115.525 ;
        RECT 38.325 115.345 38.495 116.565 ;
        RECT 38.745 116.225 39.005 116.735 ;
        RECT 37.700 115.095 38.495 115.345 ;
        RECT 38.665 115.175 39.005 116.055 ;
        RECT 39.175 115.645 40.385 116.735 ;
        RECT 38.245 115.005 38.495 115.095 ;
        RECT 37.275 114.405 38.065 114.670 ;
        RECT 38.245 114.585 38.575 115.005 ;
        RECT 38.745 114.185 39.005 115.005 ;
        RECT 39.175 114.935 39.695 115.475 ;
        RECT 39.865 115.105 40.385 115.645 ;
        RECT 40.645 115.725 40.815 116.565 ;
        RECT 40.985 116.395 42.155 116.565 ;
        RECT 40.985 115.895 41.315 116.395 ;
        RECT 41.825 116.355 42.155 116.395 ;
        RECT 42.345 116.315 42.700 116.735 ;
        RECT 41.485 116.135 41.715 116.225 ;
        RECT 42.870 116.135 43.120 116.565 ;
        RECT 41.485 115.895 43.120 116.135 ;
        RECT 43.290 115.975 43.620 116.735 ;
        RECT 43.790 115.895 44.045 116.565 ;
        RECT 40.645 115.555 43.705 115.725 ;
        RECT 40.560 115.175 40.910 115.385 ;
        RECT 41.080 115.175 41.525 115.375 ;
        RECT 41.695 115.175 42.170 115.375 ;
        RECT 39.175 114.185 40.385 114.935 ;
        RECT 40.645 114.835 41.710 115.005 ;
        RECT 40.645 114.355 40.815 114.835 ;
        RECT 40.985 114.185 41.315 114.665 ;
        RECT 41.540 114.605 41.710 114.835 ;
        RECT 41.890 114.775 42.170 115.175 ;
        RECT 42.440 115.175 42.770 115.375 ;
        RECT 42.940 115.205 43.315 115.375 ;
        RECT 42.940 115.175 43.305 115.205 ;
        RECT 42.440 114.775 42.725 115.175 ;
        RECT 43.535 115.005 43.705 115.555 ;
        RECT 42.905 114.835 43.705 115.005 ;
        RECT 42.905 114.605 43.075 114.835 ;
        RECT 43.875 114.765 44.045 115.895 ;
        RECT 43.860 114.695 44.045 114.765 ;
        RECT 43.835 114.685 44.045 114.695 ;
        RECT 41.540 114.355 43.075 114.605 ;
        RECT 43.245 114.185 43.575 114.665 ;
        RECT 43.790 114.355 44.045 114.685 ;
        RECT 45.155 115.865 45.430 116.565 ;
        RECT 45.640 116.190 45.855 116.735 ;
        RECT 46.025 116.225 46.500 116.565 ;
        RECT 46.670 116.230 47.285 116.735 ;
        RECT 46.670 116.055 46.865 116.230 ;
        RECT 45.155 114.835 45.325 115.865 ;
        RECT 45.600 115.695 46.315 115.990 ;
        RECT 46.535 115.865 46.865 116.055 ;
        RECT 47.035 115.695 47.285 116.060 ;
        RECT 45.495 115.525 47.285 115.695 ;
        RECT 45.495 115.095 45.725 115.525 ;
        RECT 45.155 114.355 45.415 114.835 ;
        RECT 45.895 114.825 46.305 115.345 ;
        RECT 45.585 114.185 45.915 114.645 ;
        RECT 46.105 114.405 46.305 114.825 ;
        RECT 46.475 114.670 46.730 115.525 ;
        RECT 47.525 115.345 47.695 116.565 ;
        RECT 47.945 116.225 48.205 116.735 ;
        RECT 48.490 116.105 48.775 116.565 ;
        RECT 48.945 116.275 49.215 116.735 ;
        RECT 46.900 115.095 47.695 115.345 ;
        RECT 47.865 115.175 48.205 116.055 ;
        RECT 48.490 115.885 49.445 116.105 ;
        RECT 48.375 115.155 49.065 115.715 ;
        RECT 47.445 115.005 47.695 115.095 ;
        RECT 46.475 114.405 47.265 114.670 ;
        RECT 47.445 114.585 47.775 115.005 ;
        RECT 47.945 114.185 48.205 115.005 ;
        RECT 49.235 114.985 49.445 115.885 ;
        RECT 48.490 114.815 49.445 114.985 ;
        RECT 49.615 115.715 50.015 116.565 ;
        RECT 50.205 116.105 50.485 116.565 ;
        RECT 51.005 116.275 51.330 116.735 ;
        RECT 50.205 115.885 51.330 116.105 ;
        RECT 49.615 115.155 50.710 115.715 ;
        RECT 50.880 115.425 51.330 115.885 ;
        RECT 51.500 115.595 51.885 116.565 ;
        RECT 48.490 114.355 48.775 114.815 ;
        RECT 48.945 114.185 49.215 114.645 ;
        RECT 49.615 114.355 50.015 115.155 ;
        RECT 50.880 115.095 51.435 115.425 ;
        RECT 50.880 114.985 51.330 115.095 ;
        RECT 50.205 114.815 51.330 114.985 ;
        RECT 51.605 114.925 51.885 115.595 ;
        RECT 52.055 115.570 52.345 116.735 ;
        RECT 52.575 115.675 52.905 116.520 ;
        RECT 53.075 115.725 53.245 116.735 ;
        RECT 53.415 116.005 53.755 116.565 ;
        RECT 53.985 116.235 54.300 116.735 ;
        RECT 54.480 116.265 55.365 116.435 ;
        RECT 52.515 115.595 52.905 115.675 ;
        RECT 53.415 115.630 54.310 116.005 ;
        RECT 50.205 114.355 50.485 114.815 ;
        RECT 51.005 114.185 51.330 114.645 ;
        RECT 51.500 114.355 51.885 114.925 ;
        RECT 52.515 115.545 52.730 115.595 ;
        RECT 52.515 114.965 52.685 115.545 ;
        RECT 53.415 115.425 53.605 115.630 ;
        RECT 54.480 115.425 54.650 116.265 ;
        RECT 55.590 116.235 55.840 116.565 ;
        RECT 52.855 115.095 53.605 115.425 ;
        RECT 53.775 115.095 54.650 115.425 ;
        RECT 52.515 114.925 52.740 114.965 ;
        RECT 53.405 114.925 53.605 115.095 ;
        RECT 52.055 114.185 52.345 114.910 ;
        RECT 52.515 114.840 52.895 114.925 ;
        RECT 52.565 114.405 52.895 114.840 ;
        RECT 53.065 114.185 53.235 114.795 ;
        RECT 53.405 114.400 53.735 114.925 ;
        RECT 53.995 114.185 54.205 114.715 ;
        RECT 54.480 114.635 54.650 115.095 ;
        RECT 54.820 115.135 55.140 116.095 ;
        RECT 55.310 115.345 55.500 116.065 ;
        RECT 55.670 115.165 55.840 116.235 ;
        RECT 56.010 115.935 56.180 116.735 ;
        RECT 56.350 116.290 57.455 116.460 ;
        RECT 56.350 115.675 56.520 116.290 ;
        RECT 57.665 116.140 57.915 116.565 ;
        RECT 58.085 116.275 58.350 116.735 ;
        RECT 56.690 115.755 57.220 116.120 ;
        RECT 57.665 116.010 57.970 116.140 ;
        RECT 56.010 115.585 56.520 115.675 ;
        RECT 56.010 115.415 56.880 115.585 ;
        RECT 56.010 115.345 56.180 115.415 ;
        RECT 56.300 115.165 56.500 115.195 ;
        RECT 54.820 114.805 55.285 115.135 ;
        RECT 55.670 114.865 56.500 115.165 ;
        RECT 55.670 114.635 55.840 114.865 ;
        RECT 54.480 114.465 55.265 114.635 ;
        RECT 55.435 114.465 55.840 114.635 ;
        RECT 56.020 114.185 56.390 114.685 ;
        RECT 56.710 114.635 56.880 115.415 ;
        RECT 57.050 115.055 57.220 115.755 ;
        RECT 57.390 115.225 57.630 115.820 ;
        RECT 57.050 114.835 57.575 115.055 ;
        RECT 57.800 114.905 57.970 116.010 ;
        RECT 57.745 114.775 57.970 114.905 ;
        RECT 58.140 114.815 58.420 115.765 ;
        RECT 57.745 114.635 57.915 114.775 ;
        RECT 56.710 114.465 57.385 114.635 ;
        RECT 57.580 114.465 57.915 114.635 ;
        RECT 58.085 114.185 58.335 114.645 ;
        RECT 58.590 114.445 58.775 116.565 ;
        RECT 58.945 116.235 59.275 116.735 ;
        RECT 59.445 116.065 59.615 116.565 ;
        RECT 58.950 115.895 59.615 116.065 ;
        RECT 58.950 114.905 59.180 115.895 ;
        RECT 59.350 115.075 59.700 115.725 ;
        RECT 59.875 115.645 61.085 116.735 ;
        RECT 59.875 114.935 60.395 115.475 ;
        RECT 60.565 115.105 61.085 115.645 ;
        RECT 61.255 115.130 61.535 116.565 ;
        RECT 61.705 115.960 62.415 116.735 ;
        RECT 62.585 115.790 62.915 116.565 ;
        RECT 61.765 115.575 62.915 115.790 ;
        RECT 58.950 114.735 59.615 114.905 ;
        RECT 58.945 114.185 59.275 114.565 ;
        RECT 59.445 114.445 59.615 114.735 ;
        RECT 59.875 114.185 61.085 114.935 ;
        RECT 61.255 114.355 61.595 115.130 ;
        RECT 61.765 115.005 62.050 115.575 ;
        RECT 62.235 115.175 62.705 115.405 ;
        RECT 63.110 115.375 63.325 116.490 ;
        RECT 63.505 116.015 63.835 116.735 ;
        RECT 63.615 115.375 63.845 115.715 ;
        RECT 64.015 115.645 65.225 116.735 ;
        RECT 62.875 115.195 63.325 115.375 ;
        RECT 62.875 115.175 63.205 115.195 ;
        RECT 63.515 115.175 63.845 115.375 ;
        RECT 61.765 114.815 62.475 115.005 ;
        RECT 62.175 114.675 62.475 114.815 ;
        RECT 62.665 114.815 63.845 115.005 ;
        RECT 62.665 114.735 62.995 114.815 ;
        RECT 62.175 114.665 62.490 114.675 ;
        RECT 62.175 114.655 62.500 114.665 ;
        RECT 62.175 114.650 62.510 114.655 ;
        RECT 61.765 114.185 61.935 114.645 ;
        RECT 62.175 114.640 62.515 114.650 ;
        RECT 62.175 114.635 62.520 114.640 ;
        RECT 62.175 114.625 62.525 114.635 ;
        RECT 62.175 114.620 62.530 114.625 ;
        RECT 62.175 114.355 62.535 114.620 ;
        RECT 63.165 114.185 63.335 114.645 ;
        RECT 63.505 114.355 63.845 114.815 ;
        RECT 64.015 114.935 64.535 115.475 ;
        RECT 64.705 115.105 65.225 115.645 ;
        RECT 65.400 115.595 65.675 116.565 ;
        RECT 65.885 115.935 66.165 116.735 ;
        RECT 66.335 116.225 67.525 116.515 ;
        RECT 66.335 115.885 67.505 116.055 ;
        RECT 66.335 115.765 66.505 115.885 ;
        RECT 65.845 115.595 66.505 115.765 ;
        RECT 64.015 114.185 65.225 114.935 ;
        RECT 65.400 114.860 65.570 115.595 ;
        RECT 65.845 115.425 66.015 115.595 ;
        RECT 66.815 115.425 67.010 115.715 ;
        RECT 67.180 115.595 67.505 115.885 ;
        RECT 67.695 115.865 67.970 116.565 ;
        RECT 68.140 116.190 68.395 116.735 ;
        RECT 68.565 116.225 69.045 116.565 ;
        RECT 69.220 116.180 69.825 116.735 ;
        RECT 69.210 116.080 69.825 116.180 ;
        RECT 69.210 116.055 69.395 116.080 ;
        RECT 65.740 115.095 66.015 115.425 ;
        RECT 66.185 115.095 67.010 115.425 ;
        RECT 67.180 115.095 67.525 115.425 ;
        RECT 65.845 114.925 66.015 115.095 ;
        RECT 65.400 114.515 65.675 114.860 ;
        RECT 65.845 114.755 67.510 114.925 ;
        RECT 65.865 114.185 66.245 114.585 ;
        RECT 66.415 114.405 66.585 114.755 ;
        RECT 66.755 114.185 67.085 114.585 ;
        RECT 67.255 114.405 67.510 114.755 ;
        RECT 67.695 114.835 67.865 115.865 ;
        RECT 68.140 115.735 68.895 115.985 ;
        RECT 69.065 115.810 69.395 116.055 ;
        RECT 68.140 115.700 68.910 115.735 ;
        RECT 68.140 115.690 68.925 115.700 ;
        RECT 68.035 115.675 68.930 115.690 ;
        RECT 68.035 115.660 68.950 115.675 ;
        RECT 68.035 115.650 68.970 115.660 ;
        RECT 68.035 115.640 68.995 115.650 ;
        RECT 68.035 115.610 69.065 115.640 ;
        RECT 68.035 115.580 69.085 115.610 ;
        RECT 68.035 115.550 69.105 115.580 ;
        RECT 68.035 115.525 69.135 115.550 ;
        RECT 68.035 115.490 69.170 115.525 ;
        RECT 68.035 115.485 69.200 115.490 ;
        RECT 68.035 115.090 68.265 115.485 ;
        RECT 68.810 115.480 69.200 115.485 ;
        RECT 68.835 115.470 69.200 115.480 ;
        RECT 68.850 115.465 69.200 115.470 ;
        RECT 68.865 115.460 69.200 115.465 ;
        RECT 69.565 115.460 69.825 115.910 ;
        RECT 68.865 115.455 69.825 115.460 ;
        RECT 68.875 115.445 69.825 115.455 ;
        RECT 68.885 115.440 69.825 115.445 ;
        RECT 68.895 115.430 69.825 115.440 ;
        RECT 68.900 115.420 69.825 115.430 ;
        RECT 68.905 115.415 69.825 115.420 ;
        RECT 68.915 115.400 69.825 115.415 ;
        RECT 68.920 115.385 69.825 115.400 ;
        RECT 68.930 115.360 69.825 115.385 ;
        RECT 68.435 114.890 68.765 115.315 ;
        RECT 68.515 114.865 68.765 114.890 ;
        RECT 67.695 114.355 67.955 114.835 ;
        RECT 68.125 114.185 68.375 114.725 ;
        RECT 68.545 114.405 68.765 114.865 ;
        RECT 68.935 115.290 69.825 115.360 ;
        RECT 69.995 115.595 70.380 116.565 ;
        RECT 70.550 116.275 70.875 116.735 ;
        RECT 71.395 116.105 71.675 116.565 ;
        RECT 70.550 115.885 71.675 116.105 ;
        RECT 68.935 114.565 69.105 115.290 ;
        RECT 69.275 114.735 69.825 115.120 ;
        RECT 69.995 114.925 70.275 115.595 ;
        RECT 70.550 115.425 71.000 115.885 ;
        RECT 71.865 115.715 72.265 116.565 ;
        RECT 72.665 116.275 72.935 116.735 ;
        RECT 73.105 116.105 73.390 116.565 ;
        RECT 70.445 115.095 71.000 115.425 ;
        RECT 71.170 115.155 72.265 115.715 ;
        RECT 70.550 114.985 71.000 115.095 ;
        RECT 68.935 114.395 69.825 114.565 ;
        RECT 69.995 114.355 70.380 114.925 ;
        RECT 70.550 114.815 71.675 114.985 ;
        RECT 70.550 114.185 70.875 114.645 ;
        RECT 71.395 114.355 71.675 114.815 ;
        RECT 71.865 114.355 72.265 115.155 ;
        RECT 72.435 115.885 73.390 116.105 ;
        RECT 73.675 115.975 74.190 116.385 ;
        RECT 74.425 115.975 74.595 116.735 ;
        RECT 74.765 116.395 76.795 116.565 ;
        RECT 72.435 114.985 72.645 115.885 ;
        RECT 72.815 115.155 73.505 115.715 ;
        RECT 73.675 115.165 74.015 115.975 ;
        RECT 74.765 115.730 74.935 116.395 ;
        RECT 75.330 116.055 76.455 116.225 ;
        RECT 74.185 115.540 74.935 115.730 ;
        RECT 75.105 115.715 76.115 115.885 ;
        RECT 73.675 114.995 74.905 115.165 ;
        RECT 72.435 114.815 73.390 114.985 ;
        RECT 72.665 114.185 72.935 114.645 ;
        RECT 73.105 114.355 73.390 114.815 ;
        RECT 73.950 114.390 74.195 114.995 ;
        RECT 74.415 114.185 74.925 114.720 ;
        RECT 75.105 114.355 75.295 115.715 ;
        RECT 75.465 114.695 75.740 115.515 ;
        RECT 75.945 114.915 76.115 115.715 ;
        RECT 76.285 114.925 76.455 116.055 ;
        RECT 76.625 115.425 76.795 116.395 ;
        RECT 76.965 115.595 77.135 116.735 ;
        RECT 77.305 115.595 77.640 116.565 ;
        RECT 76.625 115.095 76.820 115.425 ;
        RECT 77.045 115.095 77.300 115.425 ;
        RECT 77.045 114.925 77.215 115.095 ;
        RECT 77.470 114.925 77.640 115.595 ;
        RECT 77.815 115.570 78.105 116.735 ;
        RECT 78.365 116.065 78.535 116.565 ;
        RECT 78.705 116.235 79.035 116.735 ;
        RECT 78.365 115.895 79.030 116.065 ;
        RECT 78.280 115.075 78.630 115.725 ;
        RECT 76.285 114.755 77.215 114.925 ;
        RECT 76.285 114.720 76.460 114.755 ;
        RECT 75.465 114.525 75.745 114.695 ;
        RECT 75.465 114.355 75.740 114.525 ;
        RECT 75.930 114.355 76.460 114.720 ;
        RECT 76.885 114.185 77.215 114.585 ;
        RECT 77.385 114.355 77.640 114.925 ;
        RECT 77.815 114.185 78.105 114.910 ;
        RECT 78.800 114.905 79.030 115.895 ;
        RECT 78.365 114.735 79.030 114.905 ;
        RECT 78.365 114.445 78.535 114.735 ;
        RECT 78.705 114.185 79.035 114.565 ;
        RECT 79.205 114.445 79.390 116.565 ;
        RECT 79.630 116.275 79.895 116.735 ;
        RECT 80.065 116.140 80.315 116.565 ;
        RECT 80.525 116.290 81.630 116.460 ;
        RECT 80.010 116.010 80.315 116.140 ;
        RECT 79.560 114.815 79.840 115.765 ;
        RECT 80.010 114.905 80.180 116.010 ;
        RECT 80.350 115.225 80.590 115.820 ;
        RECT 80.760 115.755 81.290 116.120 ;
        RECT 80.760 115.055 80.930 115.755 ;
        RECT 81.460 115.675 81.630 116.290 ;
        RECT 81.800 115.935 81.970 116.735 ;
        RECT 82.140 116.235 82.390 116.565 ;
        RECT 82.615 116.265 83.500 116.435 ;
        RECT 81.460 115.585 81.970 115.675 ;
        RECT 80.010 114.775 80.235 114.905 ;
        RECT 80.405 114.835 80.930 115.055 ;
        RECT 81.100 115.415 81.970 115.585 ;
        RECT 79.645 114.185 79.895 114.645 ;
        RECT 80.065 114.635 80.235 114.775 ;
        RECT 81.100 114.635 81.270 115.415 ;
        RECT 81.800 115.345 81.970 115.415 ;
        RECT 81.480 115.165 81.680 115.195 ;
        RECT 82.140 115.165 82.310 116.235 ;
        RECT 82.480 115.345 82.670 116.065 ;
        RECT 81.480 114.865 82.310 115.165 ;
        RECT 82.840 115.135 83.160 116.095 ;
        RECT 80.065 114.465 80.400 114.635 ;
        RECT 80.595 114.465 81.270 114.635 ;
        RECT 81.590 114.185 81.960 114.685 ;
        RECT 82.140 114.635 82.310 114.865 ;
        RECT 82.695 114.805 83.160 115.135 ;
        RECT 83.330 115.425 83.500 116.265 ;
        RECT 83.680 116.235 83.995 116.735 ;
        RECT 84.225 116.005 84.565 116.565 ;
        RECT 83.670 115.630 84.565 116.005 ;
        RECT 84.735 115.725 84.905 116.735 ;
        RECT 84.375 115.425 84.565 115.630 ;
        RECT 85.075 115.675 85.405 116.520 ;
        RECT 85.575 115.820 85.745 116.735 ;
        RECT 86.610 115.865 86.895 116.735 ;
        RECT 87.065 116.105 87.325 116.565 ;
        RECT 87.500 116.275 87.755 116.735 ;
        RECT 87.925 116.105 88.185 116.565 ;
        RECT 87.065 115.935 88.185 116.105 ;
        RECT 88.355 115.935 88.665 116.735 ;
        RECT 87.065 115.685 87.325 115.935 ;
        RECT 88.835 115.765 89.145 116.565 ;
        RECT 85.075 115.595 85.465 115.675 ;
        RECT 85.250 115.545 85.465 115.595 ;
        RECT 83.330 115.095 84.205 115.425 ;
        RECT 84.375 115.095 85.125 115.425 ;
        RECT 83.330 114.635 83.500 115.095 ;
        RECT 84.375 114.925 84.575 115.095 ;
        RECT 85.295 114.965 85.465 115.545 ;
        RECT 85.240 114.925 85.465 114.965 ;
        RECT 82.140 114.465 82.545 114.635 ;
        RECT 82.715 114.465 83.500 114.635 ;
        RECT 83.775 114.185 83.985 114.715 ;
        RECT 84.245 114.400 84.575 114.925 ;
        RECT 85.085 114.840 85.465 114.925 ;
        RECT 86.570 115.515 87.325 115.685 ;
        RECT 88.115 115.595 89.145 115.765 ;
        RECT 89.315 115.645 92.825 116.735 ;
        RECT 92.995 115.645 94.205 116.735 ;
        RECT 94.480 116.275 94.650 116.735 ;
        RECT 94.820 116.105 95.150 116.565 ;
        RECT 86.570 115.005 86.975 115.515 ;
        RECT 88.115 115.345 88.285 115.595 ;
        RECT 87.145 115.175 88.285 115.345 ;
        RECT 84.745 114.185 84.915 114.795 ;
        RECT 85.085 114.405 85.415 114.840 ;
        RECT 86.570 114.835 88.220 115.005 ;
        RECT 88.455 114.855 88.805 115.425 ;
        RECT 85.585 114.185 85.755 114.700 ;
        RECT 86.615 114.185 86.895 114.665 ;
        RECT 87.065 114.445 87.325 114.835 ;
        RECT 87.500 114.185 87.755 114.665 ;
        RECT 87.925 114.445 88.220 114.835 ;
        RECT 88.975 114.685 89.145 115.595 ;
        RECT 88.400 114.185 88.675 114.665 ;
        RECT 88.845 114.355 89.145 114.685 ;
        RECT 89.315 114.955 90.965 115.475 ;
        RECT 91.135 115.125 92.825 115.645 ;
        RECT 89.315 114.185 92.825 114.955 ;
        RECT 92.995 114.935 93.515 115.475 ;
        RECT 93.685 115.105 94.205 115.645 ;
        RECT 94.375 115.935 95.150 116.105 ;
        RECT 95.320 115.935 95.490 116.735 ;
        RECT 92.995 114.185 94.205 114.935 ;
        RECT 94.375 114.925 94.805 115.935 ;
        RECT 96.075 115.765 96.435 115.940 ;
        RECT 94.975 115.595 96.435 115.765 ;
        RECT 96.680 115.765 96.955 116.565 ;
        RECT 97.125 115.935 97.455 116.735 ;
        RECT 97.625 116.395 98.765 116.565 ;
        RECT 97.625 115.765 97.795 116.395 ;
        RECT 94.975 115.095 95.145 115.595 ;
        RECT 94.375 114.755 95.070 114.925 ;
        RECT 95.315 114.865 95.725 115.425 ;
        RECT 94.400 114.185 94.730 114.585 ;
        RECT 94.900 114.485 95.070 114.755 ;
        RECT 95.895 114.695 96.075 115.595 ;
        RECT 96.680 115.555 97.795 115.765 ;
        RECT 97.965 115.765 98.295 116.225 ;
        RECT 98.465 115.935 98.765 116.395 ;
        RECT 97.965 115.545 98.725 115.765 ;
        RECT 99.015 115.595 99.245 116.735 ;
        RECT 99.415 115.585 99.745 116.565 ;
        RECT 99.915 115.595 100.125 116.735 ;
        RECT 101.475 116.065 101.755 116.735 ;
        RECT 101.925 115.845 102.225 116.395 ;
        RECT 102.425 116.015 102.755 116.735 ;
        RECT 102.945 116.015 103.405 116.565 ;
        RECT 96.245 115.035 96.440 115.425 ;
        RECT 96.680 115.175 97.400 115.375 ;
        RECT 97.570 115.175 98.340 115.375 ;
        RECT 96.245 114.865 96.445 115.035 ;
        RECT 98.510 115.005 98.725 115.545 ;
        RECT 98.995 115.175 99.325 115.425 ;
        RECT 95.240 114.185 95.555 114.695 ;
        RECT 95.785 114.355 96.075 114.695 ;
        RECT 96.245 114.185 96.485 114.695 ;
        RECT 96.680 114.185 96.955 115.005 ;
        RECT 97.125 114.835 98.725 115.005 ;
        RECT 97.125 114.825 98.295 114.835 ;
        RECT 97.125 114.355 97.455 114.825 ;
        RECT 97.625 114.185 97.795 114.655 ;
        RECT 97.965 114.355 98.295 114.825 ;
        RECT 98.465 114.185 98.755 114.655 ;
        RECT 99.015 114.185 99.245 115.005 ;
        RECT 99.495 114.985 99.745 115.585 ;
        RECT 101.290 115.425 101.555 115.785 ;
        RECT 101.925 115.675 102.865 115.845 ;
        RECT 102.695 115.425 102.865 115.675 ;
        RECT 101.290 115.175 101.965 115.425 ;
        RECT 102.185 115.175 102.525 115.425 ;
        RECT 102.695 115.095 102.985 115.425 ;
        RECT 102.695 115.005 102.865 115.095 ;
        RECT 99.415 114.355 99.745 114.985 ;
        RECT 99.915 114.185 100.125 115.005 ;
        RECT 101.475 114.815 102.865 115.005 ;
        RECT 101.475 114.455 101.805 114.815 ;
        RECT 103.155 114.645 103.405 116.015 ;
        RECT 103.575 115.570 103.865 116.735 ;
        RECT 104.035 115.595 104.295 116.735 ;
        RECT 104.465 115.765 104.795 116.565 ;
        RECT 104.965 115.935 105.135 116.735 ;
        RECT 105.305 115.765 105.635 116.565 ;
        RECT 105.805 115.935 106.060 116.735 ;
        RECT 104.465 115.595 106.165 115.765 ;
        RECT 106.335 115.645 109.845 116.735 ;
        RECT 110.015 115.645 111.225 116.735 ;
        RECT 111.485 116.065 111.655 116.565 ;
        RECT 111.825 116.235 112.155 116.735 ;
        RECT 111.485 115.895 112.150 116.065 ;
        RECT 104.035 115.175 104.795 115.425 ;
        RECT 104.965 115.175 105.715 115.425 ;
        RECT 105.885 115.005 106.165 115.595 ;
        RECT 102.425 114.185 102.675 114.645 ;
        RECT 102.845 114.355 103.405 114.645 ;
        RECT 103.575 114.185 103.865 114.910 ;
        RECT 104.035 114.815 105.135 114.985 ;
        RECT 104.035 114.355 104.375 114.815 ;
        RECT 104.545 114.185 104.715 114.645 ;
        RECT 104.885 114.565 105.135 114.815 ;
        RECT 105.305 114.755 106.165 115.005 ;
        RECT 106.335 114.955 107.985 115.475 ;
        RECT 108.155 115.125 109.845 115.645 ;
        RECT 105.725 114.565 106.055 114.585 ;
        RECT 104.885 114.355 106.055 114.565 ;
        RECT 106.335 114.185 109.845 114.955 ;
        RECT 110.015 114.935 110.535 115.475 ;
        RECT 110.705 115.105 111.225 115.645 ;
        RECT 111.400 115.075 111.750 115.725 ;
        RECT 110.015 114.185 111.225 114.935 ;
        RECT 111.920 114.905 112.150 115.895 ;
        RECT 111.485 114.735 112.150 114.905 ;
        RECT 111.485 114.445 111.655 114.735 ;
        RECT 111.825 114.185 112.155 114.565 ;
        RECT 112.325 114.445 112.510 116.565 ;
        RECT 112.750 116.275 113.015 116.735 ;
        RECT 113.185 116.140 113.435 116.565 ;
        RECT 113.645 116.290 114.750 116.460 ;
        RECT 113.130 116.010 113.435 116.140 ;
        RECT 112.680 114.815 112.960 115.765 ;
        RECT 113.130 114.905 113.300 116.010 ;
        RECT 113.470 115.225 113.710 115.820 ;
        RECT 113.880 115.755 114.410 116.120 ;
        RECT 113.880 115.055 114.050 115.755 ;
        RECT 114.580 115.675 114.750 116.290 ;
        RECT 114.920 115.935 115.090 116.735 ;
        RECT 115.260 116.235 115.510 116.565 ;
        RECT 115.735 116.265 116.620 116.435 ;
        RECT 114.580 115.585 115.090 115.675 ;
        RECT 113.130 114.775 113.355 114.905 ;
        RECT 113.525 114.835 114.050 115.055 ;
        RECT 114.220 115.415 115.090 115.585 ;
        RECT 112.765 114.185 113.015 114.645 ;
        RECT 113.185 114.635 113.355 114.775 ;
        RECT 114.220 114.635 114.390 115.415 ;
        RECT 114.920 115.345 115.090 115.415 ;
        RECT 114.600 115.165 114.800 115.195 ;
        RECT 115.260 115.165 115.430 116.235 ;
        RECT 115.600 115.345 115.790 116.065 ;
        RECT 114.600 114.865 115.430 115.165 ;
        RECT 115.960 115.135 116.280 116.095 ;
        RECT 113.185 114.465 113.520 114.635 ;
        RECT 113.715 114.465 114.390 114.635 ;
        RECT 114.710 114.185 115.080 114.685 ;
        RECT 115.260 114.635 115.430 114.865 ;
        RECT 115.815 114.805 116.280 115.135 ;
        RECT 116.450 115.425 116.620 116.265 ;
        RECT 116.800 116.235 117.115 116.735 ;
        RECT 117.345 116.005 117.685 116.565 ;
        RECT 116.790 115.630 117.685 116.005 ;
        RECT 117.855 115.725 118.025 116.735 ;
        RECT 117.495 115.425 117.685 115.630 ;
        RECT 118.195 115.675 118.525 116.520 ;
        RECT 118.195 115.595 118.585 115.675 ;
        RECT 118.765 115.625 119.060 116.735 ;
        RECT 118.370 115.545 118.585 115.595 ;
        RECT 116.450 115.095 117.325 115.425 ;
        RECT 117.495 115.095 118.245 115.425 ;
        RECT 116.450 114.635 116.620 115.095 ;
        RECT 117.495 114.925 117.695 115.095 ;
        RECT 118.415 114.965 118.585 115.545 ;
        RECT 119.240 115.425 119.490 116.560 ;
        RECT 119.660 115.625 119.920 116.735 ;
        RECT 120.090 115.835 120.350 116.560 ;
        RECT 120.520 116.005 120.780 116.735 ;
        RECT 120.950 115.835 121.210 116.560 ;
        RECT 121.380 116.005 121.640 116.735 ;
        RECT 121.810 115.835 122.070 116.560 ;
        RECT 122.240 116.005 122.500 116.735 ;
        RECT 122.670 115.835 122.930 116.560 ;
        RECT 123.100 116.005 123.395 116.735 ;
        RECT 120.090 115.595 123.400 115.835 ;
        RECT 124.020 115.765 124.350 116.565 ;
        RECT 124.520 115.935 124.850 116.735 ;
        RECT 125.150 115.765 125.480 116.565 ;
        RECT 126.125 115.935 126.375 116.735 ;
        RECT 124.020 115.595 126.455 115.765 ;
        RECT 126.645 115.595 126.815 116.735 ;
        RECT 126.985 115.595 127.325 116.565 ;
        RECT 127.495 115.645 129.165 116.735 ;
        RECT 118.360 114.925 118.585 114.965 ;
        RECT 115.260 114.465 115.665 114.635 ;
        RECT 115.835 114.465 116.620 114.635 ;
        RECT 116.895 114.185 117.105 114.715 ;
        RECT 117.365 114.400 117.695 114.925 ;
        RECT 118.205 114.840 118.585 114.925 ;
        RECT 117.865 114.185 118.035 114.795 ;
        RECT 118.205 114.405 118.535 114.840 ;
        RECT 118.755 114.815 119.070 115.425 ;
        RECT 119.240 115.175 122.260 115.425 ;
        RECT 118.815 114.185 119.060 114.645 ;
        RECT 119.240 114.365 119.490 115.175 ;
        RECT 122.430 115.005 123.400 115.595 ;
        RECT 123.815 115.175 124.165 115.425 ;
        RECT 120.090 114.835 123.400 115.005 ;
        RECT 124.350 114.965 124.520 115.595 ;
        RECT 124.690 115.175 125.020 115.375 ;
        RECT 125.190 115.175 125.520 115.375 ;
        RECT 125.690 115.175 126.110 115.375 ;
        RECT 126.285 115.345 126.455 115.595 ;
        RECT 126.285 115.175 126.980 115.345 ;
        RECT 119.660 114.185 119.920 114.710 ;
        RECT 120.090 114.380 120.350 114.835 ;
        RECT 120.520 114.185 120.780 114.665 ;
        RECT 120.950 114.380 121.210 114.835 ;
        RECT 121.380 114.185 121.640 114.665 ;
        RECT 121.810 114.380 122.070 114.835 ;
        RECT 122.240 114.185 122.500 114.665 ;
        RECT 122.670 114.380 122.930 114.835 ;
        RECT 123.100 114.185 123.400 114.665 ;
        RECT 124.020 114.355 124.520 114.965 ;
        RECT 125.150 114.835 126.375 115.005 ;
        RECT 127.150 114.985 127.325 115.595 ;
        RECT 125.150 114.355 125.480 114.835 ;
        RECT 125.650 114.185 125.875 114.645 ;
        RECT 126.045 114.355 126.375 114.835 ;
        RECT 126.565 114.185 126.815 114.985 ;
        RECT 126.985 114.355 127.325 114.985 ;
        RECT 127.495 114.955 128.245 115.475 ;
        RECT 128.415 115.125 129.165 115.645 ;
        RECT 129.335 115.570 129.625 116.735 ;
        RECT 129.885 116.065 130.055 116.565 ;
        RECT 130.225 116.235 130.555 116.735 ;
        RECT 129.885 115.895 130.550 116.065 ;
        RECT 129.800 115.075 130.150 115.725 ;
        RECT 127.495 114.185 129.165 114.955 ;
        RECT 129.335 114.185 129.625 114.910 ;
        RECT 130.320 114.905 130.550 115.895 ;
        RECT 129.885 114.735 130.550 114.905 ;
        RECT 129.885 114.445 130.055 114.735 ;
        RECT 130.225 114.185 130.555 114.565 ;
        RECT 130.725 114.445 130.910 116.565 ;
        RECT 131.150 116.275 131.415 116.735 ;
        RECT 131.585 116.140 131.835 116.565 ;
        RECT 132.045 116.290 133.150 116.460 ;
        RECT 131.530 116.010 131.835 116.140 ;
        RECT 131.080 114.815 131.360 115.765 ;
        RECT 131.530 114.905 131.700 116.010 ;
        RECT 131.870 115.225 132.110 115.820 ;
        RECT 132.280 115.755 132.810 116.120 ;
        RECT 132.280 115.055 132.450 115.755 ;
        RECT 132.980 115.675 133.150 116.290 ;
        RECT 133.320 115.935 133.490 116.735 ;
        RECT 133.660 116.235 133.910 116.565 ;
        RECT 134.135 116.265 135.020 116.435 ;
        RECT 132.980 115.585 133.490 115.675 ;
        RECT 131.530 114.775 131.755 114.905 ;
        RECT 131.925 114.835 132.450 115.055 ;
        RECT 132.620 115.415 133.490 115.585 ;
        RECT 131.165 114.185 131.415 114.645 ;
        RECT 131.585 114.635 131.755 114.775 ;
        RECT 132.620 114.635 132.790 115.415 ;
        RECT 133.320 115.345 133.490 115.415 ;
        RECT 133.000 115.165 133.200 115.195 ;
        RECT 133.660 115.165 133.830 116.235 ;
        RECT 134.000 115.345 134.190 116.065 ;
        RECT 133.000 114.865 133.830 115.165 ;
        RECT 134.360 115.135 134.680 116.095 ;
        RECT 131.585 114.465 131.920 114.635 ;
        RECT 132.115 114.465 132.790 114.635 ;
        RECT 133.110 114.185 133.480 114.685 ;
        RECT 133.660 114.635 133.830 114.865 ;
        RECT 134.215 114.805 134.680 115.135 ;
        RECT 134.850 115.425 135.020 116.265 ;
        RECT 135.200 116.235 135.515 116.735 ;
        RECT 135.745 116.005 136.085 116.565 ;
        RECT 135.190 115.630 136.085 116.005 ;
        RECT 136.255 115.725 136.425 116.735 ;
        RECT 135.895 115.425 136.085 115.630 ;
        RECT 136.595 115.675 136.925 116.520 ;
        RECT 136.595 115.595 136.985 115.675 ;
        RECT 136.770 115.545 136.985 115.595 ;
        RECT 134.850 115.095 135.725 115.425 ;
        RECT 135.895 115.095 136.645 115.425 ;
        RECT 134.850 114.635 135.020 115.095 ;
        RECT 135.895 114.925 136.095 115.095 ;
        RECT 136.815 114.965 136.985 115.545 ;
        RECT 137.615 115.645 138.825 116.735 ;
        RECT 137.615 115.105 138.135 115.645 ;
        RECT 136.760 114.925 136.985 114.965 ;
        RECT 138.305 114.935 138.825 115.475 ;
        RECT 133.660 114.465 134.065 114.635 ;
        RECT 134.235 114.465 135.020 114.635 ;
        RECT 135.295 114.185 135.505 114.715 ;
        RECT 135.765 114.400 136.095 114.925 ;
        RECT 136.605 114.840 136.985 114.925 ;
        RECT 136.265 114.185 136.435 114.795 ;
        RECT 136.605 114.405 136.935 114.840 ;
        RECT 137.615 114.185 138.825 114.935 ;
        RECT 13.330 114.015 138.910 114.185 ;
        RECT 13.415 113.265 14.625 114.015 ;
        RECT 13.415 112.725 13.935 113.265 ;
        RECT 14.795 113.245 17.385 114.015 ;
        RECT 18.105 113.465 18.275 113.755 ;
        RECT 18.445 113.635 18.775 114.015 ;
        RECT 18.105 113.295 18.770 113.465 ;
        RECT 14.105 112.555 14.625 113.095 ;
        RECT 14.795 112.725 16.005 113.245 ;
        RECT 16.175 112.555 17.385 113.075 ;
        RECT 13.415 111.465 14.625 112.555 ;
        RECT 14.795 111.465 17.385 112.555 ;
        RECT 18.020 112.475 18.370 113.125 ;
        RECT 18.540 112.305 18.770 113.295 ;
        RECT 18.105 112.135 18.770 112.305 ;
        RECT 18.105 111.635 18.275 112.135 ;
        RECT 18.445 111.465 18.775 111.965 ;
        RECT 18.945 111.635 19.130 113.755 ;
        RECT 19.385 113.555 19.635 114.015 ;
        RECT 19.805 113.565 20.140 113.735 ;
        RECT 20.335 113.565 21.010 113.735 ;
        RECT 19.805 113.425 19.975 113.565 ;
        RECT 19.300 112.435 19.580 113.385 ;
        RECT 19.750 113.295 19.975 113.425 ;
        RECT 19.750 112.190 19.920 113.295 ;
        RECT 20.145 113.145 20.670 113.365 ;
        RECT 20.090 112.380 20.330 112.975 ;
        RECT 20.500 112.445 20.670 113.145 ;
        RECT 20.840 112.785 21.010 113.565 ;
        RECT 21.330 113.515 21.700 114.015 ;
        RECT 21.880 113.565 22.285 113.735 ;
        RECT 22.455 113.565 23.240 113.735 ;
        RECT 21.880 113.335 22.050 113.565 ;
        RECT 21.220 113.035 22.050 113.335 ;
        RECT 22.435 113.065 22.900 113.395 ;
        RECT 21.220 113.005 21.420 113.035 ;
        RECT 21.540 112.785 21.710 112.855 ;
        RECT 20.840 112.615 21.710 112.785 ;
        RECT 21.200 112.525 21.710 112.615 ;
        RECT 19.750 112.060 20.055 112.190 ;
        RECT 20.500 112.080 21.030 112.445 ;
        RECT 19.370 111.465 19.635 111.925 ;
        RECT 19.805 111.635 20.055 112.060 ;
        RECT 21.200 111.910 21.370 112.525 ;
        RECT 20.265 111.740 21.370 111.910 ;
        RECT 21.540 111.465 21.710 112.265 ;
        RECT 21.880 111.965 22.050 113.035 ;
        RECT 22.220 112.135 22.410 112.855 ;
        RECT 22.580 112.105 22.900 113.065 ;
        RECT 23.070 113.105 23.240 113.565 ;
        RECT 23.515 113.485 23.725 114.015 ;
        RECT 23.985 113.275 24.315 113.800 ;
        RECT 24.485 113.405 24.655 114.015 ;
        RECT 24.825 113.360 25.155 113.795 ;
        RECT 24.825 113.275 25.205 113.360 ;
        RECT 24.115 113.105 24.315 113.275 ;
        RECT 24.980 113.235 25.205 113.275 ;
        RECT 23.070 112.775 23.945 113.105 ;
        RECT 24.115 112.775 24.865 113.105 ;
        RECT 21.880 111.635 22.130 111.965 ;
        RECT 23.070 111.935 23.240 112.775 ;
        RECT 24.115 112.570 24.305 112.775 ;
        RECT 25.035 112.655 25.205 113.235 ;
        RECT 25.375 113.245 27.045 114.015 ;
        RECT 27.215 113.365 27.475 113.845 ;
        RECT 27.645 113.475 27.895 114.015 ;
        RECT 25.375 112.725 26.125 113.245 ;
        RECT 24.990 112.605 25.205 112.655 ;
        RECT 23.410 112.195 24.305 112.570 ;
        RECT 24.815 112.525 25.205 112.605 ;
        RECT 26.295 112.555 27.045 113.075 ;
        RECT 22.355 111.765 23.240 111.935 ;
        RECT 23.420 111.465 23.735 111.965 ;
        RECT 23.965 111.635 24.305 112.195 ;
        RECT 24.475 111.465 24.645 112.475 ;
        RECT 24.815 111.680 25.145 112.525 ;
        RECT 25.375 111.465 27.045 112.555 ;
        RECT 27.215 112.335 27.385 113.365 ;
        RECT 28.065 113.335 28.285 113.795 ;
        RECT 28.035 113.310 28.285 113.335 ;
        RECT 27.555 112.715 27.785 113.110 ;
        RECT 27.955 112.885 28.285 113.310 ;
        RECT 28.455 113.635 29.345 113.805 ;
        RECT 28.455 112.910 28.625 113.635 ;
        RECT 29.515 113.555 30.075 113.845 ;
        RECT 30.245 113.555 30.495 114.015 ;
        RECT 28.795 113.080 29.345 113.465 ;
        RECT 28.455 112.840 29.345 112.910 ;
        RECT 28.450 112.815 29.345 112.840 ;
        RECT 28.440 112.800 29.345 112.815 ;
        RECT 28.435 112.785 29.345 112.800 ;
        RECT 28.425 112.780 29.345 112.785 ;
        RECT 28.420 112.770 29.345 112.780 ;
        RECT 28.415 112.760 29.345 112.770 ;
        RECT 28.405 112.755 29.345 112.760 ;
        RECT 28.395 112.745 29.345 112.755 ;
        RECT 28.385 112.740 29.345 112.745 ;
        RECT 28.385 112.735 28.720 112.740 ;
        RECT 28.370 112.730 28.720 112.735 ;
        RECT 28.355 112.720 28.720 112.730 ;
        RECT 28.330 112.715 28.720 112.720 ;
        RECT 27.555 112.710 28.720 112.715 ;
        RECT 27.555 112.675 28.690 112.710 ;
        RECT 27.555 112.650 28.655 112.675 ;
        RECT 27.555 112.620 28.625 112.650 ;
        RECT 27.555 112.590 28.605 112.620 ;
        RECT 27.555 112.560 28.585 112.590 ;
        RECT 27.555 112.550 28.515 112.560 ;
        RECT 27.555 112.540 28.490 112.550 ;
        RECT 27.555 112.525 28.470 112.540 ;
        RECT 27.555 112.510 28.450 112.525 ;
        RECT 27.660 112.500 28.445 112.510 ;
        RECT 27.660 112.465 28.430 112.500 ;
        RECT 27.215 111.635 27.490 112.335 ;
        RECT 27.660 112.215 28.415 112.465 ;
        RECT 28.585 112.145 28.915 112.390 ;
        RECT 29.085 112.290 29.345 112.740 ;
        RECT 28.730 112.120 28.915 112.145 ;
        RECT 29.515 112.185 29.765 113.555 ;
        RECT 31.115 113.385 31.445 113.745 ;
        RECT 31.815 113.470 37.160 114.015 ;
        RECT 30.055 113.195 31.445 113.385 ;
        RECT 30.055 113.105 30.225 113.195 ;
        RECT 29.935 112.775 30.225 113.105 ;
        RECT 30.395 112.775 30.735 113.025 ;
        RECT 30.955 112.775 31.630 113.025 ;
        RECT 30.055 112.525 30.225 112.775 ;
        RECT 30.055 112.355 30.995 112.525 ;
        RECT 31.365 112.415 31.630 112.775 ;
        RECT 33.400 112.640 33.740 113.470 ;
        RECT 37.335 113.245 39.005 114.015 ;
        RECT 39.175 113.290 39.465 114.015 ;
        RECT 39.635 113.245 41.305 114.015 ;
        RECT 42.110 113.365 42.440 113.845 ;
        RECT 42.610 113.535 42.860 114.015 ;
        RECT 43.030 113.365 43.360 113.845 ;
        RECT 43.530 113.535 43.780 114.015 ;
        RECT 43.950 113.535 44.280 113.845 ;
        RECT 43.950 113.365 44.120 113.535 ;
        RECT 44.645 113.365 44.985 113.845 ;
        RECT 28.730 112.020 29.345 112.120 ;
        RECT 27.660 111.465 27.915 112.010 ;
        RECT 28.085 111.635 28.565 111.975 ;
        RECT 28.740 111.465 29.345 112.020 ;
        RECT 29.515 111.635 29.975 112.185 ;
        RECT 30.165 111.465 30.495 112.185 ;
        RECT 30.695 111.805 30.995 112.355 ;
        RECT 31.165 111.465 31.445 112.135 ;
        RECT 35.220 111.900 35.570 113.150 ;
        RECT 37.335 112.725 38.085 113.245 ;
        RECT 38.255 112.555 39.005 113.075 ;
        RECT 39.635 112.725 40.385 113.245 ;
        RECT 42.110 113.195 44.120 113.365 ;
        RECT 44.290 113.195 44.985 113.365 ;
        RECT 31.815 111.465 37.160 111.900 ;
        RECT 37.335 111.465 39.005 112.555 ;
        RECT 39.175 111.465 39.465 112.630 ;
        RECT 40.555 112.555 41.305 113.075 ;
        RECT 41.990 112.775 42.570 113.025 ;
        RECT 42.740 112.685 43.070 113.025 ;
        RECT 43.240 112.855 43.570 113.025 ;
        RECT 39.635 111.465 41.305 112.555 ;
        RECT 42.110 111.465 42.440 112.605 ;
        RECT 42.740 111.745 43.080 112.685 ;
        RECT 43.250 111.745 43.570 112.855 ;
        RECT 43.750 112.855 44.080 113.025 ;
        RECT 43.750 111.745 44.055 112.855 ;
        RECT 44.290 112.615 44.460 113.195 ;
        RECT 44.630 112.825 44.965 113.025 ;
        RECT 44.225 111.635 44.555 112.615 ;
        RECT 44.725 111.465 44.985 112.655 ;
        RECT 45.165 111.645 45.425 113.835 ;
        RECT 45.685 113.645 46.355 114.015 ;
        RECT 46.535 113.465 46.845 113.835 ;
        RECT 45.615 113.265 46.845 113.465 ;
        RECT 45.615 112.595 45.905 113.265 ;
        RECT 47.025 113.085 47.255 113.725 ;
        RECT 47.435 113.285 47.725 114.015 ;
        RECT 47.915 113.340 48.190 113.685 ;
        RECT 48.380 113.615 48.760 114.015 ;
        RECT 48.930 113.445 49.100 113.795 ;
        RECT 49.270 113.615 49.600 114.015 ;
        RECT 49.775 113.445 49.945 113.795 ;
        RECT 50.145 113.515 50.475 114.015 ;
        RECT 46.085 112.775 46.550 113.085 ;
        RECT 46.730 112.775 47.255 113.085 ;
        RECT 47.435 112.775 47.735 113.105 ;
        RECT 47.915 112.605 48.085 113.340 ;
        RECT 48.360 113.275 49.945 113.445 ;
        RECT 48.360 113.105 48.530 113.275 ;
        RECT 50.670 113.105 50.915 113.795 ;
        RECT 51.085 113.515 51.425 114.015 ;
        RECT 51.760 113.505 52.000 114.015 ;
        RECT 52.180 113.505 52.460 113.835 ;
        RECT 52.690 113.505 52.905 114.015 ;
        RECT 48.255 112.775 48.530 113.105 ;
        RECT 48.700 112.775 49.080 113.105 ;
        RECT 48.360 112.605 48.530 112.775 ;
        RECT 45.615 112.375 46.385 112.595 ;
        RECT 45.595 111.465 45.935 112.195 ;
        RECT 46.115 111.645 46.385 112.375 ;
        RECT 46.565 112.355 47.725 112.595 ;
        RECT 46.565 111.645 46.795 112.355 ;
        RECT 46.965 111.465 47.295 112.175 ;
        RECT 47.465 111.645 47.725 112.355 ;
        RECT 47.915 111.635 48.190 112.605 ;
        RECT 48.360 112.435 49.020 112.605 ;
        RECT 49.250 112.485 49.990 113.105 ;
        RECT 50.260 112.775 50.915 113.105 ;
        RECT 51.085 112.775 51.425 113.345 ;
        RECT 51.655 112.775 52.010 113.335 ;
        RECT 48.850 112.315 49.020 112.435 ;
        RECT 50.160 112.315 50.480 112.605 ;
        RECT 48.400 111.465 48.680 112.265 ;
        RECT 48.850 112.145 50.480 112.315 ;
        RECT 50.675 112.180 50.915 112.775 ;
        RECT 52.180 112.605 52.350 113.505 ;
        RECT 52.520 112.775 52.785 113.335 ;
        RECT 53.075 113.275 53.690 113.845 ;
        RECT 53.895 113.470 59.240 114.015 ;
        RECT 59.880 113.485 60.170 113.835 ;
        RECT 60.365 113.655 60.695 114.015 ;
        RECT 60.865 113.485 61.095 113.790 ;
        RECT 53.035 112.605 53.205 113.105 ;
        RECT 48.850 111.805 50.905 111.975 ;
        RECT 48.850 111.685 50.900 111.805 ;
        RECT 51.085 111.465 51.425 112.540 ;
        RECT 51.780 112.435 53.205 112.605 ;
        RECT 51.780 112.260 52.170 112.435 ;
        RECT 52.655 111.465 52.985 112.265 ;
        RECT 53.375 112.255 53.690 113.275 ;
        RECT 55.480 112.640 55.820 113.470 ;
        RECT 59.880 113.315 61.095 113.485 ;
        RECT 61.285 113.675 61.455 113.710 ;
        RECT 61.285 113.505 61.485 113.675 ;
        RECT 53.155 111.635 53.690 112.255 ;
        RECT 57.300 111.900 57.650 113.150 ;
        RECT 61.285 113.145 61.455 113.505 ;
        RECT 59.940 112.995 60.200 113.105 ;
        RECT 59.935 112.825 60.200 112.995 ;
        RECT 59.940 112.775 60.200 112.825 ;
        RECT 60.380 112.775 60.765 113.105 ;
        RECT 60.935 112.975 61.455 113.145 ;
        RECT 61.715 113.275 62.180 113.820 ;
        RECT 53.895 111.465 59.240 111.900 ;
        RECT 59.880 111.465 60.200 112.605 ;
        RECT 60.380 111.725 60.575 112.775 ;
        RECT 60.935 112.595 61.105 112.975 ;
        RECT 60.755 112.315 61.105 112.595 ;
        RECT 61.295 112.445 61.540 112.805 ;
        RECT 61.715 112.315 61.885 113.275 ;
        RECT 62.685 113.195 62.855 114.015 ;
        RECT 63.025 113.365 63.355 113.845 ;
        RECT 63.525 113.625 63.875 114.015 ;
        RECT 64.045 113.445 64.275 113.845 ;
        RECT 63.765 113.365 64.275 113.445 ;
        RECT 63.025 113.275 64.275 113.365 ;
        RECT 64.445 113.275 64.765 113.755 ;
        RECT 64.935 113.290 65.225 114.015 ;
        RECT 63.025 113.195 63.935 113.275 ;
        RECT 62.055 112.655 62.300 113.105 ;
        RECT 62.560 112.825 63.255 113.025 ;
        RECT 63.425 112.855 64.025 113.025 ;
        RECT 63.425 112.655 63.595 112.855 ;
        RECT 64.255 112.685 64.425 113.105 ;
        RECT 62.055 112.485 63.595 112.655 ;
        RECT 63.765 112.515 64.425 112.685 ;
        RECT 63.765 112.315 63.935 112.515 ;
        RECT 64.595 112.345 64.765 113.275 ;
        RECT 65.395 113.215 66.090 113.845 ;
        RECT 66.295 113.215 66.605 114.015 ;
        RECT 66.825 113.495 67.080 113.795 ;
        RECT 67.250 113.615 67.580 114.015 ;
        RECT 66.775 113.445 67.080 113.495 ;
        RECT 67.750 113.445 67.920 113.795 ;
        RECT 68.220 113.535 68.390 114.015 ;
        RECT 68.625 113.505 68.975 113.835 ;
        RECT 69.145 113.535 69.315 114.015 ;
        RECT 66.775 113.365 67.920 113.445 ;
        RECT 66.775 113.335 68.485 113.365 ;
        RECT 66.775 113.275 68.635 113.335 ;
        RECT 65.415 112.775 65.750 113.025 ;
        RECT 60.755 111.635 61.085 112.315 ;
        RECT 61.285 111.465 61.540 112.265 ;
        RECT 61.715 112.145 63.935 112.315 ;
        RECT 64.105 112.145 64.765 112.345 ;
        RECT 61.715 111.465 62.015 111.975 ;
        RECT 62.185 111.635 62.515 112.145 ;
        RECT 64.105 111.975 64.275 112.145 ;
        RECT 62.685 111.465 63.315 111.975 ;
        RECT 63.895 111.805 64.275 111.975 ;
        RECT 64.445 111.465 64.745 111.975 ;
        RECT 64.935 111.465 65.225 112.630 ;
        RECT 65.920 112.615 66.090 113.215 ;
        RECT 66.260 112.775 66.595 113.045 ;
        RECT 65.395 111.465 65.655 112.605 ;
        RECT 65.825 111.635 66.155 112.615 ;
        RECT 66.775 112.605 66.945 113.275 ;
        RECT 67.750 113.195 68.635 113.275 ;
        RECT 68.315 113.165 68.635 113.195 ;
        RECT 67.120 112.775 67.420 113.105 ;
        RECT 66.325 111.465 66.605 112.605 ;
        RECT 66.775 112.175 67.080 112.605 ;
        RECT 67.250 112.315 67.420 112.775 ;
        RECT 67.680 112.485 68.215 113.025 ;
        RECT 68.465 112.775 68.635 113.165 ;
        RECT 68.805 112.605 68.975 113.505 ;
        RECT 69.565 113.365 69.825 113.810 ;
        RECT 68.580 112.400 68.975 112.605 ;
        RECT 69.145 113.195 69.825 113.365 ;
        RECT 67.250 112.230 68.360 112.315 ;
        RECT 69.145 112.290 69.315 113.195 ;
        RECT 70.085 113.145 70.255 113.710 ;
        RECT 70.445 113.485 70.675 113.790 ;
        RECT 70.845 113.655 71.175 114.015 ;
        RECT 71.370 113.485 71.660 113.835 ;
        RECT 70.445 113.315 71.660 113.485 ;
        RECT 71.835 113.470 77.180 114.015 ;
        RECT 77.355 113.470 82.700 114.015 ;
        RECT 69.485 112.460 69.825 113.025 ;
        RECT 70.085 112.975 70.605 113.145 ;
        RECT 70.000 112.445 70.245 112.805 ;
        RECT 70.435 112.595 70.605 112.975 ;
        RECT 70.775 112.775 71.160 113.105 ;
        RECT 71.340 112.995 71.600 113.105 ;
        RECT 71.340 112.825 71.605 112.995 ;
        RECT 71.340 112.775 71.600 112.825 ;
        RECT 70.435 112.315 70.785 112.595 ;
        RECT 69.145 112.230 69.825 112.290 ;
        RECT 67.250 112.145 69.825 112.230 ;
        RECT 68.190 112.060 69.825 112.145 ;
        RECT 66.775 111.735 67.975 111.975 ;
        RECT 68.155 111.465 68.485 111.890 ;
        RECT 69.000 111.465 69.360 111.890 ;
        RECT 69.565 111.880 69.825 112.060 ;
        RECT 70.000 111.465 70.255 112.265 ;
        RECT 70.455 111.635 70.785 112.315 ;
        RECT 70.965 111.725 71.160 112.775 ;
        RECT 73.420 112.640 73.760 113.470 ;
        RECT 71.340 111.465 71.660 112.605 ;
        RECT 75.240 111.900 75.590 113.150 ;
        RECT 78.940 112.640 79.280 113.470 ;
        RECT 83.425 113.465 83.595 113.755 ;
        RECT 83.765 113.635 84.095 114.015 ;
        RECT 83.425 113.295 84.090 113.465 ;
        RECT 80.760 111.900 81.110 113.150 ;
        RECT 83.340 112.475 83.690 113.125 ;
        RECT 83.860 112.305 84.090 113.295 ;
        RECT 83.425 112.135 84.090 112.305 ;
        RECT 71.835 111.465 77.180 111.900 ;
        RECT 77.355 111.465 82.700 111.900 ;
        RECT 83.425 111.635 83.595 112.135 ;
        RECT 83.765 111.465 84.095 111.965 ;
        RECT 84.265 111.635 84.450 113.755 ;
        RECT 84.705 113.555 84.955 114.015 ;
        RECT 85.125 113.565 85.460 113.735 ;
        RECT 85.655 113.565 86.330 113.735 ;
        RECT 85.125 113.425 85.295 113.565 ;
        RECT 84.620 112.435 84.900 113.385 ;
        RECT 85.070 113.295 85.295 113.425 ;
        RECT 85.070 112.190 85.240 113.295 ;
        RECT 85.465 113.145 85.990 113.365 ;
        RECT 85.410 112.380 85.650 112.975 ;
        RECT 85.820 112.445 85.990 113.145 ;
        RECT 86.160 112.785 86.330 113.565 ;
        RECT 86.650 113.515 87.020 114.015 ;
        RECT 87.200 113.565 87.605 113.735 ;
        RECT 87.775 113.565 88.560 113.735 ;
        RECT 87.200 113.335 87.370 113.565 ;
        RECT 86.540 113.035 87.370 113.335 ;
        RECT 87.755 113.065 88.220 113.395 ;
        RECT 86.540 113.005 86.740 113.035 ;
        RECT 86.860 112.785 87.030 112.855 ;
        RECT 86.160 112.615 87.030 112.785 ;
        RECT 86.520 112.525 87.030 112.615 ;
        RECT 85.070 112.060 85.375 112.190 ;
        RECT 85.820 112.080 86.350 112.445 ;
        RECT 84.690 111.465 84.955 111.925 ;
        RECT 85.125 111.635 85.375 112.060 ;
        RECT 86.520 111.910 86.690 112.525 ;
        RECT 85.585 111.740 86.690 111.910 ;
        RECT 86.860 111.465 87.030 112.265 ;
        RECT 87.200 111.965 87.370 113.035 ;
        RECT 87.540 112.135 87.730 112.855 ;
        RECT 87.900 112.105 88.220 113.065 ;
        RECT 88.390 113.105 88.560 113.565 ;
        RECT 88.835 113.485 89.045 114.015 ;
        RECT 89.305 113.275 89.635 113.800 ;
        RECT 89.805 113.405 89.975 114.015 ;
        RECT 90.145 113.360 90.475 113.795 ;
        RECT 90.145 113.275 90.525 113.360 ;
        RECT 90.695 113.290 90.985 114.015 ;
        RECT 89.435 113.105 89.635 113.275 ;
        RECT 90.300 113.235 90.525 113.275 ;
        RECT 88.390 112.775 89.265 113.105 ;
        RECT 89.435 112.775 90.185 113.105 ;
        RECT 87.200 111.635 87.450 111.965 ;
        RECT 88.390 111.935 88.560 112.775 ;
        RECT 89.435 112.570 89.625 112.775 ;
        RECT 90.355 112.655 90.525 113.235 ;
        RECT 90.310 112.605 90.525 112.655 ;
        RECT 88.730 112.195 89.625 112.570 ;
        RECT 90.135 112.525 90.525 112.605 ;
        RECT 87.675 111.765 88.560 111.935 ;
        RECT 88.740 111.465 89.055 111.965 ;
        RECT 89.285 111.635 89.625 112.195 ;
        RECT 89.795 111.465 89.965 112.475 ;
        RECT 90.135 111.680 90.465 112.525 ;
        RECT 90.695 111.465 90.985 112.630 ;
        RECT 91.160 112.415 91.495 113.835 ;
        RECT 91.675 113.645 92.420 114.015 ;
        RECT 92.985 113.475 93.240 113.835 ;
        RECT 93.420 113.645 93.750 114.015 ;
        RECT 93.930 113.475 94.155 113.835 ;
        RECT 91.670 113.285 94.155 113.475 ;
        RECT 94.375 113.470 99.720 114.015 ;
        RECT 91.670 112.595 91.895 113.285 ;
        RECT 92.095 112.775 92.375 113.105 ;
        RECT 92.555 112.775 93.130 113.105 ;
        RECT 93.310 112.775 93.745 113.105 ;
        RECT 93.925 112.775 94.195 113.105 ;
        RECT 95.960 112.640 96.300 113.470 ;
        RECT 99.895 113.245 101.565 114.015 ;
        RECT 91.670 112.415 94.165 112.595 ;
        RECT 91.160 111.645 91.425 112.415 ;
        RECT 91.595 111.465 91.925 112.185 ;
        RECT 92.115 112.005 93.305 112.235 ;
        RECT 92.115 111.645 92.375 112.005 ;
        RECT 92.545 111.465 92.875 111.835 ;
        RECT 93.045 111.645 93.305 112.005 ;
        RECT 93.875 111.645 94.165 112.415 ;
        RECT 97.780 111.900 98.130 113.150 ;
        RECT 99.895 112.725 100.645 113.245 ;
        RECT 102.195 113.215 102.535 113.845 ;
        RECT 102.705 113.215 102.955 114.015 ;
        RECT 103.145 113.365 103.475 113.845 ;
        RECT 103.645 113.555 103.870 114.015 ;
        RECT 104.040 113.365 104.370 113.845 ;
        RECT 100.815 112.555 101.565 113.075 ;
        RECT 94.375 111.465 99.720 111.900 ;
        RECT 99.895 111.465 101.565 112.555 ;
        RECT 102.195 112.605 102.370 113.215 ;
        RECT 103.145 113.195 104.370 113.365 ;
        RECT 105.000 113.235 105.500 113.845 ;
        RECT 105.910 113.275 106.525 113.845 ;
        RECT 106.695 113.505 106.910 114.015 ;
        RECT 107.140 113.505 107.420 113.835 ;
        RECT 107.600 113.505 107.840 114.015 ;
        RECT 102.540 112.855 103.235 113.025 ;
        RECT 103.065 112.605 103.235 112.855 ;
        RECT 103.410 112.825 103.830 113.025 ;
        RECT 104.000 112.825 104.330 113.025 ;
        RECT 104.500 112.825 104.830 113.025 ;
        RECT 105.000 112.605 105.170 113.235 ;
        RECT 105.355 112.775 105.705 113.025 ;
        RECT 102.195 111.635 102.535 112.605 ;
        RECT 102.705 111.465 102.875 112.605 ;
        RECT 103.065 112.435 105.500 112.605 ;
        RECT 103.145 111.465 103.395 112.265 ;
        RECT 104.040 111.635 104.370 112.435 ;
        RECT 104.670 111.465 105.000 112.265 ;
        RECT 105.170 111.635 105.500 112.435 ;
        RECT 105.910 112.255 106.225 113.275 ;
        RECT 106.395 112.605 106.565 113.105 ;
        RECT 106.815 112.775 107.080 113.335 ;
        RECT 107.250 112.605 107.420 113.505 ;
        RECT 107.590 112.775 107.945 113.335 ;
        RECT 108.175 113.265 109.385 114.015 ;
        RECT 109.720 113.505 109.960 114.015 ;
        RECT 110.140 113.505 110.420 113.835 ;
        RECT 110.650 113.505 110.865 114.015 ;
        RECT 108.175 112.725 108.695 113.265 ;
        RECT 106.395 112.435 107.820 112.605 ;
        RECT 108.865 112.555 109.385 113.095 ;
        RECT 109.615 112.775 109.970 113.335 ;
        RECT 110.140 112.605 110.310 113.505 ;
        RECT 110.480 112.775 110.745 113.335 ;
        RECT 111.035 113.275 111.650 113.845 ;
        RECT 110.995 112.605 111.165 113.105 ;
        RECT 105.910 111.635 106.445 112.255 ;
        RECT 106.615 111.465 106.945 112.265 ;
        RECT 107.430 112.260 107.820 112.435 ;
        RECT 108.175 111.465 109.385 112.555 ;
        RECT 109.740 112.435 111.165 112.605 ;
        RECT 109.740 112.260 110.130 112.435 ;
        RECT 110.615 111.465 110.945 112.265 ;
        RECT 111.335 112.255 111.650 113.275 ;
        RECT 111.115 111.635 111.650 112.255 ;
        RECT 111.855 113.215 112.195 113.845 ;
        RECT 112.365 113.215 112.615 114.015 ;
        RECT 112.805 113.365 113.135 113.845 ;
        RECT 113.305 113.555 113.530 114.015 ;
        RECT 113.700 113.365 114.030 113.845 ;
        RECT 111.855 112.605 112.030 113.215 ;
        RECT 112.805 113.195 114.030 113.365 ;
        RECT 114.660 113.235 115.160 113.845 ;
        RECT 116.455 113.290 116.745 114.015 ;
        RECT 116.975 113.555 117.220 114.015 ;
        RECT 112.200 112.855 112.895 113.025 ;
        RECT 112.725 112.605 112.895 112.855 ;
        RECT 113.070 112.825 113.490 113.025 ;
        RECT 113.660 112.825 113.990 113.025 ;
        RECT 114.160 112.825 114.490 113.025 ;
        RECT 114.660 112.605 114.830 113.235 ;
        RECT 115.015 112.775 115.365 113.025 ;
        RECT 116.915 112.775 117.230 113.385 ;
        RECT 117.400 113.025 117.650 113.835 ;
        RECT 117.820 113.490 118.080 114.015 ;
        RECT 118.250 113.365 118.510 113.820 ;
        RECT 118.680 113.535 118.940 114.015 ;
        RECT 119.110 113.365 119.370 113.820 ;
        RECT 119.540 113.535 119.800 114.015 ;
        RECT 119.970 113.365 120.230 113.820 ;
        RECT 120.400 113.535 120.660 114.015 ;
        RECT 120.830 113.365 121.090 113.820 ;
        RECT 121.260 113.535 121.560 114.015 ;
        RECT 118.250 113.195 121.560 113.365 ;
        RECT 117.400 112.775 120.420 113.025 ;
        RECT 111.855 111.635 112.195 112.605 ;
        RECT 112.365 111.465 112.535 112.605 ;
        RECT 112.725 112.435 115.160 112.605 ;
        RECT 112.805 111.465 113.055 112.265 ;
        RECT 113.700 111.635 114.030 112.435 ;
        RECT 114.330 111.465 114.660 112.265 ;
        RECT 114.830 111.635 115.160 112.435 ;
        RECT 116.455 111.465 116.745 112.630 ;
        RECT 116.925 111.465 117.220 112.575 ;
        RECT 117.400 111.640 117.650 112.775 ;
        RECT 120.590 112.605 121.560 113.195 ;
        RECT 121.975 113.245 123.645 114.015 ;
        RECT 121.975 112.725 122.725 113.245 ;
        RECT 124.020 113.235 124.520 113.845 ;
        RECT 117.820 111.465 118.080 112.575 ;
        RECT 118.250 112.365 121.560 112.605 ;
        RECT 122.895 112.555 123.645 113.075 ;
        RECT 123.815 112.775 124.165 113.025 ;
        RECT 124.350 112.605 124.520 113.235 ;
        RECT 125.150 113.365 125.480 113.845 ;
        RECT 125.650 113.555 125.875 114.015 ;
        RECT 126.045 113.365 126.375 113.845 ;
        RECT 125.150 113.195 126.375 113.365 ;
        RECT 126.565 113.215 126.815 114.015 ;
        RECT 126.985 113.215 127.325 113.845 ;
        RECT 127.585 113.465 127.755 113.755 ;
        RECT 127.925 113.635 128.255 114.015 ;
        RECT 127.585 113.295 128.250 113.465 ;
        RECT 124.690 112.825 125.020 113.025 ;
        RECT 125.190 112.825 125.520 113.025 ;
        RECT 125.690 112.825 126.110 113.025 ;
        RECT 126.285 112.855 126.980 113.025 ;
        RECT 126.285 112.605 126.455 112.855 ;
        RECT 127.150 112.655 127.325 113.215 ;
        RECT 127.095 112.605 127.325 112.655 ;
        RECT 118.250 111.640 118.510 112.365 ;
        RECT 118.680 111.465 118.940 112.195 ;
        RECT 119.110 111.640 119.370 112.365 ;
        RECT 119.540 111.465 119.800 112.195 ;
        RECT 119.970 111.640 120.230 112.365 ;
        RECT 120.400 111.465 120.660 112.195 ;
        RECT 120.830 111.640 121.090 112.365 ;
        RECT 121.260 111.465 121.555 112.195 ;
        RECT 121.975 111.465 123.645 112.555 ;
        RECT 124.020 112.435 126.455 112.605 ;
        RECT 124.020 111.635 124.350 112.435 ;
        RECT 124.520 111.465 124.850 112.265 ;
        RECT 125.150 111.635 125.480 112.435 ;
        RECT 126.125 111.465 126.375 112.265 ;
        RECT 126.645 111.465 126.815 112.605 ;
        RECT 126.985 111.635 127.325 112.605 ;
        RECT 127.500 112.475 127.850 113.125 ;
        RECT 128.020 112.305 128.250 113.295 ;
        RECT 127.585 112.135 128.250 112.305 ;
        RECT 127.585 111.635 127.755 112.135 ;
        RECT 127.925 111.465 128.255 111.965 ;
        RECT 128.425 111.635 128.610 113.755 ;
        RECT 128.865 113.555 129.115 114.015 ;
        RECT 129.285 113.565 129.620 113.735 ;
        RECT 129.815 113.565 130.490 113.735 ;
        RECT 129.285 113.425 129.455 113.565 ;
        RECT 128.780 112.435 129.060 113.385 ;
        RECT 129.230 113.295 129.455 113.425 ;
        RECT 129.230 112.190 129.400 113.295 ;
        RECT 129.625 113.145 130.150 113.365 ;
        RECT 129.570 112.380 129.810 112.975 ;
        RECT 129.980 112.445 130.150 113.145 ;
        RECT 130.320 112.785 130.490 113.565 ;
        RECT 130.810 113.515 131.180 114.015 ;
        RECT 131.360 113.565 131.765 113.735 ;
        RECT 131.935 113.565 132.720 113.735 ;
        RECT 131.360 113.335 131.530 113.565 ;
        RECT 130.700 113.035 131.530 113.335 ;
        RECT 131.915 113.065 132.380 113.395 ;
        RECT 130.700 113.005 130.900 113.035 ;
        RECT 131.020 112.785 131.190 112.855 ;
        RECT 130.320 112.615 131.190 112.785 ;
        RECT 130.680 112.525 131.190 112.615 ;
        RECT 129.230 112.060 129.535 112.190 ;
        RECT 129.980 112.080 130.510 112.445 ;
        RECT 128.850 111.465 129.115 111.925 ;
        RECT 129.285 111.635 129.535 112.060 ;
        RECT 130.680 111.910 130.850 112.525 ;
        RECT 129.745 111.740 130.850 111.910 ;
        RECT 131.020 111.465 131.190 112.265 ;
        RECT 131.360 111.965 131.530 113.035 ;
        RECT 131.700 112.135 131.890 112.855 ;
        RECT 132.060 112.105 132.380 113.065 ;
        RECT 132.550 113.105 132.720 113.565 ;
        RECT 132.995 113.485 133.205 114.015 ;
        RECT 133.465 113.275 133.795 113.800 ;
        RECT 133.965 113.405 134.135 114.015 ;
        RECT 134.305 113.360 134.635 113.795 ;
        RECT 135.865 113.465 136.035 113.845 ;
        RECT 136.250 113.635 136.580 114.015 ;
        RECT 134.305 113.275 134.685 113.360 ;
        RECT 135.865 113.295 136.580 113.465 ;
        RECT 133.595 113.105 133.795 113.275 ;
        RECT 134.460 113.235 134.685 113.275 ;
        RECT 132.550 112.775 133.425 113.105 ;
        RECT 133.595 112.775 134.345 113.105 ;
        RECT 131.360 111.635 131.610 111.965 ;
        RECT 132.550 111.935 132.720 112.775 ;
        RECT 133.595 112.570 133.785 112.775 ;
        RECT 134.515 112.655 134.685 113.235 ;
        RECT 135.775 112.745 136.130 113.115 ;
        RECT 136.410 113.105 136.580 113.295 ;
        RECT 136.750 113.270 137.005 113.845 ;
        RECT 136.410 112.775 136.665 113.105 ;
        RECT 134.470 112.605 134.685 112.655 ;
        RECT 132.890 112.195 133.785 112.570 ;
        RECT 134.295 112.525 134.685 112.605 ;
        RECT 136.410 112.565 136.580 112.775 ;
        RECT 131.835 111.765 132.720 111.935 ;
        RECT 132.900 111.465 133.215 111.965 ;
        RECT 133.445 111.635 133.785 112.195 ;
        RECT 133.955 111.465 134.125 112.475 ;
        RECT 134.295 111.680 134.625 112.525 ;
        RECT 135.865 112.395 136.580 112.565 ;
        RECT 136.835 112.540 137.005 113.270 ;
        RECT 137.180 113.175 137.440 114.015 ;
        RECT 137.615 113.265 138.825 114.015 ;
        RECT 135.865 111.635 136.035 112.395 ;
        RECT 136.250 111.465 136.580 112.225 ;
        RECT 136.750 111.635 137.005 112.540 ;
        RECT 137.180 111.465 137.440 112.615 ;
        RECT 137.615 112.555 138.135 113.095 ;
        RECT 138.305 112.725 138.825 113.265 ;
        RECT 137.615 111.465 138.825 112.555 ;
        RECT 13.330 111.295 138.910 111.465 ;
        RECT 13.415 110.205 14.625 111.295 ;
        RECT 14.795 110.205 17.385 111.295 ;
        RECT 17.645 110.625 17.815 111.125 ;
        RECT 17.985 110.795 18.315 111.295 ;
        RECT 17.645 110.455 18.310 110.625 ;
        RECT 13.415 109.495 13.935 110.035 ;
        RECT 14.105 109.665 14.625 110.205 ;
        RECT 14.795 109.515 16.005 110.035 ;
        RECT 16.175 109.685 17.385 110.205 ;
        RECT 17.560 109.635 17.910 110.285 ;
        RECT 13.415 108.745 14.625 109.495 ;
        RECT 14.795 108.745 17.385 109.515 ;
        RECT 18.080 109.465 18.310 110.455 ;
        RECT 17.645 109.295 18.310 109.465 ;
        RECT 17.645 109.005 17.815 109.295 ;
        RECT 17.985 108.745 18.315 109.125 ;
        RECT 18.485 109.005 18.670 111.125 ;
        RECT 18.910 110.835 19.175 111.295 ;
        RECT 19.345 110.700 19.595 111.125 ;
        RECT 19.805 110.850 20.910 111.020 ;
        RECT 19.290 110.570 19.595 110.700 ;
        RECT 18.840 109.375 19.120 110.325 ;
        RECT 19.290 109.465 19.460 110.570 ;
        RECT 19.630 109.785 19.870 110.380 ;
        RECT 20.040 110.315 20.570 110.680 ;
        RECT 20.040 109.615 20.210 110.315 ;
        RECT 20.740 110.235 20.910 110.850 ;
        RECT 21.080 110.495 21.250 111.295 ;
        RECT 21.420 110.795 21.670 111.125 ;
        RECT 21.895 110.825 22.780 110.995 ;
        RECT 20.740 110.145 21.250 110.235 ;
        RECT 19.290 109.335 19.515 109.465 ;
        RECT 19.685 109.395 20.210 109.615 ;
        RECT 20.380 109.975 21.250 110.145 ;
        RECT 18.925 108.745 19.175 109.205 ;
        RECT 19.345 109.195 19.515 109.335 ;
        RECT 20.380 109.195 20.550 109.975 ;
        RECT 21.080 109.905 21.250 109.975 ;
        RECT 20.760 109.725 20.960 109.755 ;
        RECT 21.420 109.725 21.590 110.795 ;
        RECT 21.760 109.905 21.950 110.625 ;
        RECT 20.760 109.425 21.590 109.725 ;
        RECT 22.120 109.695 22.440 110.655 ;
        RECT 19.345 109.025 19.680 109.195 ;
        RECT 19.875 109.025 20.550 109.195 ;
        RECT 20.870 108.745 21.240 109.245 ;
        RECT 21.420 109.195 21.590 109.425 ;
        RECT 21.975 109.365 22.440 109.695 ;
        RECT 22.610 109.985 22.780 110.825 ;
        RECT 22.960 110.795 23.275 111.295 ;
        RECT 23.505 110.565 23.845 111.125 ;
        RECT 22.950 110.190 23.845 110.565 ;
        RECT 24.015 110.285 24.185 111.295 ;
        RECT 23.655 109.985 23.845 110.190 ;
        RECT 24.355 110.235 24.685 111.080 ;
        RECT 24.355 110.155 24.745 110.235 ;
        RECT 24.915 110.205 26.125 111.295 ;
        RECT 24.530 110.105 24.745 110.155 ;
        RECT 22.610 109.655 23.485 109.985 ;
        RECT 23.655 109.655 24.405 109.985 ;
        RECT 22.610 109.195 22.780 109.655 ;
        RECT 23.655 109.485 23.855 109.655 ;
        RECT 24.575 109.525 24.745 110.105 ;
        RECT 24.520 109.485 24.745 109.525 ;
        RECT 21.420 109.025 21.825 109.195 ;
        RECT 21.995 109.025 22.780 109.195 ;
        RECT 23.055 108.745 23.265 109.275 ;
        RECT 23.525 108.960 23.855 109.485 ;
        RECT 24.365 109.400 24.745 109.485 ;
        RECT 24.915 109.495 25.435 110.035 ;
        RECT 25.605 109.665 26.125 110.205 ;
        RECT 26.295 110.130 26.585 111.295 ;
        RECT 26.760 110.915 27.095 111.295 ;
        RECT 24.025 108.745 24.195 109.355 ;
        RECT 24.365 108.965 24.695 109.400 ;
        RECT 24.915 108.745 26.125 109.495 ;
        RECT 26.295 108.745 26.585 109.470 ;
        RECT 26.755 109.425 26.995 110.735 ;
        RECT 27.265 110.325 27.515 111.125 ;
        RECT 27.735 110.575 28.065 111.295 ;
        RECT 28.250 110.325 28.500 111.125 ;
        RECT 28.965 110.495 29.295 111.295 ;
        RECT 29.465 110.865 29.805 111.125 ;
        RECT 27.165 110.155 29.355 110.325 ;
        RECT 27.165 109.245 27.335 110.155 ;
        RECT 29.040 109.985 29.355 110.155 ;
        RECT 26.840 108.915 27.335 109.245 ;
        RECT 27.555 109.020 27.905 109.985 ;
        RECT 28.085 109.015 28.385 109.985 ;
        RECT 28.565 109.015 28.845 109.985 ;
        RECT 29.040 109.735 29.370 109.985 ;
        RECT 29.025 108.745 29.295 109.545 ;
        RECT 29.545 109.465 29.805 110.865 ;
        RECT 29.975 110.860 35.320 111.295 ;
        RECT 35.495 110.860 40.840 111.295 ;
        RECT 29.465 108.955 29.805 109.465 ;
        RECT 31.560 109.290 31.900 110.120 ;
        RECT 33.380 109.610 33.730 110.860 ;
        RECT 37.080 109.290 37.420 110.120 ;
        RECT 38.900 109.610 39.250 110.860 ;
        RECT 41.015 110.205 42.685 111.295 ;
        RECT 41.015 109.515 41.765 110.035 ;
        RECT 41.935 109.685 42.685 110.205 ;
        RECT 42.855 110.325 43.125 111.095 ;
        RECT 43.295 110.515 43.625 111.295 ;
        RECT 43.830 110.690 44.015 111.095 ;
        RECT 44.185 110.870 44.520 111.295 ;
        RECT 43.830 110.515 44.495 110.690 ;
        RECT 42.855 110.155 43.985 110.325 ;
        RECT 29.975 108.745 35.320 109.290 ;
        RECT 35.495 108.745 40.840 109.290 ;
        RECT 41.015 108.745 42.685 109.515 ;
        RECT 42.855 109.245 43.025 110.155 ;
        RECT 43.195 109.405 43.555 109.985 ;
        RECT 43.735 109.655 43.985 110.155 ;
        RECT 44.155 109.485 44.495 110.515 ;
        RECT 44.755 110.235 45.085 111.080 ;
        RECT 45.255 110.285 45.425 111.295 ;
        RECT 45.595 110.565 45.935 111.125 ;
        RECT 46.165 110.795 46.480 111.295 ;
        RECT 46.660 110.825 47.545 110.995 ;
        RECT 43.810 109.315 44.495 109.485 ;
        RECT 44.695 110.155 45.085 110.235 ;
        RECT 45.595 110.190 46.490 110.565 ;
        RECT 44.695 110.105 44.910 110.155 ;
        RECT 44.695 109.525 44.865 110.105 ;
        RECT 45.595 109.985 45.785 110.190 ;
        RECT 46.660 109.985 46.830 110.825 ;
        RECT 47.770 110.795 48.020 111.125 ;
        RECT 45.035 109.655 45.785 109.985 ;
        RECT 45.955 109.655 46.830 109.985 ;
        RECT 44.695 109.485 44.920 109.525 ;
        RECT 45.585 109.485 45.785 109.655 ;
        RECT 44.695 109.400 45.075 109.485 ;
        RECT 42.855 108.915 43.115 109.245 ;
        RECT 43.325 108.745 43.600 109.225 ;
        RECT 43.810 108.915 44.015 109.315 ;
        RECT 44.185 108.745 44.520 109.145 ;
        RECT 44.745 108.965 45.075 109.400 ;
        RECT 45.245 108.745 45.415 109.355 ;
        RECT 45.585 108.960 45.915 109.485 ;
        RECT 46.175 108.745 46.385 109.275 ;
        RECT 46.660 109.195 46.830 109.655 ;
        RECT 47.000 109.695 47.320 110.655 ;
        RECT 47.490 109.905 47.680 110.625 ;
        RECT 47.850 109.725 48.020 110.795 ;
        RECT 48.190 110.495 48.360 111.295 ;
        RECT 48.530 110.850 49.635 111.020 ;
        RECT 48.530 110.235 48.700 110.850 ;
        RECT 49.845 110.700 50.095 111.125 ;
        RECT 50.265 110.835 50.530 111.295 ;
        RECT 48.870 110.315 49.400 110.680 ;
        RECT 49.845 110.570 50.150 110.700 ;
        RECT 48.190 110.145 48.700 110.235 ;
        RECT 48.190 109.975 49.060 110.145 ;
        RECT 48.190 109.905 48.360 109.975 ;
        RECT 48.480 109.725 48.680 109.755 ;
        RECT 47.000 109.365 47.465 109.695 ;
        RECT 47.850 109.425 48.680 109.725 ;
        RECT 47.850 109.195 48.020 109.425 ;
        RECT 46.660 109.025 47.445 109.195 ;
        RECT 47.615 109.025 48.020 109.195 ;
        RECT 48.200 108.745 48.570 109.245 ;
        RECT 48.890 109.195 49.060 109.975 ;
        RECT 49.230 109.615 49.400 110.315 ;
        RECT 49.570 109.785 49.810 110.380 ;
        RECT 49.230 109.395 49.755 109.615 ;
        RECT 49.980 109.465 50.150 110.570 ;
        RECT 49.925 109.335 50.150 109.465 ;
        RECT 50.320 109.375 50.600 110.325 ;
        RECT 49.925 109.195 50.095 109.335 ;
        RECT 48.890 109.025 49.565 109.195 ;
        RECT 49.760 109.025 50.095 109.195 ;
        RECT 50.265 108.745 50.515 109.205 ;
        RECT 50.770 109.005 50.955 111.125 ;
        RECT 51.125 110.795 51.455 111.295 ;
        RECT 51.625 110.625 51.795 111.125 ;
        RECT 51.130 110.455 51.795 110.625 ;
        RECT 51.130 109.465 51.360 110.455 ;
        RECT 51.530 109.635 51.880 110.285 ;
        RECT 52.055 110.130 52.345 111.295 ;
        RECT 52.630 110.665 52.915 111.125 ;
        RECT 53.085 110.835 53.355 111.295 ;
        RECT 52.630 110.445 53.585 110.665 ;
        RECT 52.515 109.715 53.205 110.275 ;
        RECT 53.375 109.545 53.585 110.445 ;
        RECT 51.130 109.295 51.795 109.465 ;
        RECT 51.125 108.745 51.455 109.125 ;
        RECT 51.625 109.005 51.795 109.295 ;
        RECT 52.055 108.745 52.345 109.470 ;
        RECT 52.630 109.375 53.585 109.545 ;
        RECT 53.755 110.275 54.155 111.125 ;
        RECT 54.345 110.665 54.625 111.125 ;
        RECT 55.145 110.835 55.470 111.295 ;
        RECT 54.345 110.445 55.470 110.665 ;
        RECT 53.755 109.715 54.850 110.275 ;
        RECT 55.020 109.985 55.470 110.445 ;
        RECT 55.640 110.155 56.025 111.125 ;
        RECT 56.235 110.155 56.465 111.295 ;
        RECT 52.630 108.915 52.915 109.375 ;
        RECT 53.085 108.745 53.355 109.205 ;
        RECT 53.755 108.915 54.155 109.715 ;
        RECT 55.020 109.655 55.575 109.985 ;
        RECT 55.020 109.545 55.470 109.655 ;
        RECT 54.345 109.375 55.470 109.545 ;
        RECT 55.745 109.485 56.025 110.155 ;
        RECT 56.635 110.145 56.965 111.125 ;
        RECT 57.135 110.155 57.345 111.295 ;
        RECT 57.575 110.205 61.085 111.295 ;
        RECT 56.215 109.735 56.545 109.985 ;
        RECT 54.345 108.915 54.625 109.375 ;
        RECT 55.145 108.745 55.470 109.205 ;
        RECT 55.640 108.915 56.025 109.485 ;
        RECT 56.235 108.745 56.465 109.565 ;
        RECT 56.715 109.545 56.965 110.145 ;
        RECT 56.635 108.915 56.965 109.545 ;
        RECT 57.135 108.745 57.345 109.565 ;
        RECT 57.575 109.515 59.225 110.035 ;
        RECT 59.395 109.685 61.085 110.205 ;
        RECT 61.260 110.155 61.580 111.295 ;
        RECT 61.760 109.985 61.955 111.035 ;
        RECT 62.135 110.445 62.465 111.125 ;
        RECT 62.665 110.495 62.920 111.295 ;
        RECT 63.185 110.625 63.355 111.125 ;
        RECT 63.525 110.795 63.855 111.295 ;
        RECT 63.185 110.455 63.850 110.625 ;
        RECT 62.135 110.165 62.485 110.445 ;
        RECT 61.320 109.935 61.580 109.985 ;
        RECT 61.315 109.765 61.580 109.935 ;
        RECT 61.320 109.655 61.580 109.765 ;
        RECT 61.760 109.655 62.145 109.985 ;
        RECT 62.315 109.785 62.485 110.165 ;
        RECT 62.675 109.955 62.920 110.315 ;
        RECT 62.315 109.615 62.835 109.785 ;
        RECT 63.100 109.635 63.450 110.285 ;
        RECT 57.575 108.745 61.085 109.515 ;
        RECT 61.260 109.275 62.475 109.445 ;
        RECT 61.260 108.925 61.550 109.275 ;
        RECT 61.745 108.745 62.075 109.105 ;
        RECT 62.245 108.970 62.475 109.275 ;
        RECT 62.665 109.255 62.835 109.615 ;
        RECT 63.620 109.465 63.850 110.455 ;
        RECT 63.185 109.295 63.850 109.465 ;
        RECT 62.665 109.085 62.865 109.255 ;
        RECT 62.665 109.050 62.835 109.085 ;
        RECT 63.185 109.005 63.355 109.295 ;
        RECT 63.525 108.745 63.855 109.125 ;
        RECT 64.025 109.005 64.210 111.125 ;
        RECT 64.450 110.835 64.715 111.295 ;
        RECT 64.885 110.700 65.135 111.125 ;
        RECT 65.345 110.850 66.450 111.020 ;
        RECT 64.830 110.570 65.135 110.700 ;
        RECT 64.380 109.375 64.660 110.325 ;
        RECT 64.830 109.465 65.000 110.570 ;
        RECT 65.170 109.785 65.410 110.380 ;
        RECT 65.580 110.315 66.110 110.680 ;
        RECT 65.580 109.615 65.750 110.315 ;
        RECT 66.280 110.235 66.450 110.850 ;
        RECT 66.620 110.495 66.790 111.295 ;
        RECT 66.960 110.795 67.210 111.125 ;
        RECT 67.435 110.825 68.320 110.995 ;
        RECT 66.280 110.145 66.790 110.235 ;
        RECT 64.830 109.335 65.055 109.465 ;
        RECT 65.225 109.395 65.750 109.615 ;
        RECT 65.920 109.975 66.790 110.145 ;
        RECT 64.465 108.745 64.715 109.205 ;
        RECT 64.885 109.195 65.055 109.335 ;
        RECT 65.920 109.195 66.090 109.975 ;
        RECT 66.620 109.905 66.790 109.975 ;
        RECT 66.300 109.725 66.500 109.755 ;
        RECT 66.960 109.725 67.130 110.795 ;
        RECT 67.300 109.905 67.490 110.625 ;
        RECT 66.300 109.425 67.130 109.725 ;
        RECT 67.660 109.695 67.980 110.655 ;
        RECT 64.885 109.025 65.220 109.195 ;
        RECT 65.415 109.025 66.090 109.195 ;
        RECT 66.410 108.745 66.780 109.245 ;
        RECT 66.960 109.195 67.130 109.425 ;
        RECT 67.515 109.365 67.980 109.695 ;
        RECT 68.150 109.985 68.320 110.825 ;
        RECT 68.500 110.795 68.815 111.295 ;
        RECT 69.045 110.565 69.385 111.125 ;
        RECT 68.490 110.190 69.385 110.565 ;
        RECT 69.555 110.285 69.725 111.295 ;
        RECT 69.195 109.985 69.385 110.190 ;
        RECT 69.895 110.235 70.225 111.080 ;
        RECT 70.455 110.860 75.800 111.295 ;
        RECT 69.895 110.155 70.285 110.235 ;
        RECT 70.070 110.105 70.285 110.155 ;
        RECT 68.150 109.655 69.025 109.985 ;
        RECT 69.195 109.655 69.945 109.985 ;
        RECT 68.150 109.195 68.320 109.655 ;
        RECT 69.195 109.485 69.395 109.655 ;
        RECT 70.115 109.525 70.285 110.105 ;
        RECT 70.060 109.485 70.285 109.525 ;
        RECT 66.960 109.025 67.365 109.195 ;
        RECT 67.535 109.025 68.320 109.195 ;
        RECT 68.595 108.745 68.805 109.275 ;
        RECT 69.065 108.960 69.395 109.485 ;
        RECT 69.905 109.400 70.285 109.485 ;
        RECT 69.565 108.745 69.735 109.355 ;
        RECT 69.905 108.965 70.235 109.400 ;
        RECT 72.040 109.290 72.380 110.120 ;
        RECT 73.860 109.610 74.210 110.860 ;
        RECT 75.975 110.205 77.645 111.295 ;
        RECT 75.975 109.515 76.725 110.035 ;
        RECT 76.895 109.685 77.645 110.205 ;
        RECT 77.815 110.130 78.105 111.295 ;
        RECT 78.460 110.325 78.850 110.500 ;
        RECT 79.335 110.495 79.665 111.295 ;
        RECT 79.835 110.505 80.370 111.125 ;
        RECT 78.460 110.155 79.885 110.325 ;
        RECT 70.455 108.745 75.800 109.290 ;
        RECT 75.975 108.745 77.645 109.515 ;
        RECT 77.815 108.745 78.105 109.470 ;
        RECT 78.335 109.425 78.690 109.985 ;
        RECT 78.860 109.255 79.030 110.155 ;
        RECT 79.200 109.425 79.465 109.985 ;
        RECT 79.715 109.655 79.885 110.155 ;
        RECT 80.055 109.485 80.370 110.505 ;
        RECT 80.575 110.205 82.245 111.295 ;
        RECT 78.440 108.745 78.680 109.255 ;
        RECT 78.860 108.925 79.140 109.255 ;
        RECT 79.370 108.745 79.585 109.255 ;
        RECT 79.755 108.915 80.370 109.485 ;
        RECT 80.575 109.515 81.325 110.035 ;
        RECT 81.495 109.685 82.245 110.205 ;
        RECT 82.420 110.345 82.685 111.115 ;
        RECT 82.855 110.575 83.185 111.295 ;
        RECT 83.375 110.755 83.635 111.115 ;
        RECT 83.805 110.925 84.135 111.295 ;
        RECT 84.305 110.755 84.565 111.115 ;
        RECT 83.375 110.525 84.565 110.755 ;
        RECT 85.135 110.345 85.425 111.115 ;
        RECT 86.805 110.565 87.100 111.295 ;
        RECT 87.270 110.395 87.530 111.120 ;
        RECT 87.700 110.565 87.960 111.295 ;
        RECT 88.130 110.395 88.390 111.120 ;
        RECT 88.560 110.565 88.820 111.295 ;
        RECT 88.990 110.395 89.250 111.120 ;
        RECT 89.420 110.565 89.680 111.295 ;
        RECT 89.850 110.395 90.110 111.120 ;
        RECT 80.575 108.745 82.245 109.515 ;
        RECT 82.420 108.925 82.755 110.345 ;
        RECT 82.930 110.165 85.425 110.345 ;
        RECT 82.930 109.475 83.155 110.165 ;
        RECT 86.800 110.155 90.110 110.395 ;
        RECT 90.280 110.185 90.540 111.295 ;
        RECT 83.355 109.655 83.635 109.985 ;
        RECT 83.815 109.655 84.390 109.985 ;
        RECT 84.570 109.655 85.005 109.985 ;
        RECT 85.185 109.655 85.455 109.985 ;
        RECT 86.800 109.565 87.770 110.155 ;
        RECT 90.710 109.985 90.960 111.120 ;
        RECT 91.140 110.185 91.435 111.295 ;
        RECT 91.650 110.505 92.185 111.125 ;
        RECT 87.940 109.735 90.960 109.985 ;
        RECT 82.930 109.285 85.415 109.475 ;
        RECT 86.800 109.395 90.110 109.565 ;
        RECT 82.935 108.745 83.680 109.115 ;
        RECT 84.245 108.925 84.500 109.285 ;
        RECT 84.680 108.745 85.010 109.115 ;
        RECT 85.190 108.925 85.415 109.285 ;
        RECT 86.800 108.745 87.100 109.225 ;
        RECT 87.270 108.940 87.530 109.395 ;
        RECT 87.700 108.745 87.960 109.225 ;
        RECT 88.130 108.940 88.390 109.395 ;
        RECT 88.560 108.745 88.820 109.225 ;
        RECT 88.990 108.940 89.250 109.395 ;
        RECT 89.420 108.745 89.680 109.225 ;
        RECT 89.850 108.940 90.110 109.395 ;
        RECT 90.280 108.745 90.540 109.270 ;
        RECT 90.710 108.925 90.960 109.735 ;
        RECT 91.130 109.375 91.445 109.985 ;
        RECT 91.650 109.485 91.965 110.505 ;
        RECT 92.355 110.495 92.685 111.295 ;
        RECT 93.170 110.325 93.560 110.500 ;
        RECT 92.135 110.155 93.560 110.325 ;
        RECT 93.915 110.205 97.425 111.295 ;
        RECT 92.135 109.655 92.305 110.155 ;
        RECT 91.140 108.745 91.385 109.205 ;
        RECT 91.650 108.915 92.265 109.485 ;
        RECT 92.555 109.425 92.820 109.985 ;
        RECT 92.990 109.255 93.160 110.155 ;
        RECT 93.330 109.425 93.685 109.985 ;
        RECT 93.915 109.515 95.565 110.035 ;
        RECT 95.735 109.685 97.425 110.205 ;
        RECT 97.630 110.505 98.165 111.125 ;
        RECT 92.435 108.745 92.650 109.255 ;
        RECT 92.880 108.925 93.160 109.255 ;
        RECT 93.340 108.745 93.580 109.255 ;
        RECT 93.915 108.745 97.425 109.515 ;
        RECT 97.630 109.485 97.945 110.505 ;
        RECT 98.335 110.495 98.665 111.295 ;
        RECT 99.150 110.325 99.540 110.500 ;
        RECT 98.115 110.155 99.540 110.325 ;
        RECT 100.100 110.325 100.430 111.125 ;
        RECT 100.600 110.495 100.930 111.295 ;
        RECT 101.230 110.325 101.560 111.125 ;
        RECT 102.205 110.495 102.455 111.295 ;
        RECT 100.100 110.155 102.535 110.325 ;
        RECT 102.725 110.155 102.895 111.295 ;
        RECT 103.065 110.155 103.405 111.125 ;
        RECT 98.115 109.655 98.285 110.155 ;
        RECT 97.630 108.915 98.245 109.485 ;
        RECT 98.535 109.425 98.800 109.985 ;
        RECT 98.970 109.255 99.140 110.155 ;
        RECT 99.310 109.425 99.665 109.985 ;
        RECT 99.895 109.735 100.245 109.985 ;
        RECT 100.430 109.525 100.600 110.155 ;
        RECT 100.770 109.735 101.100 109.935 ;
        RECT 101.270 109.735 101.600 109.935 ;
        RECT 101.770 109.735 102.190 109.935 ;
        RECT 102.365 109.905 102.535 110.155 ;
        RECT 102.365 109.735 103.060 109.905 ;
        RECT 103.230 109.595 103.405 110.155 ;
        RECT 103.575 110.130 103.865 111.295 ;
        RECT 104.125 110.625 104.295 111.125 ;
        RECT 104.465 110.795 104.795 111.295 ;
        RECT 104.125 110.455 104.790 110.625 ;
        RECT 104.040 109.635 104.390 110.285 ;
        RECT 98.415 108.745 98.630 109.255 ;
        RECT 98.860 108.925 99.140 109.255 ;
        RECT 99.320 108.745 99.560 109.255 ;
        RECT 100.100 108.915 100.600 109.525 ;
        RECT 101.230 109.395 102.455 109.565 ;
        RECT 103.175 109.545 103.405 109.595 ;
        RECT 101.230 108.915 101.560 109.395 ;
        RECT 101.730 108.745 101.955 109.205 ;
        RECT 102.125 108.915 102.455 109.395 ;
        RECT 102.645 108.745 102.895 109.545 ;
        RECT 103.065 108.915 103.405 109.545 ;
        RECT 103.575 108.745 103.865 109.470 ;
        RECT 104.560 109.465 104.790 110.455 ;
        RECT 104.125 109.295 104.790 109.465 ;
        RECT 104.125 109.005 104.295 109.295 ;
        RECT 104.465 108.745 104.795 109.125 ;
        RECT 104.965 109.005 105.150 111.125 ;
        RECT 105.390 110.835 105.655 111.295 ;
        RECT 105.825 110.700 106.075 111.125 ;
        RECT 106.285 110.850 107.390 111.020 ;
        RECT 105.770 110.570 106.075 110.700 ;
        RECT 105.320 109.375 105.600 110.325 ;
        RECT 105.770 109.465 105.940 110.570 ;
        RECT 106.110 109.785 106.350 110.380 ;
        RECT 106.520 110.315 107.050 110.680 ;
        RECT 106.520 109.615 106.690 110.315 ;
        RECT 107.220 110.235 107.390 110.850 ;
        RECT 107.560 110.495 107.730 111.295 ;
        RECT 107.900 110.795 108.150 111.125 ;
        RECT 108.375 110.825 109.260 110.995 ;
        RECT 107.220 110.145 107.730 110.235 ;
        RECT 105.770 109.335 105.995 109.465 ;
        RECT 106.165 109.395 106.690 109.615 ;
        RECT 106.860 109.975 107.730 110.145 ;
        RECT 105.405 108.745 105.655 109.205 ;
        RECT 105.825 109.195 105.995 109.335 ;
        RECT 106.860 109.195 107.030 109.975 ;
        RECT 107.560 109.905 107.730 109.975 ;
        RECT 107.240 109.725 107.440 109.755 ;
        RECT 107.900 109.725 108.070 110.795 ;
        RECT 108.240 109.905 108.430 110.625 ;
        RECT 107.240 109.425 108.070 109.725 ;
        RECT 108.600 109.695 108.920 110.655 ;
        RECT 105.825 109.025 106.160 109.195 ;
        RECT 106.355 109.025 107.030 109.195 ;
        RECT 107.350 108.745 107.720 109.245 ;
        RECT 107.900 109.195 108.070 109.425 ;
        RECT 108.455 109.365 108.920 109.695 ;
        RECT 109.090 109.985 109.260 110.825 ;
        RECT 109.440 110.795 109.755 111.295 ;
        RECT 109.985 110.565 110.325 111.125 ;
        RECT 109.430 110.190 110.325 110.565 ;
        RECT 110.495 110.285 110.665 111.295 ;
        RECT 110.135 109.985 110.325 110.190 ;
        RECT 110.835 110.235 111.165 111.080 ;
        RECT 111.600 110.325 111.930 111.125 ;
        RECT 112.100 110.495 112.430 111.295 ;
        RECT 112.730 110.325 113.060 111.125 ;
        RECT 113.705 110.495 113.955 111.295 ;
        RECT 110.835 110.155 111.225 110.235 ;
        RECT 111.600 110.155 114.035 110.325 ;
        RECT 114.225 110.155 114.395 111.295 ;
        RECT 114.565 110.155 114.905 111.125 ;
        RECT 115.075 110.205 118.585 111.295 ;
        RECT 118.955 110.625 119.235 111.295 ;
        RECT 119.405 110.405 119.705 110.955 ;
        RECT 119.905 110.575 120.235 111.295 ;
        RECT 120.425 110.575 120.885 111.125 ;
        RECT 111.010 110.105 111.225 110.155 ;
        RECT 109.090 109.655 109.965 109.985 ;
        RECT 110.135 109.655 110.885 109.985 ;
        RECT 109.090 109.195 109.260 109.655 ;
        RECT 110.135 109.485 110.335 109.655 ;
        RECT 111.055 109.525 111.225 110.105 ;
        RECT 111.395 109.735 111.745 109.985 ;
        RECT 111.930 109.525 112.100 110.155 ;
        RECT 112.270 109.735 112.600 109.935 ;
        RECT 112.770 109.735 113.100 109.935 ;
        RECT 113.270 109.735 113.690 109.935 ;
        RECT 113.865 109.905 114.035 110.155 ;
        RECT 113.865 109.735 114.560 109.905 ;
        RECT 111.000 109.485 111.225 109.525 ;
        RECT 107.900 109.025 108.305 109.195 ;
        RECT 108.475 109.025 109.260 109.195 ;
        RECT 109.535 108.745 109.745 109.275 ;
        RECT 110.005 108.960 110.335 109.485 ;
        RECT 110.845 109.400 111.225 109.485 ;
        RECT 110.505 108.745 110.675 109.355 ;
        RECT 110.845 108.965 111.175 109.400 ;
        RECT 111.600 108.915 112.100 109.525 ;
        RECT 112.730 109.395 113.955 109.565 ;
        RECT 114.730 109.545 114.905 110.155 ;
        RECT 112.730 108.915 113.060 109.395 ;
        RECT 113.230 108.745 113.455 109.205 ;
        RECT 113.625 108.915 113.955 109.395 ;
        RECT 114.145 108.745 114.395 109.545 ;
        RECT 114.565 108.915 114.905 109.545 ;
        RECT 115.075 109.515 116.725 110.035 ;
        RECT 116.895 109.685 118.585 110.205 ;
        RECT 118.770 109.985 119.035 110.345 ;
        RECT 119.405 110.235 120.345 110.405 ;
        RECT 120.175 109.985 120.345 110.235 ;
        RECT 118.770 109.735 119.445 109.985 ;
        RECT 119.665 109.735 120.005 109.985 ;
        RECT 120.175 109.655 120.465 109.985 ;
        RECT 120.175 109.565 120.345 109.655 ;
        RECT 115.075 108.745 118.585 109.515 ;
        RECT 118.955 109.375 120.345 109.565 ;
        RECT 118.955 109.015 119.285 109.375 ;
        RECT 120.635 109.205 120.885 110.575 ;
        RECT 119.905 108.745 120.155 109.205 ;
        RECT 120.325 108.915 120.885 109.205 ;
        RECT 121.090 110.505 121.625 111.125 ;
        RECT 121.090 109.485 121.405 110.505 ;
        RECT 121.795 110.495 122.125 111.295 ;
        RECT 122.610 110.325 123.000 110.500 ;
        RECT 121.575 110.155 123.000 110.325 ;
        RECT 123.355 110.205 125.025 111.295 ;
        RECT 121.575 109.655 121.745 110.155 ;
        RECT 121.090 108.915 121.705 109.485 ;
        RECT 121.995 109.425 122.260 109.985 ;
        RECT 122.430 109.255 122.600 110.155 ;
        RECT 122.770 109.425 123.125 109.985 ;
        RECT 123.355 109.515 124.105 110.035 ;
        RECT 124.275 109.685 125.025 110.205 ;
        RECT 125.230 110.505 125.765 111.125 ;
        RECT 121.875 108.745 122.090 109.255 ;
        RECT 122.320 108.925 122.600 109.255 ;
        RECT 122.780 108.745 123.020 109.255 ;
        RECT 123.355 108.745 125.025 109.515 ;
        RECT 125.230 109.485 125.545 110.505 ;
        RECT 125.935 110.495 126.265 111.295 ;
        RECT 126.750 110.325 127.140 110.500 ;
        RECT 125.715 110.155 127.140 110.325 ;
        RECT 127.495 110.205 129.165 111.295 ;
        RECT 125.715 109.655 125.885 110.155 ;
        RECT 125.230 108.915 125.845 109.485 ;
        RECT 126.135 109.425 126.400 109.985 ;
        RECT 126.570 109.255 126.740 110.155 ;
        RECT 126.910 109.425 127.265 109.985 ;
        RECT 127.495 109.515 128.245 110.035 ;
        RECT 128.415 109.685 129.165 110.205 ;
        RECT 129.335 110.130 129.625 111.295 ;
        RECT 129.795 110.445 130.055 111.125 ;
        RECT 130.225 110.515 130.475 111.295 ;
        RECT 130.725 110.745 130.975 111.125 ;
        RECT 131.145 110.915 131.500 111.295 ;
        RECT 132.505 110.905 132.840 111.125 ;
        RECT 132.105 110.745 132.335 110.785 ;
        RECT 130.725 110.545 132.335 110.745 ;
        RECT 130.725 110.535 131.560 110.545 ;
        RECT 132.150 110.455 132.335 110.545 ;
        RECT 126.015 108.745 126.230 109.255 ;
        RECT 126.460 108.925 126.740 109.255 ;
        RECT 126.920 108.745 127.160 109.255 ;
        RECT 127.495 108.745 129.165 109.515 ;
        RECT 129.335 108.745 129.625 109.470 ;
        RECT 129.795 109.255 129.965 110.445 ;
        RECT 131.665 110.345 131.995 110.375 ;
        RECT 130.195 110.285 131.995 110.345 ;
        RECT 132.585 110.285 132.840 110.905 ;
        RECT 130.135 110.175 132.840 110.285 ;
        RECT 134.025 110.365 134.195 111.125 ;
        RECT 134.410 110.535 134.740 111.295 ;
        RECT 134.025 110.195 134.740 110.365 ;
        RECT 134.910 110.220 135.165 111.125 ;
        RECT 130.135 110.140 130.335 110.175 ;
        RECT 130.135 109.565 130.305 110.140 ;
        RECT 131.665 110.115 132.840 110.175 ;
        RECT 130.535 109.700 130.945 110.005 ;
        RECT 131.115 109.735 131.445 109.945 ;
        RECT 130.135 109.445 130.405 109.565 ;
        RECT 130.135 109.400 130.980 109.445 ;
        RECT 130.225 109.275 130.980 109.400 ;
        RECT 131.235 109.335 131.445 109.735 ;
        RECT 131.690 109.735 132.165 109.945 ;
        RECT 132.355 109.735 132.845 109.935 ;
        RECT 131.690 109.335 131.910 109.735 ;
        RECT 133.935 109.645 134.290 110.015 ;
        RECT 134.570 109.985 134.740 110.195 ;
        RECT 134.570 109.655 134.825 109.985 ;
        RECT 129.795 109.245 130.025 109.255 ;
        RECT 129.795 108.915 130.055 109.245 ;
        RECT 130.810 109.125 130.980 109.275 ;
        RECT 130.225 108.745 130.555 109.105 ;
        RECT 130.810 108.915 132.110 109.125 ;
        RECT 132.385 108.745 132.840 109.510 ;
        RECT 134.570 109.465 134.740 109.655 ;
        RECT 134.995 109.490 135.165 110.220 ;
        RECT 135.340 110.145 135.600 111.295 ;
        RECT 135.865 110.365 136.035 111.125 ;
        RECT 136.250 110.535 136.580 111.295 ;
        RECT 135.865 110.195 136.580 110.365 ;
        RECT 136.750 110.220 137.005 111.125 ;
        RECT 135.775 109.645 136.130 110.015 ;
        RECT 136.410 109.985 136.580 110.195 ;
        RECT 136.410 109.655 136.665 109.985 ;
        RECT 134.025 109.295 134.740 109.465 ;
        RECT 134.025 108.915 134.195 109.295 ;
        RECT 134.410 108.745 134.740 109.125 ;
        RECT 134.910 108.915 135.165 109.490 ;
        RECT 135.340 108.745 135.600 109.585 ;
        RECT 136.410 109.465 136.580 109.655 ;
        RECT 136.835 109.490 137.005 110.220 ;
        RECT 137.180 110.145 137.440 111.295 ;
        RECT 137.615 110.205 138.825 111.295 ;
        RECT 137.615 109.665 138.135 110.205 ;
        RECT 135.865 109.295 136.580 109.465 ;
        RECT 135.865 108.915 136.035 109.295 ;
        RECT 136.250 108.745 136.580 109.125 ;
        RECT 136.750 108.915 137.005 109.490 ;
        RECT 137.180 108.745 137.440 109.585 ;
        RECT 138.305 109.495 138.825 110.035 ;
        RECT 137.615 108.745 138.825 109.495 ;
        RECT 13.330 108.575 138.910 108.745 ;
        RECT 13.415 107.825 14.625 108.575 ;
        RECT 13.415 107.285 13.935 107.825 ;
        RECT 14.795 107.805 17.385 108.575 ;
        RECT 17.560 108.085 17.815 108.575 ;
        RECT 17.985 108.065 19.215 108.405 ;
        RECT 14.105 107.115 14.625 107.655 ;
        RECT 14.795 107.285 16.005 107.805 ;
        RECT 16.175 107.115 17.385 107.635 ;
        RECT 17.580 107.335 17.800 107.915 ;
        RECT 17.985 107.165 18.165 108.065 ;
        RECT 18.335 107.335 18.710 107.895 ;
        RECT 18.885 107.835 19.215 108.065 ;
        RECT 19.395 107.925 19.655 108.405 ;
        RECT 19.825 108.035 20.075 108.575 ;
        RECT 18.915 107.335 19.225 107.665 ;
        RECT 13.415 106.025 14.625 107.115 ;
        RECT 14.795 106.025 17.385 107.115 ;
        RECT 17.560 106.025 17.815 107.165 ;
        RECT 17.985 106.995 19.215 107.165 ;
        RECT 17.985 106.195 18.315 106.995 ;
        RECT 18.485 106.025 18.715 106.825 ;
        RECT 18.885 106.195 19.215 106.995 ;
        RECT 19.395 106.895 19.565 107.925 ;
        RECT 20.245 107.895 20.465 108.355 ;
        RECT 20.215 107.870 20.465 107.895 ;
        RECT 19.735 107.275 19.965 107.670 ;
        RECT 20.135 107.445 20.465 107.870 ;
        RECT 20.635 108.195 21.525 108.365 ;
        RECT 20.635 107.470 20.805 108.195 ;
        RECT 20.975 107.640 21.525 108.025 ;
        RECT 21.705 107.850 22.035 108.360 ;
        RECT 22.205 108.175 22.535 108.575 ;
        RECT 23.585 108.005 23.915 108.345 ;
        RECT 24.085 108.175 24.415 108.575 ;
        RECT 20.635 107.400 21.525 107.470 ;
        RECT 20.630 107.375 21.525 107.400 ;
        RECT 20.620 107.360 21.525 107.375 ;
        RECT 20.615 107.345 21.525 107.360 ;
        RECT 20.605 107.340 21.525 107.345 ;
        RECT 20.600 107.330 21.525 107.340 ;
        RECT 20.595 107.320 21.525 107.330 ;
        RECT 20.585 107.315 21.525 107.320 ;
        RECT 20.575 107.305 21.525 107.315 ;
        RECT 20.565 107.300 21.525 107.305 ;
        RECT 20.565 107.295 20.900 107.300 ;
        RECT 20.550 107.290 20.900 107.295 ;
        RECT 20.535 107.280 20.900 107.290 ;
        RECT 20.510 107.275 20.900 107.280 ;
        RECT 19.735 107.270 20.900 107.275 ;
        RECT 19.735 107.235 20.870 107.270 ;
        RECT 19.735 107.210 20.835 107.235 ;
        RECT 19.735 107.180 20.805 107.210 ;
        RECT 19.735 107.150 20.785 107.180 ;
        RECT 19.735 107.120 20.765 107.150 ;
        RECT 19.735 107.110 20.695 107.120 ;
        RECT 19.735 107.100 20.670 107.110 ;
        RECT 19.735 107.085 20.650 107.100 ;
        RECT 19.735 107.070 20.630 107.085 ;
        RECT 19.840 107.060 20.625 107.070 ;
        RECT 19.840 107.025 20.610 107.060 ;
        RECT 19.395 106.195 19.670 106.895 ;
        RECT 19.840 106.775 20.595 107.025 ;
        RECT 20.765 106.705 21.095 106.950 ;
        RECT 21.265 106.850 21.525 107.300 ;
        RECT 21.705 107.085 21.895 107.850 ;
        RECT 22.205 107.835 24.570 108.005 ;
        RECT 24.935 107.845 25.225 108.575 ;
        RECT 22.205 107.665 22.375 107.835 ;
        RECT 22.065 107.335 22.375 107.665 ;
        RECT 22.545 107.335 22.850 107.665 ;
        RECT 20.910 106.680 21.095 106.705 ;
        RECT 20.910 106.580 21.525 106.680 ;
        RECT 19.840 106.025 20.095 106.570 ;
        RECT 20.265 106.195 20.745 106.535 ;
        RECT 20.920 106.025 21.525 106.580 ;
        RECT 21.705 106.235 22.035 107.085 ;
        RECT 22.205 106.025 22.455 107.165 ;
        RECT 22.635 107.005 22.850 107.335 ;
        RECT 23.025 107.005 23.310 107.665 ;
        RECT 23.505 107.005 23.770 107.665 ;
        RECT 23.985 107.005 24.230 107.665 ;
        RECT 24.400 106.835 24.570 107.835 ;
        RECT 24.925 107.335 25.225 107.665 ;
        RECT 25.405 107.645 25.635 108.285 ;
        RECT 25.815 108.025 26.125 108.395 ;
        RECT 26.305 108.205 26.975 108.575 ;
        RECT 25.815 107.825 27.045 108.025 ;
        RECT 25.405 107.335 25.930 107.645 ;
        RECT 26.110 107.335 26.575 107.645 ;
        RECT 26.755 107.155 27.045 107.825 ;
        RECT 22.645 106.665 23.935 106.835 ;
        RECT 22.645 106.245 22.895 106.665 ;
        RECT 23.125 106.025 23.455 106.495 ;
        RECT 23.685 106.245 23.935 106.665 ;
        RECT 24.115 106.665 24.570 106.835 ;
        RECT 24.935 106.915 26.095 107.155 ;
        RECT 24.115 106.235 24.445 106.665 ;
        RECT 24.935 106.205 25.195 106.915 ;
        RECT 25.365 106.025 25.695 106.735 ;
        RECT 25.865 106.205 26.095 106.915 ;
        RECT 26.275 106.935 27.045 107.155 ;
        RECT 26.275 106.205 26.545 106.935 ;
        RECT 26.725 106.025 27.065 106.755 ;
        RECT 27.235 106.205 27.495 108.395 ;
        RECT 27.675 108.030 33.020 108.575 ;
        RECT 33.655 108.195 34.545 108.365 ;
        RECT 29.260 107.200 29.600 108.030 ;
        RECT 31.080 106.460 31.430 107.710 ;
        RECT 33.655 107.640 34.205 108.025 ;
        RECT 34.375 107.470 34.545 108.195 ;
        RECT 33.655 107.400 34.545 107.470 ;
        RECT 34.715 107.870 34.935 108.355 ;
        RECT 35.105 108.035 35.355 108.575 ;
        RECT 35.525 107.925 35.785 108.405 ;
        RECT 34.715 107.445 35.045 107.870 ;
        RECT 33.655 107.375 34.550 107.400 ;
        RECT 33.655 107.360 34.560 107.375 ;
        RECT 33.655 107.345 34.565 107.360 ;
        RECT 33.655 107.340 34.575 107.345 ;
        RECT 33.655 107.330 34.580 107.340 ;
        RECT 33.655 107.320 34.585 107.330 ;
        RECT 33.655 107.315 34.595 107.320 ;
        RECT 33.655 107.305 34.605 107.315 ;
        RECT 33.655 107.300 34.615 107.305 ;
        RECT 33.655 106.850 33.915 107.300 ;
        RECT 34.280 107.295 34.615 107.300 ;
        RECT 34.280 107.290 34.630 107.295 ;
        RECT 34.280 107.280 34.645 107.290 ;
        RECT 34.280 107.275 34.670 107.280 ;
        RECT 35.215 107.275 35.445 107.670 ;
        RECT 34.280 107.270 35.445 107.275 ;
        RECT 34.310 107.235 35.445 107.270 ;
        RECT 34.345 107.210 35.445 107.235 ;
        RECT 34.375 107.180 35.445 107.210 ;
        RECT 34.395 107.150 35.445 107.180 ;
        RECT 34.415 107.120 35.445 107.150 ;
        RECT 34.485 107.110 35.445 107.120 ;
        RECT 34.510 107.100 35.445 107.110 ;
        RECT 34.530 107.085 35.445 107.100 ;
        RECT 34.550 107.070 35.445 107.085 ;
        RECT 34.555 107.060 35.340 107.070 ;
        RECT 34.570 107.025 35.340 107.060 ;
        RECT 34.085 106.705 34.415 106.950 ;
        RECT 34.585 106.775 35.340 107.025 ;
        RECT 35.615 106.895 35.785 107.925 ;
        RECT 34.085 106.680 34.270 106.705 ;
        RECT 33.655 106.580 34.270 106.680 ;
        RECT 27.675 106.025 33.020 106.460 ;
        RECT 33.655 106.025 34.260 106.580 ;
        RECT 34.435 106.195 34.915 106.535 ;
        RECT 35.085 106.025 35.340 106.570 ;
        RECT 35.510 106.195 35.785 106.895 ;
        RECT 35.965 106.205 36.225 108.395 ;
        RECT 36.485 108.205 37.155 108.575 ;
        RECT 37.335 108.025 37.645 108.395 ;
        RECT 36.415 107.825 37.645 108.025 ;
        RECT 36.415 107.155 36.705 107.825 ;
        RECT 37.825 107.645 38.055 108.285 ;
        RECT 38.235 107.845 38.525 108.575 ;
        RECT 39.175 107.850 39.465 108.575 ;
        RECT 39.635 107.775 40.330 108.405 ;
        RECT 40.535 107.775 40.845 108.575 ;
        RECT 41.015 107.805 43.605 108.575 ;
        RECT 44.435 107.945 44.765 108.305 ;
        RECT 45.385 108.115 45.635 108.575 ;
        RECT 45.805 108.115 46.365 108.405 ;
        RECT 36.885 107.335 37.350 107.645 ;
        RECT 37.530 107.335 38.055 107.645 ;
        RECT 38.235 107.335 38.535 107.665 ;
        RECT 39.655 107.335 39.990 107.585 ;
        RECT 36.415 106.935 37.185 107.155 ;
        RECT 36.395 106.025 36.735 106.755 ;
        RECT 36.915 106.205 37.185 106.935 ;
        RECT 37.365 106.915 38.525 107.155 ;
        RECT 37.365 106.205 37.595 106.915 ;
        RECT 37.765 106.025 38.095 106.735 ;
        RECT 38.265 106.205 38.525 106.915 ;
        RECT 39.175 106.025 39.465 107.190 ;
        RECT 40.160 107.175 40.330 107.775 ;
        RECT 40.500 107.335 40.835 107.605 ;
        RECT 41.015 107.285 42.225 107.805 ;
        RECT 44.435 107.755 45.825 107.945 ;
        RECT 45.655 107.665 45.825 107.755 ;
        RECT 39.635 106.025 39.895 107.165 ;
        RECT 40.065 106.195 40.395 107.175 ;
        RECT 40.565 106.025 40.845 107.165 ;
        RECT 42.395 107.115 43.605 107.635 ;
        RECT 41.015 106.025 43.605 107.115 ;
        RECT 44.250 107.335 44.925 107.585 ;
        RECT 45.145 107.335 45.485 107.585 ;
        RECT 45.655 107.335 45.945 107.665 ;
        RECT 44.250 106.975 44.515 107.335 ;
        RECT 45.655 107.085 45.825 107.335 ;
        RECT 44.885 106.915 45.825 107.085 ;
        RECT 44.435 106.025 44.715 106.695 ;
        RECT 44.885 106.365 45.185 106.915 ;
        RECT 46.115 106.745 46.365 108.115 ;
        RECT 46.815 107.945 47.195 108.395 ;
        RECT 46.555 106.995 46.785 107.685 ;
        RECT 46.965 107.495 47.195 107.945 ;
        RECT 47.375 107.795 47.605 108.575 ;
        RECT 47.785 107.865 48.215 108.395 ;
        RECT 47.785 107.615 48.030 107.865 ;
        RECT 48.395 107.665 48.605 108.285 ;
        RECT 48.775 107.845 49.105 108.575 ;
        RECT 49.410 107.945 49.695 108.405 ;
        RECT 49.865 108.115 50.135 108.575 ;
        RECT 49.410 107.775 50.365 107.945 ;
        RECT 46.965 106.815 47.305 107.495 ;
        RECT 45.385 106.025 45.715 106.745 ;
        RECT 45.905 106.195 46.365 106.745 ;
        RECT 46.545 106.615 47.305 106.815 ;
        RECT 47.495 107.315 48.030 107.615 ;
        RECT 48.210 107.315 48.605 107.665 ;
        RECT 48.800 107.315 49.090 107.665 ;
        RECT 46.545 106.225 46.805 106.615 ;
        RECT 46.975 106.025 47.305 106.435 ;
        RECT 47.495 106.205 47.825 107.315 ;
        RECT 47.995 106.935 49.035 107.135 ;
        RECT 49.295 107.045 49.985 107.605 ;
        RECT 47.995 106.205 48.185 106.935 ;
        RECT 48.355 106.025 48.685 106.755 ;
        RECT 48.865 106.205 49.035 106.935 ;
        RECT 50.155 106.875 50.365 107.775 ;
        RECT 49.410 106.655 50.365 106.875 ;
        RECT 50.535 107.605 50.935 108.405 ;
        RECT 51.125 107.945 51.405 108.405 ;
        RECT 51.925 108.115 52.250 108.575 ;
        RECT 51.125 107.775 52.250 107.945 ;
        RECT 52.420 107.835 52.805 108.405 ;
        RECT 53.140 108.065 53.380 108.575 ;
        RECT 53.560 108.065 53.840 108.395 ;
        RECT 54.070 108.065 54.285 108.575 ;
        RECT 51.800 107.665 52.250 107.775 ;
        RECT 50.535 107.045 51.630 107.605 ;
        RECT 51.800 107.335 52.355 107.665 ;
        RECT 49.410 106.195 49.695 106.655 ;
        RECT 49.865 106.025 50.135 106.485 ;
        RECT 50.535 106.195 50.935 107.045 ;
        RECT 51.800 106.875 52.250 107.335 ;
        RECT 52.525 107.165 52.805 107.835 ;
        RECT 53.035 107.335 53.390 107.895 ;
        RECT 53.560 107.165 53.730 108.065 ;
        RECT 53.900 107.335 54.165 107.895 ;
        RECT 54.455 107.835 55.070 108.405 ;
        RECT 54.415 107.165 54.585 107.665 ;
        RECT 51.125 106.655 52.250 106.875 ;
        RECT 51.125 106.195 51.405 106.655 ;
        RECT 51.925 106.025 52.250 106.485 ;
        RECT 52.420 106.195 52.805 107.165 ;
        RECT 53.160 106.995 54.585 107.165 ;
        RECT 53.160 106.820 53.550 106.995 ;
        RECT 54.035 106.025 54.365 106.825 ;
        RECT 54.755 106.815 55.070 107.835 ;
        RECT 54.535 106.195 55.070 106.815 ;
        RECT 55.275 107.925 55.535 108.405 ;
        RECT 55.705 108.035 55.955 108.575 ;
        RECT 55.275 106.895 55.445 107.925 ;
        RECT 56.125 107.895 56.345 108.355 ;
        RECT 56.095 107.870 56.345 107.895 ;
        RECT 55.615 107.275 55.845 107.670 ;
        RECT 56.015 107.445 56.345 107.870 ;
        RECT 56.515 108.195 57.405 108.365 ;
        RECT 56.515 107.470 56.685 108.195 ;
        RECT 56.855 107.640 57.405 108.025 ;
        RECT 57.575 107.805 61.085 108.575 ;
        RECT 61.260 108.100 61.595 108.360 ;
        RECT 61.765 108.175 62.095 108.575 ;
        RECT 62.265 108.175 63.880 108.345 ;
        RECT 56.515 107.400 57.405 107.470 ;
        RECT 56.510 107.375 57.405 107.400 ;
        RECT 56.500 107.360 57.405 107.375 ;
        RECT 56.495 107.345 57.405 107.360 ;
        RECT 56.485 107.340 57.405 107.345 ;
        RECT 56.480 107.330 57.405 107.340 ;
        RECT 56.475 107.320 57.405 107.330 ;
        RECT 56.465 107.315 57.405 107.320 ;
        RECT 56.455 107.305 57.405 107.315 ;
        RECT 56.445 107.300 57.405 107.305 ;
        RECT 56.445 107.295 56.780 107.300 ;
        RECT 56.430 107.290 56.780 107.295 ;
        RECT 56.415 107.280 56.780 107.290 ;
        RECT 56.390 107.275 56.780 107.280 ;
        RECT 55.615 107.270 56.780 107.275 ;
        RECT 55.615 107.235 56.750 107.270 ;
        RECT 55.615 107.210 56.715 107.235 ;
        RECT 55.615 107.180 56.685 107.210 ;
        RECT 55.615 107.150 56.665 107.180 ;
        RECT 55.615 107.120 56.645 107.150 ;
        RECT 55.615 107.110 56.575 107.120 ;
        RECT 55.615 107.100 56.550 107.110 ;
        RECT 55.615 107.085 56.530 107.100 ;
        RECT 55.615 107.070 56.510 107.085 ;
        RECT 55.720 107.060 56.505 107.070 ;
        RECT 55.720 107.025 56.490 107.060 ;
        RECT 55.275 106.195 55.550 106.895 ;
        RECT 55.720 106.775 56.475 107.025 ;
        RECT 56.645 106.705 56.975 106.950 ;
        RECT 57.145 106.850 57.405 107.300 ;
        RECT 57.575 107.285 59.225 107.805 ;
        RECT 59.395 107.115 61.085 107.635 ;
        RECT 56.790 106.680 56.975 106.705 ;
        RECT 56.790 106.580 57.405 106.680 ;
        RECT 55.720 106.025 55.975 106.570 ;
        RECT 56.145 106.195 56.625 106.535 ;
        RECT 56.800 106.025 57.405 106.580 ;
        RECT 57.575 106.025 61.085 107.115 ;
        RECT 61.260 106.745 61.515 108.100 ;
        RECT 62.265 108.005 62.435 108.175 ;
        RECT 61.875 107.835 62.435 108.005 ;
        RECT 61.875 107.665 62.045 107.835 ;
        RECT 61.740 107.335 62.045 107.665 ;
        RECT 62.240 107.555 62.490 107.665 ;
        RECT 62.700 107.555 62.970 107.995 ;
        RECT 63.160 107.895 63.450 107.995 ;
        RECT 63.155 107.725 63.450 107.895 ;
        RECT 62.235 107.385 62.490 107.555 ;
        RECT 62.695 107.385 62.970 107.555 ;
        RECT 62.240 107.335 62.490 107.385 ;
        RECT 62.700 107.335 62.970 107.385 ;
        RECT 63.160 107.335 63.450 107.725 ;
        RECT 63.620 107.335 64.040 108.000 ;
        RECT 64.425 107.855 64.755 108.575 ;
        RECT 64.935 107.850 65.225 108.575 ;
        RECT 65.395 107.825 66.605 108.575 ;
        RECT 66.775 107.835 67.160 108.405 ;
        RECT 67.330 108.115 67.655 108.575 ;
        RECT 68.175 107.945 68.455 108.405 ;
        RECT 64.350 107.335 64.700 107.665 ;
        RECT 61.875 107.165 62.045 107.335 ;
        RECT 64.495 107.215 64.700 107.335 ;
        RECT 65.395 107.285 65.915 107.825 ;
        RECT 61.875 106.995 64.245 107.165 ;
        RECT 64.495 107.045 64.705 107.215 ;
        RECT 61.260 106.235 61.595 106.745 ;
        RECT 61.845 106.025 62.175 106.825 ;
        RECT 62.420 106.615 63.845 106.785 ;
        RECT 62.420 106.195 62.705 106.615 ;
        RECT 62.960 106.025 63.290 106.445 ;
        RECT 63.515 106.365 63.845 106.615 ;
        RECT 64.075 106.535 64.245 106.995 ;
        RECT 64.505 106.365 64.675 106.865 ;
        RECT 63.515 106.195 64.675 106.365 ;
        RECT 64.935 106.025 65.225 107.190 ;
        RECT 66.085 107.115 66.605 107.655 ;
        RECT 65.395 106.025 66.605 107.115 ;
        RECT 66.775 107.165 67.055 107.835 ;
        RECT 67.330 107.775 68.455 107.945 ;
        RECT 67.330 107.665 67.780 107.775 ;
        RECT 67.225 107.335 67.780 107.665 ;
        RECT 68.645 107.605 69.045 108.405 ;
        RECT 69.445 108.115 69.715 108.575 ;
        RECT 69.885 107.945 70.170 108.405 ;
        RECT 66.775 106.195 67.160 107.165 ;
        RECT 67.330 106.875 67.780 107.335 ;
        RECT 67.950 107.045 69.045 107.605 ;
        RECT 67.330 106.655 68.455 106.875 ;
        RECT 67.330 106.025 67.655 106.485 ;
        RECT 68.175 106.195 68.455 106.655 ;
        RECT 68.645 106.195 69.045 107.045 ;
        RECT 69.215 107.775 70.170 107.945 ;
        RECT 70.455 107.805 73.965 108.575 ;
        RECT 74.225 108.025 74.395 108.315 ;
        RECT 74.565 108.195 74.895 108.575 ;
        RECT 74.225 107.855 74.890 108.025 ;
        RECT 69.215 106.875 69.425 107.775 ;
        RECT 69.595 107.045 70.285 107.605 ;
        RECT 70.455 107.285 72.105 107.805 ;
        RECT 72.275 107.115 73.965 107.635 ;
        RECT 69.215 106.655 70.170 106.875 ;
        RECT 69.445 106.025 69.715 106.485 ;
        RECT 69.885 106.195 70.170 106.655 ;
        RECT 70.455 106.025 73.965 107.115 ;
        RECT 74.140 107.035 74.490 107.685 ;
        RECT 74.660 106.865 74.890 107.855 ;
        RECT 74.225 106.695 74.890 106.865 ;
        RECT 74.225 106.195 74.395 106.695 ;
        RECT 74.565 106.025 74.895 106.525 ;
        RECT 75.065 106.195 75.250 108.315 ;
        RECT 75.505 108.115 75.755 108.575 ;
        RECT 75.925 108.125 76.260 108.295 ;
        RECT 76.455 108.125 77.130 108.295 ;
        RECT 75.925 107.985 76.095 108.125 ;
        RECT 75.420 106.995 75.700 107.945 ;
        RECT 75.870 107.855 76.095 107.985 ;
        RECT 75.870 106.750 76.040 107.855 ;
        RECT 76.265 107.705 76.790 107.925 ;
        RECT 76.210 106.940 76.450 107.535 ;
        RECT 76.620 107.005 76.790 107.705 ;
        RECT 76.960 107.345 77.130 108.125 ;
        RECT 77.450 108.075 77.820 108.575 ;
        RECT 78.000 108.125 78.405 108.295 ;
        RECT 78.575 108.125 79.360 108.295 ;
        RECT 78.000 107.895 78.170 108.125 ;
        RECT 77.340 107.595 78.170 107.895 ;
        RECT 78.555 107.625 79.020 107.955 ;
        RECT 77.340 107.565 77.540 107.595 ;
        RECT 77.660 107.345 77.830 107.415 ;
        RECT 76.960 107.175 77.830 107.345 ;
        RECT 77.320 107.085 77.830 107.175 ;
        RECT 75.870 106.620 76.175 106.750 ;
        RECT 76.620 106.640 77.150 107.005 ;
        RECT 75.490 106.025 75.755 106.485 ;
        RECT 75.925 106.195 76.175 106.620 ;
        RECT 77.320 106.470 77.490 107.085 ;
        RECT 76.385 106.300 77.490 106.470 ;
        RECT 77.660 106.025 77.830 106.825 ;
        RECT 78.000 106.525 78.170 107.595 ;
        RECT 78.340 106.695 78.530 107.415 ;
        RECT 78.700 106.665 79.020 107.625 ;
        RECT 79.190 107.665 79.360 108.125 ;
        RECT 79.635 108.045 79.845 108.575 ;
        RECT 80.105 107.835 80.435 108.360 ;
        RECT 80.605 107.965 80.775 108.575 ;
        RECT 80.945 107.920 81.275 108.355 ;
        RECT 80.945 107.835 81.325 107.920 ;
        RECT 80.235 107.665 80.435 107.835 ;
        RECT 81.100 107.795 81.325 107.835 ;
        RECT 79.190 107.335 80.065 107.665 ;
        RECT 80.235 107.335 80.985 107.665 ;
        RECT 78.000 106.195 78.250 106.525 ;
        RECT 79.190 106.495 79.360 107.335 ;
        RECT 80.235 107.130 80.425 107.335 ;
        RECT 81.155 107.215 81.325 107.795 ;
        RECT 81.495 107.805 85.005 108.575 ;
        RECT 81.495 107.285 83.145 107.805 ;
        RECT 85.635 107.775 85.975 108.405 ;
        RECT 86.145 107.775 86.395 108.575 ;
        RECT 86.585 107.925 86.915 108.405 ;
        RECT 87.085 108.115 87.310 108.575 ;
        RECT 87.480 107.925 87.810 108.405 ;
        RECT 81.110 107.165 81.325 107.215 ;
        RECT 79.530 106.755 80.425 107.130 ;
        RECT 80.935 107.085 81.325 107.165 ;
        RECT 83.315 107.115 85.005 107.635 ;
        RECT 78.475 106.325 79.360 106.495 ;
        RECT 79.540 106.025 79.855 106.525 ;
        RECT 80.085 106.195 80.425 106.755 ;
        RECT 80.595 106.025 80.765 107.035 ;
        RECT 80.935 106.240 81.265 107.085 ;
        RECT 81.495 106.025 85.005 107.115 ;
        RECT 85.635 107.165 85.810 107.775 ;
        RECT 86.585 107.755 87.810 107.925 ;
        RECT 88.440 107.795 88.940 108.405 ;
        RECT 89.315 107.825 90.525 108.575 ;
        RECT 90.695 107.850 90.985 108.575 ;
        RECT 91.155 108.075 91.415 108.405 ;
        RECT 91.585 108.215 91.915 108.575 ;
        RECT 92.170 108.195 93.470 108.405 ;
        RECT 91.155 108.065 91.385 108.075 ;
        RECT 85.980 107.415 86.675 107.585 ;
        RECT 86.505 107.165 86.675 107.415 ;
        RECT 86.850 107.385 87.270 107.585 ;
        RECT 87.440 107.385 87.770 107.585 ;
        RECT 87.940 107.385 88.270 107.585 ;
        RECT 88.440 107.165 88.610 107.795 ;
        RECT 88.795 107.335 89.145 107.585 ;
        RECT 89.315 107.285 89.835 107.825 ;
        RECT 85.635 106.195 85.975 107.165 ;
        RECT 86.145 106.025 86.315 107.165 ;
        RECT 86.505 106.995 88.940 107.165 ;
        RECT 90.005 107.115 90.525 107.655 ;
        RECT 86.585 106.025 86.835 106.825 ;
        RECT 87.480 106.195 87.810 106.995 ;
        RECT 88.110 106.025 88.440 106.825 ;
        RECT 88.610 106.195 88.940 106.995 ;
        RECT 89.315 106.025 90.525 107.115 ;
        RECT 90.695 106.025 90.985 107.190 ;
        RECT 91.155 106.875 91.325 108.065 ;
        RECT 92.170 108.045 92.340 108.195 ;
        RECT 91.585 107.920 92.340 108.045 ;
        RECT 91.495 107.875 92.340 107.920 ;
        RECT 91.495 107.755 91.765 107.875 ;
        RECT 91.495 107.180 91.665 107.755 ;
        RECT 91.895 107.315 92.305 107.620 ;
        RECT 92.595 107.585 92.805 107.985 ;
        RECT 92.475 107.375 92.805 107.585 ;
        RECT 93.050 107.585 93.270 107.985 ;
        RECT 93.745 107.810 94.200 108.575 ;
        RECT 94.375 108.030 99.720 108.575 ;
        RECT 93.050 107.375 93.525 107.585 ;
        RECT 93.715 107.385 94.205 107.585 ;
        RECT 91.495 107.145 91.695 107.180 ;
        RECT 93.025 107.145 94.200 107.205 ;
        RECT 95.960 107.200 96.300 108.030 ;
        RECT 99.895 107.805 102.485 108.575 ;
        RECT 103.205 108.025 103.375 108.315 ;
        RECT 103.545 108.195 103.875 108.575 ;
        RECT 103.205 107.855 103.870 108.025 ;
        RECT 91.495 107.035 94.200 107.145 ;
        RECT 91.555 106.975 93.355 107.035 ;
        RECT 93.025 106.945 93.355 106.975 ;
        RECT 91.155 106.195 91.415 106.875 ;
        RECT 91.585 106.025 91.835 106.805 ;
        RECT 92.085 106.775 92.920 106.785 ;
        RECT 93.510 106.775 93.695 106.865 ;
        RECT 92.085 106.575 93.695 106.775 ;
        RECT 92.085 106.195 92.335 106.575 ;
        RECT 93.465 106.535 93.695 106.575 ;
        RECT 93.945 106.415 94.200 107.035 ;
        RECT 97.780 106.460 98.130 107.710 ;
        RECT 99.895 107.285 101.105 107.805 ;
        RECT 101.275 107.115 102.485 107.635 ;
        RECT 92.505 106.025 92.860 106.405 ;
        RECT 93.865 106.195 94.200 106.415 ;
        RECT 94.375 106.025 99.720 106.460 ;
        RECT 99.895 106.025 102.485 107.115 ;
        RECT 103.120 107.035 103.470 107.685 ;
        RECT 103.640 106.865 103.870 107.855 ;
        RECT 103.205 106.695 103.870 106.865 ;
        RECT 103.205 106.195 103.375 106.695 ;
        RECT 103.545 106.025 103.875 106.525 ;
        RECT 104.045 106.195 104.230 108.315 ;
        RECT 104.485 108.115 104.735 108.575 ;
        RECT 104.905 108.125 105.240 108.295 ;
        RECT 105.435 108.125 106.110 108.295 ;
        RECT 104.905 107.985 105.075 108.125 ;
        RECT 104.400 106.995 104.680 107.945 ;
        RECT 104.850 107.855 105.075 107.985 ;
        RECT 104.850 106.750 105.020 107.855 ;
        RECT 105.245 107.705 105.770 107.925 ;
        RECT 105.190 106.940 105.430 107.535 ;
        RECT 105.600 107.005 105.770 107.705 ;
        RECT 105.940 107.345 106.110 108.125 ;
        RECT 106.430 108.075 106.800 108.575 ;
        RECT 106.980 108.125 107.385 108.295 ;
        RECT 107.555 108.125 108.340 108.295 ;
        RECT 106.980 107.895 107.150 108.125 ;
        RECT 106.320 107.595 107.150 107.895 ;
        RECT 107.535 107.625 108.000 107.955 ;
        RECT 106.320 107.565 106.520 107.595 ;
        RECT 106.640 107.345 106.810 107.415 ;
        RECT 105.940 107.175 106.810 107.345 ;
        RECT 106.300 107.085 106.810 107.175 ;
        RECT 104.850 106.620 105.155 106.750 ;
        RECT 105.600 106.640 106.130 107.005 ;
        RECT 104.470 106.025 104.735 106.485 ;
        RECT 104.905 106.195 105.155 106.620 ;
        RECT 106.300 106.470 106.470 107.085 ;
        RECT 105.365 106.300 106.470 106.470 ;
        RECT 106.640 106.025 106.810 106.825 ;
        RECT 106.980 106.525 107.150 107.595 ;
        RECT 107.320 106.695 107.510 107.415 ;
        RECT 107.680 106.665 108.000 107.625 ;
        RECT 108.170 107.665 108.340 108.125 ;
        RECT 108.615 108.045 108.825 108.575 ;
        RECT 109.085 107.835 109.415 108.360 ;
        RECT 109.585 107.965 109.755 108.575 ;
        RECT 109.925 107.920 110.255 108.355 ;
        RECT 109.925 107.835 110.305 107.920 ;
        RECT 109.215 107.665 109.415 107.835 ;
        RECT 110.080 107.795 110.305 107.835 ;
        RECT 108.170 107.335 109.045 107.665 ;
        RECT 109.215 107.335 109.965 107.665 ;
        RECT 106.980 106.195 107.230 106.525 ;
        RECT 108.170 106.495 108.340 107.335 ;
        RECT 109.215 107.130 109.405 107.335 ;
        RECT 110.135 107.215 110.305 107.795 ;
        RECT 110.475 107.805 113.065 108.575 ;
        RECT 113.895 107.945 114.225 108.305 ;
        RECT 114.845 108.115 115.095 108.575 ;
        RECT 115.265 108.115 115.825 108.405 ;
        RECT 110.475 107.285 111.685 107.805 ;
        RECT 113.895 107.755 115.285 107.945 ;
        RECT 115.115 107.665 115.285 107.755 ;
        RECT 110.090 107.165 110.305 107.215 ;
        RECT 108.510 106.755 109.405 107.130 ;
        RECT 109.915 107.085 110.305 107.165 ;
        RECT 111.855 107.115 113.065 107.635 ;
        RECT 107.455 106.325 108.340 106.495 ;
        RECT 108.520 106.025 108.835 106.525 ;
        RECT 109.065 106.195 109.405 106.755 ;
        RECT 109.575 106.025 109.745 107.035 ;
        RECT 109.915 106.240 110.245 107.085 ;
        RECT 110.475 106.025 113.065 107.115 ;
        RECT 113.710 107.335 114.385 107.585 ;
        RECT 114.605 107.335 114.945 107.585 ;
        RECT 115.115 107.335 115.405 107.665 ;
        RECT 113.710 106.975 113.975 107.335 ;
        RECT 115.115 107.085 115.285 107.335 ;
        RECT 114.345 106.915 115.285 107.085 ;
        RECT 113.895 106.025 114.175 106.695 ;
        RECT 114.345 106.365 114.645 106.915 ;
        RECT 115.575 106.745 115.825 108.115 ;
        RECT 116.455 107.850 116.745 108.575 ;
        RECT 116.915 108.030 122.260 108.575 ;
        RECT 118.500 107.200 118.840 108.030 ;
        RECT 122.640 107.795 123.140 108.405 ;
        RECT 114.845 106.025 115.175 106.745 ;
        RECT 115.365 106.195 115.825 106.745 ;
        RECT 116.455 106.025 116.745 107.190 ;
        RECT 120.320 106.460 120.670 107.710 ;
        RECT 122.435 107.335 122.785 107.585 ;
        RECT 122.970 107.165 123.140 107.795 ;
        RECT 123.770 107.925 124.100 108.405 ;
        RECT 124.270 108.115 124.495 108.575 ;
        RECT 124.665 107.925 124.995 108.405 ;
        RECT 123.770 107.755 124.995 107.925 ;
        RECT 125.185 107.775 125.435 108.575 ;
        RECT 125.605 107.775 125.945 108.405 ;
        RECT 126.205 108.025 126.375 108.315 ;
        RECT 126.545 108.195 126.875 108.575 ;
        RECT 126.205 107.855 126.870 108.025 ;
        RECT 125.715 107.725 125.945 107.775 ;
        RECT 123.310 107.385 123.640 107.585 ;
        RECT 123.810 107.385 124.140 107.585 ;
        RECT 124.310 107.385 124.730 107.585 ;
        RECT 124.905 107.415 125.600 107.585 ;
        RECT 124.905 107.165 125.075 107.415 ;
        RECT 125.770 107.165 125.945 107.725 ;
        RECT 122.640 106.995 125.075 107.165 ;
        RECT 116.915 106.025 122.260 106.460 ;
        RECT 122.640 106.195 122.970 106.995 ;
        RECT 123.140 106.025 123.470 106.825 ;
        RECT 123.770 106.195 124.100 106.995 ;
        RECT 124.745 106.025 124.995 106.825 ;
        RECT 125.265 106.025 125.435 107.165 ;
        RECT 125.605 106.195 125.945 107.165 ;
        RECT 126.120 107.035 126.470 107.685 ;
        RECT 126.640 106.865 126.870 107.855 ;
        RECT 126.205 106.695 126.870 106.865 ;
        RECT 126.205 106.195 126.375 106.695 ;
        RECT 126.545 106.025 126.875 106.525 ;
        RECT 127.045 106.195 127.230 108.315 ;
        RECT 127.485 108.115 127.735 108.575 ;
        RECT 127.905 108.125 128.240 108.295 ;
        RECT 128.435 108.125 129.110 108.295 ;
        RECT 127.905 107.985 128.075 108.125 ;
        RECT 127.400 106.995 127.680 107.945 ;
        RECT 127.850 107.855 128.075 107.985 ;
        RECT 127.850 106.750 128.020 107.855 ;
        RECT 128.245 107.705 128.770 107.925 ;
        RECT 128.190 106.940 128.430 107.535 ;
        RECT 128.600 107.005 128.770 107.705 ;
        RECT 128.940 107.345 129.110 108.125 ;
        RECT 129.430 108.075 129.800 108.575 ;
        RECT 129.980 108.125 130.385 108.295 ;
        RECT 130.555 108.125 131.340 108.295 ;
        RECT 129.980 107.895 130.150 108.125 ;
        RECT 129.320 107.595 130.150 107.895 ;
        RECT 130.535 107.625 131.000 107.955 ;
        RECT 129.320 107.565 129.520 107.595 ;
        RECT 129.640 107.345 129.810 107.415 ;
        RECT 128.940 107.175 129.810 107.345 ;
        RECT 129.300 107.085 129.810 107.175 ;
        RECT 127.850 106.620 128.155 106.750 ;
        RECT 128.600 106.640 129.130 107.005 ;
        RECT 127.470 106.025 127.735 106.485 ;
        RECT 127.905 106.195 128.155 106.620 ;
        RECT 129.300 106.470 129.470 107.085 ;
        RECT 128.365 106.300 129.470 106.470 ;
        RECT 129.640 106.025 129.810 106.825 ;
        RECT 129.980 106.525 130.150 107.595 ;
        RECT 130.320 106.695 130.510 107.415 ;
        RECT 130.680 106.665 131.000 107.625 ;
        RECT 131.170 107.665 131.340 108.125 ;
        RECT 131.615 108.045 131.825 108.575 ;
        RECT 132.085 107.835 132.415 108.360 ;
        RECT 132.585 107.965 132.755 108.575 ;
        RECT 132.925 107.920 133.255 108.355 ;
        RECT 133.475 108.075 133.735 108.405 ;
        RECT 133.905 108.215 134.235 108.575 ;
        RECT 134.490 108.195 135.790 108.405 ;
        RECT 132.925 107.835 133.305 107.920 ;
        RECT 132.215 107.665 132.415 107.835 ;
        RECT 133.080 107.795 133.305 107.835 ;
        RECT 131.170 107.335 132.045 107.665 ;
        RECT 132.215 107.335 132.965 107.665 ;
        RECT 129.980 106.195 130.230 106.525 ;
        RECT 131.170 106.495 131.340 107.335 ;
        RECT 132.215 107.130 132.405 107.335 ;
        RECT 133.135 107.215 133.305 107.795 ;
        RECT 133.090 107.165 133.305 107.215 ;
        RECT 131.510 106.755 132.405 107.130 ;
        RECT 132.915 107.085 133.305 107.165 ;
        RECT 130.455 106.325 131.340 106.495 ;
        RECT 131.520 106.025 131.835 106.525 ;
        RECT 132.065 106.195 132.405 106.755 ;
        RECT 132.575 106.025 132.745 107.035 ;
        RECT 132.915 106.240 133.245 107.085 ;
        RECT 133.475 106.875 133.645 108.075 ;
        RECT 134.490 108.045 134.660 108.195 ;
        RECT 133.905 107.920 134.660 108.045 ;
        RECT 133.815 107.875 134.660 107.920 ;
        RECT 133.815 107.755 134.085 107.875 ;
        RECT 133.815 107.180 133.985 107.755 ;
        RECT 134.215 107.315 134.625 107.620 ;
        RECT 134.915 107.585 135.125 107.985 ;
        RECT 134.795 107.375 135.125 107.585 ;
        RECT 135.370 107.585 135.590 107.985 ;
        RECT 136.065 107.810 136.520 108.575 ;
        RECT 137.615 107.825 138.825 108.575 ;
        RECT 135.370 107.375 135.845 107.585 ;
        RECT 136.035 107.385 136.525 107.585 ;
        RECT 133.815 107.145 134.015 107.180 ;
        RECT 135.345 107.145 136.520 107.205 ;
        RECT 133.815 107.035 136.520 107.145 ;
        RECT 133.875 106.975 135.675 107.035 ;
        RECT 135.345 106.945 135.675 106.975 ;
        RECT 133.475 106.195 133.735 106.875 ;
        RECT 133.905 106.025 134.155 106.805 ;
        RECT 134.405 106.775 135.240 106.785 ;
        RECT 135.830 106.775 136.015 106.865 ;
        RECT 134.405 106.575 136.015 106.775 ;
        RECT 134.405 106.195 134.655 106.575 ;
        RECT 135.785 106.535 136.015 106.575 ;
        RECT 136.265 106.415 136.520 107.035 ;
        RECT 134.825 106.025 135.180 106.405 ;
        RECT 136.185 106.195 136.520 106.415 ;
        RECT 137.615 107.115 138.135 107.655 ;
        RECT 138.305 107.285 138.825 107.825 ;
        RECT 137.615 106.025 138.825 107.115 ;
        RECT 13.330 105.855 138.910 106.025 ;
        RECT 13.415 104.765 14.625 105.855 ;
        RECT 14.795 105.420 20.140 105.855 ;
        RECT 13.415 104.055 13.935 104.595 ;
        RECT 14.105 104.225 14.625 104.765 ;
        RECT 13.415 103.305 14.625 104.055 ;
        RECT 16.380 103.850 16.720 104.680 ;
        RECT 18.200 104.170 18.550 105.420 ;
        RECT 20.315 104.765 21.985 105.855 ;
        RECT 20.315 104.075 21.065 104.595 ;
        RECT 21.235 104.245 21.985 104.765 ;
        RECT 22.340 104.885 22.730 105.060 ;
        RECT 23.215 105.055 23.545 105.855 ;
        RECT 23.715 105.065 24.250 105.685 ;
        RECT 22.340 104.715 23.765 104.885 ;
        RECT 14.795 103.305 20.140 103.850 ;
        RECT 20.315 103.305 21.985 104.075 ;
        RECT 22.215 103.985 22.570 104.545 ;
        RECT 22.740 103.815 22.910 104.715 ;
        RECT 23.080 103.985 23.345 104.545 ;
        RECT 23.595 104.215 23.765 104.715 ;
        RECT 23.935 104.045 24.250 105.065 ;
        RECT 24.455 104.765 26.125 105.855 ;
        RECT 22.320 103.305 22.560 103.815 ;
        RECT 22.740 103.485 23.020 103.815 ;
        RECT 23.250 103.305 23.465 103.815 ;
        RECT 23.635 103.475 24.250 104.045 ;
        RECT 24.455 104.075 25.205 104.595 ;
        RECT 25.375 104.245 26.125 104.765 ;
        RECT 26.295 104.690 26.585 105.855 ;
        RECT 26.755 104.765 30.265 105.855 ;
        RECT 30.435 104.765 31.645 105.855 ;
        RECT 26.755 104.075 28.405 104.595 ;
        RECT 28.575 104.245 30.265 104.765 ;
        RECT 24.455 103.305 26.125 104.075 ;
        RECT 26.295 103.305 26.585 104.030 ;
        RECT 26.755 103.305 30.265 104.075 ;
        RECT 30.435 104.055 30.955 104.595 ;
        RECT 31.125 104.225 31.645 104.765 ;
        RECT 31.850 105.065 32.385 105.685 ;
        RECT 30.435 103.305 31.645 104.055 ;
        RECT 31.850 104.045 32.165 105.065 ;
        RECT 32.555 105.055 32.885 105.855 ;
        RECT 34.205 105.185 34.375 105.685 ;
        RECT 34.545 105.355 34.875 105.855 ;
        RECT 33.370 104.885 33.760 105.060 ;
        RECT 34.205 105.015 34.870 105.185 ;
        RECT 32.335 104.715 33.760 104.885 ;
        RECT 32.335 104.215 32.505 104.715 ;
        RECT 31.850 103.475 32.465 104.045 ;
        RECT 32.755 103.985 33.020 104.545 ;
        RECT 33.190 103.815 33.360 104.715 ;
        RECT 33.530 103.985 33.885 104.545 ;
        RECT 34.120 104.195 34.470 104.845 ;
        RECT 34.640 104.025 34.870 105.015 ;
        RECT 34.205 103.855 34.870 104.025 ;
        RECT 32.635 103.305 32.850 103.815 ;
        RECT 33.080 103.485 33.360 103.815 ;
        RECT 33.540 103.305 33.780 103.815 ;
        RECT 34.205 103.565 34.375 103.855 ;
        RECT 34.545 103.305 34.875 103.685 ;
        RECT 35.045 103.565 35.230 105.685 ;
        RECT 35.470 105.395 35.735 105.855 ;
        RECT 35.905 105.260 36.155 105.685 ;
        RECT 36.365 105.410 37.470 105.580 ;
        RECT 35.850 105.130 36.155 105.260 ;
        RECT 35.400 103.935 35.680 104.885 ;
        RECT 35.850 104.025 36.020 105.130 ;
        RECT 36.190 104.345 36.430 104.940 ;
        RECT 36.600 104.875 37.130 105.240 ;
        RECT 36.600 104.175 36.770 104.875 ;
        RECT 37.300 104.795 37.470 105.410 ;
        RECT 37.640 105.055 37.810 105.855 ;
        RECT 37.980 105.355 38.230 105.685 ;
        RECT 38.455 105.385 39.340 105.555 ;
        RECT 37.300 104.705 37.810 104.795 ;
        RECT 35.850 103.895 36.075 104.025 ;
        RECT 36.245 103.955 36.770 104.175 ;
        RECT 36.940 104.535 37.810 104.705 ;
        RECT 35.485 103.305 35.735 103.765 ;
        RECT 35.905 103.755 36.075 103.895 ;
        RECT 36.940 103.755 37.110 104.535 ;
        RECT 37.640 104.465 37.810 104.535 ;
        RECT 37.320 104.285 37.520 104.315 ;
        RECT 37.980 104.285 38.150 105.355 ;
        RECT 38.320 104.465 38.510 105.185 ;
        RECT 37.320 103.985 38.150 104.285 ;
        RECT 38.680 104.255 39.000 105.215 ;
        RECT 35.905 103.585 36.240 103.755 ;
        RECT 36.435 103.585 37.110 103.755 ;
        RECT 37.430 103.305 37.800 103.805 ;
        RECT 37.980 103.755 38.150 103.985 ;
        RECT 38.535 103.925 39.000 104.255 ;
        RECT 39.170 104.545 39.340 105.385 ;
        RECT 39.520 105.355 39.835 105.855 ;
        RECT 40.065 105.125 40.405 105.685 ;
        RECT 39.510 104.750 40.405 105.125 ;
        RECT 40.575 104.845 40.745 105.855 ;
        RECT 40.215 104.545 40.405 104.750 ;
        RECT 40.915 104.795 41.245 105.640 ;
        RECT 41.535 104.795 41.865 105.640 ;
        RECT 42.035 104.845 42.205 105.855 ;
        RECT 42.375 105.125 42.715 105.685 ;
        RECT 42.945 105.355 43.260 105.855 ;
        RECT 43.440 105.385 44.325 105.555 ;
        RECT 40.915 104.715 41.305 104.795 ;
        RECT 41.090 104.665 41.305 104.715 ;
        RECT 39.170 104.215 40.045 104.545 ;
        RECT 40.215 104.215 40.965 104.545 ;
        RECT 39.170 103.755 39.340 104.215 ;
        RECT 40.215 104.045 40.415 104.215 ;
        RECT 41.135 104.085 41.305 104.665 ;
        RECT 41.080 104.045 41.305 104.085 ;
        RECT 37.980 103.585 38.385 103.755 ;
        RECT 38.555 103.585 39.340 103.755 ;
        RECT 39.615 103.305 39.825 103.835 ;
        RECT 40.085 103.520 40.415 104.045 ;
        RECT 40.925 103.960 41.305 104.045 ;
        RECT 41.475 104.715 41.865 104.795 ;
        RECT 42.375 104.750 43.270 105.125 ;
        RECT 41.475 104.665 41.690 104.715 ;
        RECT 41.475 104.085 41.645 104.665 ;
        RECT 42.375 104.545 42.565 104.750 ;
        RECT 43.440 104.545 43.610 105.385 ;
        RECT 44.550 105.355 44.800 105.685 ;
        RECT 41.815 104.215 42.565 104.545 ;
        RECT 42.735 104.215 43.610 104.545 ;
        RECT 41.475 104.045 41.700 104.085 ;
        RECT 42.365 104.045 42.565 104.215 ;
        RECT 41.475 103.960 41.855 104.045 ;
        RECT 40.585 103.305 40.755 103.915 ;
        RECT 40.925 103.525 41.255 103.960 ;
        RECT 41.525 103.525 41.855 103.960 ;
        RECT 42.025 103.305 42.195 103.915 ;
        RECT 42.365 103.520 42.695 104.045 ;
        RECT 42.955 103.305 43.165 103.835 ;
        RECT 43.440 103.755 43.610 104.215 ;
        RECT 43.780 104.255 44.100 105.215 ;
        RECT 44.270 104.465 44.460 105.185 ;
        RECT 44.630 104.285 44.800 105.355 ;
        RECT 44.970 105.055 45.140 105.855 ;
        RECT 45.310 105.410 46.415 105.580 ;
        RECT 45.310 104.795 45.480 105.410 ;
        RECT 46.625 105.260 46.875 105.685 ;
        RECT 47.045 105.395 47.310 105.855 ;
        RECT 45.650 104.875 46.180 105.240 ;
        RECT 46.625 105.130 46.930 105.260 ;
        RECT 44.970 104.705 45.480 104.795 ;
        RECT 44.970 104.535 45.840 104.705 ;
        RECT 44.970 104.465 45.140 104.535 ;
        RECT 45.260 104.285 45.460 104.315 ;
        RECT 43.780 103.925 44.245 104.255 ;
        RECT 44.630 103.985 45.460 104.285 ;
        RECT 44.630 103.755 44.800 103.985 ;
        RECT 43.440 103.585 44.225 103.755 ;
        RECT 44.395 103.585 44.800 103.755 ;
        RECT 44.980 103.305 45.350 103.805 ;
        RECT 45.670 103.755 45.840 104.535 ;
        RECT 46.010 104.175 46.180 104.875 ;
        RECT 46.350 104.345 46.590 104.940 ;
        RECT 46.010 103.955 46.535 104.175 ;
        RECT 46.760 104.025 46.930 105.130 ;
        RECT 46.705 103.895 46.930 104.025 ;
        RECT 47.100 103.935 47.380 104.885 ;
        RECT 46.705 103.755 46.875 103.895 ;
        RECT 45.670 103.585 46.345 103.755 ;
        RECT 46.540 103.585 46.875 103.755 ;
        RECT 47.045 103.305 47.295 103.765 ;
        RECT 47.550 103.565 47.735 105.685 ;
        RECT 47.905 105.355 48.235 105.855 ;
        RECT 48.405 105.185 48.575 105.685 ;
        RECT 48.835 105.345 49.095 105.855 ;
        RECT 47.910 105.015 48.575 105.185 ;
        RECT 47.910 104.025 48.140 105.015 ;
        RECT 48.310 104.195 48.660 104.845 ;
        RECT 48.835 104.295 49.175 105.175 ;
        RECT 49.345 104.465 49.515 105.685 ;
        RECT 49.755 105.350 50.370 105.855 ;
        RECT 49.755 104.815 50.005 105.180 ;
        RECT 50.175 105.175 50.370 105.350 ;
        RECT 50.540 105.345 51.015 105.685 ;
        RECT 51.185 105.310 51.400 105.855 ;
        RECT 50.175 104.985 50.505 105.175 ;
        RECT 50.725 104.815 51.440 105.110 ;
        RECT 51.610 104.985 51.885 105.685 ;
        RECT 49.755 104.645 51.545 104.815 ;
        RECT 49.345 104.215 50.140 104.465 ;
        RECT 49.345 104.125 49.595 104.215 ;
        RECT 47.910 103.855 48.575 104.025 ;
        RECT 47.905 103.305 48.235 103.685 ;
        RECT 48.405 103.565 48.575 103.855 ;
        RECT 48.835 103.305 49.095 104.125 ;
        RECT 49.265 103.705 49.595 104.125 ;
        RECT 50.310 103.790 50.565 104.645 ;
        RECT 49.775 103.525 50.565 103.790 ;
        RECT 50.735 103.945 51.145 104.465 ;
        RECT 51.315 104.215 51.545 104.645 ;
        RECT 51.715 103.955 51.885 104.985 ;
        RECT 52.055 104.690 52.345 105.855 ;
        RECT 52.575 104.795 52.905 105.640 ;
        RECT 53.075 104.845 53.245 105.855 ;
        RECT 53.415 105.125 53.755 105.685 ;
        RECT 53.985 105.355 54.300 105.855 ;
        RECT 54.480 105.385 55.365 105.555 ;
        RECT 52.515 104.715 52.905 104.795 ;
        RECT 53.415 104.750 54.310 105.125 ;
        RECT 52.515 104.665 52.730 104.715 ;
        RECT 52.515 104.085 52.685 104.665 ;
        RECT 53.415 104.545 53.605 104.750 ;
        RECT 54.480 104.545 54.650 105.385 ;
        RECT 55.590 105.355 55.840 105.685 ;
        RECT 52.855 104.215 53.605 104.545 ;
        RECT 53.775 104.215 54.650 104.545 ;
        RECT 52.515 104.045 52.740 104.085 ;
        RECT 53.405 104.045 53.605 104.215 ;
        RECT 50.735 103.525 50.935 103.945 ;
        RECT 51.125 103.305 51.455 103.765 ;
        RECT 51.625 103.475 51.885 103.955 ;
        RECT 52.055 103.305 52.345 104.030 ;
        RECT 52.515 103.960 52.895 104.045 ;
        RECT 52.565 103.525 52.895 103.960 ;
        RECT 53.065 103.305 53.235 103.915 ;
        RECT 53.405 103.520 53.735 104.045 ;
        RECT 53.995 103.305 54.205 103.835 ;
        RECT 54.480 103.755 54.650 104.215 ;
        RECT 54.820 104.255 55.140 105.215 ;
        RECT 55.310 104.465 55.500 105.185 ;
        RECT 55.670 104.285 55.840 105.355 ;
        RECT 56.010 105.055 56.180 105.855 ;
        RECT 56.350 105.410 57.455 105.580 ;
        RECT 56.350 104.795 56.520 105.410 ;
        RECT 57.665 105.260 57.915 105.685 ;
        RECT 58.085 105.395 58.350 105.855 ;
        RECT 56.690 104.875 57.220 105.240 ;
        RECT 57.665 105.130 57.970 105.260 ;
        RECT 56.010 104.705 56.520 104.795 ;
        RECT 56.010 104.535 56.880 104.705 ;
        RECT 56.010 104.465 56.180 104.535 ;
        RECT 56.300 104.285 56.500 104.315 ;
        RECT 54.820 103.925 55.285 104.255 ;
        RECT 55.670 103.985 56.500 104.285 ;
        RECT 55.670 103.755 55.840 103.985 ;
        RECT 54.480 103.585 55.265 103.755 ;
        RECT 55.435 103.585 55.840 103.755 ;
        RECT 56.020 103.305 56.390 103.805 ;
        RECT 56.710 103.755 56.880 104.535 ;
        RECT 57.050 104.175 57.220 104.875 ;
        RECT 57.390 104.345 57.630 104.940 ;
        RECT 57.050 103.955 57.575 104.175 ;
        RECT 57.800 104.025 57.970 105.130 ;
        RECT 57.745 103.895 57.970 104.025 ;
        RECT 58.140 103.935 58.420 104.885 ;
        RECT 57.745 103.755 57.915 103.895 ;
        RECT 56.710 103.585 57.385 103.755 ;
        RECT 57.580 103.585 57.915 103.755 ;
        RECT 58.085 103.305 58.335 103.765 ;
        RECT 58.590 103.565 58.775 105.685 ;
        RECT 58.945 105.355 59.275 105.855 ;
        RECT 59.445 105.185 59.615 105.685 ;
        RECT 58.950 105.015 59.615 105.185 ;
        RECT 60.425 105.185 60.595 105.685 ;
        RECT 60.765 105.355 61.095 105.855 ;
        RECT 60.425 105.015 61.090 105.185 ;
        RECT 58.950 104.025 59.180 105.015 ;
        RECT 59.350 104.195 59.700 104.845 ;
        RECT 60.340 104.195 60.690 104.845 ;
        RECT 60.860 104.025 61.090 105.015 ;
        RECT 58.950 103.855 59.615 104.025 ;
        RECT 58.945 103.305 59.275 103.685 ;
        RECT 59.445 103.565 59.615 103.855 ;
        RECT 60.425 103.855 61.090 104.025 ;
        RECT 60.425 103.565 60.595 103.855 ;
        RECT 60.765 103.305 61.095 103.685 ;
        RECT 61.265 103.565 61.450 105.685 ;
        RECT 61.690 105.395 61.955 105.855 ;
        RECT 62.125 105.260 62.375 105.685 ;
        RECT 62.585 105.410 63.690 105.580 ;
        RECT 62.070 105.130 62.375 105.260 ;
        RECT 61.620 103.935 61.900 104.885 ;
        RECT 62.070 104.025 62.240 105.130 ;
        RECT 62.410 104.345 62.650 104.940 ;
        RECT 62.820 104.875 63.350 105.240 ;
        RECT 62.820 104.175 62.990 104.875 ;
        RECT 63.520 104.795 63.690 105.410 ;
        RECT 63.860 105.055 64.030 105.855 ;
        RECT 64.200 105.355 64.450 105.685 ;
        RECT 64.675 105.385 65.560 105.555 ;
        RECT 63.520 104.705 64.030 104.795 ;
        RECT 62.070 103.895 62.295 104.025 ;
        RECT 62.465 103.955 62.990 104.175 ;
        RECT 63.160 104.535 64.030 104.705 ;
        RECT 61.705 103.305 61.955 103.765 ;
        RECT 62.125 103.755 62.295 103.895 ;
        RECT 63.160 103.755 63.330 104.535 ;
        RECT 63.860 104.465 64.030 104.535 ;
        RECT 63.540 104.285 63.740 104.315 ;
        RECT 64.200 104.285 64.370 105.355 ;
        RECT 64.540 104.465 64.730 105.185 ;
        RECT 63.540 103.985 64.370 104.285 ;
        RECT 64.900 104.255 65.220 105.215 ;
        RECT 62.125 103.585 62.460 103.755 ;
        RECT 62.655 103.585 63.330 103.755 ;
        RECT 63.650 103.305 64.020 103.805 ;
        RECT 64.200 103.755 64.370 103.985 ;
        RECT 64.755 103.925 65.220 104.255 ;
        RECT 65.390 104.545 65.560 105.385 ;
        RECT 65.740 105.355 66.055 105.855 ;
        RECT 66.285 105.125 66.625 105.685 ;
        RECT 65.730 104.750 66.625 105.125 ;
        RECT 66.795 104.845 66.965 105.855 ;
        RECT 66.435 104.545 66.625 104.750 ;
        RECT 67.135 104.795 67.465 105.640 ;
        RECT 67.695 105.420 73.040 105.855 ;
        RECT 67.135 104.715 67.525 104.795 ;
        RECT 67.310 104.665 67.525 104.715 ;
        RECT 65.390 104.215 66.265 104.545 ;
        RECT 66.435 104.215 67.185 104.545 ;
        RECT 65.390 103.755 65.560 104.215 ;
        RECT 66.435 104.045 66.635 104.215 ;
        RECT 67.355 104.085 67.525 104.665 ;
        RECT 67.300 104.045 67.525 104.085 ;
        RECT 64.200 103.585 64.605 103.755 ;
        RECT 64.775 103.585 65.560 103.755 ;
        RECT 65.835 103.305 66.045 103.835 ;
        RECT 66.305 103.520 66.635 104.045 ;
        RECT 67.145 103.960 67.525 104.045 ;
        RECT 66.805 103.305 66.975 103.915 ;
        RECT 67.145 103.525 67.475 103.960 ;
        RECT 69.280 103.850 69.620 104.680 ;
        RECT 71.100 104.170 71.450 105.420 ;
        RECT 73.215 104.765 74.885 105.855 ;
        RECT 73.215 104.075 73.965 104.595 ;
        RECT 74.135 104.245 74.885 104.765 ;
        RECT 75.550 105.065 76.085 105.685 ;
        RECT 67.695 103.305 73.040 103.850 ;
        RECT 73.215 103.305 74.885 104.075 ;
        RECT 75.550 104.045 75.865 105.065 ;
        RECT 76.255 105.055 76.585 105.855 ;
        RECT 77.070 104.885 77.460 105.060 ;
        RECT 76.035 104.715 77.460 104.885 ;
        RECT 76.035 104.215 76.205 104.715 ;
        RECT 75.550 103.475 76.165 104.045 ;
        RECT 76.455 103.985 76.720 104.545 ;
        RECT 76.890 103.815 77.060 104.715 ;
        RECT 77.815 104.690 78.105 105.855 ;
        RECT 78.275 104.715 78.615 105.685 ;
        RECT 78.785 104.715 78.955 105.855 ;
        RECT 79.225 105.055 79.475 105.855 ;
        RECT 80.120 104.885 80.450 105.685 ;
        RECT 80.750 105.055 81.080 105.855 ;
        RECT 81.250 104.885 81.580 105.685 ;
        RECT 79.145 104.715 81.580 104.885 ;
        RECT 82.420 104.905 82.685 105.675 ;
        RECT 82.855 105.135 83.185 105.855 ;
        RECT 83.375 105.315 83.635 105.675 ;
        RECT 83.805 105.485 84.135 105.855 ;
        RECT 84.305 105.315 84.565 105.675 ;
        RECT 83.375 105.085 84.565 105.315 ;
        RECT 85.135 104.905 85.425 105.675 ;
        RECT 85.725 105.185 85.895 105.685 ;
        RECT 86.065 105.355 86.395 105.855 ;
        RECT 85.725 105.015 86.390 105.185 ;
        RECT 77.230 103.985 77.585 104.545 ;
        RECT 78.275 104.105 78.450 104.715 ;
        RECT 79.145 104.465 79.315 104.715 ;
        RECT 78.620 104.295 79.315 104.465 ;
        RECT 79.490 104.295 79.910 104.495 ;
        RECT 80.080 104.295 80.410 104.495 ;
        RECT 80.580 104.295 80.910 104.495 ;
        RECT 76.335 103.305 76.550 103.815 ;
        RECT 76.780 103.485 77.060 103.815 ;
        RECT 77.240 103.305 77.480 103.815 ;
        RECT 77.815 103.305 78.105 104.030 ;
        RECT 78.275 103.475 78.615 104.105 ;
        RECT 78.785 103.305 79.035 104.105 ;
        RECT 79.225 103.955 80.450 104.125 ;
        RECT 79.225 103.475 79.555 103.955 ;
        RECT 79.725 103.305 79.950 103.765 ;
        RECT 80.120 103.475 80.450 103.955 ;
        RECT 81.080 104.085 81.250 104.715 ;
        RECT 81.435 104.295 81.785 104.545 ;
        RECT 81.080 103.475 81.580 104.085 ;
        RECT 82.420 103.485 82.755 104.905 ;
        RECT 82.930 104.725 85.425 104.905 ;
        RECT 82.930 104.035 83.155 104.725 ;
        RECT 83.355 104.215 83.635 104.545 ;
        RECT 83.815 104.215 84.390 104.545 ;
        RECT 84.570 104.215 85.005 104.545 ;
        RECT 85.185 104.215 85.455 104.545 ;
        RECT 85.640 104.195 85.990 104.845 ;
        RECT 82.930 103.845 85.415 104.035 ;
        RECT 86.160 104.025 86.390 105.015 ;
        RECT 82.935 103.305 83.680 103.675 ;
        RECT 84.245 103.485 84.500 103.845 ;
        RECT 84.680 103.305 85.010 103.675 ;
        RECT 85.190 103.485 85.415 103.845 ;
        RECT 85.725 103.855 86.390 104.025 ;
        RECT 85.725 103.565 85.895 103.855 ;
        RECT 86.065 103.305 86.395 103.685 ;
        RECT 86.565 103.565 86.750 105.685 ;
        RECT 86.990 105.395 87.255 105.855 ;
        RECT 87.425 105.260 87.675 105.685 ;
        RECT 87.885 105.410 88.990 105.580 ;
        RECT 87.370 105.130 87.675 105.260 ;
        RECT 86.920 103.935 87.200 104.885 ;
        RECT 87.370 104.025 87.540 105.130 ;
        RECT 87.710 104.345 87.950 104.940 ;
        RECT 88.120 104.875 88.650 105.240 ;
        RECT 88.120 104.175 88.290 104.875 ;
        RECT 88.820 104.795 88.990 105.410 ;
        RECT 89.160 105.055 89.330 105.855 ;
        RECT 89.500 105.355 89.750 105.685 ;
        RECT 89.975 105.385 90.860 105.555 ;
        RECT 88.820 104.705 89.330 104.795 ;
        RECT 87.370 103.895 87.595 104.025 ;
        RECT 87.765 103.955 88.290 104.175 ;
        RECT 88.460 104.535 89.330 104.705 ;
        RECT 87.005 103.305 87.255 103.765 ;
        RECT 87.425 103.755 87.595 103.895 ;
        RECT 88.460 103.755 88.630 104.535 ;
        RECT 89.160 104.465 89.330 104.535 ;
        RECT 88.840 104.285 89.040 104.315 ;
        RECT 89.500 104.285 89.670 105.355 ;
        RECT 89.840 104.465 90.030 105.185 ;
        RECT 88.840 103.985 89.670 104.285 ;
        RECT 90.200 104.255 90.520 105.215 ;
        RECT 87.425 103.585 87.760 103.755 ;
        RECT 87.955 103.585 88.630 103.755 ;
        RECT 88.950 103.305 89.320 103.805 ;
        RECT 89.500 103.755 89.670 103.985 ;
        RECT 90.055 103.925 90.520 104.255 ;
        RECT 90.690 104.545 90.860 105.385 ;
        RECT 91.040 105.355 91.355 105.855 ;
        RECT 91.585 105.125 91.925 105.685 ;
        RECT 91.030 104.750 91.925 105.125 ;
        RECT 92.095 104.845 92.265 105.855 ;
        RECT 91.735 104.545 91.925 104.750 ;
        RECT 92.435 104.795 92.765 105.640 ;
        RECT 93.030 105.065 93.565 105.685 ;
        RECT 92.435 104.715 92.825 104.795 ;
        RECT 92.610 104.665 92.825 104.715 ;
        RECT 90.690 104.215 91.565 104.545 ;
        RECT 91.735 104.215 92.485 104.545 ;
        RECT 90.690 103.755 90.860 104.215 ;
        RECT 91.735 104.045 91.935 104.215 ;
        RECT 92.655 104.085 92.825 104.665 ;
        RECT 92.600 104.045 92.825 104.085 ;
        RECT 89.500 103.585 89.905 103.755 ;
        RECT 90.075 103.585 90.860 103.755 ;
        RECT 91.135 103.305 91.345 103.835 ;
        RECT 91.605 103.520 91.935 104.045 ;
        RECT 92.445 103.960 92.825 104.045 ;
        RECT 93.030 104.045 93.345 105.065 ;
        RECT 93.735 105.055 94.065 105.855 ;
        RECT 94.550 104.885 94.940 105.060 ;
        RECT 93.515 104.715 94.940 104.885 ;
        RECT 95.755 104.715 96.015 105.855 ;
        RECT 96.185 104.885 96.515 105.685 ;
        RECT 96.685 105.055 96.855 105.855 ;
        RECT 97.025 104.885 97.355 105.685 ;
        RECT 97.525 105.055 97.780 105.855 ;
        RECT 98.055 105.135 98.515 105.685 ;
        RECT 98.705 105.135 99.035 105.855 ;
        RECT 96.185 104.715 97.885 104.885 ;
        RECT 93.515 104.215 93.685 104.715 ;
        RECT 92.105 103.305 92.275 103.915 ;
        RECT 92.445 103.525 92.775 103.960 ;
        RECT 93.030 103.475 93.645 104.045 ;
        RECT 93.935 103.985 94.200 104.545 ;
        RECT 94.370 103.815 94.540 104.715 ;
        RECT 94.710 103.985 95.065 104.545 ;
        RECT 95.755 104.295 96.515 104.545 ;
        RECT 96.685 104.295 97.435 104.545 ;
        RECT 97.605 104.125 97.885 104.715 ;
        RECT 95.755 103.935 96.855 104.105 ;
        RECT 93.815 103.305 94.030 103.815 ;
        RECT 94.260 103.485 94.540 103.815 ;
        RECT 94.720 103.305 94.960 103.815 ;
        RECT 95.755 103.475 96.095 103.935 ;
        RECT 96.265 103.305 96.435 103.765 ;
        RECT 96.605 103.685 96.855 103.935 ;
        RECT 97.025 103.875 97.885 104.125 ;
        RECT 98.055 103.765 98.305 105.135 ;
        RECT 99.235 104.965 99.535 105.515 ;
        RECT 99.705 105.185 99.985 105.855 ;
        RECT 98.595 104.795 99.535 104.965 ;
        RECT 98.595 104.545 98.765 104.795 ;
        RECT 99.905 104.545 100.170 104.905 ;
        RECT 100.355 104.765 102.945 105.855 ;
        RECT 98.475 104.215 98.765 104.545 ;
        RECT 98.935 104.295 99.275 104.545 ;
        RECT 99.495 104.295 100.170 104.545 ;
        RECT 98.595 104.125 98.765 104.215 ;
        RECT 98.595 103.935 99.985 104.125 ;
        RECT 97.445 103.685 97.775 103.705 ;
        RECT 96.605 103.475 97.775 103.685 ;
        RECT 98.055 103.475 98.615 103.765 ;
        RECT 98.785 103.305 99.035 103.765 ;
        RECT 99.655 103.575 99.985 103.935 ;
        RECT 100.355 104.075 101.565 104.595 ;
        RECT 101.735 104.245 102.945 104.765 ;
        RECT 103.575 104.690 103.865 105.855 ;
        RECT 104.035 104.765 107.545 105.855 ;
        RECT 107.715 104.765 108.925 105.855 ;
        RECT 104.035 104.075 105.685 104.595 ;
        RECT 105.855 104.245 107.545 104.765 ;
        RECT 100.355 103.305 102.945 104.075 ;
        RECT 103.575 103.305 103.865 104.030 ;
        RECT 104.035 103.305 107.545 104.075 ;
        RECT 107.715 104.055 108.235 104.595 ;
        RECT 108.405 104.225 108.925 104.765 ;
        RECT 109.095 104.715 109.355 105.855 ;
        RECT 109.525 104.885 109.855 105.685 ;
        RECT 110.025 105.055 110.195 105.855 ;
        RECT 110.365 104.885 110.695 105.685 ;
        RECT 110.865 105.055 111.120 105.855 ;
        RECT 111.485 105.185 111.655 105.685 ;
        RECT 111.825 105.355 112.155 105.855 ;
        RECT 111.485 105.015 112.150 105.185 ;
        RECT 109.525 104.715 111.225 104.885 ;
        RECT 109.095 104.295 109.855 104.545 ;
        RECT 110.025 104.295 110.775 104.545 ;
        RECT 110.945 104.125 111.225 104.715 ;
        RECT 111.400 104.195 111.750 104.845 ;
        RECT 107.715 103.305 108.925 104.055 ;
        RECT 109.095 103.935 110.195 104.105 ;
        RECT 109.095 103.475 109.435 103.935 ;
        RECT 109.605 103.305 109.775 103.765 ;
        RECT 109.945 103.685 110.195 103.935 ;
        RECT 110.365 103.875 111.225 104.125 ;
        RECT 111.920 104.025 112.150 105.015 ;
        RECT 111.485 103.855 112.150 104.025 ;
        RECT 110.785 103.685 111.115 103.705 ;
        RECT 109.945 103.475 111.115 103.685 ;
        RECT 111.485 103.565 111.655 103.855 ;
        RECT 111.825 103.305 112.155 103.685 ;
        RECT 112.325 103.565 112.510 105.685 ;
        RECT 112.750 105.395 113.015 105.855 ;
        RECT 113.185 105.260 113.435 105.685 ;
        RECT 113.645 105.410 114.750 105.580 ;
        RECT 113.130 105.130 113.435 105.260 ;
        RECT 112.680 103.935 112.960 104.885 ;
        RECT 113.130 104.025 113.300 105.130 ;
        RECT 113.470 104.345 113.710 104.940 ;
        RECT 113.880 104.875 114.410 105.240 ;
        RECT 113.880 104.175 114.050 104.875 ;
        RECT 114.580 104.795 114.750 105.410 ;
        RECT 114.920 105.055 115.090 105.855 ;
        RECT 115.260 105.355 115.510 105.685 ;
        RECT 115.735 105.385 116.620 105.555 ;
        RECT 114.580 104.705 115.090 104.795 ;
        RECT 113.130 103.895 113.355 104.025 ;
        RECT 113.525 103.955 114.050 104.175 ;
        RECT 114.220 104.535 115.090 104.705 ;
        RECT 112.765 103.305 113.015 103.765 ;
        RECT 113.185 103.755 113.355 103.895 ;
        RECT 114.220 103.755 114.390 104.535 ;
        RECT 114.920 104.465 115.090 104.535 ;
        RECT 114.600 104.285 114.800 104.315 ;
        RECT 115.260 104.285 115.430 105.355 ;
        RECT 115.600 104.465 115.790 105.185 ;
        RECT 114.600 103.985 115.430 104.285 ;
        RECT 115.960 104.255 116.280 105.215 ;
        RECT 113.185 103.585 113.520 103.755 ;
        RECT 113.715 103.585 114.390 103.755 ;
        RECT 114.710 103.305 115.080 103.805 ;
        RECT 115.260 103.755 115.430 103.985 ;
        RECT 115.815 103.925 116.280 104.255 ;
        RECT 116.450 104.545 116.620 105.385 ;
        RECT 116.800 105.355 117.115 105.855 ;
        RECT 117.345 105.125 117.685 105.685 ;
        RECT 116.790 104.750 117.685 105.125 ;
        RECT 117.855 104.845 118.025 105.855 ;
        RECT 117.495 104.545 117.685 104.750 ;
        RECT 118.195 104.795 118.525 105.640 ;
        RECT 118.755 105.420 124.100 105.855 ;
        RECT 118.195 104.715 118.585 104.795 ;
        RECT 118.370 104.665 118.585 104.715 ;
        RECT 116.450 104.215 117.325 104.545 ;
        RECT 117.495 104.215 118.245 104.545 ;
        RECT 116.450 103.755 116.620 104.215 ;
        RECT 117.495 104.045 117.695 104.215 ;
        RECT 118.415 104.085 118.585 104.665 ;
        RECT 118.360 104.045 118.585 104.085 ;
        RECT 115.260 103.585 115.665 103.755 ;
        RECT 115.835 103.585 116.620 103.755 ;
        RECT 116.895 103.305 117.105 103.835 ;
        RECT 117.365 103.520 117.695 104.045 ;
        RECT 118.205 103.960 118.585 104.045 ;
        RECT 117.865 103.305 118.035 103.915 ;
        RECT 118.205 103.525 118.535 103.960 ;
        RECT 120.340 103.850 120.680 104.680 ;
        RECT 122.160 104.170 122.510 105.420 ;
        RECT 124.770 105.065 125.305 105.685 ;
        RECT 124.770 104.045 125.085 105.065 ;
        RECT 125.475 105.055 125.805 105.855 ;
        RECT 127.070 105.065 127.605 105.685 ;
        RECT 126.290 104.885 126.680 105.060 ;
        RECT 125.255 104.715 126.680 104.885 ;
        RECT 125.255 104.215 125.425 104.715 ;
        RECT 118.755 103.305 124.100 103.850 ;
        RECT 124.770 103.475 125.385 104.045 ;
        RECT 125.675 103.985 125.940 104.545 ;
        RECT 126.110 103.815 126.280 104.715 ;
        RECT 126.450 103.985 126.805 104.545 ;
        RECT 127.070 104.045 127.385 105.065 ;
        RECT 127.775 105.055 128.105 105.855 ;
        RECT 128.590 104.885 128.980 105.060 ;
        RECT 127.555 104.715 128.980 104.885 ;
        RECT 127.555 104.215 127.725 104.715 ;
        RECT 125.555 103.305 125.770 103.815 ;
        RECT 126.000 103.485 126.280 103.815 ;
        RECT 126.460 103.305 126.700 103.815 ;
        RECT 127.070 103.475 127.685 104.045 ;
        RECT 127.975 103.985 128.240 104.545 ;
        RECT 128.410 103.815 128.580 104.715 ;
        RECT 129.335 104.690 129.625 105.855 ;
        RECT 129.795 105.005 130.055 105.685 ;
        RECT 130.225 105.075 130.475 105.855 ;
        RECT 130.725 105.305 130.975 105.685 ;
        RECT 131.145 105.475 131.500 105.855 ;
        RECT 132.505 105.465 132.840 105.685 ;
        RECT 132.105 105.305 132.335 105.345 ;
        RECT 130.725 105.105 132.335 105.305 ;
        RECT 130.725 105.095 131.560 105.105 ;
        RECT 132.150 105.015 132.335 105.105 ;
        RECT 128.750 103.985 129.105 104.545 ;
        RECT 127.855 103.305 128.070 103.815 ;
        RECT 128.300 103.485 128.580 103.815 ;
        RECT 128.760 103.305 129.000 103.815 ;
        RECT 129.335 103.305 129.625 104.030 ;
        RECT 129.795 103.815 129.965 105.005 ;
        RECT 131.665 104.905 131.995 104.935 ;
        RECT 130.195 104.845 131.995 104.905 ;
        RECT 132.585 104.845 132.840 105.465 ;
        RECT 130.135 104.735 132.840 104.845 ;
        RECT 130.135 104.700 130.335 104.735 ;
        RECT 130.135 104.125 130.305 104.700 ;
        RECT 131.665 104.675 132.840 104.735 ;
        RECT 133.200 104.885 133.590 105.060 ;
        RECT 134.075 105.055 134.405 105.855 ;
        RECT 134.575 105.065 135.110 105.685 ;
        RECT 133.200 104.715 134.625 104.885 ;
        RECT 130.535 104.260 130.945 104.565 ;
        RECT 131.115 104.295 131.445 104.505 ;
        RECT 130.135 104.005 130.405 104.125 ;
        RECT 130.135 103.960 130.980 104.005 ;
        RECT 130.225 103.835 130.980 103.960 ;
        RECT 131.235 103.895 131.445 104.295 ;
        RECT 131.690 104.295 132.165 104.505 ;
        RECT 132.355 104.295 132.845 104.495 ;
        RECT 131.690 103.895 131.910 104.295 ;
        RECT 129.795 103.805 130.025 103.815 ;
        RECT 129.795 103.475 130.055 103.805 ;
        RECT 130.810 103.685 130.980 103.835 ;
        RECT 130.225 103.305 130.555 103.665 ;
        RECT 130.810 103.475 132.110 103.685 ;
        RECT 132.385 103.305 132.840 104.070 ;
        RECT 133.075 103.985 133.430 104.545 ;
        RECT 133.600 103.815 133.770 104.715 ;
        RECT 133.940 103.985 134.205 104.545 ;
        RECT 134.455 104.215 134.625 104.715 ;
        RECT 134.795 104.045 135.110 105.065 ;
        RECT 135.865 104.925 136.035 105.685 ;
        RECT 136.250 105.095 136.580 105.855 ;
        RECT 135.865 104.755 136.580 104.925 ;
        RECT 136.750 104.780 137.005 105.685 ;
        RECT 135.775 104.205 136.130 104.575 ;
        RECT 136.410 104.545 136.580 104.755 ;
        RECT 136.410 104.215 136.665 104.545 ;
        RECT 133.180 103.305 133.420 103.815 ;
        RECT 133.600 103.485 133.880 103.815 ;
        RECT 134.110 103.305 134.325 103.815 ;
        RECT 134.495 103.475 135.110 104.045 ;
        RECT 136.410 104.025 136.580 104.215 ;
        RECT 136.835 104.050 137.005 104.780 ;
        RECT 137.180 104.705 137.440 105.855 ;
        RECT 137.615 104.765 138.825 105.855 ;
        RECT 137.615 104.225 138.135 104.765 ;
        RECT 135.865 103.855 136.580 104.025 ;
        RECT 135.865 103.475 136.035 103.855 ;
        RECT 136.250 103.305 136.580 103.685 ;
        RECT 136.750 103.475 137.005 104.050 ;
        RECT 137.180 103.305 137.440 104.145 ;
        RECT 138.305 104.055 138.825 104.595 ;
        RECT 137.615 103.305 138.825 104.055 ;
        RECT 13.330 103.135 138.910 103.305 ;
        RECT 13.415 102.385 14.625 103.135 ;
        RECT 13.415 101.845 13.935 102.385 ;
        RECT 14.795 102.365 17.385 103.135 ;
        RECT 14.105 101.675 14.625 102.215 ;
        RECT 14.795 101.845 16.005 102.365 ;
        RECT 17.555 102.335 17.865 103.135 ;
        RECT 18.070 102.335 18.765 102.965 ;
        RECT 18.955 102.445 19.195 102.965 ;
        RECT 19.365 102.640 19.760 103.135 ;
        RECT 20.325 102.805 20.495 102.950 ;
        RECT 20.120 102.610 20.495 102.805 ;
        RECT 16.175 101.675 17.385 102.195 ;
        RECT 17.565 101.895 17.900 102.165 ;
        RECT 18.070 101.735 18.240 102.335 ;
        RECT 18.410 101.895 18.745 102.145 ;
        RECT 13.415 100.585 14.625 101.675 ;
        RECT 14.795 100.585 17.385 101.675 ;
        RECT 17.555 100.585 17.835 101.725 ;
        RECT 18.005 100.755 18.335 101.735 ;
        RECT 18.505 100.585 18.765 101.725 ;
        RECT 18.955 101.640 19.130 102.445 ;
        RECT 20.120 102.275 20.290 102.610 ;
        RECT 20.775 102.565 21.015 102.940 ;
        RECT 21.185 102.630 21.520 103.135 ;
        RECT 20.775 102.415 20.995 102.565 ;
        RECT 21.745 102.480 22.075 102.915 ;
        RECT 22.245 102.525 22.415 103.135 ;
        RECT 19.305 101.915 20.290 102.275 ;
        RECT 20.460 102.085 20.995 102.415 ;
        RECT 19.305 101.895 20.590 101.915 ;
        RECT 19.730 101.745 20.590 101.895 ;
        RECT 18.955 100.855 19.260 101.640 ;
        RECT 19.435 101.265 20.130 101.575 ;
        RECT 19.440 100.585 20.125 101.055 ;
        RECT 20.305 100.800 20.590 101.745 ;
        RECT 20.760 101.435 20.995 102.085 ;
        RECT 21.165 101.605 21.465 102.455 ;
        RECT 21.695 102.395 22.075 102.480 ;
        RECT 22.585 102.395 22.915 102.920 ;
        RECT 23.175 102.605 23.385 103.135 ;
        RECT 23.660 102.685 24.445 102.855 ;
        RECT 24.615 102.685 25.020 102.855 ;
        RECT 21.695 102.355 21.920 102.395 ;
        RECT 21.695 101.775 21.865 102.355 ;
        RECT 22.585 102.225 22.785 102.395 ;
        RECT 23.660 102.225 23.830 102.685 ;
        RECT 22.035 101.895 22.785 102.225 ;
        RECT 22.955 101.895 23.830 102.225 ;
        RECT 21.695 101.725 21.910 101.775 ;
        RECT 21.695 101.645 22.085 101.725 ;
        RECT 20.760 101.205 21.435 101.435 ;
        RECT 20.765 100.585 21.095 101.035 ;
        RECT 21.265 100.775 21.435 101.205 ;
        RECT 21.755 100.800 22.085 101.645 ;
        RECT 22.595 101.690 22.785 101.895 ;
        RECT 22.255 100.585 22.425 101.595 ;
        RECT 22.595 101.315 23.490 101.690 ;
        RECT 22.595 100.755 22.935 101.315 ;
        RECT 23.165 100.585 23.480 101.085 ;
        RECT 23.660 101.055 23.830 101.895 ;
        RECT 24.000 102.185 24.465 102.515 ;
        RECT 24.850 102.455 25.020 102.685 ;
        RECT 25.200 102.635 25.570 103.135 ;
        RECT 25.890 102.685 26.565 102.855 ;
        RECT 26.760 102.685 27.095 102.855 ;
        RECT 24.000 101.225 24.320 102.185 ;
        RECT 24.850 102.155 25.680 102.455 ;
        RECT 24.490 101.255 24.680 101.975 ;
        RECT 24.850 101.085 25.020 102.155 ;
        RECT 25.480 102.125 25.680 102.155 ;
        RECT 25.190 101.905 25.360 101.975 ;
        RECT 25.890 101.905 26.060 102.685 ;
        RECT 26.925 102.545 27.095 102.685 ;
        RECT 27.265 102.675 27.515 103.135 ;
        RECT 25.190 101.735 26.060 101.905 ;
        RECT 26.230 102.265 26.755 102.485 ;
        RECT 26.925 102.415 27.150 102.545 ;
        RECT 25.190 101.645 25.700 101.735 ;
        RECT 23.660 100.885 24.545 101.055 ;
        RECT 24.770 100.755 25.020 101.085 ;
        RECT 25.190 100.585 25.360 101.385 ;
        RECT 25.530 101.030 25.700 101.645 ;
        RECT 26.230 101.565 26.400 102.265 ;
        RECT 25.870 101.200 26.400 101.565 ;
        RECT 26.570 101.500 26.810 102.095 ;
        RECT 26.980 101.310 27.150 102.415 ;
        RECT 27.320 101.555 27.600 102.505 ;
        RECT 26.845 101.180 27.150 101.310 ;
        RECT 25.530 100.860 26.635 101.030 ;
        RECT 26.845 100.755 27.095 101.180 ;
        RECT 27.265 100.585 27.530 101.045 ;
        RECT 27.770 100.755 27.955 102.875 ;
        RECT 28.125 102.755 28.455 103.135 ;
        RECT 28.625 102.585 28.795 102.875 ;
        RECT 28.130 102.415 28.795 102.585 ;
        RECT 29.055 102.485 29.315 102.965 ;
        RECT 29.485 102.595 29.735 103.135 ;
        RECT 28.130 101.425 28.360 102.415 ;
        RECT 28.530 101.595 28.880 102.245 ;
        RECT 29.055 101.455 29.225 102.485 ;
        RECT 29.905 102.430 30.125 102.915 ;
        RECT 29.395 101.835 29.625 102.230 ;
        RECT 29.795 102.005 30.125 102.430 ;
        RECT 30.295 102.755 31.185 102.925 ;
        RECT 30.295 102.030 30.465 102.755 ;
        RECT 30.635 102.200 31.185 102.585 ;
        RECT 31.355 102.365 34.865 103.135 ;
        RECT 35.495 102.485 35.755 102.965 ;
        RECT 35.925 102.675 36.255 103.135 ;
        RECT 36.445 102.495 36.645 102.915 ;
        RECT 30.295 101.960 31.185 102.030 ;
        RECT 30.290 101.935 31.185 101.960 ;
        RECT 30.280 101.920 31.185 101.935 ;
        RECT 30.275 101.905 31.185 101.920 ;
        RECT 30.265 101.900 31.185 101.905 ;
        RECT 30.260 101.890 31.185 101.900 ;
        RECT 30.255 101.880 31.185 101.890 ;
        RECT 30.245 101.875 31.185 101.880 ;
        RECT 30.235 101.865 31.185 101.875 ;
        RECT 30.225 101.860 31.185 101.865 ;
        RECT 30.225 101.855 30.560 101.860 ;
        RECT 30.210 101.850 30.560 101.855 ;
        RECT 30.195 101.840 30.560 101.850 ;
        RECT 30.170 101.835 30.560 101.840 ;
        RECT 29.395 101.830 30.560 101.835 ;
        RECT 29.395 101.795 30.530 101.830 ;
        RECT 29.395 101.770 30.495 101.795 ;
        RECT 29.395 101.740 30.465 101.770 ;
        RECT 29.395 101.710 30.445 101.740 ;
        RECT 29.395 101.680 30.425 101.710 ;
        RECT 29.395 101.670 30.355 101.680 ;
        RECT 29.395 101.660 30.330 101.670 ;
        RECT 29.395 101.645 30.310 101.660 ;
        RECT 29.395 101.630 30.290 101.645 ;
        RECT 29.500 101.620 30.285 101.630 ;
        RECT 29.500 101.585 30.270 101.620 ;
        RECT 28.130 101.255 28.795 101.425 ;
        RECT 28.125 100.585 28.455 101.085 ;
        RECT 28.625 100.755 28.795 101.255 ;
        RECT 29.055 100.755 29.330 101.455 ;
        RECT 29.500 101.335 30.255 101.585 ;
        RECT 30.425 101.265 30.755 101.510 ;
        RECT 30.925 101.410 31.185 101.860 ;
        RECT 31.355 101.845 33.005 102.365 ;
        RECT 33.175 101.675 34.865 102.195 ;
        RECT 30.570 101.240 30.755 101.265 ;
        RECT 30.570 101.140 31.185 101.240 ;
        RECT 29.500 100.585 29.755 101.130 ;
        RECT 29.925 100.755 30.405 101.095 ;
        RECT 30.580 100.585 31.185 101.140 ;
        RECT 31.355 100.585 34.865 101.675 ;
        RECT 35.495 101.455 35.665 102.485 ;
        RECT 35.835 101.795 36.065 102.225 ;
        RECT 36.235 101.975 36.645 102.495 ;
        RECT 36.815 102.650 37.605 102.915 ;
        RECT 36.815 101.795 37.070 102.650 ;
        RECT 37.785 102.315 38.115 102.735 ;
        RECT 38.285 102.315 38.545 103.135 ;
        RECT 39.175 102.410 39.465 103.135 ;
        RECT 39.635 102.755 40.525 102.925 ;
        RECT 37.785 102.225 38.035 102.315 ;
        RECT 37.240 101.975 38.035 102.225 ;
        RECT 39.635 102.200 40.185 102.585 ;
        RECT 35.835 101.625 37.625 101.795 ;
        RECT 35.495 100.755 35.770 101.455 ;
        RECT 35.940 101.330 36.655 101.625 ;
        RECT 36.875 101.265 37.205 101.455 ;
        RECT 35.980 100.585 36.195 101.130 ;
        RECT 36.365 100.755 36.840 101.095 ;
        RECT 37.010 101.090 37.205 101.265 ;
        RECT 37.375 101.260 37.625 101.625 ;
        RECT 37.010 100.585 37.625 101.090 ;
        RECT 37.865 100.755 38.035 101.975 ;
        RECT 38.205 101.265 38.545 102.145 ;
        RECT 40.355 102.030 40.525 102.755 ;
        RECT 39.635 101.960 40.525 102.030 ;
        RECT 40.695 102.430 40.915 102.915 ;
        RECT 41.085 102.595 41.335 103.135 ;
        RECT 41.505 102.485 41.765 102.965 ;
        RECT 40.695 102.005 41.025 102.430 ;
        RECT 39.635 101.935 40.530 101.960 ;
        RECT 39.635 101.920 40.540 101.935 ;
        RECT 39.635 101.905 40.545 101.920 ;
        RECT 39.635 101.900 40.555 101.905 ;
        RECT 39.635 101.890 40.560 101.900 ;
        RECT 39.635 101.880 40.565 101.890 ;
        RECT 39.635 101.875 40.575 101.880 ;
        RECT 39.635 101.865 40.585 101.875 ;
        RECT 39.635 101.860 40.595 101.865 ;
        RECT 38.285 100.585 38.545 101.095 ;
        RECT 39.175 100.585 39.465 101.750 ;
        RECT 39.635 101.410 39.895 101.860 ;
        RECT 40.260 101.855 40.595 101.860 ;
        RECT 40.260 101.850 40.610 101.855 ;
        RECT 40.260 101.840 40.625 101.850 ;
        RECT 40.260 101.835 40.650 101.840 ;
        RECT 41.195 101.835 41.425 102.230 ;
        RECT 40.260 101.830 41.425 101.835 ;
        RECT 40.290 101.795 41.425 101.830 ;
        RECT 40.325 101.770 41.425 101.795 ;
        RECT 40.355 101.740 41.425 101.770 ;
        RECT 40.375 101.710 41.425 101.740 ;
        RECT 40.395 101.680 41.425 101.710 ;
        RECT 40.465 101.670 41.425 101.680 ;
        RECT 40.490 101.660 41.425 101.670 ;
        RECT 40.510 101.645 41.425 101.660 ;
        RECT 40.530 101.630 41.425 101.645 ;
        RECT 40.535 101.620 41.320 101.630 ;
        RECT 40.550 101.585 41.320 101.620 ;
        RECT 40.065 101.265 40.395 101.510 ;
        RECT 40.565 101.335 41.320 101.585 ;
        RECT 41.595 101.455 41.765 102.485 ;
        RECT 41.935 102.365 44.525 103.135 ;
        RECT 45.320 102.625 45.560 103.135 ;
        RECT 45.740 102.625 46.020 102.955 ;
        RECT 46.250 102.625 46.465 103.135 ;
        RECT 41.935 101.845 43.145 102.365 ;
        RECT 43.315 101.675 44.525 102.195 ;
        RECT 45.215 101.895 45.570 102.455 ;
        RECT 45.740 101.725 45.910 102.625 ;
        RECT 46.080 101.895 46.345 102.455 ;
        RECT 46.635 102.395 47.250 102.965 ;
        RECT 47.505 102.480 47.835 102.915 ;
        RECT 48.005 102.525 48.175 103.135 ;
        RECT 46.595 101.725 46.765 102.225 ;
        RECT 40.065 101.240 40.250 101.265 ;
        RECT 39.635 101.140 40.250 101.240 ;
        RECT 39.635 100.585 40.240 101.140 ;
        RECT 40.415 100.755 40.895 101.095 ;
        RECT 41.065 100.585 41.320 101.130 ;
        RECT 41.490 100.755 41.765 101.455 ;
        RECT 41.935 100.585 44.525 101.675 ;
        RECT 45.340 101.555 46.765 101.725 ;
        RECT 45.340 101.380 45.730 101.555 ;
        RECT 46.215 100.585 46.545 101.385 ;
        RECT 46.935 101.375 47.250 102.395 ;
        RECT 47.455 102.395 47.835 102.480 ;
        RECT 48.345 102.395 48.675 102.920 ;
        RECT 48.935 102.605 49.145 103.135 ;
        RECT 49.420 102.685 50.205 102.855 ;
        RECT 50.375 102.685 50.780 102.855 ;
        RECT 47.455 102.355 47.680 102.395 ;
        RECT 47.455 101.775 47.625 102.355 ;
        RECT 48.345 102.225 48.545 102.395 ;
        RECT 49.420 102.225 49.590 102.685 ;
        RECT 47.795 101.895 48.545 102.225 ;
        RECT 48.715 101.895 49.590 102.225 ;
        RECT 47.455 101.725 47.670 101.775 ;
        RECT 47.455 101.645 47.845 101.725 ;
        RECT 46.715 100.755 47.250 101.375 ;
        RECT 47.515 100.800 47.845 101.645 ;
        RECT 48.355 101.690 48.545 101.895 ;
        RECT 48.015 100.585 48.185 101.595 ;
        RECT 48.355 101.315 49.250 101.690 ;
        RECT 48.355 100.755 48.695 101.315 ;
        RECT 48.925 100.585 49.240 101.085 ;
        RECT 49.420 101.055 49.590 101.895 ;
        RECT 49.760 102.185 50.225 102.515 ;
        RECT 50.610 102.455 50.780 102.685 ;
        RECT 50.960 102.635 51.330 103.135 ;
        RECT 51.650 102.685 52.325 102.855 ;
        RECT 52.520 102.685 52.855 102.855 ;
        RECT 49.760 101.225 50.080 102.185 ;
        RECT 50.610 102.155 51.440 102.455 ;
        RECT 50.250 101.255 50.440 101.975 ;
        RECT 50.610 101.085 50.780 102.155 ;
        RECT 51.240 102.125 51.440 102.155 ;
        RECT 50.950 101.905 51.120 101.975 ;
        RECT 51.650 101.905 51.820 102.685 ;
        RECT 52.685 102.545 52.855 102.685 ;
        RECT 53.025 102.675 53.275 103.135 ;
        RECT 50.950 101.735 51.820 101.905 ;
        RECT 51.990 102.265 52.515 102.485 ;
        RECT 52.685 102.415 52.910 102.545 ;
        RECT 50.950 101.645 51.460 101.735 ;
        RECT 49.420 100.885 50.305 101.055 ;
        RECT 50.530 100.755 50.780 101.085 ;
        RECT 50.950 100.585 51.120 101.385 ;
        RECT 51.290 101.030 51.460 101.645 ;
        RECT 51.990 101.565 52.160 102.265 ;
        RECT 51.630 101.200 52.160 101.565 ;
        RECT 52.330 101.500 52.570 102.095 ;
        RECT 52.740 101.310 52.910 102.415 ;
        RECT 53.080 101.555 53.360 102.505 ;
        RECT 52.605 101.180 52.910 101.310 ;
        RECT 51.290 100.860 52.395 101.030 ;
        RECT 52.605 100.755 52.855 101.180 ;
        RECT 53.025 100.585 53.290 101.045 ;
        RECT 53.530 100.755 53.715 102.875 ;
        RECT 53.885 102.755 54.215 103.135 ;
        RECT 54.385 102.585 54.555 102.875 ;
        RECT 54.815 102.590 60.160 103.135 ;
        RECT 53.890 102.415 54.555 102.585 ;
        RECT 53.890 101.425 54.120 102.415 ;
        RECT 54.290 101.595 54.640 102.245 ;
        RECT 56.400 101.760 56.740 102.590 ;
        RECT 60.335 102.365 63.845 103.135 ;
        RECT 64.935 102.410 65.225 103.135 ;
        RECT 65.395 102.590 70.740 103.135 ;
        RECT 53.890 101.255 54.555 101.425 ;
        RECT 53.885 100.585 54.215 101.085 ;
        RECT 54.385 100.755 54.555 101.255 ;
        RECT 58.220 101.020 58.570 102.270 ;
        RECT 60.335 101.845 61.985 102.365 ;
        RECT 62.155 101.675 63.845 102.195 ;
        RECT 66.980 101.760 67.320 102.590 ;
        RECT 70.915 102.365 73.505 103.135 ;
        RECT 54.815 100.585 60.160 101.020 ;
        RECT 60.335 100.585 63.845 101.675 ;
        RECT 64.935 100.585 65.225 101.750 ;
        RECT 68.800 101.020 69.150 102.270 ;
        RECT 70.915 101.845 72.125 102.365 ;
        RECT 74.135 102.335 74.475 102.965 ;
        RECT 74.645 102.335 74.895 103.135 ;
        RECT 75.085 102.485 75.415 102.965 ;
        RECT 75.585 102.675 75.810 103.135 ;
        RECT 75.980 102.485 76.310 102.965 ;
        RECT 72.295 101.675 73.505 102.195 ;
        RECT 65.395 100.585 70.740 101.020 ;
        RECT 70.915 100.585 73.505 101.675 ;
        RECT 74.135 101.725 74.310 102.335 ;
        RECT 75.085 102.315 76.310 102.485 ;
        RECT 76.940 102.355 77.440 102.965 ;
        RECT 77.850 102.395 78.465 102.965 ;
        RECT 78.635 102.625 78.850 103.135 ;
        RECT 79.080 102.625 79.360 102.955 ;
        RECT 79.540 102.625 79.780 103.135 ;
        RECT 74.480 101.975 75.175 102.145 ;
        RECT 75.005 101.725 75.175 101.975 ;
        RECT 75.350 101.945 75.770 102.145 ;
        RECT 75.940 101.945 76.270 102.145 ;
        RECT 76.440 101.945 76.770 102.145 ;
        RECT 76.940 101.725 77.110 102.355 ;
        RECT 77.295 101.895 77.645 102.145 ;
        RECT 74.135 100.755 74.475 101.725 ;
        RECT 74.645 100.585 74.815 101.725 ;
        RECT 75.005 101.555 77.440 101.725 ;
        RECT 75.085 100.585 75.335 101.385 ;
        RECT 75.980 100.755 76.310 101.555 ;
        RECT 76.610 100.585 76.940 101.385 ;
        RECT 77.110 100.755 77.440 101.555 ;
        RECT 77.850 101.375 78.165 102.395 ;
        RECT 78.335 101.725 78.505 102.225 ;
        RECT 78.755 101.895 79.020 102.455 ;
        RECT 79.190 101.725 79.360 102.625 ;
        RECT 79.530 101.895 79.885 102.455 ;
        RECT 80.115 102.365 82.705 103.135 ;
        RECT 80.115 101.845 81.325 102.365 ;
        RECT 78.335 101.555 79.760 101.725 ;
        RECT 81.495 101.675 82.705 102.195 ;
        RECT 77.850 100.755 78.385 101.375 ;
        RECT 78.555 100.585 78.885 101.385 ;
        RECT 79.370 101.380 79.760 101.555 ;
        RECT 80.115 100.585 82.705 101.675 ;
        RECT 82.880 101.535 83.215 102.955 ;
        RECT 83.395 102.765 84.140 103.135 ;
        RECT 84.705 102.595 84.960 102.955 ;
        RECT 85.140 102.765 85.470 103.135 ;
        RECT 85.650 102.595 85.875 102.955 ;
        RECT 83.390 102.405 85.875 102.595 ;
        RECT 83.390 101.715 83.615 102.405 ;
        RECT 86.555 102.335 86.895 102.965 ;
        RECT 87.065 102.335 87.315 103.135 ;
        RECT 87.505 102.485 87.835 102.965 ;
        RECT 88.005 102.675 88.230 103.135 ;
        RECT 88.400 102.485 88.730 102.965 ;
        RECT 83.815 101.895 84.095 102.225 ;
        RECT 84.275 101.895 84.850 102.225 ;
        RECT 85.030 101.895 85.465 102.225 ;
        RECT 85.645 101.895 85.915 102.225 ;
        RECT 86.555 101.725 86.730 102.335 ;
        RECT 87.505 102.315 88.730 102.485 ;
        RECT 89.360 102.355 89.860 102.965 ;
        RECT 90.695 102.410 90.985 103.135 ;
        RECT 91.155 102.590 96.500 103.135 ;
        RECT 86.900 101.975 87.595 102.145 ;
        RECT 87.425 101.725 87.595 101.975 ;
        RECT 87.770 101.945 88.190 102.145 ;
        RECT 88.360 101.945 88.690 102.145 ;
        RECT 88.860 101.945 89.190 102.145 ;
        RECT 89.360 101.725 89.530 102.355 ;
        RECT 89.715 101.895 90.065 102.145 ;
        RECT 92.740 101.760 93.080 102.590 ;
        RECT 96.675 102.365 98.345 103.135 ;
        RECT 98.605 102.585 98.775 102.875 ;
        RECT 98.945 102.755 99.275 103.135 ;
        RECT 98.605 102.415 99.270 102.585 ;
        RECT 83.390 101.535 85.885 101.715 ;
        RECT 82.880 100.765 83.145 101.535 ;
        RECT 83.315 100.585 83.645 101.305 ;
        RECT 83.835 101.125 85.025 101.355 ;
        RECT 83.835 100.765 84.095 101.125 ;
        RECT 84.265 100.585 84.595 100.955 ;
        RECT 84.765 100.765 85.025 101.125 ;
        RECT 85.595 100.765 85.885 101.535 ;
        RECT 86.555 100.755 86.895 101.725 ;
        RECT 87.065 100.585 87.235 101.725 ;
        RECT 87.425 101.555 89.860 101.725 ;
        RECT 87.505 100.585 87.755 101.385 ;
        RECT 88.400 100.755 88.730 101.555 ;
        RECT 89.030 100.585 89.360 101.385 ;
        RECT 89.530 100.755 89.860 101.555 ;
        RECT 90.695 100.585 90.985 101.750 ;
        RECT 94.560 101.020 94.910 102.270 ;
        RECT 96.675 101.845 97.425 102.365 ;
        RECT 97.595 101.675 98.345 102.195 ;
        RECT 91.155 100.585 96.500 101.020 ;
        RECT 96.675 100.585 98.345 101.675 ;
        RECT 98.520 101.595 98.870 102.245 ;
        RECT 99.040 101.425 99.270 102.415 ;
        RECT 98.605 101.255 99.270 101.425 ;
        RECT 98.605 100.755 98.775 101.255 ;
        RECT 98.945 100.585 99.275 101.085 ;
        RECT 99.445 100.755 99.630 102.875 ;
        RECT 99.885 102.675 100.135 103.135 ;
        RECT 100.305 102.685 100.640 102.855 ;
        RECT 100.835 102.685 101.510 102.855 ;
        RECT 100.305 102.545 100.475 102.685 ;
        RECT 99.800 101.555 100.080 102.505 ;
        RECT 100.250 102.415 100.475 102.545 ;
        RECT 100.250 101.310 100.420 102.415 ;
        RECT 100.645 102.265 101.170 102.485 ;
        RECT 100.590 101.500 100.830 102.095 ;
        RECT 101.000 101.565 101.170 102.265 ;
        RECT 101.340 101.905 101.510 102.685 ;
        RECT 101.830 102.635 102.200 103.135 ;
        RECT 102.380 102.685 102.785 102.855 ;
        RECT 102.955 102.685 103.740 102.855 ;
        RECT 102.380 102.455 102.550 102.685 ;
        RECT 101.720 102.155 102.550 102.455 ;
        RECT 102.935 102.185 103.400 102.515 ;
        RECT 101.720 102.125 101.920 102.155 ;
        RECT 102.040 101.905 102.210 101.975 ;
        RECT 101.340 101.735 102.210 101.905 ;
        RECT 101.700 101.645 102.210 101.735 ;
        RECT 100.250 101.180 100.555 101.310 ;
        RECT 101.000 101.200 101.530 101.565 ;
        RECT 99.870 100.585 100.135 101.045 ;
        RECT 100.305 100.755 100.555 101.180 ;
        RECT 101.700 101.030 101.870 101.645 ;
        RECT 100.765 100.860 101.870 101.030 ;
        RECT 102.040 100.585 102.210 101.385 ;
        RECT 102.380 101.085 102.550 102.155 ;
        RECT 102.720 101.255 102.910 101.975 ;
        RECT 103.080 101.225 103.400 102.185 ;
        RECT 103.570 102.225 103.740 102.685 ;
        RECT 104.015 102.605 104.225 103.135 ;
        RECT 104.485 102.395 104.815 102.920 ;
        RECT 104.985 102.525 105.155 103.135 ;
        RECT 105.325 102.480 105.655 102.915 ;
        RECT 105.325 102.395 105.705 102.480 ;
        RECT 104.615 102.225 104.815 102.395 ;
        RECT 105.480 102.355 105.705 102.395 ;
        RECT 103.570 101.895 104.445 102.225 ;
        RECT 104.615 101.895 105.365 102.225 ;
        RECT 102.380 100.755 102.630 101.085 ;
        RECT 103.570 101.055 103.740 101.895 ;
        RECT 104.615 101.690 104.805 101.895 ;
        RECT 105.535 101.775 105.705 102.355 ;
        RECT 105.875 102.365 107.545 103.135 ;
        RECT 107.715 102.635 107.975 102.965 ;
        RECT 108.145 102.775 108.475 103.135 ;
        RECT 108.730 102.755 110.030 102.965 ;
        RECT 105.875 101.845 106.625 102.365 ;
        RECT 105.490 101.725 105.705 101.775 ;
        RECT 103.910 101.315 104.805 101.690 ;
        RECT 105.315 101.645 105.705 101.725 ;
        RECT 106.795 101.675 107.545 102.195 ;
        RECT 102.855 100.885 103.740 101.055 ;
        RECT 103.920 100.585 104.235 101.085 ;
        RECT 104.465 100.755 104.805 101.315 ;
        RECT 104.975 100.585 105.145 101.595 ;
        RECT 105.315 100.800 105.645 101.645 ;
        RECT 105.875 100.585 107.545 101.675 ;
        RECT 107.715 101.435 107.885 102.635 ;
        RECT 108.730 102.605 108.900 102.755 ;
        RECT 108.145 102.480 108.900 102.605 ;
        RECT 108.055 102.435 108.900 102.480 ;
        RECT 108.055 102.315 108.325 102.435 ;
        RECT 108.055 101.740 108.225 102.315 ;
        RECT 108.455 101.875 108.865 102.180 ;
        RECT 109.155 102.145 109.365 102.545 ;
        RECT 109.035 101.935 109.365 102.145 ;
        RECT 109.610 102.145 109.830 102.545 ;
        RECT 110.305 102.370 110.760 103.135 ;
        RECT 110.935 102.365 112.605 103.135 ;
        RECT 109.610 101.935 110.085 102.145 ;
        RECT 110.275 101.945 110.765 102.145 ;
        RECT 110.935 101.845 111.685 102.365 ;
        RECT 112.775 102.335 113.115 102.965 ;
        RECT 113.285 102.335 113.535 103.135 ;
        RECT 113.725 102.485 114.055 102.965 ;
        RECT 114.225 102.675 114.450 103.135 ;
        RECT 114.620 102.485 114.950 102.965 ;
        RECT 108.055 101.705 108.255 101.740 ;
        RECT 109.585 101.705 110.760 101.765 ;
        RECT 108.055 101.595 110.760 101.705 ;
        RECT 111.855 101.675 112.605 102.195 ;
        RECT 108.115 101.535 109.915 101.595 ;
        RECT 109.585 101.505 109.915 101.535 ;
        RECT 107.715 100.755 107.975 101.435 ;
        RECT 108.145 100.585 108.395 101.365 ;
        RECT 108.645 101.335 109.480 101.345 ;
        RECT 110.070 101.335 110.255 101.425 ;
        RECT 108.645 101.135 110.255 101.335 ;
        RECT 108.645 100.755 108.895 101.135 ;
        RECT 110.025 101.095 110.255 101.135 ;
        RECT 110.505 100.975 110.760 101.595 ;
        RECT 109.065 100.585 109.420 100.965 ;
        RECT 110.425 100.755 110.760 100.975 ;
        RECT 110.935 100.585 112.605 101.675 ;
        RECT 112.775 101.775 112.950 102.335 ;
        RECT 113.725 102.315 114.950 102.485 ;
        RECT 115.580 102.355 116.080 102.965 ;
        RECT 116.455 102.410 116.745 103.135 ;
        RECT 117.005 102.585 117.175 102.875 ;
        RECT 117.345 102.755 117.675 103.135 ;
        RECT 117.005 102.415 117.670 102.585 ;
        RECT 113.120 101.975 113.815 102.145 ;
        RECT 112.775 101.725 113.005 101.775 ;
        RECT 113.645 101.725 113.815 101.975 ;
        RECT 113.990 101.945 114.410 102.145 ;
        RECT 114.580 101.945 114.910 102.145 ;
        RECT 115.080 101.945 115.410 102.145 ;
        RECT 115.580 101.725 115.750 102.355 ;
        RECT 115.935 101.895 116.285 102.145 ;
        RECT 112.775 100.755 113.115 101.725 ;
        RECT 113.285 100.585 113.455 101.725 ;
        RECT 113.645 101.555 116.080 101.725 ;
        RECT 113.725 100.585 113.975 101.385 ;
        RECT 114.620 100.755 114.950 101.555 ;
        RECT 115.250 100.585 115.580 101.385 ;
        RECT 115.750 100.755 116.080 101.555 ;
        RECT 116.455 100.585 116.745 101.750 ;
        RECT 116.920 101.595 117.270 102.245 ;
        RECT 117.440 101.425 117.670 102.415 ;
        RECT 117.005 101.255 117.670 101.425 ;
        RECT 117.005 100.755 117.175 101.255 ;
        RECT 117.345 100.585 117.675 101.085 ;
        RECT 117.845 100.755 118.030 102.875 ;
        RECT 118.285 102.675 118.535 103.135 ;
        RECT 118.705 102.685 119.040 102.855 ;
        RECT 119.235 102.685 119.910 102.855 ;
        RECT 118.705 102.545 118.875 102.685 ;
        RECT 118.200 101.555 118.480 102.505 ;
        RECT 118.650 102.415 118.875 102.545 ;
        RECT 118.650 101.310 118.820 102.415 ;
        RECT 119.045 102.265 119.570 102.485 ;
        RECT 118.990 101.500 119.230 102.095 ;
        RECT 119.400 101.565 119.570 102.265 ;
        RECT 119.740 101.905 119.910 102.685 ;
        RECT 120.230 102.635 120.600 103.135 ;
        RECT 120.780 102.685 121.185 102.855 ;
        RECT 121.355 102.685 122.140 102.855 ;
        RECT 120.780 102.455 120.950 102.685 ;
        RECT 120.120 102.155 120.950 102.455 ;
        RECT 121.335 102.185 121.800 102.515 ;
        RECT 120.120 102.125 120.320 102.155 ;
        RECT 120.440 101.905 120.610 101.975 ;
        RECT 119.740 101.735 120.610 101.905 ;
        RECT 120.100 101.645 120.610 101.735 ;
        RECT 118.650 101.180 118.955 101.310 ;
        RECT 119.400 101.200 119.930 101.565 ;
        RECT 118.270 100.585 118.535 101.045 ;
        RECT 118.705 100.755 118.955 101.180 ;
        RECT 120.100 101.030 120.270 101.645 ;
        RECT 119.165 100.860 120.270 101.030 ;
        RECT 120.440 100.585 120.610 101.385 ;
        RECT 120.780 101.085 120.950 102.155 ;
        RECT 121.120 101.255 121.310 101.975 ;
        RECT 121.480 101.225 121.800 102.185 ;
        RECT 121.970 102.225 122.140 102.685 ;
        RECT 122.415 102.605 122.625 103.135 ;
        RECT 122.885 102.395 123.215 102.920 ;
        RECT 123.385 102.525 123.555 103.135 ;
        RECT 123.725 102.480 124.055 102.915 ;
        RECT 123.725 102.395 124.105 102.480 ;
        RECT 123.015 102.225 123.215 102.395 ;
        RECT 123.880 102.355 124.105 102.395 ;
        RECT 124.940 102.355 125.440 102.965 ;
        RECT 121.970 101.895 122.845 102.225 ;
        RECT 123.015 101.895 123.765 102.225 ;
        RECT 120.780 100.755 121.030 101.085 ;
        RECT 121.970 101.055 122.140 101.895 ;
        RECT 123.015 101.690 123.205 101.895 ;
        RECT 123.935 101.775 124.105 102.355 ;
        RECT 124.735 101.895 125.085 102.145 ;
        RECT 123.890 101.725 124.105 101.775 ;
        RECT 125.270 101.725 125.440 102.355 ;
        RECT 126.070 102.485 126.400 102.965 ;
        RECT 126.570 102.675 126.795 103.135 ;
        RECT 126.965 102.485 127.295 102.965 ;
        RECT 126.070 102.315 127.295 102.485 ;
        RECT 127.485 102.335 127.735 103.135 ;
        RECT 127.905 102.335 128.245 102.965 ;
        RECT 128.505 102.585 128.675 102.875 ;
        RECT 128.845 102.755 129.175 103.135 ;
        RECT 128.505 102.415 129.170 102.585 ;
        RECT 125.610 101.945 125.940 102.145 ;
        RECT 126.110 101.945 126.440 102.145 ;
        RECT 126.610 101.945 127.030 102.145 ;
        RECT 127.205 101.975 127.900 102.145 ;
        RECT 127.205 101.725 127.375 101.975 ;
        RECT 128.070 101.725 128.245 102.335 ;
        RECT 122.310 101.315 123.205 101.690 ;
        RECT 123.715 101.645 124.105 101.725 ;
        RECT 121.255 100.885 122.140 101.055 ;
        RECT 122.320 100.585 122.635 101.085 ;
        RECT 122.865 100.755 123.205 101.315 ;
        RECT 123.375 100.585 123.545 101.595 ;
        RECT 123.715 100.800 124.045 101.645 ;
        RECT 124.940 101.555 127.375 101.725 ;
        RECT 124.940 100.755 125.270 101.555 ;
        RECT 125.440 100.585 125.770 101.385 ;
        RECT 126.070 100.755 126.400 101.555 ;
        RECT 127.045 100.585 127.295 101.385 ;
        RECT 127.565 100.585 127.735 101.725 ;
        RECT 127.905 100.755 128.245 101.725 ;
        RECT 128.420 101.595 128.770 102.245 ;
        RECT 128.940 101.425 129.170 102.415 ;
        RECT 128.505 101.255 129.170 101.425 ;
        RECT 128.505 100.755 128.675 101.255 ;
        RECT 128.845 100.585 129.175 101.085 ;
        RECT 129.345 100.755 129.530 102.875 ;
        RECT 129.785 102.675 130.035 103.135 ;
        RECT 130.205 102.685 130.540 102.855 ;
        RECT 130.735 102.685 131.410 102.855 ;
        RECT 130.205 102.545 130.375 102.685 ;
        RECT 129.700 101.555 129.980 102.505 ;
        RECT 130.150 102.415 130.375 102.545 ;
        RECT 130.150 101.310 130.320 102.415 ;
        RECT 130.545 102.265 131.070 102.485 ;
        RECT 130.490 101.500 130.730 102.095 ;
        RECT 130.900 101.565 131.070 102.265 ;
        RECT 131.240 101.905 131.410 102.685 ;
        RECT 131.730 102.635 132.100 103.135 ;
        RECT 132.280 102.685 132.685 102.855 ;
        RECT 132.855 102.685 133.640 102.855 ;
        RECT 132.280 102.455 132.450 102.685 ;
        RECT 131.620 102.155 132.450 102.455 ;
        RECT 132.835 102.185 133.300 102.515 ;
        RECT 131.620 102.125 131.820 102.155 ;
        RECT 131.940 101.905 132.110 101.975 ;
        RECT 131.240 101.735 132.110 101.905 ;
        RECT 131.600 101.645 132.110 101.735 ;
        RECT 130.150 101.180 130.455 101.310 ;
        RECT 130.900 101.200 131.430 101.565 ;
        RECT 129.770 100.585 130.035 101.045 ;
        RECT 130.205 100.755 130.455 101.180 ;
        RECT 131.600 101.030 131.770 101.645 ;
        RECT 130.665 100.860 131.770 101.030 ;
        RECT 131.940 100.585 132.110 101.385 ;
        RECT 132.280 101.085 132.450 102.155 ;
        RECT 132.620 101.255 132.810 101.975 ;
        RECT 132.980 101.225 133.300 102.185 ;
        RECT 133.470 102.225 133.640 102.685 ;
        RECT 133.915 102.605 134.125 103.135 ;
        RECT 134.385 102.395 134.715 102.920 ;
        RECT 134.885 102.525 135.055 103.135 ;
        RECT 135.225 102.480 135.555 102.915 ;
        RECT 135.865 102.585 136.035 102.965 ;
        RECT 136.250 102.755 136.580 103.135 ;
        RECT 135.225 102.395 135.605 102.480 ;
        RECT 135.865 102.415 136.580 102.585 ;
        RECT 134.515 102.225 134.715 102.395 ;
        RECT 135.380 102.355 135.605 102.395 ;
        RECT 133.470 101.895 134.345 102.225 ;
        RECT 134.515 101.895 135.265 102.225 ;
        RECT 132.280 100.755 132.530 101.085 ;
        RECT 133.470 101.055 133.640 101.895 ;
        RECT 134.515 101.690 134.705 101.895 ;
        RECT 135.435 101.775 135.605 102.355 ;
        RECT 135.775 101.865 136.130 102.235 ;
        RECT 136.410 102.225 136.580 102.415 ;
        RECT 136.750 102.390 137.005 102.965 ;
        RECT 136.410 101.895 136.665 102.225 ;
        RECT 135.390 101.725 135.605 101.775 ;
        RECT 133.810 101.315 134.705 101.690 ;
        RECT 135.215 101.645 135.605 101.725 ;
        RECT 136.410 101.685 136.580 101.895 ;
        RECT 132.755 100.885 133.640 101.055 ;
        RECT 133.820 100.585 134.135 101.085 ;
        RECT 134.365 100.755 134.705 101.315 ;
        RECT 134.875 100.585 135.045 101.595 ;
        RECT 135.215 100.800 135.545 101.645 ;
        RECT 135.865 101.515 136.580 101.685 ;
        RECT 136.835 101.660 137.005 102.390 ;
        RECT 137.180 102.295 137.440 103.135 ;
        RECT 137.615 102.385 138.825 103.135 ;
        RECT 135.865 100.755 136.035 101.515 ;
        RECT 136.250 100.585 136.580 101.345 ;
        RECT 136.750 100.755 137.005 101.660 ;
        RECT 137.180 100.585 137.440 101.735 ;
        RECT 137.615 101.675 138.135 102.215 ;
        RECT 138.305 101.845 138.825 102.385 ;
        RECT 137.615 100.585 138.825 101.675 ;
        RECT 13.330 100.415 138.910 100.585 ;
        RECT 13.415 99.325 14.625 100.415 ;
        RECT 14.795 99.325 18.305 100.415 ;
        RECT 18.565 99.745 18.735 100.245 ;
        RECT 18.905 99.915 19.235 100.415 ;
        RECT 18.565 99.575 19.230 99.745 ;
        RECT 13.415 98.615 13.935 99.155 ;
        RECT 14.105 98.785 14.625 99.325 ;
        RECT 14.795 98.635 16.445 99.155 ;
        RECT 16.615 98.805 18.305 99.325 ;
        RECT 18.480 98.755 18.830 99.405 ;
        RECT 13.415 97.865 14.625 98.615 ;
        RECT 14.795 97.865 18.305 98.635 ;
        RECT 19.000 98.585 19.230 99.575 ;
        RECT 18.565 98.415 19.230 98.585 ;
        RECT 18.565 98.125 18.735 98.415 ;
        RECT 18.905 97.865 19.235 98.245 ;
        RECT 19.405 98.125 19.590 100.245 ;
        RECT 19.830 99.955 20.095 100.415 ;
        RECT 20.265 99.820 20.515 100.245 ;
        RECT 20.725 99.970 21.830 100.140 ;
        RECT 20.210 99.690 20.515 99.820 ;
        RECT 19.760 98.495 20.040 99.445 ;
        RECT 20.210 98.585 20.380 99.690 ;
        RECT 20.550 98.905 20.790 99.500 ;
        RECT 20.960 99.435 21.490 99.800 ;
        RECT 20.960 98.735 21.130 99.435 ;
        RECT 21.660 99.355 21.830 99.970 ;
        RECT 22.000 99.615 22.170 100.415 ;
        RECT 22.340 99.915 22.590 100.245 ;
        RECT 22.815 99.945 23.700 100.115 ;
        RECT 21.660 99.265 22.170 99.355 ;
        RECT 20.210 98.455 20.435 98.585 ;
        RECT 20.605 98.515 21.130 98.735 ;
        RECT 21.300 99.095 22.170 99.265 ;
        RECT 19.845 97.865 20.095 98.325 ;
        RECT 20.265 98.315 20.435 98.455 ;
        RECT 21.300 98.315 21.470 99.095 ;
        RECT 22.000 99.025 22.170 99.095 ;
        RECT 21.680 98.845 21.880 98.875 ;
        RECT 22.340 98.845 22.510 99.915 ;
        RECT 22.680 99.025 22.870 99.745 ;
        RECT 21.680 98.545 22.510 98.845 ;
        RECT 23.040 98.815 23.360 99.775 ;
        RECT 20.265 98.145 20.600 98.315 ;
        RECT 20.795 98.145 21.470 98.315 ;
        RECT 21.790 97.865 22.160 98.365 ;
        RECT 22.340 98.315 22.510 98.545 ;
        RECT 22.895 98.485 23.360 98.815 ;
        RECT 23.530 99.105 23.700 99.945 ;
        RECT 23.880 99.915 24.195 100.415 ;
        RECT 24.425 99.685 24.765 100.245 ;
        RECT 23.870 99.310 24.765 99.685 ;
        RECT 24.935 99.405 25.105 100.415 ;
        RECT 24.575 99.105 24.765 99.310 ;
        RECT 25.275 99.355 25.605 100.200 ;
        RECT 25.275 99.275 25.665 99.355 ;
        RECT 25.450 99.225 25.665 99.275 ;
        RECT 26.295 99.250 26.585 100.415 ;
        RECT 26.755 99.980 32.100 100.415 ;
        RECT 32.275 99.980 37.620 100.415 ;
        RECT 37.795 99.980 43.140 100.415 ;
        RECT 43.315 99.980 48.660 100.415 ;
        RECT 23.530 98.775 24.405 99.105 ;
        RECT 24.575 98.775 25.325 99.105 ;
        RECT 23.530 98.315 23.700 98.775 ;
        RECT 24.575 98.605 24.775 98.775 ;
        RECT 25.495 98.645 25.665 99.225 ;
        RECT 25.440 98.605 25.665 98.645 ;
        RECT 22.340 98.145 22.745 98.315 ;
        RECT 22.915 98.145 23.700 98.315 ;
        RECT 23.975 97.865 24.185 98.395 ;
        RECT 24.445 98.080 24.775 98.605 ;
        RECT 25.285 98.520 25.665 98.605 ;
        RECT 24.945 97.865 25.115 98.475 ;
        RECT 25.285 98.085 25.615 98.520 ;
        RECT 26.295 97.865 26.585 98.590 ;
        RECT 28.340 98.410 28.680 99.240 ;
        RECT 30.160 98.730 30.510 99.980 ;
        RECT 33.860 98.410 34.200 99.240 ;
        RECT 35.680 98.730 36.030 99.980 ;
        RECT 39.380 98.410 39.720 99.240 ;
        RECT 41.200 98.730 41.550 99.980 ;
        RECT 44.900 98.410 45.240 99.240 ;
        RECT 46.720 98.730 47.070 99.980 ;
        RECT 48.835 99.275 49.095 100.415 ;
        RECT 49.265 99.265 49.595 100.245 ;
        RECT 49.765 99.275 50.045 100.415 ;
        RECT 50.215 99.325 51.885 100.415 ;
        RECT 48.855 98.855 49.190 99.105 ;
        RECT 49.360 98.665 49.530 99.265 ;
        RECT 49.700 98.835 50.035 99.105 ;
        RECT 26.755 97.865 32.100 98.410 ;
        RECT 32.275 97.865 37.620 98.410 ;
        RECT 37.795 97.865 43.140 98.410 ;
        RECT 43.315 97.865 48.660 98.410 ;
        RECT 48.835 98.035 49.530 98.665 ;
        RECT 49.735 97.865 50.045 98.665 ;
        RECT 50.215 98.635 50.965 99.155 ;
        RECT 51.135 98.805 51.885 99.325 ;
        RECT 52.055 99.250 52.345 100.415 ;
        RECT 52.515 99.980 57.860 100.415 ;
        RECT 58.035 99.980 63.380 100.415 ;
        RECT 63.555 99.980 68.900 100.415 ;
        RECT 50.215 97.865 51.885 98.635 ;
        RECT 52.055 97.865 52.345 98.590 ;
        RECT 54.100 98.410 54.440 99.240 ;
        RECT 55.920 98.730 56.270 99.980 ;
        RECT 59.620 98.410 59.960 99.240 ;
        RECT 61.440 98.730 61.790 99.980 ;
        RECT 65.140 98.410 65.480 99.240 ;
        RECT 66.960 98.730 67.310 99.980 ;
        RECT 69.075 99.325 70.285 100.415 ;
        RECT 70.545 99.745 70.715 100.245 ;
        RECT 70.885 99.915 71.215 100.415 ;
        RECT 70.545 99.575 71.210 99.745 ;
        RECT 69.075 98.615 69.595 99.155 ;
        RECT 69.765 98.785 70.285 99.325 ;
        RECT 70.460 98.755 70.810 99.405 ;
        RECT 52.515 97.865 57.860 98.410 ;
        RECT 58.035 97.865 63.380 98.410 ;
        RECT 63.555 97.865 68.900 98.410 ;
        RECT 69.075 97.865 70.285 98.615 ;
        RECT 70.980 98.585 71.210 99.575 ;
        RECT 70.545 98.415 71.210 98.585 ;
        RECT 70.545 98.125 70.715 98.415 ;
        RECT 70.885 97.865 71.215 98.245 ;
        RECT 71.385 98.125 71.570 100.245 ;
        RECT 71.810 99.955 72.075 100.415 ;
        RECT 72.245 99.820 72.495 100.245 ;
        RECT 72.705 99.970 73.810 100.140 ;
        RECT 72.190 99.690 72.495 99.820 ;
        RECT 71.740 98.495 72.020 99.445 ;
        RECT 72.190 98.585 72.360 99.690 ;
        RECT 72.530 98.905 72.770 99.500 ;
        RECT 72.940 99.435 73.470 99.800 ;
        RECT 72.940 98.735 73.110 99.435 ;
        RECT 73.640 99.355 73.810 99.970 ;
        RECT 73.980 99.615 74.150 100.415 ;
        RECT 74.320 99.915 74.570 100.245 ;
        RECT 74.795 99.945 75.680 100.115 ;
        RECT 73.640 99.265 74.150 99.355 ;
        RECT 72.190 98.455 72.415 98.585 ;
        RECT 72.585 98.515 73.110 98.735 ;
        RECT 73.280 99.095 74.150 99.265 ;
        RECT 71.825 97.865 72.075 98.325 ;
        RECT 72.245 98.315 72.415 98.455 ;
        RECT 73.280 98.315 73.450 99.095 ;
        RECT 73.980 99.025 74.150 99.095 ;
        RECT 73.660 98.845 73.860 98.875 ;
        RECT 74.320 98.845 74.490 99.915 ;
        RECT 74.660 99.025 74.850 99.745 ;
        RECT 73.660 98.545 74.490 98.845 ;
        RECT 75.020 98.815 75.340 99.775 ;
        RECT 72.245 98.145 72.580 98.315 ;
        RECT 72.775 98.145 73.450 98.315 ;
        RECT 73.770 97.865 74.140 98.365 ;
        RECT 74.320 98.315 74.490 98.545 ;
        RECT 74.875 98.485 75.340 98.815 ;
        RECT 75.510 99.105 75.680 99.945 ;
        RECT 75.860 99.915 76.175 100.415 ;
        RECT 76.405 99.685 76.745 100.245 ;
        RECT 75.850 99.310 76.745 99.685 ;
        RECT 76.915 99.405 77.085 100.415 ;
        RECT 76.555 99.105 76.745 99.310 ;
        RECT 77.255 99.355 77.585 100.200 ;
        RECT 77.255 99.275 77.645 99.355 ;
        RECT 77.430 99.225 77.645 99.275 ;
        RECT 77.815 99.250 78.105 100.415 ;
        RECT 78.275 99.275 78.615 100.245 ;
        RECT 78.785 99.275 78.955 100.415 ;
        RECT 79.225 99.615 79.475 100.415 ;
        RECT 80.120 99.445 80.450 100.245 ;
        RECT 80.750 99.615 81.080 100.415 ;
        RECT 81.250 99.445 81.580 100.245 ;
        RECT 79.145 99.275 81.580 99.445 ;
        RECT 82.505 99.485 82.675 100.245 ;
        RECT 82.890 99.655 83.220 100.415 ;
        RECT 82.505 99.315 83.220 99.485 ;
        RECT 83.390 99.340 83.645 100.245 ;
        RECT 75.510 98.775 76.385 99.105 ;
        RECT 76.555 98.775 77.305 99.105 ;
        RECT 75.510 98.315 75.680 98.775 ;
        RECT 76.555 98.605 76.755 98.775 ;
        RECT 77.475 98.645 77.645 99.225 ;
        RECT 77.420 98.605 77.645 98.645 ;
        RECT 74.320 98.145 74.725 98.315 ;
        RECT 74.895 98.145 75.680 98.315 ;
        RECT 75.955 97.865 76.165 98.395 ;
        RECT 76.425 98.080 76.755 98.605 ;
        RECT 77.265 98.520 77.645 98.605 ;
        RECT 78.275 98.665 78.450 99.275 ;
        RECT 79.145 99.025 79.315 99.275 ;
        RECT 78.620 98.855 79.315 99.025 ;
        RECT 79.490 98.855 79.910 99.055 ;
        RECT 80.080 98.855 80.410 99.055 ;
        RECT 80.580 98.855 80.910 99.055 ;
        RECT 76.925 97.865 77.095 98.475 ;
        RECT 77.265 98.085 77.595 98.520 ;
        RECT 77.815 97.865 78.105 98.590 ;
        RECT 78.275 98.035 78.615 98.665 ;
        RECT 78.785 97.865 79.035 98.665 ;
        RECT 79.225 98.515 80.450 98.685 ;
        RECT 79.225 98.035 79.555 98.515 ;
        RECT 79.725 97.865 79.950 98.325 ;
        RECT 80.120 98.035 80.450 98.515 ;
        RECT 81.080 98.645 81.250 99.275 ;
        RECT 81.435 98.855 81.785 99.105 ;
        RECT 82.415 98.765 82.770 99.135 ;
        RECT 83.050 99.105 83.220 99.315 ;
        RECT 83.050 98.775 83.305 99.105 ;
        RECT 81.080 98.035 81.580 98.645 ;
        RECT 83.050 98.585 83.220 98.775 ;
        RECT 83.475 98.610 83.645 99.340 ;
        RECT 83.820 99.265 84.080 100.415 ;
        RECT 84.255 99.325 86.845 100.415 ;
        RECT 82.505 98.415 83.220 98.585 ;
        RECT 82.505 98.035 82.675 98.415 ;
        RECT 82.890 97.865 83.220 98.245 ;
        RECT 83.390 98.035 83.645 98.610 ;
        RECT 83.820 97.865 84.080 98.705 ;
        RECT 84.255 98.635 85.465 99.155 ;
        RECT 85.635 98.805 86.845 99.325 ;
        RECT 87.015 99.565 87.275 100.245 ;
        RECT 87.445 99.635 87.695 100.415 ;
        RECT 87.945 99.865 88.195 100.245 ;
        RECT 88.365 100.035 88.720 100.415 ;
        RECT 89.725 100.025 90.060 100.245 ;
        RECT 89.325 99.865 89.555 99.905 ;
        RECT 87.945 99.665 89.555 99.865 ;
        RECT 87.945 99.655 88.780 99.665 ;
        RECT 89.370 99.575 89.555 99.665 ;
        RECT 84.255 97.865 86.845 98.635 ;
        RECT 87.015 98.365 87.185 99.565 ;
        RECT 88.885 99.465 89.215 99.495 ;
        RECT 87.415 99.405 89.215 99.465 ;
        RECT 89.805 99.405 90.060 100.025 ;
        RECT 90.235 99.980 95.580 100.415 ;
        RECT 87.355 99.295 90.060 99.405 ;
        RECT 87.355 99.260 87.555 99.295 ;
        RECT 87.355 98.685 87.525 99.260 ;
        RECT 88.885 99.235 90.060 99.295 ;
        RECT 87.755 98.820 88.165 99.125 ;
        RECT 88.335 98.855 88.665 99.065 ;
        RECT 87.355 98.565 87.625 98.685 ;
        RECT 87.355 98.520 88.200 98.565 ;
        RECT 87.445 98.395 88.200 98.520 ;
        RECT 88.455 98.455 88.665 98.855 ;
        RECT 88.910 98.855 89.385 99.065 ;
        RECT 89.575 98.855 90.065 99.055 ;
        RECT 88.910 98.455 89.130 98.855 ;
        RECT 87.015 98.035 87.275 98.365 ;
        RECT 88.030 98.245 88.200 98.395 ;
        RECT 87.445 97.865 87.775 98.225 ;
        RECT 88.030 98.035 89.330 98.245 ;
        RECT 89.605 97.865 90.060 98.630 ;
        RECT 91.820 98.410 92.160 99.240 ;
        RECT 93.640 98.730 93.990 99.980 ;
        RECT 95.755 99.325 97.425 100.415 ;
        RECT 95.755 98.635 96.505 99.155 ;
        RECT 96.675 98.805 97.425 99.325 ;
        RECT 98.055 99.275 98.395 100.245 ;
        RECT 98.565 99.275 98.735 100.415 ;
        RECT 99.005 99.615 99.255 100.415 ;
        RECT 99.900 99.445 100.230 100.245 ;
        RECT 100.530 99.615 100.860 100.415 ;
        RECT 101.030 99.445 101.360 100.245 ;
        RECT 98.925 99.275 101.360 99.445 ;
        RECT 98.055 98.665 98.230 99.275 ;
        RECT 98.925 99.025 99.095 99.275 ;
        RECT 98.400 98.855 99.095 99.025 ;
        RECT 99.270 98.855 99.690 99.055 ;
        RECT 99.860 98.855 100.190 99.055 ;
        RECT 100.360 98.855 100.690 99.055 ;
        RECT 90.235 97.865 95.580 98.410 ;
        RECT 95.755 97.865 97.425 98.635 ;
        RECT 98.055 98.035 98.395 98.665 ;
        RECT 98.565 97.865 98.815 98.665 ;
        RECT 99.005 98.515 100.230 98.685 ;
        RECT 99.005 98.035 99.335 98.515 ;
        RECT 99.505 97.865 99.730 98.325 ;
        RECT 99.900 98.035 100.230 98.515 ;
        RECT 100.860 98.645 101.030 99.275 ;
        RECT 101.740 99.265 102.000 100.415 ;
        RECT 102.175 99.340 102.430 100.245 ;
        RECT 102.600 99.655 102.930 100.415 ;
        RECT 103.145 99.485 103.315 100.245 ;
        RECT 101.215 98.855 101.565 99.105 ;
        RECT 100.860 98.035 101.360 98.645 ;
        RECT 101.740 97.865 102.000 98.705 ;
        RECT 102.175 98.610 102.345 99.340 ;
        RECT 102.600 99.315 103.315 99.485 ;
        RECT 102.600 99.105 102.770 99.315 ;
        RECT 103.575 99.250 103.865 100.415 ;
        RECT 104.070 99.625 104.605 100.245 ;
        RECT 102.515 98.775 102.770 99.105 ;
        RECT 102.175 98.035 102.430 98.610 ;
        RECT 102.600 98.585 102.770 98.775 ;
        RECT 103.050 98.765 103.405 99.135 ;
        RECT 104.070 98.605 104.385 99.625 ;
        RECT 104.775 99.615 105.105 100.415 ;
        RECT 106.335 99.980 111.680 100.415 ;
        RECT 105.590 99.445 105.980 99.620 ;
        RECT 104.555 99.275 105.980 99.445 ;
        RECT 104.555 98.775 104.725 99.275 ;
        RECT 102.600 98.415 103.315 98.585 ;
        RECT 102.600 97.865 102.930 98.245 ;
        RECT 103.145 98.035 103.315 98.415 ;
        RECT 103.575 97.865 103.865 98.590 ;
        RECT 104.070 98.035 104.685 98.605 ;
        RECT 104.975 98.545 105.240 99.105 ;
        RECT 105.410 98.375 105.580 99.275 ;
        RECT 105.750 98.545 106.105 99.105 ;
        RECT 107.920 98.410 108.260 99.240 ;
        RECT 109.740 98.730 110.090 99.980 ;
        RECT 111.855 99.325 113.525 100.415 ;
        RECT 111.855 98.635 112.605 99.155 ;
        RECT 112.775 98.805 113.525 99.325 ;
        RECT 114.340 99.445 114.730 99.620 ;
        RECT 115.215 99.615 115.545 100.415 ;
        RECT 115.715 99.625 116.250 100.245 ;
        RECT 114.340 99.275 115.765 99.445 ;
        RECT 104.855 97.865 105.070 98.375 ;
        RECT 105.300 98.045 105.580 98.375 ;
        RECT 105.760 97.865 106.000 98.375 ;
        RECT 106.335 97.865 111.680 98.410 ;
        RECT 111.855 97.865 113.525 98.635 ;
        RECT 114.215 98.545 114.570 99.105 ;
        RECT 114.740 98.375 114.910 99.275 ;
        RECT 115.080 98.545 115.345 99.105 ;
        RECT 115.595 98.775 115.765 99.275 ;
        RECT 115.935 98.605 116.250 99.625 ;
        RECT 116.545 99.485 116.715 100.245 ;
        RECT 116.930 99.655 117.260 100.415 ;
        RECT 116.545 99.315 117.260 99.485 ;
        RECT 117.430 99.340 117.685 100.245 ;
        RECT 116.455 98.765 116.810 99.135 ;
        RECT 117.090 99.105 117.260 99.315 ;
        RECT 117.090 98.775 117.345 99.105 ;
        RECT 114.320 97.865 114.560 98.375 ;
        RECT 114.740 98.045 115.020 98.375 ;
        RECT 115.250 97.865 115.465 98.375 ;
        RECT 115.635 98.035 116.250 98.605 ;
        RECT 117.090 98.585 117.260 98.775 ;
        RECT 117.515 98.610 117.685 99.340 ;
        RECT 117.860 99.265 118.120 100.415 ;
        RECT 118.295 99.980 123.640 100.415 ;
        RECT 116.545 98.415 117.260 98.585 ;
        RECT 116.545 98.035 116.715 98.415 ;
        RECT 116.930 97.865 117.260 98.245 ;
        RECT 117.430 98.035 117.685 98.610 ;
        RECT 117.860 97.865 118.120 98.705 ;
        RECT 119.880 98.410 120.220 99.240 ;
        RECT 121.700 98.730 122.050 99.980 ;
        RECT 123.815 99.325 125.485 100.415 ;
        RECT 123.815 98.635 124.565 99.155 ;
        RECT 124.735 98.805 125.485 99.325 ;
        RECT 125.860 99.445 126.190 100.245 ;
        RECT 126.360 99.615 126.690 100.415 ;
        RECT 126.990 99.445 127.320 100.245 ;
        RECT 127.965 99.615 128.215 100.415 ;
        RECT 125.860 99.275 128.295 99.445 ;
        RECT 128.485 99.275 128.655 100.415 ;
        RECT 128.825 99.275 129.165 100.245 ;
        RECT 125.655 98.855 126.005 99.105 ;
        RECT 126.190 98.645 126.360 99.275 ;
        RECT 126.530 98.855 126.860 99.055 ;
        RECT 127.030 98.855 127.360 99.055 ;
        RECT 127.530 98.855 127.950 99.055 ;
        RECT 128.125 99.025 128.295 99.275 ;
        RECT 128.125 98.855 128.820 99.025 ;
        RECT 128.990 98.715 129.165 99.275 ;
        RECT 129.335 99.250 129.625 100.415 ;
        RECT 129.885 99.745 130.055 100.245 ;
        RECT 130.225 99.915 130.555 100.415 ;
        RECT 129.885 99.575 130.550 99.745 ;
        RECT 129.800 98.755 130.150 99.405 ;
        RECT 118.295 97.865 123.640 98.410 ;
        RECT 123.815 97.865 125.485 98.635 ;
        RECT 125.860 98.035 126.360 98.645 ;
        RECT 126.990 98.515 128.215 98.685 ;
        RECT 128.935 98.665 129.165 98.715 ;
        RECT 126.990 98.035 127.320 98.515 ;
        RECT 127.490 97.865 127.715 98.325 ;
        RECT 127.885 98.035 128.215 98.515 ;
        RECT 128.405 97.865 128.655 98.665 ;
        RECT 128.825 98.035 129.165 98.665 ;
        RECT 129.335 97.865 129.625 98.590 ;
        RECT 130.320 98.585 130.550 99.575 ;
        RECT 129.885 98.415 130.550 98.585 ;
        RECT 129.885 98.125 130.055 98.415 ;
        RECT 130.225 97.865 130.555 98.245 ;
        RECT 130.725 98.125 130.910 100.245 ;
        RECT 131.150 99.955 131.415 100.415 ;
        RECT 131.585 99.820 131.835 100.245 ;
        RECT 132.045 99.970 133.150 100.140 ;
        RECT 131.530 99.690 131.835 99.820 ;
        RECT 131.080 98.495 131.360 99.445 ;
        RECT 131.530 98.585 131.700 99.690 ;
        RECT 131.870 98.905 132.110 99.500 ;
        RECT 132.280 99.435 132.810 99.800 ;
        RECT 132.280 98.735 132.450 99.435 ;
        RECT 132.980 99.355 133.150 99.970 ;
        RECT 133.320 99.615 133.490 100.415 ;
        RECT 133.660 99.915 133.910 100.245 ;
        RECT 134.135 99.945 135.020 100.115 ;
        RECT 132.980 99.265 133.490 99.355 ;
        RECT 131.530 98.455 131.755 98.585 ;
        RECT 131.925 98.515 132.450 98.735 ;
        RECT 132.620 99.095 133.490 99.265 ;
        RECT 131.165 97.865 131.415 98.325 ;
        RECT 131.585 98.315 131.755 98.455 ;
        RECT 132.620 98.315 132.790 99.095 ;
        RECT 133.320 99.025 133.490 99.095 ;
        RECT 133.000 98.845 133.200 98.875 ;
        RECT 133.660 98.845 133.830 99.915 ;
        RECT 134.000 99.025 134.190 99.745 ;
        RECT 133.000 98.545 133.830 98.845 ;
        RECT 134.360 98.815 134.680 99.775 ;
        RECT 131.585 98.145 131.920 98.315 ;
        RECT 132.115 98.145 132.790 98.315 ;
        RECT 133.110 97.865 133.480 98.365 ;
        RECT 133.660 98.315 133.830 98.545 ;
        RECT 134.215 98.485 134.680 98.815 ;
        RECT 134.850 99.105 135.020 99.945 ;
        RECT 135.200 99.915 135.515 100.415 ;
        RECT 135.745 99.685 136.085 100.245 ;
        RECT 135.190 99.310 136.085 99.685 ;
        RECT 136.255 99.405 136.425 100.415 ;
        RECT 135.895 99.105 136.085 99.310 ;
        RECT 136.595 99.355 136.925 100.200 ;
        RECT 136.595 99.275 136.985 99.355 ;
        RECT 136.770 99.225 136.985 99.275 ;
        RECT 134.850 98.775 135.725 99.105 ;
        RECT 135.895 98.775 136.645 99.105 ;
        RECT 134.850 98.315 135.020 98.775 ;
        RECT 135.895 98.605 136.095 98.775 ;
        RECT 136.815 98.645 136.985 99.225 ;
        RECT 137.615 99.325 138.825 100.415 ;
        RECT 137.615 98.785 138.135 99.325 ;
        RECT 136.760 98.605 136.985 98.645 ;
        RECT 138.305 98.615 138.825 99.155 ;
        RECT 133.660 98.145 134.065 98.315 ;
        RECT 134.235 98.145 135.020 98.315 ;
        RECT 135.295 97.865 135.505 98.395 ;
        RECT 135.765 98.080 136.095 98.605 ;
        RECT 136.605 98.520 136.985 98.605 ;
        RECT 136.265 97.865 136.435 98.475 ;
        RECT 136.605 98.085 136.935 98.520 ;
        RECT 137.615 97.865 138.825 98.615 ;
        RECT 13.330 97.695 138.910 97.865 ;
        RECT 13.415 96.945 14.625 97.695 ;
        RECT 14.795 97.150 20.140 97.695 ;
        RECT 20.315 97.150 25.660 97.695 ;
        RECT 25.835 97.150 31.180 97.695 ;
        RECT 31.355 97.150 36.700 97.695 ;
        RECT 13.415 96.405 13.935 96.945 ;
        RECT 14.105 96.235 14.625 96.775 ;
        RECT 16.380 96.320 16.720 97.150 ;
        RECT 13.415 95.145 14.625 96.235 ;
        RECT 18.200 95.580 18.550 96.830 ;
        RECT 21.900 96.320 22.240 97.150 ;
        RECT 23.720 95.580 24.070 96.830 ;
        RECT 27.420 96.320 27.760 97.150 ;
        RECT 29.240 95.580 29.590 96.830 ;
        RECT 32.940 96.320 33.280 97.150 ;
        RECT 36.875 96.925 38.545 97.695 ;
        RECT 39.175 96.970 39.465 97.695 ;
        RECT 39.635 97.150 44.980 97.695 ;
        RECT 45.155 97.150 50.500 97.695 ;
        RECT 50.675 97.150 56.020 97.695 ;
        RECT 56.195 97.150 61.540 97.695 ;
        RECT 34.760 95.580 35.110 96.830 ;
        RECT 36.875 96.405 37.625 96.925 ;
        RECT 37.795 96.235 38.545 96.755 ;
        RECT 41.220 96.320 41.560 97.150 ;
        RECT 14.795 95.145 20.140 95.580 ;
        RECT 20.315 95.145 25.660 95.580 ;
        RECT 25.835 95.145 31.180 95.580 ;
        RECT 31.355 95.145 36.700 95.580 ;
        RECT 36.875 95.145 38.545 96.235 ;
        RECT 39.175 95.145 39.465 96.310 ;
        RECT 43.040 95.580 43.390 96.830 ;
        RECT 46.740 96.320 47.080 97.150 ;
        RECT 48.560 95.580 48.910 96.830 ;
        RECT 52.260 96.320 52.600 97.150 ;
        RECT 54.080 95.580 54.430 96.830 ;
        RECT 57.780 96.320 58.120 97.150 ;
        RECT 61.715 96.925 64.305 97.695 ;
        RECT 64.935 96.970 65.225 97.695 ;
        RECT 65.395 97.150 70.740 97.695 ;
        RECT 59.600 95.580 59.950 96.830 ;
        RECT 61.715 96.405 62.925 96.925 ;
        RECT 63.095 96.235 64.305 96.755 ;
        RECT 66.980 96.320 67.320 97.150 ;
        RECT 71.005 97.145 71.175 97.435 ;
        RECT 71.345 97.315 71.675 97.695 ;
        RECT 71.005 96.975 71.670 97.145 ;
        RECT 39.635 95.145 44.980 95.580 ;
        RECT 45.155 95.145 50.500 95.580 ;
        RECT 50.675 95.145 56.020 95.580 ;
        RECT 56.195 95.145 61.540 95.580 ;
        RECT 61.715 95.145 64.305 96.235 ;
        RECT 64.935 95.145 65.225 96.310 ;
        RECT 68.800 95.580 69.150 96.830 ;
        RECT 70.920 96.155 71.270 96.805 ;
        RECT 71.440 95.985 71.670 96.975 ;
        RECT 71.005 95.815 71.670 95.985 ;
        RECT 65.395 95.145 70.740 95.580 ;
        RECT 71.005 95.315 71.175 95.815 ;
        RECT 71.345 95.145 71.675 95.645 ;
        RECT 71.845 95.315 72.030 97.435 ;
        RECT 72.285 97.235 72.535 97.695 ;
        RECT 72.705 97.245 73.040 97.415 ;
        RECT 73.235 97.245 73.910 97.415 ;
        RECT 72.705 97.105 72.875 97.245 ;
        RECT 72.200 96.115 72.480 97.065 ;
        RECT 72.650 96.975 72.875 97.105 ;
        RECT 72.650 95.870 72.820 96.975 ;
        RECT 73.045 96.825 73.570 97.045 ;
        RECT 72.990 96.060 73.230 96.655 ;
        RECT 73.400 96.125 73.570 96.825 ;
        RECT 73.740 96.465 73.910 97.245 ;
        RECT 74.230 97.195 74.600 97.695 ;
        RECT 74.780 97.245 75.185 97.415 ;
        RECT 75.355 97.245 76.140 97.415 ;
        RECT 74.780 97.015 74.950 97.245 ;
        RECT 74.120 96.715 74.950 97.015 ;
        RECT 75.335 96.745 75.800 97.075 ;
        RECT 74.120 96.685 74.320 96.715 ;
        RECT 74.440 96.465 74.610 96.535 ;
        RECT 73.740 96.295 74.610 96.465 ;
        RECT 74.100 96.205 74.610 96.295 ;
        RECT 72.650 95.740 72.955 95.870 ;
        RECT 73.400 95.760 73.930 96.125 ;
        RECT 72.270 95.145 72.535 95.605 ;
        RECT 72.705 95.315 72.955 95.740 ;
        RECT 74.100 95.590 74.270 96.205 ;
        RECT 73.165 95.420 74.270 95.590 ;
        RECT 74.440 95.145 74.610 95.945 ;
        RECT 74.780 95.645 74.950 96.715 ;
        RECT 75.120 95.815 75.310 96.535 ;
        RECT 75.480 95.785 75.800 96.745 ;
        RECT 75.970 96.785 76.140 97.245 ;
        RECT 76.415 97.165 76.625 97.695 ;
        RECT 76.885 96.955 77.215 97.480 ;
        RECT 77.385 97.085 77.555 97.695 ;
        RECT 77.725 97.040 78.055 97.475 ;
        RECT 77.725 96.955 78.105 97.040 ;
        RECT 77.015 96.785 77.215 96.955 ;
        RECT 77.880 96.915 78.105 96.955 ;
        RECT 75.970 96.455 76.845 96.785 ;
        RECT 77.015 96.455 77.765 96.785 ;
        RECT 74.780 95.315 75.030 95.645 ;
        RECT 75.970 95.615 76.140 96.455 ;
        RECT 77.015 96.250 77.205 96.455 ;
        RECT 77.935 96.335 78.105 96.915 ;
        RECT 78.275 96.945 79.485 97.695 ;
        RECT 78.275 96.405 78.795 96.945 ;
        RECT 79.655 96.895 79.995 97.525 ;
        RECT 80.165 96.895 80.415 97.695 ;
        RECT 80.605 97.045 80.935 97.525 ;
        RECT 81.105 97.235 81.330 97.695 ;
        RECT 81.500 97.045 81.830 97.525 ;
        RECT 77.890 96.285 78.105 96.335 ;
        RECT 76.310 95.875 77.205 96.250 ;
        RECT 77.715 96.205 78.105 96.285 ;
        RECT 78.965 96.235 79.485 96.775 ;
        RECT 75.255 95.445 76.140 95.615 ;
        RECT 76.320 95.145 76.635 95.645 ;
        RECT 76.865 95.315 77.205 95.875 ;
        RECT 77.375 95.145 77.545 96.155 ;
        RECT 77.715 95.360 78.045 96.205 ;
        RECT 78.275 95.145 79.485 96.235 ;
        RECT 79.655 96.285 79.830 96.895 ;
        RECT 80.605 96.875 81.830 97.045 ;
        RECT 82.460 96.915 82.960 97.525 ;
        RECT 80.000 96.535 80.695 96.705 ;
        RECT 80.525 96.285 80.695 96.535 ;
        RECT 80.870 96.505 81.290 96.705 ;
        RECT 81.460 96.505 81.790 96.705 ;
        RECT 81.960 96.505 82.290 96.705 ;
        RECT 82.460 96.285 82.630 96.915 ;
        RECT 83.335 96.895 83.675 97.525 ;
        RECT 83.845 96.895 84.095 97.695 ;
        RECT 84.285 97.045 84.615 97.525 ;
        RECT 84.785 97.235 85.010 97.695 ;
        RECT 85.180 97.045 85.510 97.525 ;
        RECT 82.815 96.455 83.165 96.705 ;
        RECT 83.335 96.285 83.510 96.895 ;
        RECT 84.285 96.875 85.510 97.045 ;
        RECT 86.140 96.915 86.640 97.525 ;
        RECT 87.015 97.195 87.275 97.525 ;
        RECT 87.445 97.335 87.775 97.695 ;
        RECT 88.030 97.315 89.330 97.525 ;
        RECT 83.680 96.535 84.375 96.705 ;
        RECT 84.205 96.285 84.375 96.535 ;
        RECT 84.550 96.505 84.970 96.705 ;
        RECT 85.140 96.505 85.470 96.705 ;
        RECT 85.640 96.505 85.970 96.705 ;
        RECT 86.140 96.285 86.310 96.915 ;
        RECT 86.495 96.455 86.845 96.705 ;
        RECT 79.655 95.315 79.995 96.285 ;
        RECT 80.165 95.145 80.335 96.285 ;
        RECT 80.525 96.115 82.960 96.285 ;
        RECT 80.605 95.145 80.855 95.945 ;
        RECT 81.500 95.315 81.830 96.115 ;
        RECT 82.130 95.145 82.460 95.945 ;
        RECT 82.630 95.315 82.960 96.115 ;
        RECT 83.335 95.315 83.675 96.285 ;
        RECT 83.845 95.145 84.015 96.285 ;
        RECT 84.205 96.115 86.640 96.285 ;
        RECT 84.285 95.145 84.535 95.945 ;
        RECT 85.180 95.315 85.510 96.115 ;
        RECT 85.810 95.145 86.140 95.945 ;
        RECT 86.310 95.315 86.640 96.115 ;
        RECT 87.015 95.995 87.185 97.195 ;
        RECT 88.030 97.165 88.200 97.315 ;
        RECT 87.445 97.040 88.200 97.165 ;
        RECT 87.355 96.995 88.200 97.040 ;
        RECT 87.355 96.875 87.625 96.995 ;
        RECT 87.355 96.300 87.525 96.875 ;
        RECT 87.755 96.435 88.165 96.740 ;
        RECT 88.455 96.705 88.665 97.105 ;
        RECT 88.335 96.495 88.665 96.705 ;
        RECT 88.910 96.705 89.130 97.105 ;
        RECT 89.605 96.930 90.060 97.695 ;
        RECT 90.695 96.970 90.985 97.695 ;
        RECT 91.320 97.185 91.560 97.695 ;
        RECT 91.740 97.185 92.020 97.515 ;
        RECT 92.250 97.185 92.465 97.695 ;
        RECT 88.910 96.495 89.385 96.705 ;
        RECT 89.575 96.505 90.065 96.705 ;
        RECT 91.215 96.455 91.570 97.015 ;
        RECT 87.355 96.265 87.555 96.300 ;
        RECT 88.885 96.265 90.060 96.325 ;
        RECT 87.355 96.155 90.060 96.265 ;
        RECT 87.415 96.095 89.215 96.155 ;
        RECT 88.885 96.065 89.215 96.095 ;
        RECT 87.015 95.315 87.275 95.995 ;
        RECT 87.445 95.145 87.695 95.925 ;
        RECT 87.945 95.895 88.780 95.905 ;
        RECT 89.370 95.895 89.555 95.985 ;
        RECT 87.945 95.695 89.555 95.895 ;
        RECT 87.945 95.315 88.195 95.695 ;
        RECT 89.325 95.655 89.555 95.695 ;
        RECT 89.805 95.535 90.060 96.155 ;
        RECT 88.365 95.145 88.720 95.525 ;
        RECT 89.725 95.315 90.060 95.535 ;
        RECT 90.695 95.145 90.985 96.310 ;
        RECT 91.740 96.285 91.910 97.185 ;
        RECT 92.080 96.455 92.345 97.015 ;
        RECT 92.635 96.955 93.250 97.525 ;
        RECT 92.595 96.285 92.765 96.785 ;
        RECT 91.340 96.115 92.765 96.285 ;
        RECT 91.340 95.940 91.730 96.115 ;
        RECT 92.215 95.145 92.545 95.945 ;
        RECT 92.935 95.935 93.250 96.955 ;
        RECT 93.660 96.915 94.160 97.525 ;
        RECT 93.455 96.455 93.805 96.705 ;
        RECT 93.990 96.285 94.160 96.915 ;
        RECT 94.790 97.045 95.120 97.525 ;
        RECT 95.290 97.235 95.515 97.695 ;
        RECT 95.685 97.045 96.015 97.525 ;
        RECT 94.790 96.875 96.015 97.045 ;
        RECT 96.205 96.895 96.455 97.695 ;
        RECT 96.625 96.895 96.965 97.525 ;
        RECT 94.330 96.505 94.660 96.705 ;
        RECT 94.830 96.505 95.160 96.705 ;
        RECT 95.330 96.505 95.750 96.705 ;
        RECT 95.925 96.535 96.620 96.705 ;
        RECT 95.925 96.285 96.095 96.535 ;
        RECT 96.790 96.285 96.965 96.895 ;
        RECT 97.135 96.945 98.345 97.695 ;
        RECT 98.605 97.145 98.775 97.435 ;
        RECT 98.945 97.315 99.275 97.695 ;
        RECT 98.605 96.975 99.270 97.145 ;
        RECT 97.135 96.405 97.655 96.945 ;
        RECT 92.715 95.315 93.250 95.935 ;
        RECT 93.660 96.115 96.095 96.285 ;
        RECT 93.660 95.315 93.990 96.115 ;
        RECT 94.160 95.145 94.490 95.945 ;
        RECT 94.790 95.315 95.120 96.115 ;
        RECT 95.765 95.145 96.015 95.945 ;
        RECT 96.285 95.145 96.455 96.285 ;
        RECT 96.625 95.315 96.965 96.285 ;
        RECT 97.825 96.235 98.345 96.775 ;
        RECT 97.135 95.145 98.345 96.235 ;
        RECT 98.520 96.155 98.870 96.805 ;
        RECT 99.040 95.985 99.270 96.975 ;
        RECT 98.605 95.815 99.270 95.985 ;
        RECT 98.605 95.315 98.775 95.815 ;
        RECT 98.945 95.145 99.275 95.645 ;
        RECT 99.445 95.315 99.630 97.435 ;
        RECT 99.885 97.235 100.135 97.695 ;
        RECT 100.305 97.245 100.640 97.415 ;
        RECT 100.835 97.245 101.510 97.415 ;
        RECT 100.305 97.105 100.475 97.245 ;
        RECT 99.800 96.115 100.080 97.065 ;
        RECT 100.250 96.975 100.475 97.105 ;
        RECT 100.250 95.870 100.420 96.975 ;
        RECT 100.645 96.825 101.170 97.045 ;
        RECT 100.590 96.060 100.830 96.655 ;
        RECT 101.000 96.125 101.170 96.825 ;
        RECT 101.340 96.465 101.510 97.245 ;
        RECT 101.830 97.195 102.200 97.695 ;
        RECT 102.380 97.245 102.785 97.415 ;
        RECT 102.955 97.245 103.740 97.415 ;
        RECT 102.380 97.015 102.550 97.245 ;
        RECT 101.720 96.715 102.550 97.015 ;
        RECT 102.935 96.745 103.400 97.075 ;
        RECT 101.720 96.685 101.920 96.715 ;
        RECT 102.040 96.465 102.210 96.535 ;
        RECT 101.340 96.295 102.210 96.465 ;
        RECT 101.700 96.205 102.210 96.295 ;
        RECT 100.250 95.740 100.555 95.870 ;
        RECT 101.000 95.760 101.530 96.125 ;
        RECT 99.870 95.145 100.135 95.605 ;
        RECT 100.305 95.315 100.555 95.740 ;
        RECT 101.700 95.590 101.870 96.205 ;
        RECT 100.765 95.420 101.870 95.590 ;
        RECT 102.040 95.145 102.210 95.945 ;
        RECT 102.380 95.645 102.550 96.715 ;
        RECT 102.720 95.815 102.910 96.535 ;
        RECT 103.080 95.785 103.400 96.745 ;
        RECT 103.570 96.785 103.740 97.245 ;
        RECT 104.015 97.165 104.225 97.695 ;
        RECT 104.485 96.955 104.815 97.480 ;
        RECT 104.985 97.085 105.155 97.695 ;
        RECT 105.325 97.040 105.655 97.475 ;
        RECT 105.325 96.955 105.705 97.040 ;
        RECT 104.615 96.785 104.815 96.955 ;
        RECT 105.480 96.915 105.705 96.955 ;
        RECT 103.570 96.455 104.445 96.785 ;
        RECT 104.615 96.455 105.365 96.785 ;
        RECT 102.380 95.315 102.630 95.645 ;
        RECT 103.570 95.615 103.740 96.455 ;
        RECT 104.615 96.250 104.805 96.455 ;
        RECT 105.535 96.335 105.705 96.915 ;
        RECT 105.490 96.285 105.705 96.335 ;
        RECT 103.910 95.875 104.805 96.250 ;
        RECT 105.315 96.205 105.705 96.285 ;
        RECT 105.875 96.895 106.215 97.525 ;
        RECT 106.385 96.895 106.635 97.695 ;
        RECT 106.825 97.045 107.155 97.525 ;
        RECT 107.325 97.235 107.550 97.695 ;
        RECT 107.720 97.045 108.050 97.525 ;
        RECT 105.875 96.285 106.050 96.895 ;
        RECT 106.825 96.875 108.050 97.045 ;
        RECT 108.680 96.915 109.180 97.525 ;
        RECT 109.560 96.930 110.015 97.695 ;
        RECT 110.290 97.315 111.590 97.525 ;
        RECT 111.845 97.335 112.175 97.695 ;
        RECT 111.420 97.165 111.590 97.315 ;
        RECT 112.345 97.195 112.605 97.525 ;
        RECT 106.220 96.535 106.915 96.705 ;
        RECT 106.745 96.285 106.915 96.535 ;
        RECT 107.090 96.505 107.510 96.705 ;
        RECT 107.680 96.505 108.010 96.705 ;
        RECT 108.180 96.505 108.510 96.705 ;
        RECT 108.680 96.285 108.850 96.915 ;
        RECT 110.490 96.705 110.710 97.105 ;
        RECT 109.035 96.455 109.385 96.705 ;
        RECT 109.555 96.505 110.045 96.705 ;
        RECT 110.235 96.495 110.710 96.705 ;
        RECT 110.955 96.705 111.165 97.105 ;
        RECT 111.420 97.040 112.175 97.165 ;
        RECT 111.420 96.995 112.265 97.040 ;
        RECT 111.995 96.875 112.265 96.995 ;
        RECT 110.955 96.495 111.285 96.705 ;
        RECT 111.455 96.435 111.865 96.740 ;
        RECT 102.855 95.445 103.740 95.615 ;
        RECT 103.920 95.145 104.235 95.645 ;
        RECT 104.465 95.315 104.805 95.875 ;
        RECT 104.975 95.145 105.145 96.155 ;
        RECT 105.315 95.360 105.645 96.205 ;
        RECT 105.875 95.315 106.215 96.285 ;
        RECT 106.385 95.145 106.555 96.285 ;
        RECT 106.745 96.115 109.180 96.285 ;
        RECT 106.825 95.145 107.075 95.945 ;
        RECT 107.720 95.315 108.050 96.115 ;
        RECT 108.350 95.145 108.680 95.945 ;
        RECT 108.850 95.315 109.180 96.115 ;
        RECT 109.560 96.265 110.735 96.325 ;
        RECT 112.095 96.300 112.265 96.875 ;
        RECT 112.065 96.265 112.265 96.300 ;
        RECT 109.560 96.155 112.265 96.265 ;
        RECT 109.560 95.535 109.815 96.155 ;
        RECT 110.405 96.095 112.205 96.155 ;
        RECT 110.405 96.065 110.735 96.095 ;
        RECT 112.435 95.995 112.605 97.195 ;
        RECT 112.775 96.945 113.985 97.695 ;
        RECT 114.320 97.185 114.560 97.695 ;
        RECT 114.740 97.185 115.020 97.515 ;
        RECT 115.250 97.185 115.465 97.695 ;
        RECT 112.775 96.405 113.295 96.945 ;
        RECT 113.465 96.235 113.985 96.775 ;
        RECT 114.215 96.455 114.570 97.015 ;
        RECT 114.740 96.285 114.910 97.185 ;
        RECT 115.080 96.455 115.345 97.015 ;
        RECT 115.635 96.955 116.250 97.525 ;
        RECT 116.455 96.970 116.745 97.695 ;
        RECT 115.595 96.285 115.765 96.785 ;
        RECT 110.065 95.895 110.250 95.985 ;
        RECT 110.840 95.895 111.675 95.905 ;
        RECT 110.065 95.695 111.675 95.895 ;
        RECT 110.065 95.655 110.295 95.695 ;
        RECT 109.560 95.315 109.895 95.535 ;
        RECT 110.900 95.145 111.255 95.525 ;
        RECT 111.425 95.315 111.675 95.695 ;
        RECT 111.925 95.145 112.175 95.925 ;
        RECT 112.345 95.315 112.605 95.995 ;
        RECT 112.775 95.145 113.985 96.235 ;
        RECT 114.340 96.115 115.765 96.285 ;
        RECT 114.340 95.940 114.730 96.115 ;
        RECT 115.215 95.145 115.545 95.945 ;
        RECT 115.935 95.935 116.250 96.955 ;
        RECT 117.120 96.915 117.620 97.525 ;
        RECT 116.915 96.455 117.265 96.705 ;
        RECT 115.715 95.315 116.250 95.935 ;
        RECT 116.455 95.145 116.745 96.310 ;
        RECT 117.450 96.285 117.620 96.915 ;
        RECT 118.250 97.045 118.580 97.525 ;
        RECT 118.750 97.235 118.975 97.695 ;
        RECT 119.145 97.045 119.475 97.525 ;
        RECT 118.250 96.875 119.475 97.045 ;
        RECT 119.665 96.895 119.915 97.695 ;
        RECT 120.085 96.895 120.425 97.525 ;
        RECT 117.790 96.505 118.120 96.705 ;
        RECT 118.290 96.505 118.620 96.705 ;
        RECT 118.790 96.505 119.210 96.705 ;
        RECT 119.385 96.535 120.080 96.705 ;
        RECT 119.385 96.285 119.555 96.535 ;
        RECT 120.250 96.285 120.425 96.895 ;
        RECT 117.120 96.115 119.555 96.285 ;
        RECT 117.120 95.315 117.450 96.115 ;
        RECT 117.620 95.145 117.950 95.945 ;
        RECT 118.250 95.315 118.580 96.115 ;
        RECT 119.225 95.145 119.475 95.945 ;
        RECT 119.745 95.145 119.915 96.285 ;
        RECT 120.085 95.315 120.425 96.285 ;
        RECT 121.055 96.895 121.395 97.525 ;
        RECT 121.565 96.895 121.815 97.695 ;
        RECT 122.005 97.045 122.335 97.525 ;
        RECT 122.505 97.235 122.730 97.695 ;
        RECT 122.900 97.045 123.230 97.525 ;
        RECT 121.055 96.285 121.230 96.895 ;
        RECT 122.005 96.875 123.230 97.045 ;
        RECT 123.860 96.915 124.360 97.525 ;
        RECT 125.245 97.040 125.575 97.475 ;
        RECT 125.745 97.085 125.915 97.695 ;
        RECT 125.195 96.955 125.575 97.040 ;
        RECT 126.085 96.955 126.415 97.480 ;
        RECT 126.675 97.165 126.885 97.695 ;
        RECT 127.160 97.245 127.945 97.415 ;
        RECT 128.115 97.245 128.520 97.415 ;
        RECT 125.195 96.915 125.420 96.955 ;
        RECT 121.400 96.535 122.095 96.705 ;
        RECT 121.925 96.285 122.095 96.535 ;
        RECT 122.270 96.505 122.690 96.705 ;
        RECT 122.860 96.505 123.190 96.705 ;
        RECT 123.360 96.505 123.690 96.705 ;
        RECT 123.860 96.285 124.030 96.915 ;
        RECT 124.215 96.455 124.565 96.705 ;
        RECT 125.195 96.335 125.365 96.915 ;
        RECT 126.085 96.785 126.285 96.955 ;
        RECT 127.160 96.785 127.330 97.245 ;
        RECT 125.535 96.455 126.285 96.785 ;
        RECT 126.455 96.455 127.330 96.785 ;
        RECT 125.195 96.285 125.410 96.335 ;
        RECT 121.055 95.315 121.395 96.285 ;
        RECT 121.565 95.145 121.735 96.285 ;
        RECT 121.925 96.115 124.360 96.285 ;
        RECT 125.195 96.205 125.585 96.285 ;
        RECT 122.005 95.145 122.255 95.945 ;
        RECT 122.900 95.315 123.230 96.115 ;
        RECT 123.530 95.145 123.860 95.945 ;
        RECT 124.030 95.315 124.360 96.115 ;
        RECT 125.255 95.360 125.585 96.205 ;
        RECT 126.095 96.250 126.285 96.455 ;
        RECT 125.755 95.145 125.925 96.155 ;
        RECT 126.095 95.875 126.990 96.250 ;
        RECT 126.095 95.315 126.435 95.875 ;
        RECT 126.665 95.145 126.980 95.645 ;
        RECT 127.160 95.615 127.330 96.455 ;
        RECT 127.500 96.745 127.965 97.075 ;
        RECT 128.350 97.015 128.520 97.245 ;
        RECT 128.700 97.195 129.070 97.695 ;
        RECT 129.390 97.245 130.065 97.415 ;
        RECT 130.260 97.245 130.595 97.415 ;
        RECT 127.500 95.785 127.820 96.745 ;
        RECT 128.350 96.715 129.180 97.015 ;
        RECT 127.990 95.815 128.180 96.535 ;
        RECT 128.350 95.645 128.520 96.715 ;
        RECT 128.980 96.685 129.180 96.715 ;
        RECT 128.690 96.465 128.860 96.535 ;
        RECT 129.390 96.465 129.560 97.245 ;
        RECT 130.425 97.105 130.595 97.245 ;
        RECT 130.765 97.235 131.015 97.695 ;
        RECT 128.690 96.295 129.560 96.465 ;
        RECT 129.730 96.825 130.255 97.045 ;
        RECT 130.425 96.975 130.650 97.105 ;
        RECT 128.690 96.205 129.200 96.295 ;
        RECT 127.160 95.445 128.045 95.615 ;
        RECT 128.270 95.315 128.520 95.645 ;
        RECT 128.690 95.145 128.860 95.945 ;
        RECT 129.030 95.590 129.200 96.205 ;
        RECT 129.730 96.125 129.900 96.825 ;
        RECT 129.370 95.760 129.900 96.125 ;
        RECT 130.070 96.060 130.310 96.655 ;
        RECT 130.480 95.870 130.650 96.975 ;
        RECT 130.820 96.115 131.100 97.065 ;
        RECT 130.345 95.740 130.650 95.870 ;
        RECT 129.030 95.420 130.135 95.590 ;
        RECT 130.345 95.315 130.595 95.740 ;
        RECT 130.765 95.145 131.030 95.605 ;
        RECT 131.270 95.315 131.455 97.435 ;
        RECT 131.625 97.315 131.955 97.695 ;
        RECT 132.125 97.145 132.295 97.435 ;
        RECT 131.630 96.975 132.295 97.145 ;
        RECT 131.630 95.985 131.860 96.975 ;
        RECT 132.555 96.945 133.765 97.695 ;
        RECT 134.025 97.145 134.195 97.525 ;
        RECT 134.410 97.315 134.740 97.695 ;
        RECT 134.025 96.975 134.740 97.145 ;
        RECT 132.030 96.155 132.380 96.805 ;
        RECT 132.555 96.405 133.075 96.945 ;
        RECT 133.245 96.235 133.765 96.775 ;
        RECT 133.935 96.425 134.290 96.795 ;
        RECT 134.570 96.785 134.740 96.975 ;
        RECT 134.910 96.950 135.165 97.525 ;
        RECT 134.570 96.455 134.825 96.785 ;
        RECT 134.570 96.245 134.740 96.455 ;
        RECT 131.630 95.815 132.295 95.985 ;
        RECT 131.625 95.145 131.955 95.645 ;
        RECT 132.125 95.315 132.295 95.815 ;
        RECT 132.555 95.145 133.765 96.235 ;
        RECT 134.025 96.075 134.740 96.245 ;
        RECT 134.995 96.220 135.165 96.950 ;
        RECT 135.340 96.855 135.600 97.695 ;
        RECT 135.865 97.145 136.035 97.525 ;
        RECT 136.250 97.315 136.580 97.695 ;
        RECT 135.865 96.975 136.580 97.145 ;
        RECT 135.775 96.425 136.130 96.795 ;
        RECT 136.410 96.785 136.580 96.975 ;
        RECT 136.750 96.950 137.005 97.525 ;
        RECT 136.410 96.455 136.665 96.785 ;
        RECT 134.025 95.315 134.195 96.075 ;
        RECT 134.410 95.145 134.740 95.905 ;
        RECT 134.910 95.315 135.165 96.220 ;
        RECT 135.340 95.145 135.600 96.295 ;
        RECT 136.410 96.245 136.580 96.455 ;
        RECT 135.865 96.075 136.580 96.245 ;
        RECT 136.835 96.220 137.005 96.950 ;
        RECT 137.180 96.855 137.440 97.695 ;
        RECT 137.615 96.945 138.825 97.695 ;
        RECT 135.865 95.315 136.035 96.075 ;
        RECT 136.250 95.145 136.580 95.905 ;
        RECT 136.750 95.315 137.005 96.220 ;
        RECT 137.180 95.145 137.440 96.295 ;
        RECT 137.615 96.235 138.135 96.775 ;
        RECT 138.305 96.405 138.825 96.945 ;
        RECT 137.615 95.145 138.825 96.235 ;
        RECT 13.330 94.975 138.910 95.145 ;
        RECT 13.415 93.885 14.625 94.975 ;
        RECT 14.795 94.540 20.140 94.975 ;
        RECT 20.315 94.540 25.660 94.975 ;
        RECT 13.415 93.175 13.935 93.715 ;
        RECT 14.105 93.345 14.625 93.885 ;
        RECT 13.415 92.425 14.625 93.175 ;
        RECT 16.380 92.970 16.720 93.800 ;
        RECT 18.200 93.290 18.550 94.540 ;
        RECT 21.900 92.970 22.240 93.800 ;
        RECT 23.720 93.290 24.070 94.540 ;
        RECT 26.295 93.810 26.585 94.975 ;
        RECT 26.755 94.540 32.100 94.975 ;
        RECT 32.275 94.540 37.620 94.975 ;
        RECT 37.795 94.540 43.140 94.975 ;
        RECT 43.315 94.540 48.660 94.975 ;
        RECT 14.795 92.425 20.140 92.970 ;
        RECT 20.315 92.425 25.660 92.970 ;
        RECT 26.295 92.425 26.585 93.150 ;
        RECT 28.340 92.970 28.680 93.800 ;
        RECT 30.160 93.290 30.510 94.540 ;
        RECT 33.860 92.970 34.200 93.800 ;
        RECT 35.680 93.290 36.030 94.540 ;
        RECT 39.380 92.970 39.720 93.800 ;
        RECT 41.200 93.290 41.550 94.540 ;
        RECT 44.900 92.970 45.240 93.800 ;
        RECT 46.720 93.290 47.070 94.540 ;
        RECT 48.835 93.885 51.425 94.975 ;
        RECT 48.835 93.195 50.045 93.715 ;
        RECT 50.215 93.365 51.425 93.885 ;
        RECT 52.055 93.810 52.345 94.975 ;
        RECT 52.515 94.540 57.860 94.975 ;
        RECT 58.035 94.540 63.380 94.975 ;
        RECT 63.555 94.540 68.900 94.975 ;
        RECT 69.075 94.540 74.420 94.975 ;
        RECT 26.755 92.425 32.100 92.970 ;
        RECT 32.275 92.425 37.620 92.970 ;
        RECT 37.795 92.425 43.140 92.970 ;
        RECT 43.315 92.425 48.660 92.970 ;
        RECT 48.835 92.425 51.425 93.195 ;
        RECT 52.055 92.425 52.345 93.150 ;
        RECT 54.100 92.970 54.440 93.800 ;
        RECT 55.920 93.290 56.270 94.540 ;
        RECT 59.620 92.970 59.960 93.800 ;
        RECT 61.440 93.290 61.790 94.540 ;
        RECT 65.140 92.970 65.480 93.800 ;
        RECT 66.960 93.290 67.310 94.540 ;
        RECT 70.660 92.970 71.000 93.800 ;
        RECT 72.480 93.290 72.830 94.540 ;
        RECT 74.595 93.885 77.185 94.975 ;
        RECT 74.595 93.195 75.805 93.715 ;
        RECT 75.975 93.365 77.185 93.885 ;
        RECT 77.815 93.810 78.105 94.975 ;
        RECT 78.365 94.305 78.535 94.805 ;
        RECT 78.705 94.475 79.035 94.975 ;
        RECT 78.365 94.135 79.030 94.305 ;
        RECT 78.280 93.315 78.630 93.965 ;
        RECT 52.515 92.425 57.860 92.970 ;
        RECT 58.035 92.425 63.380 92.970 ;
        RECT 63.555 92.425 68.900 92.970 ;
        RECT 69.075 92.425 74.420 92.970 ;
        RECT 74.595 92.425 77.185 93.195 ;
        RECT 77.815 92.425 78.105 93.150 ;
        RECT 78.800 93.145 79.030 94.135 ;
        RECT 78.365 92.975 79.030 93.145 ;
        RECT 78.365 92.685 78.535 92.975 ;
        RECT 78.705 92.425 79.035 92.805 ;
        RECT 79.205 92.685 79.390 94.805 ;
        RECT 79.630 94.515 79.895 94.975 ;
        RECT 80.065 94.380 80.315 94.805 ;
        RECT 80.525 94.530 81.630 94.700 ;
        RECT 80.010 94.250 80.315 94.380 ;
        RECT 79.560 93.055 79.840 94.005 ;
        RECT 80.010 93.145 80.180 94.250 ;
        RECT 80.350 93.465 80.590 94.060 ;
        RECT 80.760 93.995 81.290 94.360 ;
        RECT 80.760 93.295 80.930 93.995 ;
        RECT 81.460 93.915 81.630 94.530 ;
        RECT 81.800 94.175 81.970 94.975 ;
        RECT 82.140 94.475 82.390 94.805 ;
        RECT 82.615 94.505 83.500 94.675 ;
        RECT 81.460 93.825 81.970 93.915 ;
        RECT 80.010 93.015 80.235 93.145 ;
        RECT 80.405 93.075 80.930 93.295 ;
        RECT 81.100 93.655 81.970 93.825 ;
        RECT 79.645 92.425 79.895 92.885 ;
        RECT 80.065 92.875 80.235 93.015 ;
        RECT 81.100 92.875 81.270 93.655 ;
        RECT 81.800 93.585 81.970 93.655 ;
        RECT 81.480 93.405 81.680 93.435 ;
        RECT 82.140 93.405 82.310 94.475 ;
        RECT 82.480 93.585 82.670 94.305 ;
        RECT 81.480 93.105 82.310 93.405 ;
        RECT 82.840 93.375 83.160 94.335 ;
        RECT 80.065 92.705 80.400 92.875 ;
        RECT 80.595 92.705 81.270 92.875 ;
        RECT 81.590 92.425 81.960 92.925 ;
        RECT 82.140 92.875 82.310 93.105 ;
        RECT 82.695 93.045 83.160 93.375 ;
        RECT 83.330 93.665 83.500 94.505 ;
        RECT 83.680 94.475 83.995 94.975 ;
        RECT 84.225 94.245 84.565 94.805 ;
        RECT 83.670 93.870 84.565 94.245 ;
        RECT 84.735 93.965 84.905 94.975 ;
        RECT 84.375 93.665 84.565 93.870 ;
        RECT 85.075 93.915 85.405 94.760 ;
        RECT 85.075 93.835 85.465 93.915 ;
        RECT 85.635 93.885 86.845 94.975 ;
        RECT 87.105 94.305 87.275 94.805 ;
        RECT 87.445 94.475 87.775 94.975 ;
        RECT 87.105 94.135 87.770 94.305 ;
        RECT 85.250 93.785 85.465 93.835 ;
        RECT 83.330 93.335 84.205 93.665 ;
        RECT 84.375 93.335 85.125 93.665 ;
        RECT 83.330 92.875 83.500 93.335 ;
        RECT 84.375 93.165 84.575 93.335 ;
        RECT 85.295 93.205 85.465 93.785 ;
        RECT 85.240 93.165 85.465 93.205 ;
        RECT 82.140 92.705 82.545 92.875 ;
        RECT 82.715 92.705 83.500 92.875 ;
        RECT 83.775 92.425 83.985 92.955 ;
        RECT 84.245 92.640 84.575 93.165 ;
        RECT 85.085 93.080 85.465 93.165 ;
        RECT 85.635 93.175 86.155 93.715 ;
        RECT 86.325 93.345 86.845 93.885 ;
        RECT 87.020 93.315 87.370 93.965 ;
        RECT 84.745 92.425 84.915 93.035 ;
        RECT 85.085 92.645 85.415 93.080 ;
        RECT 85.635 92.425 86.845 93.175 ;
        RECT 87.540 93.145 87.770 94.135 ;
        RECT 87.105 92.975 87.770 93.145 ;
        RECT 87.105 92.685 87.275 92.975 ;
        RECT 87.445 92.425 87.775 92.805 ;
        RECT 87.945 92.685 88.130 94.805 ;
        RECT 88.370 94.515 88.635 94.975 ;
        RECT 88.805 94.380 89.055 94.805 ;
        RECT 89.265 94.530 90.370 94.700 ;
        RECT 88.750 94.250 89.055 94.380 ;
        RECT 88.300 93.055 88.580 94.005 ;
        RECT 88.750 93.145 88.920 94.250 ;
        RECT 89.090 93.465 89.330 94.060 ;
        RECT 89.500 93.995 90.030 94.360 ;
        RECT 89.500 93.295 89.670 93.995 ;
        RECT 90.200 93.915 90.370 94.530 ;
        RECT 90.540 94.175 90.710 94.975 ;
        RECT 90.880 94.475 91.130 94.805 ;
        RECT 91.355 94.505 92.240 94.675 ;
        RECT 90.200 93.825 90.710 93.915 ;
        RECT 88.750 93.015 88.975 93.145 ;
        RECT 89.145 93.075 89.670 93.295 ;
        RECT 89.840 93.655 90.710 93.825 ;
        RECT 88.385 92.425 88.635 92.885 ;
        RECT 88.805 92.875 88.975 93.015 ;
        RECT 89.840 92.875 90.010 93.655 ;
        RECT 90.540 93.585 90.710 93.655 ;
        RECT 90.220 93.405 90.420 93.435 ;
        RECT 90.880 93.405 91.050 94.475 ;
        RECT 91.220 93.585 91.410 94.305 ;
        RECT 90.220 93.105 91.050 93.405 ;
        RECT 91.580 93.375 91.900 94.335 ;
        RECT 88.805 92.705 89.140 92.875 ;
        RECT 89.335 92.705 90.010 92.875 ;
        RECT 90.330 92.425 90.700 92.925 ;
        RECT 90.880 92.875 91.050 93.105 ;
        RECT 91.435 93.045 91.900 93.375 ;
        RECT 92.070 93.665 92.240 94.505 ;
        RECT 92.420 94.475 92.735 94.975 ;
        RECT 92.965 94.245 93.305 94.805 ;
        RECT 92.410 93.870 93.305 94.245 ;
        RECT 93.475 93.965 93.645 94.975 ;
        RECT 93.115 93.665 93.305 93.870 ;
        RECT 93.815 93.915 94.145 94.760 ;
        RECT 94.465 94.305 94.635 94.805 ;
        RECT 94.805 94.475 95.135 94.975 ;
        RECT 94.465 94.135 95.130 94.305 ;
        RECT 93.815 93.835 94.205 93.915 ;
        RECT 93.990 93.785 94.205 93.835 ;
        RECT 92.070 93.335 92.945 93.665 ;
        RECT 93.115 93.335 93.865 93.665 ;
        RECT 92.070 92.875 92.240 93.335 ;
        RECT 93.115 93.165 93.315 93.335 ;
        RECT 94.035 93.205 94.205 93.785 ;
        RECT 94.380 93.315 94.730 93.965 ;
        RECT 93.980 93.165 94.205 93.205 ;
        RECT 90.880 92.705 91.285 92.875 ;
        RECT 91.455 92.705 92.240 92.875 ;
        RECT 92.515 92.425 92.725 92.955 ;
        RECT 92.985 92.640 93.315 93.165 ;
        RECT 93.825 93.080 94.205 93.165 ;
        RECT 94.900 93.145 95.130 94.135 ;
        RECT 93.485 92.425 93.655 93.035 ;
        RECT 93.825 92.645 94.155 93.080 ;
        RECT 94.465 92.975 95.130 93.145 ;
        RECT 94.465 92.685 94.635 92.975 ;
        RECT 94.805 92.425 95.135 92.805 ;
        RECT 95.305 92.685 95.490 94.805 ;
        RECT 95.730 94.515 95.995 94.975 ;
        RECT 96.165 94.380 96.415 94.805 ;
        RECT 96.625 94.530 97.730 94.700 ;
        RECT 96.110 94.250 96.415 94.380 ;
        RECT 95.660 93.055 95.940 94.005 ;
        RECT 96.110 93.145 96.280 94.250 ;
        RECT 96.450 93.465 96.690 94.060 ;
        RECT 96.860 93.995 97.390 94.360 ;
        RECT 96.860 93.295 97.030 93.995 ;
        RECT 97.560 93.915 97.730 94.530 ;
        RECT 97.900 94.175 98.070 94.975 ;
        RECT 98.240 94.475 98.490 94.805 ;
        RECT 98.715 94.505 99.600 94.675 ;
        RECT 97.560 93.825 98.070 93.915 ;
        RECT 96.110 93.015 96.335 93.145 ;
        RECT 96.505 93.075 97.030 93.295 ;
        RECT 97.200 93.655 98.070 93.825 ;
        RECT 95.745 92.425 95.995 92.885 ;
        RECT 96.165 92.875 96.335 93.015 ;
        RECT 97.200 92.875 97.370 93.655 ;
        RECT 97.900 93.585 98.070 93.655 ;
        RECT 97.580 93.405 97.780 93.435 ;
        RECT 98.240 93.405 98.410 94.475 ;
        RECT 98.580 93.585 98.770 94.305 ;
        RECT 97.580 93.105 98.410 93.405 ;
        RECT 98.940 93.375 99.260 94.335 ;
        RECT 96.165 92.705 96.500 92.875 ;
        RECT 96.695 92.705 97.370 92.875 ;
        RECT 97.690 92.425 98.060 92.925 ;
        RECT 98.240 92.875 98.410 93.105 ;
        RECT 98.795 93.045 99.260 93.375 ;
        RECT 99.430 93.665 99.600 94.505 ;
        RECT 99.780 94.475 100.095 94.975 ;
        RECT 100.325 94.245 100.665 94.805 ;
        RECT 99.770 93.870 100.665 94.245 ;
        RECT 100.835 93.965 101.005 94.975 ;
        RECT 100.475 93.665 100.665 93.870 ;
        RECT 101.175 93.915 101.505 94.760 ;
        RECT 101.735 94.005 102.005 94.775 ;
        RECT 102.175 94.195 102.505 94.975 ;
        RECT 102.710 94.370 102.895 94.775 ;
        RECT 103.065 94.550 103.400 94.975 ;
        RECT 102.710 94.195 103.375 94.370 ;
        RECT 101.175 93.835 101.565 93.915 ;
        RECT 101.350 93.785 101.565 93.835 ;
        RECT 99.430 93.335 100.305 93.665 ;
        RECT 100.475 93.335 101.225 93.665 ;
        RECT 99.430 92.875 99.600 93.335 ;
        RECT 100.475 93.165 100.675 93.335 ;
        RECT 101.395 93.205 101.565 93.785 ;
        RECT 101.340 93.165 101.565 93.205 ;
        RECT 98.240 92.705 98.645 92.875 ;
        RECT 98.815 92.705 99.600 92.875 ;
        RECT 99.875 92.425 100.085 92.955 ;
        RECT 100.345 92.640 100.675 93.165 ;
        RECT 101.185 93.080 101.565 93.165 ;
        RECT 101.735 93.835 102.865 94.005 ;
        RECT 100.845 92.425 101.015 93.035 ;
        RECT 101.185 92.645 101.515 93.080 ;
        RECT 101.735 92.925 101.905 93.835 ;
        RECT 102.075 93.085 102.435 93.665 ;
        RECT 102.615 93.335 102.865 93.835 ;
        RECT 103.035 93.165 103.375 94.195 ;
        RECT 103.575 93.810 103.865 94.975 ;
        RECT 104.035 93.835 104.375 94.805 ;
        RECT 104.545 93.835 104.715 94.975 ;
        RECT 104.985 94.175 105.235 94.975 ;
        RECT 105.880 94.005 106.210 94.805 ;
        RECT 106.510 94.175 106.840 94.975 ;
        RECT 107.010 94.005 107.340 94.805 ;
        RECT 104.905 93.835 107.340 94.005 ;
        RECT 107.720 94.585 108.055 94.805 ;
        RECT 109.060 94.595 109.415 94.975 ;
        RECT 107.720 93.965 107.975 94.585 ;
        RECT 108.225 94.425 108.455 94.465 ;
        RECT 109.585 94.425 109.835 94.805 ;
        RECT 108.225 94.225 109.835 94.425 ;
        RECT 108.225 94.135 108.410 94.225 ;
        RECT 109.000 94.215 109.835 94.225 ;
        RECT 110.085 94.195 110.335 94.975 ;
        RECT 110.505 94.125 110.765 94.805 ;
        RECT 108.565 94.025 108.895 94.055 ;
        RECT 108.565 93.965 110.365 94.025 ;
        RECT 107.720 93.855 110.425 93.965 ;
        RECT 102.690 92.995 103.375 93.165 ;
        RECT 104.035 93.225 104.210 93.835 ;
        RECT 104.905 93.585 105.075 93.835 ;
        RECT 104.380 93.415 105.075 93.585 ;
        RECT 105.250 93.415 105.670 93.615 ;
        RECT 105.840 93.415 106.170 93.615 ;
        RECT 106.340 93.415 106.670 93.615 ;
        RECT 101.735 92.595 101.995 92.925 ;
        RECT 102.205 92.425 102.480 92.905 ;
        RECT 102.690 92.595 102.895 92.995 ;
        RECT 103.065 92.425 103.400 92.825 ;
        RECT 103.575 92.425 103.865 93.150 ;
        RECT 104.035 92.595 104.375 93.225 ;
        RECT 104.545 92.425 104.795 93.225 ;
        RECT 104.985 93.075 106.210 93.245 ;
        RECT 104.985 92.595 105.315 93.075 ;
        RECT 105.485 92.425 105.710 92.885 ;
        RECT 105.880 92.595 106.210 93.075 ;
        RECT 106.840 93.205 107.010 93.835 ;
        RECT 107.720 93.795 108.895 93.855 ;
        RECT 110.225 93.820 110.425 93.855 ;
        RECT 107.195 93.415 107.545 93.665 ;
        RECT 107.715 93.415 108.205 93.615 ;
        RECT 108.395 93.415 108.870 93.625 ;
        RECT 106.840 92.595 107.340 93.205 ;
        RECT 107.720 92.425 108.175 93.190 ;
        RECT 108.650 93.015 108.870 93.415 ;
        RECT 109.115 93.415 109.445 93.625 ;
        RECT 109.115 93.015 109.325 93.415 ;
        RECT 109.615 93.380 110.025 93.685 ;
        RECT 110.255 93.245 110.425 93.820 ;
        RECT 110.155 93.125 110.425 93.245 ;
        RECT 109.580 93.080 110.425 93.125 ;
        RECT 109.580 92.955 110.335 93.080 ;
        RECT 109.580 92.805 109.750 92.955 ;
        RECT 110.595 92.935 110.765 94.125 ;
        RECT 111.455 93.915 111.785 94.760 ;
        RECT 111.955 93.965 112.125 94.975 ;
        RECT 112.295 94.245 112.635 94.805 ;
        RECT 112.865 94.475 113.180 94.975 ;
        RECT 113.360 94.505 114.245 94.675 ;
        RECT 111.395 93.835 111.785 93.915 ;
        RECT 112.295 93.870 113.190 94.245 ;
        RECT 111.395 93.785 111.610 93.835 ;
        RECT 111.395 93.205 111.565 93.785 ;
        RECT 112.295 93.665 112.485 93.870 ;
        RECT 113.360 93.665 113.530 94.505 ;
        RECT 114.470 94.475 114.720 94.805 ;
        RECT 111.735 93.335 112.485 93.665 ;
        RECT 112.655 93.335 113.530 93.665 ;
        RECT 111.395 93.165 111.620 93.205 ;
        RECT 112.285 93.165 112.485 93.335 ;
        RECT 111.395 93.080 111.775 93.165 ;
        RECT 110.535 92.925 110.765 92.935 ;
        RECT 108.450 92.595 109.750 92.805 ;
        RECT 110.005 92.425 110.335 92.785 ;
        RECT 110.505 92.595 110.765 92.925 ;
        RECT 111.445 92.645 111.775 93.080 ;
        RECT 111.945 92.425 112.115 93.035 ;
        RECT 112.285 92.640 112.615 93.165 ;
        RECT 112.875 92.425 113.085 92.955 ;
        RECT 113.360 92.875 113.530 93.335 ;
        RECT 113.700 93.375 114.020 94.335 ;
        RECT 114.190 93.585 114.380 94.305 ;
        RECT 114.550 93.405 114.720 94.475 ;
        RECT 114.890 94.175 115.060 94.975 ;
        RECT 115.230 94.530 116.335 94.700 ;
        RECT 115.230 93.915 115.400 94.530 ;
        RECT 116.545 94.380 116.795 94.805 ;
        RECT 116.965 94.515 117.230 94.975 ;
        RECT 115.570 93.995 116.100 94.360 ;
        RECT 116.545 94.250 116.850 94.380 ;
        RECT 114.890 93.825 115.400 93.915 ;
        RECT 114.890 93.655 115.760 93.825 ;
        RECT 114.890 93.585 115.060 93.655 ;
        RECT 115.180 93.405 115.380 93.435 ;
        RECT 113.700 93.045 114.165 93.375 ;
        RECT 114.550 93.105 115.380 93.405 ;
        RECT 114.550 92.875 114.720 93.105 ;
        RECT 113.360 92.705 114.145 92.875 ;
        RECT 114.315 92.705 114.720 92.875 ;
        RECT 114.900 92.425 115.270 92.925 ;
        RECT 115.590 92.875 115.760 93.655 ;
        RECT 115.930 93.295 116.100 93.995 ;
        RECT 116.270 93.465 116.510 94.060 ;
        RECT 115.930 93.075 116.455 93.295 ;
        RECT 116.680 93.145 116.850 94.250 ;
        RECT 116.625 93.015 116.850 93.145 ;
        RECT 117.020 93.055 117.300 94.005 ;
        RECT 116.625 92.875 116.795 93.015 ;
        RECT 115.590 92.705 116.265 92.875 ;
        RECT 116.460 92.705 116.795 92.875 ;
        RECT 116.965 92.425 117.215 92.885 ;
        RECT 117.470 92.685 117.655 94.805 ;
        RECT 117.825 94.475 118.155 94.975 ;
        RECT 118.325 94.305 118.495 94.805 ;
        RECT 117.830 94.135 118.495 94.305 ;
        RECT 118.845 94.305 119.015 94.805 ;
        RECT 119.185 94.475 119.515 94.975 ;
        RECT 118.845 94.135 119.510 94.305 ;
        RECT 117.830 93.145 118.060 94.135 ;
        RECT 118.230 93.315 118.580 93.965 ;
        RECT 118.760 93.315 119.110 93.965 ;
        RECT 119.280 93.145 119.510 94.135 ;
        RECT 117.830 92.975 118.495 93.145 ;
        RECT 117.825 92.425 118.155 92.805 ;
        RECT 118.325 92.685 118.495 92.975 ;
        RECT 118.845 92.975 119.510 93.145 ;
        RECT 118.845 92.685 119.015 92.975 ;
        RECT 119.185 92.425 119.515 92.805 ;
        RECT 119.685 92.685 119.870 94.805 ;
        RECT 120.110 94.515 120.375 94.975 ;
        RECT 120.545 94.380 120.795 94.805 ;
        RECT 121.005 94.530 122.110 94.700 ;
        RECT 120.490 94.250 120.795 94.380 ;
        RECT 120.040 93.055 120.320 94.005 ;
        RECT 120.490 93.145 120.660 94.250 ;
        RECT 120.830 93.465 121.070 94.060 ;
        RECT 121.240 93.995 121.770 94.360 ;
        RECT 121.240 93.295 121.410 93.995 ;
        RECT 121.940 93.915 122.110 94.530 ;
        RECT 122.280 94.175 122.450 94.975 ;
        RECT 122.620 94.475 122.870 94.805 ;
        RECT 123.095 94.505 123.980 94.675 ;
        RECT 121.940 93.825 122.450 93.915 ;
        RECT 120.490 93.015 120.715 93.145 ;
        RECT 120.885 93.075 121.410 93.295 ;
        RECT 121.580 93.655 122.450 93.825 ;
        RECT 120.125 92.425 120.375 92.885 ;
        RECT 120.545 92.875 120.715 93.015 ;
        RECT 121.580 92.875 121.750 93.655 ;
        RECT 122.280 93.585 122.450 93.655 ;
        RECT 121.960 93.405 122.160 93.435 ;
        RECT 122.620 93.405 122.790 94.475 ;
        RECT 122.960 93.585 123.150 94.305 ;
        RECT 121.960 93.105 122.790 93.405 ;
        RECT 123.320 93.375 123.640 94.335 ;
        RECT 120.545 92.705 120.880 92.875 ;
        RECT 121.075 92.705 121.750 92.875 ;
        RECT 122.070 92.425 122.440 92.925 ;
        RECT 122.620 92.875 122.790 93.105 ;
        RECT 123.175 93.045 123.640 93.375 ;
        RECT 123.810 93.665 123.980 94.505 ;
        RECT 124.160 94.475 124.475 94.975 ;
        RECT 124.705 94.245 125.045 94.805 ;
        RECT 124.150 93.870 125.045 94.245 ;
        RECT 125.215 93.965 125.385 94.975 ;
        RECT 124.855 93.665 125.045 93.870 ;
        RECT 125.555 93.915 125.885 94.760 ;
        RECT 126.150 94.185 126.685 94.805 ;
        RECT 125.555 93.835 125.945 93.915 ;
        RECT 125.730 93.785 125.945 93.835 ;
        RECT 123.810 93.335 124.685 93.665 ;
        RECT 124.855 93.335 125.605 93.665 ;
        RECT 123.810 92.875 123.980 93.335 ;
        RECT 124.855 93.165 125.055 93.335 ;
        RECT 125.775 93.205 125.945 93.785 ;
        RECT 125.720 93.165 125.945 93.205 ;
        RECT 122.620 92.705 123.025 92.875 ;
        RECT 123.195 92.705 123.980 92.875 ;
        RECT 124.255 92.425 124.465 92.955 ;
        RECT 124.725 92.640 125.055 93.165 ;
        RECT 125.565 93.080 125.945 93.165 ;
        RECT 126.150 93.165 126.465 94.185 ;
        RECT 126.855 94.175 127.185 94.975 ;
        RECT 127.670 94.005 128.060 94.180 ;
        RECT 126.635 93.835 128.060 94.005 ;
        RECT 126.635 93.335 126.805 93.835 ;
        RECT 125.225 92.425 125.395 93.035 ;
        RECT 125.565 92.645 125.895 93.080 ;
        RECT 126.150 92.595 126.765 93.165 ;
        RECT 127.055 93.105 127.320 93.665 ;
        RECT 127.490 92.935 127.660 93.835 ;
        RECT 129.335 93.810 129.625 94.975 ;
        RECT 130.000 94.005 130.330 94.805 ;
        RECT 130.500 94.175 130.830 94.975 ;
        RECT 131.130 94.005 131.460 94.805 ;
        RECT 132.105 94.175 132.355 94.975 ;
        RECT 130.000 93.835 132.435 94.005 ;
        RECT 132.625 93.835 132.795 94.975 ;
        RECT 132.965 93.835 133.305 94.805 ;
        RECT 133.475 93.885 135.145 94.975 ;
        RECT 127.830 93.105 128.185 93.665 ;
        RECT 129.795 93.415 130.145 93.665 ;
        RECT 130.330 93.205 130.500 93.835 ;
        RECT 130.670 93.415 131.000 93.615 ;
        RECT 131.170 93.415 131.500 93.615 ;
        RECT 131.670 93.415 132.090 93.615 ;
        RECT 132.265 93.585 132.435 93.835 ;
        RECT 132.265 93.415 132.960 93.585 ;
        RECT 126.935 92.425 127.150 92.935 ;
        RECT 127.380 92.605 127.660 92.935 ;
        RECT 127.840 92.425 128.080 92.935 ;
        RECT 129.335 92.425 129.625 93.150 ;
        RECT 130.000 92.595 130.500 93.205 ;
        RECT 131.130 93.075 132.355 93.245 ;
        RECT 133.130 93.225 133.305 93.835 ;
        RECT 131.130 92.595 131.460 93.075 ;
        RECT 131.630 92.425 131.855 92.885 ;
        RECT 132.025 92.595 132.355 93.075 ;
        RECT 132.545 92.425 132.795 93.225 ;
        RECT 132.965 92.595 133.305 93.225 ;
        RECT 133.475 93.195 134.225 93.715 ;
        RECT 134.395 93.365 135.145 93.885 ;
        RECT 135.865 94.045 136.035 94.805 ;
        RECT 136.250 94.215 136.580 94.975 ;
        RECT 135.865 93.875 136.580 94.045 ;
        RECT 136.750 93.900 137.005 94.805 ;
        RECT 135.775 93.325 136.130 93.695 ;
        RECT 136.410 93.665 136.580 93.875 ;
        RECT 136.410 93.335 136.665 93.665 ;
        RECT 133.475 92.425 135.145 93.195 ;
        RECT 136.410 93.145 136.580 93.335 ;
        RECT 136.835 93.170 137.005 93.900 ;
        RECT 137.180 93.825 137.440 94.975 ;
        RECT 137.615 93.885 138.825 94.975 ;
        RECT 137.615 93.345 138.135 93.885 ;
        RECT 135.865 92.975 136.580 93.145 ;
        RECT 135.865 92.595 136.035 92.975 ;
        RECT 136.250 92.425 136.580 92.805 ;
        RECT 136.750 92.595 137.005 93.170 ;
        RECT 137.180 92.425 137.440 93.265 ;
        RECT 138.305 93.175 138.825 93.715 ;
        RECT 137.615 92.425 138.825 93.175 ;
        RECT 13.330 92.255 138.910 92.425 ;
        RECT 13.415 91.505 14.625 92.255 ;
        RECT 14.795 91.710 20.140 92.255 ;
        RECT 20.315 91.710 25.660 92.255 ;
        RECT 25.835 91.710 31.180 92.255 ;
        RECT 31.355 91.710 36.700 92.255 ;
        RECT 13.415 90.965 13.935 91.505 ;
        RECT 14.105 90.795 14.625 91.335 ;
        RECT 16.380 90.880 16.720 91.710 ;
        RECT 13.415 89.705 14.625 90.795 ;
        RECT 18.200 90.140 18.550 91.390 ;
        RECT 21.900 90.880 22.240 91.710 ;
        RECT 23.720 90.140 24.070 91.390 ;
        RECT 27.420 90.880 27.760 91.710 ;
        RECT 29.240 90.140 29.590 91.390 ;
        RECT 32.940 90.880 33.280 91.710 ;
        RECT 36.875 91.485 38.545 92.255 ;
        RECT 39.175 91.530 39.465 92.255 ;
        RECT 39.635 91.710 44.980 92.255 ;
        RECT 45.155 91.710 50.500 92.255 ;
        RECT 50.675 91.710 56.020 92.255 ;
        RECT 56.195 91.710 61.540 92.255 ;
        RECT 34.760 90.140 35.110 91.390 ;
        RECT 36.875 90.965 37.625 91.485 ;
        RECT 37.795 90.795 38.545 91.315 ;
        RECT 41.220 90.880 41.560 91.710 ;
        RECT 14.795 89.705 20.140 90.140 ;
        RECT 20.315 89.705 25.660 90.140 ;
        RECT 25.835 89.705 31.180 90.140 ;
        RECT 31.355 89.705 36.700 90.140 ;
        RECT 36.875 89.705 38.545 90.795 ;
        RECT 39.175 89.705 39.465 90.870 ;
        RECT 43.040 90.140 43.390 91.390 ;
        RECT 46.740 90.880 47.080 91.710 ;
        RECT 48.560 90.140 48.910 91.390 ;
        RECT 52.260 90.880 52.600 91.710 ;
        RECT 54.080 90.140 54.430 91.390 ;
        RECT 57.780 90.880 58.120 91.710 ;
        RECT 61.715 91.485 64.305 92.255 ;
        RECT 64.935 91.530 65.225 92.255 ;
        RECT 65.395 91.710 70.740 92.255 ;
        RECT 70.915 91.710 76.260 92.255 ;
        RECT 59.600 90.140 59.950 91.390 ;
        RECT 61.715 90.965 62.925 91.485 ;
        RECT 63.095 90.795 64.305 91.315 ;
        RECT 66.980 90.880 67.320 91.710 ;
        RECT 39.635 89.705 44.980 90.140 ;
        RECT 45.155 89.705 50.500 90.140 ;
        RECT 50.675 89.705 56.020 90.140 ;
        RECT 56.195 89.705 61.540 90.140 ;
        RECT 61.715 89.705 64.305 90.795 ;
        RECT 64.935 89.705 65.225 90.870 ;
        RECT 68.800 90.140 69.150 91.390 ;
        RECT 72.500 90.880 72.840 91.710 ;
        RECT 76.525 91.705 76.695 91.995 ;
        RECT 76.865 91.875 77.195 92.255 ;
        RECT 76.525 91.535 77.190 91.705 ;
        RECT 74.320 90.140 74.670 91.390 ;
        RECT 76.440 90.715 76.790 91.365 ;
        RECT 76.960 90.545 77.190 91.535 ;
        RECT 76.525 90.375 77.190 90.545 ;
        RECT 65.395 89.705 70.740 90.140 ;
        RECT 70.915 89.705 76.260 90.140 ;
        RECT 76.525 89.875 76.695 90.375 ;
        RECT 76.865 89.705 77.195 90.205 ;
        RECT 77.365 89.875 77.550 91.995 ;
        RECT 77.805 91.795 78.055 92.255 ;
        RECT 78.225 91.805 78.560 91.975 ;
        RECT 78.755 91.805 79.430 91.975 ;
        RECT 78.225 91.665 78.395 91.805 ;
        RECT 77.720 90.675 78.000 91.625 ;
        RECT 78.170 91.535 78.395 91.665 ;
        RECT 78.170 90.430 78.340 91.535 ;
        RECT 78.565 91.385 79.090 91.605 ;
        RECT 78.510 90.620 78.750 91.215 ;
        RECT 78.920 90.685 79.090 91.385 ;
        RECT 79.260 91.025 79.430 91.805 ;
        RECT 79.750 91.755 80.120 92.255 ;
        RECT 80.300 91.805 80.705 91.975 ;
        RECT 80.875 91.805 81.660 91.975 ;
        RECT 80.300 91.575 80.470 91.805 ;
        RECT 79.640 91.275 80.470 91.575 ;
        RECT 80.855 91.305 81.320 91.635 ;
        RECT 79.640 91.245 79.840 91.275 ;
        RECT 79.960 91.025 80.130 91.095 ;
        RECT 79.260 90.855 80.130 91.025 ;
        RECT 79.620 90.765 80.130 90.855 ;
        RECT 78.170 90.300 78.475 90.430 ;
        RECT 78.920 90.320 79.450 90.685 ;
        RECT 77.790 89.705 78.055 90.165 ;
        RECT 78.225 89.875 78.475 90.300 ;
        RECT 79.620 90.150 79.790 90.765 ;
        RECT 78.685 89.980 79.790 90.150 ;
        RECT 79.960 89.705 80.130 90.505 ;
        RECT 80.300 90.205 80.470 91.275 ;
        RECT 80.640 90.375 80.830 91.095 ;
        RECT 81.000 90.345 81.320 91.305 ;
        RECT 81.490 91.345 81.660 91.805 ;
        RECT 81.935 91.725 82.145 92.255 ;
        RECT 82.405 91.515 82.735 92.040 ;
        RECT 82.905 91.645 83.075 92.255 ;
        RECT 83.245 91.600 83.575 92.035 ;
        RECT 83.245 91.515 83.625 91.600 ;
        RECT 82.535 91.345 82.735 91.515 ;
        RECT 83.400 91.475 83.625 91.515 ;
        RECT 81.490 91.015 82.365 91.345 ;
        RECT 82.535 91.015 83.285 91.345 ;
        RECT 80.300 89.875 80.550 90.205 ;
        RECT 81.490 90.175 81.660 91.015 ;
        RECT 82.535 90.810 82.725 91.015 ;
        RECT 83.455 90.895 83.625 91.475 ;
        RECT 83.410 90.845 83.625 90.895 ;
        RECT 81.830 90.435 82.725 90.810 ;
        RECT 83.235 90.765 83.625 90.845 ;
        RECT 83.830 91.515 84.445 92.085 ;
        RECT 84.615 91.745 84.830 92.255 ;
        RECT 85.060 91.745 85.340 92.075 ;
        RECT 85.520 91.745 85.760 92.255 ;
        RECT 80.775 90.005 81.660 90.175 ;
        RECT 81.840 89.705 82.155 90.205 ;
        RECT 82.385 89.875 82.725 90.435 ;
        RECT 82.895 89.705 83.065 90.715 ;
        RECT 83.235 89.920 83.565 90.765 ;
        RECT 83.830 90.495 84.145 91.515 ;
        RECT 84.315 90.845 84.485 91.345 ;
        RECT 84.735 91.015 85.000 91.575 ;
        RECT 85.170 90.845 85.340 91.745 ;
        RECT 85.510 91.015 85.865 91.575 ;
        RECT 86.130 91.515 86.745 92.085 ;
        RECT 86.915 91.745 87.130 92.255 ;
        RECT 87.360 91.745 87.640 92.075 ;
        RECT 87.820 91.745 88.060 92.255 ;
        RECT 84.315 90.675 85.740 90.845 ;
        RECT 83.830 89.875 84.365 90.495 ;
        RECT 84.535 89.705 84.865 90.505 ;
        RECT 85.350 90.500 85.740 90.675 ;
        RECT 86.130 90.495 86.445 91.515 ;
        RECT 86.615 90.845 86.785 91.345 ;
        RECT 87.035 91.015 87.300 91.575 ;
        RECT 87.470 90.845 87.640 91.745 ;
        RECT 87.810 91.015 88.165 91.575 ;
        RECT 88.395 91.485 90.065 92.255 ;
        RECT 90.695 91.530 90.985 92.255 ;
        RECT 88.395 90.965 89.145 91.485 ;
        RECT 91.155 91.455 91.495 92.085 ;
        RECT 91.665 91.455 91.915 92.255 ;
        RECT 92.105 91.605 92.435 92.085 ;
        RECT 92.605 91.795 92.830 92.255 ;
        RECT 93.000 91.605 93.330 92.085 ;
        RECT 86.615 90.675 88.040 90.845 ;
        RECT 89.315 90.795 90.065 91.315 ;
        RECT 86.130 89.875 86.665 90.495 ;
        RECT 86.835 89.705 87.165 90.505 ;
        RECT 87.650 90.500 88.040 90.675 ;
        RECT 88.395 89.705 90.065 90.795 ;
        RECT 90.695 89.705 90.985 90.870 ;
        RECT 91.155 90.845 91.330 91.455 ;
        RECT 92.105 91.435 93.330 91.605 ;
        RECT 93.960 91.475 94.460 92.085 ;
        RECT 95.330 91.515 95.945 92.085 ;
        RECT 96.115 91.745 96.330 92.255 ;
        RECT 96.560 91.745 96.840 92.075 ;
        RECT 97.020 91.745 97.260 92.255 ;
        RECT 91.500 91.095 92.195 91.265 ;
        RECT 92.025 90.845 92.195 91.095 ;
        RECT 92.370 91.065 92.790 91.265 ;
        RECT 92.960 91.065 93.290 91.265 ;
        RECT 93.460 91.065 93.790 91.265 ;
        RECT 93.960 90.845 94.130 91.475 ;
        RECT 94.315 91.015 94.665 91.265 ;
        RECT 91.155 89.875 91.495 90.845 ;
        RECT 91.665 89.705 91.835 90.845 ;
        RECT 92.025 90.675 94.460 90.845 ;
        RECT 92.105 89.705 92.355 90.505 ;
        RECT 93.000 89.875 93.330 90.675 ;
        RECT 93.630 89.705 93.960 90.505 ;
        RECT 94.130 89.875 94.460 90.675 ;
        RECT 95.330 90.495 95.645 91.515 ;
        RECT 95.815 90.845 95.985 91.345 ;
        RECT 96.235 91.015 96.500 91.575 ;
        RECT 96.670 90.845 96.840 91.745 ;
        RECT 97.645 91.600 97.975 92.035 ;
        RECT 98.145 91.645 98.315 92.255 ;
        RECT 97.010 91.015 97.365 91.575 ;
        RECT 97.595 91.515 97.975 91.600 ;
        RECT 98.485 91.515 98.815 92.040 ;
        RECT 99.075 91.725 99.285 92.255 ;
        RECT 99.560 91.805 100.345 91.975 ;
        RECT 100.515 91.805 100.920 91.975 ;
        RECT 97.595 91.475 97.820 91.515 ;
        RECT 97.595 90.895 97.765 91.475 ;
        RECT 98.485 91.345 98.685 91.515 ;
        RECT 99.560 91.345 99.730 91.805 ;
        RECT 97.935 91.015 98.685 91.345 ;
        RECT 98.855 91.015 99.730 91.345 ;
        RECT 97.595 90.845 97.810 90.895 ;
        RECT 95.815 90.675 97.240 90.845 ;
        RECT 97.595 90.765 97.985 90.845 ;
        RECT 95.330 89.875 95.865 90.495 ;
        RECT 96.035 89.705 96.365 90.505 ;
        RECT 96.850 90.500 97.240 90.675 ;
        RECT 97.655 89.920 97.985 90.765 ;
        RECT 98.495 90.810 98.685 91.015 ;
        RECT 98.155 89.705 98.325 90.715 ;
        RECT 98.495 90.435 99.390 90.810 ;
        RECT 98.495 89.875 98.835 90.435 ;
        RECT 99.065 89.705 99.380 90.205 ;
        RECT 99.560 90.175 99.730 91.015 ;
        RECT 99.900 91.305 100.365 91.635 ;
        RECT 100.750 91.575 100.920 91.805 ;
        RECT 101.100 91.755 101.470 92.255 ;
        RECT 101.790 91.805 102.465 91.975 ;
        RECT 102.660 91.805 102.995 91.975 ;
        RECT 99.900 90.345 100.220 91.305 ;
        RECT 100.750 91.275 101.580 91.575 ;
        RECT 100.390 90.375 100.580 91.095 ;
        RECT 100.750 90.205 100.920 91.275 ;
        RECT 101.380 91.245 101.580 91.275 ;
        RECT 101.090 91.025 101.260 91.095 ;
        RECT 101.790 91.025 101.960 91.805 ;
        RECT 102.825 91.665 102.995 91.805 ;
        RECT 103.165 91.795 103.415 92.255 ;
        RECT 101.090 90.855 101.960 91.025 ;
        RECT 102.130 91.385 102.655 91.605 ;
        RECT 102.825 91.535 103.050 91.665 ;
        RECT 101.090 90.765 101.600 90.855 ;
        RECT 99.560 90.005 100.445 90.175 ;
        RECT 100.670 89.875 100.920 90.205 ;
        RECT 101.090 89.705 101.260 90.505 ;
        RECT 101.430 90.150 101.600 90.765 ;
        RECT 102.130 90.685 102.300 91.385 ;
        RECT 101.770 90.320 102.300 90.685 ;
        RECT 102.470 90.620 102.710 91.215 ;
        RECT 102.880 90.430 103.050 91.535 ;
        RECT 103.220 90.675 103.500 91.625 ;
        RECT 102.745 90.300 103.050 90.430 ;
        RECT 101.430 89.980 102.535 90.150 ;
        RECT 102.745 89.875 102.995 90.300 ;
        RECT 103.165 89.705 103.430 90.165 ;
        RECT 103.670 89.875 103.855 91.995 ;
        RECT 104.025 91.875 104.355 92.255 ;
        RECT 104.525 91.705 104.695 91.995 ;
        RECT 105.120 91.745 105.360 92.255 ;
        RECT 105.540 91.745 105.820 92.075 ;
        RECT 106.050 91.745 106.265 92.255 ;
        RECT 104.030 91.535 104.695 91.705 ;
        RECT 104.030 90.545 104.260 91.535 ;
        RECT 104.430 90.715 104.780 91.365 ;
        RECT 105.015 91.015 105.370 91.575 ;
        RECT 105.540 90.845 105.710 91.745 ;
        RECT 105.880 91.015 106.145 91.575 ;
        RECT 106.435 91.515 107.050 92.085 ;
        RECT 106.395 90.845 106.565 91.345 ;
        RECT 105.140 90.675 106.565 90.845 ;
        RECT 104.030 90.375 104.695 90.545 ;
        RECT 105.140 90.500 105.530 90.675 ;
        RECT 104.025 89.705 104.355 90.205 ;
        RECT 104.525 89.875 104.695 90.375 ;
        RECT 106.015 89.705 106.345 90.505 ;
        RECT 106.735 90.495 107.050 91.515 ;
        RECT 107.255 91.485 108.925 92.255 ;
        RECT 109.095 91.755 109.355 92.085 ;
        RECT 109.525 91.895 109.855 92.255 ;
        RECT 110.110 91.875 111.410 92.085 ;
        RECT 109.095 91.745 109.325 91.755 ;
        RECT 107.255 90.965 108.005 91.485 ;
        RECT 108.175 90.795 108.925 91.315 ;
        RECT 106.515 89.875 107.050 90.495 ;
        RECT 107.255 89.705 108.925 90.795 ;
        RECT 109.095 90.555 109.265 91.745 ;
        RECT 110.110 91.725 110.280 91.875 ;
        RECT 109.525 91.600 110.280 91.725 ;
        RECT 109.435 91.555 110.280 91.600 ;
        RECT 109.435 91.435 109.705 91.555 ;
        RECT 109.435 90.860 109.605 91.435 ;
        RECT 109.835 90.995 110.245 91.300 ;
        RECT 110.535 91.265 110.745 91.665 ;
        RECT 110.415 91.055 110.745 91.265 ;
        RECT 110.990 91.265 111.210 91.665 ;
        RECT 111.685 91.490 112.140 92.255 ;
        RECT 112.320 91.490 112.775 92.255 ;
        RECT 113.050 91.875 114.350 92.085 ;
        RECT 114.605 91.895 114.935 92.255 ;
        RECT 114.180 91.725 114.350 91.875 ;
        RECT 115.105 91.755 115.365 92.085 ;
        RECT 115.135 91.745 115.365 91.755 ;
        RECT 113.250 91.265 113.470 91.665 ;
        RECT 110.990 91.055 111.465 91.265 ;
        RECT 111.655 91.065 112.145 91.265 ;
        RECT 112.315 91.065 112.805 91.265 ;
        RECT 112.995 91.055 113.470 91.265 ;
        RECT 113.715 91.265 113.925 91.665 ;
        RECT 114.180 91.600 114.935 91.725 ;
        RECT 114.180 91.555 115.025 91.600 ;
        RECT 114.755 91.435 115.025 91.555 ;
        RECT 113.715 91.055 114.045 91.265 ;
        RECT 114.215 90.995 114.625 91.300 ;
        RECT 109.435 90.825 109.635 90.860 ;
        RECT 110.965 90.825 112.140 90.885 ;
        RECT 109.435 90.715 112.140 90.825 ;
        RECT 109.495 90.655 111.295 90.715 ;
        RECT 110.965 90.625 111.295 90.655 ;
        RECT 109.095 89.875 109.355 90.555 ;
        RECT 109.525 89.705 109.775 90.485 ;
        RECT 110.025 90.455 110.860 90.465 ;
        RECT 111.450 90.455 111.635 90.545 ;
        RECT 110.025 90.255 111.635 90.455 ;
        RECT 110.025 89.875 110.275 90.255 ;
        RECT 111.405 90.215 111.635 90.255 ;
        RECT 111.885 90.095 112.140 90.715 ;
        RECT 110.445 89.705 110.800 90.085 ;
        RECT 111.805 89.875 112.140 90.095 ;
        RECT 112.320 90.825 113.495 90.885 ;
        RECT 114.855 90.860 115.025 91.435 ;
        RECT 114.825 90.825 115.025 90.860 ;
        RECT 112.320 90.715 115.025 90.825 ;
        RECT 112.320 90.095 112.575 90.715 ;
        RECT 113.165 90.655 114.965 90.715 ;
        RECT 113.165 90.625 113.495 90.655 ;
        RECT 115.195 90.555 115.365 91.745 ;
        RECT 116.455 91.530 116.745 92.255 ;
        RECT 116.915 91.455 117.255 92.085 ;
        RECT 117.425 91.455 117.675 92.255 ;
        RECT 117.865 91.605 118.195 92.085 ;
        RECT 118.365 91.795 118.590 92.255 ;
        RECT 118.760 91.605 119.090 92.085 ;
        RECT 112.825 90.455 113.010 90.545 ;
        RECT 113.600 90.455 114.435 90.465 ;
        RECT 112.825 90.255 114.435 90.455 ;
        RECT 112.825 90.215 113.055 90.255 ;
        RECT 112.320 89.875 112.655 90.095 ;
        RECT 113.660 89.705 114.015 90.085 ;
        RECT 114.185 89.875 114.435 90.255 ;
        RECT 114.685 89.705 114.935 90.485 ;
        RECT 115.105 89.875 115.365 90.555 ;
        RECT 116.455 89.705 116.745 90.870 ;
        RECT 116.915 90.845 117.090 91.455 ;
        RECT 117.865 91.435 119.090 91.605 ;
        RECT 119.720 91.475 120.220 92.085 ;
        RECT 121.145 91.705 121.315 91.995 ;
        RECT 121.485 91.875 121.815 92.255 ;
        RECT 121.145 91.535 121.810 91.705 ;
        RECT 117.260 91.095 117.955 91.265 ;
        RECT 117.785 90.845 117.955 91.095 ;
        RECT 118.130 91.065 118.550 91.265 ;
        RECT 118.720 91.065 119.050 91.265 ;
        RECT 119.220 91.065 119.550 91.265 ;
        RECT 119.720 90.845 119.890 91.475 ;
        RECT 120.075 91.015 120.425 91.265 ;
        RECT 116.915 89.875 117.255 90.845 ;
        RECT 117.425 89.705 117.595 90.845 ;
        RECT 117.785 90.675 120.220 90.845 ;
        RECT 121.060 90.715 121.410 91.365 ;
        RECT 117.865 89.705 118.115 90.505 ;
        RECT 118.760 89.875 119.090 90.675 ;
        RECT 119.390 89.705 119.720 90.505 ;
        RECT 119.890 89.875 120.220 90.675 ;
        RECT 121.580 90.545 121.810 91.535 ;
        RECT 121.145 90.375 121.810 90.545 ;
        RECT 121.145 89.875 121.315 90.375 ;
        RECT 121.485 89.705 121.815 90.205 ;
        RECT 121.985 89.875 122.170 91.995 ;
        RECT 122.425 91.795 122.675 92.255 ;
        RECT 122.845 91.805 123.180 91.975 ;
        RECT 123.375 91.805 124.050 91.975 ;
        RECT 122.845 91.665 123.015 91.805 ;
        RECT 122.340 90.675 122.620 91.625 ;
        RECT 122.790 91.535 123.015 91.665 ;
        RECT 122.790 90.430 122.960 91.535 ;
        RECT 123.185 91.385 123.710 91.605 ;
        RECT 123.130 90.620 123.370 91.215 ;
        RECT 123.540 90.685 123.710 91.385 ;
        RECT 123.880 91.025 124.050 91.805 ;
        RECT 124.370 91.755 124.740 92.255 ;
        RECT 124.920 91.805 125.325 91.975 ;
        RECT 125.495 91.805 126.280 91.975 ;
        RECT 124.920 91.575 125.090 91.805 ;
        RECT 124.260 91.275 125.090 91.575 ;
        RECT 125.475 91.305 125.940 91.635 ;
        RECT 124.260 91.245 124.460 91.275 ;
        RECT 124.580 91.025 124.750 91.095 ;
        RECT 123.880 90.855 124.750 91.025 ;
        RECT 124.240 90.765 124.750 90.855 ;
        RECT 122.790 90.300 123.095 90.430 ;
        RECT 123.540 90.320 124.070 90.685 ;
        RECT 122.410 89.705 122.675 90.165 ;
        RECT 122.845 89.875 123.095 90.300 ;
        RECT 124.240 90.150 124.410 90.765 ;
        RECT 123.305 89.980 124.410 90.150 ;
        RECT 124.580 89.705 124.750 90.505 ;
        RECT 124.920 90.205 125.090 91.275 ;
        RECT 125.260 90.375 125.450 91.095 ;
        RECT 125.620 90.345 125.940 91.305 ;
        RECT 126.110 91.345 126.280 91.805 ;
        RECT 126.555 91.725 126.765 92.255 ;
        RECT 127.025 91.515 127.355 92.040 ;
        RECT 127.525 91.645 127.695 92.255 ;
        RECT 127.865 91.600 128.195 92.035 ;
        RECT 128.580 91.745 128.820 92.255 ;
        RECT 129.000 91.745 129.280 92.075 ;
        RECT 129.510 91.745 129.725 92.255 ;
        RECT 127.865 91.515 128.245 91.600 ;
        RECT 127.155 91.345 127.355 91.515 ;
        RECT 128.020 91.475 128.245 91.515 ;
        RECT 126.110 91.015 126.985 91.345 ;
        RECT 127.155 91.015 127.905 91.345 ;
        RECT 124.920 89.875 125.170 90.205 ;
        RECT 126.110 90.175 126.280 91.015 ;
        RECT 127.155 90.810 127.345 91.015 ;
        RECT 128.075 90.895 128.245 91.475 ;
        RECT 128.475 91.015 128.830 91.575 ;
        RECT 128.030 90.845 128.245 90.895 ;
        RECT 129.000 90.845 129.170 91.745 ;
        RECT 129.340 91.015 129.605 91.575 ;
        RECT 129.895 91.515 130.510 92.085 ;
        RECT 129.855 90.845 130.025 91.345 ;
        RECT 126.450 90.435 127.345 90.810 ;
        RECT 127.855 90.765 128.245 90.845 ;
        RECT 125.395 90.005 126.280 90.175 ;
        RECT 126.460 89.705 126.775 90.205 ;
        RECT 127.005 89.875 127.345 90.435 ;
        RECT 127.515 89.705 127.685 90.715 ;
        RECT 127.855 89.920 128.185 90.765 ;
        RECT 128.600 90.675 130.025 90.845 ;
        RECT 128.600 90.500 128.990 90.675 ;
        RECT 129.475 89.705 129.805 90.505 ;
        RECT 130.195 90.495 130.510 91.515 ;
        RECT 130.715 91.485 134.225 92.255 ;
        RECT 134.395 91.505 135.605 92.255 ;
        RECT 135.865 91.705 136.035 92.085 ;
        RECT 136.250 91.875 136.580 92.255 ;
        RECT 135.865 91.535 136.580 91.705 ;
        RECT 130.715 90.965 132.365 91.485 ;
        RECT 132.535 90.795 134.225 91.315 ;
        RECT 134.395 90.965 134.915 91.505 ;
        RECT 135.085 90.795 135.605 91.335 ;
        RECT 135.775 90.985 136.130 91.355 ;
        RECT 136.410 91.345 136.580 91.535 ;
        RECT 136.750 91.510 137.005 92.085 ;
        RECT 136.410 91.015 136.665 91.345 ;
        RECT 136.410 90.805 136.580 91.015 ;
        RECT 129.975 89.875 130.510 90.495 ;
        RECT 130.715 89.705 134.225 90.795 ;
        RECT 134.395 89.705 135.605 90.795 ;
        RECT 135.865 90.635 136.580 90.805 ;
        RECT 136.835 90.780 137.005 91.510 ;
        RECT 137.180 91.415 137.440 92.255 ;
        RECT 137.615 91.505 138.825 92.255 ;
        RECT 135.865 89.875 136.035 90.635 ;
        RECT 136.250 89.705 136.580 90.465 ;
        RECT 136.750 89.875 137.005 90.780 ;
        RECT 137.180 89.705 137.440 90.855 ;
        RECT 137.615 90.795 138.135 91.335 ;
        RECT 138.305 90.965 138.825 91.505 ;
        RECT 137.615 89.705 138.825 90.795 ;
        RECT 13.330 89.535 138.910 89.705 ;
        RECT 13.415 88.445 14.625 89.535 ;
        RECT 14.795 89.100 20.140 89.535 ;
        RECT 20.315 89.100 25.660 89.535 ;
        RECT 13.415 87.735 13.935 88.275 ;
        RECT 14.105 87.905 14.625 88.445 ;
        RECT 13.415 86.985 14.625 87.735 ;
        RECT 16.380 87.530 16.720 88.360 ;
        RECT 18.200 87.850 18.550 89.100 ;
        RECT 21.900 87.530 22.240 88.360 ;
        RECT 23.720 87.850 24.070 89.100 ;
        RECT 26.295 88.370 26.585 89.535 ;
        RECT 26.755 89.100 32.100 89.535 ;
        RECT 32.275 89.100 37.620 89.535 ;
        RECT 14.795 86.985 20.140 87.530 ;
        RECT 20.315 86.985 25.660 87.530 ;
        RECT 26.295 86.985 26.585 87.710 ;
        RECT 28.340 87.530 28.680 88.360 ;
        RECT 30.160 87.850 30.510 89.100 ;
        RECT 33.860 87.530 34.200 88.360 ;
        RECT 35.680 87.850 36.030 89.100 ;
        RECT 37.795 88.445 39.005 89.535 ;
        RECT 37.795 87.735 38.315 88.275 ;
        RECT 38.485 87.905 39.005 88.445 ;
        RECT 39.175 88.370 39.465 89.535 ;
        RECT 39.635 89.100 44.980 89.535 ;
        RECT 45.155 89.100 50.500 89.535 ;
        RECT 26.755 86.985 32.100 87.530 ;
        RECT 32.275 86.985 37.620 87.530 ;
        RECT 37.795 86.985 39.005 87.735 ;
        RECT 39.175 86.985 39.465 87.710 ;
        RECT 41.220 87.530 41.560 88.360 ;
        RECT 43.040 87.850 43.390 89.100 ;
        RECT 46.740 87.530 47.080 88.360 ;
        RECT 48.560 87.850 48.910 89.100 ;
        RECT 50.675 88.445 51.885 89.535 ;
        RECT 50.675 87.735 51.195 88.275 ;
        RECT 51.365 87.905 51.885 88.445 ;
        RECT 52.055 88.370 52.345 89.535 ;
        RECT 52.515 89.100 57.860 89.535 ;
        RECT 39.635 86.985 44.980 87.530 ;
        RECT 45.155 86.985 50.500 87.530 ;
        RECT 50.675 86.985 51.885 87.735 ;
        RECT 52.055 86.985 52.345 87.710 ;
        RECT 54.100 87.530 54.440 88.360 ;
        RECT 55.920 87.850 56.270 89.100 ;
        RECT 58.035 88.445 59.705 89.535 ;
        RECT 58.035 87.755 58.785 88.275 ;
        RECT 58.955 87.925 59.705 88.445 ;
        RECT 59.965 88.605 60.135 89.365 ;
        RECT 60.350 88.775 60.680 89.535 ;
        RECT 59.965 88.435 60.680 88.605 ;
        RECT 60.850 88.460 61.105 89.365 ;
        RECT 59.875 87.885 60.230 88.255 ;
        RECT 60.510 88.225 60.680 88.435 ;
        RECT 60.510 87.895 60.765 88.225 ;
        RECT 52.515 86.985 57.860 87.530 ;
        RECT 58.035 86.985 59.705 87.755 ;
        RECT 60.510 87.705 60.680 87.895 ;
        RECT 60.935 87.730 61.105 88.460 ;
        RECT 61.280 88.385 61.540 89.535 ;
        RECT 61.715 88.445 64.305 89.535 ;
        RECT 59.965 87.535 60.680 87.705 ;
        RECT 59.965 87.155 60.135 87.535 ;
        RECT 60.350 86.985 60.680 87.365 ;
        RECT 60.850 87.155 61.105 87.730 ;
        RECT 61.280 86.985 61.540 87.825 ;
        RECT 61.715 87.755 62.925 88.275 ;
        RECT 63.095 87.925 64.305 88.445 ;
        RECT 64.935 88.370 65.225 89.535 ;
        RECT 66.320 88.385 66.580 89.535 ;
        RECT 66.755 88.460 67.010 89.365 ;
        RECT 67.180 88.775 67.510 89.535 ;
        RECT 67.725 88.605 67.895 89.365 ;
        RECT 61.715 86.985 64.305 87.755 ;
        RECT 64.935 86.985 65.225 87.710 ;
        RECT 66.320 86.985 66.580 87.825 ;
        RECT 66.755 87.730 66.925 88.460 ;
        RECT 67.180 88.435 67.895 88.605 ;
        RECT 68.155 88.445 69.365 89.535 ;
        RECT 69.535 88.940 69.970 89.365 ;
        RECT 70.140 89.110 70.525 89.535 ;
        RECT 69.535 88.770 70.525 88.940 ;
        RECT 67.180 88.225 67.350 88.435 ;
        RECT 67.095 87.895 67.350 88.225 ;
        RECT 66.755 87.155 67.010 87.730 ;
        RECT 67.180 87.705 67.350 87.895 ;
        RECT 67.630 87.885 67.985 88.255 ;
        RECT 68.155 87.735 68.675 88.275 ;
        RECT 68.845 87.905 69.365 88.445 ;
        RECT 69.535 87.895 70.020 88.600 ;
        RECT 70.190 88.225 70.525 88.770 ;
        RECT 70.695 88.575 71.120 89.365 ;
        RECT 71.290 88.940 71.565 89.365 ;
        RECT 71.735 89.110 72.120 89.535 ;
        RECT 71.290 88.745 72.120 88.940 ;
        RECT 70.695 88.395 71.600 88.575 ;
        RECT 70.190 87.895 70.600 88.225 ;
        RECT 70.770 87.895 71.600 88.395 ;
        RECT 71.770 88.225 72.120 88.745 ;
        RECT 72.290 88.575 72.535 89.365 ;
        RECT 72.725 88.940 72.980 89.365 ;
        RECT 73.150 89.110 73.535 89.535 ;
        RECT 72.725 88.745 73.535 88.940 ;
        RECT 72.290 88.395 73.015 88.575 ;
        RECT 71.770 87.895 72.195 88.225 ;
        RECT 72.365 87.895 73.015 88.395 ;
        RECT 73.185 88.225 73.535 88.745 ;
        RECT 73.705 88.395 73.965 89.365 ;
        RECT 73.185 87.895 73.610 88.225 ;
        RECT 67.180 87.535 67.895 87.705 ;
        RECT 67.180 86.985 67.510 87.365 ;
        RECT 67.725 87.155 67.895 87.535 ;
        RECT 68.155 86.985 69.365 87.735 ;
        RECT 70.190 87.725 70.525 87.895 ;
        RECT 70.770 87.725 71.120 87.895 ;
        RECT 71.770 87.725 72.120 87.895 ;
        RECT 72.365 87.725 72.535 87.895 ;
        RECT 73.185 87.725 73.535 87.895 ;
        RECT 73.780 87.725 73.965 88.395 ;
        RECT 74.140 88.385 74.400 89.535 ;
        RECT 74.575 88.460 74.830 89.365 ;
        RECT 75.000 88.775 75.330 89.535 ;
        RECT 75.545 88.605 75.715 89.365 ;
        RECT 69.535 87.555 70.525 87.725 ;
        RECT 69.535 87.155 69.970 87.555 ;
        RECT 70.140 86.985 70.525 87.385 ;
        RECT 70.695 87.155 71.120 87.725 ;
        RECT 71.310 87.555 72.120 87.725 ;
        RECT 71.310 87.155 71.565 87.555 ;
        RECT 71.735 86.985 72.120 87.385 ;
        RECT 72.290 87.155 72.535 87.725 ;
        RECT 72.725 87.555 73.535 87.725 ;
        RECT 72.725 87.155 72.980 87.555 ;
        RECT 73.150 86.985 73.535 87.385 ;
        RECT 73.705 87.155 73.965 87.725 ;
        RECT 74.140 86.985 74.400 87.825 ;
        RECT 74.575 87.730 74.745 88.460 ;
        RECT 75.000 88.435 75.715 88.605 ;
        RECT 75.000 88.225 75.170 88.435 ;
        RECT 75.980 88.385 76.240 89.535 ;
        RECT 76.415 88.460 76.670 89.365 ;
        RECT 76.840 88.775 77.170 89.535 ;
        RECT 77.385 88.605 77.555 89.365 ;
        RECT 74.915 87.895 75.170 88.225 ;
        RECT 74.575 87.155 74.830 87.730 ;
        RECT 75.000 87.705 75.170 87.895 ;
        RECT 75.450 87.885 75.805 88.255 ;
        RECT 75.000 87.535 75.715 87.705 ;
        RECT 75.000 86.985 75.330 87.365 ;
        RECT 75.545 87.155 75.715 87.535 ;
        RECT 75.980 86.985 76.240 87.825 ;
        RECT 76.415 87.730 76.585 88.460 ;
        RECT 76.840 88.435 77.555 88.605 ;
        RECT 76.840 88.225 77.010 88.435 ;
        RECT 77.815 88.370 78.105 89.535 ;
        RECT 79.200 88.385 79.460 89.535 ;
        RECT 79.635 88.460 79.890 89.365 ;
        RECT 80.060 88.775 80.390 89.535 ;
        RECT 80.605 88.605 80.775 89.365 ;
        RECT 76.755 87.895 77.010 88.225 ;
        RECT 76.415 87.155 76.670 87.730 ;
        RECT 76.840 87.705 77.010 87.895 ;
        RECT 77.290 87.885 77.645 88.255 ;
        RECT 76.840 87.535 77.555 87.705 ;
        RECT 76.840 86.985 77.170 87.365 ;
        RECT 77.385 87.155 77.555 87.535 ;
        RECT 77.815 86.985 78.105 87.710 ;
        RECT 79.200 86.985 79.460 87.825 ;
        RECT 79.635 87.730 79.805 88.460 ;
        RECT 80.060 88.435 80.775 88.605 ;
        RECT 81.035 88.445 82.245 89.535 ;
        RECT 80.060 88.225 80.230 88.435 ;
        RECT 79.975 87.895 80.230 88.225 ;
        RECT 79.635 87.155 79.890 87.730 ;
        RECT 80.060 87.705 80.230 87.895 ;
        RECT 80.510 87.885 80.865 88.255 ;
        RECT 81.035 87.735 81.555 88.275 ;
        RECT 81.725 87.905 82.245 88.445 ;
        RECT 82.420 88.385 82.680 89.535 ;
        RECT 82.855 88.460 83.110 89.365 ;
        RECT 83.280 88.775 83.610 89.535 ;
        RECT 83.825 88.605 83.995 89.365 ;
        RECT 80.060 87.535 80.775 87.705 ;
        RECT 80.060 86.985 80.390 87.365 ;
        RECT 80.605 87.155 80.775 87.535 ;
        RECT 81.035 86.985 82.245 87.735 ;
        RECT 82.420 86.985 82.680 87.825 ;
        RECT 82.855 87.730 83.025 88.460 ;
        RECT 83.280 88.435 83.995 88.605 ;
        RECT 84.255 88.445 85.465 89.535 ;
        RECT 83.280 88.225 83.450 88.435 ;
        RECT 83.195 87.895 83.450 88.225 ;
        RECT 82.855 87.155 83.110 87.730 ;
        RECT 83.280 87.705 83.450 87.895 ;
        RECT 83.730 87.885 84.085 88.255 ;
        RECT 84.255 87.735 84.775 88.275 ;
        RECT 84.945 87.905 85.465 88.445 ;
        RECT 85.640 88.385 85.900 89.535 ;
        RECT 86.075 88.460 86.330 89.365 ;
        RECT 86.500 88.775 86.830 89.535 ;
        RECT 87.045 88.605 87.215 89.365 ;
        RECT 83.280 87.535 83.995 87.705 ;
        RECT 83.280 86.985 83.610 87.365 ;
        RECT 83.825 87.155 83.995 87.535 ;
        RECT 84.255 86.985 85.465 87.735 ;
        RECT 85.640 86.985 85.900 87.825 ;
        RECT 86.075 87.730 86.245 88.460 ;
        RECT 86.500 88.435 87.215 88.605 ;
        RECT 87.475 88.445 88.685 89.535 ;
        RECT 86.500 88.225 86.670 88.435 ;
        RECT 86.415 87.895 86.670 88.225 ;
        RECT 86.075 87.155 86.330 87.730 ;
        RECT 86.500 87.705 86.670 87.895 ;
        RECT 86.950 87.885 87.305 88.255 ;
        RECT 87.475 87.735 87.995 88.275 ;
        RECT 88.165 87.905 88.685 88.445 ;
        RECT 88.860 88.385 89.120 89.535 ;
        RECT 89.295 88.460 89.550 89.365 ;
        RECT 89.720 88.775 90.050 89.535 ;
        RECT 90.265 88.605 90.435 89.365 ;
        RECT 86.500 87.535 87.215 87.705 ;
        RECT 86.500 86.985 86.830 87.365 ;
        RECT 87.045 87.155 87.215 87.535 ;
        RECT 87.475 86.985 88.685 87.735 ;
        RECT 88.860 86.985 89.120 87.825 ;
        RECT 89.295 87.730 89.465 88.460 ;
        RECT 89.720 88.435 90.435 88.605 ;
        RECT 89.720 88.225 89.890 88.435 ;
        RECT 90.695 88.370 90.985 89.535 ;
        RECT 92.080 88.385 92.340 89.535 ;
        RECT 92.515 88.460 92.770 89.365 ;
        RECT 92.940 88.775 93.270 89.535 ;
        RECT 93.485 88.605 93.655 89.365 ;
        RECT 89.635 87.895 89.890 88.225 ;
        RECT 89.295 87.155 89.550 87.730 ;
        RECT 89.720 87.705 89.890 87.895 ;
        RECT 90.170 87.885 90.525 88.255 ;
        RECT 89.720 87.535 90.435 87.705 ;
        RECT 89.720 86.985 90.050 87.365 ;
        RECT 90.265 87.155 90.435 87.535 ;
        RECT 90.695 86.985 90.985 87.710 ;
        RECT 92.080 86.985 92.340 87.825 ;
        RECT 92.515 87.730 92.685 88.460 ;
        RECT 92.940 88.435 93.655 88.605 ;
        RECT 93.915 88.445 95.125 89.535 ;
        RECT 92.940 88.225 93.110 88.435 ;
        RECT 92.855 87.895 93.110 88.225 ;
        RECT 92.515 87.155 92.770 87.730 ;
        RECT 92.940 87.705 93.110 87.895 ;
        RECT 93.390 87.885 93.745 88.255 ;
        RECT 93.915 87.735 94.435 88.275 ;
        RECT 94.605 87.905 95.125 88.445 ;
        RECT 95.300 88.385 95.560 89.535 ;
        RECT 95.735 88.460 95.990 89.365 ;
        RECT 96.160 88.775 96.490 89.535 ;
        RECT 96.705 88.605 96.875 89.365 ;
        RECT 92.940 87.535 93.655 87.705 ;
        RECT 92.940 86.985 93.270 87.365 ;
        RECT 93.485 87.155 93.655 87.535 ;
        RECT 93.915 86.985 95.125 87.735 ;
        RECT 95.300 86.985 95.560 87.825 ;
        RECT 95.735 87.730 95.905 88.460 ;
        RECT 96.160 88.435 96.875 88.605 ;
        RECT 96.160 88.225 96.330 88.435 ;
        RECT 98.060 88.385 98.320 89.535 ;
        RECT 98.495 88.460 98.750 89.365 ;
        RECT 98.920 88.775 99.250 89.535 ;
        RECT 99.465 88.605 99.635 89.365 ;
        RECT 96.075 87.895 96.330 88.225 ;
        RECT 95.735 87.155 95.990 87.730 ;
        RECT 96.160 87.705 96.330 87.895 ;
        RECT 96.610 87.885 96.965 88.255 ;
        RECT 96.160 87.535 96.875 87.705 ;
        RECT 96.160 86.985 96.490 87.365 ;
        RECT 96.705 87.155 96.875 87.535 ;
        RECT 98.060 86.985 98.320 87.825 ;
        RECT 98.495 87.730 98.665 88.460 ;
        RECT 98.920 88.435 99.635 88.605 ;
        RECT 100.080 88.565 100.470 88.740 ;
        RECT 100.955 88.735 101.285 89.535 ;
        RECT 101.455 88.745 101.990 89.365 ;
        RECT 98.920 88.225 99.090 88.435 ;
        RECT 100.080 88.395 101.505 88.565 ;
        RECT 98.835 87.895 99.090 88.225 ;
        RECT 98.495 87.155 98.750 87.730 ;
        RECT 98.920 87.705 99.090 87.895 ;
        RECT 99.370 87.885 99.725 88.255 ;
        RECT 98.920 87.535 99.635 87.705 ;
        RECT 99.955 87.665 100.310 88.225 ;
        RECT 98.920 86.985 99.250 87.365 ;
        RECT 99.465 87.155 99.635 87.535 ;
        RECT 100.480 87.495 100.650 88.395 ;
        RECT 100.820 87.665 101.085 88.225 ;
        RECT 101.335 87.895 101.505 88.395 ;
        RECT 101.675 87.725 101.990 88.745 ;
        RECT 102.195 88.445 103.405 89.535 ;
        RECT 100.060 86.985 100.300 87.495 ;
        RECT 100.480 87.165 100.760 87.495 ;
        RECT 100.990 86.985 101.205 87.495 ;
        RECT 101.375 87.155 101.990 87.725 ;
        RECT 102.195 87.735 102.715 88.275 ;
        RECT 102.885 87.905 103.405 88.445 ;
        RECT 103.575 88.370 103.865 89.535 ;
        RECT 104.040 88.385 104.300 89.535 ;
        RECT 104.475 88.460 104.730 89.365 ;
        RECT 104.900 88.775 105.230 89.535 ;
        RECT 105.445 88.605 105.615 89.365 ;
        RECT 102.195 86.985 103.405 87.735 ;
        RECT 103.575 86.985 103.865 87.710 ;
        RECT 104.040 86.985 104.300 87.825 ;
        RECT 104.475 87.730 104.645 88.460 ;
        RECT 104.900 88.435 105.615 88.605 ;
        RECT 104.900 88.225 105.070 88.435 ;
        RECT 105.880 88.385 106.140 89.535 ;
        RECT 106.315 88.460 106.570 89.365 ;
        RECT 106.740 88.775 107.070 89.535 ;
        RECT 107.285 88.605 107.455 89.365 ;
        RECT 104.815 87.895 105.070 88.225 ;
        RECT 104.475 87.155 104.730 87.730 ;
        RECT 104.900 87.705 105.070 87.895 ;
        RECT 105.350 87.885 105.705 88.255 ;
        RECT 104.900 87.535 105.615 87.705 ;
        RECT 104.900 86.985 105.230 87.365 ;
        RECT 105.445 87.155 105.615 87.535 ;
        RECT 105.880 86.985 106.140 87.825 ;
        RECT 106.315 87.730 106.485 88.460 ;
        RECT 106.740 88.435 107.455 88.605 ;
        RECT 106.740 88.225 106.910 88.435 ;
        RECT 108.180 88.385 108.440 89.535 ;
        RECT 108.615 88.460 108.870 89.365 ;
        RECT 109.040 88.775 109.370 89.535 ;
        RECT 109.585 88.605 109.755 89.365 ;
        RECT 106.655 87.895 106.910 88.225 ;
        RECT 106.315 87.155 106.570 87.730 ;
        RECT 106.740 87.705 106.910 87.895 ;
        RECT 107.190 87.885 107.545 88.255 ;
        RECT 106.740 87.535 107.455 87.705 ;
        RECT 106.740 86.985 107.070 87.365 ;
        RECT 107.285 87.155 107.455 87.535 ;
        RECT 108.180 86.985 108.440 87.825 ;
        RECT 108.615 87.730 108.785 88.460 ;
        RECT 109.040 88.435 109.755 88.605 ;
        RECT 110.015 88.445 111.225 89.535 ;
        RECT 109.040 88.225 109.210 88.435 ;
        RECT 108.955 87.895 109.210 88.225 ;
        RECT 108.615 87.155 108.870 87.730 ;
        RECT 109.040 87.705 109.210 87.895 ;
        RECT 109.490 87.885 109.845 88.255 ;
        RECT 110.015 87.735 110.535 88.275 ;
        RECT 110.705 87.905 111.225 88.445 ;
        RECT 111.485 88.605 111.655 89.365 ;
        RECT 111.870 88.775 112.200 89.535 ;
        RECT 111.485 88.435 112.200 88.605 ;
        RECT 112.370 88.460 112.625 89.365 ;
        RECT 111.395 87.885 111.750 88.255 ;
        RECT 112.030 88.225 112.200 88.435 ;
        RECT 112.030 87.895 112.285 88.225 ;
        RECT 109.040 87.535 109.755 87.705 ;
        RECT 109.040 86.985 109.370 87.365 ;
        RECT 109.585 87.155 109.755 87.535 ;
        RECT 110.015 86.985 111.225 87.735 ;
        RECT 112.030 87.705 112.200 87.895 ;
        RECT 112.455 87.730 112.625 88.460 ;
        RECT 112.800 88.385 113.060 89.535 ;
        RECT 113.880 88.565 114.270 88.740 ;
        RECT 114.755 88.735 115.085 89.535 ;
        RECT 115.255 88.745 115.790 89.365 ;
        RECT 113.880 88.395 115.305 88.565 ;
        RECT 111.485 87.535 112.200 87.705 ;
        RECT 111.485 87.155 111.655 87.535 ;
        RECT 111.870 86.985 112.200 87.365 ;
        RECT 112.370 87.155 112.625 87.730 ;
        RECT 112.800 86.985 113.060 87.825 ;
        RECT 113.755 87.665 114.110 88.225 ;
        RECT 114.280 87.495 114.450 88.395 ;
        RECT 114.620 87.665 114.885 88.225 ;
        RECT 115.135 87.895 115.305 88.395 ;
        RECT 115.475 87.725 115.790 88.745 ;
        RECT 116.455 88.370 116.745 89.535 ;
        RECT 117.005 88.605 117.175 89.365 ;
        RECT 117.390 88.775 117.720 89.535 ;
        RECT 117.005 88.435 117.720 88.605 ;
        RECT 117.890 88.460 118.145 89.365 ;
        RECT 116.915 87.885 117.270 88.255 ;
        RECT 117.550 88.225 117.720 88.435 ;
        RECT 117.550 87.895 117.805 88.225 ;
        RECT 113.860 86.985 114.100 87.495 ;
        RECT 114.280 87.165 114.560 87.495 ;
        RECT 114.790 86.985 115.005 87.495 ;
        RECT 115.175 87.155 115.790 87.725 ;
        RECT 116.455 86.985 116.745 87.710 ;
        RECT 117.550 87.705 117.720 87.895 ;
        RECT 117.975 87.730 118.145 88.460 ;
        RECT 118.320 88.385 118.580 89.535 ;
        RECT 118.845 88.605 119.015 89.365 ;
        RECT 119.230 88.775 119.560 89.535 ;
        RECT 118.845 88.435 119.560 88.605 ;
        RECT 119.730 88.460 119.985 89.365 ;
        RECT 118.755 87.885 119.110 88.255 ;
        RECT 119.390 88.225 119.560 88.435 ;
        RECT 119.390 87.895 119.645 88.225 ;
        RECT 117.005 87.535 117.720 87.705 ;
        RECT 117.005 87.155 117.175 87.535 ;
        RECT 117.390 86.985 117.720 87.365 ;
        RECT 117.890 87.155 118.145 87.730 ;
        RECT 118.320 86.985 118.580 87.825 ;
        RECT 119.390 87.705 119.560 87.895 ;
        RECT 119.815 87.730 119.985 88.460 ;
        RECT 120.160 88.385 120.420 89.535 ;
        RECT 121.060 88.385 121.320 89.535 ;
        RECT 121.495 88.460 121.750 89.365 ;
        RECT 121.920 88.775 122.250 89.535 ;
        RECT 122.465 88.605 122.635 89.365 ;
        RECT 118.845 87.535 119.560 87.705 ;
        RECT 118.845 87.155 119.015 87.535 ;
        RECT 119.230 86.985 119.560 87.365 ;
        RECT 119.730 87.155 119.985 87.730 ;
        RECT 120.160 86.985 120.420 87.825 ;
        RECT 121.060 86.985 121.320 87.825 ;
        RECT 121.495 87.730 121.665 88.460 ;
        RECT 121.920 88.435 122.635 88.605 ;
        RECT 122.895 88.445 124.105 89.535 ;
        RECT 121.920 88.225 122.090 88.435 ;
        RECT 121.835 87.895 122.090 88.225 ;
        RECT 121.495 87.155 121.750 87.730 ;
        RECT 121.920 87.705 122.090 87.895 ;
        RECT 122.370 87.885 122.725 88.255 ;
        RECT 122.895 87.735 123.415 88.275 ;
        RECT 123.585 87.905 124.105 88.445 ;
        RECT 124.365 88.605 124.535 89.365 ;
        RECT 124.750 88.775 125.080 89.535 ;
        RECT 124.365 88.435 125.080 88.605 ;
        RECT 125.250 88.460 125.505 89.365 ;
        RECT 124.275 87.885 124.630 88.255 ;
        RECT 124.910 88.225 125.080 88.435 ;
        RECT 124.910 87.895 125.165 88.225 ;
        RECT 121.920 87.535 122.635 87.705 ;
        RECT 121.920 86.985 122.250 87.365 ;
        RECT 122.465 87.155 122.635 87.535 ;
        RECT 122.895 86.985 124.105 87.735 ;
        RECT 124.910 87.705 125.080 87.895 ;
        RECT 125.335 87.730 125.505 88.460 ;
        RECT 125.680 88.385 125.940 89.535 ;
        RECT 126.115 88.445 127.325 89.535 ;
        RECT 124.365 87.535 125.080 87.705 ;
        RECT 124.365 87.155 124.535 87.535 ;
        RECT 124.750 86.985 125.080 87.365 ;
        RECT 125.250 87.155 125.505 87.730 ;
        RECT 125.680 86.985 125.940 87.825 ;
        RECT 126.115 87.735 126.635 88.275 ;
        RECT 126.805 87.905 127.325 88.445 ;
        RECT 127.585 88.605 127.755 89.365 ;
        RECT 127.970 88.775 128.300 89.535 ;
        RECT 127.585 88.435 128.300 88.605 ;
        RECT 128.470 88.460 128.725 89.365 ;
        RECT 127.495 87.885 127.850 88.255 ;
        RECT 128.130 88.225 128.300 88.435 ;
        RECT 128.130 87.895 128.385 88.225 ;
        RECT 126.115 86.985 127.325 87.735 ;
        RECT 128.130 87.705 128.300 87.895 ;
        RECT 128.555 87.730 128.725 88.460 ;
        RECT 128.900 88.385 129.160 89.535 ;
        RECT 129.335 88.370 129.625 89.535 ;
        RECT 130.720 88.385 130.980 89.535 ;
        RECT 131.155 88.460 131.410 89.365 ;
        RECT 131.580 88.775 131.910 89.535 ;
        RECT 132.125 88.605 132.295 89.365 ;
        RECT 127.585 87.535 128.300 87.705 ;
        RECT 127.585 87.155 127.755 87.535 ;
        RECT 127.970 86.985 128.300 87.365 ;
        RECT 128.470 87.155 128.725 87.730 ;
        RECT 128.900 86.985 129.160 87.825 ;
        RECT 129.335 86.985 129.625 87.710 ;
        RECT 130.720 86.985 130.980 87.825 ;
        RECT 131.155 87.730 131.325 88.460 ;
        RECT 131.580 88.435 132.295 88.605 ;
        RECT 132.555 88.445 136.065 89.535 ;
        RECT 136.235 88.445 137.445 89.535 ;
        RECT 131.580 88.225 131.750 88.435 ;
        RECT 131.495 87.895 131.750 88.225 ;
        RECT 131.155 87.155 131.410 87.730 ;
        RECT 131.580 87.705 131.750 87.895 ;
        RECT 132.030 87.885 132.385 88.255 ;
        RECT 132.555 87.755 134.205 88.275 ;
        RECT 134.375 87.925 136.065 88.445 ;
        RECT 131.580 87.535 132.295 87.705 ;
        RECT 131.580 86.985 131.910 87.365 ;
        RECT 132.125 87.155 132.295 87.535 ;
        RECT 132.555 86.985 136.065 87.755 ;
        RECT 136.235 87.735 136.755 88.275 ;
        RECT 136.925 87.905 137.445 88.445 ;
        RECT 137.615 88.445 138.825 89.535 ;
        RECT 137.615 87.905 138.135 88.445 ;
        RECT 138.305 87.735 138.825 88.275 ;
        RECT 136.235 86.985 137.445 87.735 ;
        RECT 137.615 86.985 138.825 87.735 ;
        RECT 13.330 86.815 138.910 86.985 ;
        RECT 12.920 51.555 48.800 51.725 ;
        RECT 13.005 50.465 14.215 51.555 ;
        RECT 14.385 51.120 19.730 51.555 ;
        RECT 13.005 49.755 13.525 50.295 ;
        RECT 13.695 49.925 14.215 50.465 ;
        RECT 13.005 49.005 14.215 49.755 ;
        RECT 15.970 49.550 16.310 50.380 ;
        RECT 17.790 49.870 18.140 51.120 ;
        RECT 20.915 50.625 21.085 51.385 ;
        RECT 21.300 50.795 21.630 51.555 ;
        RECT 20.915 50.455 21.630 50.625 ;
        RECT 21.800 50.480 22.055 51.385 ;
        RECT 20.825 49.905 21.180 50.275 ;
        RECT 21.460 50.245 21.630 50.455 ;
        RECT 21.460 49.915 21.715 50.245 ;
        RECT 21.460 49.725 21.630 49.915 ;
        RECT 21.885 49.750 22.055 50.480 ;
        RECT 22.230 50.405 22.490 51.555 ;
        RECT 22.675 50.755 23.005 51.555 ;
        RECT 23.185 51.215 24.615 51.385 ;
        RECT 23.185 50.585 23.435 51.215 ;
        RECT 22.665 50.415 23.435 50.585 ;
        RECT 20.915 49.555 21.630 49.725 ;
        RECT 14.385 49.005 19.730 49.550 ;
        RECT 20.915 49.175 21.085 49.555 ;
        RECT 21.300 49.005 21.630 49.385 ;
        RECT 21.800 49.175 22.055 49.750 ;
        RECT 22.230 49.005 22.490 49.845 ;
        RECT 22.665 49.745 22.835 50.415 ;
        RECT 23.005 49.915 23.410 50.245 ;
        RECT 23.625 49.915 23.875 51.045 ;
        RECT 24.075 50.245 24.275 51.045 ;
        RECT 24.445 50.535 24.615 51.215 ;
        RECT 24.785 50.705 25.100 51.555 ;
        RECT 25.275 50.755 25.715 51.385 ;
        RECT 24.445 50.365 25.235 50.535 ;
        RECT 24.075 49.915 24.320 50.245 ;
        RECT 24.505 49.915 24.895 50.195 ;
        RECT 25.065 49.915 25.235 50.365 ;
        RECT 25.405 49.745 25.715 50.755 ;
        RECT 25.885 50.390 26.175 51.555 ;
        RECT 27.380 50.925 27.665 51.385 ;
        RECT 27.835 51.095 28.105 51.555 ;
        RECT 27.380 50.705 28.335 50.925 ;
        RECT 27.265 49.975 27.955 50.535 ;
        RECT 28.125 49.805 28.335 50.705 ;
        RECT 22.665 49.175 23.155 49.745 ;
        RECT 23.325 49.575 24.485 49.745 ;
        RECT 23.325 49.175 23.555 49.575 ;
        RECT 23.725 49.005 24.145 49.405 ;
        RECT 24.315 49.175 24.485 49.575 ;
        RECT 24.655 49.005 25.105 49.745 ;
        RECT 25.275 49.185 25.715 49.745 ;
        RECT 25.885 49.005 26.175 49.730 ;
        RECT 27.380 49.635 28.335 49.805 ;
        RECT 28.505 50.535 28.905 51.385 ;
        RECT 29.095 50.925 29.375 51.385 ;
        RECT 29.895 51.095 30.220 51.555 ;
        RECT 29.095 50.705 30.220 50.925 ;
        RECT 28.505 49.975 29.600 50.535 ;
        RECT 29.770 50.245 30.220 50.705 ;
        RECT 30.390 50.415 30.775 51.385 ;
        RECT 27.380 49.175 27.665 49.635 ;
        RECT 27.835 49.005 28.105 49.465 ;
        RECT 28.505 49.175 28.905 49.975 ;
        RECT 29.770 49.915 30.325 50.245 ;
        RECT 29.770 49.805 30.220 49.915 ;
        RECT 29.095 49.635 30.220 49.805 ;
        RECT 30.495 49.745 30.775 50.415 ;
        RECT 31.870 50.405 32.130 51.555 ;
        RECT 32.305 50.480 32.560 51.385 ;
        RECT 32.730 50.795 33.060 51.555 ;
        RECT 33.275 50.625 33.445 51.385 ;
        RECT 33.820 50.925 34.105 51.385 ;
        RECT 34.275 51.095 34.545 51.555 ;
        RECT 33.820 50.705 34.775 50.925 ;
        RECT 29.095 49.175 29.375 49.635 ;
        RECT 29.895 49.005 30.220 49.465 ;
        RECT 30.390 49.175 30.775 49.745 ;
        RECT 31.870 49.005 32.130 49.845 ;
        RECT 32.305 49.750 32.475 50.480 ;
        RECT 32.730 50.455 33.445 50.625 ;
        RECT 32.730 50.245 32.900 50.455 ;
        RECT 32.645 49.915 32.900 50.245 ;
        RECT 32.305 49.175 32.560 49.750 ;
        RECT 32.730 49.725 32.900 49.915 ;
        RECT 33.180 49.905 33.535 50.275 ;
        RECT 33.705 49.975 34.395 50.535 ;
        RECT 34.565 49.805 34.775 50.705 ;
        RECT 32.730 49.555 33.445 49.725 ;
        RECT 32.730 49.005 33.060 49.385 ;
        RECT 33.275 49.175 33.445 49.555 ;
        RECT 33.820 49.635 34.775 49.805 ;
        RECT 34.945 50.535 35.345 51.385 ;
        RECT 35.535 50.925 35.815 51.385 ;
        RECT 36.335 51.095 36.660 51.555 ;
        RECT 35.535 50.705 36.660 50.925 ;
        RECT 34.945 49.975 36.040 50.535 ;
        RECT 36.210 50.245 36.660 50.705 ;
        RECT 36.830 50.415 37.215 51.385 ;
        RECT 37.465 50.625 37.645 51.385 ;
        RECT 37.825 50.795 38.155 51.555 ;
        RECT 37.465 50.455 38.140 50.625 ;
        RECT 38.325 50.480 38.595 51.385 ;
        RECT 33.820 49.175 34.105 49.635 ;
        RECT 34.275 49.005 34.545 49.465 ;
        RECT 34.945 49.175 35.345 49.975 ;
        RECT 36.210 49.915 36.765 50.245 ;
        RECT 36.210 49.805 36.660 49.915 ;
        RECT 35.535 49.635 36.660 49.805 ;
        RECT 36.935 49.745 37.215 50.415 ;
        RECT 37.970 50.310 38.140 50.455 ;
        RECT 37.405 49.905 37.745 50.275 ;
        RECT 37.970 49.980 38.245 50.310 ;
        RECT 35.535 49.175 35.815 49.635 ;
        RECT 36.335 49.005 36.660 49.465 ;
        RECT 36.830 49.175 37.215 49.745 ;
        RECT 37.970 49.725 38.140 49.980 ;
        RECT 37.475 49.555 38.140 49.725 ;
        RECT 38.415 49.680 38.595 50.480 ;
        RECT 38.765 50.390 39.055 51.555 ;
        RECT 40.150 50.405 40.410 51.555 ;
        RECT 40.585 50.480 40.840 51.385 ;
        RECT 41.010 50.795 41.340 51.555 ;
        RECT 41.555 50.625 41.725 51.385 ;
        RECT 37.475 49.175 37.645 49.555 ;
        RECT 37.825 49.005 38.155 49.385 ;
        RECT 38.335 49.175 38.595 49.680 ;
        RECT 38.765 49.005 39.055 49.730 ;
        RECT 40.150 49.005 40.410 49.845 ;
        RECT 40.585 49.750 40.755 50.480 ;
        RECT 41.010 50.455 41.725 50.625 ;
        RECT 41.985 50.465 43.195 51.555 ;
        RECT 41.010 50.245 41.180 50.455 ;
        RECT 40.925 49.915 41.180 50.245 ;
        RECT 40.585 49.175 40.840 49.750 ;
        RECT 41.010 49.725 41.180 49.915 ;
        RECT 41.460 49.905 41.815 50.275 ;
        RECT 41.985 49.755 42.505 50.295 ;
        RECT 42.675 49.925 43.195 50.465 ;
        RECT 43.365 50.480 43.635 51.385 ;
        RECT 43.805 50.795 44.135 51.555 ;
        RECT 44.315 50.625 44.485 51.385 ;
        RECT 41.010 49.555 41.725 49.725 ;
        RECT 41.010 49.005 41.340 49.385 ;
        RECT 41.555 49.175 41.725 49.555 ;
        RECT 41.985 49.005 43.195 49.755 ;
        RECT 43.365 49.680 43.535 50.480 ;
        RECT 43.820 50.455 44.485 50.625 ;
        RECT 44.745 50.480 45.015 51.385 ;
        RECT 45.185 50.795 45.515 51.555 ;
        RECT 45.695 50.625 45.865 51.385 ;
        RECT 43.820 50.310 43.990 50.455 ;
        RECT 43.705 49.980 43.990 50.310 ;
        RECT 43.820 49.725 43.990 49.980 ;
        RECT 44.225 49.905 44.555 50.275 ;
        RECT 43.365 49.175 43.625 49.680 ;
        RECT 43.820 49.555 44.485 49.725 ;
        RECT 43.805 49.005 44.135 49.385 ;
        RECT 44.315 49.175 44.485 49.555 ;
        RECT 44.745 49.680 44.915 50.480 ;
        RECT 45.200 50.455 45.865 50.625 ;
        RECT 46.125 50.480 46.395 51.385 ;
        RECT 46.565 50.795 46.895 51.555 ;
        RECT 47.075 50.625 47.255 51.385 ;
        RECT 45.200 50.310 45.370 50.455 ;
        RECT 45.085 49.980 45.370 50.310 ;
        RECT 45.200 49.725 45.370 49.980 ;
        RECT 45.605 49.905 45.935 50.275 ;
        RECT 44.745 49.175 45.005 49.680 ;
        RECT 45.200 49.555 45.865 49.725 ;
        RECT 45.185 49.005 45.515 49.385 ;
        RECT 45.695 49.175 45.865 49.555 ;
        RECT 46.125 49.680 46.305 50.480 ;
        RECT 46.580 50.455 47.255 50.625 ;
        RECT 47.505 50.465 48.715 51.555 ;
        RECT 46.580 50.310 46.750 50.455 ;
        RECT 46.475 49.980 46.750 50.310 ;
        RECT 46.580 49.725 46.750 49.980 ;
        RECT 46.975 49.905 47.315 50.275 ;
        RECT 47.505 49.925 48.025 50.465 ;
        RECT 48.195 49.755 48.715 50.295 ;
        RECT 46.125 49.175 46.385 49.680 ;
        RECT 46.580 49.555 47.245 49.725 ;
        RECT 46.565 49.005 46.895 49.385 ;
        RECT 47.075 49.175 47.245 49.555 ;
        RECT 47.505 49.005 48.715 49.755 ;
        RECT 12.920 48.835 48.800 49.005 ;
        RECT 13.005 48.085 14.215 48.835 ;
        RECT 13.005 47.545 13.525 48.085 ;
        RECT 14.385 48.065 17.895 48.835 ;
        RECT 18.575 48.180 18.905 48.615 ;
        RECT 19.075 48.225 19.245 48.835 ;
        RECT 18.525 48.095 18.905 48.180 ;
        RECT 19.415 48.095 19.745 48.620 ;
        RECT 20.005 48.305 20.215 48.835 ;
        RECT 20.490 48.385 21.275 48.555 ;
        RECT 21.445 48.385 21.850 48.555 ;
        RECT 13.695 47.375 14.215 47.915 ;
        RECT 14.385 47.545 16.035 48.065 ;
        RECT 18.525 48.055 18.750 48.095 ;
        RECT 16.205 47.375 17.895 47.895 ;
        RECT 13.005 46.285 14.215 47.375 ;
        RECT 14.385 46.285 17.895 47.375 ;
        RECT 18.525 47.475 18.695 48.055 ;
        RECT 19.415 47.925 19.615 48.095 ;
        RECT 20.490 47.925 20.660 48.385 ;
        RECT 18.865 47.595 19.615 47.925 ;
        RECT 19.785 47.595 20.660 47.925 ;
        RECT 18.525 47.425 18.740 47.475 ;
        RECT 18.525 47.345 18.915 47.425 ;
        RECT 18.585 46.500 18.915 47.345 ;
        RECT 19.425 47.390 19.615 47.595 ;
        RECT 19.085 46.285 19.255 47.295 ;
        RECT 19.425 47.015 20.320 47.390 ;
        RECT 19.425 46.455 19.765 47.015 ;
        RECT 19.995 46.285 20.310 46.785 ;
        RECT 20.490 46.755 20.660 47.595 ;
        RECT 20.830 47.885 21.295 48.215 ;
        RECT 21.680 48.155 21.850 48.385 ;
        RECT 22.030 48.335 22.400 48.835 ;
        RECT 22.720 48.385 23.395 48.555 ;
        RECT 23.590 48.385 23.925 48.555 ;
        RECT 20.830 46.925 21.150 47.885 ;
        RECT 21.680 47.855 22.510 48.155 ;
        RECT 21.320 46.955 21.510 47.675 ;
        RECT 21.680 46.785 21.850 47.855 ;
        RECT 22.310 47.825 22.510 47.855 ;
        RECT 22.020 47.605 22.190 47.675 ;
        RECT 22.720 47.605 22.890 48.385 ;
        RECT 23.755 48.245 23.925 48.385 ;
        RECT 24.095 48.375 24.345 48.835 ;
        RECT 22.020 47.435 22.890 47.605 ;
        RECT 23.060 47.965 23.585 48.185 ;
        RECT 23.755 48.115 23.980 48.245 ;
        RECT 22.020 47.345 22.530 47.435 ;
        RECT 20.490 46.585 21.375 46.755 ;
        RECT 21.600 46.455 21.850 46.785 ;
        RECT 22.020 46.285 22.190 47.085 ;
        RECT 22.360 46.730 22.530 47.345 ;
        RECT 23.060 47.265 23.230 47.965 ;
        RECT 22.700 46.900 23.230 47.265 ;
        RECT 23.400 47.200 23.640 47.795 ;
        RECT 23.810 47.010 23.980 48.115 ;
        RECT 24.150 47.255 24.430 48.205 ;
        RECT 23.675 46.880 23.980 47.010 ;
        RECT 22.360 46.560 23.465 46.730 ;
        RECT 23.675 46.455 23.925 46.880 ;
        RECT 24.095 46.285 24.360 46.745 ;
        RECT 24.600 46.455 24.785 48.575 ;
        RECT 24.955 48.455 25.285 48.835 ;
        RECT 25.455 48.285 25.625 48.575 ;
        RECT 24.960 48.115 25.625 48.285 ;
        RECT 25.975 48.285 26.145 48.575 ;
        RECT 26.315 48.455 26.645 48.835 ;
        RECT 25.975 48.115 26.640 48.285 ;
        RECT 24.960 47.125 25.190 48.115 ;
        RECT 25.360 47.295 25.710 47.945 ;
        RECT 25.890 47.295 26.240 47.945 ;
        RECT 26.410 47.125 26.640 48.115 ;
        RECT 24.960 46.955 25.625 47.125 ;
        RECT 24.955 46.285 25.285 46.785 ;
        RECT 25.455 46.455 25.625 46.955 ;
        RECT 25.975 46.955 26.640 47.125 ;
        RECT 25.975 46.455 26.145 46.955 ;
        RECT 26.315 46.285 26.645 46.785 ;
        RECT 26.815 46.455 27.000 48.575 ;
        RECT 27.255 48.375 27.505 48.835 ;
        RECT 27.675 48.385 28.010 48.555 ;
        RECT 28.205 48.385 28.880 48.555 ;
        RECT 27.675 48.245 27.845 48.385 ;
        RECT 27.170 47.255 27.450 48.205 ;
        RECT 27.620 48.115 27.845 48.245 ;
        RECT 27.620 47.010 27.790 48.115 ;
        RECT 28.015 47.965 28.540 48.185 ;
        RECT 27.960 47.200 28.200 47.795 ;
        RECT 28.370 47.265 28.540 47.965 ;
        RECT 28.710 47.605 28.880 48.385 ;
        RECT 29.200 48.335 29.570 48.835 ;
        RECT 29.750 48.385 30.155 48.555 ;
        RECT 30.325 48.385 31.110 48.555 ;
        RECT 29.750 48.155 29.920 48.385 ;
        RECT 29.090 47.855 29.920 48.155 ;
        RECT 30.305 47.885 30.770 48.215 ;
        RECT 29.090 47.825 29.290 47.855 ;
        RECT 29.410 47.605 29.580 47.675 ;
        RECT 28.710 47.435 29.580 47.605 ;
        RECT 29.070 47.345 29.580 47.435 ;
        RECT 27.620 46.880 27.925 47.010 ;
        RECT 28.370 46.900 28.900 47.265 ;
        RECT 27.240 46.285 27.505 46.745 ;
        RECT 27.675 46.455 27.925 46.880 ;
        RECT 29.070 46.730 29.240 47.345 ;
        RECT 28.135 46.560 29.240 46.730 ;
        RECT 29.410 46.285 29.580 47.085 ;
        RECT 29.750 46.785 29.920 47.855 ;
        RECT 30.090 46.955 30.280 47.675 ;
        RECT 30.450 46.925 30.770 47.885 ;
        RECT 30.940 47.925 31.110 48.385 ;
        RECT 31.385 48.305 31.595 48.835 ;
        RECT 31.855 48.095 32.185 48.620 ;
        RECT 32.355 48.225 32.525 48.835 ;
        RECT 32.695 48.180 33.025 48.615 ;
        RECT 32.695 48.095 33.075 48.180 ;
        RECT 31.985 47.925 32.185 48.095 ;
        RECT 32.850 48.055 33.075 48.095 ;
        RECT 30.940 47.595 31.815 47.925 ;
        RECT 31.985 47.595 32.735 47.925 ;
        RECT 29.750 46.455 30.000 46.785 ;
        RECT 30.940 46.755 31.110 47.595 ;
        RECT 31.985 47.390 32.175 47.595 ;
        RECT 32.905 47.475 33.075 48.055 ;
        RECT 32.860 47.425 33.075 47.475 ;
        RECT 31.280 47.015 32.175 47.390 ;
        RECT 32.685 47.345 33.075 47.425 ;
        RECT 33.280 48.095 33.895 48.665 ;
        RECT 34.065 48.325 34.280 48.835 ;
        RECT 34.510 48.325 34.790 48.655 ;
        RECT 34.970 48.325 35.210 48.835 ;
        RECT 30.225 46.585 31.110 46.755 ;
        RECT 31.290 46.285 31.605 46.785 ;
        RECT 31.835 46.455 32.175 47.015 ;
        RECT 32.345 46.285 32.515 47.295 ;
        RECT 32.685 46.500 33.015 47.345 ;
        RECT 33.280 47.075 33.595 48.095 ;
        RECT 33.765 47.425 33.935 47.925 ;
        RECT 34.185 47.595 34.450 48.155 ;
        RECT 34.620 47.425 34.790 48.325 ;
        RECT 35.635 48.285 35.805 48.665 ;
        RECT 36.020 48.455 36.350 48.835 ;
        RECT 34.960 47.595 35.315 48.155 ;
        RECT 35.635 48.115 36.350 48.285 ;
        RECT 35.545 47.565 35.900 47.935 ;
        RECT 36.180 47.925 36.350 48.115 ;
        RECT 36.520 48.090 36.775 48.665 ;
        RECT 36.180 47.595 36.435 47.925 ;
        RECT 33.765 47.255 35.190 47.425 ;
        RECT 36.180 47.385 36.350 47.595 ;
        RECT 33.280 46.455 33.815 47.075 ;
        RECT 33.985 46.285 34.315 47.085 ;
        RECT 34.800 47.080 35.190 47.255 ;
        RECT 35.635 47.215 36.350 47.385 ;
        RECT 36.605 47.360 36.775 48.090 ;
        RECT 36.950 47.995 37.210 48.835 ;
        RECT 37.425 48.015 37.655 48.835 ;
        RECT 37.825 48.035 38.155 48.665 ;
        RECT 37.405 47.595 37.735 47.845 ;
        RECT 37.905 47.435 38.155 48.035 ;
        RECT 38.325 48.015 38.535 48.835 ;
        RECT 38.765 48.110 39.055 48.835 ;
        RECT 39.225 48.095 39.665 48.655 ;
        RECT 39.835 48.095 40.285 48.835 ;
        RECT 40.455 48.265 40.625 48.665 ;
        RECT 40.795 48.435 41.215 48.835 ;
        RECT 41.385 48.265 41.615 48.665 ;
        RECT 40.455 48.095 41.615 48.265 ;
        RECT 41.785 48.095 42.275 48.665 ;
        RECT 35.635 46.455 35.805 47.215 ;
        RECT 36.020 46.285 36.350 47.045 ;
        RECT 36.520 46.455 36.775 47.360 ;
        RECT 36.950 46.285 37.210 47.435 ;
        RECT 37.425 46.285 37.655 47.425 ;
        RECT 37.825 46.455 38.155 47.435 ;
        RECT 38.325 46.285 38.535 47.425 ;
        RECT 38.765 46.285 39.055 47.450 ;
        RECT 39.225 47.085 39.535 48.095 ;
        RECT 39.705 47.475 39.875 47.925 ;
        RECT 40.045 47.645 40.435 47.925 ;
        RECT 40.620 47.595 40.865 47.925 ;
        RECT 39.705 47.305 40.495 47.475 ;
        RECT 39.225 46.455 39.665 47.085 ;
        RECT 39.840 46.285 40.155 47.135 ;
        RECT 40.325 46.625 40.495 47.305 ;
        RECT 40.665 46.795 40.865 47.595 ;
        RECT 41.065 46.795 41.315 47.925 ;
        RECT 41.530 47.595 41.935 47.925 ;
        RECT 42.105 47.425 42.275 48.095 ;
        RECT 42.560 48.205 42.845 48.665 ;
        RECT 43.015 48.375 43.285 48.835 ;
        RECT 42.560 48.035 43.515 48.205 ;
        RECT 41.505 47.255 42.275 47.425 ;
        RECT 42.445 47.305 43.135 47.865 ;
        RECT 41.505 46.625 41.755 47.255 ;
        RECT 43.305 47.135 43.515 48.035 ;
        RECT 40.325 46.455 41.755 46.625 ;
        RECT 41.935 46.285 42.265 47.085 ;
        RECT 42.560 46.915 43.515 47.135 ;
        RECT 43.685 47.865 44.085 48.665 ;
        RECT 44.275 48.205 44.555 48.665 ;
        RECT 45.075 48.375 45.400 48.835 ;
        RECT 44.275 48.035 45.400 48.205 ;
        RECT 45.570 48.095 45.955 48.665 ;
        RECT 44.950 47.925 45.400 48.035 ;
        RECT 43.685 47.305 44.780 47.865 ;
        RECT 44.950 47.595 45.505 47.925 ;
        RECT 42.560 46.455 42.845 46.915 ;
        RECT 43.015 46.285 43.285 46.745 ;
        RECT 43.685 46.455 44.085 47.305 ;
        RECT 44.950 47.135 45.400 47.595 ;
        RECT 45.675 47.425 45.955 48.095 ;
        RECT 44.275 46.915 45.400 47.135 ;
        RECT 44.275 46.455 44.555 46.915 ;
        RECT 45.075 46.285 45.400 46.745 ;
        RECT 45.570 46.455 45.955 47.425 ;
        RECT 46.125 48.160 46.385 48.665 ;
        RECT 46.565 48.455 46.895 48.835 ;
        RECT 47.075 48.285 47.245 48.665 ;
        RECT 46.125 47.360 46.305 48.160 ;
        RECT 46.580 48.115 47.245 48.285 ;
        RECT 46.580 47.860 46.750 48.115 ;
        RECT 47.505 48.085 48.715 48.835 ;
        RECT 46.475 47.530 46.750 47.860 ;
        RECT 46.975 47.565 47.315 47.935 ;
        RECT 46.580 47.385 46.750 47.530 ;
        RECT 46.125 46.455 46.395 47.360 ;
        RECT 46.580 47.215 47.255 47.385 ;
        RECT 46.565 46.285 46.895 47.045 ;
        RECT 47.075 46.455 47.255 47.215 ;
        RECT 47.505 47.375 48.025 47.915 ;
        RECT 48.195 47.545 48.715 48.085 ;
        RECT 47.505 46.285 48.715 47.375 ;
        RECT 12.920 46.115 48.800 46.285 ;
        RECT 13.005 45.025 14.215 46.115 ;
        RECT 14.475 45.445 14.645 45.945 ;
        RECT 14.815 45.615 15.145 46.115 ;
        RECT 14.475 45.275 15.140 45.445 ;
        RECT 13.005 44.315 13.525 44.855 ;
        RECT 13.695 44.485 14.215 45.025 ;
        RECT 14.390 44.455 14.740 45.105 ;
        RECT 13.005 43.565 14.215 44.315 ;
        RECT 14.910 44.285 15.140 45.275 ;
        RECT 14.475 44.115 15.140 44.285 ;
        RECT 14.475 43.825 14.645 44.115 ;
        RECT 14.815 43.565 15.145 43.945 ;
        RECT 15.315 43.825 15.500 45.945 ;
        RECT 15.740 45.655 16.005 46.115 ;
        RECT 16.175 45.520 16.425 45.945 ;
        RECT 16.635 45.670 17.740 45.840 ;
        RECT 16.120 45.390 16.425 45.520 ;
        RECT 15.670 44.195 15.950 45.145 ;
        RECT 16.120 44.285 16.290 45.390 ;
        RECT 16.460 44.605 16.700 45.200 ;
        RECT 16.870 45.135 17.400 45.500 ;
        RECT 16.870 44.435 17.040 45.135 ;
        RECT 17.570 45.055 17.740 45.670 ;
        RECT 17.910 45.315 18.080 46.115 ;
        RECT 18.250 45.615 18.500 45.945 ;
        RECT 18.725 45.645 19.610 45.815 ;
        RECT 17.570 44.965 18.080 45.055 ;
        RECT 16.120 44.155 16.345 44.285 ;
        RECT 16.515 44.215 17.040 44.435 ;
        RECT 17.210 44.795 18.080 44.965 ;
        RECT 15.755 43.565 16.005 44.025 ;
        RECT 16.175 44.015 16.345 44.155 ;
        RECT 17.210 44.015 17.380 44.795 ;
        RECT 17.910 44.725 18.080 44.795 ;
        RECT 17.590 44.545 17.790 44.575 ;
        RECT 18.250 44.545 18.420 45.615 ;
        RECT 18.590 44.725 18.780 45.445 ;
        RECT 17.590 44.245 18.420 44.545 ;
        RECT 18.950 44.515 19.270 45.475 ;
        RECT 16.175 43.845 16.510 44.015 ;
        RECT 16.705 43.845 17.380 44.015 ;
        RECT 17.700 43.565 18.070 44.065 ;
        RECT 18.250 44.015 18.420 44.245 ;
        RECT 18.805 44.185 19.270 44.515 ;
        RECT 19.440 44.805 19.610 45.645 ;
        RECT 19.790 45.615 20.105 46.115 ;
        RECT 20.335 45.385 20.675 45.945 ;
        RECT 19.780 45.010 20.675 45.385 ;
        RECT 20.845 45.105 21.015 46.115 ;
        RECT 20.485 44.805 20.675 45.010 ;
        RECT 21.185 45.055 21.515 45.900 ;
        RECT 21.185 44.975 21.575 45.055 ;
        RECT 21.360 44.925 21.575 44.975 ;
        RECT 19.440 44.475 20.315 44.805 ;
        RECT 20.485 44.475 21.235 44.805 ;
        RECT 19.440 44.015 19.610 44.475 ;
        RECT 20.485 44.305 20.685 44.475 ;
        RECT 21.405 44.345 21.575 44.925 ;
        RECT 21.350 44.305 21.575 44.345 ;
        RECT 18.250 43.845 18.655 44.015 ;
        RECT 18.825 43.845 19.610 44.015 ;
        RECT 19.885 43.565 20.095 44.095 ;
        RECT 20.355 43.780 20.685 44.305 ;
        RECT 21.195 44.220 21.575 44.305 ;
        RECT 21.745 44.975 22.130 45.945 ;
        RECT 22.300 45.655 22.625 46.115 ;
        RECT 23.145 45.485 23.425 45.945 ;
        RECT 22.300 45.265 23.425 45.485 ;
        RECT 21.745 44.305 22.025 44.975 ;
        RECT 22.300 44.805 22.750 45.265 ;
        RECT 23.615 45.095 24.015 45.945 ;
        RECT 24.415 45.655 24.685 46.115 ;
        RECT 24.855 45.485 25.140 45.945 ;
        RECT 22.195 44.475 22.750 44.805 ;
        RECT 22.920 44.535 24.015 45.095 ;
        RECT 22.300 44.365 22.750 44.475 ;
        RECT 20.855 43.565 21.025 44.175 ;
        RECT 21.195 43.785 21.525 44.220 ;
        RECT 21.745 43.735 22.130 44.305 ;
        RECT 22.300 44.195 23.425 44.365 ;
        RECT 22.300 43.565 22.625 44.025 ;
        RECT 23.145 43.735 23.425 44.195 ;
        RECT 23.615 43.735 24.015 44.535 ;
        RECT 24.185 45.265 25.140 45.485 ;
        RECT 24.185 44.365 24.395 45.265 ;
        RECT 24.565 44.535 25.255 45.095 ;
        RECT 25.885 44.950 26.175 46.115 ;
        RECT 26.350 44.975 26.685 45.945 ;
        RECT 26.855 44.975 27.025 46.115 ;
        RECT 27.195 45.775 29.225 45.945 ;
        RECT 24.185 44.195 25.140 44.365 ;
        RECT 26.350 44.305 26.520 44.975 ;
        RECT 27.195 44.805 27.365 45.775 ;
        RECT 26.690 44.475 26.945 44.805 ;
        RECT 27.170 44.475 27.365 44.805 ;
        RECT 27.535 45.435 28.660 45.605 ;
        RECT 26.775 44.305 26.945 44.475 ;
        RECT 27.535 44.305 27.705 45.435 ;
        RECT 24.415 43.565 24.685 44.025 ;
        RECT 24.855 43.735 25.140 44.195 ;
        RECT 25.885 43.565 26.175 44.290 ;
        RECT 26.350 43.735 26.605 44.305 ;
        RECT 26.775 44.135 27.705 44.305 ;
        RECT 27.875 45.095 28.885 45.265 ;
        RECT 27.875 44.295 28.045 45.095 ;
        RECT 28.250 44.755 28.525 44.895 ;
        RECT 28.245 44.585 28.525 44.755 ;
        RECT 27.530 44.100 27.705 44.135 ;
        RECT 26.775 43.565 27.105 43.965 ;
        RECT 27.530 43.735 28.060 44.100 ;
        RECT 28.250 43.735 28.525 44.585 ;
        RECT 28.695 43.735 28.885 45.095 ;
        RECT 29.055 45.110 29.225 45.775 ;
        RECT 29.395 45.355 29.565 46.115 ;
        RECT 29.800 45.355 30.315 45.765 ;
        RECT 29.055 44.920 29.805 45.110 ;
        RECT 29.975 44.545 30.315 45.355 ;
        RECT 31.130 45.145 31.520 45.320 ;
        RECT 32.005 45.315 32.335 46.115 ;
        RECT 32.505 45.325 33.040 45.945 ;
        RECT 31.130 44.975 32.555 45.145 ;
        RECT 29.085 44.375 30.315 44.545 ;
        RECT 29.065 43.565 29.575 44.100 ;
        RECT 29.795 43.770 30.040 44.375 ;
        RECT 31.005 44.245 31.360 44.805 ;
        RECT 31.530 44.075 31.700 44.975 ;
        RECT 31.870 44.245 32.135 44.805 ;
        RECT 32.385 44.475 32.555 44.975 ;
        RECT 32.725 44.305 33.040 45.325 ;
        RECT 33.305 44.975 33.515 46.115 ;
        RECT 33.685 44.965 34.015 45.945 ;
        RECT 34.185 44.975 34.415 46.115 ;
        RECT 34.715 45.445 34.885 45.945 ;
        RECT 35.055 45.615 35.385 46.115 ;
        RECT 34.715 45.275 35.380 45.445 ;
        RECT 31.110 43.565 31.350 44.075 ;
        RECT 31.530 43.745 31.810 44.075 ;
        RECT 32.040 43.565 32.255 44.075 ;
        RECT 32.425 43.735 33.040 44.305 ;
        RECT 33.305 43.565 33.515 44.385 ;
        RECT 33.685 44.365 33.935 44.965 ;
        RECT 34.105 44.555 34.435 44.805 ;
        RECT 34.630 44.455 34.980 45.105 ;
        RECT 33.685 43.735 34.015 44.365 ;
        RECT 34.185 43.565 34.415 44.385 ;
        RECT 35.150 44.285 35.380 45.275 ;
        RECT 34.715 44.115 35.380 44.285 ;
        RECT 34.715 43.825 34.885 44.115 ;
        RECT 35.055 43.565 35.385 43.945 ;
        RECT 35.555 43.825 35.740 45.945 ;
        RECT 35.980 45.655 36.245 46.115 ;
        RECT 36.415 45.520 36.665 45.945 ;
        RECT 36.875 45.670 37.980 45.840 ;
        RECT 36.360 45.390 36.665 45.520 ;
        RECT 35.910 44.195 36.190 45.145 ;
        RECT 36.360 44.285 36.530 45.390 ;
        RECT 36.700 44.605 36.940 45.200 ;
        RECT 37.110 45.135 37.640 45.500 ;
        RECT 37.110 44.435 37.280 45.135 ;
        RECT 37.810 45.055 37.980 45.670 ;
        RECT 38.150 45.315 38.320 46.115 ;
        RECT 38.490 45.615 38.740 45.945 ;
        RECT 38.965 45.645 39.850 45.815 ;
        RECT 37.810 44.965 38.320 45.055 ;
        RECT 36.360 44.155 36.585 44.285 ;
        RECT 36.755 44.215 37.280 44.435 ;
        RECT 37.450 44.795 38.320 44.965 ;
        RECT 35.995 43.565 36.245 44.025 ;
        RECT 36.415 44.015 36.585 44.155 ;
        RECT 37.450 44.015 37.620 44.795 ;
        RECT 38.150 44.725 38.320 44.795 ;
        RECT 37.830 44.545 38.030 44.575 ;
        RECT 38.490 44.545 38.660 45.615 ;
        RECT 38.830 44.725 39.020 45.445 ;
        RECT 37.830 44.245 38.660 44.545 ;
        RECT 39.190 44.515 39.510 45.475 ;
        RECT 36.415 43.845 36.750 44.015 ;
        RECT 36.945 43.845 37.620 44.015 ;
        RECT 37.940 43.565 38.310 44.065 ;
        RECT 38.490 44.015 38.660 44.245 ;
        RECT 39.045 44.185 39.510 44.515 ;
        RECT 39.680 44.805 39.850 45.645 ;
        RECT 40.030 45.615 40.345 46.115 ;
        RECT 40.575 45.385 40.915 45.945 ;
        RECT 40.020 45.010 40.915 45.385 ;
        RECT 41.085 45.105 41.255 46.115 ;
        RECT 40.725 44.805 40.915 45.010 ;
        RECT 41.425 45.055 41.755 45.900 ;
        RECT 42.630 45.145 43.020 45.320 ;
        RECT 43.505 45.315 43.835 46.115 ;
        RECT 44.005 45.325 44.540 45.945 ;
        RECT 41.425 44.975 41.815 45.055 ;
        RECT 42.630 44.975 44.055 45.145 ;
        RECT 41.600 44.925 41.815 44.975 ;
        RECT 39.680 44.475 40.555 44.805 ;
        RECT 40.725 44.475 41.475 44.805 ;
        RECT 39.680 44.015 39.850 44.475 ;
        RECT 40.725 44.305 40.925 44.475 ;
        RECT 41.645 44.345 41.815 44.925 ;
        RECT 41.590 44.305 41.815 44.345 ;
        RECT 38.490 43.845 38.895 44.015 ;
        RECT 39.065 43.845 39.850 44.015 ;
        RECT 40.125 43.565 40.335 44.095 ;
        RECT 40.595 43.780 40.925 44.305 ;
        RECT 41.435 44.220 41.815 44.305 ;
        RECT 42.505 44.245 42.860 44.805 ;
        RECT 41.095 43.565 41.265 44.175 ;
        RECT 41.435 43.785 41.765 44.220 ;
        RECT 43.030 44.075 43.200 44.975 ;
        RECT 43.370 44.245 43.635 44.805 ;
        RECT 43.885 44.475 44.055 44.975 ;
        RECT 44.225 44.305 44.540 45.325 ;
        RECT 44.835 45.185 45.005 45.945 ;
        RECT 45.185 45.355 45.515 46.115 ;
        RECT 44.835 45.015 45.500 45.185 ;
        RECT 45.685 45.040 45.955 45.945 ;
        RECT 45.330 44.870 45.500 45.015 ;
        RECT 44.765 44.465 45.095 44.835 ;
        RECT 45.330 44.540 45.615 44.870 ;
        RECT 42.610 43.565 42.850 44.075 ;
        RECT 43.030 43.745 43.310 44.075 ;
        RECT 43.540 43.565 43.755 44.075 ;
        RECT 43.925 43.735 44.540 44.305 ;
        RECT 45.330 44.285 45.500 44.540 ;
        RECT 44.835 44.115 45.500 44.285 ;
        RECT 45.785 44.240 45.955 45.040 ;
        RECT 44.835 43.735 45.005 44.115 ;
        RECT 45.185 43.565 45.515 43.945 ;
        RECT 45.695 43.735 45.955 44.240 ;
        RECT 46.125 45.040 46.395 45.945 ;
        RECT 46.565 45.355 46.895 46.115 ;
        RECT 47.075 45.185 47.255 45.945 ;
        RECT 46.125 44.240 46.305 45.040 ;
        RECT 46.580 45.015 47.255 45.185 ;
        RECT 47.505 45.025 48.715 46.115 ;
        RECT 46.580 44.870 46.750 45.015 ;
        RECT 46.475 44.540 46.750 44.870 ;
        RECT 46.580 44.285 46.750 44.540 ;
        RECT 46.975 44.465 47.315 44.835 ;
        RECT 47.505 44.485 48.025 45.025 ;
        RECT 48.195 44.315 48.715 44.855 ;
        RECT 46.125 43.735 46.385 44.240 ;
        RECT 46.580 44.115 47.245 44.285 ;
        RECT 46.565 43.565 46.895 43.945 ;
        RECT 47.075 43.735 47.245 44.115 ;
        RECT 47.505 43.565 48.715 44.315 ;
        RECT 12.920 43.395 48.800 43.565 ;
        RECT 13.005 42.645 14.215 43.395 ;
        RECT 13.005 42.105 13.525 42.645 ;
        RECT 14.390 42.555 14.650 43.395 ;
        RECT 14.825 42.650 15.080 43.225 ;
        RECT 15.250 43.015 15.580 43.395 ;
        RECT 15.795 42.845 15.965 43.225 ;
        RECT 15.250 42.675 15.965 42.845 ;
        RECT 13.695 41.935 14.215 42.475 ;
        RECT 13.005 40.845 14.215 41.935 ;
        RECT 14.390 40.845 14.650 41.995 ;
        RECT 14.825 41.920 14.995 42.650 ;
        RECT 15.250 42.485 15.420 42.675 ;
        RECT 16.230 42.655 16.485 43.225 ;
        RECT 16.655 42.995 16.985 43.395 ;
        RECT 17.410 42.860 17.940 43.225 ;
        RECT 18.130 43.055 18.405 43.225 ;
        RECT 18.125 42.885 18.405 43.055 ;
        RECT 17.410 42.825 17.585 42.860 ;
        RECT 16.655 42.655 17.585 42.825 ;
        RECT 15.165 42.155 15.420 42.485 ;
        RECT 15.250 41.945 15.420 42.155 ;
        RECT 15.700 42.125 16.055 42.495 ;
        RECT 16.230 41.985 16.400 42.655 ;
        RECT 16.655 42.485 16.825 42.655 ;
        RECT 16.570 42.155 16.825 42.485 ;
        RECT 17.050 42.155 17.245 42.485 ;
        RECT 14.825 41.015 15.080 41.920 ;
        RECT 15.250 41.775 15.965 41.945 ;
        RECT 15.250 40.845 15.580 41.605 ;
        RECT 15.795 41.015 15.965 41.775 ;
        RECT 16.230 41.015 16.565 41.985 ;
        RECT 16.735 40.845 16.905 41.985 ;
        RECT 17.075 41.185 17.245 42.155 ;
        RECT 17.415 41.525 17.585 42.655 ;
        RECT 17.755 41.865 17.925 42.665 ;
        RECT 18.130 42.065 18.405 42.885 ;
        RECT 18.575 41.865 18.765 43.225 ;
        RECT 18.945 42.860 19.455 43.395 ;
        RECT 19.675 42.585 19.920 43.190 ;
        RECT 20.365 42.645 21.575 43.395 ;
        RECT 21.835 42.915 22.135 43.395 ;
        RECT 22.305 42.745 22.565 43.200 ;
        RECT 22.735 42.915 22.995 43.395 ;
        RECT 23.175 42.745 23.435 43.200 ;
        RECT 23.605 42.915 23.855 43.395 ;
        RECT 24.035 42.745 24.295 43.200 ;
        RECT 24.465 42.915 24.715 43.395 ;
        RECT 24.895 42.745 25.155 43.200 ;
        RECT 25.325 42.915 25.570 43.395 ;
        RECT 25.740 42.745 26.015 43.200 ;
        RECT 26.185 42.915 26.430 43.395 ;
        RECT 26.600 42.745 26.860 43.200 ;
        RECT 27.030 42.915 27.290 43.395 ;
        RECT 27.460 42.745 27.720 43.200 ;
        RECT 27.890 42.915 28.150 43.395 ;
        RECT 28.320 42.745 28.580 43.200 ;
        RECT 28.750 42.835 29.010 43.395 ;
        RECT 18.965 42.415 20.195 42.585 ;
        RECT 17.755 41.695 18.765 41.865 ;
        RECT 18.935 41.850 19.685 42.040 ;
        RECT 17.415 41.355 18.540 41.525 ;
        RECT 18.935 41.185 19.105 41.850 ;
        RECT 19.855 41.605 20.195 42.415 ;
        RECT 20.365 42.105 20.885 42.645 ;
        RECT 21.835 42.575 28.580 42.745 ;
        RECT 21.055 41.935 21.575 42.475 ;
        RECT 17.075 41.015 19.105 41.185 ;
        RECT 19.275 40.845 19.445 41.605 ;
        RECT 19.680 41.195 20.195 41.605 ;
        RECT 20.365 40.845 21.575 41.935 ;
        RECT 21.835 41.985 23.000 42.575 ;
        RECT 29.180 42.405 29.430 43.215 ;
        RECT 29.610 42.870 29.870 43.395 ;
        RECT 30.040 42.405 30.290 43.215 ;
        RECT 30.470 42.885 30.775 43.395 ;
        RECT 23.170 42.155 30.290 42.405 ;
        RECT 30.460 42.155 30.775 42.715 ;
        RECT 30.945 42.655 31.330 43.225 ;
        RECT 31.500 42.935 31.825 43.395 ;
        RECT 32.345 42.765 32.625 43.225 ;
        RECT 21.835 41.760 28.580 41.985 ;
        RECT 21.835 40.845 22.105 41.590 ;
        RECT 22.275 41.020 22.565 41.760 ;
        RECT 23.175 41.745 28.580 41.760 ;
        RECT 22.735 40.850 22.990 41.575 ;
        RECT 23.175 41.020 23.435 41.745 ;
        RECT 23.605 40.850 23.850 41.575 ;
        RECT 24.035 41.020 24.295 41.745 ;
        RECT 24.465 40.850 24.710 41.575 ;
        RECT 24.895 41.020 25.155 41.745 ;
        RECT 25.325 40.850 25.570 41.575 ;
        RECT 25.740 41.020 26.000 41.745 ;
        RECT 26.170 40.850 26.430 41.575 ;
        RECT 26.600 41.020 26.860 41.745 ;
        RECT 27.030 40.850 27.290 41.575 ;
        RECT 27.460 41.020 27.720 41.745 ;
        RECT 27.890 40.850 28.150 41.575 ;
        RECT 28.320 41.020 28.580 41.745 ;
        RECT 28.750 40.850 29.010 41.645 ;
        RECT 29.180 41.020 29.430 42.155 ;
        RECT 22.735 40.845 29.010 40.850 ;
        RECT 29.610 40.845 29.870 41.655 ;
        RECT 30.045 41.015 30.290 42.155 ;
        RECT 30.945 41.985 31.225 42.655 ;
        RECT 31.500 42.595 32.625 42.765 ;
        RECT 31.500 42.485 31.950 42.595 ;
        RECT 31.395 42.155 31.950 42.485 ;
        RECT 32.815 42.425 33.215 43.225 ;
        RECT 33.615 42.935 33.885 43.395 ;
        RECT 34.055 42.765 34.340 43.225 ;
        RECT 30.470 40.845 30.765 41.655 ;
        RECT 30.945 41.015 31.330 41.985 ;
        RECT 31.500 41.695 31.950 42.155 ;
        RECT 32.120 41.865 33.215 42.425 ;
        RECT 31.500 41.475 32.625 41.695 ;
        RECT 31.500 40.845 31.825 41.305 ;
        RECT 32.345 41.015 32.625 41.475 ;
        RECT 32.815 41.015 33.215 41.865 ;
        RECT 33.385 42.595 34.340 42.765 ;
        RECT 34.625 42.645 35.835 43.395 ;
        RECT 36.015 42.895 36.345 43.395 ;
        RECT 36.545 42.825 36.715 43.175 ;
        RECT 36.915 42.995 37.245 43.395 ;
        RECT 37.415 42.825 37.585 43.175 ;
        RECT 37.755 42.995 38.135 43.395 ;
        RECT 33.385 41.695 33.595 42.595 ;
        RECT 33.765 41.865 34.455 42.425 ;
        RECT 34.625 42.105 35.145 42.645 ;
        RECT 35.315 41.935 35.835 42.475 ;
        RECT 36.010 42.155 36.360 42.725 ;
        RECT 36.545 42.655 38.155 42.825 ;
        RECT 38.325 42.720 38.595 43.065 ;
        RECT 37.985 42.485 38.155 42.655 ;
        RECT 33.385 41.475 34.340 41.695 ;
        RECT 33.615 40.845 33.885 41.305 ;
        RECT 34.055 41.015 34.340 41.475 ;
        RECT 34.625 40.845 35.835 41.935 ;
        RECT 36.010 41.695 36.330 41.985 ;
        RECT 36.530 41.865 37.240 42.485 ;
        RECT 37.410 42.155 37.815 42.485 ;
        RECT 37.985 42.155 38.255 42.485 ;
        RECT 37.985 41.985 38.155 42.155 ;
        RECT 38.425 41.985 38.595 42.720 ;
        RECT 38.765 42.670 39.055 43.395 ;
        RECT 39.225 42.655 39.585 43.030 ;
        RECT 39.850 42.655 40.020 43.395 ;
        RECT 40.300 42.825 40.470 43.030 ;
        RECT 40.300 42.655 40.840 42.825 ;
        RECT 37.430 41.815 38.155 41.985 ;
        RECT 37.430 41.695 37.600 41.815 ;
        RECT 36.010 41.525 37.600 41.695 ;
        RECT 36.010 41.065 37.665 41.355 ;
        RECT 37.835 40.845 38.115 41.645 ;
        RECT 38.325 41.015 38.595 41.985 ;
        RECT 38.765 40.845 39.055 42.010 ;
        RECT 39.225 42.000 39.480 42.655 ;
        RECT 39.650 42.155 40.000 42.485 ;
        RECT 40.170 42.155 40.500 42.485 ;
        RECT 39.225 41.015 39.565 42.000 ;
        RECT 39.735 41.615 40.000 42.155 ;
        RECT 40.670 41.955 40.840 42.655 ;
        RECT 40.215 41.785 40.840 41.955 ;
        RECT 41.010 42.025 41.180 43.225 ;
        RECT 41.410 42.745 41.740 43.225 ;
        RECT 41.910 42.925 42.080 43.395 ;
        RECT 42.250 42.745 42.580 43.210 ;
        RECT 41.410 42.575 42.580 42.745 ;
        RECT 42.905 42.655 43.265 43.030 ;
        RECT 43.530 42.655 43.700 43.395 ;
        RECT 43.980 42.825 44.150 43.030 ;
        RECT 43.980 42.655 44.520 42.825 ;
        RECT 41.350 42.195 41.920 42.405 ;
        RECT 42.090 42.195 42.735 42.405 ;
        RECT 41.010 41.615 41.715 42.025 ;
        RECT 42.905 42.000 43.160 42.655 ;
        RECT 43.330 42.155 43.680 42.485 ;
        RECT 43.850 42.155 44.180 42.485 ;
        RECT 39.735 41.445 41.715 41.615 ;
        RECT 39.735 40.845 40.145 41.275 ;
        RECT 40.890 40.845 41.220 41.265 ;
        RECT 41.390 41.015 41.715 41.445 ;
        RECT 42.190 40.845 42.520 41.945 ;
        RECT 42.905 41.015 43.245 42.000 ;
        RECT 43.415 41.615 43.680 42.155 ;
        RECT 44.350 41.955 44.520 42.655 ;
        RECT 43.895 41.785 44.520 41.955 ;
        RECT 44.690 42.025 44.860 43.225 ;
        RECT 45.090 42.745 45.420 43.225 ;
        RECT 45.590 42.925 45.760 43.395 ;
        RECT 45.930 42.745 46.260 43.210 ;
        RECT 45.090 42.575 46.260 42.745 ;
        RECT 47.505 42.645 48.715 43.395 ;
        RECT 45.030 42.195 45.600 42.405 ;
        RECT 45.770 42.195 46.415 42.405 ;
        RECT 44.690 41.615 45.395 42.025 ;
        RECT 43.415 41.445 45.395 41.615 ;
        RECT 43.415 40.845 43.825 41.275 ;
        RECT 44.570 40.845 44.900 41.265 ;
        RECT 45.070 41.015 45.395 41.445 ;
        RECT 45.870 40.845 46.200 41.945 ;
        RECT 47.505 41.935 48.025 42.475 ;
        RECT 48.195 42.105 48.715 42.645 ;
        RECT 47.505 40.845 48.715 41.935 ;
        RECT 12.920 40.675 48.800 40.845 ;
        RECT 13.005 39.585 14.215 40.675 ;
        RECT 13.005 38.875 13.525 39.415 ;
        RECT 13.695 39.045 14.215 39.585 ;
        RECT 14.390 39.535 14.725 40.505 ;
        RECT 14.895 39.535 15.065 40.675 ;
        RECT 15.235 40.335 17.265 40.505 ;
        RECT 13.005 38.125 14.215 38.875 ;
        RECT 14.390 38.865 14.560 39.535 ;
        RECT 15.235 39.365 15.405 40.335 ;
        RECT 14.730 39.035 14.985 39.365 ;
        RECT 15.210 39.035 15.405 39.365 ;
        RECT 15.575 39.995 16.700 40.165 ;
        RECT 14.815 38.865 14.985 39.035 ;
        RECT 15.575 38.865 15.745 39.995 ;
        RECT 14.390 38.295 14.645 38.865 ;
        RECT 14.815 38.695 15.745 38.865 ;
        RECT 15.915 39.655 16.925 39.825 ;
        RECT 15.915 38.855 16.085 39.655 ;
        RECT 15.570 38.660 15.745 38.695 ;
        RECT 14.815 38.125 15.145 38.525 ;
        RECT 15.570 38.295 16.100 38.660 ;
        RECT 16.290 38.635 16.565 39.455 ;
        RECT 16.285 38.465 16.565 38.635 ;
        RECT 16.290 38.295 16.565 38.465 ;
        RECT 16.735 38.295 16.925 39.655 ;
        RECT 17.095 39.670 17.265 40.335 ;
        RECT 17.435 39.915 17.605 40.675 ;
        RECT 17.840 39.915 18.355 40.325 ;
        RECT 17.095 39.480 17.845 39.670 ;
        RECT 18.015 39.105 18.355 39.915 ;
        RECT 18.615 40.005 18.785 40.505 ;
        RECT 18.955 40.175 19.285 40.675 ;
        RECT 18.615 39.835 19.280 40.005 ;
        RECT 17.125 38.935 18.355 39.105 ;
        RECT 18.530 39.015 18.880 39.665 ;
        RECT 17.105 38.125 17.615 38.660 ;
        RECT 17.835 38.330 18.080 38.935 ;
        RECT 19.050 38.845 19.280 39.835 ;
        RECT 18.615 38.675 19.280 38.845 ;
        RECT 18.615 38.385 18.785 38.675 ;
        RECT 18.955 38.125 19.285 38.505 ;
        RECT 19.455 38.385 19.640 40.505 ;
        RECT 19.880 40.215 20.145 40.675 ;
        RECT 20.315 40.080 20.565 40.505 ;
        RECT 20.775 40.230 21.880 40.400 ;
        RECT 20.260 39.950 20.565 40.080 ;
        RECT 19.810 38.755 20.090 39.705 ;
        RECT 20.260 38.845 20.430 39.950 ;
        RECT 20.600 39.165 20.840 39.760 ;
        RECT 21.010 39.695 21.540 40.060 ;
        RECT 21.010 38.995 21.180 39.695 ;
        RECT 21.710 39.615 21.880 40.230 ;
        RECT 22.050 39.875 22.220 40.675 ;
        RECT 22.390 40.175 22.640 40.505 ;
        RECT 22.865 40.205 23.750 40.375 ;
        RECT 21.710 39.525 22.220 39.615 ;
        RECT 20.260 38.715 20.485 38.845 ;
        RECT 20.655 38.775 21.180 38.995 ;
        RECT 21.350 39.355 22.220 39.525 ;
        RECT 19.895 38.125 20.145 38.585 ;
        RECT 20.315 38.575 20.485 38.715 ;
        RECT 21.350 38.575 21.520 39.355 ;
        RECT 22.050 39.285 22.220 39.355 ;
        RECT 21.730 39.105 21.930 39.135 ;
        RECT 22.390 39.105 22.560 40.175 ;
        RECT 22.730 39.285 22.920 40.005 ;
        RECT 21.730 38.805 22.560 39.105 ;
        RECT 23.090 39.075 23.410 40.035 ;
        RECT 20.315 38.405 20.650 38.575 ;
        RECT 20.845 38.405 21.520 38.575 ;
        RECT 21.840 38.125 22.210 38.625 ;
        RECT 22.390 38.575 22.560 38.805 ;
        RECT 22.945 38.745 23.410 39.075 ;
        RECT 23.580 39.365 23.750 40.205 ;
        RECT 23.930 40.175 24.245 40.675 ;
        RECT 24.475 39.945 24.815 40.505 ;
        RECT 23.920 39.570 24.815 39.945 ;
        RECT 24.985 39.665 25.155 40.675 ;
        RECT 24.625 39.365 24.815 39.570 ;
        RECT 25.325 39.615 25.655 40.460 ;
        RECT 25.325 39.535 25.715 39.615 ;
        RECT 25.500 39.485 25.715 39.535 ;
        RECT 25.885 39.510 26.175 40.675 ;
        RECT 26.435 40.005 26.605 40.505 ;
        RECT 26.775 40.175 27.105 40.675 ;
        RECT 26.435 39.835 27.100 40.005 ;
        RECT 23.580 39.035 24.455 39.365 ;
        RECT 24.625 39.035 25.375 39.365 ;
        RECT 23.580 38.575 23.750 39.035 ;
        RECT 24.625 38.865 24.825 39.035 ;
        RECT 25.545 38.905 25.715 39.485 ;
        RECT 26.350 39.015 26.700 39.665 ;
        RECT 25.490 38.865 25.715 38.905 ;
        RECT 22.390 38.405 22.795 38.575 ;
        RECT 22.965 38.405 23.750 38.575 ;
        RECT 24.025 38.125 24.235 38.655 ;
        RECT 24.495 38.340 24.825 38.865 ;
        RECT 25.335 38.780 25.715 38.865 ;
        RECT 24.995 38.125 25.165 38.735 ;
        RECT 25.335 38.345 25.665 38.780 ;
        RECT 25.885 38.125 26.175 38.850 ;
        RECT 26.870 38.845 27.100 39.835 ;
        RECT 26.435 38.675 27.100 38.845 ;
        RECT 26.435 38.385 26.605 38.675 ;
        RECT 26.775 38.125 27.105 38.505 ;
        RECT 27.275 38.385 27.460 40.505 ;
        RECT 27.700 40.215 27.965 40.675 ;
        RECT 28.135 40.080 28.385 40.505 ;
        RECT 28.595 40.230 29.700 40.400 ;
        RECT 28.080 39.950 28.385 40.080 ;
        RECT 27.630 38.755 27.910 39.705 ;
        RECT 28.080 38.845 28.250 39.950 ;
        RECT 28.420 39.165 28.660 39.760 ;
        RECT 28.830 39.695 29.360 40.060 ;
        RECT 28.830 38.995 29.000 39.695 ;
        RECT 29.530 39.615 29.700 40.230 ;
        RECT 29.870 39.875 30.040 40.675 ;
        RECT 30.210 40.175 30.460 40.505 ;
        RECT 30.685 40.205 31.570 40.375 ;
        RECT 29.530 39.525 30.040 39.615 ;
        RECT 28.080 38.715 28.305 38.845 ;
        RECT 28.475 38.775 29.000 38.995 ;
        RECT 29.170 39.355 30.040 39.525 ;
        RECT 27.715 38.125 27.965 38.585 ;
        RECT 28.135 38.575 28.305 38.715 ;
        RECT 29.170 38.575 29.340 39.355 ;
        RECT 29.870 39.285 30.040 39.355 ;
        RECT 29.550 39.105 29.750 39.135 ;
        RECT 30.210 39.105 30.380 40.175 ;
        RECT 30.550 39.285 30.740 40.005 ;
        RECT 29.550 38.805 30.380 39.105 ;
        RECT 30.910 39.075 31.230 40.035 ;
        RECT 28.135 38.405 28.470 38.575 ;
        RECT 28.665 38.405 29.340 38.575 ;
        RECT 29.660 38.125 30.030 38.625 ;
        RECT 30.210 38.575 30.380 38.805 ;
        RECT 30.765 38.745 31.230 39.075 ;
        RECT 31.400 39.365 31.570 40.205 ;
        RECT 31.750 40.175 32.065 40.675 ;
        RECT 32.295 39.945 32.635 40.505 ;
        RECT 31.740 39.570 32.635 39.945 ;
        RECT 32.805 39.665 32.975 40.675 ;
        RECT 32.445 39.365 32.635 39.570 ;
        RECT 33.145 39.615 33.475 40.460 ;
        RECT 34.165 39.720 34.435 40.675 ;
        RECT 34.620 39.620 34.925 40.405 ;
        RECT 35.105 40.205 35.790 40.675 ;
        RECT 35.100 39.685 35.795 39.995 ;
        RECT 33.145 39.535 33.535 39.615 ;
        RECT 33.320 39.485 33.535 39.535 ;
        RECT 31.400 39.035 32.275 39.365 ;
        RECT 32.445 39.035 33.195 39.365 ;
        RECT 31.400 38.575 31.570 39.035 ;
        RECT 32.445 38.865 32.645 39.035 ;
        RECT 33.365 38.905 33.535 39.485 ;
        RECT 33.310 38.865 33.535 38.905 ;
        RECT 30.210 38.405 30.615 38.575 ;
        RECT 30.785 38.405 31.570 38.575 ;
        RECT 31.845 38.125 32.055 38.655 ;
        RECT 32.315 38.340 32.645 38.865 ;
        RECT 33.155 38.780 33.535 38.865 ;
        RECT 34.620 38.815 34.795 39.620 ;
        RECT 35.970 39.515 36.255 40.460 ;
        RECT 36.455 40.225 36.785 40.675 ;
        RECT 36.955 40.055 37.125 40.485 ;
        RECT 35.395 39.365 36.255 39.515 ;
        RECT 34.965 39.345 36.255 39.365 ;
        RECT 36.445 39.825 37.125 40.055 ;
        RECT 38.305 39.875 38.745 40.505 ;
        RECT 34.965 38.985 35.955 39.345 ;
        RECT 36.445 39.175 36.680 39.825 ;
        RECT 32.815 38.125 32.985 38.735 ;
        RECT 33.155 38.345 33.485 38.780 ;
        RECT 34.165 38.125 34.435 38.760 ;
        RECT 34.620 38.295 34.855 38.815 ;
        RECT 35.785 38.650 35.955 38.985 ;
        RECT 36.125 38.845 36.680 39.175 ;
        RECT 36.465 38.695 36.680 38.845 ;
        RECT 36.850 38.975 37.150 39.655 ;
        RECT 36.850 38.805 37.155 38.975 ;
        RECT 38.305 38.865 38.615 39.875 ;
        RECT 38.920 39.825 39.235 40.675 ;
        RECT 39.405 40.335 40.835 40.505 ;
        RECT 39.405 39.655 39.575 40.335 ;
        RECT 38.785 39.485 39.575 39.655 ;
        RECT 38.785 39.035 38.955 39.485 ;
        RECT 39.745 39.365 39.945 40.165 ;
        RECT 39.125 39.035 39.515 39.315 ;
        RECT 39.700 39.035 39.945 39.365 ;
        RECT 40.145 39.035 40.395 40.165 ;
        RECT 40.585 39.705 40.835 40.335 ;
        RECT 41.015 39.875 41.345 40.675 ;
        RECT 41.535 39.705 41.865 40.490 ;
        RECT 40.585 39.535 41.355 39.705 ;
        RECT 41.535 39.535 42.215 39.705 ;
        RECT 42.395 39.535 42.725 40.675 ;
        RECT 40.610 39.035 41.015 39.365 ;
        RECT 41.185 38.865 41.355 39.535 ;
        RECT 41.525 39.115 41.875 39.365 ;
        RECT 42.045 38.935 42.215 39.535 ;
        RECT 43.365 39.520 43.705 40.505 ;
        RECT 43.875 40.245 44.285 40.675 ;
        RECT 45.030 40.255 45.360 40.675 ;
        RECT 45.530 40.075 45.855 40.505 ;
        RECT 43.875 39.905 45.855 40.075 ;
        RECT 42.385 39.115 42.735 39.365 ;
        RECT 35.025 38.125 35.425 38.620 ;
        RECT 35.785 38.455 36.185 38.650 ;
        RECT 36.015 38.310 36.185 38.455 ;
        RECT 36.465 38.320 36.705 38.695 ;
        RECT 36.875 38.125 37.205 38.630 ;
        RECT 38.305 38.305 38.745 38.865 ;
        RECT 38.915 38.125 39.365 38.865 ;
        RECT 39.535 38.695 40.695 38.865 ;
        RECT 39.535 38.295 39.705 38.695 ;
        RECT 39.875 38.125 40.295 38.525 ;
        RECT 40.465 38.295 40.695 38.695 ;
        RECT 40.865 38.295 41.355 38.865 ;
        RECT 41.545 38.125 41.785 38.935 ;
        RECT 41.955 38.295 42.285 38.935 ;
        RECT 42.455 38.125 42.725 38.935 ;
        RECT 43.365 38.865 43.620 39.520 ;
        RECT 43.875 39.365 44.140 39.905 ;
        RECT 44.355 39.565 44.980 39.735 ;
        RECT 43.790 39.035 44.140 39.365 ;
        RECT 44.310 39.035 44.640 39.365 ;
        RECT 44.810 38.865 44.980 39.565 ;
        RECT 43.365 38.490 43.725 38.865 ;
        RECT 43.990 38.125 44.160 38.865 ;
        RECT 44.440 38.695 44.980 38.865 ;
        RECT 45.150 39.495 45.855 39.905 ;
        RECT 46.330 39.575 46.660 40.675 ;
        RECT 47.505 39.585 48.715 40.675 ;
        RECT 44.440 38.490 44.610 38.695 ;
        RECT 45.150 38.295 45.320 39.495 ;
        RECT 45.490 39.115 46.060 39.325 ;
        RECT 46.230 39.115 46.875 39.325 ;
        RECT 47.505 39.045 48.025 39.585 ;
        RECT 45.550 38.775 46.720 38.945 ;
        RECT 48.195 38.875 48.715 39.415 ;
        RECT 45.550 38.295 45.880 38.775 ;
        RECT 46.050 38.125 46.220 38.595 ;
        RECT 46.390 38.310 46.720 38.775 ;
        RECT 47.505 38.125 48.715 38.875 ;
        RECT 12.920 37.955 48.800 38.125 ;
        RECT 13.005 37.205 14.215 37.955 ;
        RECT 14.435 37.300 14.765 37.735 ;
        RECT 14.935 37.345 15.105 37.955 ;
        RECT 14.385 37.215 14.765 37.300 ;
        RECT 15.275 37.215 15.605 37.740 ;
        RECT 15.865 37.425 16.075 37.955 ;
        RECT 16.350 37.505 17.135 37.675 ;
        RECT 17.305 37.505 17.710 37.675 ;
        RECT 13.005 36.665 13.525 37.205 ;
        RECT 14.385 37.175 14.610 37.215 ;
        RECT 13.695 36.495 14.215 37.035 ;
        RECT 13.005 35.405 14.215 36.495 ;
        RECT 14.385 36.595 14.555 37.175 ;
        RECT 15.275 37.045 15.475 37.215 ;
        RECT 16.350 37.045 16.520 37.505 ;
        RECT 14.725 36.715 15.475 37.045 ;
        RECT 15.645 36.715 16.520 37.045 ;
        RECT 14.385 36.545 14.600 36.595 ;
        RECT 14.385 36.465 14.775 36.545 ;
        RECT 14.445 35.620 14.775 36.465 ;
        RECT 15.285 36.510 15.475 36.715 ;
        RECT 14.945 35.405 15.115 36.415 ;
        RECT 15.285 36.135 16.180 36.510 ;
        RECT 15.285 35.575 15.625 36.135 ;
        RECT 15.855 35.405 16.170 35.905 ;
        RECT 16.350 35.875 16.520 36.715 ;
        RECT 16.690 37.005 17.155 37.335 ;
        RECT 17.540 37.275 17.710 37.505 ;
        RECT 17.890 37.455 18.260 37.955 ;
        RECT 18.580 37.505 19.255 37.675 ;
        RECT 19.450 37.505 19.785 37.675 ;
        RECT 16.690 36.045 17.010 37.005 ;
        RECT 17.540 36.975 18.370 37.275 ;
        RECT 17.180 36.075 17.370 36.795 ;
        RECT 17.540 35.905 17.710 36.975 ;
        RECT 18.170 36.945 18.370 36.975 ;
        RECT 17.880 36.725 18.050 36.795 ;
        RECT 18.580 36.725 18.750 37.505 ;
        RECT 19.615 37.365 19.785 37.505 ;
        RECT 19.955 37.495 20.205 37.955 ;
        RECT 17.880 36.555 18.750 36.725 ;
        RECT 18.920 37.085 19.445 37.305 ;
        RECT 19.615 37.235 19.840 37.365 ;
        RECT 17.880 36.465 18.390 36.555 ;
        RECT 16.350 35.705 17.235 35.875 ;
        RECT 17.460 35.575 17.710 35.905 ;
        RECT 17.880 35.405 18.050 36.205 ;
        RECT 18.220 35.850 18.390 36.465 ;
        RECT 18.920 36.385 19.090 37.085 ;
        RECT 18.560 36.020 19.090 36.385 ;
        RECT 19.260 36.320 19.500 36.915 ;
        RECT 19.670 36.130 19.840 37.235 ;
        RECT 20.010 36.375 20.290 37.325 ;
        RECT 19.535 36.000 19.840 36.130 ;
        RECT 18.220 35.680 19.325 35.850 ;
        RECT 19.535 35.575 19.785 36.000 ;
        RECT 19.955 35.405 20.220 35.865 ;
        RECT 20.460 35.575 20.645 37.695 ;
        RECT 20.815 37.575 21.145 37.955 ;
        RECT 21.315 37.405 21.485 37.695 ;
        RECT 20.820 37.235 21.485 37.405 ;
        RECT 20.820 36.245 21.050 37.235 ;
        RECT 21.745 37.185 24.335 37.955 ;
        RECT 24.965 37.445 25.270 37.955 ;
        RECT 21.220 36.415 21.570 37.065 ;
        RECT 21.745 36.665 22.955 37.185 ;
        RECT 23.125 36.495 24.335 37.015 ;
        RECT 24.965 36.715 25.280 37.275 ;
        RECT 25.450 36.965 25.700 37.775 ;
        RECT 25.870 37.430 26.130 37.955 ;
        RECT 26.310 36.965 26.560 37.775 ;
        RECT 26.730 37.395 26.990 37.955 ;
        RECT 27.160 37.305 27.420 37.760 ;
        RECT 27.590 37.475 27.850 37.955 ;
        RECT 28.020 37.305 28.280 37.760 ;
        RECT 28.450 37.475 28.710 37.955 ;
        RECT 28.880 37.305 29.140 37.760 ;
        RECT 29.310 37.475 29.555 37.955 ;
        RECT 29.725 37.305 30.000 37.760 ;
        RECT 30.170 37.475 30.415 37.955 ;
        RECT 30.585 37.305 30.845 37.760 ;
        RECT 31.025 37.475 31.275 37.955 ;
        RECT 31.445 37.305 31.705 37.760 ;
        RECT 31.885 37.475 32.135 37.955 ;
        RECT 32.305 37.305 32.565 37.760 ;
        RECT 32.745 37.475 33.005 37.955 ;
        RECT 33.175 37.305 33.435 37.760 ;
        RECT 33.605 37.475 33.905 37.955 ;
        RECT 27.160 37.135 33.905 37.305 ;
        RECT 25.450 36.715 32.570 36.965 ;
        RECT 20.820 36.075 21.485 36.245 ;
        RECT 20.815 35.405 21.145 35.905 ;
        RECT 21.315 35.575 21.485 36.075 ;
        RECT 21.745 35.405 24.335 36.495 ;
        RECT 24.975 35.405 25.270 36.215 ;
        RECT 25.450 35.575 25.695 36.715 ;
        RECT 25.870 35.405 26.130 36.215 ;
        RECT 26.310 35.580 26.560 36.715 ;
        RECT 32.740 36.545 33.905 37.135 ;
        RECT 27.160 36.320 33.905 36.545 ;
        RECT 34.165 37.215 34.550 37.785 ;
        RECT 34.720 37.495 35.045 37.955 ;
        RECT 35.565 37.325 35.845 37.785 ;
        RECT 34.165 36.545 34.445 37.215 ;
        RECT 34.720 37.155 35.845 37.325 ;
        RECT 34.720 37.045 35.170 37.155 ;
        RECT 34.615 36.715 35.170 37.045 ;
        RECT 36.035 36.985 36.435 37.785 ;
        RECT 36.835 37.495 37.105 37.955 ;
        RECT 37.275 37.325 37.560 37.785 ;
        RECT 27.160 36.305 32.565 36.320 ;
        RECT 26.730 35.410 26.990 36.205 ;
        RECT 27.160 35.580 27.420 36.305 ;
        RECT 27.590 35.410 27.850 36.135 ;
        RECT 28.020 35.580 28.280 36.305 ;
        RECT 28.450 35.410 28.710 36.135 ;
        RECT 28.880 35.580 29.140 36.305 ;
        RECT 29.310 35.410 29.570 36.135 ;
        RECT 29.740 35.580 30.000 36.305 ;
        RECT 30.170 35.410 30.415 36.135 ;
        RECT 30.585 35.580 30.845 36.305 ;
        RECT 31.030 35.410 31.275 36.135 ;
        RECT 31.445 35.580 31.705 36.305 ;
        RECT 31.890 35.410 32.135 36.135 ;
        RECT 32.305 35.580 32.565 36.305 ;
        RECT 32.750 35.410 33.005 36.135 ;
        RECT 33.175 35.580 33.465 36.320 ;
        RECT 26.730 35.405 33.005 35.410 ;
        RECT 33.635 35.405 33.905 36.150 ;
        RECT 34.165 35.575 34.550 36.545 ;
        RECT 34.720 36.255 35.170 36.715 ;
        RECT 35.340 36.425 36.435 36.985 ;
        RECT 34.720 36.035 35.845 36.255 ;
        RECT 34.720 35.405 35.045 35.865 ;
        RECT 35.565 35.575 35.845 36.035 ;
        RECT 36.035 35.575 36.435 36.425 ;
        RECT 36.605 37.155 37.560 37.325 ;
        RECT 38.765 37.230 39.055 37.955 ;
        RECT 39.240 37.385 39.495 37.735 ;
        RECT 39.665 37.555 39.995 37.955 ;
        RECT 40.165 37.385 40.335 37.735 ;
        RECT 40.505 37.555 40.885 37.955 ;
        RECT 39.240 37.215 40.905 37.385 ;
        RECT 41.075 37.280 41.350 37.625 ;
        RECT 36.605 36.255 36.815 37.155 ;
        RECT 40.735 37.045 40.905 37.215 ;
        RECT 36.985 36.425 37.675 36.985 ;
        RECT 39.225 36.715 39.570 37.045 ;
        RECT 39.740 36.715 40.565 37.045 ;
        RECT 40.735 36.715 41.010 37.045 ;
        RECT 36.605 36.035 37.560 36.255 ;
        RECT 36.835 35.405 37.105 35.865 ;
        RECT 37.275 35.575 37.560 36.035 ;
        RECT 38.765 35.405 39.055 36.570 ;
        RECT 39.245 36.255 39.570 36.545 ;
        RECT 39.740 36.425 39.935 36.715 ;
        RECT 40.735 36.545 40.905 36.715 ;
        RECT 41.180 36.545 41.350 37.280 ;
        RECT 41.525 37.185 44.115 37.955 ;
        RECT 41.525 36.665 42.735 37.185 ;
        RECT 44.755 37.145 45.025 37.955 ;
        RECT 45.195 37.145 45.525 37.785 ;
        RECT 45.695 37.145 45.935 37.955 ;
        RECT 46.125 37.280 46.385 37.785 ;
        RECT 46.565 37.575 46.895 37.955 ;
        RECT 47.075 37.405 47.245 37.785 ;
        RECT 40.245 36.375 40.905 36.545 ;
        RECT 40.245 36.255 40.415 36.375 ;
        RECT 39.245 36.085 40.415 36.255 ;
        RECT 39.225 35.625 40.415 35.915 ;
        RECT 40.585 35.405 40.865 36.205 ;
        RECT 41.075 35.575 41.350 36.545 ;
        RECT 42.905 36.495 44.115 37.015 ;
        RECT 44.745 36.715 45.095 36.965 ;
        RECT 45.265 36.545 45.435 37.145 ;
        RECT 45.605 36.715 45.955 36.965 ;
        RECT 41.525 35.405 44.115 36.495 ;
        RECT 44.755 35.405 45.085 36.545 ;
        RECT 45.265 36.375 45.945 36.545 ;
        RECT 45.615 35.590 45.945 36.375 ;
        RECT 46.125 36.480 46.295 37.280 ;
        RECT 46.580 37.235 47.245 37.405 ;
        RECT 46.580 36.980 46.750 37.235 ;
        RECT 47.505 37.205 48.715 37.955 ;
        RECT 46.465 36.650 46.750 36.980 ;
        RECT 46.985 36.685 47.315 37.055 ;
        RECT 46.580 36.505 46.750 36.650 ;
        RECT 46.125 35.575 46.395 36.480 ;
        RECT 46.580 36.335 47.245 36.505 ;
        RECT 46.565 35.405 46.895 36.165 ;
        RECT 47.075 35.575 47.245 36.335 ;
        RECT 47.505 36.495 48.025 37.035 ;
        RECT 48.195 36.665 48.715 37.205 ;
        RECT 47.505 35.405 48.715 36.495 ;
        RECT 12.920 35.235 48.800 35.405 ;
        RECT 13.005 34.145 14.215 35.235 ;
        RECT 14.385 34.145 15.595 35.235 ;
        RECT 15.880 34.605 16.165 35.065 ;
        RECT 16.335 34.775 16.605 35.235 ;
        RECT 15.880 34.385 16.835 34.605 ;
        RECT 13.005 33.435 13.525 33.975 ;
        RECT 13.695 33.605 14.215 34.145 ;
        RECT 14.385 33.435 14.905 33.975 ;
        RECT 15.075 33.605 15.595 34.145 ;
        RECT 15.765 33.655 16.455 34.215 ;
        RECT 16.625 33.485 16.835 34.385 ;
        RECT 13.005 32.685 14.215 33.435 ;
        RECT 14.385 32.685 15.595 33.435 ;
        RECT 15.880 33.315 16.835 33.485 ;
        RECT 17.005 34.215 17.405 35.065 ;
        RECT 17.595 34.605 17.875 35.065 ;
        RECT 18.395 34.775 18.720 35.235 ;
        RECT 17.595 34.385 18.720 34.605 ;
        RECT 17.005 33.655 18.100 34.215 ;
        RECT 18.270 33.925 18.720 34.385 ;
        RECT 18.890 34.095 19.275 35.065 ;
        RECT 15.880 32.855 16.165 33.315 ;
        RECT 16.335 32.685 16.605 33.145 ;
        RECT 17.005 32.855 17.405 33.655 ;
        RECT 18.270 33.595 18.825 33.925 ;
        RECT 18.270 33.485 18.720 33.595 ;
        RECT 17.595 33.315 18.720 33.485 ;
        RECT 18.995 33.425 19.275 34.095 ;
        RECT 17.595 32.855 17.875 33.315 ;
        RECT 18.395 32.685 18.720 33.145 ;
        RECT 18.890 32.855 19.275 33.425 ;
        RECT 19.445 34.095 19.830 35.065 ;
        RECT 20.000 34.775 20.325 35.235 ;
        RECT 20.845 34.605 21.125 35.065 ;
        RECT 20.000 34.385 21.125 34.605 ;
        RECT 19.445 33.425 19.725 34.095 ;
        RECT 20.000 33.925 20.450 34.385 ;
        RECT 21.315 34.215 21.715 35.065 ;
        RECT 22.115 34.775 22.385 35.235 ;
        RECT 22.555 34.605 22.840 35.065 ;
        RECT 19.895 33.595 20.450 33.925 ;
        RECT 20.620 33.655 21.715 34.215 ;
        RECT 20.000 33.485 20.450 33.595 ;
        RECT 19.445 32.855 19.830 33.425 ;
        RECT 20.000 33.315 21.125 33.485 ;
        RECT 20.000 32.685 20.325 33.145 ;
        RECT 20.845 32.855 21.125 33.315 ;
        RECT 21.315 32.855 21.715 33.655 ;
        RECT 21.885 34.385 22.840 34.605 ;
        RECT 21.885 33.485 22.095 34.385 ;
        RECT 22.265 33.655 22.955 34.215 ;
        RECT 23.125 34.145 25.715 35.235 ;
        RECT 21.885 33.315 22.840 33.485 ;
        RECT 22.115 32.685 22.385 33.145 ;
        RECT 22.555 32.855 22.840 33.315 ;
        RECT 23.125 33.455 24.335 33.975 ;
        RECT 24.505 33.625 25.715 34.145 ;
        RECT 25.885 34.070 26.175 35.235 ;
        RECT 26.355 34.095 26.685 35.235 ;
        RECT 27.215 34.265 27.545 35.050 ;
        RECT 26.865 34.095 27.545 34.265 ;
        RECT 27.845 34.115 28.175 35.235 ;
        RECT 26.345 33.675 26.695 33.925 ;
        RECT 26.865 33.495 27.035 34.095 ;
        RECT 27.205 33.675 27.555 33.925 ;
        RECT 27.785 33.675 28.295 33.925 ;
        RECT 28.505 33.675 28.875 34.990 ;
        RECT 29.045 33.675 29.375 34.990 ;
        RECT 29.585 33.675 29.915 34.990 ;
        RECT 30.185 34.345 30.435 35.065 ;
        RECT 30.605 34.515 30.935 35.235 ;
        RECT 30.185 34.055 30.935 34.345 ;
        RECT 31.170 34.055 31.695 35.065 ;
        RECT 30.675 33.885 30.935 34.055 ;
        RECT 30.085 33.675 30.505 33.885 ;
        RECT 30.675 33.675 31.255 33.885 ;
        RECT 30.675 33.505 31.045 33.675 ;
        RECT 23.125 32.685 25.715 33.455 ;
        RECT 25.885 32.685 26.175 33.410 ;
        RECT 26.355 32.685 26.625 33.495 ;
        RECT 26.795 32.855 27.125 33.495 ;
        RECT 27.295 32.685 27.535 33.495 ;
        RECT 27.825 33.335 30.125 33.505 ;
        RECT 27.825 32.855 28.155 33.335 ;
        RECT 28.325 32.685 28.655 33.145 ;
        RECT 28.870 32.855 29.200 33.335 ;
        RECT 29.400 32.685 29.730 33.145 ;
        RECT 29.955 33.015 30.125 33.335 ;
        RECT 30.295 33.315 31.045 33.505 ;
        RECT 31.425 33.485 31.695 34.055 ;
        RECT 30.295 32.870 30.625 33.315 ;
        RECT 30.895 32.685 31.065 33.145 ;
        RECT 31.355 32.855 31.695 33.485 ;
        RECT 31.865 34.095 32.250 35.065 ;
        RECT 32.420 34.775 32.745 35.235 ;
        RECT 33.265 34.605 33.545 35.065 ;
        RECT 32.420 34.385 33.545 34.605 ;
        RECT 31.865 33.425 32.145 34.095 ;
        RECT 32.420 33.925 32.870 34.385 ;
        RECT 33.735 34.215 34.135 35.065 ;
        RECT 34.535 34.775 34.805 35.235 ;
        RECT 34.975 34.605 35.260 35.065 ;
        RECT 32.315 33.595 32.870 33.925 ;
        RECT 33.040 33.655 34.135 34.215 ;
        RECT 32.420 33.485 32.870 33.595 ;
        RECT 31.865 32.855 32.250 33.425 ;
        RECT 32.420 33.315 33.545 33.485 ;
        RECT 32.420 32.685 32.745 33.145 ;
        RECT 33.265 32.855 33.545 33.315 ;
        RECT 33.735 32.855 34.135 33.655 ;
        RECT 34.305 34.385 35.260 34.605 ;
        RECT 34.305 33.485 34.515 34.385 ;
        RECT 34.685 33.655 35.375 34.215 ;
        RECT 35.545 34.145 36.755 35.235 ;
        RECT 34.305 33.315 35.260 33.485 ;
        RECT 34.535 32.685 34.805 33.145 ;
        RECT 34.975 32.855 35.260 33.315 ;
        RECT 35.545 33.435 36.065 33.975 ;
        RECT 36.235 33.605 36.755 34.145 ;
        RECT 36.925 34.095 37.200 35.065 ;
        RECT 37.410 34.435 37.690 35.235 ;
        RECT 37.860 34.725 39.910 35.015 ;
        RECT 37.860 34.385 39.490 34.555 ;
        RECT 37.860 34.265 38.030 34.385 ;
        RECT 37.370 34.095 38.030 34.265 ;
        RECT 35.545 32.685 36.755 33.435 ;
        RECT 36.925 33.360 37.095 34.095 ;
        RECT 37.370 33.925 37.540 34.095 ;
        RECT 37.265 33.595 37.540 33.925 ;
        RECT 37.710 33.595 38.090 33.925 ;
        RECT 38.260 33.595 39.000 34.215 ;
        RECT 39.170 34.095 39.490 34.385 ;
        RECT 39.685 33.925 39.925 34.520 ;
        RECT 40.095 34.160 40.435 35.235 ;
        RECT 40.615 34.265 40.945 35.050 ;
        RECT 40.615 34.095 41.295 34.265 ;
        RECT 41.475 34.095 41.805 35.235 ;
        RECT 42.065 34.305 42.245 35.065 ;
        RECT 42.425 34.475 42.755 35.235 ;
        RECT 42.065 34.135 42.740 34.305 ;
        RECT 42.925 34.160 43.195 35.065 ;
        RECT 39.270 33.595 39.925 33.925 ;
        RECT 37.370 33.425 37.540 33.595 ;
        RECT 36.925 33.015 37.200 33.360 ;
        RECT 37.370 33.255 38.955 33.425 ;
        RECT 37.390 32.685 37.770 33.085 ;
        RECT 37.940 32.905 38.110 33.255 ;
        RECT 38.280 32.685 38.610 33.085 ;
        RECT 38.785 32.905 38.955 33.255 ;
        RECT 39.155 32.685 39.485 33.185 ;
        RECT 39.680 32.905 39.925 33.595 ;
        RECT 40.095 33.355 40.435 33.925 ;
        RECT 40.605 33.675 40.955 33.925 ;
        RECT 41.125 33.495 41.295 34.095 ;
        RECT 42.570 33.990 42.740 34.135 ;
        RECT 41.465 33.675 41.815 33.925 ;
        RECT 42.005 33.585 42.345 33.955 ;
        RECT 42.570 33.660 42.845 33.990 ;
        RECT 40.095 32.685 40.435 33.185 ;
        RECT 40.625 32.685 40.865 33.495 ;
        RECT 41.035 32.855 41.365 33.495 ;
        RECT 41.535 32.685 41.805 33.495 ;
        RECT 42.570 33.405 42.740 33.660 ;
        RECT 42.075 33.235 42.740 33.405 ;
        RECT 43.015 33.360 43.195 34.160 ;
        RECT 43.580 34.135 43.910 35.235 ;
        RECT 44.385 34.635 44.710 35.065 ;
        RECT 44.880 34.815 45.210 35.235 ;
        RECT 45.955 34.805 46.365 35.235 ;
        RECT 44.385 34.465 46.365 34.635 ;
        RECT 44.385 34.055 45.090 34.465 ;
        RECT 43.365 33.675 44.010 33.885 ;
        RECT 44.180 33.675 44.750 33.885 ;
        RECT 42.075 32.855 42.245 33.235 ;
        RECT 42.425 32.685 42.755 33.065 ;
        RECT 42.935 32.855 43.195 33.360 ;
        RECT 43.520 33.335 44.690 33.505 ;
        RECT 43.520 32.870 43.850 33.335 ;
        RECT 44.020 32.685 44.190 33.155 ;
        RECT 44.360 32.855 44.690 33.335 ;
        RECT 44.920 32.855 45.090 34.055 ;
        RECT 45.260 34.125 45.885 34.295 ;
        RECT 45.260 33.425 45.430 34.125 ;
        RECT 46.100 33.925 46.365 34.465 ;
        RECT 46.535 34.080 46.875 35.065 ;
        RECT 45.600 33.595 45.930 33.925 ;
        RECT 46.100 33.595 46.450 33.925 ;
        RECT 46.620 33.425 46.875 34.080 ;
        RECT 47.505 34.145 48.715 35.235 ;
        RECT 47.505 33.605 48.025 34.145 ;
        RECT 48.195 33.435 48.715 33.975 ;
        RECT 45.260 33.255 45.800 33.425 ;
        RECT 45.630 33.050 45.800 33.255 ;
        RECT 46.080 32.685 46.250 33.425 ;
        RECT 46.515 33.050 46.875 33.425 ;
        RECT 47.505 32.685 48.715 33.435 ;
        RECT 12.920 32.515 48.800 32.685 ;
        RECT 13.005 31.765 14.215 32.515 ;
        RECT 13.005 31.225 13.525 31.765 ;
        RECT 14.390 31.675 14.650 32.515 ;
        RECT 14.825 31.770 15.080 32.345 ;
        RECT 15.250 32.135 15.580 32.515 ;
        RECT 15.795 31.965 15.965 32.345 ;
        RECT 15.250 31.795 15.965 31.965 ;
        RECT 13.695 31.055 14.215 31.595 ;
        RECT 13.005 29.965 14.215 31.055 ;
        RECT 14.390 29.965 14.650 31.115 ;
        RECT 14.825 31.040 14.995 31.770 ;
        RECT 15.250 31.605 15.420 31.795 ;
        RECT 16.690 31.775 16.945 32.345 ;
        RECT 17.115 32.115 17.445 32.515 ;
        RECT 17.870 31.980 18.400 32.345 ;
        RECT 18.590 32.175 18.865 32.345 ;
        RECT 18.585 32.005 18.865 32.175 ;
        RECT 17.870 31.945 18.045 31.980 ;
        RECT 17.115 31.775 18.045 31.945 ;
        RECT 15.165 31.275 15.420 31.605 ;
        RECT 15.250 31.065 15.420 31.275 ;
        RECT 15.700 31.245 16.055 31.615 ;
        RECT 16.690 31.105 16.860 31.775 ;
        RECT 17.115 31.605 17.285 31.775 ;
        RECT 17.030 31.275 17.285 31.605 ;
        RECT 17.510 31.275 17.705 31.605 ;
        RECT 14.825 30.135 15.080 31.040 ;
        RECT 15.250 30.895 15.965 31.065 ;
        RECT 15.250 29.965 15.580 30.725 ;
        RECT 15.795 30.135 15.965 30.895 ;
        RECT 16.690 30.135 17.025 31.105 ;
        RECT 17.195 29.965 17.365 31.105 ;
        RECT 17.535 30.305 17.705 31.275 ;
        RECT 17.875 30.645 18.045 31.775 ;
        RECT 18.215 30.985 18.385 31.785 ;
        RECT 18.590 31.185 18.865 32.005 ;
        RECT 19.035 30.985 19.225 32.345 ;
        RECT 19.405 31.980 19.915 32.515 ;
        RECT 20.135 31.705 20.380 32.310 ;
        RECT 20.915 31.965 21.085 32.255 ;
        RECT 21.255 32.135 21.585 32.515 ;
        RECT 20.915 31.795 21.580 31.965 ;
        RECT 19.425 31.535 20.655 31.705 ;
        RECT 18.215 30.815 19.225 30.985 ;
        RECT 19.395 30.970 20.145 31.160 ;
        RECT 17.875 30.475 19.000 30.645 ;
        RECT 19.395 30.305 19.565 30.970 ;
        RECT 20.315 30.725 20.655 31.535 ;
        RECT 20.830 30.975 21.180 31.625 ;
        RECT 21.350 30.805 21.580 31.795 ;
        RECT 17.535 30.135 19.565 30.305 ;
        RECT 19.735 29.965 19.905 30.725 ;
        RECT 20.140 30.315 20.655 30.725 ;
        RECT 20.915 30.635 21.580 30.805 ;
        RECT 20.915 30.135 21.085 30.635 ;
        RECT 21.255 29.965 21.585 30.465 ;
        RECT 21.755 30.135 21.940 32.255 ;
        RECT 22.195 32.055 22.445 32.515 ;
        RECT 22.615 32.065 22.950 32.235 ;
        RECT 23.145 32.065 23.820 32.235 ;
        RECT 22.615 31.925 22.785 32.065 ;
        RECT 22.110 30.935 22.390 31.885 ;
        RECT 22.560 31.795 22.785 31.925 ;
        RECT 22.560 30.690 22.730 31.795 ;
        RECT 22.955 31.645 23.480 31.865 ;
        RECT 22.900 30.880 23.140 31.475 ;
        RECT 23.310 30.945 23.480 31.645 ;
        RECT 23.650 31.285 23.820 32.065 ;
        RECT 24.140 32.015 24.510 32.515 ;
        RECT 24.690 32.065 25.095 32.235 ;
        RECT 25.265 32.065 26.050 32.235 ;
        RECT 24.690 31.835 24.860 32.065 ;
        RECT 24.030 31.535 24.860 31.835 ;
        RECT 25.245 31.565 25.710 31.895 ;
        RECT 24.030 31.505 24.230 31.535 ;
        RECT 24.350 31.285 24.520 31.355 ;
        RECT 23.650 31.115 24.520 31.285 ;
        RECT 24.010 31.025 24.520 31.115 ;
        RECT 22.560 30.560 22.865 30.690 ;
        RECT 23.310 30.580 23.840 30.945 ;
        RECT 22.180 29.965 22.445 30.425 ;
        RECT 22.615 30.135 22.865 30.560 ;
        RECT 24.010 30.410 24.180 31.025 ;
        RECT 23.075 30.240 24.180 30.410 ;
        RECT 24.350 29.965 24.520 30.765 ;
        RECT 24.690 30.465 24.860 31.535 ;
        RECT 25.030 30.635 25.220 31.355 ;
        RECT 25.390 30.605 25.710 31.565 ;
        RECT 25.880 31.605 26.050 32.065 ;
        RECT 26.325 31.985 26.535 32.515 ;
        RECT 26.795 31.775 27.125 32.300 ;
        RECT 27.295 31.905 27.465 32.515 ;
        RECT 27.635 31.860 27.965 32.295 ;
        RECT 27.635 31.775 28.015 31.860 ;
        RECT 26.925 31.605 27.125 31.775 ;
        RECT 27.790 31.735 28.015 31.775 ;
        RECT 25.880 31.275 26.755 31.605 ;
        RECT 26.925 31.275 27.675 31.605 ;
        RECT 24.690 30.135 24.940 30.465 ;
        RECT 25.880 30.435 26.050 31.275 ;
        RECT 26.925 31.070 27.115 31.275 ;
        RECT 27.845 31.155 28.015 31.735 ;
        RECT 27.800 31.105 28.015 31.155 ;
        RECT 26.220 30.695 27.115 31.070 ;
        RECT 27.625 31.025 28.015 31.105 ;
        RECT 28.190 31.775 28.445 32.345 ;
        RECT 28.615 32.115 28.945 32.515 ;
        RECT 29.370 31.980 29.900 32.345 ;
        RECT 29.370 31.945 29.545 31.980 ;
        RECT 28.615 31.775 29.545 31.945 ;
        RECT 28.190 31.105 28.360 31.775 ;
        RECT 28.615 31.605 28.785 31.775 ;
        RECT 28.530 31.275 28.785 31.605 ;
        RECT 29.010 31.275 29.205 31.605 ;
        RECT 25.165 30.265 26.050 30.435 ;
        RECT 26.230 29.965 26.545 30.465 ;
        RECT 26.775 30.135 27.115 30.695 ;
        RECT 27.285 29.965 27.455 30.975 ;
        RECT 27.625 30.180 27.955 31.025 ;
        RECT 28.190 30.135 28.525 31.105 ;
        RECT 28.695 29.965 28.865 31.105 ;
        RECT 29.035 30.305 29.205 31.275 ;
        RECT 29.375 30.645 29.545 31.775 ;
        RECT 29.715 30.985 29.885 31.785 ;
        RECT 30.090 31.495 30.365 32.345 ;
        RECT 30.085 31.325 30.365 31.495 ;
        RECT 30.090 31.185 30.365 31.325 ;
        RECT 30.535 30.985 30.725 32.345 ;
        RECT 30.905 31.980 31.415 32.515 ;
        RECT 31.635 31.705 31.880 32.310 ;
        RECT 32.325 31.775 32.710 32.345 ;
        RECT 32.880 32.055 33.205 32.515 ;
        RECT 33.725 31.885 34.005 32.345 ;
        RECT 30.925 31.535 32.155 31.705 ;
        RECT 29.715 30.815 30.725 30.985 ;
        RECT 30.895 30.970 31.645 31.160 ;
        RECT 29.375 30.475 30.500 30.645 ;
        RECT 30.895 30.305 31.065 30.970 ;
        RECT 31.815 30.725 32.155 31.535 ;
        RECT 29.035 30.135 31.065 30.305 ;
        RECT 31.235 29.965 31.405 30.725 ;
        RECT 31.640 30.315 32.155 30.725 ;
        RECT 32.325 31.105 32.605 31.775 ;
        RECT 32.880 31.715 34.005 31.885 ;
        RECT 32.880 31.605 33.330 31.715 ;
        RECT 32.775 31.275 33.330 31.605 ;
        RECT 34.195 31.545 34.595 32.345 ;
        RECT 34.995 32.055 35.265 32.515 ;
        RECT 35.435 31.885 35.720 32.345 ;
        RECT 32.325 30.135 32.710 31.105 ;
        RECT 32.880 30.815 33.330 31.275 ;
        RECT 33.500 30.985 34.595 31.545 ;
        RECT 32.880 30.595 34.005 30.815 ;
        RECT 32.880 29.965 33.205 30.425 ;
        RECT 33.725 30.135 34.005 30.595 ;
        RECT 34.195 30.135 34.595 30.985 ;
        RECT 34.765 31.715 35.720 31.885 ;
        RECT 36.005 31.745 38.595 32.515 ;
        RECT 38.765 31.790 39.055 32.515 ;
        RECT 39.555 32.115 39.885 32.515 ;
        RECT 40.055 31.945 40.385 32.285 ;
        RECT 41.435 32.115 41.765 32.515 ;
        RECT 39.400 31.775 41.765 31.945 ;
        RECT 41.935 31.790 42.265 32.300 ;
        RECT 34.765 30.815 34.975 31.715 ;
        RECT 35.145 30.985 35.835 31.545 ;
        RECT 36.005 31.225 37.215 31.745 ;
        RECT 37.385 31.055 38.595 31.575 ;
        RECT 34.765 30.595 35.720 30.815 ;
        RECT 34.995 29.965 35.265 30.425 ;
        RECT 35.435 30.135 35.720 30.595 ;
        RECT 36.005 29.965 38.595 31.055 ;
        RECT 38.765 29.965 39.055 31.130 ;
        RECT 39.400 30.775 39.570 31.775 ;
        RECT 41.595 31.605 41.765 31.775 ;
        RECT 39.740 30.945 39.985 31.605 ;
        RECT 40.200 30.945 40.465 31.605 ;
        RECT 40.660 30.945 40.945 31.605 ;
        RECT 41.120 31.275 41.425 31.605 ;
        RECT 41.595 31.275 41.905 31.605 ;
        RECT 41.120 30.945 41.335 31.275 ;
        RECT 39.400 30.605 39.855 30.775 ;
        RECT 39.525 30.175 39.855 30.605 ;
        RECT 40.035 30.605 41.325 30.775 ;
        RECT 40.035 30.185 40.285 30.605 ;
        RECT 40.515 29.965 40.845 30.435 ;
        RECT 41.075 30.185 41.325 30.605 ;
        RECT 41.515 29.965 41.765 31.105 ;
        RECT 42.075 31.025 42.265 31.790 ;
        RECT 43.520 31.865 43.850 32.330 ;
        RECT 44.020 32.045 44.190 32.515 ;
        RECT 44.360 31.865 44.690 32.345 ;
        RECT 43.520 31.695 44.690 31.865 ;
        RECT 43.365 31.315 44.010 31.525 ;
        RECT 44.180 31.315 44.750 31.525 ;
        RECT 44.920 31.145 45.090 32.345 ;
        RECT 45.630 31.945 45.800 32.150 ;
        RECT 41.935 30.175 42.265 31.025 ;
        RECT 43.580 29.965 43.910 31.065 ;
        RECT 44.385 30.735 45.090 31.145 ;
        RECT 45.260 31.775 45.800 31.945 ;
        RECT 46.080 31.775 46.250 32.515 ;
        RECT 46.645 32.150 46.815 32.175 ;
        RECT 46.515 31.775 46.875 32.150 ;
        RECT 45.260 31.075 45.430 31.775 ;
        RECT 45.600 31.275 45.930 31.605 ;
        RECT 46.100 31.275 46.450 31.605 ;
        RECT 45.260 30.905 45.885 31.075 ;
        RECT 46.100 30.735 46.365 31.275 ;
        RECT 46.620 31.120 46.875 31.775 ;
        RECT 47.505 31.765 48.715 32.515 ;
        RECT 44.385 30.565 46.365 30.735 ;
        RECT 44.385 30.135 44.710 30.565 ;
        RECT 44.880 29.965 45.210 30.385 ;
        RECT 45.955 29.965 46.365 30.395 ;
        RECT 46.535 30.135 46.875 31.120 ;
        RECT 47.505 31.055 48.025 31.595 ;
        RECT 48.195 31.225 48.715 31.765 ;
        RECT 47.505 29.965 48.715 31.055 ;
        RECT 12.920 29.795 48.800 29.965 ;
        RECT 13.005 28.705 14.215 29.795 ;
        RECT 14.475 29.125 14.645 29.625 ;
        RECT 14.815 29.295 15.145 29.795 ;
        RECT 14.475 28.955 15.140 29.125 ;
        RECT 13.005 27.995 13.525 28.535 ;
        RECT 13.695 28.165 14.215 28.705 ;
        RECT 14.390 28.135 14.740 28.785 ;
        RECT 13.005 27.245 14.215 27.995 ;
        RECT 14.910 27.965 15.140 28.955 ;
        RECT 14.475 27.795 15.140 27.965 ;
        RECT 14.475 27.505 14.645 27.795 ;
        RECT 14.815 27.245 15.145 27.625 ;
        RECT 15.315 27.505 15.500 29.625 ;
        RECT 15.740 29.335 16.005 29.795 ;
        RECT 16.175 29.200 16.425 29.625 ;
        RECT 16.635 29.350 17.740 29.520 ;
        RECT 16.120 29.070 16.425 29.200 ;
        RECT 15.670 27.875 15.950 28.825 ;
        RECT 16.120 27.965 16.290 29.070 ;
        RECT 16.460 28.285 16.700 28.880 ;
        RECT 16.870 28.815 17.400 29.180 ;
        RECT 16.870 28.115 17.040 28.815 ;
        RECT 17.570 28.735 17.740 29.350 ;
        RECT 17.910 28.995 18.080 29.795 ;
        RECT 18.250 29.295 18.500 29.625 ;
        RECT 18.725 29.325 19.610 29.495 ;
        RECT 17.570 28.645 18.080 28.735 ;
        RECT 16.120 27.835 16.345 27.965 ;
        RECT 16.515 27.895 17.040 28.115 ;
        RECT 17.210 28.475 18.080 28.645 ;
        RECT 15.755 27.245 16.005 27.705 ;
        RECT 16.175 27.695 16.345 27.835 ;
        RECT 17.210 27.695 17.380 28.475 ;
        RECT 17.910 28.405 18.080 28.475 ;
        RECT 17.590 28.225 17.790 28.255 ;
        RECT 18.250 28.225 18.420 29.295 ;
        RECT 18.590 28.405 18.780 29.125 ;
        RECT 17.590 27.925 18.420 28.225 ;
        RECT 18.950 28.195 19.270 29.155 ;
        RECT 16.175 27.525 16.510 27.695 ;
        RECT 16.705 27.525 17.380 27.695 ;
        RECT 17.700 27.245 18.070 27.745 ;
        RECT 18.250 27.695 18.420 27.925 ;
        RECT 18.805 27.865 19.270 28.195 ;
        RECT 19.440 28.485 19.610 29.325 ;
        RECT 19.790 29.295 20.105 29.795 ;
        RECT 20.335 29.065 20.675 29.625 ;
        RECT 19.780 28.690 20.675 29.065 ;
        RECT 20.845 28.785 21.015 29.795 ;
        RECT 20.485 28.485 20.675 28.690 ;
        RECT 21.185 28.735 21.515 29.580 ;
        RECT 21.185 28.655 21.575 28.735 ;
        RECT 21.745 28.705 25.255 29.795 ;
        RECT 21.360 28.605 21.575 28.655 ;
        RECT 19.440 28.155 20.315 28.485 ;
        RECT 20.485 28.155 21.235 28.485 ;
        RECT 19.440 27.695 19.610 28.155 ;
        RECT 20.485 27.985 20.685 28.155 ;
        RECT 21.405 28.025 21.575 28.605 ;
        RECT 21.350 27.985 21.575 28.025 ;
        RECT 18.250 27.525 18.655 27.695 ;
        RECT 18.825 27.525 19.610 27.695 ;
        RECT 19.885 27.245 20.095 27.775 ;
        RECT 20.355 27.460 20.685 27.985 ;
        RECT 21.195 27.900 21.575 27.985 ;
        RECT 21.745 28.015 23.395 28.535 ;
        RECT 23.565 28.185 25.255 28.705 ;
        RECT 25.885 28.630 26.175 29.795 ;
        RECT 26.435 29.125 26.605 29.625 ;
        RECT 26.775 29.295 27.105 29.795 ;
        RECT 26.435 28.955 27.100 29.125 ;
        RECT 26.350 28.135 26.700 28.785 ;
        RECT 20.855 27.245 21.025 27.855 ;
        RECT 21.195 27.465 21.525 27.900 ;
        RECT 21.745 27.245 25.255 28.015 ;
        RECT 25.885 27.245 26.175 27.970 ;
        RECT 26.870 27.965 27.100 28.955 ;
        RECT 26.435 27.795 27.100 27.965 ;
        RECT 26.435 27.505 26.605 27.795 ;
        RECT 26.775 27.245 27.105 27.625 ;
        RECT 27.275 27.505 27.460 29.625 ;
        RECT 27.700 29.335 27.965 29.795 ;
        RECT 28.135 29.200 28.385 29.625 ;
        RECT 28.595 29.350 29.700 29.520 ;
        RECT 28.080 29.070 28.385 29.200 ;
        RECT 27.630 27.875 27.910 28.825 ;
        RECT 28.080 27.965 28.250 29.070 ;
        RECT 28.420 28.285 28.660 28.880 ;
        RECT 28.830 28.815 29.360 29.180 ;
        RECT 28.830 28.115 29.000 28.815 ;
        RECT 29.530 28.735 29.700 29.350 ;
        RECT 29.870 28.995 30.040 29.795 ;
        RECT 30.210 29.295 30.460 29.625 ;
        RECT 30.685 29.325 31.570 29.495 ;
        RECT 29.530 28.645 30.040 28.735 ;
        RECT 28.080 27.835 28.305 27.965 ;
        RECT 28.475 27.895 29.000 28.115 ;
        RECT 29.170 28.475 30.040 28.645 ;
        RECT 27.715 27.245 27.965 27.705 ;
        RECT 28.135 27.695 28.305 27.835 ;
        RECT 29.170 27.695 29.340 28.475 ;
        RECT 29.870 28.405 30.040 28.475 ;
        RECT 29.550 28.225 29.750 28.255 ;
        RECT 30.210 28.225 30.380 29.295 ;
        RECT 30.550 28.405 30.740 29.125 ;
        RECT 29.550 27.925 30.380 28.225 ;
        RECT 30.910 28.195 31.230 29.155 ;
        RECT 28.135 27.525 28.470 27.695 ;
        RECT 28.665 27.525 29.340 27.695 ;
        RECT 29.660 27.245 30.030 27.745 ;
        RECT 30.210 27.695 30.380 27.925 ;
        RECT 30.765 27.865 31.230 28.195 ;
        RECT 31.400 28.485 31.570 29.325 ;
        RECT 31.750 29.295 32.065 29.795 ;
        RECT 32.295 29.065 32.635 29.625 ;
        RECT 31.740 28.690 32.635 29.065 ;
        RECT 32.805 28.785 32.975 29.795 ;
        RECT 32.445 28.485 32.635 28.690 ;
        RECT 33.145 28.735 33.475 29.580 ;
        RECT 33.795 29.175 33.965 29.605 ;
        RECT 34.135 29.345 34.465 29.795 ;
        RECT 33.795 28.945 34.475 29.175 ;
        RECT 33.145 28.655 33.535 28.735 ;
        RECT 33.320 28.605 33.535 28.655 ;
        RECT 33.765 28.605 34.070 28.775 ;
        RECT 31.400 28.155 32.275 28.485 ;
        RECT 32.445 28.155 33.195 28.485 ;
        RECT 31.400 27.695 31.570 28.155 ;
        RECT 32.445 27.985 32.645 28.155 ;
        RECT 33.365 28.025 33.535 28.605 ;
        RECT 33.310 27.985 33.535 28.025 ;
        RECT 30.210 27.525 30.615 27.695 ;
        RECT 30.785 27.525 31.570 27.695 ;
        RECT 31.845 27.245 32.055 27.775 ;
        RECT 32.315 27.460 32.645 27.985 ;
        RECT 33.155 27.900 33.535 27.985 ;
        RECT 33.770 27.925 34.070 28.605 ;
        RECT 34.240 28.295 34.475 28.945 ;
        RECT 34.665 28.635 34.950 29.580 ;
        RECT 35.130 29.325 35.815 29.795 ;
        RECT 35.125 28.805 35.820 29.115 ;
        RECT 35.995 28.740 36.300 29.525 ;
        RECT 36.485 28.840 36.755 29.795 ;
        RECT 34.665 28.485 35.525 28.635 ;
        RECT 34.665 28.465 35.955 28.485 ;
        RECT 34.240 27.965 34.795 28.295 ;
        RECT 34.965 28.105 35.955 28.465 ;
        RECT 32.815 27.245 32.985 27.855 ;
        RECT 33.155 27.465 33.485 27.900 ;
        RECT 34.240 27.815 34.455 27.965 ;
        RECT 33.715 27.245 34.045 27.750 ;
        RECT 34.215 27.440 34.455 27.815 ;
        RECT 34.965 27.770 35.135 28.105 ;
        RECT 36.125 27.935 36.300 28.740 ;
        RECT 36.925 28.705 39.515 29.795 ;
        RECT 40.260 29.165 40.545 29.625 ;
        RECT 40.715 29.335 40.985 29.795 ;
        RECT 40.260 28.945 41.215 29.165 ;
        RECT 34.735 27.575 35.135 27.770 ;
        RECT 34.735 27.430 34.905 27.575 ;
        RECT 35.495 27.245 35.895 27.740 ;
        RECT 36.065 27.415 36.300 27.935 ;
        RECT 36.925 28.015 38.135 28.535 ;
        RECT 38.305 28.185 39.515 28.705 ;
        RECT 40.145 28.215 40.835 28.775 ;
        RECT 41.005 28.045 41.215 28.945 ;
        RECT 36.485 27.245 36.755 27.880 ;
        RECT 36.925 27.245 39.515 28.015 ;
        RECT 40.260 27.875 41.215 28.045 ;
        RECT 41.385 28.775 41.785 29.625 ;
        RECT 41.975 29.165 42.255 29.625 ;
        RECT 42.775 29.335 43.100 29.795 ;
        RECT 41.975 28.945 43.100 29.165 ;
        RECT 41.385 28.215 42.480 28.775 ;
        RECT 42.650 28.485 43.100 28.945 ;
        RECT 43.270 28.655 43.655 29.625 ;
        RECT 40.260 27.415 40.545 27.875 ;
        RECT 40.715 27.245 40.985 27.705 ;
        RECT 41.385 27.415 41.785 28.215 ;
        RECT 42.650 28.155 43.205 28.485 ;
        RECT 42.650 28.045 43.100 28.155 ;
        RECT 41.975 27.875 43.100 28.045 ;
        RECT 43.375 27.985 43.655 28.655 ;
        RECT 41.975 27.415 42.255 27.875 ;
        RECT 42.775 27.245 43.100 27.705 ;
        RECT 43.270 27.415 43.655 27.985 ;
        RECT 43.825 28.995 44.265 29.625 ;
        RECT 43.825 27.985 44.135 28.995 ;
        RECT 44.440 28.945 44.755 29.795 ;
        RECT 44.925 29.455 46.355 29.625 ;
        RECT 44.925 28.775 45.095 29.455 ;
        RECT 44.305 28.605 45.095 28.775 ;
        RECT 44.305 28.155 44.475 28.605 ;
        RECT 45.265 28.485 45.465 29.285 ;
        RECT 44.645 28.155 45.035 28.435 ;
        RECT 45.220 28.155 45.465 28.485 ;
        RECT 45.665 28.155 45.915 29.285 ;
        RECT 46.105 28.825 46.355 29.455 ;
        RECT 46.535 28.995 46.865 29.795 ;
        RECT 46.105 28.655 46.875 28.825 ;
        RECT 46.130 28.155 46.535 28.485 ;
        RECT 46.705 27.985 46.875 28.655 ;
        RECT 47.505 28.705 48.715 29.795 ;
        RECT 47.505 28.165 48.025 28.705 ;
        RECT 48.195 27.995 48.715 28.535 ;
        RECT 43.825 27.425 44.265 27.985 ;
        RECT 44.435 27.245 44.885 27.985 ;
        RECT 45.055 27.815 46.215 27.985 ;
        RECT 45.055 27.415 45.225 27.815 ;
        RECT 45.395 27.245 45.815 27.645 ;
        RECT 45.985 27.415 46.215 27.815 ;
        RECT 46.385 27.415 46.875 27.985 ;
        RECT 47.505 27.245 48.715 27.995 ;
        RECT 12.920 27.075 48.800 27.245 ;
        RECT 13.005 26.325 14.215 27.075 ;
        RECT 13.005 25.785 13.525 26.325 ;
        RECT 14.390 26.235 14.650 27.075 ;
        RECT 14.825 26.330 15.080 26.905 ;
        RECT 15.250 26.695 15.580 27.075 ;
        RECT 15.795 26.525 15.965 26.905 ;
        RECT 15.250 26.355 15.965 26.525 ;
        RECT 17.260 26.445 17.545 26.905 ;
        RECT 17.715 26.615 17.985 27.075 ;
        RECT 13.695 25.615 14.215 26.155 ;
        RECT 13.005 24.525 14.215 25.615 ;
        RECT 14.390 24.525 14.650 25.675 ;
        RECT 14.825 25.600 14.995 26.330 ;
        RECT 15.250 26.165 15.420 26.355 ;
        RECT 17.260 26.275 18.215 26.445 ;
        RECT 15.165 25.835 15.420 26.165 ;
        RECT 15.250 25.625 15.420 25.835 ;
        RECT 15.700 25.805 16.055 26.175 ;
        RECT 14.825 24.695 15.080 25.600 ;
        RECT 15.250 25.455 15.965 25.625 ;
        RECT 17.145 25.545 17.835 26.105 ;
        RECT 15.250 24.525 15.580 25.285 ;
        RECT 15.795 24.695 15.965 25.455 ;
        RECT 18.005 25.375 18.215 26.275 ;
        RECT 17.260 25.155 18.215 25.375 ;
        RECT 18.385 26.105 18.785 26.905 ;
        RECT 18.975 26.445 19.255 26.905 ;
        RECT 19.775 26.615 20.100 27.075 ;
        RECT 18.975 26.275 20.100 26.445 ;
        RECT 20.270 26.335 20.655 26.905 ;
        RECT 19.650 26.165 20.100 26.275 ;
        RECT 18.385 25.545 19.480 26.105 ;
        RECT 19.650 25.835 20.205 26.165 ;
        RECT 17.260 24.695 17.545 25.155 ;
        RECT 17.715 24.525 17.985 24.985 ;
        RECT 18.385 24.695 18.785 25.545 ;
        RECT 19.650 25.375 20.100 25.835 ;
        RECT 20.375 25.665 20.655 26.335 ;
        RECT 21.860 26.445 22.145 26.905 ;
        RECT 22.315 26.615 22.585 27.075 ;
        RECT 21.860 26.275 22.815 26.445 ;
        RECT 18.975 25.155 20.100 25.375 ;
        RECT 18.975 24.695 19.255 25.155 ;
        RECT 19.775 24.525 20.100 24.985 ;
        RECT 20.270 24.695 20.655 25.665 ;
        RECT 21.745 25.545 22.435 26.105 ;
        RECT 22.605 25.375 22.815 26.275 ;
        RECT 21.860 25.155 22.815 25.375 ;
        RECT 22.985 26.105 23.385 26.905 ;
        RECT 23.575 26.445 23.855 26.905 ;
        RECT 24.375 26.615 24.700 27.075 ;
        RECT 23.575 26.275 24.700 26.445 ;
        RECT 24.870 26.335 25.255 26.905 ;
        RECT 24.250 26.165 24.700 26.275 ;
        RECT 22.985 25.545 24.080 26.105 ;
        RECT 24.250 25.835 24.805 26.165 ;
        RECT 21.860 24.695 22.145 25.155 ;
        RECT 22.315 24.525 22.585 24.985 ;
        RECT 22.985 24.695 23.385 25.545 ;
        RECT 24.250 25.375 24.700 25.835 ;
        RECT 24.975 25.665 25.255 26.335 ;
        RECT 25.700 26.265 25.945 26.870 ;
        RECT 26.165 26.540 26.675 27.075 ;
        RECT 23.575 25.155 24.700 25.375 ;
        RECT 23.575 24.695 23.855 25.155 ;
        RECT 24.375 24.525 24.700 24.985 ;
        RECT 24.870 24.695 25.255 25.665 ;
        RECT 25.425 26.095 26.655 26.265 ;
        RECT 25.425 25.285 25.765 26.095 ;
        RECT 25.935 25.530 26.685 25.720 ;
        RECT 25.425 24.875 25.940 25.285 ;
        RECT 26.175 24.525 26.345 25.285 ;
        RECT 26.515 24.865 26.685 25.530 ;
        RECT 26.855 25.545 27.045 26.905 ;
        RECT 27.215 26.055 27.490 26.905 ;
        RECT 27.680 26.540 28.210 26.905 ;
        RECT 28.635 26.675 28.965 27.075 ;
        RECT 28.035 26.505 28.210 26.540 ;
        RECT 27.215 25.885 27.495 26.055 ;
        RECT 27.215 25.745 27.490 25.885 ;
        RECT 27.695 25.545 27.865 26.345 ;
        RECT 26.855 25.375 27.865 25.545 ;
        RECT 28.035 26.335 28.965 26.505 ;
        RECT 29.135 26.335 29.390 26.905 ;
        RECT 28.035 25.205 28.205 26.335 ;
        RECT 28.795 26.165 28.965 26.335 ;
        RECT 27.080 25.035 28.205 25.205 ;
        RECT 28.375 25.835 28.570 26.165 ;
        RECT 28.795 25.835 29.050 26.165 ;
        RECT 28.375 24.865 28.545 25.835 ;
        RECT 29.220 25.665 29.390 26.335 ;
        RECT 29.565 26.305 31.235 27.075 ;
        RECT 31.495 26.525 31.665 26.815 ;
        RECT 31.835 26.695 32.165 27.075 ;
        RECT 31.495 26.355 32.160 26.525 ;
        RECT 29.565 25.785 30.315 26.305 ;
        RECT 26.515 24.695 28.545 24.865 ;
        RECT 28.715 24.525 28.885 25.665 ;
        RECT 29.055 24.695 29.390 25.665 ;
        RECT 30.485 25.615 31.235 26.135 ;
        RECT 29.565 24.525 31.235 25.615 ;
        RECT 31.410 25.535 31.760 26.185 ;
        RECT 31.930 25.365 32.160 26.355 ;
        RECT 31.495 25.195 32.160 25.365 ;
        RECT 31.495 24.695 31.665 25.195 ;
        RECT 31.835 24.525 32.165 25.025 ;
        RECT 32.335 24.695 32.520 26.815 ;
        RECT 32.775 26.615 33.025 27.075 ;
        RECT 33.195 26.625 33.530 26.795 ;
        RECT 33.725 26.625 34.400 26.795 ;
        RECT 33.195 26.485 33.365 26.625 ;
        RECT 32.690 25.495 32.970 26.445 ;
        RECT 33.140 26.355 33.365 26.485 ;
        RECT 33.140 25.250 33.310 26.355 ;
        RECT 33.535 26.205 34.060 26.425 ;
        RECT 33.480 25.440 33.720 26.035 ;
        RECT 33.890 25.505 34.060 26.205 ;
        RECT 34.230 25.845 34.400 26.625 ;
        RECT 34.720 26.575 35.090 27.075 ;
        RECT 35.270 26.625 35.675 26.795 ;
        RECT 35.845 26.625 36.630 26.795 ;
        RECT 35.270 26.395 35.440 26.625 ;
        RECT 34.610 26.095 35.440 26.395 ;
        RECT 35.825 26.125 36.290 26.455 ;
        RECT 34.610 26.065 34.810 26.095 ;
        RECT 34.930 25.845 35.100 25.915 ;
        RECT 34.230 25.675 35.100 25.845 ;
        RECT 34.590 25.585 35.100 25.675 ;
        RECT 33.140 25.120 33.445 25.250 ;
        RECT 33.890 25.140 34.420 25.505 ;
        RECT 32.760 24.525 33.025 24.985 ;
        RECT 33.195 24.695 33.445 25.120 ;
        RECT 34.590 24.970 34.760 25.585 ;
        RECT 33.655 24.800 34.760 24.970 ;
        RECT 34.930 24.525 35.100 25.325 ;
        RECT 35.270 25.025 35.440 26.095 ;
        RECT 35.610 25.195 35.800 25.915 ;
        RECT 35.970 25.165 36.290 26.125 ;
        RECT 36.460 26.165 36.630 26.625 ;
        RECT 36.905 26.545 37.115 27.075 ;
        RECT 37.375 26.335 37.705 26.860 ;
        RECT 37.875 26.465 38.045 27.075 ;
        RECT 38.215 26.420 38.545 26.855 ;
        RECT 38.215 26.335 38.595 26.420 ;
        RECT 38.765 26.350 39.055 27.075 ;
        RECT 37.505 26.165 37.705 26.335 ;
        RECT 38.370 26.295 38.595 26.335 ;
        RECT 36.460 25.835 37.335 26.165 ;
        RECT 37.505 25.835 38.255 26.165 ;
        RECT 35.270 24.695 35.520 25.025 ;
        RECT 36.460 24.995 36.630 25.835 ;
        RECT 37.505 25.630 37.695 25.835 ;
        RECT 38.425 25.715 38.595 26.295 ;
        RECT 38.380 25.665 38.595 25.715 ;
        RECT 39.230 26.335 39.485 26.905 ;
        RECT 39.655 26.675 39.985 27.075 ;
        RECT 40.410 26.540 40.940 26.905 ;
        RECT 41.130 26.735 41.405 26.905 ;
        RECT 41.125 26.565 41.405 26.735 ;
        RECT 40.410 26.505 40.585 26.540 ;
        RECT 39.655 26.335 40.585 26.505 ;
        RECT 36.800 25.255 37.695 25.630 ;
        RECT 38.205 25.585 38.595 25.665 ;
        RECT 35.745 24.825 36.630 24.995 ;
        RECT 36.810 24.525 37.125 25.025 ;
        RECT 37.355 24.695 37.695 25.255 ;
        RECT 37.865 24.525 38.035 25.535 ;
        RECT 38.205 24.740 38.535 25.585 ;
        RECT 38.765 24.525 39.055 25.690 ;
        RECT 39.230 25.665 39.400 26.335 ;
        RECT 39.655 26.165 39.825 26.335 ;
        RECT 39.570 25.835 39.825 26.165 ;
        RECT 40.050 25.835 40.245 26.165 ;
        RECT 39.230 24.695 39.565 25.665 ;
        RECT 39.735 24.525 39.905 25.665 ;
        RECT 40.075 24.865 40.245 25.835 ;
        RECT 40.415 25.205 40.585 26.335 ;
        RECT 40.755 25.545 40.925 26.345 ;
        RECT 41.130 25.745 41.405 26.565 ;
        RECT 41.575 25.545 41.765 26.905 ;
        RECT 41.945 26.540 42.455 27.075 ;
        RECT 42.675 26.265 42.920 26.870 ;
        RECT 43.455 26.525 43.625 26.905 ;
        RECT 43.805 26.695 44.135 27.075 ;
        RECT 43.455 26.355 44.120 26.525 ;
        RECT 44.315 26.400 44.575 26.905 ;
        RECT 41.965 26.095 43.195 26.265 ;
        RECT 40.755 25.375 41.765 25.545 ;
        RECT 41.935 25.530 42.685 25.720 ;
        RECT 40.415 25.035 41.540 25.205 ;
        RECT 41.935 24.865 42.105 25.530 ;
        RECT 42.855 25.285 43.195 26.095 ;
        RECT 43.385 25.805 43.715 26.175 ;
        RECT 43.950 26.100 44.120 26.355 ;
        RECT 43.950 25.770 44.235 26.100 ;
        RECT 43.950 25.625 44.120 25.770 ;
        RECT 40.075 24.695 42.105 24.865 ;
        RECT 42.275 24.525 42.445 25.285 ;
        RECT 42.680 24.875 43.195 25.285 ;
        RECT 43.455 25.455 44.120 25.625 ;
        RECT 44.405 25.600 44.575 26.400 ;
        RECT 43.455 24.695 43.625 25.455 ;
        RECT 43.805 24.525 44.135 25.285 ;
        RECT 44.305 24.695 44.575 25.600 ;
        RECT 44.745 26.400 45.015 26.745 ;
        RECT 45.205 26.675 45.585 27.075 ;
        RECT 45.755 26.505 45.925 26.855 ;
        RECT 46.095 26.675 46.425 27.075 ;
        RECT 46.625 26.505 46.795 26.855 ;
        RECT 46.995 26.575 47.325 27.075 ;
        RECT 44.745 25.665 44.915 26.400 ;
        RECT 45.185 26.335 46.795 26.505 ;
        RECT 45.185 26.165 45.355 26.335 ;
        RECT 45.085 25.835 45.355 26.165 ;
        RECT 45.525 25.835 45.930 26.165 ;
        RECT 45.185 25.665 45.355 25.835 ;
        RECT 44.745 24.695 45.015 25.665 ;
        RECT 45.185 25.495 45.910 25.665 ;
        RECT 46.100 25.545 46.810 26.165 ;
        RECT 46.980 25.835 47.330 26.405 ;
        RECT 47.505 26.325 48.715 27.075 ;
        RECT 45.740 25.375 45.910 25.495 ;
        RECT 47.010 25.375 47.330 25.665 ;
        RECT 45.225 24.525 45.505 25.325 ;
        RECT 45.740 25.205 47.330 25.375 ;
        RECT 47.505 25.615 48.025 26.155 ;
        RECT 48.195 25.785 48.715 26.325 ;
        RECT 45.675 24.745 47.330 25.035 ;
        RECT 47.505 24.525 48.715 25.615 ;
        RECT 12.920 24.355 48.800 24.525 ;
        RECT 13.005 23.265 14.215 24.355 ;
        RECT 14.445 23.295 14.775 24.140 ;
        RECT 14.945 23.345 15.115 24.355 ;
        RECT 15.285 23.625 15.625 24.185 ;
        RECT 15.855 23.855 16.170 24.355 ;
        RECT 16.350 23.885 17.235 24.055 ;
        RECT 13.005 22.555 13.525 23.095 ;
        RECT 13.695 22.725 14.215 23.265 ;
        RECT 14.385 23.215 14.775 23.295 ;
        RECT 15.285 23.250 16.180 23.625 ;
        RECT 14.385 23.165 14.600 23.215 ;
        RECT 14.385 22.585 14.555 23.165 ;
        RECT 15.285 23.045 15.475 23.250 ;
        RECT 16.350 23.045 16.520 23.885 ;
        RECT 17.460 23.855 17.710 24.185 ;
        RECT 14.725 22.715 15.475 23.045 ;
        RECT 15.645 22.715 16.520 23.045 ;
        RECT 13.005 21.805 14.215 22.555 ;
        RECT 14.385 22.545 14.610 22.585 ;
        RECT 15.275 22.545 15.475 22.715 ;
        RECT 14.385 22.460 14.765 22.545 ;
        RECT 14.435 22.025 14.765 22.460 ;
        RECT 14.935 21.805 15.105 22.415 ;
        RECT 15.275 22.020 15.605 22.545 ;
        RECT 15.865 21.805 16.075 22.335 ;
        RECT 16.350 22.255 16.520 22.715 ;
        RECT 16.690 22.755 17.010 23.715 ;
        RECT 17.180 22.965 17.370 23.685 ;
        RECT 17.540 22.785 17.710 23.855 ;
        RECT 17.880 23.555 18.050 24.355 ;
        RECT 18.220 23.910 19.325 24.080 ;
        RECT 18.220 23.295 18.390 23.910 ;
        RECT 19.535 23.760 19.785 24.185 ;
        RECT 19.955 23.895 20.220 24.355 ;
        RECT 18.560 23.375 19.090 23.740 ;
        RECT 19.535 23.630 19.840 23.760 ;
        RECT 17.880 23.205 18.390 23.295 ;
        RECT 17.880 23.035 18.750 23.205 ;
        RECT 17.880 22.965 18.050 23.035 ;
        RECT 18.170 22.785 18.370 22.815 ;
        RECT 16.690 22.425 17.155 22.755 ;
        RECT 17.540 22.485 18.370 22.785 ;
        RECT 17.540 22.255 17.710 22.485 ;
        RECT 16.350 22.085 17.135 22.255 ;
        RECT 17.305 22.085 17.710 22.255 ;
        RECT 17.890 21.805 18.260 22.305 ;
        RECT 18.580 22.255 18.750 23.035 ;
        RECT 18.920 22.675 19.090 23.375 ;
        RECT 19.260 22.845 19.500 23.440 ;
        RECT 18.920 22.455 19.445 22.675 ;
        RECT 19.670 22.525 19.840 23.630 ;
        RECT 19.615 22.395 19.840 22.525 ;
        RECT 20.010 22.435 20.290 23.385 ;
        RECT 19.615 22.255 19.785 22.395 ;
        RECT 18.580 22.085 19.255 22.255 ;
        RECT 19.450 22.085 19.785 22.255 ;
        RECT 19.955 21.805 20.205 22.265 ;
        RECT 20.460 22.065 20.645 24.185 ;
        RECT 20.815 23.855 21.145 24.355 ;
        RECT 21.315 23.685 21.485 24.185 ;
        RECT 20.820 23.515 21.485 23.685 ;
        RECT 20.820 22.525 21.050 23.515 ;
        RECT 21.220 22.695 21.570 23.345 ;
        RECT 21.745 23.265 25.255 24.355 ;
        RECT 21.745 22.575 23.395 23.095 ;
        RECT 23.565 22.745 25.255 23.265 ;
        RECT 25.885 23.190 26.175 24.355 ;
        RECT 26.355 23.545 26.650 24.355 ;
        RECT 26.830 23.045 27.075 24.185 ;
        RECT 27.250 23.545 27.510 24.355 ;
        RECT 28.110 24.350 34.385 24.355 ;
        RECT 27.690 23.045 27.940 24.180 ;
        RECT 28.110 23.555 28.370 24.350 ;
        RECT 28.540 23.455 28.800 24.180 ;
        RECT 28.970 23.625 29.230 24.350 ;
        RECT 29.400 23.455 29.660 24.180 ;
        RECT 29.830 23.625 30.090 24.350 ;
        RECT 30.260 23.455 30.520 24.180 ;
        RECT 30.690 23.625 30.950 24.350 ;
        RECT 31.120 23.455 31.380 24.180 ;
        RECT 31.550 23.625 31.795 24.350 ;
        RECT 31.965 23.455 32.225 24.180 ;
        RECT 32.410 23.625 32.655 24.350 ;
        RECT 32.825 23.455 33.085 24.180 ;
        RECT 33.270 23.625 33.515 24.350 ;
        RECT 33.685 23.455 33.945 24.180 ;
        RECT 34.130 23.625 34.385 24.350 ;
        RECT 28.540 23.440 33.945 23.455 ;
        RECT 34.555 23.440 34.845 24.180 ;
        RECT 35.015 23.610 35.285 24.355 ;
        RECT 28.540 23.215 35.285 23.440 ;
        RECT 35.545 23.265 36.755 24.355 ;
        RECT 20.820 22.355 21.485 22.525 ;
        RECT 20.815 21.805 21.145 22.185 ;
        RECT 21.315 22.065 21.485 22.355 ;
        RECT 21.745 21.805 25.255 22.575 ;
        RECT 25.885 21.805 26.175 22.530 ;
        RECT 26.345 22.485 26.660 23.045 ;
        RECT 26.830 22.795 33.950 23.045 ;
        RECT 26.345 21.805 26.650 22.315 ;
        RECT 26.830 21.985 27.080 22.795 ;
        RECT 27.250 21.805 27.510 22.330 ;
        RECT 27.690 21.985 27.940 22.795 ;
        RECT 34.120 22.625 35.285 23.215 ;
        RECT 28.540 22.455 35.285 22.625 ;
        RECT 35.545 22.555 36.065 23.095 ;
        RECT 36.235 22.725 36.755 23.265 ;
        RECT 37.015 23.425 37.185 24.185 ;
        RECT 37.365 23.595 37.695 24.355 ;
        RECT 37.015 23.255 37.680 23.425 ;
        RECT 37.865 23.280 38.135 24.185 ;
        RECT 37.510 23.110 37.680 23.255 ;
        RECT 36.945 22.705 37.275 23.075 ;
        RECT 37.510 22.780 37.795 23.110 ;
        RECT 28.110 21.805 28.370 22.365 ;
        RECT 28.540 22.000 28.800 22.455 ;
        RECT 28.970 21.805 29.230 22.285 ;
        RECT 29.400 22.000 29.660 22.455 ;
        RECT 29.830 21.805 30.090 22.285 ;
        RECT 30.260 22.000 30.520 22.455 ;
        RECT 30.690 21.805 30.935 22.285 ;
        RECT 31.105 22.000 31.380 22.455 ;
        RECT 31.550 21.805 31.795 22.285 ;
        RECT 31.965 22.000 32.225 22.455 ;
        RECT 32.405 21.805 32.655 22.285 ;
        RECT 32.825 22.000 33.085 22.455 ;
        RECT 33.265 21.805 33.515 22.285 ;
        RECT 33.685 22.000 33.945 22.455 ;
        RECT 34.125 21.805 34.385 22.285 ;
        RECT 34.555 22.000 34.815 22.455 ;
        RECT 34.985 21.805 35.285 22.285 ;
        RECT 35.545 21.805 36.755 22.555 ;
        RECT 37.510 22.525 37.680 22.780 ;
        RECT 37.015 22.355 37.680 22.525 ;
        RECT 37.965 22.480 38.135 23.280 ;
        RECT 38.395 23.425 38.565 24.185 ;
        RECT 38.745 23.595 39.075 24.355 ;
        RECT 38.395 23.255 39.060 23.425 ;
        RECT 39.245 23.280 39.515 24.185 ;
        RECT 38.890 23.110 39.060 23.255 ;
        RECT 38.325 22.705 38.655 23.075 ;
        RECT 38.890 22.780 39.175 23.110 ;
        RECT 38.890 22.525 39.060 22.780 ;
        RECT 37.015 21.975 37.185 22.355 ;
        RECT 37.365 21.805 37.695 22.185 ;
        RECT 37.875 21.975 38.135 22.480 ;
        RECT 38.395 22.355 39.060 22.525 ;
        RECT 39.345 22.480 39.515 23.280 ;
        RECT 39.775 23.425 39.945 24.185 ;
        RECT 40.125 23.595 40.455 24.355 ;
        RECT 39.775 23.255 40.440 23.425 ;
        RECT 40.625 23.280 40.895 24.185 ;
        RECT 40.270 23.110 40.440 23.255 ;
        RECT 39.705 22.705 40.035 23.075 ;
        RECT 40.270 22.780 40.555 23.110 ;
        RECT 40.270 22.525 40.440 22.780 ;
        RECT 38.395 21.975 38.565 22.355 ;
        RECT 38.745 21.805 39.075 22.185 ;
        RECT 39.255 21.975 39.515 22.480 ;
        RECT 39.775 22.355 40.440 22.525 ;
        RECT 40.725 22.480 40.895 23.280 ;
        RECT 41.155 23.425 41.325 24.185 ;
        RECT 41.505 23.595 41.835 24.355 ;
        RECT 41.155 23.255 41.820 23.425 ;
        RECT 42.005 23.280 42.275 24.185 ;
        RECT 41.650 23.110 41.820 23.255 ;
        RECT 41.085 22.705 41.415 23.075 ;
        RECT 41.650 22.780 41.935 23.110 ;
        RECT 41.650 22.525 41.820 22.780 ;
        RECT 39.775 21.975 39.945 22.355 ;
        RECT 40.125 21.805 40.455 22.185 ;
        RECT 40.635 21.975 40.895 22.480 ;
        RECT 41.155 22.355 41.820 22.525 ;
        RECT 42.105 22.480 42.275 23.280 ;
        RECT 42.455 23.215 42.785 24.355 ;
        RECT 43.315 23.385 43.645 24.170 ;
        RECT 42.965 23.215 43.645 23.385 ;
        RECT 42.445 22.795 42.795 23.045 ;
        RECT 42.965 22.615 43.135 23.215 ;
        RECT 43.825 23.200 44.165 24.185 ;
        RECT 44.335 23.925 44.745 24.355 ;
        RECT 45.490 23.935 45.820 24.355 ;
        RECT 45.990 23.755 46.315 24.185 ;
        RECT 44.335 23.585 46.315 23.755 ;
        RECT 43.305 22.795 43.655 23.045 ;
        RECT 41.155 21.975 41.325 22.355 ;
        RECT 41.505 21.805 41.835 22.185 ;
        RECT 42.015 21.975 42.275 22.480 ;
        RECT 42.455 21.805 42.725 22.615 ;
        RECT 42.895 21.975 43.225 22.615 ;
        RECT 43.395 21.805 43.635 22.615 ;
        RECT 43.825 22.545 44.080 23.200 ;
        RECT 44.335 23.045 44.600 23.585 ;
        RECT 44.815 23.245 45.440 23.415 ;
        RECT 44.250 22.715 44.600 23.045 ;
        RECT 44.770 22.715 45.100 23.045 ;
        RECT 45.270 22.545 45.440 23.245 ;
        RECT 43.825 22.170 44.185 22.545 ;
        RECT 44.450 21.805 44.620 22.545 ;
        RECT 44.900 22.375 45.440 22.545 ;
        RECT 45.610 23.175 46.315 23.585 ;
        RECT 46.790 23.255 47.120 24.355 ;
        RECT 47.505 23.265 48.715 24.355 ;
        RECT 44.900 22.170 45.070 22.375 ;
        RECT 45.610 21.975 45.780 23.175 ;
        RECT 45.950 22.795 46.520 23.005 ;
        RECT 46.690 22.795 47.335 23.005 ;
        RECT 47.505 22.725 48.025 23.265 ;
        RECT 46.010 22.455 47.180 22.625 ;
        RECT 48.195 22.555 48.715 23.095 ;
        RECT 46.010 21.975 46.340 22.455 ;
        RECT 46.510 21.805 46.680 22.275 ;
        RECT 46.850 21.990 47.180 22.455 ;
        RECT 47.505 21.805 48.715 22.555 ;
        RECT 12.920 21.635 48.800 21.805 ;
        RECT 13.005 20.885 14.215 21.635 ;
        RECT 13.005 20.345 13.525 20.885 ;
        RECT 14.390 20.795 14.650 21.635 ;
        RECT 14.825 20.890 15.080 21.465 ;
        RECT 15.250 21.255 15.580 21.635 ;
        RECT 15.795 21.085 15.965 21.465 ;
        RECT 15.250 20.915 15.965 21.085 ;
        RECT 13.695 20.175 14.215 20.715 ;
        RECT 13.005 19.085 14.215 20.175 ;
        RECT 14.390 19.085 14.650 20.235 ;
        RECT 14.825 20.160 14.995 20.890 ;
        RECT 15.250 20.725 15.420 20.915 ;
        RECT 17.150 20.895 17.405 21.465 ;
        RECT 17.575 21.235 17.905 21.635 ;
        RECT 18.330 21.100 18.860 21.465 ;
        RECT 19.050 21.295 19.325 21.465 ;
        RECT 19.045 21.125 19.325 21.295 ;
        RECT 18.330 21.065 18.505 21.100 ;
        RECT 17.575 20.895 18.505 21.065 ;
        RECT 15.165 20.395 15.420 20.725 ;
        RECT 15.250 20.185 15.420 20.395 ;
        RECT 15.700 20.365 16.055 20.735 ;
        RECT 17.150 20.225 17.320 20.895 ;
        RECT 17.575 20.725 17.745 20.895 ;
        RECT 17.490 20.395 17.745 20.725 ;
        RECT 17.970 20.395 18.165 20.725 ;
        RECT 14.825 19.255 15.080 20.160 ;
        RECT 15.250 20.015 15.965 20.185 ;
        RECT 15.250 19.085 15.580 19.845 ;
        RECT 15.795 19.255 15.965 20.015 ;
        RECT 17.150 19.255 17.485 20.225 ;
        RECT 17.655 19.085 17.825 20.225 ;
        RECT 17.995 19.425 18.165 20.395 ;
        RECT 18.335 19.765 18.505 20.895 ;
        RECT 18.675 20.105 18.845 20.905 ;
        RECT 19.050 20.305 19.325 21.125 ;
        RECT 19.495 20.105 19.685 21.465 ;
        RECT 19.865 21.100 20.375 21.635 ;
        RECT 20.595 20.825 20.840 21.430 ;
        RECT 21.285 20.865 24.795 21.635 ;
        RECT 24.965 20.885 26.175 21.635 ;
        RECT 26.395 20.980 26.725 21.415 ;
        RECT 26.895 21.025 27.065 21.635 ;
        RECT 26.345 20.895 26.725 20.980 ;
        RECT 27.235 20.895 27.565 21.420 ;
        RECT 27.825 21.105 28.035 21.635 ;
        RECT 28.310 21.185 29.095 21.355 ;
        RECT 29.265 21.185 29.670 21.355 ;
        RECT 19.885 20.655 21.115 20.825 ;
        RECT 18.675 19.935 19.685 20.105 ;
        RECT 19.855 20.090 20.605 20.280 ;
        RECT 18.335 19.595 19.460 19.765 ;
        RECT 19.855 19.425 20.025 20.090 ;
        RECT 20.775 19.845 21.115 20.655 ;
        RECT 21.285 20.345 22.935 20.865 ;
        RECT 23.105 20.175 24.795 20.695 ;
        RECT 24.965 20.345 25.485 20.885 ;
        RECT 26.345 20.855 26.570 20.895 ;
        RECT 25.655 20.175 26.175 20.715 ;
        RECT 17.995 19.255 20.025 19.425 ;
        RECT 20.195 19.085 20.365 19.845 ;
        RECT 20.600 19.435 21.115 19.845 ;
        RECT 21.285 19.085 24.795 20.175 ;
        RECT 24.965 19.085 26.175 20.175 ;
        RECT 26.345 20.275 26.515 20.855 ;
        RECT 27.235 20.725 27.435 20.895 ;
        RECT 28.310 20.725 28.480 21.185 ;
        RECT 26.685 20.395 27.435 20.725 ;
        RECT 27.605 20.395 28.480 20.725 ;
        RECT 26.345 20.225 26.560 20.275 ;
        RECT 26.345 20.145 26.735 20.225 ;
        RECT 26.405 19.300 26.735 20.145 ;
        RECT 27.245 20.190 27.435 20.395 ;
        RECT 26.905 19.085 27.075 20.095 ;
        RECT 27.245 19.815 28.140 20.190 ;
        RECT 27.245 19.255 27.585 19.815 ;
        RECT 27.815 19.085 28.130 19.585 ;
        RECT 28.310 19.555 28.480 20.395 ;
        RECT 28.650 20.685 29.115 21.015 ;
        RECT 29.500 20.955 29.670 21.185 ;
        RECT 29.850 21.135 30.220 21.635 ;
        RECT 30.540 21.185 31.215 21.355 ;
        RECT 31.410 21.185 31.745 21.355 ;
        RECT 28.650 19.725 28.970 20.685 ;
        RECT 29.500 20.655 30.330 20.955 ;
        RECT 29.140 19.755 29.330 20.475 ;
        RECT 29.500 19.585 29.670 20.655 ;
        RECT 30.130 20.625 30.330 20.655 ;
        RECT 29.840 20.405 30.010 20.475 ;
        RECT 30.540 20.405 30.710 21.185 ;
        RECT 31.575 21.045 31.745 21.185 ;
        RECT 31.915 21.175 32.165 21.635 ;
        RECT 29.840 20.235 30.710 20.405 ;
        RECT 30.880 20.765 31.405 20.985 ;
        RECT 31.575 20.915 31.800 21.045 ;
        RECT 29.840 20.145 30.350 20.235 ;
        RECT 28.310 19.385 29.195 19.555 ;
        RECT 29.420 19.255 29.670 19.585 ;
        RECT 29.840 19.085 30.010 19.885 ;
        RECT 30.180 19.530 30.350 20.145 ;
        RECT 30.880 20.065 31.050 20.765 ;
        RECT 30.520 19.700 31.050 20.065 ;
        RECT 31.220 20.000 31.460 20.595 ;
        RECT 31.630 19.810 31.800 20.915 ;
        RECT 31.970 20.055 32.250 21.005 ;
        RECT 31.495 19.680 31.800 19.810 ;
        RECT 30.180 19.360 31.285 19.530 ;
        RECT 31.495 19.255 31.745 19.680 ;
        RECT 31.915 19.085 32.180 19.545 ;
        RECT 32.420 19.255 32.605 21.375 ;
        RECT 32.775 21.255 33.105 21.635 ;
        RECT 33.275 21.085 33.445 21.375 ;
        RECT 32.780 20.915 33.445 21.085 ;
        RECT 32.780 19.925 33.010 20.915 ;
        RECT 33.710 20.895 33.965 21.465 ;
        RECT 34.135 21.235 34.465 21.635 ;
        RECT 34.890 21.100 35.420 21.465 ;
        RECT 34.890 21.065 35.065 21.100 ;
        RECT 34.135 20.895 35.065 21.065 ;
        RECT 33.180 20.095 33.530 20.745 ;
        RECT 33.710 20.225 33.880 20.895 ;
        RECT 34.135 20.725 34.305 20.895 ;
        RECT 34.050 20.395 34.305 20.725 ;
        RECT 34.530 20.395 34.725 20.725 ;
        RECT 32.780 19.755 33.445 19.925 ;
        RECT 32.775 19.085 33.105 19.585 ;
        RECT 33.275 19.255 33.445 19.755 ;
        RECT 33.710 19.255 34.045 20.225 ;
        RECT 34.215 19.085 34.385 20.225 ;
        RECT 34.555 19.425 34.725 20.395 ;
        RECT 34.895 19.765 35.065 20.895 ;
        RECT 35.235 20.105 35.405 20.905 ;
        RECT 35.610 20.615 35.885 21.465 ;
        RECT 35.605 20.445 35.885 20.615 ;
        RECT 35.610 20.305 35.885 20.445 ;
        RECT 36.055 20.105 36.245 21.465 ;
        RECT 36.425 21.100 36.935 21.635 ;
        RECT 37.155 20.825 37.400 21.430 ;
        RECT 38.765 20.910 39.055 21.635 ;
        RECT 39.225 20.895 39.610 21.465 ;
        RECT 39.780 21.175 40.105 21.635 ;
        RECT 40.625 21.005 40.905 21.465 ;
        RECT 36.445 20.655 37.675 20.825 ;
        RECT 35.235 19.935 36.245 20.105 ;
        RECT 36.415 20.090 37.165 20.280 ;
        RECT 34.895 19.595 36.020 19.765 ;
        RECT 36.415 19.425 36.585 20.090 ;
        RECT 37.335 19.845 37.675 20.655 ;
        RECT 34.555 19.255 36.585 19.425 ;
        RECT 36.755 19.085 36.925 19.845 ;
        RECT 37.160 19.435 37.675 19.845 ;
        RECT 38.765 19.085 39.055 20.250 ;
        RECT 39.225 20.225 39.505 20.895 ;
        RECT 39.780 20.835 40.905 21.005 ;
        RECT 39.780 20.725 40.230 20.835 ;
        RECT 39.675 20.395 40.230 20.725 ;
        RECT 41.095 20.665 41.495 21.465 ;
        RECT 41.895 21.175 42.165 21.635 ;
        RECT 42.335 21.005 42.620 21.465 ;
        RECT 39.225 19.255 39.610 20.225 ;
        RECT 39.780 19.935 40.230 20.395 ;
        RECT 40.400 20.105 41.495 20.665 ;
        RECT 39.780 19.715 40.905 19.935 ;
        RECT 39.780 19.085 40.105 19.545 ;
        RECT 40.625 19.255 40.905 19.715 ;
        RECT 41.095 19.255 41.495 20.105 ;
        RECT 41.665 20.835 42.620 21.005 ;
        RECT 43.825 21.005 44.165 21.465 ;
        RECT 44.335 21.175 44.505 21.635 ;
        RECT 45.135 21.200 45.495 21.465 ;
        RECT 45.140 21.195 45.495 21.200 ;
        RECT 45.145 21.185 45.495 21.195 ;
        RECT 45.150 21.180 45.495 21.185 ;
        RECT 45.155 21.170 45.495 21.180 ;
        RECT 45.735 21.175 45.905 21.635 ;
        RECT 45.160 21.165 45.495 21.170 ;
        RECT 45.170 21.155 45.495 21.165 ;
        RECT 45.180 21.145 45.495 21.155 ;
        RECT 44.675 21.005 45.005 21.085 ;
        RECT 41.665 19.935 41.875 20.835 ;
        RECT 43.825 20.815 45.005 21.005 ;
        RECT 45.195 21.005 45.495 21.145 ;
        RECT 45.195 20.815 45.905 21.005 ;
        RECT 42.045 20.105 42.735 20.665 ;
        RECT 43.825 20.445 44.155 20.645 ;
        RECT 44.465 20.625 44.795 20.645 ;
        RECT 44.345 20.445 44.795 20.625 ;
        RECT 43.825 20.105 44.055 20.445 ;
        RECT 41.665 19.715 42.620 19.935 ;
        RECT 41.895 19.085 42.165 19.545 ;
        RECT 42.335 19.255 42.620 19.715 ;
        RECT 43.835 19.085 44.165 19.805 ;
        RECT 44.345 19.330 44.560 20.445 ;
        RECT 44.965 20.415 45.435 20.645 ;
        RECT 45.620 20.245 45.905 20.815 ;
        RECT 46.075 20.690 46.415 21.465 ;
        RECT 47.505 20.885 48.715 21.635 ;
        RECT 44.755 20.030 45.905 20.245 ;
        RECT 44.755 19.255 45.085 20.030 ;
        RECT 45.255 19.085 45.965 19.860 ;
        RECT 46.135 19.255 46.415 20.690 ;
        RECT 47.505 20.175 48.025 20.715 ;
        RECT 48.195 20.345 48.715 20.885 ;
        RECT 47.505 19.085 48.715 20.175 ;
        RECT 12.920 18.915 48.800 19.085 ;
        RECT 13.005 17.825 14.215 18.915 ;
        RECT 14.385 18.480 19.730 18.915 ;
        RECT 13.005 17.115 13.525 17.655 ;
        RECT 13.695 17.285 14.215 17.825 ;
        RECT 13.005 16.365 14.215 17.115 ;
        RECT 15.970 16.910 16.310 17.740 ;
        RECT 17.790 17.230 18.140 18.480 ;
        RECT 19.905 17.825 23.415 18.915 ;
        RECT 19.905 17.135 21.555 17.655 ;
        RECT 21.725 17.305 23.415 17.825 ;
        RECT 24.135 17.985 24.305 18.745 ;
        RECT 24.520 18.155 24.850 18.915 ;
        RECT 24.135 17.815 24.850 17.985 ;
        RECT 25.020 17.840 25.275 18.745 ;
        RECT 24.045 17.265 24.400 17.635 ;
        RECT 24.680 17.605 24.850 17.815 ;
        RECT 24.680 17.275 24.935 17.605 ;
        RECT 14.385 16.365 19.730 16.910 ;
        RECT 19.905 16.365 23.415 17.135 ;
        RECT 24.680 17.085 24.850 17.275 ;
        RECT 25.105 17.110 25.275 17.840 ;
        RECT 25.450 17.765 25.710 18.915 ;
        RECT 25.885 17.750 26.175 18.915 ;
        RECT 26.810 17.765 27.070 18.915 ;
        RECT 27.245 17.840 27.500 18.745 ;
        RECT 27.670 18.155 28.000 18.915 ;
        RECT 28.215 17.985 28.385 18.745 ;
        RECT 28.735 18.245 28.905 18.745 ;
        RECT 29.075 18.415 29.405 18.915 ;
        RECT 28.735 18.075 29.400 18.245 ;
        RECT 24.135 16.915 24.850 17.085 ;
        RECT 24.135 16.535 24.305 16.915 ;
        RECT 24.520 16.365 24.850 16.745 ;
        RECT 25.020 16.535 25.275 17.110 ;
        RECT 25.450 16.365 25.710 17.205 ;
        RECT 25.885 16.365 26.175 17.090 ;
        RECT 26.810 16.365 27.070 17.205 ;
        RECT 27.245 17.110 27.415 17.840 ;
        RECT 27.670 17.815 28.385 17.985 ;
        RECT 27.670 17.605 27.840 17.815 ;
        RECT 27.585 17.275 27.840 17.605 ;
        RECT 27.245 16.535 27.500 17.110 ;
        RECT 27.670 17.085 27.840 17.275 ;
        RECT 28.120 17.265 28.475 17.635 ;
        RECT 28.650 17.255 29.000 17.905 ;
        RECT 29.170 17.085 29.400 18.075 ;
        RECT 27.670 16.915 28.385 17.085 ;
        RECT 27.670 16.365 28.000 16.745 ;
        RECT 28.215 16.535 28.385 16.915 ;
        RECT 28.735 16.915 29.400 17.085 ;
        RECT 28.735 16.625 28.905 16.915 ;
        RECT 29.075 16.365 29.405 16.745 ;
        RECT 29.575 16.625 29.760 18.745 ;
        RECT 30.000 18.455 30.265 18.915 ;
        RECT 30.435 18.320 30.685 18.745 ;
        RECT 30.895 18.470 32.000 18.640 ;
        RECT 30.380 18.190 30.685 18.320 ;
        RECT 29.930 16.995 30.210 17.945 ;
        RECT 30.380 17.085 30.550 18.190 ;
        RECT 30.720 17.405 30.960 18.000 ;
        RECT 31.130 17.935 31.660 18.300 ;
        RECT 31.130 17.235 31.300 17.935 ;
        RECT 31.830 17.855 32.000 18.470 ;
        RECT 32.170 18.115 32.340 18.915 ;
        RECT 32.510 18.415 32.760 18.745 ;
        RECT 32.985 18.445 33.870 18.615 ;
        RECT 31.830 17.765 32.340 17.855 ;
        RECT 30.380 16.955 30.605 17.085 ;
        RECT 30.775 17.015 31.300 17.235 ;
        RECT 31.470 17.595 32.340 17.765 ;
        RECT 30.015 16.365 30.265 16.825 ;
        RECT 30.435 16.815 30.605 16.955 ;
        RECT 31.470 16.815 31.640 17.595 ;
        RECT 32.170 17.525 32.340 17.595 ;
        RECT 31.850 17.345 32.050 17.375 ;
        RECT 32.510 17.345 32.680 18.415 ;
        RECT 32.850 17.525 33.040 18.245 ;
        RECT 31.850 17.045 32.680 17.345 ;
        RECT 33.210 17.315 33.530 18.275 ;
        RECT 30.435 16.645 30.770 16.815 ;
        RECT 30.965 16.645 31.640 16.815 ;
        RECT 31.960 16.365 32.330 16.865 ;
        RECT 32.510 16.815 32.680 17.045 ;
        RECT 33.065 16.985 33.530 17.315 ;
        RECT 33.700 17.605 33.870 18.445 ;
        RECT 34.050 18.415 34.365 18.915 ;
        RECT 34.595 18.185 34.935 18.745 ;
        RECT 34.040 17.810 34.935 18.185 ;
        RECT 35.105 17.905 35.275 18.915 ;
        RECT 34.745 17.605 34.935 17.810 ;
        RECT 35.445 17.855 35.775 18.700 ;
        RECT 35.445 17.775 35.835 17.855 ;
        RECT 35.620 17.725 35.835 17.775 ;
        RECT 36.010 17.765 36.270 18.915 ;
        RECT 36.445 17.840 36.700 18.745 ;
        RECT 36.870 18.155 37.200 18.915 ;
        RECT 37.415 17.985 37.585 18.745 ;
        RECT 33.700 17.275 34.575 17.605 ;
        RECT 34.745 17.275 35.495 17.605 ;
        RECT 33.700 16.815 33.870 17.275 ;
        RECT 34.745 17.105 34.945 17.275 ;
        RECT 35.665 17.145 35.835 17.725 ;
        RECT 35.610 17.105 35.835 17.145 ;
        RECT 32.510 16.645 32.915 16.815 ;
        RECT 33.085 16.645 33.870 16.815 ;
        RECT 34.145 16.365 34.355 16.895 ;
        RECT 34.615 16.580 34.945 17.105 ;
        RECT 35.455 17.020 35.835 17.105 ;
        RECT 35.115 16.365 35.285 16.975 ;
        RECT 35.455 16.585 35.785 17.020 ;
        RECT 36.010 16.365 36.270 17.205 ;
        RECT 36.445 17.110 36.615 17.840 ;
        RECT 36.870 17.815 37.585 17.985 ;
        RECT 36.870 17.605 37.040 17.815 ;
        RECT 38.765 17.750 39.055 18.915 ;
        RECT 40.235 17.985 40.405 18.745 ;
        RECT 40.620 18.155 40.950 18.915 ;
        RECT 40.235 17.815 40.950 17.985 ;
        RECT 41.120 17.840 41.375 18.745 ;
        RECT 36.785 17.275 37.040 17.605 ;
        RECT 36.445 16.535 36.700 17.110 ;
        RECT 36.870 17.085 37.040 17.275 ;
        RECT 37.320 17.265 37.675 17.635 ;
        RECT 40.145 17.265 40.500 17.635 ;
        RECT 40.780 17.605 40.950 17.815 ;
        RECT 40.780 17.275 41.035 17.605 ;
        RECT 36.870 16.915 37.585 17.085 ;
        RECT 36.870 16.365 37.200 16.745 ;
        RECT 37.415 16.535 37.585 16.915 ;
        RECT 38.765 16.365 39.055 17.090 ;
        RECT 40.780 17.085 40.950 17.275 ;
        RECT 41.205 17.110 41.375 17.840 ;
        RECT 41.550 17.765 41.810 18.915 ;
        RECT 41.985 17.840 42.255 18.745 ;
        RECT 42.425 18.155 42.755 18.915 ;
        RECT 42.935 17.985 43.115 18.745 ;
        RECT 44.375 18.295 44.545 18.725 ;
        RECT 44.715 18.465 45.045 18.915 ;
        RECT 44.375 18.065 45.050 18.295 ;
        RECT 40.235 16.915 40.950 17.085 ;
        RECT 40.235 16.535 40.405 16.915 ;
        RECT 40.620 16.365 40.950 16.745 ;
        RECT 41.120 16.535 41.375 17.110 ;
        RECT 41.550 16.365 41.810 17.205 ;
        RECT 41.985 17.040 42.165 17.840 ;
        RECT 42.440 17.815 43.115 17.985 ;
        RECT 42.440 17.670 42.610 17.815 ;
        RECT 42.335 17.340 42.610 17.670 ;
        RECT 42.440 17.085 42.610 17.340 ;
        RECT 42.835 17.265 43.175 17.635 ;
        RECT 41.985 16.535 42.245 17.040 ;
        RECT 42.440 16.915 43.105 17.085 ;
        RECT 44.345 17.045 44.645 17.895 ;
        RECT 44.815 17.415 45.050 18.065 ;
        RECT 45.220 17.755 45.505 18.700 ;
        RECT 45.685 18.445 46.370 18.915 ;
        RECT 45.680 17.925 46.375 18.235 ;
        RECT 46.550 17.860 46.855 18.645 ;
        RECT 45.220 17.605 46.080 17.755 ;
        RECT 45.220 17.585 46.505 17.605 ;
        RECT 44.815 17.085 45.350 17.415 ;
        RECT 45.520 17.225 46.505 17.585 ;
        RECT 44.815 16.935 45.035 17.085 ;
        RECT 42.425 16.365 42.755 16.745 ;
        RECT 42.935 16.535 43.105 16.915 ;
        RECT 44.290 16.365 44.625 16.870 ;
        RECT 44.795 16.560 45.035 16.935 ;
        RECT 45.520 16.890 45.690 17.225 ;
        RECT 46.680 17.055 46.855 17.860 ;
        RECT 47.505 17.825 48.715 18.915 ;
        RECT 47.505 17.285 48.025 17.825 ;
        RECT 48.195 17.115 48.715 17.655 ;
        RECT 45.315 16.695 45.690 16.890 ;
        RECT 45.315 16.550 45.485 16.695 ;
        RECT 46.050 16.365 46.445 16.860 ;
        RECT 46.615 16.535 46.855 17.055 ;
        RECT 47.505 16.365 48.715 17.115 ;
        RECT 12.920 16.195 48.800 16.365 ;
      LAYER met1 ;
        RECT 13.330 211.780 138.910 212.260 ;
        RECT 72.280 211.580 72.600 211.640 ;
        RECT 73.215 211.580 73.505 211.625 ;
        RECT 72.280 211.440 73.505 211.580 ;
        RECT 72.280 211.380 72.600 211.440 ;
        RECT 73.215 211.395 73.505 211.440 ;
        RECT 73.660 210.900 73.980 210.960 ;
        RECT 74.135 210.900 74.425 210.945 ;
        RECT 73.660 210.760 74.425 210.900 ;
        RECT 73.660 210.700 73.980 210.760 ;
        RECT 74.135 210.715 74.425 210.760 ;
        RECT 13.330 209.060 138.910 209.540 ;
        RECT 13.330 206.340 138.910 206.820 ;
        RECT 13.330 203.620 138.910 204.100 ;
        RECT 13.330 200.900 138.910 201.380 ;
        RECT 54.800 200.020 55.120 200.080 ;
        RECT 64.015 200.020 64.305 200.065 ;
        RECT 54.800 199.880 64.305 200.020 ;
        RECT 54.800 199.820 55.120 199.880 ;
        RECT 64.015 199.835 64.305 199.880 ;
        RECT 66.315 200.020 66.605 200.065 ;
        RECT 67.220 200.020 67.540 200.080 ;
        RECT 68.140 200.065 68.460 200.080 ;
        RECT 66.315 199.880 67.540 200.020 ;
        RECT 66.315 199.835 66.605 199.880 ;
        RECT 67.220 199.820 67.540 199.880 ;
        RECT 68.110 199.835 68.460 200.065 ;
        RECT 68.140 199.820 68.460 199.835 ;
        RECT 77.340 200.020 77.660 200.080 ;
        RECT 79.655 200.020 79.945 200.065 ;
        RECT 77.340 199.880 79.945 200.020 ;
        RECT 77.340 199.820 77.660 199.880 ;
        RECT 79.655 199.835 79.945 199.880 ;
        RECT 114.615 200.020 114.905 200.065 ;
        RECT 116.440 200.020 116.760 200.080 ;
        RECT 114.615 199.880 116.760 200.020 ;
        RECT 114.615 199.835 114.905 199.880 ;
        RECT 116.440 199.820 116.760 199.880 ;
        RECT 66.760 199.480 67.080 199.740 ;
        RECT 67.655 199.680 67.945 199.725 ;
        RECT 68.845 199.680 69.135 199.725 ;
        RECT 71.365 199.680 71.655 199.725 ;
        RECT 67.655 199.540 71.655 199.680 ;
        RECT 67.655 199.495 67.945 199.540 ;
        RECT 68.845 199.495 69.135 199.540 ;
        RECT 71.365 199.495 71.655 199.540 ;
        RECT 74.580 199.680 74.900 199.740 ;
        RECT 76.895 199.680 77.185 199.725 ;
        RECT 74.580 199.540 77.185 199.680 ;
        RECT 74.580 199.480 74.900 199.540 ;
        RECT 76.895 199.495 77.185 199.540 ;
        RECT 62.160 199.340 62.480 199.400 ;
        RECT 65.855 199.340 66.145 199.385 ;
        RECT 62.160 199.200 66.145 199.340 ;
        RECT 62.160 199.140 62.480 199.200 ;
        RECT 65.855 199.155 66.145 199.200 ;
        RECT 67.260 199.340 67.550 199.385 ;
        RECT 69.360 199.340 69.650 199.385 ;
        RECT 70.930 199.340 71.220 199.385 ;
        RECT 67.260 199.200 71.220 199.340 ;
        RECT 67.260 199.155 67.550 199.200 ;
        RECT 69.360 199.155 69.650 199.200 ;
        RECT 70.930 199.155 71.220 199.200 ;
        RECT 73.660 199.140 73.980 199.400 ;
        RECT 63.080 198.800 63.400 199.060 ;
        RECT 74.120 198.800 74.440 199.060 ;
        RECT 79.180 198.800 79.500 199.060 ;
        RECT 113.680 198.800 114.000 199.060 ;
        RECT 13.330 198.180 138.910 198.660 ;
        RECT 74.120 197.980 74.440 198.040 ;
        RECT 99.895 197.980 100.185 198.025 ;
        RECT 68.230 197.840 74.440 197.980 ;
        RECT 64.475 196.960 64.765 197.005 ;
        RECT 64.920 196.960 65.240 197.020 ;
        RECT 64.475 196.820 65.240 196.960 ;
        RECT 64.475 196.775 64.765 196.820 ;
        RECT 64.920 196.760 65.240 196.820 ;
        RECT 65.855 196.775 66.145 197.005 ;
        RECT 66.300 196.960 66.620 197.020 ;
        RECT 68.230 197.005 68.370 197.840 ;
        RECT 74.120 197.780 74.440 197.840 ;
        RECT 98.590 197.840 100.185 197.980 ;
        RECT 70.440 197.640 70.760 197.700 ;
        RECT 68.690 197.500 70.760 197.640 ;
        RECT 68.690 197.345 68.830 197.500 ;
        RECT 70.440 197.440 70.760 197.500 ;
        RECT 70.940 197.640 71.230 197.685 ;
        RECT 73.040 197.640 73.330 197.685 ;
        RECT 74.610 197.640 74.900 197.685 ;
        RECT 70.940 197.500 74.900 197.640 ;
        RECT 70.940 197.455 71.230 197.500 ;
        RECT 73.040 197.455 73.330 197.500 ;
        RECT 74.610 197.455 74.900 197.500 ;
        RECT 94.360 197.640 94.650 197.685 ;
        RECT 95.930 197.640 96.220 197.685 ;
        RECT 98.030 197.640 98.320 197.685 ;
        RECT 94.360 197.500 98.320 197.640 ;
        RECT 94.360 197.455 94.650 197.500 ;
        RECT 95.930 197.455 96.220 197.500 ;
        RECT 98.030 197.455 98.320 197.500 ;
        RECT 68.615 197.115 68.905 197.345 ;
        RECT 71.335 197.300 71.625 197.345 ;
        RECT 72.525 197.300 72.815 197.345 ;
        RECT 75.045 197.300 75.335 197.345 ;
        RECT 69.150 197.160 71.175 197.300 ;
        RECT 66.775 196.960 67.065 197.005 ;
        RECT 66.300 196.820 67.065 196.960 ;
        RECT 65.930 196.620 66.070 196.775 ;
        RECT 66.300 196.760 66.620 196.820 ;
        RECT 66.775 196.775 67.065 196.820 ;
        RECT 68.155 196.775 68.445 197.005 ;
        RECT 67.220 196.620 67.540 196.680 ;
        RECT 65.930 196.480 67.540 196.620 ;
        RECT 67.220 196.420 67.540 196.480 ;
        RECT 69.150 196.340 69.290 197.160 ;
        RECT 69.520 196.960 69.840 197.020 ;
        RECT 70.455 196.960 70.745 197.005 ;
        RECT 69.520 196.820 70.745 196.960 ;
        RECT 71.035 196.960 71.175 197.160 ;
        RECT 71.335 197.160 75.335 197.300 ;
        RECT 71.335 197.115 71.625 197.160 ;
        RECT 72.525 197.115 72.815 197.160 ;
        RECT 75.045 197.115 75.335 197.160 ;
        RECT 93.925 197.300 94.215 197.345 ;
        RECT 96.445 197.300 96.735 197.345 ;
        RECT 97.635 197.300 97.925 197.345 ;
        RECT 98.590 197.300 98.730 197.840 ;
        RECT 99.895 197.795 100.185 197.840 ;
        RECT 111.380 197.640 111.670 197.685 ;
        RECT 112.950 197.640 113.240 197.685 ;
        RECT 115.050 197.640 115.340 197.685 ;
        RECT 111.380 197.500 115.340 197.640 ;
        RECT 111.380 197.455 111.670 197.500 ;
        RECT 112.950 197.455 113.240 197.500 ;
        RECT 115.050 197.455 115.340 197.500 ;
        RECT 118.740 197.640 119.030 197.685 ;
        RECT 120.310 197.640 120.600 197.685 ;
        RECT 122.410 197.640 122.700 197.685 ;
        RECT 118.740 197.500 122.700 197.640 ;
        RECT 118.740 197.455 119.030 197.500 ;
        RECT 120.310 197.455 120.600 197.500 ;
        RECT 122.410 197.455 122.700 197.500 ;
        RECT 93.925 197.160 97.925 197.300 ;
        RECT 93.925 197.115 94.215 197.160 ;
        RECT 96.445 197.115 96.735 197.160 ;
        RECT 97.635 197.115 97.925 197.160 ;
        RECT 98.130 197.160 98.730 197.300 ;
        RECT 78.275 196.960 78.565 197.005 ;
        RECT 71.035 196.820 78.565 196.960 ;
        RECT 69.520 196.760 69.840 196.820 ;
        RECT 70.455 196.775 70.745 196.820 ;
        RECT 78.275 196.775 78.565 196.820 ;
        RECT 89.315 196.775 89.605 197.005 ;
        RECT 90.235 196.960 90.525 197.005 ;
        RECT 95.740 196.960 96.060 197.020 ;
        RECT 90.235 196.820 96.060 196.960 ;
        RECT 90.235 196.775 90.525 196.820 ;
        RECT 71.680 196.620 71.970 196.665 ;
        RECT 70.070 196.480 71.970 196.620 ;
        RECT 61.255 196.280 61.545 196.325 ;
        RECT 62.620 196.280 62.940 196.340 ;
        RECT 61.255 196.140 62.940 196.280 ;
        RECT 61.255 196.095 61.545 196.140 ;
        RECT 62.620 196.080 62.940 196.140 ;
        RECT 66.315 196.280 66.605 196.325 ;
        RECT 69.060 196.280 69.380 196.340 ;
        RECT 70.070 196.325 70.210 196.480 ;
        RECT 71.680 196.435 71.970 196.480 ;
        RECT 73.660 196.620 73.980 196.680 ;
        RECT 79.195 196.620 79.485 196.665 ;
        RECT 73.660 196.480 79.485 196.620 ;
        RECT 89.390 196.620 89.530 196.775 ;
        RECT 95.740 196.760 96.060 196.820 ;
        RECT 97.235 196.960 97.525 197.005 ;
        RECT 98.130 196.960 98.270 197.160 ;
        RECT 99.895 197.115 100.185 197.345 ;
        RECT 100.355 197.300 100.645 197.345 ;
        RECT 102.655 197.300 102.945 197.345 ;
        RECT 104.020 197.300 104.340 197.360 ;
        RECT 100.355 197.160 101.950 197.300 ;
        RECT 100.355 197.115 100.645 197.160 ;
        RECT 97.235 196.820 98.270 196.960 ;
        RECT 97.235 196.775 97.525 196.820 ;
        RECT 98.500 196.760 98.820 197.020 ;
        RECT 98.975 196.620 99.265 196.665 ;
        RECT 99.420 196.620 99.740 196.680 ;
        RECT 89.390 196.480 99.740 196.620 ;
        RECT 73.660 196.420 73.980 196.480 ;
        RECT 79.195 196.435 79.485 196.480 ;
        RECT 98.975 196.435 99.265 196.480 ;
        RECT 99.420 196.420 99.740 196.480 ;
        RECT 66.315 196.140 69.380 196.280 ;
        RECT 66.315 196.095 66.605 196.140 ;
        RECT 69.060 196.080 69.380 196.140 ;
        RECT 69.995 196.095 70.285 196.325 ;
        RECT 74.580 196.280 74.900 196.340 ;
        RECT 77.355 196.280 77.645 196.325 ;
        RECT 74.580 196.140 77.645 196.280 ;
        RECT 74.580 196.080 74.900 196.140 ;
        RECT 77.355 196.095 77.645 196.140 ;
        RECT 80.100 196.080 80.420 196.340 ;
        RECT 89.775 196.280 90.065 196.325 ;
        RECT 90.680 196.280 91.000 196.340 ;
        RECT 89.775 196.140 91.000 196.280 ;
        RECT 89.775 196.095 90.065 196.140 ;
        RECT 90.680 196.080 91.000 196.140 ;
        RECT 91.600 196.080 91.920 196.340 ;
        RECT 97.120 196.280 97.440 196.340 ;
        RECT 99.970 196.280 100.110 197.115 ;
        RECT 100.815 196.775 101.105 197.005 ;
        RECT 97.120 196.140 100.110 196.280 ;
        RECT 100.890 196.280 101.030 196.775 ;
        RECT 101.260 196.760 101.580 197.020 ;
        RECT 101.810 197.005 101.950 197.160 ;
        RECT 102.655 197.160 104.340 197.300 ;
        RECT 102.655 197.115 102.945 197.160 ;
        RECT 104.020 197.100 104.340 197.160 ;
        RECT 110.945 197.300 111.235 197.345 ;
        RECT 113.465 197.300 113.755 197.345 ;
        RECT 114.655 197.300 114.945 197.345 ;
        RECT 110.945 197.160 114.945 197.300 ;
        RECT 110.945 197.115 111.235 197.160 ;
        RECT 113.465 197.115 113.755 197.160 ;
        RECT 114.655 197.115 114.945 197.160 ;
        RECT 118.305 197.300 118.595 197.345 ;
        RECT 120.825 197.300 121.115 197.345 ;
        RECT 122.015 197.300 122.305 197.345 ;
        RECT 118.305 197.160 122.305 197.300 ;
        RECT 118.305 197.115 118.595 197.160 ;
        RECT 120.825 197.115 121.115 197.160 ;
        RECT 122.015 197.115 122.305 197.160 ;
        RECT 101.735 196.960 102.025 197.005 ;
        RECT 106.320 196.960 106.640 197.020 ;
        RECT 101.735 196.820 106.640 196.960 ;
        RECT 101.735 196.775 102.025 196.820 ;
        RECT 106.320 196.760 106.640 196.820 ;
        RECT 115.535 196.960 115.825 197.005 ;
        RECT 122.895 196.960 123.185 197.005 ;
        RECT 124.720 196.960 125.040 197.020 ;
        RECT 115.535 196.820 125.040 196.960 ;
        RECT 115.535 196.775 115.825 196.820 ;
        RECT 122.895 196.775 123.185 196.820 ;
        RECT 124.720 196.760 125.040 196.820 ;
        RECT 105.860 196.620 106.180 196.680 ;
        RECT 102.270 196.480 106.180 196.620 ;
        RECT 102.270 196.280 102.410 196.480 ;
        RECT 105.860 196.420 106.180 196.480 ;
        RECT 113.220 196.620 113.540 196.680 ;
        RECT 114.200 196.620 114.490 196.665 ;
        RECT 113.220 196.480 114.490 196.620 ;
        RECT 113.220 196.420 113.540 196.480 ;
        RECT 114.200 196.435 114.490 196.480 ;
        RECT 115.060 196.620 115.380 196.680 ;
        RECT 121.560 196.620 121.850 196.665 ;
        RECT 115.060 196.480 121.850 196.620 ;
        RECT 115.060 196.420 115.380 196.480 ;
        RECT 121.560 196.435 121.850 196.480 ;
        RECT 100.890 196.140 102.410 196.280 ;
        RECT 102.655 196.280 102.945 196.325 ;
        RECT 104.940 196.280 105.260 196.340 ;
        RECT 102.655 196.140 105.260 196.280 ;
        RECT 97.120 196.080 97.440 196.140 ;
        RECT 102.655 196.095 102.945 196.140 ;
        RECT 104.940 196.080 105.260 196.140 ;
        RECT 108.620 196.080 108.940 196.340 ;
        RECT 115.995 196.280 116.285 196.325 ;
        RECT 116.440 196.280 116.760 196.340 ;
        RECT 115.995 196.140 116.760 196.280 ;
        RECT 115.995 196.095 116.285 196.140 ;
        RECT 116.440 196.080 116.760 196.140 ;
        RECT 13.330 195.460 138.910 195.940 ;
        RECT 54.800 195.260 55.120 195.320 ;
        RECT 51.670 195.120 55.120 195.260 ;
        RECT 51.670 194.965 51.810 195.120 ;
        RECT 54.800 195.060 55.120 195.120 ;
        RECT 66.760 195.060 67.080 195.320 ;
        RECT 67.220 195.260 67.540 195.320 ;
        RECT 69.980 195.260 70.300 195.320 ;
        RECT 72.295 195.260 72.585 195.305 ;
        RECT 67.220 195.120 72.585 195.260 ;
        RECT 67.220 195.060 67.540 195.120 ;
        RECT 69.980 195.060 70.300 195.120 ;
        RECT 72.295 195.075 72.585 195.120 ;
        RECT 114.615 195.260 114.905 195.305 ;
        RECT 115.060 195.260 115.380 195.320 ;
        RECT 114.615 195.120 115.380 195.260 ;
        RECT 114.615 195.075 114.905 195.120 ;
        RECT 115.060 195.060 115.380 195.120 ;
        RECT 51.595 194.735 51.885 194.965 ;
        RECT 66.850 194.920 66.990 195.060 ;
        RECT 69.520 194.920 69.840 194.980 ;
        RECT 61.790 194.780 69.840 194.920 ;
        RECT 60.320 194.625 60.640 194.640 ;
        RECT 61.790 194.625 61.930 194.780 ;
        RECT 60.320 194.395 60.670 194.625 ;
        RECT 61.715 194.395 62.005 194.625 ;
        RECT 60.320 194.380 60.640 194.395 ;
        RECT 62.160 194.380 62.480 194.640 ;
        RECT 62.620 194.380 62.940 194.640 ;
        RECT 65.470 194.625 65.610 194.780 ;
        RECT 69.520 194.720 69.840 194.780 ;
        RECT 75.975 194.920 76.265 194.965 ;
        RECT 80.100 194.920 80.420 194.980 ;
        RECT 75.975 194.780 80.420 194.920 ;
        RECT 75.975 194.735 76.265 194.780 ;
        RECT 80.100 194.720 80.420 194.780 ;
        RECT 90.220 194.920 90.540 194.980 ;
        RECT 98.500 194.920 98.820 194.980 ;
        RECT 90.220 194.780 98.820 194.920 ;
        RECT 90.220 194.720 90.540 194.780 ;
        RECT 65.395 194.395 65.685 194.625 ;
        RECT 66.730 194.580 67.020 194.625 ;
        RECT 68.600 194.580 68.920 194.640 ;
        RECT 66.730 194.440 68.920 194.580 ;
        RECT 66.730 194.395 67.020 194.440 ;
        RECT 68.600 194.380 68.920 194.440 ;
        RECT 70.440 194.580 70.760 194.640 ;
        RECT 74.135 194.580 74.425 194.625 ;
        RECT 77.800 194.580 78.120 194.640 ;
        RECT 70.440 194.440 78.120 194.580 ;
        RECT 70.440 194.380 70.760 194.440 ;
        RECT 74.135 194.395 74.425 194.440 ;
        RECT 77.800 194.380 78.120 194.440 ;
        RECT 80.560 194.380 80.880 194.640 ;
        RECT 81.480 194.380 81.800 194.640 ;
        RECT 96.775 194.580 97.065 194.625 ;
        RECT 97.580 194.580 97.900 194.640 ;
        RECT 98.130 194.625 98.270 194.780 ;
        RECT 98.500 194.720 98.820 194.780 ;
        RECT 96.775 194.440 97.900 194.580 ;
        RECT 96.775 194.395 97.065 194.440 ;
        RECT 97.580 194.380 97.900 194.440 ;
        RECT 98.055 194.580 98.345 194.625 ;
        RECT 103.115 194.580 103.405 194.625 ;
        RECT 98.055 194.440 103.405 194.580 ;
        RECT 98.055 194.395 98.345 194.440 ;
        RECT 103.115 194.395 103.405 194.440 ;
        RECT 103.560 194.580 103.880 194.640 ;
        RECT 104.395 194.580 104.685 194.625 ;
        RECT 103.560 194.440 104.685 194.580 ;
        RECT 103.560 194.380 103.880 194.440 ;
        RECT 104.395 194.395 104.685 194.440 ;
        RECT 110.920 194.580 111.240 194.640 ;
        RECT 112.315 194.580 112.605 194.625 ;
        RECT 110.920 194.440 112.605 194.580 ;
        RECT 110.920 194.380 111.240 194.440 ;
        RECT 112.315 194.395 112.605 194.440 ;
        RECT 112.760 194.380 113.080 194.640 ;
        RECT 32.275 194.055 32.565 194.285 ;
        RECT 30.880 193.900 31.200 193.960 ;
        RECT 32.350 193.900 32.490 194.055 ;
        RECT 33.640 194.040 33.960 194.300 ;
        RECT 34.100 194.040 34.420 194.300 ;
        RECT 34.700 194.240 34.990 194.285 ;
        RECT 37.780 194.240 38.100 194.300 ;
        RECT 34.700 194.100 38.100 194.240 ;
        RECT 34.700 194.055 34.990 194.100 ;
        RECT 37.780 194.040 38.100 194.100 ;
        RECT 57.125 194.240 57.415 194.285 ;
        RECT 59.645 194.240 59.935 194.285 ;
        RECT 60.835 194.240 61.125 194.285 ;
        RECT 57.125 194.100 61.125 194.240 ;
        RECT 57.125 194.055 57.415 194.100 ;
        RECT 59.645 194.055 59.935 194.100 ;
        RECT 60.835 194.055 61.125 194.100 ;
        RECT 63.540 194.040 63.860 194.300 ;
        RECT 64.000 194.040 64.320 194.300 ;
        RECT 66.275 194.240 66.565 194.285 ;
        RECT 67.465 194.240 67.755 194.285 ;
        RECT 69.985 194.240 70.275 194.285 ;
        RECT 66.275 194.100 70.275 194.240 ;
        RECT 66.275 194.055 66.565 194.100 ;
        RECT 67.465 194.055 67.755 194.100 ;
        RECT 69.985 194.055 70.275 194.100 ;
        RECT 73.675 194.240 73.965 194.285 ;
        RECT 74.580 194.240 74.900 194.300 ;
        RECT 73.675 194.100 74.900 194.240 ;
        RECT 73.675 194.055 73.965 194.100 ;
        RECT 74.580 194.040 74.900 194.100 ;
        RECT 75.500 194.040 75.820 194.300 ;
        RECT 79.195 194.055 79.485 194.285 ;
        RECT 57.560 193.900 57.850 193.945 ;
        RECT 59.130 193.900 59.420 193.945 ;
        RECT 61.230 193.900 61.520 193.945 ;
        RECT 30.880 193.760 35.250 193.900 ;
        RECT 30.880 193.700 31.200 193.760 ;
        RECT 35.110 193.620 35.250 193.760 ;
        RECT 57.560 193.760 61.520 193.900 ;
        RECT 57.560 193.715 57.850 193.760 ;
        RECT 59.130 193.715 59.420 193.760 ;
        RECT 61.230 193.715 61.520 193.760 ;
        RECT 65.880 193.900 66.170 193.945 ;
        RECT 67.980 193.900 68.270 193.945 ;
        RECT 69.550 193.900 69.840 193.945 ;
        RECT 65.880 193.760 69.840 193.900 ;
        RECT 74.670 193.900 74.810 194.040 ;
        RECT 79.270 193.900 79.410 194.055 ;
        RECT 88.840 194.040 89.160 194.300 ;
        RECT 93.465 194.240 93.755 194.285 ;
        RECT 95.985 194.240 96.275 194.285 ;
        RECT 97.175 194.240 97.465 194.285 ;
        RECT 93.465 194.100 97.465 194.240 ;
        RECT 93.465 194.055 93.755 194.100 ;
        RECT 95.985 194.055 96.275 194.100 ;
        RECT 97.175 194.055 97.465 194.100 ;
        RECT 98.515 194.055 98.805 194.285 ;
        RECT 103.995 194.240 104.285 194.285 ;
        RECT 105.185 194.240 105.475 194.285 ;
        RECT 107.705 194.240 107.995 194.285 ;
        RECT 103.995 194.100 107.995 194.240 ;
        RECT 103.995 194.055 104.285 194.100 ;
        RECT 105.185 194.055 105.475 194.100 ;
        RECT 107.705 194.055 107.995 194.100 ;
        RECT 111.855 194.240 112.145 194.285 ;
        RECT 113.680 194.240 114.000 194.300 ;
        RECT 111.855 194.100 114.000 194.240 ;
        RECT 111.855 194.055 112.145 194.100 ;
        RECT 74.670 193.760 79.410 193.900 ;
        RECT 93.900 193.900 94.190 193.945 ;
        RECT 95.470 193.900 95.760 193.945 ;
        RECT 97.570 193.900 97.860 193.945 ;
        RECT 93.900 193.760 97.860 193.900 ;
        RECT 65.880 193.715 66.170 193.760 ;
        RECT 67.980 193.715 68.270 193.760 ;
        RECT 69.550 193.715 69.840 193.760 ;
        RECT 93.900 193.715 94.190 193.760 ;
        RECT 95.470 193.715 95.760 193.760 ;
        RECT 97.570 193.715 97.860 193.760 ;
        RECT 35.020 193.360 35.340 193.620 ;
        RECT 35.480 193.360 35.800 193.620 ;
        RECT 51.120 193.360 51.440 193.620 ;
        RECT 64.460 193.360 64.780 193.620 ;
        RECT 72.740 193.360 73.060 193.620 ;
        RECT 73.200 193.560 73.520 193.620 ;
        RECT 76.435 193.560 76.725 193.605 ;
        RECT 73.200 193.420 76.725 193.560 ;
        RECT 73.200 193.360 73.520 193.420 ;
        RECT 76.435 193.375 76.725 193.420 ;
        RECT 76.880 193.560 77.200 193.620 ;
        RECT 81.495 193.560 81.785 193.605 ;
        RECT 76.880 193.420 81.785 193.560 ;
        RECT 76.880 193.360 77.200 193.420 ;
        RECT 81.495 193.375 81.785 193.420 ;
        RECT 85.620 193.560 85.940 193.620 ;
        RECT 86.095 193.560 86.385 193.605 ;
        RECT 85.620 193.420 86.385 193.560 ;
        RECT 85.620 193.360 85.940 193.420 ;
        RECT 86.095 193.375 86.385 193.420 ;
        RECT 91.140 193.560 91.460 193.620 ;
        RECT 96.660 193.560 96.980 193.620 ;
        RECT 98.590 193.560 98.730 194.055 ;
        RECT 113.680 194.040 114.000 194.100 ;
        RECT 103.600 193.900 103.890 193.945 ;
        RECT 105.700 193.900 105.990 193.945 ;
        RECT 107.270 193.900 107.560 193.945 ;
        RECT 103.600 193.760 107.560 193.900 ;
        RECT 103.600 193.715 103.890 193.760 ;
        RECT 105.700 193.715 105.990 193.760 ;
        RECT 107.270 193.715 107.560 193.760 ;
        RECT 91.140 193.420 98.730 193.560 ;
        RECT 101.260 193.560 101.580 193.620 ;
        RECT 101.735 193.560 102.025 193.605 ;
        RECT 101.260 193.420 102.025 193.560 ;
        RECT 91.140 193.360 91.460 193.420 ;
        RECT 96.660 193.360 96.980 193.420 ;
        RECT 101.260 193.360 101.580 193.420 ;
        RECT 101.735 193.375 102.025 193.420 ;
        RECT 109.080 193.560 109.400 193.620 ;
        RECT 110.015 193.560 110.305 193.605 ;
        RECT 109.080 193.420 110.305 193.560 ;
        RECT 109.080 193.360 109.400 193.420 ;
        RECT 110.015 193.375 110.305 193.420 ;
        RECT 13.330 192.740 138.910 193.220 ;
        RECT 34.100 192.540 34.420 192.600 ;
        RECT 50.200 192.540 50.520 192.600 ;
        RECT 32.840 192.400 50.520 192.540 ;
        RECT 19.420 192.200 19.710 192.245 ;
        RECT 21.520 192.200 21.810 192.245 ;
        RECT 23.090 192.200 23.380 192.245 ;
        RECT 19.420 192.060 23.380 192.200 ;
        RECT 19.420 192.015 19.710 192.060 ;
        RECT 21.520 192.015 21.810 192.060 ;
        RECT 23.090 192.015 23.380 192.060 ;
        RECT 25.820 192.000 26.140 192.260 ;
        RECT 26.280 192.200 26.600 192.260 ;
        RECT 32.840 192.200 32.980 192.400 ;
        RECT 34.100 192.340 34.420 192.400 ;
        RECT 50.200 192.340 50.520 192.400 ;
        RECT 60.320 192.340 60.640 192.600 ;
        RECT 64.475 192.540 64.765 192.585 ;
        RECT 66.300 192.540 66.620 192.600 ;
        RECT 67.680 192.540 68.000 192.600 ;
        RECT 63.170 192.400 68.000 192.540 ;
        RECT 26.280 192.060 32.980 192.200 ;
        RECT 33.220 192.200 33.510 192.245 ;
        RECT 35.320 192.200 35.610 192.245 ;
        RECT 36.890 192.200 37.180 192.245 ;
        RECT 33.220 192.060 37.180 192.200 ;
        RECT 26.280 192.000 26.600 192.060 ;
        RECT 19.815 191.860 20.105 191.905 ;
        RECT 21.005 191.860 21.295 191.905 ;
        RECT 23.525 191.860 23.815 191.905 ;
        RECT 19.815 191.720 23.815 191.860 ;
        RECT 19.815 191.675 20.105 191.720 ;
        RECT 21.005 191.675 21.295 191.720 ;
        RECT 23.525 191.675 23.815 191.720 ;
        RECT 23.980 191.860 24.300 191.920 ;
        RECT 29.055 191.860 29.345 191.905 ;
        RECT 29.960 191.860 30.280 191.920 ;
        RECT 30.970 191.905 31.110 192.060 ;
        RECT 33.220 192.015 33.510 192.060 ;
        RECT 35.320 192.015 35.610 192.060 ;
        RECT 36.890 192.015 37.180 192.060 ;
        RECT 44.260 192.200 44.550 192.245 ;
        RECT 46.360 192.200 46.650 192.245 ;
        RECT 47.930 192.200 48.220 192.245 ;
        RECT 44.260 192.060 48.220 192.200 ;
        RECT 44.260 192.015 44.550 192.060 ;
        RECT 46.360 192.015 46.650 192.060 ;
        RECT 47.930 192.015 48.220 192.060 ;
        RECT 53.000 192.200 53.290 192.245 ;
        RECT 55.100 192.200 55.390 192.245 ;
        RECT 56.670 192.200 56.960 192.245 ;
        RECT 53.000 192.060 56.960 192.200 ;
        RECT 53.000 192.015 53.290 192.060 ;
        RECT 55.100 192.015 55.390 192.060 ;
        RECT 56.670 192.015 56.960 192.060 ;
        RECT 31.340 191.905 31.660 191.920 ;
        RECT 23.980 191.720 30.280 191.860 ;
        RECT 23.980 191.660 24.300 191.720 ;
        RECT 29.055 191.675 29.345 191.720 ;
        RECT 29.960 191.660 30.280 191.720 ;
        RECT 30.895 191.675 31.185 191.905 ;
        RECT 31.340 191.675 31.770 191.905 ;
        RECT 33.615 191.860 33.905 191.905 ;
        RECT 34.805 191.860 35.095 191.905 ;
        RECT 37.325 191.860 37.615 191.905 ;
        RECT 33.615 191.720 37.615 191.860 ;
        RECT 33.615 191.675 33.905 191.720 ;
        RECT 34.805 191.675 35.095 191.720 ;
        RECT 37.325 191.675 37.615 191.720 ;
        RECT 44.655 191.860 44.945 191.905 ;
        RECT 45.845 191.860 46.135 191.905 ;
        RECT 48.365 191.860 48.655 191.905 ;
        RECT 44.655 191.720 48.655 191.860 ;
        RECT 44.655 191.675 44.945 191.720 ;
        RECT 45.845 191.675 46.135 191.720 ;
        RECT 48.365 191.675 48.655 191.720 ;
        RECT 53.395 191.860 53.685 191.905 ;
        RECT 54.585 191.860 54.875 191.905 ;
        RECT 57.105 191.860 57.395 191.905 ;
        RECT 53.395 191.720 57.395 191.860 ;
        RECT 53.395 191.675 53.685 191.720 ;
        RECT 54.585 191.675 54.875 191.720 ;
        RECT 57.105 191.675 57.395 191.720 ;
        RECT 61.255 191.860 61.545 191.905 ;
        RECT 62.160 191.860 62.480 191.920 ;
        RECT 61.255 191.720 62.480 191.860 ;
        RECT 61.255 191.675 61.545 191.720 ;
        RECT 31.340 191.660 31.660 191.675 ;
        RECT 62.160 191.660 62.480 191.720 ;
        RECT 17.540 191.520 17.860 191.580 ;
        RECT 18.935 191.520 19.225 191.565 ;
        RECT 32.735 191.520 33.025 191.565 ;
        RECT 17.540 191.380 19.225 191.520 ;
        RECT 17.540 191.320 17.860 191.380 ;
        RECT 18.935 191.335 19.225 191.380 ;
        RECT 30.970 191.380 33.025 191.520 ;
        RECT 30.970 191.240 31.110 191.380 ;
        RECT 32.735 191.335 33.025 191.380 ;
        RECT 34.070 191.520 34.360 191.565 ;
        RECT 35.480 191.520 35.800 191.580 ;
        RECT 34.070 191.380 35.800 191.520 ;
        RECT 34.070 191.335 34.360 191.380 ;
        RECT 35.480 191.320 35.800 191.380 ;
        RECT 43.775 191.520 44.065 191.565 ;
        RECT 49.280 191.520 49.600 191.580 ;
        RECT 52.515 191.520 52.805 191.565 ;
        RECT 43.775 191.380 52.805 191.520 ;
        RECT 43.775 191.335 44.065 191.380 ;
        RECT 49.280 191.320 49.600 191.380 ;
        RECT 52.515 191.335 52.805 191.380 ;
        RECT 61.715 191.520 62.005 191.565 ;
        RECT 63.170 191.520 63.310 192.400 ;
        RECT 64.475 192.355 64.765 192.400 ;
        RECT 66.300 192.340 66.620 192.400 ;
        RECT 67.680 192.340 68.000 192.400 ;
        RECT 68.600 192.340 68.920 192.600 ;
        RECT 69.980 192.540 70.300 192.600 ;
        RECT 74.135 192.540 74.425 192.585 ;
        RECT 76.420 192.540 76.740 192.600 ;
        RECT 69.980 192.400 76.740 192.540 ;
        RECT 69.980 192.340 70.300 192.400 ;
        RECT 74.135 192.355 74.425 192.400 ;
        RECT 76.420 192.340 76.740 192.400 ;
        RECT 76.895 192.540 77.185 192.585 ;
        RECT 77.800 192.540 78.120 192.600 ;
        RECT 76.895 192.400 78.120 192.540 ;
        RECT 76.895 192.355 77.185 192.400 ;
        RECT 77.800 192.340 78.120 192.400 ;
        RECT 91.600 192.540 91.920 192.600 ;
        RECT 101.275 192.540 101.565 192.585 ;
        RECT 91.600 192.400 96.890 192.540 ;
        RECT 91.600 192.340 91.920 192.400 ;
        RECT 64.920 192.200 65.240 192.260 ;
        RECT 65.840 192.200 66.160 192.260 ;
        RECT 64.090 192.060 66.160 192.200 ;
        RECT 64.090 191.565 64.230 192.060 ;
        RECT 64.920 192.000 65.240 192.060 ;
        RECT 65.840 192.000 66.160 192.060 ;
        RECT 68.140 192.200 68.460 192.260 ;
        RECT 69.075 192.200 69.365 192.245 ;
        RECT 68.140 192.060 69.365 192.200 ;
        RECT 68.140 192.000 68.460 192.060 ;
        RECT 69.075 192.015 69.365 192.060 ;
        RECT 70.455 192.200 70.745 192.245 ;
        RECT 81.020 192.200 81.340 192.260 ;
        RECT 70.455 192.060 81.340 192.200 ;
        RECT 70.455 192.015 70.745 192.060 ;
        RECT 81.020 192.000 81.340 192.060 ;
        RECT 81.940 192.200 82.230 192.245 ;
        RECT 83.510 192.200 83.800 192.245 ;
        RECT 85.610 192.200 85.900 192.245 ;
        RECT 81.940 192.060 85.900 192.200 ;
        RECT 81.940 192.015 82.230 192.060 ;
        RECT 83.510 192.015 83.800 192.060 ;
        RECT 85.610 192.015 85.900 192.060 ;
        RECT 90.720 192.200 91.010 192.245 ;
        RECT 92.820 192.200 93.110 192.245 ;
        RECT 94.390 192.200 94.680 192.245 ;
        RECT 90.720 192.060 94.680 192.200 ;
        RECT 90.720 192.015 91.010 192.060 ;
        RECT 92.820 192.015 93.110 192.060 ;
        RECT 94.390 192.015 94.680 192.060 ;
        RECT 64.460 191.860 64.780 191.920 ;
        RECT 65.395 191.860 65.685 191.905 ;
        RECT 73.200 191.860 73.520 191.920 ;
        RECT 76.880 191.860 77.200 191.920 ;
        RECT 64.460 191.720 65.685 191.860 ;
        RECT 64.460 191.660 64.780 191.720 ;
        RECT 65.395 191.675 65.685 191.720 ;
        RECT 70.070 191.720 73.520 191.860 ;
        RECT 61.715 191.380 63.310 191.520 ;
        RECT 61.715 191.335 62.005 191.380 ;
        RECT 64.015 191.335 64.305 191.565 ;
        RECT 64.975 191.490 65.265 191.535 ;
        RECT 68.140 191.520 68.460 191.580 ;
        RECT 69.520 191.520 69.840 191.580 ;
        RECT 70.070 191.565 70.210 191.720 ;
        RECT 73.200 191.660 73.520 191.720 ;
        RECT 74.210 191.720 77.200 191.860 ;
        RECT 64.975 191.350 65.610 191.490 ;
        RECT 20.300 191.225 20.620 191.240 ;
        RECT 20.270 190.995 20.620 191.225 ;
        RECT 20.300 190.980 20.620 190.995 ;
        RECT 30.880 190.980 31.200 191.240 ;
        RECT 33.640 191.180 33.960 191.240 ;
        RECT 31.890 191.040 33.960 191.180 ;
        RECT 20.760 190.840 21.080 190.900 ;
        RECT 30.435 190.840 30.725 190.885 ;
        RECT 31.890 190.840 32.030 191.040 ;
        RECT 33.640 190.980 33.960 191.040 ;
        RECT 42.840 191.180 43.160 191.240 ;
        RECT 45.000 191.180 45.290 191.225 ;
        RECT 42.840 191.040 45.290 191.180 ;
        RECT 42.840 190.980 43.160 191.040 ;
        RECT 45.000 190.995 45.290 191.040 ;
        RECT 51.580 191.180 51.900 191.240 ;
        RECT 53.740 191.180 54.030 191.225 ;
        RECT 51.580 191.040 54.030 191.180 ;
        RECT 51.580 190.980 51.900 191.040 ;
        RECT 53.740 190.995 54.030 191.040 ;
        RECT 63.080 190.980 63.400 191.240 ;
        RECT 63.540 190.980 63.860 191.240 ;
        RECT 20.760 190.700 32.030 190.840 ;
        RECT 20.760 190.640 21.080 190.700 ;
        RECT 30.435 190.655 30.725 190.700 ;
        RECT 32.260 190.640 32.580 190.900 ;
        RECT 39.620 190.640 39.940 190.900 ;
        RECT 41.000 190.840 41.320 190.900 ;
        RECT 50.675 190.840 50.965 190.885 ;
        RECT 52.960 190.840 53.280 190.900 ;
        RECT 41.000 190.700 53.280 190.840 ;
        RECT 41.000 190.640 41.320 190.700 ;
        RECT 50.675 190.655 50.965 190.700 ;
        RECT 52.960 190.640 53.280 190.700 ;
        RECT 59.415 190.840 59.705 190.885 ;
        RECT 64.090 190.840 64.230 191.335 ;
        RECT 64.975 191.305 65.265 191.350 ;
        RECT 59.415 190.700 64.230 190.840 ;
        RECT 65.470 190.840 65.610 191.350 ;
        RECT 68.140 191.380 69.840 191.520 ;
        RECT 68.140 191.320 68.460 191.380 ;
        RECT 69.520 191.320 69.840 191.380 ;
        RECT 69.995 191.335 70.285 191.565 ;
        RECT 70.440 191.520 70.760 191.580 ;
        RECT 70.915 191.520 71.205 191.565 ;
        RECT 70.440 191.380 71.205 191.520 ;
        RECT 70.440 191.320 70.760 191.380 ;
        RECT 70.915 191.335 71.205 191.380 ;
        RECT 71.360 191.320 71.680 191.580 ;
        RECT 72.295 191.520 72.585 191.565 ;
        RECT 72.740 191.520 73.060 191.580 ;
        RECT 74.210 191.565 74.350 191.720 ;
        RECT 76.880 191.660 77.200 191.720 ;
        RECT 81.505 191.860 81.795 191.905 ;
        RECT 84.025 191.860 84.315 191.905 ;
        RECT 85.215 191.860 85.505 191.905 ;
        RECT 90.220 191.860 90.540 191.920 ;
        RECT 81.505 191.720 85.505 191.860 ;
        RECT 81.505 191.675 81.795 191.720 ;
        RECT 84.025 191.675 84.315 191.720 ;
        RECT 85.215 191.675 85.505 191.720 ;
        RECT 86.170 191.720 90.540 191.860 ;
        RECT 86.170 191.580 86.310 191.720 ;
        RECT 90.220 191.660 90.540 191.720 ;
        RECT 91.115 191.860 91.405 191.905 ;
        RECT 92.305 191.860 92.595 191.905 ;
        RECT 94.825 191.860 95.115 191.905 ;
        RECT 91.115 191.720 95.115 191.860 ;
        RECT 96.750 191.860 96.890 192.400 ;
        RECT 100.430 192.400 101.565 192.540 ;
        RECT 100.430 191.905 100.570 192.400 ;
        RECT 101.275 192.355 101.565 192.400 ;
        RECT 103.560 192.540 103.880 192.600 ;
        RECT 104.035 192.540 104.325 192.585 ;
        RECT 103.560 192.400 104.325 192.540 ;
        RECT 103.560 192.340 103.880 192.400 ;
        RECT 104.035 192.355 104.325 192.400 ;
        RECT 105.860 192.540 106.180 192.600 ;
        RECT 105.860 192.400 109.770 192.540 ;
        RECT 105.860 192.340 106.180 192.400 ;
        RECT 106.320 192.200 106.640 192.260 ;
        RECT 107.715 192.200 108.005 192.245 ;
        RECT 106.320 192.060 108.005 192.200 ;
        RECT 109.630 192.200 109.770 192.400 ;
        RECT 113.220 192.340 113.540 192.600 ;
        RECT 115.520 192.540 115.840 192.600 ;
        RECT 113.770 192.400 115.840 192.540 ;
        RECT 113.770 192.200 113.910 192.400 ;
        RECT 115.520 192.340 115.840 192.400 ;
        RECT 109.630 192.060 113.910 192.200 ;
        RECT 114.140 192.200 114.460 192.260 ;
        RECT 118.740 192.200 119.060 192.260 ;
        RECT 136.235 192.200 136.525 192.245 ;
        RECT 114.140 192.060 118.510 192.200 ;
        RECT 106.320 192.000 106.640 192.060 ;
        RECT 107.715 192.015 108.005 192.060 ;
        RECT 114.140 192.000 114.460 192.060 ;
        RECT 100.355 191.860 100.645 191.905 ;
        RECT 101.735 191.860 102.025 191.905 ;
        RECT 103.560 191.860 103.880 191.920 ;
        RECT 110.460 191.860 110.780 191.920 ;
        RECT 112.760 191.860 113.080 191.920 ;
        RECT 116.455 191.860 116.745 191.905 ;
        RECT 96.750 191.720 100.645 191.860 ;
        RECT 91.115 191.675 91.405 191.720 ;
        RECT 92.305 191.675 92.595 191.720 ;
        RECT 94.825 191.675 95.115 191.720 ;
        RECT 100.355 191.675 100.645 191.720 ;
        RECT 100.890 191.720 103.880 191.860 ;
        RECT 72.295 191.380 73.060 191.520 ;
        RECT 72.295 191.335 72.585 191.380 ;
        RECT 72.740 191.320 73.060 191.380 ;
        RECT 74.135 191.335 74.425 191.565 ;
        RECT 74.580 191.320 74.900 191.580 ;
        RECT 76.420 191.320 76.740 191.580 ;
        RECT 77.355 191.335 77.645 191.565 ;
        RECT 84.815 191.520 85.105 191.565 ;
        RECT 85.620 191.520 85.940 191.580 ;
        RECT 84.815 191.380 85.940 191.520 ;
        RECT 84.815 191.335 85.105 191.380 ;
        RECT 73.660 191.180 73.980 191.240 ;
        RECT 77.430 191.180 77.570 191.335 ;
        RECT 85.620 191.320 85.940 191.380 ;
        RECT 86.080 191.320 86.400 191.580 ;
        RECT 86.555 191.335 86.845 191.565 ;
        RECT 90.680 191.520 91.000 191.580 ;
        RECT 91.515 191.520 91.805 191.565 ;
        RECT 90.680 191.380 91.805 191.520 ;
        RECT 73.660 191.040 77.570 191.180 ;
        RECT 73.660 190.980 73.980 191.040 ;
        RECT 74.580 190.840 74.900 190.900 ;
        RECT 65.470 190.700 74.900 190.840 ;
        RECT 59.415 190.655 59.705 190.700 ;
        RECT 74.580 190.640 74.900 190.700 ;
        RECT 75.975 190.840 76.265 190.885 ;
        RECT 76.420 190.840 76.740 190.900 ;
        RECT 75.975 190.700 76.740 190.840 ;
        RECT 75.975 190.655 76.265 190.700 ;
        RECT 76.420 190.640 76.740 190.700 ;
        RECT 79.195 190.840 79.485 190.885 ;
        RECT 80.560 190.840 80.880 190.900 ;
        RECT 86.630 190.840 86.770 191.335 ;
        RECT 90.680 191.320 91.000 191.380 ;
        RECT 91.515 191.335 91.805 191.380 ;
        RECT 96.660 191.520 96.980 191.580 ;
        RECT 100.890 191.520 101.030 191.720 ;
        RECT 101.735 191.675 102.025 191.720 ;
        RECT 103.560 191.660 103.880 191.720 ;
        RECT 106.410 191.720 110.780 191.860 ;
        RECT 96.660 191.380 101.030 191.520 ;
        RECT 101.275 191.520 101.565 191.565 ;
        RECT 102.640 191.520 102.960 191.580 ;
        RECT 101.275 191.380 102.960 191.520 ;
        RECT 96.660 191.320 96.980 191.380 ;
        RECT 101.275 191.335 101.565 191.380 ;
        RECT 102.640 191.320 102.960 191.380 ;
        RECT 104.940 191.320 105.260 191.580 ;
        RECT 106.410 191.565 106.550 191.720 ;
        RECT 110.460 191.660 110.780 191.720 ;
        RECT 112.390 191.720 116.745 191.860 ;
        RECT 105.415 191.335 105.705 191.565 ;
        RECT 106.335 191.335 106.625 191.565 ;
        RECT 100.800 191.180 101.120 191.240 ;
        RECT 97.210 191.040 101.120 191.180 ;
        RECT 79.195 190.700 86.770 190.840 ;
        RECT 87.920 190.840 88.240 190.900 ;
        RECT 89.775 190.840 90.065 190.885 ;
        RECT 87.920 190.700 90.065 190.840 ;
        RECT 79.195 190.655 79.485 190.700 ;
        RECT 80.560 190.640 80.880 190.700 ;
        RECT 87.920 190.640 88.240 190.700 ;
        RECT 89.775 190.655 90.065 190.700 ;
        RECT 92.980 190.840 93.300 190.900 ;
        RECT 97.210 190.885 97.350 191.040 ;
        RECT 100.800 190.980 101.120 191.040 ;
        RECT 97.135 190.840 97.425 190.885 ;
        RECT 92.980 190.700 97.425 190.840 ;
        RECT 92.980 190.640 93.300 190.700 ;
        RECT 97.135 190.655 97.425 190.700 ;
        RECT 97.580 190.640 97.900 190.900 ;
        RECT 103.100 190.640 103.420 190.900 ;
        RECT 105.030 190.840 105.170 191.320 ;
        RECT 105.490 191.180 105.630 191.335 ;
        RECT 106.780 191.320 107.100 191.580 ;
        RECT 107.715 191.335 108.005 191.565 ;
        RECT 108.620 191.520 108.940 191.580 ;
        RECT 112.390 191.565 112.530 191.720 ;
        RECT 112.760 191.660 113.080 191.720 ;
        RECT 116.455 191.675 116.745 191.720 ;
        RECT 110.015 191.520 110.305 191.565 ;
        RECT 108.620 191.380 110.305 191.520 ;
        RECT 107.790 191.180 107.930 191.335 ;
        RECT 108.620 191.320 108.940 191.380 ;
        RECT 110.015 191.335 110.305 191.380 ;
        RECT 112.315 191.335 112.605 191.565 ;
        RECT 113.680 191.320 114.000 191.580 ;
        RECT 114.140 191.520 114.460 191.580 ;
        RECT 115.535 191.520 115.825 191.565 ;
        RECT 114.140 191.380 115.825 191.520 ;
        RECT 114.140 191.320 114.460 191.380 ;
        RECT 115.535 191.335 115.825 191.380 ;
        RECT 115.980 191.320 116.300 191.580 ;
        RECT 116.900 191.320 117.220 191.580 ;
        RECT 118.370 191.565 118.510 192.060 ;
        RECT 118.740 192.060 136.525 192.200 ;
        RECT 118.740 192.000 119.060 192.060 ;
        RECT 136.235 192.015 136.525 192.060 ;
        RECT 117.375 191.335 117.665 191.565 ;
        RECT 118.295 191.335 118.585 191.565 ;
        RECT 109.080 191.180 109.400 191.240 ;
        RECT 110.920 191.225 111.240 191.240 ;
        RECT 110.705 191.180 111.240 191.225 ;
        RECT 105.490 191.040 109.400 191.180 ;
        RECT 109.080 190.980 109.400 191.040 ;
        RECT 109.630 191.040 111.240 191.180 ;
        RECT 109.630 190.840 109.770 191.040 ;
        RECT 110.705 190.995 111.240 191.040 ;
        RECT 111.395 190.995 111.685 191.225 ;
        RECT 110.920 190.980 111.240 190.995 ;
        RECT 105.030 190.700 109.770 190.840 ;
        RECT 111.470 190.840 111.610 190.995 ;
        RECT 111.840 190.980 112.160 191.240 ;
        RECT 113.770 191.180 113.910 191.320 ;
        RECT 114.615 191.180 114.905 191.225 ;
        RECT 113.770 191.040 114.905 191.180 ;
        RECT 114.615 190.995 114.905 191.040 ;
        RECT 116.440 191.180 116.760 191.240 ;
        RECT 117.450 191.180 117.590 191.335 ;
        RECT 133.920 191.320 134.240 191.580 ;
        RECT 137.140 191.320 137.460 191.580 ;
        RECT 116.440 191.040 117.590 191.180 ;
        RECT 116.440 190.980 116.760 191.040 ;
        RECT 113.680 190.840 114.000 190.900 ;
        RECT 111.470 190.700 114.000 190.840 ;
        RECT 113.680 190.640 114.000 190.700 ;
        RECT 117.360 190.640 117.680 190.900 ;
        RECT 134.855 190.840 135.145 190.885 ;
        RECT 135.760 190.840 136.080 190.900 ;
        RECT 134.855 190.700 136.080 190.840 ;
        RECT 134.855 190.655 135.145 190.700 ;
        RECT 135.760 190.640 136.080 190.700 ;
        RECT 13.330 190.020 138.910 190.500 ;
        RECT 20.300 189.620 20.620 189.880 ;
        RECT 20.760 189.820 21.080 189.880 ;
        RECT 22.155 189.820 22.445 189.865 ;
        RECT 32.720 189.820 33.040 189.880 ;
        RECT 20.760 189.680 22.445 189.820 ;
        RECT 20.760 189.620 21.080 189.680 ;
        RECT 22.155 189.635 22.445 189.680 ;
        RECT 28.670 189.680 33.040 189.820 ;
        RECT 28.670 189.525 28.810 189.680 ;
        RECT 32.720 189.620 33.040 189.680 ;
        RECT 34.100 189.820 34.420 189.880 ;
        RECT 34.100 189.680 41.690 189.820 ;
        RECT 34.100 189.620 34.420 189.680 ;
        RECT 28.595 189.295 28.885 189.525 ;
        RECT 29.595 189.480 29.885 189.525 ;
        RECT 29.130 189.340 29.885 189.480 ;
        RECT 21.110 189.140 21.400 189.185 ;
        RECT 21.110 189.000 24.210 189.140 ;
        RECT 21.110 188.955 21.400 189.000 ;
        RECT 21.680 188.600 22.000 188.860 ;
        RECT 23.520 188.600 23.840 188.860 ;
        RECT 24.070 188.845 24.210 189.000 ;
        RECT 25.820 188.940 26.140 189.200 ;
        RECT 29.130 189.140 29.270 189.340 ;
        RECT 29.595 189.295 29.885 189.340 ;
        RECT 31.800 189.280 32.120 189.540 ;
        RECT 41.000 189.480 41.320 189.540 ;
        RECT 40.630 189.340 41.320 189.480 ;
        RECT 41.550 189.480 41.690 189.680 ;
        RECT 42.840 189.620 43.160 189.880 ;
        RECT 65.840 189.820 66.160 189.880 ;
        RECT 73.660 189.820 73.980 189.880 ;
        RECT 43.390 189.680 50.890 189.820 ;
        RECT 43.390 189.480 43.530 189.680 ;
        RECT 41.550 189.340 43.530 189.480 ;
        RECT 44.235 189.480 44.525 189.525 ;
        RECT 47.440 189.480 47.760 189.540 ;
        RECT 44.235 189.340 47.760 189.480 ;
        RECT 26.830 189.000 29.270 189.140 ;
        RECT 31.890 189.130 32.030 189.280 ;
        RECT 40.630 189.185 40.770 189.340 ;
        RECT 41.000 189.280 41.320 189.340 ;
        RECT 44.235 189.295 44.525 189.340 ;
        RECT 47.440 189.280 47.760 189.340 ;
        RECT 50.750 189.200 50.890 189.680 ;
        RECT 65.840 189.680 73.980 189.820 ;
        RECT 65.840 189.620 66.160 189.680 ;
        RECT 73.660 189.620 73.980 189.680 ;
        RECT 81.480 189.820 81.800 189.880 ;
        RECT 82.415 189.820 82.705 189.865 ;
        RECT 81.480 189.680 82.705 189.820 ;
        RECT 81.480 189.620 81.800 189.680 ;
        RECT 82.415 189.635 82.705 189.680 ;
        RECT 86.555 189.820 86.845 189.865 ;
        RECT 88.840 189.820 89.160 189.880 ;
        RECT 97.135 189.820 97.425 189.865 ;
        RECT 86.555 189.680 89.160 189.820 ;
        RECT 86.555 189.635 86.845 189.680 ;
        RECT 88.840 189.620 89.160 189.680 ;
        RECT 93.530 189.680 97.425 189.820 ;
        RECT 51.120 189.480 51.440 189.540 ;
        RECT 51.595 189.480 51.885 189.525 ;
        RECT 51.120 189.340 51.885 189.480 ;
        RECT 51.120 189.280 51.440 189.340 ;
        RECT 51.595 189.295 51.885 189.340 ;
        RECT 68.615 189.480 68.905 189.525 ;
        RECT 69.980 189.480 70.300 189.540 ;
        RECT 68.615 189.340 70.300 189.480 ;
        RECT 68.615 189.295 68.905 189.340 ;
        RECT 69.980 189.280 70.300 189.340 ;
        RECT 76.850 189.480 77.140 189.525 ;
        RECT 77.340 189.480 77.660 189.540 ;
        RECT 93.530 189.525 93.670 189.680 ;
        RECT 97.135 189.635 97.425 189.680 ;
        RECT 98.040 189.820 98.360 189.880 ;
        RECT 98.515 189.820 98.805 189.865 ;
        RECT 111.065 189.820 111.355 189.865 ;
        RECT 111.840 189.820 112.160 189.880 ;
        RECT 114.155 189.820 114.445 189.865 ;
        RECT 117.360 189.820 117.680 189.880 ;
        RECT 98.040 189.680 98.805 189.820 ;
        RECT 98.040 189.620 98.360 189.680 ;
        RECT 98.515 189.635 98.805 189.680 ;
        RECT 105.490 189.680 108.850 189.820 ;
        RECT 93.900 189.525 94.220 189.540 ;
        RECT 93.455 189.480 93.745 189.525 ;
        RECT 76.850 189.340 77.660 189.480 ;
        RECT 76.850 189.295 77.140 189.340 ;
        RECT 77.340 189.280 77.660 189.340 ;
        RECT 88.930 189.340 93.745 189.480 ;
        RECT 32.230 189.130 32.520 189.185 ;
        RECT 26.830 188.860 26.970 189.000 ;
        RECT 31.890 188.990 32.520 189.130 ;
        RECT 32.230 188.955 32.520 188.990 ;
        RECT 40.555 188.955 40.845 189.185 ;
        RECT 44.695 189.140 44.985 189.185 ;
        RECT 46.980 189.140 47.300 189.200 ;
        RECT 44.695 189.000 47.300 189.140 ;
        RECT 44.695 188.955 44.985 189.000 ;
        RECT 46.980 188.940 47.300 189.000 ;
        RECT 50.200 188.940 50.520 189.200 ;
        RECT 50.660 188.940 50.980 189.200 ;
        RECT 64.475 188.955 64.765 189.185 ;
        RECT 67.235 188.955 67.525 189.185 ;
        RECT 23.995 188.615 24.285 188.845 ;
        RECT 26.295 188.800 26.585 188.845 ;
        RECT 26.740 188.800 27.060 188.860 ;
        RECT 26.295 188.660 27.060 188.800 ;
        RECT 26.295 188.615 26.585 188.660 ;
        RECT 26.740 188.600 27.060 188.660 ;
        RECT 30.880 188.600 31.200 188.860 ;
        RECT 31.775 188.800 32.065 188.845 ;
        RECT 32.965 188.800 33.255 188.845 ;
        RECT 35.485 188.800 35.775 188.845 ;
        RECT 31.775 188.660 35.775 188.800 ;
        RECT 31.775 188.615 32.065 188.660 ;
        RECT 32.965 188.615 33.255 188.660 ;
        RECT 35.485 188.615 35.775 188.660 ;
        RECT 41.015 188.800 41.305 188.845 ;
        RECT 41.920 188.800 42.240 188.860 ;
        RECT 41.015 188.660 42.240 188.800 ;
        RECT 41.015 188.615 41.305 188.660 ;
        RECT 41.920 188.600 42.240 188.660 ;
        RECT 42.395 188.800 42.685 188.845 ;
        RECT 43.650 188.800 43.940 188.845 ;
        RECT 42.395 188.660 43.940 188.800 ;
        RECT 42.395 188.615 42.685 188.660 ;
        RECT 43.650 188.615 43.940 188.660 ;
        RECT 46.075 188.800 46.365 188.845 ;
        RECT 46.520 188.800 46.840 188.860 ;
        RECT 63.080 188.800 63.400 188.860 ;
        RECT 46.075 188.660 63.400 188.800 ;
        RECT 46.075 188.615 46.365 188.660 ;
        RECT 46.520 188.600 46.840 188.660 ;
        RECT 63.080 188.600 63.400 188.660 ;
        RECT 17.540 188.460 17.860 188.520 ;
        RECT 30.970 188.460 31.110 188.600 ;
        RECT 17.540 188.320 31.110 188.460 ;
        RECT 31.380 188.460 31.670 188.505 ;
        RECT 33.480 188.460 33.770 188.505 ;
        RECT 35.050 188.460 35.340 188.505 ;
        RECT 31.380 188.320 35.340 188.460 ;
        RECT 17.540 188.260 17.860 188.320 ;
        RECT 31.380 188.275 31.670 188.320 ;
        RECT 33.480 188.275 33.770 188.320 ;
        RECT 35.050 188.275 35.340 188.320 ;
        RECT 51.580 188.260 51.900 188.520 ;
        RECT 64.550 188.460 64.690 188.955 ;
        RECT 64.920 188.800 65.240 188.860 ;
        RECT 66.775 188.800 67.065 188.845 ;
        RECT 64.920 188.660 67.065 188.800 ;
        RECT 67.310 188.800 67.450 188.955 ;
        RECT 67.680 188.940 68.000 189.200 ;
        RECT 87.920 188.940 88.240 189.200 ;
        RECT 88.380 188.940 88.700 189.200 ;
        RECT 88.930 189.185 89.070 189.340 ;
        RECT 93.455 189.295 93.745 189.340 ;
        RECT 93.900 189.295 94.330 189.525 ;
        RECT 97.580 189.480 97.900 189.540 ;
        RECT 99.895 189.480 100.185 189.525 ;
        RECT 97.580 189.340 100.185 189.480 ;
        RECT 93.900 189.280 94.220 189.295 ;
        RECT 97.580 189.280 97.900 189.340 ;
        RECT 99.895 189.295 100.185 189.340 ;
        RECT 100.800 189.480 101.120 189.540 ;
        RECT 105.490 189.480 105.630 189.680 ;
        RECT 100.800 189.340 105.630 189.480 ;
        RECT 100.800 189.280 101.120 189.340 ;
        RECT 88.855 188.955 89.145 189.185 ;
        RECT 89.775 189.140 90.065 189.185 ;
        RECT 99.420 189.140 99.740 189.200 ;
        RECT 89.775 189.000 91.370 189.140 ;
        RECT 89.775 188.955 90.065 189.000 ;
        RECT 68.140 188.800 68.460 188.860 ;
        RECT 75.515 188.800 75.805 188.845 ;
        RECT 67.310 188.660 67.910 188.800 ;
        RECT 64.920 188.600 65.240 188.660 ;
        RECT 66.775 188.615 67.065 188.660 ;
        RECT 65.395 188.460 65.685 188.505 ;
        RECT 64.550 188.320 65.685 188.460 ;
        RECT 67.770 188.460 67.910 188.660 ;
        RECT 68.140 188.660 75.805 188.800 ;
        RECT 68.140 188.600 68.460 188.660 ;
        RECT 75.515 188.615 75.805 188.660 ;
        RECT 76.395 188.800 76.685 188.845 ;
        RECT 77.585 188.800 77.875 188.845 ;
        RECT 80.105 188.800 80.395 188.845 ;
        RECT 76.395 188.660 80.395 188.800 ;
        RECT 76.395 188.615 76.685 188.660 ;
        RECT 77.585 188.615 77.875 188.660 ;
        RECT 80.105 188.615 80.395 188.660 ;
        RECT 85.620 188.800 85.940 188.860 ;
        RECT 88.930 188.800 89.070 188.955 ;
        RECT 91.230 188.860 91.370 189.000 ;
        RECT 94.910 189.000 99.740 189.140 ;
        RECT 85.620 188.660 89.070 188.800 ;
        RECT 91.140 188.800 91.460 188.860 ;
        RECT 91.615 188.800 91.905 188.845 ;
        RECT 91.140 188.660 91.905 188.800 ;
        RECT 85.620 188.600 85.940 188.660 ;
        RECT 91.140 188.600 91.460 188.660 ;
        RECT 91.615 188.615 91.905 188.660 ;
        RECT 69.060 188.460 69.380 188.520 ;
        RECT 67.770 188.320 69.380 188.460 ;
        RECT 65.395 188.275 65.685 188.320 ;
        RECT 69.060 188.260 69.380 188.320 ;
        RECT 76.000 188.460 76.290 188.505 ;
        RECT 78.100 188.460 78.390 188.505 ;
        RECT 79.670 188.460 79.960 188.505 ;
        RECT 76.000 188.320 79.960 188.460 ;
        RECT 76.000 188.275 76.290 188.320 ;
        RECT 78.100 188.275 78.390 188.320 ;
        RECT 79.670 188.275 79.960 188.320 ;
        RECT 25.820 188.120 26.140 188.180 ;
        RECT 29.515 188.120 29.805 188.165 ;
        RECT 25.820 187.980 29.805 188.120 ;
        RECT 25.820 187.920 26.140 187.980 ;
        RECT 29.515 187.935 29.805 187.980 ;
        RECT 30.435 188.120 30.725 188.165 ;
        RECT 30.880 188.120 31.200 188.180 ;
        RECT 30.435 187.980 31.200 188.120 ;
        RECT 30.435 187.935 30.725 187.980 ;
        RECT 30.880 187.920 31.200 187.980 ;
        RECT 32.260 188.120 32.580 188.180 ;
        RECT 34.560 188.120 34.880 188.180 ;
        RECT 37.795 188.120 38.085 188.165 ;
        RECT 32.260 187.980 38.085 188.120 ;
        RECT 32.260 187.920 32.580 187.980 ;
        RECT 34.560 187.920 34.880 187.980 ;
        RECT 37.795 187.935 38.085 187.980 ;
        RECT 64.015 188.120 64.305 188.165 ;
        RECT 66.300 188.120 66.620 188.180 ;
        RECT 64.015 187.980 66.620 188.120 ;
        RECT 64.015 187.935 64.305 187.980 ;
        RECT 66.300 187.920 66.620 187.980 ;
        RECT 67.220 187.920 67.540 188.180 ;
        RECT 67.680 188.120 68.000 188.180 ;
        RECT 69.535 188.120 69.825 188.165 ;
        RECT 67.680 187.980 69.825 188.120 ;
        RECT 67.680 187.920 68.000 187.980 ;
        RECT 69.535 187.935 69.825 187.980 ;
        RECT 76.880 188.120 77.200 188.180 ;
        RECT 85.160 188.120 85.480 188.180 ;
        RECT 76.880 187.980 85.480 188.120 ;
        RECT 91.690 188.120 91.830 188.615 ;
        RECT 92.980 188.600 93.300 188.860 ;
        RECT 94.910 188.505 95.050 189.000 ;
        RECT 99.420 188.940 99.740 189.000 ;
        RECT 100.355 188.955 100.645 189.185 ;
        RECT 95.740 188.800 96.060 188.860 ;
        RECT 100.430 188.800 100.570 188.955 ;
        RECT 101.260 188.940 101.580 189.200 ;
        RECT 102.640 188.940 102.960 189.200 ;
        RECT 103.560 189.140 103.880 189.200 ;
        RECT 104.035 189.140 104.325 189.185 ;
        RECT 103.560 189.000 104.325 189.140 ;
        RECT 103.560 188.940 103.880 189.000 ;
        RECT 104.035 188.955 104.325 189.000 ;
        RECT 104.480 188.940 104.800 189.200 ;
        RECT 105.490 189.185 105.630 189.340 ;
        RECT 105.860 189.480 106.180 189.540 ;
        RECT 108.710 189.525 108.850 189.680 ;
        RECT 111.065 189.680 117.680 189.820 ;
        RECT 111.065 189.635 111.355 189.680 ;
        RECT 111.840 189.620 112.160 189.680 ;
        RECT 114.155 189.635 114.445 189.680 ;
        RECT 117.360 189.620 117.680 189.680 ;
        RECT 131.635 189.635 131.925 189.865 ;
        RECT 106.335 189.480 106.625 189.525 ;
        RECT 105.860 189.340 106.625 189.480 ;
        RECT 105.860 189.280 106.180 189.340 ;
        RECT 106.335 189.295 106.625 189.340 ;
        RECT 107.485 189.310 107.775 189.355 ;
        RECT 105.415 188.955 105.705 189.185 ;
        RECT 107.485 189.140 107.850 189.310 ;
        RECT 108.635 189.295 108.925 189.525 ;
        RECT 109.540 189.480 109.860 189.540 ;
        RECT 110.015 189.480 110.305 189.525 ;
        RECT 109.540 189.340 110.305 189.480 ;
        RECT 109.540 189.280 109.860 189.340 ;
        RECT 110.015 189.295 110.305 189.340 ;
        RECT 111.840 189.140 112.160 189.200 ;
        RECT 107.485 189.125 112.160 189.140 ;
        RECT 107.710 189.000 112.160 189.125 ;
        RECT 111.840 188.940 112.160 189.000 ;
        RECT 124.735 189.140 125.025 189.185 ;
        RECT 125.180 189.140 125.500 189.200 ;
        RECT 124.735 189.000 125.500 189.140 ;
        RECT 124.735 188.955 125.025 189.000 ;
        RECT 125.180 188.940 125.500 189.000 ;
        RECT 126.070 189.140 126.360 189.185 ;
        RECT 129.780 189.140 130.100 189.200 ;
        RECT 126.070 189.000 130.100 189.140 ;
        RECT 131.710 189.140 131.850 189.635 ;
        RECT 133.920 189.140 134.240 189.200 ;
        RECT 134.855 189.140 135.145 189.185 ;
        RECT 131.710 189.000 135.145 189.140 ;
        RECT 126.070 188.955 126.360 189.000 ;
        RECT 129.780 188.940 130.100 189.000 ;
        RECT 133.920 188.940 134.240 189.000 ;
        RECT 134.855 188.955 135.145 189.000 ;
        RECT 135.760 188.940 136.080 189.200 ;
        RECT 95.740 188.660 100.570 188.800 ;
        RECT 95.740 188.600 96.060 188.660 ;
        RECT 94.835 188.275 95.125 188.505 ;
        RECT 95.295 188.275 95.585 188.505 ;
        RECT 96.200 188.460 96.520 188.520 ;
        RECT 101.735 188.460 102.025 188.505 ;
        RECT 104.570 188.460 104.710 188.940 ;
        RECT 104.940 188.800 105.260 188.860 ;
        RECT 115.980 188.800 116.300 188.860 ;
        RECT 104.940 188.660 116.300 188.800 ;
        RECT 104.940 188.600 105.260 188.660 ;
        RECT 115.980 188.600 116.300 188.660 ;
        RECT 125.615 188.800 125.905 188.845 ;
        RECT 126.805 188.800 127.095 188.845 ;
        RECT 129.325 188.800 129.615 188.845 ;
        RECT 125.615 188.660 129.615 188.800 ;
        RECT 125.615 188.615 125.905 188.660 ;
        RECT 126.805 188.615 127.095 188.660 ;
        RECT 129.325 188.615 129.615 188.660 ;
        RECT 131.620 188.800 131.940 188.860 ;
        RECT 132.095 188.800 132.385 188.845 ;
        RECT 131.620 188.660 132.385 188.800 ;
        RECT 131.620 188.600 131.940 188.660 ;
        RECT 132.095 188.615 132.385 188.660 ;
        RECT 109.540 188.460 109.860 188.520 ;
        RECT 112.315 188.460 112.605 188.505 ;
        RECT 113.220 188.460 113.540 188.520 ;
        RECT 96.200 188.320 102.025 188.460 ;
        RECT 95.370 188.120 95.510 188.275 ;
        RECT 96.200 188.260 96.520 188.320 ;
        RECT 101.735 188.275 102.025 188.320 ;
        RECT 103.190 188.320 107.930 188.460 ;
        RECT 91.690 187.980 95.510 188.120 ;
        RECT 76.880 187.920 77.200 187.980 ;
        RECT 85.160 187.920 85.480 187.980 ;
        RECT 97.120 187.920 97.440 188.180 ;
        RECT 98.055 188.120 98.345 188.165 ;
        RECT 103.190 188.120 103.330 188.320 ;
        RECT 107.790 188.180 107.930 188.320 ;
        RECT 109.540 188.320 113.540 188.460 ;
        RECT 109.540 188.260 109.860 188.320 ;
        RECT 112.315 188.275 112.605 188.320 ;
        RECT 113.220 188.260 113.540 188.320 ;
        RECT 125.220 188.460 125.510 188.505 ;
        RECT 127.320 188.460 127.610 188.505 ;
        RECT 128.890 188.460 129.180 188.505 ;
        RECT 125.220 188.320 129.180 188.460 ;
        RECT 125.220 188.275 125.510 188.320 ;
        RECT 127.320 188.275 127.610 188.320 ;
        RECT 128.890 188.275 129.180 188.320 ;
        RECT 98.055 187.980 103.330 188.120 ;
        RECT 98.055 187.935 98.345 187.980 ;
        RECT 103.560 187.920 103.880 188.180 ;
        RECT 105.400 188.120 105.720 188.180 ;
        RECT 106.780 188.120 107.100 188.180 ;
        RECT 105.400 187.980 107.100 188.120 ;
        RECT 105.400 187.920 105.720 187.980 ;
        RECT 106.780 187.920 107.100 187.980 ;
        RECT 107.700 187.920 108.020 188.180 ;
        RECT 110.935 188.120 111.225 188.165 ;
        RECT 111.380 188.120 111.700 188.180 ;
        RECT 110.935 187.980 111.700 188.120 ;
        RECT 110.935 187.935 111.225 187.980 ;
        RECT 111.380 187.920 111.700 187.980 ;
        RECT 111.855 188.120 112.145 188.165 ;
        RECT 112.760 188.120 113.080 188.180 ;
        RECT 111.855 187.980 113.080 188.120 ;
        RECT 111.855 187.935 112.145 187.980 ;
        RECT 112.760 187.920 113.080 187.980 ;
        RECT 113.680 188.120 114.000 188.180 ;
        RECT 114.155 188.120 114.445 188.165 ;
        RECT 114.600 188.120 114.920 188.180 ;
        RECT 113.680 187.980 114.920 188.120 ;
        RECT 113.680 187.920 114.000 187.980 ;
        RECT 114.155 187.935 114.445 187.980 ;
        RECT 114.600 187.920 114.920 187.980 ;
        RECT 115.060 187.920 115.380 188.180 ;
        RECT 136.680 187.920 137.000 188.180 ;
        RECT 13.330 187.300 138.910 187.780 ;
        RECT 25.820 187.100 26.140 187.160 ;
        RECT 30.420 187.100 30.740 187.160 ;
        RECT 25.820 186.960 30.740 187.100 ;
        RECT 25.820 186.900 26.140 186.960 ;
        RECT 30.420 186.900 30.740 186.960 ;
        RECT 31.340 187.100 31.660 187.160 ;
        RECT 31.815 187.100 32.105 187.145 ;
        RECT 31.340 186.960 32.105 187.100 ;
        RECT 31.340 186.900 31.660 186.960 ;
        RECT 31.815 186.915 32.105 186.960 ;
        RECT 35.020 187.100 35.340 187.160 ;
        RECT 95.755 187.100 96.045 187.145 ;
        RECT 97.120 187.100 97.440 187.160 ;
        RECT 35.020 186.960 45.830 187.100 ;
        RECT 35.020 186.900 35.340 186.960 ;
        RECT 21.680 186.760 22.000 186.820 ;
        RECT 26.280 186.760 26.600 186.820 ;
        RECT 21.680 186.620 26.600 186.760 ;
        RECT 21.680 186.560 22.000 186.620 ;
        RECT 26.280 186.560 26.600 186.620 ;
        RECT 26.740 186.760 27.060 186.820 ;
        RECT 33.640 186.760 33.960 186.820 ;
        RECT 26.740 186.620 33.960 186.760 ;
        RECT 26.740 186.560 27.060 186.620 ;
        RECT 33.640 186.560 33.960 186.620 ;
        RECT 34.115 186.760 34.405 186.805 ;
        RECT 39.620 186.760 39.940 186.820 ;
        RECT 34.115 186.620 39.940 186.760 ;
        RECT 34.115 186.575 34.405 186.620 ;
        RECT 39.620 186.560 39.940 186.620 ;
        RECT 45.690 186.760 45.830 186.960 ;
        RECT 95.755 186.960 97.440 187.100 ;
        RECT 95.755 186.915 96.045 186.960 ;
        RECT 97.120 186.900 97.440 186.960 ;
        RECT 97.595 187.100 97.885 187.145 ;
        RECT 102.640 187.100 102.960 187.160 ;
        RECT 97.595 186.960 102.960 187.100 ;
        RECT 97.595 186.915 97.885 186.960 ;
        RECT 102.640 186.900 102.960 186.960 ;
        RECT 104.480 187.100 104.800 187.160 ;
        RECT 105.860 187.100 106.180 187.160 ;
        RECT 104.480 186.960 106.180 187.100 ;
        RECT 104.480 186.900 104.800 186.960 ;
        RECT 105.860 186.900 106.180 186.960 ;
        RECT 108.175 187.100 108.465 187.145 ;
        RECT 108.620 187.100 108.940 187.160 ;
        RECT 114.600 187.100 114.920 187.160 ;
        RECT 108.175 186.960 111.150 187.100 ;
        RECT 108.175 186.915 108.465 186.960 ;
        RECT 108.620 186.900 108.940 186.960 ;
        RECT 51.120 186.760 51.440 186.820 ;
        RECT 69.060 186.760 69.380 186.820 ;
        RECT 90.235 186.760 90.525 186.805 ;
        RECT 93.915 186.760 94.205 186.805 ;
        RECT 45.690 186.620 51.440 186.760 ;
        RECT 20.300 186.220 20.620 186.480 ;
        RECT 21.770 186.420 21.910 186.560 ;
        RECT 20.850 186.280 21.910 186.420 ;
        RECT 31.430 186.280 36.630 186.420 ;
        RECT 19.840 186.080 20.160 186.140 ;
        RECT 20.850 186.080 20.990 186.280 ;
        RECT 19.840 185.940 20.990 186.080 ;
        RECT 21.220 186.080 21.540 186.140 ;
        RECT 21.695 186.080 21.985 186.125 ;
        RECT 23.520 186.080 23.840 186.140 ;
        RECT 21.220 185.940 23.840 186.080 ;
        RECT 19.840 185.880 20.160 185.940 ;
        RECT 21.220 185.880 21.540 185.940 ;
        RECT 21.695 185.895 21.985 185.940 ;
        RECT 23.520 185.880 23.840 185.940 ;
        RECT 30.880 186.080 31.200 186.140 ;
        RECT 31.430 186.080 31.570 186.280 ;
        RECT 30.880 185.940 31.570 186.080 ;
        RECT 30.880 185.880 31.200 185.940 ;
        RECT 31.815 185.895 32.105 186.125 ;
        RECT 19.270 185.740 19.560 185.785 ;
        RECT 25.820 185.740 26.140 185.800 ;
        RECT 19.270 185.600 26.140 185.740 ;
        RECT 19.270 185.555 19.560 185.600 ;
        RECT 25.820 185.540 26.140 185.600 ;
        RECT 18.460 185.200 18.780 185.460 ;
        RECT 31.890 185.400 32.030 185.895 ;
        RECT 32.260 185.880 32.580 186.140 ;
        RECT 33.180 185.880 33.500 186.140 ;
        RECT 33.640 186.080 33.960 186.140 ;
        RECT 35.955 186.080 36.245 186.125 ;
        RECT 33.640 185.940 36.245 186.080 ;
        RECT 33.640 185.880 33.960 185.940 ;
        RECT 35.955 185.895 36.245 185.940 ;
        RECT 33.270 185.740 33.410 185.880 ;
        RECT 35.495 185.740 35.785 185.785 ;
        RECT 33.270 185.600 35.785 185.740 ;
        RECT 36.490 185.740 36.630 186.280 ;
        RECT 37.780 186.220 38.100 186.480 ;
        RECT 45.690 186.465 45.830 186.620 ;
        RECT 51.120 186.560 51.440 186.620 ;
        RECT 60.410 186.620 69.380 186.760 ;
        RECT 39.175 186.420 39.465 186.465 ;
        RECT 45.615 186.420 45.905 186.465 ;
        RECT 38.330 186.280 39.465 186.420 ;
        RECT 45.505 186.280 45.905 186.420 ;
        RECT 37.320 185.880 37.640 186.140 ;
        RECT 38.330 186.125 38.470 186.280 ;
        RECT 39.175 186.235 39.465 186.280 ;
        RECT 45.615 186.235 45.905 186.280 ;
        RECT 59.875 186.420 60.165 186.465 ;
        RECT 60.410 186.420 60.550 186.620 ;
        RECT 69.060 186.560 69.380 186.620 ;
        RECT 88.470 186.620 94.205 186.760 ;
        RECT 88.470 186.480 88.610 186.620 ;
        RECT 90.235 186.575 90.525 186.620 ;
        RECT 93.915 186.575 94.205 186.620 ;
        RECT 94.360 186.760 94.680 186.820 ;
        RECT 99.895 186.760 100.185 186.805 ;
        RECT 104.940 186.760 105.260 186.820 ;
        RECT 111.010 186.805 111.150 186.960 ;
        RECT 112.390 186.960 114.920 187.100 ;
        RECT 94.360 186.620 105.260 186.760 ;
        RECT 94.360 186.560 94.680 186.620 ;
        RECT 99.895 186.575 100.185 186.620 ;
        RECT 104.940 186.560 105.260 186.620 ;
        RECT 110.935 186.575 111.225 186.805 ;
        RECT 111.380 186.760 111.700 186.820 ;
        RECT 112.390 186.760 112.530 186.960 ;
        RECT 114.600 186.900 114.920 186.960 ;
        RECT 115.520 187.100 115.840 187.160 ;
        RECT 117.360 187.100 117.680 187.160 ;
        RECT 115.520 186.960 117.680 187.100 ;
        RECT 115.520 186.900 115.840 186.960 ;
        RECT 117.360 186.900 117.680 186.960 ;
        RECT 120.135 186.915 120.425 187.145 ;
        RECT 111.380 186.620 112.530 186.760 ;
        RECT 113.235 186.760 113.525 186.805 ;
        RECT 113.680 186.760 114.000 186.820 ;
        RECT 113.235 186.620 114.000 186.760 ;
        RECT 114.690 186.760 114.830 186.900 ;
        RECT 117.835 186.760 118.125 186.805 ;
        RECT 114.690 186.620 118.125 186.760 ;
        RECT 59.875 186.280 60.550 186.420 ;
        RECT 60.795 186.420 61.085 186.465 ;
        RECT 62.175 186.420 62.465 186.465 ;
        RECT 60.795 186.280 62.465 186.420 ;
        RECT 59.875 186.235 60.165 186.280 ;
        RECT 60.795 186.235 61.085 186.280 ;
        RECT 62.175 186.235 62.465 186.280 ;
        RECT 63.540 186.420 63.860 186.480 ;
        RECT 63.540 186.280 66.990 186.420 ;
        RECT 63.540 186.220 63.860 186.280 ;
        RECT 38.255 185.895 38.545 186.125 ;
        RECT 38.715 185.895 39.005 186.125 ;
        RECT 38.790 185.740 38.930 185.895 ;
        RECT 39.620 185.880 39.940 186.140 ;
        RECT 43.300 186.080 43.620 186.140 ;
        RECT 49.295 186.080 49.585 186.125 ;
        RECT 43.300 185.940 49.585 186.080 ;
        RECT 43.300 185.880 43.620 185.940 ;
        RECT 49.295 185.895 49.585 185.940 ;
        RECT 50.215 186.080 50.505 186.125 ;
        RECT 53.420 186.080 53.740 186.140 ;
        RECT 50.215 185.940 53.740 186.080 ;
        RECT 50.215 185.895 50.505 185.940 ;
        RECT 53.420 185.880 53.740 185.940 ;
        RECT 60.335 185.895 60.625 186.125 ;
        RECT 61.255 185.895 61.545 186.125 ;
        RECT 64.000 186.080 64.320 186.140 ;
        RECT 64.920 186.080 65.240 186.140 ;
        RECT 64.000 185.940 65.240 186.080 ;
        RECT 36.490 185.600 38.930 185.740 ;
        RECT 48.040 185.740 48.330 185.785 ;
        RECT 49.755 185.740 50.045 185.785 ;
        RECT 48.040 185.600 50.045 185.740 ;
        RECT 35.495 185.555 35.785 185.600 ;
        RECT 48.040 185.555 48.330 185.600 ;
        RECT 49.755 185.555 50.045 185.600 ;
        RECT 32.765 185.400 33.055 185.445 ;
        RECT 31.890 185.260 33.055 185.400 ;
        RECT 32.765 185.215 33.055 185.260 ;
        RECT 34.560 185.400 34.880 185.460 ;
        RECT 35.035 185.400 35.325 185.445 ;
        RECT 34.560 185.260 35.325 185.400 ;
        RECT 34.560 185.200 34.880 185.260 ;
        RECT 35.035 185.215 35.325 185.260 ;
        RECT 36.875 185.400 37.165 185.445 ;
        RECT 37.320 185.400 37.640 185.460 ;
        RECT 41.920 185.400 42.240 185.460 ;
        RECT 36.875 185.260 42.240 185.400 ;
        RECT 36.875 185.215 37.165 185.260 ;
        RECT 37.320 185.200 37.640 185.260 ;
        RECT 41.920 185.200 42.240 185.260 ;
        RECT 46.980 185.200 47.300 185.460 ;
        RECT 47.440 185.200 47.760 185.460 ;
        RECT 48.820 185.200 49.140 185.460 ;
        RECT 58.480 185.400 58.800 185.460 ;
        RECT 58.955 185.400 59.245 185.445 ;
        RECT 58.480 185.260 59.245 185.400 ;
        RECT 60.410 185.400 60.550 185.895 ;
        RECT 61.330 185.740 61.470 185.895 ;
        RECT 64.000 185.880 64.320 185.940 ;
        RECT 64.920 185.880 65.240 185.940 ;
        RECT 66.300 185.740 66.620 185.800 ;
        RECT 61.330 185.600 66.620 185.740 ;
        RECT 66.850 185.740 66.990 186.280 ;
        RECT 68.690 186.280 70.670 186.420 ;
        RECT 67.220 186.080 67.540 186.140 ;
        RECT 68.690 186.125 68.830 186.280 ;
        RECT 70.530 186.140 70.670 186.280 ;
        RECT 88.380 186.220 88.700 186.480 ;
        RECT 91.140 186.420 91.460 186.480 ;
        RECT 92.535 186.420 92.825 186.465 ;
        RECT 98.040 186.420 98.360 186.480 ;
        RECT 109.540 186.420 109.860 186.480 ;
        RECT 91.140 186.280 92.825 186.420 ;
        RECT 91.140 186.220 91.460 186.280 ;
        RECT 92.535 186.235 92.825 186.280 ;
        RECT 96.290 186.280 98.360 186.420 ;
        RECT 68.615 186.080 68.905 186.125 ;
        RECT 67.220 185.940 68.905 186.080 ;
        RECT 67.220 185.880 67.540 185.940 ;
        RECT 68.615 185.895 68.905 185.940 ;
        RECT 69.520 185.880 69.840 186.140 ;
        RECT 70.440 185.880 70.760 186.140 ;
        RECT 70.915 185.895 71.205 186.125 ;
        RECT 69.995 185.740 70.285 185.785 ;
        RECT 70.990 185.740 71.130 185.895 ;
        RECT 71.820 185.880 72.140 186.140 ;
        RECT 75.500 186.080 75.820 186.140 ;
        RECT 78.275 186.080 78.565 186.125 ;
        RECT 75.500 185.940 78.565 186.080 ;
        RECT 75.500 185.880 75.820 185.940 ;
        RECT 78.275 185.895 78.565 185.940 ;
        RECT 85.620 186.080 85.940 186.140 ;
        RECT 87.935 186.080 88.225 186.125 ;
        RECT 85.620 185.940 88.225 186.080 ;
        RECT 88.470 186.080 88.610 186.220 ;
        RECT 88.855 186.080 89.145 186.125 ;
        RECT 88.470 185.940 89.145 186.080 ;
        RECT 85.620 185.880 85.940 185.940 ;
        RECT 87.935 185.895 88.225 185.940 ;
        RECT 88.855 185.895 89.145 185.940 ;
        RECT 89.315 185.895 89.605 186.125 ;
        RECT 90.235 186.080 90.525 186.125 ;
        RECT 92.980 186.080 93.300 186.140 ;
        RECT 93.900 186.080 94.220 186.140 ;
        RECT 95.740 186.080 96.060 186.140 ;
        RECT 96.290 186.125 96.430 186.280 ;
        RECT 98.040 186.220 98.360 186.280 ;
        RECT 108.170 186.280 109.860 186.420 ;
        RECT 111.010 186.420 111.150 186.575 ;
        RECT 111.380 186.560 111.700 186.620 ;
        RECT 113.235 186.575 113.525 186.620 ;
        RECT 113.680 186.560 114.000 186.620 ;
        RECT 117.835 186.575 118.125 186.620 ;
        RECT 114.140 186.420 114.460 186.480 ;
        RECT 114.615 186.420 114.905 186.465 ;
        RECT 111.010 186.280 114.905 186.420 ;
        RECT 90.235 185.940 93.670 186.080 ;
        RECT 90.235 185.895 90.525 185.940 ;
        RECT 66.850 185.600 71.130 185.740 ;
        RECT 89.390 185.740 89.530 185.895 ;
        RECT 92.980 185.880 93.300 185.940 ;
        RECT 91.600 185.740 91.920 185.800 ;
        RECT 89.390 185.600 91.920 185.740 ;
        RECT 93.530 185.740 93.670 185.940 ;
        RECT 93.900 185.940 96.060 186.080 ;
        RECT 93.900 185.880 94.220 185.940 ;
        RECT 95.740 185.880 96.060 185.940 ;
        RECT 96.215 185.895 96.505 186.125 ;
        RECT 97.135 185.895 97.425 186.125 ;
        RECT 101.270 185.895 101.560 186.125 ;
        RECT 101.735 186.080 102.025 186.125 ;
        RECT 103.100 186.080 103.420 186.140 ;
        RECT 101.735 185.940 103.420 186.080 ;
        RECT 108.170 185.955 108.310 186.280 ;
        RECT 109.540 186.220 109.860 186.280 ;
        RECT 114.140 186.220 114.460 186.280 ;
        RECT 114.615 186.235 114.905 186.280 ;
        RECT 115.535 186.420 115.825 186.465 ;
        RECT 118.280 186.420 118.600 186.480 ;
        RECT 115.535 186.280 118.600 186.420 ;
        RECT 115.535 186.235 115.825 186.280 ;
        RECT 118.280 186.220 118.600 186.280 ;
        RECT 118.755 186.420 119.045 186.465 ;
        RECT 120.210 186.420 120.350 186.915 ;
        RECT 129.780 186.900 130.100 187.160 ;
        RECT 121.500 186.420 121.820 186.480 ;
        RECT 118.755 186.280 121.820 186.420 ;
        RECT 118.755 186.235 119.045 186.280 ;
        RECT 121.500 186.220 121.820 186.280 ;
        RECT 125.180 186.420 125.500 186.480 ;
        RECT 132.555 186.420 132.845 186.465 ;
        RECT 125.180 186.280 132.845 186.420 ;
        RECT 125.180 186.220 125.500 186.280 ;
        RECT 132.555 186.235 132.845 186.280 ;
        RECT 110.920 186.080 111.240 186.140 ;
        RECT 101.735 185.895 102.025 185.940 ;
        RECT 97.210 185.740 97.350 185.895 ;
        RECT 93.530 185.600 97.350 185.740 ;
        RECT 101.350 185.740 101.490 185.895 ;
        RECT 103.100 185.880 103.420 185.940 ;
        RECT 106.320 185.740 106.640 185.800 ;
        RECT 101.350 185.600 106.640 185.740 ;
        RECT 107.945 185.770 108.310 185.955 ;
        RECT 109.170 185.940 111.240 186.080 ;
        RECT 109.170 185.785 109.310 185.940 ;
        RECT 110.920 185.880 111.240 185.940 ;
        RECT 111.840 186.080 112.160 186.140 ;
        RECT 111.840 185.940 114.830 186.080 ;
        RECT 111.840 185.880 112.160 185.940 ;
        RECT 107.945 185.725 108.235 185.770 ;
        RECT 66.300 185.540 66.620 185.600 ;
        RECT 69.995 185.555 70.285 185.600 ;
        RECT 91.600 185.540 91.920 185.600 ;
        RECT 106.320 185.540 106.640 185.600 ;
        RECT 109.095 185.555 109.385 185.785 ;
        RECT 63.540 185.400 63.860 185.460 ;
        RECT 60.410 185.260 63.860 185.400 ;
        RECT 58.480 185.200 58.800 185.260 ;
        RECT 58.955 185.215 59.245 185.260 ;
        RECT 63.540 185.200 63.860 185.260 ;
        RECT 65.855 185.400 66.145 185.445 ;
        RECT 67.220 185.400 67.540 185.460 ;
        RECT 65.855 185.260 67.540 185.400 ;
        RECT 65.855 185.215 66.145 185.260 ;
        RECT 67.220 185.200 67.540 185.260 ;
        RECT 71.375 185.400 71.665 185.445 ;
        RECT 73.660 185.400 73.980 185.460 ;
        RECT 71.375 185.260 73.980 185.400 ;
        RECT 71.375 185.215 71.665 185.260 ;
        RECT 73.660 185.200 73.980 185.260 ;
        RECT 80.100 185.400 80.420 185.460 ;
        RECT 81.020 185.400 81.340 185.460 ;
        RECT 81.495 185.400 81.785 185.445 ;
        RECT 80.100 185.260 81.785 185.400 ;
        RECT 80.100 185.200 80.420 185.260 ;
        RECT 81.020 185.200 81.340 185.260 ;
        RECT 81.495 185.215 81.785 185.260 ;
        RECT 88.395 185.400 88.685 185.445 ;
        RECT 93.900 185.400 94.220 185.460 ;
        RECT 88.395 185.260 94.220 185.400 ;
        RECT 88.395 185.215 88.685 185.260 ;
        RECT 93.900 185.200 94.220 185.260 ;
        RECT 94.835 185.400 95.125 185.445 ;
        RECT 106.780 185.400 107.100 185.460 ;
        RECT 94.835 185.260 107.100 185.400 ;
        RECT 94.835 185.215 95.125 185.260 ;
        RECT 106.780 185.200 107.100 185.260 ;
        RECT 107.240 185.200 107.560 185.460 ;
        RECT 111.840 185.200 112.160 185.460 ;
        RECT 112.390 185.445 112.530 185.940 ;
        RECT 114.690 185.800 114.830 185.940 ;
        RECT 115.075 186.050 115.365 186.125 ;
        RECT 115.075 186.030 115.750 186.050 ;
        RECT 115.075 185.910 115.840 186.030 ;
        RECT 115.075 185.895 115.365 185.910 ;
        RECT 114.600 185.540 114.920 185.800 ;
        RECT 115.520 185.770 115.840 185.910 ;
        RECT 117.375 185.895 117.665 186.125 ;
        RECT 118.370 186.080 118.510 186.220 ;
        RECT 119.215 186.080 119.505 186.125 ;
        RECT 118.370 185.940 119.505 186.080 ;
        RECT 119.215 185.895 119.505 185.940 ;
        RECT 117.450 185.740 117.590 185.895 ;
        RECT 131.620 185.880 131.940 186.140 ;
        RECT 133.935 185.895 134.225 186.125 ;
        RECT 116.070 185.600 117.590 185.740 ;
        RECT 126.100 185.740 126.420 185.800 ;
        RECT 134.010 185.740 134.150 185.895 ;
        RECT 135.760 185.880 136.080 186.140 ;
        RECT 126.100 185.600 134.150 185.740 ;
        RECT 112.315 185.215 112.605 185.445 ;
        RECT 113.680 185.400 114.000 185.460 ;
        RECT 116.070 185.400 116.210 185.600 ;
        RECT 126.100 185.540 126.420 185.600 ;
        RECT 113.680 185.260 116.210 185.400 ;
        RECT 116.915 185.400 117.205 185.445 ;
        RECT 117.820 185.400 118.140 185.460 ;
        RECT 116.915 185.260 118.140 185.400 ;
        RECT 113.680 185.200 114.000 185.260 ;
        RECT 116.915 185.215 117.205 185.260 ;
        RECT 117.820 185.200 118.140 185.260 ;
        RECT 118.755 185.400 119.045 185.445 ;
        RECT 119.660 185.400 119.980 185.460 ;
        RECT 118.755 185.260 119.980 185.400 ;
        RECT 118.755 185.215 119.045 185.260 ;
        RECT 119.660 185.200 119.980 185.260 ;
        RECT 127.480 185.400 127.800 185.460 ;
        RECT 132.095 185.400 132.385 185.445 ;
        RECT 127.480 185.260 132.385 185.400 ;
        RECT 127.480 185.200 127.800 185.260 ;
        RECT 132.095 185.215 132.385 185.260 ;
        RECT 134.840 185.200 135.160 185.460 ;
        RECT 136.695 185.400 136.985 185.445 ;
        RECT 137.600 185.400 137.920 185.460 ;
        RECT 136.695 185.260 137.920 185.400 ;
        RECT 136.695 185.215 136.985 185.260 ;
        RECT 137.600 185.200 137.920 185.260 ;
        RECT 13.330 184.580 138.910 185.060 ;
        RECT 25.820 184.180 26.140 184.440 ;
        RECT 42.380 184.380 42.700 184.440 ;
        RECT 44.775 184.380 45.065 184.425 ;
        RECT 42.010 184.240 45.065 184.380 ;
        RECT 18.460 184.040 18.780 184.100 ;
        RECT 19.240 184.040 19.530 184.085 ;
        RECT 18.460 183.900 19.530 184.040 ;
        RECT 18.460 183.840 18.780 183.900 ;
        RECT 19.240 183.855 19.530 183.900 ;
        RECT 12.020 183.700 12.340 183.760 ;
        RECT 14.795 183.700 15.085 183.745 ;
        RECT 12.020 183.560 15.085 183.700 ;
        RECT 12.020 183.500 12.340 183.560 ;
        RECT 14.795 183.515 15.085 183.560 ;
        RECT 24.440 183.700 24.760 183.760 ;
        RECT 25.375 183.700 25.665 183.745 ;
        RECT 24.440 183.560 25.665 183.700 ;
        RECT 24.440 183.500 24.760 183.560 ;
        RECT 25.375 183.515 25.665 183.560 ;
        RECT 26.295 183.700 26.585 183.745 ;
        RECT 26.740 183.700 27.060 183.760 ;
        RECT 42.010 183.745 42.150 184.240 ;
        RECT 42.380 184.180 42.700 184.240 ;
        RECT 44.775 184.195 45.065 184.240 ;
        RECT 45.615 184.380 45.905 184.425 ;
        RECT 53.420 184.380 53.740 184.440 ;
        RECT 45.615 184.240 53.740 184.380 ;
        RECT 45.615 184.195 45.905 184.240 ;
        RECT 53.420 184.180 53.740 184.240 ;
        RECT 64.475 184.380 64.765 184.425 ;
        RECT 66.760 184.380 67.080 184.440 ;
        RECT 64.475 184.240 67.080 184.380 ;
        RECT 64.475 184.195 64.765 184.240 ;
        RECT 66.760 184.180 67.080 184.240 ;
        RECT 67.220 184.180 67.540 184.440 ;
        RECT 69.060 184.380 69.380 184.440 ;
        RECT 71.820 184.380 72.140 184.440 ;
        RECT 69.060 184.240 72.140 184.380 ;
        RECT 69.060 184.180 69.380 184.240 ;
        RECT 71.820 184.180 72.140 184.240 ;
        RECT 75.500 184.180 75.820 184.440 ;
        RECT 118.740 184.380 119.060 184.440 ;
        RECT 110.090 184.240 119.060 184.380 ;
        RECT 43.775 183.855 44.065 184.085 ;
        RECT 49.280 184.040 49.600 184.100 ;
        RECT 46.150 183.900 49.600 184.040 ;
        RECT 26.295 183.560 27.060 183.700 ;
        RECT 26.295 183.515 26.585 183.560 ;
        RECT 26.740 183.500 27.060 183.560 ;
        RECT 41.935 183.515 42.225 183.745 ;
        RECT 42.395 183.515 42.685 183.745 ;
        RECT 42.840 183.700 43.160 183.760 ;
        RECT 43.315 183.700 43.605 183.745 ;
        RECT 43.850 183.700 43.990 183.855 ;
        RECT 46.150 183.745 46.290 183.900 ;
        RECT 49.280 183.840 49.600 183.900 ;
        RECT 71.360 184.040 71.680 184.100 ;
        RECT 75.040 184.040 75.360 184.100 ;
        RECT 71.360 183.900 75.360 184.040 ;
        RECT 71.360 183.840 71.680 183.900 ;
        RECT 75.040 183.840 75.360 183.900 ;
        RECT 42.840 183.560 43.990 183.700 ;
        RECT 17.540 183.360 17.860 183.420 ;
        RECT 18.015 183.360 18.305 183.405 ;
        RECT 17.540 183.220 18.305 183.360 ;
        RECT 17.540 183.160 17.860 183.220 ;
        RECT 18.015 183.175 18.305 183.220 ;
        RECT 18.895 183.360 19.185 183.405 ;
        RECT 20.085 183.360 20.375 183.405 ;
        RECT 22.605 183.360 22.895 183.405 ;
        RECT 18.895 183.220 22.895 183.360 ;
        RECT 18.895 183.175 19.185 183.220 ;
        RECT 20.085 183.175 20.375 183.220 ;
        RECT 22.605 183.175 22.895 183.220 ;
        RECT 41.460 183.360 41.780 183.420 ;
        RECT 42.010 183.360 42.150 183.515 ;
        RECT 41.460 183.220 42.150 183.360 ;
        RECT 41.460 183.160 41.780 183.220 ;
        RECT 18.500 183.020 18.790 183.065 ;
        RECT 20.600 183.020 20.890 183.065 ;
        RECT 22.170 183.020 22.460 183.065 ;
        RECT 18.500 182.880 22.460 183.020 ;
        RECT 18.500 182.835 18.790 182.880 ;
        RECT 20.600 182.835 20.890 182.880 ;
        RECT 22.170 182.835 22.460 182.880 ;
        RECT 15.715 182.680 16.005 182.725 ;
        RECT 23.980 182.680 24.300 182.740 ;
        RECT 15.715 182.540 24.300 182.680 ;
        RECT 15.715 182.495 16.005 182.540 ;
        RECT 23.980 182.480 24.300 182.540 ;
        RECT 24.900 182.480 25.220 182.740 ;
        RECT 40.080 182.680 40.400 182.740 ;
        RECT 41.000 182.680 41.320 182.740 ;
        RECT 42.470 182.680 42.610 183.515 ;
        RECT 42.840 183.500 43.160 183.560 ;
        RECT 43.315 183.515 43.605 183.560 ;
        RECT 43.300 182.820 43.620 183.080 ;
        RECT 43.850 183.020 43.990 183.560 ;
        RECT 46.075 183.515 46.365 183.745 ;
        RECT 47.410 183.700 47.700 183.745 ;
        RECT 48.820 183.700 49.140 183.760 ;
        RECT 47.410 183.560 49.140 183.700 ;
        RECT 47.410 183.515 47.700 183.560 ;
        RECT 48.820 183.500 49.140 183.560 ;
        RECT 58.910 183.700 59.200 183.745 ;
        RECT 65.395 183.700 65.685 183.745 ;
        RECT 58.910 183.560 65.685 183.700 ;
        RECT 58.910 183.515 59.200 183.560 ;
        RECT 65.395 183.515 65.685 183.560 ;
        RECT 66.300 183.500 66.620 183.760 ;
        RECT 67.680 183.500 68.000 183.760 ;
        RECT 68.140 183.500 68.460 183.760 ;
        RECT 69.490 183.700 69.780 183.745 ;
        RECT 72.280 183.700 72.600 183.760 ;
        RECT 69.490 183.560 72.600 183.700 ;
        RECT 69.490 183.515 69.780 183.560 ;
        RECT 72.280 183.500 72.600 183.560 ;
        RECT 46.955 183.360 47.245 183.405 ;
        RECT 48.145 183.360 48.435 183.405 ;
        RECT 50.665 183.360 50.955 183.405 ;
        RECT 46.955 183.220 50.955 183.360 ;
        RECT 46.955 183.175 47.245 183.220 ;
        RECT 48.145 183.175 48.435 183.220 ;
        RECT 50.665 183.175 50.955 183.220 ;
        RECT 55.720 183.360 56.040 183.420 ;
        RECT 57.575 183.360 57.865 183.405 ;
        RECT 55.720 183.220 57.865 183.360 ;
        RECT 55.720 183.160 56.040 183.220 ;
        RECT 57.575 183.175 57.865 183.220 ;
        RECT 58.455 183.360 58.745 183.405 ;
        RECT 59.645 183.360 59.935 183.405 ;
        RECT 62.165 183.360 62.455 183.405 ;
        RECT 58.455 183.220 62.455 183.360 ;
        RECT 58.455 183.175 58.745 183.220 ;
        RECT 59.645 183.175 59.935 183.220 ;
        RECT 62.165 183.175 62.455 183.220 ;
        RECT 69.035 183.360 69.325 183.405 ;
        RECT 70.225 183.360 70.515 183.405 ;
        RECT 72.745 183.360 73.035 183.405 ;
        RECT 69.035 183.220 73.035 183.360 ;
        RECT 69.035 183.175 69.325 183.220 ;
        RECT 70.225 183.175 70.515 183.220 ;
        RECT 72.745 183.175 73.035 183.220 ;
        RECT 46.560 183.020 46.850 183.065 ;
        RECT 48.660 183.020 48.950 183.065 ;
        RECT 50.230 183.020 50.520 183.065 ;
        RECT 43.850 182.880 46.290 183.020 ;
        RECT 44.695 182.680 44.985 182.725 ;
        RECT 40.080 182.540 44.985 182.680 ;
        RECT 46.150 182.680 46.290 182.880 ;
        RECT 46.560 182.880 50.520 183.020 ;
        RECT 46.560 182.835 46.850 182.880 ;
        RECT 48.660 182.835 48.950 182.880 ;
        RECT 50.230 182.835 50.520 182.880 ;
        RECT 58.060 183.020 58.350 183.065 ;
        RECT 60.160 183.020 60.450 183.065 ;
        RECT 61.730 183.020 62.020 183.065 ;
        RECT 58.060 182.880 62.020 183.020 ;
        RECT 58.060 182.835 58.350 182.880 ;
        RECT 60.160 182.835 60.450 182.880 ;
        RECT 61.730 182.835 62.020 182.880 ;
        RECT 68.640 183.020 68.930 183.065 ;
        RECT 70.740 183.020 71.030 183.065 ;
        RECT 72.310 183.020 72.600 183.065 ;
        RECT 75.590 183.020 75.730 184.180 ;
        RECT 109.555 184.040 109.845 184.085 ;
        RECT 68.640 182.880 72.600 183.020 ;
        RECT 68.640 182.835 68.930 182.880 ;
        RECT 70.740 182.835 71.030 182.880 ;
        RECT 72.310 182.835 72.600 182.880 ;
        RECT 74.670 182.880 75.730 183.020 ;
        RECT 76.050 183.900 86.770 184.040 ;
        RECT 52.975 182.680 53.265 182.725 ;
        RECT 55.260 182.680 55.580 182.740 ;
        RECT 46.150 182.540 55.580 182.680 ;
        RECT 40.080 182.480 40.400 182.540 ;
        RECT 41.000 182.480 41.320 182.540 ;
        RECT 44.695 182.495 44.985 182.540 ;
        RECT 52.975 182.495 53.265 182.540 ;
        RECT 55.260 182.480 55.580 182.540 ;
        RECT 69.060 182.680 69.380 182.740 ;
        RECT 74.670 182.680 74.810 182.880 ;
        RECT 76.050 182.740 76.190 183.900 ;
        RECT 81.135 183.700 81.425 183.745 ;
        RECT 81.940 183.700 82.260 183.760 ;
        RECT 81.135 183.560 82.260 183.700 ;
        RECT 81.135 183.515 81.425 183.560 ;
        RECT 81.940 183.500 82.260 183.560 ;
        RECT 82.415 183.700 82.705 183.745 ;
        RECT 86.080 183.700 86.400 183.760 ;
        RECT 82.415 183.560 86.400 183.700 ;
        RECT 82.415 183.515 82.705 183.560 ;
        RECT 86.080 183.500 86.400 183.560 ;
        RECT 77.825 183.360 78.115 183.405 ;
        RECT 80.345 183.360 80.635 183.405 ;
        RECT 81.535 183.360 81.825 183.405 ;
        RECT 77.825 183.220 81.825 183.360 ;
        RECT 77.825 183.175 78.115 183.220 ;
        RECT 80.345 183.175 80.635 183.220 ;
        RECT 81.535 183.175 81.825 183.220 ;
        RECT 85.635 183.360 85.925 183.405 ;
        RECT 86.630 183.360 86.770 183.900 ;
        RECT 107.790 183.900 109.845 184.040 ;
        RECT 107.790 183.760 107.930 183.900 ;
        RECT 109.555 183.855 109.845 183.900 ;
        RECT 106.795 183.700 107.085 183.745 ;
        RECT 107.700 183.700 108.020 183.760 ;
        RECT 106.795 183.560 108.020 183.700 ;
        RECT 106.795 183.515 107.085 183.560 ;
        RECT 107.700 183.500 108.020 183.560 ;
        RECT 108.175 183.700 108.465 183.745 ;
        RECT 110.090 183.700 110.230 184.240 ;
        RECT 118.740 184.180 119.060 184.240 ;
        RECT 120.135 184.380 120.425 184.425 ;
        RECT 124.720 184.380 125.040 184.440 ;
        RECT 133.475 184.380 133.765 184.425 ;
        RECT 120.135 184.240 125.040 184.380 ;
        RECT 120.135 184.195 120.425 184.240 ;
        RECT 124.720 184.180 125.040 184.240 ;
        RECT 125.270 184.240 133.765 184.380 ;
        RECT 112.760 184.040 113.080 184.100 ;
        RECT 115.535 184.040 115.825 184.085 ;
        RECT 119.200 184.040 119.520 184.100 ;
        RECT 112.760 183.900 120.810 184.040 ;
        RECT 112.760 183.840 113.080 183.900 ;
        RECT 115.535 183.855 115.825 183.900 ;
        RECT 119.200 183.840 119.520 183.900 ;
        RECT 108.175 183.560 110.230 183.700 ;
        RECT 108.175 183.515 108.465 183.560 ;
        RECT 110.460 183.500 110.780 183.760 ;
        RECT 111.855 183.700 112.145 183.745 ;
        RECT 113.680 183.700 114.000 183.760 ;
        RECT 111.855 183.560 114.000 183.700 ;
        RECT 111.855 183.515 112.145 183.560 ;
        RECT 113.680 183.500 114.000 183.560 ;
        RECT 114.140 183.700 114.460 183.760 ;
        RECT 114.615 183.700 114.905 183.745 ;
        RECT 116.440 183.700 116.760 183.760 ;
        RECT 114.140 183.560 116.760 183.700 ;
        RECT 114.140 183.500 114.460 183.560 ;
        RECT 114.615 183.515 114.905 183.560 ;
        RECT 116.440 183.500 116.760 183.560 ;
        RECT 116.915 183.700 117.205 183.745 ;
        RECT 117.360 183.700 117.680 183.760 ;
        RECT 116.915 183.560 117.680 183.700 ;
        RECT 116.915 183.515 117.205 183.560 ;
        RECT 117.360 183.500 117.680 183.560 ;
        RECT 117.820 183.500 118.140 183.760 ;
        RECT 120.670 183.745 120.810 183.900 ;
        RECT 118.295 183.515 118.585 183.745 ;
        RECT 118.755 183.515 119.045 183.745 ;
        RECT 120.595 183.515 120.885 183.745 ;
        RECT 121.975 183.700 122.265 183.745 ;
        RECT 123.800 183.700 124.120 183.760 ;
        RECT 125.270 183.745 125.410 184.240 ;
        RECT 133.475 184.195 133.765 184.240 ;
        RECT 121.975 183.560 124.120 183.700 ;
        RECT 121.975 183.515 122.265 183.560 ;
        RECT 85.635 183.220 86.770 183.360 ;
        RECT 107.240 183.360 107.560 183.420 ;
        RECT 109.540 183.360 109.860 183.420 ;
        RECT 107.240 183.220 109.860 183.360 ;
        RECT 85.635 183.175 85.925 183.220 ;
        RECT 107.240 183.160 107.560 183.220 ;
        RECT 109.540 183.160 109.860 183.220 ;
        RECT 111.380 183.360 111.700 183.420 ;
        RECT 112.315 183.360 112.605 183.405 ;
        RECT 111.380 183.220 112.605 183.360 ;
        RECT 111.380 183.160 111.700 183.220 ;
        RECT 112.315 183.175 112.605 183.220 ;
        RECT 113.235 183.360 113.525 183.405 ;
        RECT 115.980 183.360 116.300 183.420 ;
        RECT 118.370 183.360 118.510 183.515 ;
        RECT 113.235 183.220 114.370 183.360 ;
        RECT 113.235 183.175 113.525 183.220 ;
        RECT 78.260 183.020 78.550 183.065 ;
        RECT 79.830 183.020 80.120 183.065 ;
        RECT 81.930 183.020 82.220 183.065 ;
        RECT 78.260 182.880 82.220 183.020 ;
        RECT 78.260 182.835 78.550 182.880 ;
        RECT 79.830 182.835 80.120 182.880 ;
        RECT 81.930 182.835 82.220 182.880 ;
        RECT 107.700 182.820 108.020 183.080 ;
        RECT 113.680 183.020 114.000 183.080 ;
        RECT 108.250 182.880 114.000 183.020 ;
        RECT 114.230 183.020 114.370 183.220 ;
        RECT 115.980 183.220 118.510 183.360 ;
        RECT 115.980 183.160 116.300 183.220 ;
        RECT 116.900 183.020 117.220 183.080 ;
        RECT 118.830 183.020 118.970 183.515 ;
        RECT 123.800 183.500 124.120 183.560 ;
        RECT 125.195 183.515 125.485 183.745 ;
        RECT 125.640 183.700 125.960 183.760 ;
        RECT 126.560 183.700 126.880 183.760 ;
        RECT 127.940 183.745 128.260 183.760 ;
        RECT 125.640 183.560 126.880 183.700 ;
        RECT 125.640 183.500 125.960 183.560 ;
        RECT 126.560 183.500 126.880 183.560 ;
        RECT 127.910 183.515 128.260 183.745 ;
        RECT 133.550 183.700 133.690 184.195 ;
        RECT 136.695 183.700 136.985 183.745 ;
        RECT 133.550 183.560 136.985 183.700 ;
        RECT 136.695 183.515 136.985 183.560 ;
        RECT 127.940 183.500 128.260 183.515 ;
        RECT 122.420 183.160 122.740 183.420 ;
        RECT 127.455 183.360 127.745 183.405 ;
        RECT 128.645 183.360 128.935 183.405 ;
        RECT 131.165 183.360 131.455 183.405 ;
        RECT 127.455 183.220 131.455 183.360 ;
        RECT 127.455 183.175 127.745 183.220 ;
        RECT 128.645 183.175 128.935 183.220 ;
        RECT 131.165 183.175 131.455 183.220 ;
        RECT 114.230 182.880 115.750 183.020 ;
        RECT 69.060 182.540 74.810 182.680 ;
        RECT 75.055 182.680 75.345 182.725 ;
        RECT 75.960 182.680 76.280 182.740 ;
        RECT 75.055 182.540 76.280 182.680 ;
        RECT 69.060 182.480 69.380 182.540 ;
        RECT 75.055 182.495 75.345 182.540 ;
        RECT 75.960 182.480 76.280 182.540 ;
        RECT 76.880 182.680 77.200 182.740 ;
        RECT 82.875 182.680 83.165 182.725 ;
        RECT 76.880 182.540 83.165 182.680 ;
        RECT 76.880 182.480 77.200 182.540 ;
        RECT 82.875 182.495 83.165 182.540 ;
        RECT 103.560 182.680 103.880 182.740 ;
        RECT 108.250 182.680 108.390 182.880 ;
        RECT 113.680 182.820 114.000 182.880 ;
        RECT 103.560 182.540 108.390 182.680 ;
        RECT 108.620 182.680 108.940 182.740 ;
        RECT 109.095 182.680 109.385 182.725 ;
        RECT 108.620 182.540 109.385 182.680 ;
        RECT 103.560 182.480 103.880 182.540 ;
        RECT 108.620 182.480 108.940 182.540 ;
        RECT 109.095 182.495 109.385 182.540 ;
        RECT 110.935 182.680 111.225 182.725 ;
        RECT 111.840 182.680 112.160 182.740 ;
        RECT 110.935 182.540 112.160 182.680 ;
        RECT 110.935 182.495 111.225 182.540 ;
        RECT 111.840 182.480 112.160 182.540 ;
        RECT 112.775 182.680 113.065 182.725 ;
        RECT 113.220 182.680 113.540 182.740 ;
        RECT 112.775 182.540 113.540 182.680 ;
        RECT 112.775 182.495 113.065 182.540 ;
        RECT 113.220 182.480 113.540 182.540 ;
        RECT 114.140 182.480 114.460 182.740 ;
        RECT 115.610 182.680 115.750 182.880 ;
        RECT 116.900 182.880 118.970 183.020 ;
        RECT 116.900 182.820 117.220 182.880 ;
        RECT 126.100 182.820 126.420 183.080 ;
        RECT 127.060 183.020 127.350 183.065 ;
        RECT 129.160 183.020 129.450 183.065 ;
        RECT 130.730 183.020 131.020 183.065 ;
        RECT 127.060 182.880 131.020 183.020 ;
        RECT 127.060 182.835 127.350 182.880 ;
        RECT 129.160 182.835 129.450 182.880 ;
        RECT 130.730 182.835 131.020 182.880 ;
        RECT 120.580 182.680 120.900 182.740 ;
        RECT 115.610 182.540 120.900 182.680 ;
        RECT 120.580 182.480 120.900 182.540 ;
        RECT 133.920 182.480 134.240 182.740 ;
        RECT 13.330 181.860 138.910 182.340 ;
        RECT 24.440 181.460 24.760 181.720 ;
        RECT 33.655 181.660 33.945 181.705 ;
        RECT 34.560 181.660 34.880 181.720 ;
        RECT 33.655 181.520 34.880 181.660 ;
        RECT 33.655 181.475 33.945 181.520 ;
        RECT 17.580 181.320 17.870 181.365 ;
        RECT 19.680 181.320 19.970 181.365 ;
        RECT 21.250 181.320 21.540 181.365 ;
        RECT 17.580 181.180 21.540 181.320 ;
        RECT 17.580 181.135 17.870 181.180 ;
        RECT 19.680 181.135 19.970 181.180 ;
        RECT 21.250 181.135 21.540 181.180 ;
        RECT 17.975 180.980 18.265 181.025 ;
        RECT 19.165 180.980 19.455 181.025 ;
        RECT 21.685 180.980 21.975 181.025 ;
        RECT 17.975 180.840 21.975 180.980 ;
        RECT 17.975 180.795 18.265 180.840 ;
        RECT 19.165 180.795 19.455 180.840 ;
        RECT 21.685 180.795 21.975 180.840 ;
        RECT 23.980 180.980 24.300 181.040 ;
        RECT 33.730 180.980 33.870 181.475 ;
        RECT 34.560 181.460 34.880 181.520 ;
        RECT 64.000 181.460 64.320 181.720 ;
        RECT 67.680 181.660 68.000 181.720 ;
        RECT 71.360 181.660 71.680 181.720 ;
        RECT 67.680 181.520 71.680 181.660 ;
        RECT 67.680 181.460 68.000 181.520 ;
        RECT 71.360 181.460 71.680 181.520 ;
        RECT 71.820 181.660 72.140 181.720 ;
        RECT 74.595 181.660 74.885 181.705 ;
        RECT 71.820 181.520 74.885 181.660 ;
        RECT 71.820 181.460 72.140 181.520 ;
        RECT 74.595 181.475 74.885 181.520 ;
        RECT 75.040 181.660 75.360 181.720 ;
        RECT 75.515 181.660 75.805 181.705 ;
        RECT 78.260 181.660 78.580 181.720 ;
        RECT 75.040 181.520 78.580 181.660 ;
        RECT 75.040 181.460 75.360 181.520 ;
        RECT 75.515 181.475 75.805 181.520 ;
        RECT 78.260 181.460 78.580 181.520 ;
        RECT 81.940 181.660 82.260 181.720 ;
        RECT 82.415 181.660 82.705 181.705 ;
        RECT 81.940 181.520 82.705 181.660 ;
        RECT 81.940 181.460 82.260 181.520 ;
        RECT 82.415 181.475 82.705 181.520 ;
        RECT 107.700 181.660 108.020 181.720 ;
        RECT 109.555 181.660 109.845 181.705 ;
        RECT 107.700 181.520 109.845 181.660 ;
        RECT 107.700 181.460 108.020 181.520 ;
        RECT 35.495 181.320 35.785 181.365 ;
        RECT 36.400 181.320 36.720 181.380 ;
        RECT 35.495 181.180 36.720 181.320 ;
        RECT 35.495 181.135 35.785 181.180 ;
        RECT 36.400 181.120 36.720 181.180 ;
        RECT 36.860 181.320 37.180 181.380 ;
        RECT 41.000 181.320 41.320 181.380 ;
        RECT 47.440 181.320 47.730 181.365 ;
        RECT 49.010 181.320 49.300 181.365 ;
        RECT 51.110 181.320 51.400 181.365 ;
        RECT 36.860 181.180 44.450 181.320 ;
        RECT 36.860 181.120 37.180 181.180 ;
        RECT 41.000 181.120 41.320 181.180 ;
        RECT 38.255 180.980 38.545 181.025 ;
        RECT 39.620 180.980 39.940 181.040 ;
        RECT 23.980 180.840 29.270 180.980 ;
        RECT 23.980 180.780 24.300 180.840 ;
        RECT 17.095 180.640 17.385 180.685 ;
        RECT 17.540 180.640 17.860 180.700 ;
        RECT 19.840 180.640 20.160 180.700 ;
        RECT 17.095 180.500 20.160 180.640 ;
        RECT 17.095 180.455 17.385 180.500 ;
        RECT 17.540 180.440 17.860 180.500 ;
        RECT 19.840 180.440 20.160 180.500 ;
        RECT 22.140 180.640 22.460 180.700 ;
        RECT 24.455 180.640 24.745 180.685 ;
        RECT 22.140 180.500 24.745 180.640 ;
        RECT 22.140 180.440 22.460 180.500 ;
        RECT 24.455 180.455 24.745 180.500 ;
        RECT 24.900 180.640 25.220 180.700 ;
        RECT 25.375 180.640 25.665 180.685 ;
        RECT 28.120 180.640 28.440 180.700 ;
        RECT 29.130 180.685 29.270 180.840 ;
        RECT 32.810 180.840 33.870 180.980 ;
        RECT 34.650 180.840 39.940 180.980 ;
        RECT 32.810 180.685 32.950 180.840 ;
        RECT 34.650 180.685 34.790 180.840 ;
        RECT 38.255 180.795 38.545 180.840 ;
        RECT 39.620 180.780 39.940 180.840 ;
        RECT 40.080 180.980 40.400 181.040 ;
        RECT 43.775 180.980 44.065 181.025 ;
        RECT 40.080 180.840 44.065 180.980 ;
        RECT 40.080 180.780 40.400 180.840 ;
        RECT 43.775 180.795 44.065 180.840 ;
        RECT 24.900 180.500 28.440 180.640 ;
        RECT 24.900 180.440 25.220 180.500 ;
        RECT 25.375 180.455 25.665 180.500 ;
        RECT 28.120 180.440 28.440 180.500 ;
        RECT 29.055 180.455 29.345 180.685 ;
        RECT 32.270 180.455 32.560 180.685 ;
        RECT 32.735 180.455 33.025 180.685 ;
        RECT 33.195 180.455 33.485 180.685 ;
        RECT 34.575 180.455 34.865 180.685 ;
        RECT 18.460 180.345 18.780 180.360 ;
        RECT 18.430 180.115 18.780 180.345 ;
        RECT 31.800 180.300 32.120 180.360 ;
        RECT 32.305 180.300 32.445 180.455 ;
        RECT 33.270 180.300 33.410 180.455 ;
        RECT 36.860 180.440 37.180 180.700 ;
        RECT 37.335 180.640 37.625 180.685 ;
        RECT 37.780 180.640 38.100 180.700 ;
        RECT 37.335 180.500 38.100 180.640 ;
        RECT 37.335 180.455 37.625 180.500 ;
        RECT 37.780 180.440 38.100 180.500 ;
        RECT 38.715 180.640 39.005 180.685 ;
        RECT 39.175 180.640 39.465 180.685 ;
        RECT 40.540 180.640 40.860 180.700 ;
        RECT 38.715 180.500 40.860 180.640 ;
        RECT 38.715 180.455 39.005 180.500 ;
        RECT 39.175 180.455 39.465 180.500 ;
        RECT 40.540 180.440 40.860 180.500 ;
        RECT 42.855 180.640 43.145 180.685 ;
        RECT 44.310 180.640 44.450 181.180 ;
        RECT 47.440 181.180 51.400 181.320 ;
        RECT 47.440 181.135 47.730 181.180 ;
        RECT 49.010 181.135 49.300 181.180 ;
        RECT 51.110 181.135 51.400 181.180 ;
        RECT 55.260 181.120 55.580 181.380 ;
        RECT 57.600 181.320 57.890 181.365 ;
        RECT 59.700 181.320 59.990 181.365 ;
        RECT 61.270 181.320 61.560 181.365 ;
        RECT 57.600 181.180 61.560 181.320 ;
        RECT 57.600 181.135 57.890 181.180 ;
        RECT 59.700 181.135 59.990 181.180 ;
        RECT 61.270 181.135 61.560 181.180 ;
        RECT 68.690 181.180 70.670 181.320 ;
        RECT 47.005 180.980 47.295 181.025 ;
        RECT 49.525 180.980 49.815 181.025 ;
        RECT 50.715 180.980 51.005 181.025 ;
        RECT 47.005 180.840 51.005 180.980 ;
        RECT 47.005 180.795 47.295 180.840 ;
        RECT 49.525 180.795 49.815 180.840 ;
        RECT 50.715 180.795 51.005 180.840 ;
        RECT 57.995 180.980 58.285 181.025 ;
        RECT 59.185 180.980 59.475 181.025 ;
        RECT 61.705 180.980 61.995 181.025 ;
        RECT 68.690 180.980 68.830 181.180 ;
        RECT 57.995 180.840 61.995 180.980 ;
        RECT 57.995 180.795 58.285 180.840 ;
        RECT 59.185 180.795 59.475 180.840 ;
        RECT 61.705 180.795 61.995 180.840 ;
        RECT 64.550 180.840 68.830 180.980 ;
        RECT 70.530 180.980 70.670 181.180 ;
        RECT 70.900 181.120 71.220 181.380 ;
        RECT 79.640 181.320 79.960 181.380 ;
        RECT 108.175 181.320 108.465 181.365 ;
        RECT 79.640 181.180 84.010 181.320 ;
        RECT 79.640 181.120 79.960 181.180 ;
        RECT 71.360 180.980 71.680 181.040 ;
        RECT 72.295 180.980 72.585 181.025 ;
        RECT 70.530 180.840 72.585 180.980 ;
        RECT 51.595 180.640 51.885 180.685 ;
        RECT 55.720 180.640 56.040 180.700 ;
        RECT 58.480 180.685 58.800 180.700 ;
        RECT 64.550 180.685 64.690 180.840 ;
        RECT 71.360 180.780 71.680 180.840 ;
        RECT 72.295 180.795 72.585 180.840 ;
        RECT 72.740 180.780 73.060 181.040 ;
        RECT 73.215 180.980 73.505 181.025 ;
        RECT 75.040 180.980 75.360 181.040 ;
        RECT 73.215 180.840 75.360 180.980 ;
        RECT 73.215 180.795 73.505 180.840 ;
        RECT 75.040 180.780 75.360 180.840 ;
        RECT 75.960 180.780 76.280 181.040 ;
        RECT 79.180 180.780 79.500 181.040 ;
        RECT 80.100 180.780 80.420 181.040 ;
        RECT 83.335 180.980 83.625 181.025 ;
        RECT 80.650 180.840 83.625 180.980 ;
        RECT 57.115 180.640 57.405 180.685 ;
        RECT 58.450 180.640 58.800 180.685 ;
        RECT 42.855 180.500 44.450 180.640 ;
        RECT 49.370 180.500 57.405 180.640 ;
        RECT 58.285 180.500 58.800 180.640 ;
        RECT 42.855 180.455 43.145 180.500 ;
        RECT 49.370 180.360 49.510 180.500 ;
        RECT 51.595 180.455 51.885 180.500 ;
        RECT 55.720 180.440 56.040 180.500 ;
        RECT 57.115 180.455 57.405 180.500 ;
        RECT 58.450 180.455 58.800 180.500 ;
        RECT 64.475 180.455 64.765 180.685 ;
        RECT 65.395 180.640 65.685 180.685 ;
        RECT 68.600 180.640 68.920 180.700 ;
        RECT 65.395 180.500 68.920 180.640 ;
        RECT 65.395 180.455 65.685 180.500 ;
        RECT 58.480 180.440 58.800 180.455 ;
        RECT 68.600 180.440 68.920 180.500 ;
        RECT 69.980 180.440 70.300 180.700 ;
        RECT 71.820 180.440 72.140 180.700 ;
        RECT 74.090 180.640 74.380 180.685 ;
        RECT 73.750 180.500 74.380 180.640 ;
        RECT 41.015 180.300 41.305 180.345 ;
        RECT 18.460 180.100 18.780 180.115 ;
        RECT 30.050 180.160 41.305 180.300 ;
        RECT 23.980 179.760 24.300 180.020 ;
        RECT 30.050 180.005 30.190 180.160 ;
        RECT 31.800 180.100 32.120 180.160 ;
        RECT 41.015 180.115 41.305 180.160 ;
        RECT 41.460 180.300 41.780 180.360 ;
        RECT 41.460 180.160 45.370 180.300 ;
        RECT 41.460 180.100 41.780 180.160 ;
        RECT 29.975 179.775 30.265 180.005 ;
        RECT 30.880 179.760 31.200 180.020 ;
        RECT 35.940 179.760 36.260 180.020 ;
        RECT 41.920 179.760 42.240 180.020 ;
        RECT 44.680 179.760 45.000 180.020 ;
        RECT 45.230 179.960 45.370 180.160 ;
        RECT 49.280 180.100 49.600 180.360 ;
        RECT 49.740 180.300 50.060 180.360 ;
        RECT 50.260 180.300 50.550 180.345 ;
        RECT 49.740 180.160 50.550 180.300 ;
        RECT 49.740 180.100 50.060 180.160 ;
        RECT 50.260 180.115 50.550 180.160 ;
        RECT 52.500 180.100 52.820 180.360 ;
        RECT 52.960 180.300 53.280 180.360 ;
        RECT 53.895 180.300 54.185 180.345 ;
        RECT 52.960 180.160 54.185 180.300 ;
        RECT 52.960 180.100 53.280 180.160 ;
        RECT 53.895 180.115 54.185 180.160 ;
        RECT 53.435 179.960 53.725 180.005 ;
        RECT 45.230 179.820 53.725 179.960 ;
        RECT 53.435 179.775 53.725 179.820 ;
        RECT 54.340 179.760 54.660 180.020 ;
        RECT 65.380 179.760 65.700 180.020 ;
        RECT 67.220 179.760 67.540 180.020 ;
        RECT 68.690 179.960 68.830 180.440 ;
        RECT 73.750 179.960 73.890 180.500 ;
        RECT 74.090 180.455 74.380 180.500 ;
        RECT 76.420 180.640 76.740 180.700 ;
        RECT 77.355 180.640 77.645 180.685 ;
        RECT 80.650 180.640 80.790 180.840 ;
        RECT 83.335 180.795 83.625 180.840 ;
        RECT 76.420 180.500 80.790 180.640 ;
        RECT 76.420 180.440 76.740 180.500 ;
        RECT 77.355 180.455 77.645 180.500 ;
        RECT 82.860 180.440 83.180 180.700 ;
        RECT 83.870 180.685 84.010 181.180 ;
        RECT 93.990 181.180 108.465 181.320 ;
        RECT 93.990 181.025 94.130 181.180 ;
        RECT 108.175 181.135 108.465 181.180 ;
        RECT 93.915 180.795 94.205 181.025 ;
        RECT 94.820 180.980 95.140 181.040 ;
        RECT 98.975 180.980 99.265 181.025 ;
        RECT 94.820 180.840 99.265 180.980 ;
        RECT 94.820 180.780 95.140 180.840 ;
        RECT 98.975 180.795 99.265 180.840 ;
        RECT 103.100 180.980 103.420 181.040 ;
        RECT 108.710 180.980 108.850 181.520 ;
        RECT 109.555 181.475 109.845 181.520 ;
        RECT 111.380 181.460 111.700 181.720 ;
        RECT 113.680 181.660 114.000 181.720 ;
        RECT 112.850 181.520 114.000 181.660 ;
        RECT 110.920 181.320 111.240 181.380 ;
        RECT 112.850 181.320 112.990 181.520 ;
        RECT 113.680 181.460 114.000 181.520 ;
        RECT 116.915 181.660 117.205 181.705 ;
        RECT 119.200 181.660 119.520 181.720 ;
        RECT 116.915 181.520 119.520 181.660 ;
        RECT 116.915 181.475 117.205 181.520 ;
        RECT 119.200 181.460 119.520 181.520 ;
        RECT 124.735 181.660 125.025 181.705 ;
        RECT 127.480 181.660 127.800 181.720 ;
        RECT 124.735 181.520 127.800 181.660 ;
        RECT 124.735 181.475 125.025 181.520 ;
        RECT 127.480 181.460 127.800 181.520 ;
        RECT 127.940 181.660 128.260 181.720 ;
        RECT 128.875 181.660 129.165 181.705 ;
        RECT 127.940 181.520 129.165 181.660 ;
        RECT 127.940 181.460 128.260 181.520 ;
        RECT 128.875 181.475 129.165 181.520 ;
        RECT 110.090 181.180 111.240 181.320 ;
        RECT 110.090 181.025 110.230 181.180 ;
        RECT 110.920 181.120 111.240 181.180 ;
        RECT 111.470 181.180 112.990 181.320 ;
        RECT 103.100 180.840 108.850 180.980 ;
        RECT 103.100 180.780 103.420 180.840 ;
        RECT 83.795 180.455 84.085 180.685 ;
        RECT 92.995 180.640 93.285 180.685 ;
        RECT 94.360 180.640 94.680 180.700 ;
        RECT 92.995 180.500 94.680 180.640 ;
        RECT 92.995 180.455 93.285 180.500 ;
        RECT 94.360 180.440 94.680 180.500 ;
        RECT 95.280 180.640 95.600 180.700 ;
        RECT 105.030 180.685 105.170 180.840 ;
        RECT 110.015 180.795 110.305 181.025 ;
        RECT 98.055 180.640 98.345 180.685 ;
        RECT 95.280 180.500 98.345 180.640 ;
        RECT 95.280 180.440 95.600 180.500 ;
        RECT 98.055 180.455 98.345 180.500 ;
        RECT 104.955 180.455 105.245 180.685 ;
        RECT 105.415 180.455 105.705 180.685 ;
        RECT 80.575 180.300 80.865 180.345 ;
        RECT 103.560 180.300 103.880 180.360 ;
        RECT 105.490 180.300 105.630 180.455 ;
        RECT 106.320 180.440 106.640 180.700 ;
        RECT 107.240 180.440 107.560 180.700 ;
        RECT 107.715 180.455 108.005 180.685 ;
        RECT 80.575 180.160 84.010 180.300 ;
        RECT 80.575 180.115 80.865 180.160 ;
        RECT 83.870 180.020 84.010 180.160 ;
        RECT 103.560 180.160 105.630 180.300 ;
        RECT 107.790 180.300 107.930 180.455 ;
        RECT 108.620 180.440 108.940 180.700 ;
        RECT 109.540 180.440 109.860 180.700 ;
        RECT 110.920 180.640 111.240 180.700 ;
        RECT 111.470 180.640 111.610 181.180 ;
        RECT 112.850 180.980 112.990 181.180 ;
        RECT 114.600 181.320 114.920 181.380 ;
        RECT 115.980 181.320 116.300 181.380 ;
        RECT 114.600 181.180 116.300 181.320 ;
        RECT 114.600 181.120 114.920 181.180 ;
        RECT 115.980 181.120 116.300 181.180 ;
        RECT 130.280 181.320 130.570 181.365 ;
        RECT 132.380 181.320 132.670 181.365 ;
        RECT 133.950 181.320 134.240 181.365 ;
        RECT 130.280 181.180 134.240 181.320 ;
        RECT 130.280 181.135 130.570 181.180 ;
        RECT 132.380 181.135 132.670 181.180 ;
        RECT 133.950 181.135 134.240 181.180 ;
        RECT 113.695 180.980 113.985 181.025 ;
        RECT 112.850 180.840 113.985 180.980 ;
        RECT 113.695 180.795 113.985 180.840 ;
        RECT 115.535 180.980 115.825 181.025 ;
        RECT 125.655 180.980 125.945 181.025 ;
        RECT 115.535 180.840 125.945 180.980 ;
        RECT 115.535 180.795 115.825 180.840 ;
        RECT 125.655 180.795 125.945 180.840 ;
        RECT 126.560 180.980 126.880 181.040 ;
        RECT 129.795 180.980 130.085 181.025 ;
        RECT 126.560 180.840 130.085 180.980 ;
        RECT 126.560 180.780 126.880 180.840 ;
        RECT 129.795 180.795 130.085 180.840 ;
        RECT 130.675 180.980 130.965 181.025 ;
        RECT 131.865 180.980 132.155 181.025 ;
        RECT 134.385 180.980 134.675 181.025 ;
        RECT 130.675 180.840 134.675 180.980 ;
        RECT 130.675 180.795 130.965 180.840 ;
        RECT 131.865 180.795 132.155 180.840 ;
        RECT 134.385 180.795 134.675 180.840 ;
        RECT 110.920 180.500 111.610 180.640 ;
        RECT 110.920 180.440 111.240 180.500 ;
        RECT 111.840 180.440 112.160 180.700 ;
        RECT 112.760 180.440 113.080 180.700 ;
        RECT 113.235 180.650 113.525 180.685 ;
        RECT 114.140 180.650 114.460 180.700 ;
        RECT 113.235 180.510 114.460 180.650 ;
        RECT 113.235 180.455 113.525 180.510 ;
        RECT 114.140 180.440 114.460 180.510 ;
        RECT 114.600 180.440 114.920 180.700 ;
        RECT 115.995 180.640 116.285 180.685 ;
        RECT 116.440 180.640 116.760 180.700 ;
        RECT 115.995 180.500 116.760 180.640 ;
        RECT 115.995 180.455 116.285 180.500 ;
        RECT 116.440 180.440 116.760 180.500 ;
        RECT 116.915 180.640 117.205 180.685 ;
        RECT 120.135 180.640 120.425 180.685 ;
        RECT 121.975 180.640 122.265 180.685 ;
        RECT 116.915 180.500 119.430 180.640 ;
        RECT 116.915 180.455 117.205 180.500 ;
        RECT 119.290 180.360 119.430 180.500 ;
        RECT 120.135 180.500 122.265 180.640 ;
        RECT 120.135 180.455 120.425 180.500 ;
        RECT 121.975 180.455 122.265 180.500 ;
        RECT 122.420 180.640 122.740 180.700 ;
        RECT 122.895 180.640 123.185 180.685 ;
        RECT 122.420 180.500 123.185 180.640 ;
        RECT 122.420 180.440 122.740 180.500 ;
        RECT 122.895 180.455 123.185 180.500 ;
        RECT 123.800 180.440 124.120 180.700 ;
        RECT 127.035 180.640 127.325 180.685 ;
        RECT 133.920 180.640 134.240 180.700 ;
        RECT 127.035 180.500 134.240 180.640 ;
        RECT 127.035 180.455 127.325 180.500 ;
        RECT 133.920 180.440 134.240 180.500 ;
        RECT 111.380 180.300 111.700 180.360 ;
        RECT 115.520 180.300 115.840 180.360 ;
        RECT 118.295 180.300 118.585 180.345 ;
        RECT 107.790 180.160 111.700 180.300 ;
        RECT 103.560 180.100 103.880 180.160 ;
        RECT 111.380 180.100 111.700 180.160 ;
        RECT 115.175 180.160 118.585 180.300 ;
        RECT 68.690 179.820 73.890 179.960 ;
        RECT 83.780 179.760 84.100 180.020 ;
        RECT 91.140 179.760 91.460 180.020 ;
        RECT 93.455 179.960 93.745 180.005 ;
        RECT 95.295 179.960 95.585 180.005 ;
        RECT 93.455 179.820 95.585 179.960 ;
        RECT 93.455 179.775 93.745 179.820 ;
        RECT 95.295 179.775 95.585 179.820 ;
        RECT 101.260 179.960 101.580 180.020 ;
        RECT 102.195 179.960 102.485 180.005 ;
        RECT 101.260 179.820 102.485 179.960 ;
        RECT 101.260 179.760 101.580 179.820 ;
        RECT 102.195 179.775 102.485 179.820 ;
        RECT 104.940 179.960 105.260 180.020 ;
        RECT 105.415 179.960 105.705 180.005 ;
        RECT 104.940 179.820 105.705 179.960 ;
        RECT 104.940 179.760 105.260 179.820 ;
        RECT 105.415 179.775 105.705 179.820 ;
        RECT 106.780 179.960 107.100 180.020 ;
        RECT 115.175 179.960 115.315 180.160 ;
        RECT 115.520 180.100 115.840 180.160 ;
        RECT 118.295 180.115 118.585 180.160 ;
        RECT 119.200 180.300 119.520 180.360 ;
        RECT 120.580 180.300 120.900 180.360 ;
        RECT 131.160 180.345 131.480 180.360 ;
        RECT 119.200 180.160 120.900 180.300 ;
        RECT 119.200 180.100 119.520 180.160 ;
        RECT 120.580 180.100 120.900 180.160 ;
        RECT 123.355 180.115 123.645 180.345 ;
        RECT 131.130 180.115 131.480 180.345 ;
        RECT 106.780 179.820 115.315 179.960 ;
        RECT 106.780 179.760 107.100 179.820 ;
        RECT 117.820 179.760 118.140 180.020 ;
        RECT 121.040 179.960 121.360 180.020 ;
        RECT 123.430 179.960 123.570 180.115 ;
        RECT 131.160 180.100 131.480 180.115 ;
        RECT 121.040 179.820 123.570 179.960 ;
        RECT 126.100 179.960 126.420 180.020 ;
        RECT 126.575 179.960 126.865 180.005 ;
        RECT 126.100 179.820 126.865 179.960 ;
        RECT 121.040 179.760 121.360 179.820 ;
        RECT 126.100 179.760 126.420 179.820 ;
        RECT 126.575 179.775 126.865 179.820 ;
        RECT 136.680 179.760 137.000 180.020 ;
        RECT 13.330 179.140 138.910 179.620 ;
        RECT 18.015 178.940 18.305 178.985 ;
        RECT 18.460 178.940 18.780 179.000 ;
        RECT 18.015 178.800 18.780 178.940 ;
        RECT 18.015 178.755 18.305 178.800 ;
        RECT 18.460 178.740 18.780 178.800 ;
        RECT 19.380 178.740 19.700 179.000 ;
        RECT 19.840 178.940 20.160 179.000 ;
        RECT 44.680 178.940 45.000 179.000 ;
        RECT 54.340 178.940 54.660 179.000 ;
        RECT 70.440 178.940 70.760 179.000 ;
        RECT 72.280 178.940 72.600 179.000 ;
        RECT 72.755 178.940 73.045 178.985 ;
        RECT 19.840 178.800 34.790 178.940 ;
        RECT 19.840 178.740 20.160 178.800 ;
        RECT 21.680 178.600 22.000 178.660 ;
        RECT 22.455 178.600 22.745 178.645 ;
        RECT 21.680 178.460 22.745 178.600 ;
        RECT 21.680 178.400 22.000 178.460 ;
        RECT 22.455 178.415 22.745 178.460 ;
        RECT 23.535 178.600 23.825 178.645 ;
        RECT 23.980 178.600 24.300 178.660 ;
        RECT 24.915 178.600 25.205 178.645 ;
        RECT 23.535 178.460 25.205 178.600 ;
        RECT 23.535 178.415 23.825 178.460 ;
        RECT 23.980 178.400 24.300 178.460 ;
        RECT 24.915 178.415 25.205 178.460 ;
        RECT 26.740 178.400 27.060 178.660 ;
        RECT 28.120 178.600 28.440 178.660 ;
        RECT 34.650 178.645 34.790 178.800 ;
        RECT 44.680 178.800 56.870 178.940 ;
        RECT 44.680 178.740 45.000 178.800 ;
        RECT 54.340 178.740 54.660 178.800 ;
        RECT 34.575 178.600 34.865 178.645 ;
        RECT 49.280 178.600 49.600 178.660 ;
        RECT 51.135 178.600 51.425 178.645 ;
        RECT 52.960 178.600 53.280 178.660 ;
        RECT 28.120 178.460 32.030 178.600 ;
        RECT 28.120 178.400 28.440 178.460 ;
        RECT 16.635 178.075 16.925 178.305 ;
        RECT 16.710 177.580 16.850 178.075 ;
        RECT 17.540 178.060 17.860 178.320 ;
        RECT 19.855 178.260 20.145 178.305 ;
        RECT 20.300 178.260 20.620 178.320 ;
        RECT 19.855 178.120 20.620 178.260 ;
        RECT 19.855 178.075 20.145 178.120 ;
        RECT 20.300 178.060 20.620 178.120 ;
        RECT 21.220 178.060 21.540 178.320 ;
        RECT 25.375 178.075 25.665 178.305 ;
        RECT 17.095 177.920 17.385 177.965 ;
        RECT 18.810 177.920 19.100 177.965 ;
        RECT 17.095 177.780 19.100 177.920 ;
        RECT 17.095 177.735 17.385 177.780 ;
        RECT 18.810 177.735 19.100 177.780 ;
        RECT 23.995 177.920 24.285 177.965 ;
        RECT 24.900 177.920 25.220 177.980 ;
        RECT 23.995 177.780 25.220 177.920 ;
        RECT 23.995 177.735 24.285 177.780 ;
        RECT 24.900 177.720 25.220 177.780 ;
        RECT 21.695 177.580 21.985 177.625 ;
        RECT 22.140 177.580 22.460 177.640 ;
        RECT 16.710 177.440 22.460 177.580 ;
        RECT 21.695 177.395 21.985 177.440 ;
        RECT 22.140 177.380 22.460 177.440 ;
        RECT 18.920 177.240 19.240 177.300 ;
        RECT 22.615 177.240 22.905 177.285 ;
        RECT 25.450 177.240 25.590 178.075 ;
        RECT 25.820 178.060 26.140 178.320 ;
        RECT 29.975 178.260 30.265 178.305 ;
        RECT 30.420 178.260 30.740 178.320 ;
        RECT 29.975 178.120 30.740 178.260 ;
        RECT 29.975 178.075 30.265 178.120 ;
        RECT 30.420 178.060 30.740 178.120 ;
        RECT 30.880 178.060 31.200 178.320 ;
        RECT 31.340 178.060 31.660 178.320 ;
        RECT 31.890 178.305 32.030 178.460 ;
        RECT 34.575 178.460 39.850 178.600 ;
        RECT 34.575 178.415 34.865 178.460 ;
        RECT 39.710 178.305 39.850 178.460 ;
        RECT 49.280 178.460 53.280 178.600 ;
        RECT 49.280 178.400 49.600 178.460 ;
        RECT 51.135 178.415 51.425 178.460 ;
        RECT 52.960 178.400 53.280 178.460 ;
        RECT 53.420 178.600 53.740 178.660 ;
        RECT 53.420 178.460 55.950 178.600 ;
        RECT 53.420 178.400 53.740 178.460 ;
        RECT 55.810 178.305 55.950 178.460 ;
        RECT 56.730 178.305 56.870 178.800 ;
        RECT 70.440 178.800 72.050 178.940 ;
        RECT 70.440 178.740 70.760 178.800 ;
        RECT 69.980 178.600 70.300 178.660 ;
        RECT 70.900 178.645 71.220 178.660 ;
        RECT 70.900 178.600 71.250 178.645 ;
        RECT 71.910 178.600 72.050 178.800 ;
        RECT 72.280 178.800 73.045 178.940 ;
        RECT 72.280 178.740 72.600 178.800 ;
        RECT 72.755 178.755 73.045 178.800 ;
        RECT 74.595 178.940 74.885 178.985 ;
        RECT 76.880 178.940 77.200 179.000 ;
        RECT 74.595 178.800 77.200 178.940 ;
        RECT 74.595 178.755 74.885 178.800 ;
        RECT 76.880 178.740 77.200 178.800 ;
        RECT 77.800 178.740 78.120 179.000 ;
        RECT 83.780 178.740 84.100 179.000 ;
        RECT 86.095 178.940 86.385 178.985 ;
        RECT 91.155 178.940 91.445 178.985 ;
        RECT 94.820 178.940 95.140 179.000 ;
        RECT 86.095 178.800 95.140 178.940 ;
        RECT 86.095 178.755 86.385 178.800 ;
        RECT 91.155 178.755 91.445 178.800 ;
        RECT 94.820 178.740 95.140 178.800 ;
        RECT 98.515 178.755 98.805 178.985 ;
        RECT 106.780 178.940 107.100 179.000 ;
        RECT 99.510 178.800 107.100 178.940 ;
        RECT 76.435 178.600 76.725 178.645 ;
        RECT 69.980 178.460 70.670 178.600 ;
        RECT 69.980 178.400 70.300 178.460 ;
        RECT 31.815 178.075 32.105 178.305 ;
        RECT 38.715 178.075 39.005 178.305 ;
        RECT 39.635 178.075 39.925 178.305 ;
        RECT 55.275 178.075 55.565 178.305 ;
        RECT 55.735 178.075 56.025 178.305 ;
        RECT 56.655 178.075 56.945 178.305 ;
        RECT 70.530 178.260 70.670 178.460 ;
        RECT 70.900 178.460 71.415 178.600 ;
        RECT 71.910 178.460 76.725 178.600 ;
        RECT 70.900 178.415 71.250 178.460 ;
        RECT 76.435 178.415 76.725 178.460 ;
        RECT 77.355 178.600 77.645 178.645 ;
        RECT 78.260 178.600 78.580 178.660 ;
        RECT 82.860 178.600 83.180 178.660 ;
        RECT 77.355 178.460 78.580 178.600 ;
        RECT 77.355 178.415 77.645 178.460 ;
        RECT 70.900 178.400 71.220 178.415 ;
        RECT 78.260 178.400 78.580 178.460 ;
        RECT 78.810 178.460 83.180 178.600 ;
        RECT 70.530 178.120 72.970 178.260 ;
        RECT 30.510 177.920 30.650 178.060 ;
        RECT 33.180 177.920 33.500 177.980 ;
        RECT 30.510 177.780 33.500 177.920 ;
        RECT 38.790 177.920 38.930 178.075 ;
        RECT 55.350 177.920 55.490 178.075 ;
        RECT 60.320 177.920 60.640 177.980 ;
        RECT 38.790 177.780 60.640 177.920 ;
        RECT 33.180 177.720 33.500 177.780 ;
        RECT 60.320 177.720 60.640 177.780 ;
        RECT 67.705 177.920 67.995 177.965 ;
        RECT 70.225 177.920 70.515 177.965 ;
        RECT 71.415 177.920 71.705 177.965 ;
        RECT 67.705 177.780 71.705 177.920 ;
        RECT 67.705 177.735 67.995 177.780 ;
        RECT 70.225 177.735 70.515 177.780 ;
        RECT 71.415 177.735 71.705 177.780 ;
        RECT 72.280 177.720 72.600 177.980 ;
        RECT 72.830 177.920 72.970 178.120 ;
        RECT 73.660 178.060 73.980 178.320 ;
        RECT 75.040 178.060 75.360 178.320 ;
        RECT 75.500 178.260 75.820 178.320 ;
        RECT 78.810 178.305 78.950 178.460 ;
        RECT 82.860 178.400 83.180 178.460 ;
        RECT 96.830 178.600 97.120 178.645 ;
        RECT 98.590 178.600 98.730 178.755 ;
        RECT 96.830 178.460 98.730 178.600 ;
        RECT 96.830 178.415 97.120 178.460 ;
        RECT 78.735 178.260 79.025 178.305 ;
        RECT 75.500 178.120 79.025 178.260 ;
        RECT 75.500 178.060 75.820 178.120 ;
        RECT 78.735 178.075 79.025 178.120 ;
        RECT 79.640 178.060 79.960 178.320 ;
        RECT 84.700 178.260 85.020 178.320 ;
        RECT 85.635 178.260 85.925 178.305 ;
        RECT 94.360 178.260 94.680 178.320 ;
        RECT 99.510 178.305 99.650 178.800 ;
        RECT 106.780 178.740 107.100 178.800 ;
        RECT 110.920 178.940 111.240 179.000 ;
        RECT 112.775 178.940 113.065 178.985 ;
        RECT 110.920 178.800 113.065 178.940 ;
        RECT 110.920 178.740 111.240 178.800 ;
        RECT 112.775 178.755 113.065 178.800 ;
        RECT 114.600 178.740 114.920 179.000 ;
        RECT 122.420 178.940 122.740 179.000 ;
        RECT 122.050 178.800 122.740 178.940 ;
        RECT 100.355 178.600 100.645 178.645 ;
        RECT 101.735 178.600 102.025 178.645 ;
        RECT 104.940 178.600 105.260 178.660 ;
        RECT 118.740 178.600 119.060 178.660 ;
        RECT 122.050 178.645 122.190 178.800 ;
        RECT 122.420 178.740 122.740 178.800 ;
        RECT 123.340 178.940 123.660 179.000 ;
        RECT 126.100 178.940 126.420 179.000 ;
        RECT 127.035 178.940 127.325 178.985 ;
        RECT 123.340 178.800 125.870 178.940 ;
        RECT 123.340 178.740 123.660 178.800 ;
        RECT 100.355 178.460 102.025 178.600 ;
        RECT 100.355 178.415 100.645 178.460 ;
        RECT 101.735 178.415 102.025 178.460 ;
        RECT 102.270 178.460 105.260 178.600 ;
        RECT 84.700 178.120 85.925 178.260 ;
        RECT 84.700 178.060 85.020 178.120 ;
        RECT 85.635 178.075 85.925 178.120 ;
        RECT 87.090 178.120 94.680 178.260 ;
        RECT 79.730 177.920 79.870 178.060 ;
        RECT 72.830 177.780 79.870 177.920 ;
        RECT 80.100 177.720 80.420 177.980 ;
        RECT 87.090 177.965 87.230 178.120 ;
        RECT 94.360 178.060 94.680 178.120 ;
        RECT 99.435 178.075 99.725 178.305 ;
        RECT 99.895 178.075 100.185 178.305 ;
        RECT 87.015 177.735 87.305 177.965 ;
        RECT 93.465 177.920 93.755 177.965 ;
        RECT 95.985 177.920 96.275 177.965 ;
        RECT 97.175 177.920 97.465 177.965 ;
        RECT 93.465 177.780 97.465 177.920 ;
        RECT 93.465 177.735 93.755 177.780 ;
        RECT 95.985 177.735 96.275 177.780 ;
        RECT 97.175 177.735 97.465 177.780 ;
        RECT 98.040 177.720 98.360 177.980 ;
        RECT 99.970 177.920 100.110 178.075 ;
        RECT 101.260 178.060 101.580 178.320 ;
        RECT 102.270 177.920 102.410 178.460 ;
        RECT 104.940 178.400 105.260 178.460 ;
        RECT 114.690 178.460 119.060 178.600 ;
        RECT 102.655 178.075 102.945 178.305 ;
        RECT 103.115 178.075 103.405 178.305 ;
        RECT 99.970 177.780 102.410 177.920 ;
        RECT 68.140 177.580 68.430 177.625 ;
        RECT 69.710 177.580 70.000 177.625 ;
        RECT 71.810 177.580 72.100 177.625 ;
        RECT 74.580 177.580 74.900 177.640 ;
        RECT 68.140 177.440 72.100 177.580 ;
        RECT 68.140 177.395 68.430 177.440 ;
        RECT 69.710 177.395 70.000 177.440 ;
        RECT 71.810 177.395 72.100 177.440 ;
        RECT 72.370 177.440 74.900 177.580 ;
        RECT 18.920 177.100 25.590 177.240 ;
        RECT 33.195 177.240 33.485 177.285 ;
        RECT 33.640 177.240 33.960 177.300 ;
        RECT 33.195 177.100 33.960 177.240 ;
        RECT 18.920 177.040 19.240 177.100 ;
        RECT 22.615 177.055 22.905 177.100 ;
        RECT 33.195 177.055 33.485 177.100 ;
        RECT 33.640 177.040 33.960 177.100 ;
        RECT 51.120 177.240 51.440 177.300 ;
        RECT 55.735 177.240 56.025 177.285 ;
        RECT 51.120 177.100 56.025 177.240 ;
        RECT 51.120 177.040 51.440 177.100 ;
        RECT 55.735 177.055 56.025 177.100 ;
        RECT 65.395 177.240 65.685 177.285 ;
        RECT 70.440 177.240 70.760 177.300 ;
        RECT 72.370 177.240 72.510 177.440 ;
        RECT 74.580 177.380 74.900 177.440 ;
        RECT 83.335 177.580 83.625 177.625 ;
        RECT 84.240 177.580 84.560 177.640 ;
        RECT 83.335 177.440 84.560 177.580 ;
        RECT 83.335 177.395 83.625 177.440 ;
        RECT 84.240 177.380 84.560 177.440 ;
        RECT 93.900 177.580 94.190 177.625 ;
        RECT 95.470 177.580 95.760 177.625 ;
        RECT 97.570 177.580 97.860 177.625 ;
        RECT 93.900 177.440 97.860 177.580 ;
        RECT 102.730 177.580 102.870 178.075 ;
        RECT 103.190 177.920 103.330 178.075 ;
        RECT 104.020 178.060 104.340 178.320 ;
        RECT 104.480 178.260 104.800 178.320 ;
        RECT 106.320 178.260 106.640 178.320 ;
        RECT 104.480 178.120 106.640 178.260 ;
        RECT 104.480 178.060 104.800 178.120 ;
        RECT 106.320 178.060 106.640 178.120 ;
        RECT 108.620 178.260 108.940 178.320 ;
        RECT 110.475 178.260 110.765 178.305 ;
        RECT 108.620 178.120 110.765 178.260 ;
        RECT 108.620 178.060 108.940 178.120 ;
        RECT 110.475 178.075 110.765 178.120 ;
        RECT 110.935 178.075 111.225 178.305 ;
        RECT 112.315 178.260 112.605 178.305 ;
        RECT 112.315 178.120 112.990 178.260 ;
        RECT 112.315 178.075 112.605 178.120 ;
        RECT 107.240 177.920 107.560 177.980 ;
        RECT 103.190 177.780 107.560 177.920 ;
        RECT 107.240 177.720 107.560 177.780 ;
        RECT 106.780 177.580 107.100 177.640 ;
        RECT 102.730 177.440 107.100 177.580 ;
        RECT 93.900 177.395 94.190 177.440 ;
        RECT 95.470 177.395 95.760 177.440 ;
        RECT 97.570 177.395 97.860 177.440 ;
        RECT 106.780 177.380 107.100 177.440 ;
        RECT 110.460 177.580 110.780 177.640 ;
        RECT 111.010 177.580 111.150 178.075 ;
        RECT 111.380 177.920 111.700 177.980 ;
        RECT 111.855 177.920 112.145 177.965 ;
        RECT 111.380 177.780 112.145 177.920 ;
        RECT 111.380 177.720 111.700 177.780 ;
        RECT 111.855 177.735 112.145 177.780 ;
        RECT 110.460 177.440 111.150 177.580 ;
        RECT 112.850 177.580 112.990 178.120 ;
        RECT 113.695 178.250 113.985 178.305 ;
        RECT 114.690 178.260 114.830 178.460 ;
        RECT 118.740 178.400 119.060 178.460 ;
        RECT 121.975 178.600 122.265 178.645 ;
        RECT 125.195 178.600 125.485 178.645 ;
        RECT 121.975 178.460 125.485 178.600 ;
        RECT 125.730 178.600 125.870 178.800 ;
        RECT 126.100 178.800 127.325 178.940 ;
        RECT 126.100 178.740 126.420 178.800 ;
        RECT 127.035 178.755 127.325 178.800 ;
        RECT 131.160 178.740 131.480 179.000 ;
        RECT 132.555 178.940 132.845 178.985 ;
        RECT 135.760 178.940 136.080 179.000 ;
        RECT 132.555 178.800 136.080 178.940 ;
        RECT 132.555 178.755 132.845 178.800 ;
        RECT 135.760 178.740 136.080 178.800 ;
        RECT 129.335 178.600 129.625 178.645 ;
        RECT 133.015 178.600 133.305 178.645 ;
        RECT 125.730 178.460 126.330 178.600 ;
        RECT 121.975 178.415 122.265 178.460 ;
        RECT 125.195 178.415 125.485 178.460 ;
        RECT 114.230 178.250 114.830 178.260 ;
        RECT 113.695 178.120 114.830 178.250 ;
        RECT 115.075 178.260 115.365 178.305 ;
        RECT 115.980 178.260 116.300 178.320 ;
        RECT 115.075 178.120 116.300 178.260 ;
        RECT 113.695 178.110 114.370 178.120 ;
        RECT 113.695 178.075 113.985 178.110 ;
        RECT 115.075 178.075 115.365 178.120 ;
        RECT 115.980 178.060 116.300 178.120 ;
        RECT 116.915 178.260 117.205 178.305 ;
        RECT 117.360 178.260 117.680 178.320 ;
        RECT 116.915 178.120 117.680 178.260 ;
        RECT 116.915 178.075 117.205 178.120 ;
        RECT 117.360 178.060 117.680 178.120 ;
        RECT 117.835 178.075 118.125 178.305 ;
        RECT 113.220 177.920 113.540 177.980 ;
        RECT 117.910 177.920 118.050 178.075 ;
        RECT 118.280 178.060 118.600 178.320 ;
        RECT 119.675 178.075 119.965 178.305 ;
        RECT 120.120 178.260 120.440 178.320 ;
        RECT 121.055 178.260 121.345 178.305 ;
        RECT 122.435 178.260 122.725 178.305 ;
        RECT 120.120 178.120 121.345 178.260 ;
        RECT 113.220 177.780 118.050 177.920 ;
        RECT 113.220 177.720 113.540 177.780 ;
        RECT 118.740 177.720 119.060 177.980 ;
        RECT 114.140 177.580 114.460 177.640 ;
        RECT 117.820 177.580 118.140 177.640 ;
        RECT 119.750 177.580 119.890 178.075 ;
        RECT 120.120 178.060 120.440 178.120 ;
        RECT 121.055 178.075 121.345 178.120 ;
        RECT 122.050 178.120 122.725 178.260 ;
        RECT 122.050 177.980 122.190 178.120 ;
        RECT 122.435 178.075 122.725 178.120 ;
        RECT 122.895 178.260 123.185 178.305 ;
        RECT 123.340 178.260 123.660 178.320 ;
        RECT 122.895 178.120 123.660 178.260 ;
        RECT 122.895 178.075 123.185 178.120 ;
        RECT 123.340 178.060 123.660 178.120 ;
        RECT 124.260 178.060 124.580 178.320 ;
        RECT 125.640 178.060 125.960 178.320 ;
        RECT 126.190 178.305 126.330 178.460 ;
        RECT 129.335 178.460 133.305 178.600 ;
        RECT 129.335 178.415 129.625 178.460 ;
        RECT 133.015 178.415 133.305 178.460 ;
        RECT 126.115 178.075 126.405 178.305 ;
        RECT 131.635 178.260 131.925 178.305 ;
        RECT 136.235 178.260 136.525 178.305 ;
        RECT 136.680 178.260 137.000 178.320 ;
        RECT 131.635 178.120 137.000 178.260 ;
        RECT 131.635 178.075 131.925 178.120 ;
        RECT 136.235 178.075 136.525 178.120 ;
        RECT 136.680 178.060 137.000 178.120 ;
        RECT 121.960 177.720 122.280 177.980 ;
        RECT 127.955 177.920 128.245 177.965 ;
        RECT 123.430 177.780 128.245 177.920 ;
        RECT 112.850 177.440 119.890 177.580 ;
        RECT 120.595 177.580 120.885 177.625 ;
        RECT 123.430 177.580 123.570 177.780 ;
        RECT 127.955 177.735 128.245 177.780 ;
        RECT 128.875 177.735 129.165 177.965 ;
        RECT 120.595 177.440 123.570 177.580 ;
        RECT 123.815 177.580 124.105 177.625 ;
        RECT 128.950 177.580 129.090 177.735 ;
        RECT 123.815 177.440 129.090 177.580 ;
        RECT 110.460 177.380 110.780 177.440 ;
        RECT 65.395 177.100 72.510 177.240 ;
        RECT 72.740 177.240 73.060 177.300 ;
        RECT 75.040 177.240 75.360 177.300 ;
        RECT 75.515 177.240 75.805 177.285 ;
        RECT 72.740 177.100 75.805 177.240 ;
        RECT 65.395 177.055 65.685 177.100 ;
        RECT 70.440 177.040 70.760 177.100 ;
        RECT 72.740 177.040 73.060 177.100 ;
        RECT 75.040 177.040 75.360 177.100 ;
        RECT 75.515 177.055 75.805 177.100 ;
        RECT 79.180 177.240 79.500 177.300 ;
        RECT 83.780 177.240 84.100 177.300 ;
        RECT 79.180 177.100 84.100 177.240 ;
        RECT 79.180 177.040 79.500 177.100 ;
        RECT 83.780 177.040 84.100 177.100 ;
        RECT 109.540 177.040 109.860 177.300 ;
        RECT 111.010 177.240 111.150 177.440 ;
        RECT 114.140 177.380 114.460 177.440 ;
        RECT 117.820 177.380 118.140 177.440 ;
        RECT 120.595 177.395 120.885 177.440 ;
        RECT 123.815 177.395 124.105 177.440 ;
        RECT 123.340 177.240 123.660 177.300 ;
        RECT 111.010 177.100 123.660 177.240 ;
        RECT 123.340 177.040 123.660 177.100 ;
        RECT 13.330 176.420 138.910 176.900 ;
        RECT 17.540 176.220 17.860 176.280 ;
        RECT 22.615 176.220 22.905 176.265 ;
        RECT 17.540 176.080 22.905 176.220 ;
        RECT 17.540 176.020 17.860 176.080 ;
        RECT 22.615 176.035 22.905 176.080 ;
        RECT 23.980 176.220 24.300 176.280 ;
        RECT 26.740 176.220 27.060 176.280 ;
        RECT 29.055 176.220 29.345 176.265 ;
        RECT 23.980 176.080 29.345 176.220 ;
        RECT 23.980 176.020 24.300 176.080 ;
        RECT 26.740 176.020 27.060 176.080 ;
        RECT 29.055 176.035 29.345 176.080 ;
        RECT 39.635 176.220 39.925 176.265 ;
        RECT 41.920 176.220 42.240 176.280 ;
        RECT 39.635 176.080 42.240 176.220 ;
        RECT 39.635 176.035 39.925 176.080 ;
        RECT 41.920 176.020 42.240 176.080 ;
        RECT 49.740 176.020 50.060 176.280 ;
        RECT 78.735 176.220 79.025 176.265 ;
        RECT 80.100 176.220 80.420 176.280 ;
        RECT 78.735 176.080 80.420 176.220 ;
        RECT 78.735 176.035 79.025 176.080 ;
        RECT 80.100 176.020 80.420 176.080 ;
        RECT 92.995 176.220 93.285 176.265 ;
        RECT 93.440 176.220 93.760 176.280 ;
        RECT 95.280 176.220 95.600 176.280 ;
        RECT 92.995 176.080 95.600 176.220 ;
        RECT 92.995 176.035 93.285 176.080 ;
        RECT 93.440 176.020 93.760 176.080 ;
        RECT 95.280 176.020 95.600 176.080 ;
        RECT 104.940 176.220 105.260 176.280 ;
        RECT 111.840 176.220 112.160 176.280 ;
        RECT 117.360 176.220 117.680 176.280 ;
        RECT 104.940 176.080 111.610 176.220 ;
        RECT 104.940 176.020 105.260 176.080 ;
        RECT 30.895 175.695 31.185 175.925 ;
        RECT 49.280 175.880 49.600 175.940 ;
        RECT 50.200 175.880 50.520 175.940 ;
        RECT 48.450 175.740 50.520 175.880 ;
        RECT 25.820 175.540 26.140 175.600 ;
        RECT 21.770 175.400 26.140 175.540 ;
        RECT 21.770 175.260 21.910 175.400 ;
        RECT 25.820 175.340 26.140 175.400 ;
        RECT 28.120 175.540 28.440 175.600 ;
        RECT 29.515 175.540 29.805 175.585 ;
        RECT 28.120 175.400 29.805 175.540 ;
        RECT 30.970 175.540 31.110 175.695 ;
        RECT 30.970 175.400 34.790 175.540 ;
        RECT 28.120 175.340 28.440 175.400 ;
        RECT 29.515 175.355 29.805 175.400 ;
        RECT 21.235 175.200 21.525 175.245 ;
        RECT 21.680 175.200 22.000 175.260 ;
        RECT 21.235 175.060 22.000 175.200 ;
        RECT 21.235 175.015 21.525 175.060 ;
        RECT 21.680 175.000 22.000 175.060 ;
        RECT 22.615 175.200 22.905 175.245 ;
        RECT 23.980 175.200 24.300 175.260 ;
        RECT 22.615 175.060 24.300 175.200 ;
        RECT 22.615 175.015 22.905 175.060 ;
        RECT 23.980 175.000 24.300 175.060 ;
        RECT 27.200 175.200 27.520 175.260 ;
        RECT 29.055 175.200 29.345 175.245 ;
        RECT 27.200 175.060 29.345 175.200 ;
        RECT 27.200 175.000 27.520 175.060 ;
        RECT 29.055 175.015 29.345 175.060 ;
        RECT 30.880 175.200 31.200 175.260 ;
        RECT 32.275 175.200 32.565 175.245 ;
        RECT 30.880 175.060 32.565 175.200 ;
        RECT 30.880 175.000 31.200 175.060 ;
        RECT 32.275 175.015 32.565 175.060 ;
        RECT 33.180 175.000 33.500 175.260 ;
        RECT 33.640 175.000 33.960 175.260 ;
        RECT 34.650 175.245 34.790 175.400 ;
        RECT 36.030 175.400 40.310 175.540 ;
        RECT 36.030 175.260 36.170 175.400 ;
        RECT 34.575 175.015 34.865 175.245 ;
        RECT 35.035 175.015 35.325 175.245 ;
        RECT 35.495 175.200 35.785 175.245 ;
        RECT 35.940 175.200 36.260 175.260 ;
        RECT 35.495 175.060 36.260 175.200 ;
        RECT 35.495 175.015 35.785 175.060 ;
        RECT 35.110 174.860 35.250 175.015 ;
        RECT 35.940 175.000 36.260 175.060 ;
        RECT 36.400 175.200 36.720 175.260 ;
        RECT 40.170 175.245 40.310 175.400 ;
        RECT 46.520 175.340 46.840 175.600 ;
        RECT 48.450 175.585 48.590 175.740 ;
        RECT 49.280 175.680 49.600 175.740 ;
        RECT 50.200 175.680 50.520 175.740 ;
        RECT 81.480 175.880 81.770 175.925 ;
        RECT 83.050 175.880 83.340 175.925 ;
        RECT 85.150 175.880 85.440 175.925 ;
        RECT 81.480 175.740 85.440 175.880 ;
        RECT 81.480 175.695 81.770 175.740 ;
        RECT 83.050 175.695 83.340 175.740 ;
        RECT 85.150 175.695 85.440 175.740 ;
        RECT 86.580 175.880 86.870 175.925 ;
        RECT 88.680 175.880 88.970 175.925 ;
        RECT 90.250 175.880 90.540 175.925 ;
        RECT 86.580 175.740 90.540 175.880 ;
        RECT 86.580 175.695 86.870 175.740 ;
        RECT 88.680 175.695 88.970 175.740 ;
        RECT 90.250 175.695 90.540 175.740 ;
        RECT 98.040 175.880 98.330 175.925 ;
        RECT 99.610 175.880 99.900 175.925 ;
        RECT 101.710 175.880 102.000 175.925 ;
        RECT 98.040 175.740 102.000 175.880 ;
        RECT 98.040 175.695 98.330 175.740 ;
        RECT 99.610 175.695 99.900 175.740 ;
        RECT 101.710 175.695 102.000 175.740 ;
        RECT 104.480 175.880 104.800 175.940 ;
        RECT 109.095 175.880 109.385 175.925 ;
        RECT 104.480 175.740 109.385 175.880 ;
        RECT 104.480 175.680 104.800 175.740 ;
        RECT 109.095 175.695 109.385 175.740 ;
        RECT 48.375 175.355 48.665 175.585 ;
        RECT 52.500 175.540 52.820 175.600 ;
        RECT 50.290 175.400 52.820 175.540 ;
        RECT 50.290 175.260 50.430 175.400 ;
        RECT 52.500 175.340 52.820 175.400 ;
        RECT 81.045 175.540 81.335 175.585 ;
        RECT 83.565 175.540 83.855 175.585 ;
        RECT 84.755 175.540 85.045 175.585 ;
        RECT 81.045 175.400 85.045 175.540 ;
        RECT 81.045 175.355 81.335 175.400 ;
        RECT 83.565 175.355 83.855 175.400 ;
        RECT 84.755 175.355 85.045 175.400 ;
        RECT 85.635 175.540 85.925 175.585 ;
        RECT 86.080 175.540 86.400 175.600 ;
        RECT 85.635 175.400 86.400 175.540 ;
        RECT 85.635 175.355 85.925 175.400 ;
        RECT 86.080 175.340 86.400 175.400 ;
        RECT 86.975 175.540 87.265 175.585 ;
        RECT 88.165 175.540 88.455 175.585 ;
        RECT 90.685 175.540 90.975 175.585 ;
        RECT 86.975 175.400 90.975 175.540 ;
        RECT 86.975 175.355 87.265 175.400 ;
        RECT 88.165 175.355 88.455 175.400 ;
        RECT 90.685 175.355 90.975 175.400 ;
        RECT 97.605 175.540 97.895 175.585 ;
        RECT 100.125 175.540 100.415 175.585 ;
        RECT 101.315 175.540 101.605 175.585 ;
        RECT 97.605 175.400 101.605 175.540 ;
        RECT 97.605 175.355 97.895 175.400 ;
        RECT 100.125 175.355 100.415 175.400 ;
        RECT 101.315 175.355 101.605 175.400 ;
        RECT 103.100 175.540 103.420 175.600 ;
        RECT 109.555 175.540 109.845 175.585 ;
        RECT 103.100 175.400 109.845 175.540 ;
        RECT 103.100 175.340 103.420 175.400 ;
        RECT 109.555 175.355 109.845 175.400 ;
        RECT 110.935 175.355 111.225 175.585 ;
        RECT 38.255 175.200 38.545 175.245 ;
        RECT 36.400 175.060 38.545 175.200 ;
        RECT 36.400 175.000 36.720 175.060 ;
        RECT 38.255 175.015 38.545 175.060 ;
        RECT 40.095 175.200 40.385 175.245 ;
        RECT 41.475 175.200 41.765 175.245 ;
        RECT 40.095 175.060 41.765 175.200 ;
        RECT 40.095 175.015 40.385 175.060 ;
        RECT 41.475 175.015 41.765 175.060 ;
        RECT 50.200 175.000 50.520 175.260 ;
        RECT 51.120 175.000 51.440 175.260 ;
        RECT 52.960 175.000 53.280 175.260 ;
        RECT 60.320 175.200 60.640 175.260 ;
        RECT 63.080 175.200 63.400 175.260 ;
        RECT 60.320 175.060 63.400 175.200 ;
        RECT 60.320 175.000 60.640 175.060 ;
        RECT 63.080 175.000 63.400 175.060 ;
        RECT 64.475 175.200 64.765 175.245 ;
        RECT 65.380 175.200 65.700 175.260 ;
        RECT 66.315 175.200 66.605 175.245 ;
        RECT 68.140 175.200 68.460 175.260 ;
        RECT 72.280 175.200 72.600 175.260 ;
        RECT 64.475 175.060 72.600 175.200 ;
        RECT 64.475 175.015 64.765 175.060 ;
        RECT 65.380 175.000 65.700 175.060 ;
        RECT 66.315 175.015 66.605 175.060 ;
        RECT 68.140 175.000 68.460 175.060 ;
        RECT 72.280 175.000 72.600 175.060 ;
        RECT 76.435 175.015 76.725 175.245 ;
        RECT 77.355 175.200 77.645 175.245 ;
        RECT 78.260 175.200 78.580 175.260 ;
        RECT 77.355 175.060 78.580 175.200 ;
        RECT 77.355 175.015 77.645 175.060 ;
        RECT 40.555 174.860 40.845 174.905 ;
        RECT 41.920 174.860 42.240 174.920 ;
        RECT 35.110 174.720 42.240 174.860 ;
        RECT 40.555 174.675 40.845 174.720 ;
        RECT 41.920 174.660 42.240 174.720 ;
        RECT 48.960 174.860 49.250 174.905 ;
        RECT 50.675 174.860 50.965 174.905 ;
        RECT 48.960 174.720 50.965 174.860 ;
        RECT 48.960 174.675 49.250 174.720 ;
        RECT 50.675 174.675 50.965 174.720 ;
        RECT 64.920 174.860 65.240 174.920 ;
        RECT 67.220 174.860 67.540 174.920 ;
        RECT 76.510 174.860 76.650 175.015 ;
        RECT 78.260 175.000 78.580 175.060 ;
        RECT 87.430 175.200 87.720 175.245 ;
        RECT 91.140 175.200 91.460 175.260 ;
        RECT 87.430 175.060 91.460 175.200 ;
        RECT 87.430 175.015 87.720 175.060 ;
        RECT 91.140 175.000 91.460 175.060 ;
        RECT 98.040 175.200 98.360 175.260 ;
        RECT 102.195 175.200 102.485 175.245 ;
        RECT 98.040 175.060 102.485 175.200 ;
        RECT 98.040 175.000 98.360 175.060 ;
        RECT 102.195 175.015 102.485 175.060 ;
        RECT 104.020 175.000 104.340 175.260 ;
        RECT 107.240 175.200 107.560 175.260 ;
        RECT 108.635 175.200 108.925 175.245 ;
        RECT 107.240 175.060 108.925 175.200 ;
        RECT 107.240 175.000 107.560 175.060 ;
        RECT 108.635 175.015 108.925 175.060 ;
        RECT 110.015 175.200 110.305 175.245 ;
        RECT 111.010 175.200 111.150 175.355 ;
        RECT 110.015 175.060 111.150 175.200 ;
        RECT 111.470 175.200 111.610 176.080 ;
        RECT 111.840 176.080 117.680 176.220 ;
        RECT 111.840 176.020 112.160 176.080 ;
        RECT 117.360 176.020 117.680 176.080 ;
        RECT 118.740 176.020 119.060 176.280 ;
        RECT 112.760 175.880 113.080 175.940 ;
        RECT 111.930 175.740 113.080 175.880 ;
        RECT 111.930 175.585 112.070 175.740 ;
        RECT 112.760 175.680 113.080 175.740 ;
        RECT 114.600 175.880 114.920 175.940 ;
        RECT 118.295 175.880 118.585 175.925 ;
        RECT 124.260 175.880 124.580 175.940 ;
        RECT 114.600 175.740 116.670 175.880 ;
        RECT 114.600 175.680 114.920 175.740 ;
        RECT 111.855 175.355 112.145 175.585 ;
        RECT 112.315 175.540 112.605 175.585 ;
        RECT 113.680 175.540 114.000 175.600 ;
        RECT 112.315 175.400 114.000 175.540 ;
        RECT 112.315 175.355 112.605 175.400 ;
        RECT 113.680 175.340 114.000 175.400 ;
        RECT 112.760 175.200 113.080 175.260 ;
        RECT 111.470 175.060 113.080 175.200 ;
        RECT 110.015 175.015 110.305 175.060 ;
        RECT 112.760 175.000 113.080 175.060 ;
        RECT 113.235 175.200 113.525 175.245 ;
        RECT 114.600 175.200 114.920 175.260 ;
        RECT 115.980 175.200 116.300 175.260 ;
        RECT 116.530 175.245 116.670 175.740 ;
        RECT 118.295 175.740 124.580 175.880 ;
        RECT 118.295 175.695 118.585 175.740 ;
        RECT 124.260 175.680 124.580 175.740 ;
        RECT 120.120 175.540 120.440 175.600 ;
        RECT 132.555 175.540 132.845 175.585 ;
        RECT 120.120 175.400 132.845 175.540 ;
        RECT 120.120 175.340 120.440 175.400 ;
        RECT 132.555 175.355 132.845 175.400 ;
        RECT 113.235 175.060 113.910 175.200 ;
        RECT 113.235 175.015 113.525 175.060 ;
        RECT 64.920 174.720 76.650 174.860 ;
        RECT 81.940 174.860 82.260 174.920 ;
        RECT 84.300 174.860 84.590 174.905 ;
        RECT 81.940 174.720 84.590 174.860 ;
        RECT 64.920 174.660 65.240 174.720 ;
        RECT 67.220 174.660 67.540 174.720 ;
        RECT 81.940 174.660 82.260 174.720 ;
        RECT 84.300 174.675 84.590 174.720 ;
        RECT 100.970 174.860 101.260 174.905 ;
        RECT 107.715 174.860 108.005 174.905 ;
        RECT 100.970 174.720 108.005 174.860 ;
        RECT 100.970 174.675 101.260 174.720 ;
        RECT 107.715 174.675 108.005 174.720 ;
        RECT 18.920 174.520 19.240 174.580 ;
        RECT 21.695 174.520 21.985 174.565 ;
        RECT 18.920 174.380 21.985 174.520 ;
        RECT 18.920 174.320 19.240 174.380 ;
        RECT 21.695 174.335 21.985 174.380 ;
        RECT 33.195 174.520 33.485 174.565 ;
        RECT 35.940 174.520 36.260 174.580 ;
        RECT 33.195 174.380 36.260 174.520 ;
        RECT 33.195 174.335 33.485 174.380 ;
        RECT 35.940 174.320 36.260 174.380 ;
        RECT 36.860 174.320 37.180 174.580 ;
        RECT 37.320 174.320 37.640 174.580 ;
        RECT 42.380 174.320 42.700 174.580 ;
        RECT 47.915 174.520 48.205 174.565 ;
        RECT 51.120 174.520 51.440 174.580 ;
        RECT 47.915 174.380 51.440 174.520 ;
        RECT 47.915 174.335 48.205 174.380 ;
        RECT 51.120 174.320 51.440 174.380 ;
        RECT 76.880 174.320 77.200 174.580 ;
        RECT 95.295 174.520 95.585 174.565 ;
        RECT 99.420 174.520 99.740 174.580 ;
        RECT 104.020 174.520 104.340 174.580 ;
        RECT 95.295 174.380 104.340 174.520 ;
        RECT 95.295 174.335 95.585 174.380 ;
        RECT 99.420 174.320 99.740 174.380 ;
        RECT 104.020 174.320 104.340 174.380 ;
        RECT 107.255 174.520 107.545 174.565 ;
        RECT 113.770 174.520 113.910 175.060 ;
        RECT 114.600 175.060 116.300 175.200 ;
        RECT 114.600 175.000 114.920 175.060 ;
        RECT 115.980 175.000 116.300 175.060 ;
        RECT 116.455 175.015 116.745 175.245 ;
        RECT 117.375 175.200 117.665 175.245 ;
        RECT 118.280 175.200 118.600 175.260 ;
        RECT 119.200 175.200 119.520 175.260 ;
        RECT 117.375 175.060 119.520 175.200 ;
        RECT 117.375 175.015 117.665 175.060 ;
        RECT 118.280 175.000 118.600 175.060 ;
        RECT 119.200 175.000 119.520 175.060 ;
        RECT 120.580 175.000 120.900 175.260 ;
        RECT 127.480 175.000 127.800 175.260 ;
        RECT 134.380 175.200 134.700 175.260 ;
        RECT 136.695 175.200 136.985 175.245 ;
        RECT 134.380 175.060 136.985 175.200 ;
        RECT 134.380 175.000 134.700 175.060 ;
        RECT 136.695 175.015 136.985 175.060 ;
        RECT 119.660 174.660 119.980 174.920 ;
        RECT 131.635 174.860 131.925 174.905 ;
        RECT 133.935 174.860 134.225 174.905 ;
        RECT 131.635 174.720 134.225 174.860 ;
        RECT 131.635 174.675 131.925 174.720 ;
        RECT 133.935 174.675 134.225 174.720 ;
        RECT 107.255 174.380 113.910 174.520 ;
        RECT 114.140 174.520 114.460 174.580 ;
        RECT 116.900 174.520 117.220 174.580 ;
        RECT 114.140 174.380 117.220 174.520 ;
        RECT 107.255 174.335 107.545 174.380 ;
        RECT 114.140 174.320 114.460 174.380 ;
        RECT 116.900 174.320 117.220 174.380 ;
        RECT 125.640 174.520 125.960 174.580 ;
        RECT 127.020 174.520 127.340 174.580 ;
        RECT 125.640 174.380 127.340 174.520 ;
        RECT 125.640 174.320 125.960 174.380 ;
        RECT 127.020 174.320 127.340 174.380 ;
        RECT 128.400 174.320 128.720 174.580 ;
        RECT 129.780 174.320 130.100 174.580 ;
        RECT 130.240 174.520 130.560 174.580 ;
        RECT 132.095 174.520 132.385 174.565 ;
        RECT 130.240 174.380 132.385 174.520 ;
        RECT 130.240 174.320 130.560 174.380 ;
        RECT 132.095 174.335 132.385 174.380 ;
        RECT 13.330 173.700 138.910 174.180 ;
        RECT 69.980 173.500 70.300 173.560 ;
        RECT 72.295 173.500 72.585 173.545 ;
        RECT 69.980 173.360 72.585 173.500 ;
        RECT 69.980 173.300 70.300 173.360 ;
        RECT 72.295 173.315 72.585 173.360 ;
        RECT 77.340 173.300 77.660 173.560 ;
        RECT 79.655 173.500 79.945 173.545 ;
        RECT 80.100 173.500 80.420 173.560 ;
        RECT 79.655 173.360 80.420 173.500 ;
        RECT 79.655 173.315 79.945 173.360 ;
        RECT 80.100 173.300 80.420 173.360 ;
        RECT 81.940 173.300 82.260 173.560 ;
        RECT 103.100 173.300 103.420 173.560 ;
        RECT 112.760 173.500 113.080 173.560 ;
        RECT 114.025 173.500 114.315 173.545 ;
        RECT 118.740 173.500 119.060 173.560 ;
        RECT 112.760 173.360 114.315 173.500 ;
        RECT 112.760 173.300 113.080 173.360 ;
        RECT 114.025 173.315 114.315 173.360 ;
        RECT 115.150 173.360 119.060 173.500 ;
        RECT 19.380 173.160 19.700 173.220 ;
        RECT 23.520 173.160 23.840 173.220 ;
        RECT 36.860 173.160 37.180 173.220 ;
        RECT 46.980 173.160 47.300 173.220 ;
        RECT 48.820 173.160 49.140 173.220 ;
        RECT 52.975 173.160 53.265 173.205 ;
        RECT 19.380 173.020 21.450 173.160 ;
        RECT 19.380 172.960 19.700 173.020 ;
        RECT 18.920 172.620 19.240 172.880 ;
        RECT 21.310 172.865 21.450 173.020 ;
        RECT 21.770 173.020 23.840 173.160 ;
        RECT 21.235 172.820 21.525 172.865 ;
        RECT 21.770 172.820 21.910 173.020 ;
        RECT 23.520 172.960 23.840 173.020 ;
        RECT 24.070 173.020 36.170 173.160 ;
        RECT 21.235 172.680 21.910 172.820 ;
        RECT 22.155 172.820 22.445 172.865 ;
        RECT 24.070 172.820 24.210 173.020 ;
        RECT 22.155 172.680 24.210 172.820 ;
        RECT 21.235 172.635 21.525 172.680 ;
        RECT 22.155 172.635 22.445 172.680 ;
        RECT 26.740 172.620 27.060 172.880 ;
        RECT 28.120 172.820 28.440 172.880 ;
        RECT 29.975 172.820 30.265 172.865 ;
        RECT 28.120 172.680 30.265 172.820 ;
        RECT 28.120 172.620 28.440 172.680 ;
        RECT 29.975 172.635 30.265 172.680 ;
        RECT 31.340 172.820 31.660 172.880 ;
        RECT 35.495 172.820 35.785 172.865 ;
        RECT 31.340 172.680 35.785 172.820 ;
        RECT 31.340 172.620 31.660 172.680 ;
        RECT 35.495 172.635 35.785 172.680 ;
        RECT 19.395 172.480 19.685 172.525 ;
        RECT 21.680 172.480 22.000 172.540 ;
        RECT 19.395 172.340 22.000 172.480 ;
        RECT 19.395 172.295 19.685 172.340 ;
        RECT 21.680 172.280 22.000 172.340 ;
        RECT 27.200 172.280 27.520 172.540 ;
        RECT 30.435 172.480 30.725 172.525 ;
        RECT 30.880 172.480 31.200 172.540 ;
        RECT 30.435 172.340 31.200 172.480 ;
        RECT 30.435 172.295 30.725 172.340 ;
        RECT 30.880 172.280 31.200 172.340 ;
        RECT 28.595 172.140 28.885 172.185 ;
        RECT 31.430 172.140 31.570 172.620 ;
        RECT 28.595 172.000 31.570 172.140 ;
        RECT 36.030 172.140 36.170 173.020 ;
        RECT 36.860 173.020 40.310 173.160 ;
        RECT 36.860 172.960 37.180 173.020 ;
        RECT 36.415 172.820 36.705 172.865 ;
        RECT 37.320 172.820 37.640 172.880 ;
        RECT 36.415 172.680 37.640 172.820 ;
        RECT 36.415 172.635 36.705 172.680 ;
        RECT 37.320 172.620 37.640 172.680 ;
        RECT 37.780 172.820 38.100 172.880 ;
        RECT 40.170 172.865 40.310 173.020 ;
        RECT 46.980 173.020 53.265 173.160 ;
        RECT 46.980 172.960 47.300 173.020 ;
        RECT 48.820 172.960 49.140 173.020 ;
        RECT 52.975 172.975 53.265 173.020 ;
        RECT 62.635 173.160 62.925 173.205 ;
        RECT 66.620 173.160 66.910 173.205 ;
        RECT 104.940 173.160 105.260 173.220 ;
        RECT 115.150 173.205 115.290 173.360 ;
        RECT 118.740 173.300 119.060 173.360 ;
        RECT 120.120 173.300 120.440 173.560 ;
        RECT 126.575 173.500 126.865 173.545 ;
        RECT 127.480 173.500 127.800 173.560 ;
        RECT 133.935 173.500 134.225 173.545 ;
        RECT 134.380 173.500 134.700 173.560 ;
        RECT 126.575 173.360 127.800 173.500 ;
        RECT 126.575 173.315 126.865 173.360 ;
        RECT 127.480 173.300 127.800 173.360 ;
        RECT 128.030 173.360 134.700 173.500 ;
        RECT 62.635 173.020 66.910 173.160 ;
        RECT 62.635 172.975 62.925 173.020 ;
        RECT 66.620 172.975 66.910 173.020 ;
        RECT 102.270 173.020 105.260 173.160 ;
        RECT 39.635 172.820 39.925 172.865 ;
        RECT 37.780 172.680 39.925 172.820 ;
        RECT 37.780 172.620 38.100 172.680 ;
        RECT 39.635 172.635 39.925 172.680 ;
        RECT 40.100 172.635 40.390 172.865 ;
        RECT 40.540 172.820 40.860 172.880 ;
        RECT 42.380 172.865 42.700 172.880 ;
        RECT 41.015 172.820 41.305 172.865 ;
        RECT 40.540 172.680 41.305 172.820 ;
        RECT 40.540 172.620 40.860 172.680 ;
        RECT 41.015 172.635 41.305 172.680 ;
        RECT 41.475 172.635 41.765 172.865 ;
        RECT 42.165 172.635 42.700 172.865 ;
        RECT 37.410 172.480 37.550 172.620 ;
        RECT 41.550 172.480 41.690 172.635 ;
        RECT 42.380 172.620 42.700 172.635 ;
        RECT 49.740 172.620 50.060 172.880 ;
        RECT 61.255 172.820 61.545 172.865 ;
        RECT 64.920 172.820 65.240 172.880 ;
        RECT 61.255 172.680 65.240 172.820 ;
        RECT 61.255 172.635 61.545 172.680 ;
        RECT 64.920 172.620 65.240 172.680 ;
        RECT 65.380 172.620 65.700 172.880 ;
        RECT 78.260 172.820 78.580 172.880 ;
        RECT 80.115 172.820 80.405 172.865 ;
        RECT 78.260 172.680 80.405 172.820 ;
        RECT 78.260 172.620 78.580 172.680 ;
        RECT 80.115 172.635 80.405 172.680 ;
        RECT 83.795 172.820 84.085 172.865 ;
        RECT 91.140 172.820 91.460 172.880 ;
        RECT 83.795 172.680 91.460 172.820 ;
        RECT 83.795 172.635 84.085 172.680 ;
        RECT 91.140 172.620 91.460 172.680 ;
        RECT 93.900 172.620 94.220 172.880 ;
        RECT 102.270 172.865 102.410 173.020 ;
        RECT 104.940 172.960 105.260 173.020 ;
        RECT 115.075 172.975 115.365 173.205 ;
        RECT 115.980 173.160 116.300 173.220 ;
        RECT 128.030 173.160 128.170 173.360 ;
        RECT 133.935 173.315 134.225 173.360 ;
        RECT 134.380 173.300 134.700 173.360 ;
        RECT 136.680 173.300 137.000 173.560 ;
        RECT 115.980 173.020 118.510 173.160 ;
        RECT 115.980 172.960 116.300 173.020 ;
        RECT 102.195 172.635 102.485 172.865 ;
        RECT 103.115 172.820 103.405 172.865 ;
        RECT 104.020 172.820 104.340 172.880 ;
        RECT 103.115 172.680 104.340 172.820 ;
        RECT 103.115 172.635 103.405 172.680 ;
        RECT 104.020 172.620 104.340 172.680 ;
        RECT 116.915 172.820 117.205 172.865 ;
        RECT 117.360 172.820 117.680 172.880 ;
        RECT 118.370 172.865 118.510 173.020 ;
        RECT 125.730 173.020 128.170 173.160 ;
        RECT 128.370 173.160 128.660 173.205 ;
        RECT 129.780 173.160 130.100 173.220 ;
        RECT 128.370 173.020 130.100 173.160 ;
        RECT 125.730 172.865 125.870 173.020 ;
        RECT 128.370 172.975 128.660 173.020 ;
        RECT 129.780 172.960 130.100 173.020 ;
        RECT 132.080 173.160 132.400 173.220 ;
        RECT 132.080 173.020 135.990 173.160 ;
        RECT 132.080 172.960 132.400 173.020 ;
        RECT 116.915 172.680 117.680 172.820 ;
        RECT 116.915 172.635 117.205 172.680 ;
        RECT 117.360 172.620 117.680 172.680 ;
        RECT 117.835 172.635 118.125 172.865 ;
        RECT 118.295 172.635 118.585 172.865 ;
        RECT 118.755 172.635 119.045 172.865 ;
        RECT 125.655 172.635 125.945 172.865 ;
        RECT 126.560 172.820 126.880 172.880 ;
        RECT 127.035 172.820 127.325 172.865 ;
        RECT 126.560 172.680 127.325 172.820 ;
        RECT 37.410 172.340 41.690 172.480 ;
        RECT 50.200 172.280 50.520 172.540 ;
        RECT 51.120 172.480 51.440 172.540 ;
        RECT 52.055 172.480 52.345 172.525 ;
        RECT 51.120 172.340 52.345 172.480 ;
        RECT 51.120 172.280 51.440 172.340 ;
        RECT 52.055 172.295 52.345 172.340 ;
        RECT 62.635 172.295 62.925 172.525 ;
        RECT 66.275 172.480 66.565 172.525 ;
        RECT 67.465 172.480 67.755 172.525 ;
        RECT 69.985 172.480 70.275 172.525 ;
        RECT 66.275 172.340 70.275 172.480 ;
        RECT 66.275 172.295 66.565 172.340 ;
        RECT 67.465 172.295 67.755 172.340 ;
        RECT 69.985 172.295 70.275 172.340 ;
        RECT 45.140 172.140 45.460 172.200 ;
        RECT 47.440 172.140 47.760 172.200 ;
        RECT 48.360 172.140 48.680 172.200 ;
        RECT 59.860 172.140 60.180 172.200 ;
        RECT 36.030 172.000 60.180 172.140 ;
        RECT 28.595 171.955 28.885 172.000 ;
        RECT 45.140 171.940 45.460 172.000 ;
        RECT 47.440 171.940 47.760 172.000 ;
        RECT 48.360 171.940 48.680 172.000 ;
        RECT 59.860 171.940 60.180 172.000 ;
        RECT 20.760 171.600 21.080 171.860 ;
        RECT 31.355 171.800 31.645 171.845 ;
        RECT 31.800 171.800 32.120 171.860 ;
        RECT 35.495 171.800 35.785 171.845 ;
        RECT 31.355 171.660 35.785 171.800 ;
        RECT 31.355 171.615 31.645 171.660 ;
        RECT 31.800 171.600 32.120 171.660 ;
        RECT 35.495 171.615 35.785 171.660 ;
        RECT 37.335 171.800 37.625 171.845 ;
        RECT 37.780 171.800 38.100 171.860 ;
        RECT 37.335 171.660 38.100 171.800 ;
        RECT 37.335 171.615 37.625 171.660 ;
        RECT 37.780 171.600 38.100 171.660 ;
        RECT 42.840 171.600 43.160 171.860 ;
        RECT 51.595 171.800 51.885 171.845 ;
        RECT 59.400 171.800 59.720 171.860 ;
        RECT 51.595 171.660 59.720 171.800 ;
        RECT 51.595 171.615 51.885 171.660 ;
        RECT 59.400 171.600 59.720 171.660 ;
        RECT 61.700 171.600 62.020 171.860 ;
        RECT 62.710 171.800 62.850 172.295 ;
        RECT 74.120 172.280 74.440 172.540 ;
        RECT 75.960 172.480 76.280 172.540 ;
        RECT 80.575 172.480 80.865 172.525 ;
        RECT 75.960 172.340 80.865 172.480 ;
        RECT 75.960 172.280 76.280 172.340 ;
        RECT 80.575 172.295 80.865 172.340 ;
        RECT 84.240 172.280 84.560 172.540 ;
        RECT 85.160 172.280 85.480 172.540 ;
        RECT 86.080 172.480 86.400 172.540 ;
        RECT 97.595 172.480 97.885 172.525 ;
        RECT 98.040 172.480 98.360 172.540 ;
        RECT 86.080 172.340 98.360 172.480 ;
        RECT 117.910 172.480 118.050 172.635 ;
        RECT 117.910 172.340 118.280 172.480 ;
        RECT 86.080 172.280 86.400 172.340 ;
        RECT 97.595 172.295 97.885 172.340 ;
        RECT 98.040 172.280 98.360 172.340 ;
        RECT 118.140 172.200 118.280 172.340 ;
        RECT 65.880 172.140 66.170 172.185 ;
        RECT 67.980 172.140 68.270 172.185 ;
        RECT 69.550 172.140 69.840 172.185 ;
        RECT 76.880 172.140 77.200 172.200 ;
        RECT 65.880 172.000 69.840 172.140 ;
        RECT 65.880 171.955 66.170 172.000 ;
        RECT 67.980 171.955 68.270 172.000 ;
        RECT 69.550 171.955 69.840 172.000 ;
        RECT 71.910 172.000 77.200 172.140 ;
        RECT 118.140 172.000 118.600 172.200 ;
        RECT 71.910 171.800 72.050 172.000 ;
        RECT 76.880 171.940 77.200 172.000 ;
        RECT 118.280 171.940 118.600 172.000 ;
        RECT 62.710 171.660 72.050 171.800 ;
        RECT 77.800 171.600 78.120 171.860 ;
        RECT 113.220 171.600 113.540 171.860 ;
        RECT 113.680 171.800 114.000 171.860 ;
        RECT 114.155 171.800 114.445 171.845 ;
        RECT 113.680 171.660 114.445 171.800 ;
        RECT 113.680 171.600 114.000 171.660 ;
        RECT 114.155 171.615 114.445 171.660 ;
        RECT 115.520 171.800 115.840 171.860 ;
        RECT 117.820 171.800 118.140 171.860 ;
        RECT 118.830 171.800 118.970 172.635 ;
        RECT 126.560 172.620 126.880 172.680 ;
        RECT 127.035 172.635 127.325 172.680 ;
        RECT 135.300 172.620 135.620 172.880 ;
        RECT 135.850 172.865 135.990 173.020 ;
        RECT 135.775 172.635 136.065 172.865 ;
        RECT 127.915 172.480 128.205 172.525 ;
        RECT 129.105 172.480 129.395 172.525 ;
        RECT 131.625 172.480 131.915 172.525 ;
        RECT 127.915 172.340 131.915 172.480 ;
        RECT 127.915 172.295 128.205 172.340 ;
        RECT 129.105 172.295 129.395 172.340 ;
        RECT 131.625 172.295 131.915 172.340 ;
        RECT 127.520 172.140 127.810 172.185 ;
        RECT 129.620 172.140 129.910 172.185 ;
        RECT 131.190 172.140 131.480 172.185 ;
        RECT 127.520 172.000 131.480 172.140 ;
        RECT 127.520 171.955 127.810 172.000 ;
        RECT 129.620 171.955 129.910 172.000 ;
        RECT 131.190 171.955 131.480 172.000 ;
        RECT 120.580 171.800 120.900 171.860 ;
        RECT 115.520 171.660 120.900 171.800 ;
        RECT 115.520 171.600 115.840 171.660 ;
        RECT 117.820 171.600 118.140 171.660 ;
        RECT 120.580 171.600 120.900 171.660 ;
        RECT 134.380 171.600 134.700 171.860 ;
        RECT 13.330 170.980 138.910 171.460 ;
        RECT 15.715 170.780 16.005 170.825 ;
        RECT 28.580 170.780 28.900 170.840 ;
        RECT 15.715 170.640 28.900 170.780 ;
        RECT 15.715 170.595 16.005 170.640 ;
        RECT 28.580 170.580 28.900 170.640 ;
        RECT 33.180 170.780 33.500 170.840 ;
        RECT 35.035 170.780 35.325 170.825 ;
        RECT 60.320 170.780 60.640 170.840 ;
        RECT 33.180 170.640 35.325 170.780 ;
        RECT 33.180 170.580 33.500 170.640 ;
        RECT 35.035 170.595 35.325 170.640 ;
        RECT 35.555 170.640 60.640 170.780 ;
        RECT 21.220 170.440 21.540 170.500 ;
        RECT 35.555 170.440 35.695 170.640 ;
        RECT 60.320 170.580 60.640 170.640 ;
        RECT 66.315 170.780 66.605 170.825 ;
        RECT 69.075 170.780 69.365 170.825 ;
        RECT 70.440 170.780 70.760 170.840 ;
        RECT 66.315 170.640 70.760 170.780 ;
        RECT 66.315 170.595 66.605 170.640 ;
        RECT 69.075 170.595 69.365 170.640 ;
        RECT 70.440 170.580 70.760 170.640 ;
        RECT 76.880 170.580 77.200 170.840 ;
        RECT 91.140 170.580 91.460 170.840 ;
        RECT 115.535 170.780 115.825 170.825 ;
        RECT 120.120 170.780 120.440 170.840 ;
        RECT 115.535 170.640 120.440 170.780 ;
        RECT 115.535 170.595 115.825 170.640 ;
        RECT 120.120 170.580 120.440 170.640 ;
        RECT 126.115 170.780 126.405 170.825 ;
        RECT 130.240 170.780 130.560 170.840 ;
        RECT 126.115 170.640 130.560 170.780 ;
        RECT 126.115 170.595 126.405 170.640 ;
        RECT 130.240 170.580 130.560 170.640 ;
        RECT 21.220 170.300 35.695 170.440 ;
        RECT 46.980 170.440 47.300 170.500 ;
        RECT 50.200 170.440 50.520 170.500 ;
        RECT 55.260 170.440 55.550 170.485 ;
        RECT 56.830 170.440 57.120 170.485 ;
        RECT 58.930 170.440 59.220 170.485 ;
        RECT 46.980 170.300 50.890 170.440 ;
        RECT 21.220 170.240 21.540 170.300 ;
        RECT 18.935 170.100 19.225 170.145 ;
        RECT 20.300 170.100 20.620 170.160 ;
        RECT 18.935 169.960 20.620 170.100 ;
        RECT 18.935 169.915 19.225 169.960 ;
        RECT 20.300 169.900 20.620 169.960 ;
        RECT 20.760 170.100 21.080 170.160 ;
        RECT 22.950 170.100 23.240 170.145 ;
        RECT 20.760 169.960 23.240 170.100 ;
        RECT 20.760 169.900 21.080 169.960 ;
        RECT 22.950 169.915 23.240 169.960 ;
        RECT 23.520 169.900 23.840 170.160 ;
        RECT 25.450 170.145 25.590 170.300 ;
        RECT 46.980 170.240 47.300 170.300 ;
        RECT 50.200 170.240 50.520 170.300 ;
        RECT 25.375 169.915 25.665 170.145 ;
        RECT 35.940 169.900 36.260 170.160 ;
        RECT 36.400 170.100 36.720 170.160 ;
        RECT 41.460 170.100 41.780 170.160 ;
        RECT 36.400 169.960 48.130 170.100 ;
        RECT 36.400 169.900 36.720 169.960 ;
        RECT 12.020 169.760 12.340 169.820 ;
        RECT 14.795 169.760 15.085 169.805 ;
        RECT 12.020 169.620 15.085 169.760 ;
        RECT 12.020 169.560 12.340 169.620 ;
        RECT 14.795 169.575 15.085 169.620 ;
        RECT 18.475 169.760 18.765 169.805 ;
        RECT 19.380 169.760 19.700 169.820 ;
        RECT 18.475 169.620 19.700 169.760 ;
        RECT 20.390 169.760 20.530 169.900 ;
        RECT 23.995 169.760 24.285 169.805 ;
        RECT 20.390 169.620 24.285 169.760 ;
        RECT 18.475 169.575 18.765 169.620 ;
        RECT 19.380 169.560 19.700 169.620 ;
        RECT 23.995 169.575 24.285 169.620 ;
        RECT 26.740 169.760 27.060 169.820 ;
        RECT 27.215 169.760 27.505 169.805 ;
        RECT 26.740 169.620 27.505 169.760 ;
        RECT 26.740 169.560 27.060 169.620 ;
        RECT 27.215 169.575 27.505 169.620 ;
        RECT 28.120 169.560 28.440 169.820 ;
        RECT 31.340 169.560 31.660 169.820 ;
        RECT 31.800 169.560 32.120 169.820 ;
        RECT 32.735 169.575 33.025 169.805 ;
        RECT 21.235 169.420 21.525 169.465 ;
        RECT 21.680 169.420 22.000 169.480 ;
        RECT 21.235 169.280 22.000 169.420 ;
        RECT 32.810 169.420 32.950 169.575 ;
        RECT 33.180 169.560 33.500 169.820 ;
        RECT 34.560 169.805 34.880 169.820 ;
        RECT 34.515 169.575 34.880 169.805 ;
        RECT 34.560 169.560 34.880 169.575 ;
        RECT 36.860 169.560 37.180 169.820 ;
        RECT 40.540 169.760 40.860 169.820 ;
        RECT 41.090 169.805 41.230 169.960 ;
        RECT 41.460 169.900 41.780 169.960 ;
        RECT 37.410 169.620 40.860 169.760 ;
        RECT 35.480 169.420 35.800 169.480 ;
        RECT 37.410 169.420 37.550 169.620 ;
        RECT 40.540 169.560 40.860 169.620 ;
        RECT 41.015 169.575 41.305 169.805 ;
        RECT 44.680 169.760 45.000 169.820 ;
        RECT 47.990 169.805 48.130 169.960 ;
        RECT 49.740 169.900 50.060 170.160 ;
        RECT 50.750 170.145 50.890 170.300 ;
        RECT 55.260 170.300 59.220 170.440 ;
        RECT 55.260 170.255 55.550 170.300 ;
        RECT 56.830 170.255 57.120 170.300 ;
        RECT 58.930 170.255 59.220 170.300 ;
        RECT 61.700 170.440 62.020 170.500 ;
        RECT 69.980 170.440 70.300 170.500 ;
        RECT 61.700 170.300 70.300 170.440 ;
        RECT 61.700 170.240 62.020 170.300 ;
        RECT 69.980 170.240 70.300 170.300 ;
        RECT 50.675 169.915 50.965 170.145 ;
        RECT 54.825 170.100 55.115 170.145 ;
        RECT 57.345 170.100 57.635 170.145 ;
        RECT 58.535 170.100 58.825 170.145 ;
        RECT 54.825 169.960 58.825 170.100 ;
        RECT 54.825 169.915 55.115 169.960 ;
        RECT 57.345 169.915 57.635 169.960 ;
        RECT 58.535 169.915 58.825 169.960 ;
        RECT 69.520 170.100 69.840 170.160 ;
        RECT 70.530 170.100 70.670 170.580 ;
        RECT 74.135 170.255 74.425 170.485 ;
        RECT 120.580 170.440 120.900 170.500 ;
        RECT 120.580 170.300 121.730 170.440 ;
        RECT 69.520 169.900 69.980 170.100 ;
        RECT 70.530 169.960 72.510 170.100 ;
        RECT 46.535 169.760 46.825 169.805 ;
        RECT 44.680 169.620 46.825 169.760 ;
        RECT 44.680 169.560 45.000 169.620 ;
        RECT 46.535 169.575 46.825 169.620 ;
        RECT 47.915 169.575 48.205 169.805 ;
        RECT 49.295 169.575 49.585 169.805 ;
        RECT 50.215 169.760 50.505 169.805 ;
        RECT 52.500 169.760 52.820 169.820 ;
        RECT 50.215 169.620 52.820 169.760 ;
        RECT 50.215 169.575 50.505 169.620 ;
        RECT 32.810 169.280 35.800 169.420 ;
        RECT 21.235 169.235 21.525 169.280 ;
        RECT 21.680 169.220 22.000 169.280 ;
        RECT 35.480 169.220 35.800 169.280 ;
        RECT 36.950 169.280 37.550 169.420 ;
        RECT 17.540 168.880 17.860 169.140 ;
        RECT 22.140 168.880 22.460 169.140 ;
        RECT 27.675 169.080 27.965 169.125 ;
        RECT 29.960 169.080 30.280 169.140 ;
        RECT 27.675 168.940 30.280 169.080 ;
        RECT 27.675 168.895 27.965 168.940 ;
        RECT 29.960 168.880 30.280 168.940 ;
        RECT 34.115 169.080 34.405 169.125 ;
        RECT 36.950 169.080 37.090 169.280 ;
        RECT 40.080 169.220 40.400 169.480 ;
        RECT 49.370 169.420 49.510 169.575 ;
        RECT 52.500 169.560 52.820 169.620 ;
        RECT 58.940 169.760 59.260 169.820 ;
        RECT 59.415 169.760 59.705 169.805 ;
        RECT 69.840 169.760 69.980 169.900 ;
        RECT 72.370 169.805 72.510 169.960 ;
        RECT 71.835 169.760 72.125 169.805 ;
        RECT 58.940 169.620 59.705 169.760 ;
        RECT 58.940 169.560 59.260 169.620 ;
        RECT 59.415 169.575 59.705 169.620 ;
        RECT 68.230 169.620 72.125 169.760 ;
        RECT 68.230 169.480 68.370 169.620 ;
        RECT 71.835 169.575 72.125 169.620 ;
        RECT 72.295 169.575 72.585 169.805 ;
        RECT 72.755 169.760 73.045 169.805 ;
        RECT 73.200 169.760 73.520 169.820 ;
        RECT 72.755 169.620 73.520 169.760 ;
        RECT 72.755 169.575 73.045 169.620 ;
        RECT 73.200 169.560 73.520 169.620 ;
        RECT 73.675 169.760 73.965 169.805 ;
        RECT 74.210 169.760 74.350 170.255 ;
        RECT 120.580 170.240 120.900 170.300 ;
        RECT 74.580 170.100 74.900 170.160 ;
        RECT 75.515 170.100 75.805 170.145 ;
        RECT 74.580 169.960 75.805 170.100 ;
        RECT 74.580 169.900 74.900 169.960 ;
        RECT 75.515 169.915 75.805 169.960 ;
        RECT 83.780 169.900 84.100 170.160 ;
        RECT 93.440 169.900 93.760 170.160 ;
        RECT 94.360 169.900 94.680 170.160 ;
        RECT 117.820 170.100 118.140 170.160 ;
        RECT 117.820 169.960 121.270 170.100 ;
        RECT 117.820 169.900 118.140 169.960 ;
        RECT 73.675 169.620 74.350 169.760 ;
        RECT 73.675 169.575 73.965 169.620 ;
        RECT 75.055 169.575 75.345 169.805 ;
        RECT 75.960 169.760 76.280 169.820 ;
        RECT 77.355 169.760 77.645 169.805 ;
        RECT 75.960 169.620 77.645 169.760 ;
        RECT 56.180 169.420 56.500 169.480 ;
        RECT 58.080 169.420 58.370 169.465 ;
        RECT 45.230 169.280 52.730 169.420 ;
        RECT 34.115 168.940 37.090 169.080 ;
        RECT 37.320 169.080 37.640 169.140 ;
        RECT 37.795 169.080 38.085 169.125 ;
        RECT 37.320 168.940 38.085 169.080 ;
        RECT 34.115 168.895 34.405 168.940 ;
        RECT 37.320 168.880 37.640 168.940 ;
        RECT 37.795 168.895 38.085 168.940 ;
        RECT 39.160 168.880 39.480 169.140 ;
        RECT 40.170 169.080 40.310 169.220 ;
        RECT 45.230 169.080 45.370 169.280 ;
        RECT 40.170 168.940 45.370 169.080 ;
        RECT 45.600 168.880 45.920 169.140 ;
        RECT 47.455 169.080 47.745 169.125 ;
        RECT 49.740 169.080 50.060 169.140 ;
        RECT 47.455 168.940 50.060 169.080 ;
        RECT 47.455 168.895 47.745 168.940 ;
        RECT 49.740 168.880 50.060 168.940 ;
        RECT 51.580 168.880 51.900 169.140 ;
        RECT 52.590 169.125 52.730 169.280 ;
        RECT 56.180 169.280 58.370 169.420 ;
        RECT 56.180 169.220 56.500 169.280 ;
        RECT 58.080 169.235 58.370 169.280 ;
        RECT 65.395 169.420 65.685 169.465 ;
        RECT 68.140 169.420 68.460 169.480 ;
        RECT 65.395 169.280 68.460 169.420 ;
        RECT 65.395 169.235 65.685 169.280 ;
        RECT 68.140 169.220 68.460 169.280 ;
        RECT 69.060 169.465 69.380 169.480 ;
        RECT 69.060 169.235 69.445 169.465 ;
        RECT 75.130 169.420 75.270 169.575 ;
        RECT 75.960 169.560 76.280 169.620 ;
        RECT 77.355 169.575 77.645 169.620 ;
        RECT 79.655 169.760 79.945 169.805 ;
        RECT 80.100 169.760 80.420 169.820 ;
        RECT 79.655 169.620 80.420 169.760 ;
        RECT 79.655 169.575 79.945 169.620 ;
        RECT 80.100 169.560 80.420 169.620 ;
        RECT 80.560 169.760 80.880 169.820 ;
        RECT 87.015 169.760 87.305 169.805 ;
        RECT 80.560 169.620 87.305 169.760 ;
        RECT 80.560 169.560 80.880 169.620 ;
        RECT 87.015 169.575 87.305 169.620 ;
        RECT 92.060 169.760 92.380 169.820 ;
        RECT 96.675 169.760 96.965 169.805 ;
        RECT 92.060 169.620 96.965 169.760 ;
        RECT 92.060 169.560 92.380 169.620 ;
        RECT 96.675 169.575 96.965 169.620 ;
        RECT 111.380 169.760 111.700 169.820 ;
        RECT 113.695 169.760 113.985 169.805 ;
        RECT 111.380 169.620 113.985 169.760 ;
        RECT 111.380 169.560 111.700 169.620 ;
        RECT 113.695 169.575 113.985 169.620 ;
        RECT 114.615 169.760 114.905 169.805 ;
        RECT 115.060 169.760 115.380 169.820 ;
        RECT 114.615 169.620 115.380 169.760 ;
        RECT 114.615 169.575 114.905 169.620 ;
        RECT 115.060 169.560 115.380 169.620 ;
        RECT 115.520 169.760 115.840 169.820 ;
        RECT 115.520 169.755 116.670 169.760 ;
        RECT 116.915 169.755 117.205 169.805 ;
        RECT 115.520 169.620 117.205 169.755 ;
        RECT 115.520 169.560 115.840 169.620 ;
        RECT 116.530 169.615 117.205 169.620 ;
        RECT 116.915 169.575 117.205 169.615 ;
        RECT 70.070 169.280 75.270 169.420 ;
        RECT 84.715 169.420 85.005 169.465 ;
        RECT 97.120 169.420 97.440 169.480 ;
        RECT 117.375 169.465 117.665 169.695 ;
        RECT 119.200 169.560 119.520 169.820 ;
        RECT 119.660 169.560 119.980 169.820 ;
        RECT 121.130 169.805 121.270 169.960 ;
        RECT 121.590 169.805 121.730 170.300 ;
        RECT 125.640 170.100 125.960 170.160 ;
        RECT 132.555 170.100 132.845 170.145 ;
        RECT 125.640 169.960 132.845 170.100 ;
        RECT 125.640 169.900 125.960 169.960 ;
        RECT 132.555 169.915 132.845 169.960 ;
        RECT 120.595 169.760 120.885 169.805 ;
        RECT 120.210 169.620 120.885 169.760 ;
        RECT 84.715 169.280 97.440 169.420 ;
        RECT 69.060 169.220 69.380 169.235 ;
        RECT 66.300 169.125 66.620 169.140 ;
        RECT 52.515 168.895 52.805 169.125 ;
        RECT 66.300 168.895 66.685 169.125 ;
        RECT 66.300 168.880 66.620 168.895 ;
        RECT 67.220 168.880 67.540 169.140 ;
        RECT 70.070 169.125 70.210 169.280 ;
        RECT 84.715 169.235 85.005 169.280 ;
        RECT 97.120 169.220 97.440 169.280 ;
        RECT 69.995 168.895 70.285 169.125 ;
        RECT 70.455 169.080 70.745 169.125 ;
        RECT 72.740 169.080 73.060 169.140 ;
        RECT 70.455 168.940 73.060 169.080 ;
        RECT 70.455 168.895 70.745 168.940 ;
        RECT 72.740 168.880 73.060 168.940 ;
        RECT 82.415 169.080 82.705 169.125 ;
        RECT 84.255 169.080 84.545 169.125 ;
        RECT 82.415 168.940 84.545 169.080 ;
        RECT 82.415 168.895 82.705 168.940 ;
        RECT 84.255 168.895 84.545 168.940 ;
        RECT 85.620 169.080 85.940 169.140 ;
        RECT 86.555 169.080 86.845 169.125 ;
        RECT 85.620 168.940 86.845 169.080 ;
        RECT 85.620 168.880 85.940 168.940 ;
        RECT 86.555 168.895 86.845 168.940 ;
        RECT 87.920 169.080 88.240 169.140 ;
        RECT 90.235 169.080 90.525 169.125 ;
        RECT 87.920 168.940 90.525 169.080 ;
        RECT 87.920 168.880 88.240 168.940 ;
        RECT 90.235 168.895 90.525 168.940 ;
        RECT 92.995 169.080 93.285 169.125 ;
        RECT 93.440 169.080 93.760 169.140 ;
        RECT 92.995 168.940 93.760 169.080 ;
        RECT 92.995 168.895 93.285 168.940 ;
        RECT 93.440 168.880 93.760 168.940 ;
        RECT 99.895 169.080 100.185 169.125 ;
        RECT 100.800 169.080 101.120 169.140 ;
        RECT 99.895 168.940 101.120 169.080 ;
        RECT 99.895 168.895 100.185 168.940 ;
        RECT 100.800 168.880 101.120 168.940 ;
        RECT 105.860 169.080 106.180 169.140 ;
        RECT 109.080 169.080 109.400 169.140 ;
        RECT 114.600 169.080 114.920 169.140 ;
        RECT 105.860 168.940 114.920 169.080 ;
        RECT 105.860 168.880 106.180 168.940 ;
        RECT 109.080 168.880 109.400 168.940 ;
        RECT 114.600 168.880 114.920 168.940 ;
        RECT 115.980 168.880 116.300 169.140 ;
        RECT 116.900 169.080 117.220 169.140 ;
        RECT 117.450 169.080 117.590 169.465 ;
        RECT 118.740 169.220 119.060 169.480 ;
        RECT 116.900 168.940 117.590 169.080 ;
        RECT 117.820 169.080 118.140 169.140 ;
        RECT 120.210 169.080 120.350 169.620 ;
        RECT 120.595 169.575 120.885 169.620 ;
        RECT 121.055 169.575 121.345 169.805 ;
        RECT 121.515 169.575 121.805 169.805 ;
        RECT 123.355 169.760 123.645 169.805 ;
        RECT 123.800 169.760 124.120 169.820 ;
        RECT 123.355 169.620 124.120 169.760 ;
        RECT 123.355 169.575 123.645 169.620 ;
        RECT 123.800 169.560 124.120 169.620 ;
        RECT 125.195 169.760 125.485 169.805 ;
        RECT 126.100 169.760 126.420 169.820 ;
        RECT 125.195 169.620 126.420 169.760 ;
        RECT 125.195 169.575 125.485 169.620 ;
        RECT 126.100 169.560 126.420 169.620 ;
        RECT 133.460 169.760 133.780 169.820 ;
        RECT 135.300 169.760 135.620 169.820 ;
        RECT 136.695 169.760 136.985 169.805 ;
        RECT 133.460 169.620 136.985 169.760 ;
        RECT 133.460 169.560 133.780 169.620 ;
        RECT 135.300 169.560 135.620 169.620 ;
        RECT 136.695 169.575 136.985 169.620 ;
        RECT 122.420 169.420 122.740 169.480 ;
        RECT 124.275 169.420 124.565 169.465 ;
        RECT 122.420 169.280 124.565 169.420 ;
        RECT 122.420 169.220 122.740 169.280 ;
        RECT 124.275 169.235 124.565 169.280 ;
        RECT 124.735 169.420 125.025 169.465 ;
        RECT 128.860 169.420 129.180 169.480 ;
        RECT 124.735 169.280 129.180 169.420 ;
        RECT 124.735 169.235 125.025 169.280 ;
        RECT 128.860 169.220 129.180 169.280 ;
        RECT 131.635 169.420 131.925 169.465 ;
        RECT 133.935 169.420 134.225 169.465 ;
        RECT 131.635 169.280 134.225 169.420 ;
        RECT 131.635 169.235 131.925 169.280 ;
        RECT 133.935 169.235 134.225 169.280 ;
        RECT 117.820 168.940 120.350 169.080 ;
        RECT 122.895 169.080 123.185 169.125 ;
        RECT 129.320 169.080 129.640 169.140 ;
        RECT 122.895 168.940 129.640 169.080 ;
        RECT 116.900 168.880 117.220 168.940 ;
        RECT 117.820 168.880 118.140 168.940 ;
        RECT 122.895 168.895 123.185 168.940 ;
        RECT 129.320 168.880 129.640 168.940 ;
        RECT 129.780 168.880 130.100 169.140 ;
        RECT 130.700 169.080 131.020 169.140 ;
        RECT 132.095 169.080 132.385 169.125 ;
        RECT 130.700 168.940 132.385 169.080 ;
        RECT 130.700 168.880 131.020 168.940 ;
        RECT 132.095 168.895 132.385 168.940 ;
        RECT 13.330 168.260 138.910 168.740 ;
        RECT 17.095 168.060 17.385 168.105 ;
        RECT 18.920 168.060 19.240 168.120 ;
        RECT 28.120 168.060 28.440 168.120 ;
        RECT 32.735 168.060 33.025 168.105 ;
        RECT 34.100 168.060 34.420 168.120 ;
        RECT 17.095 167.920 31.570 168.060 ;
        RECT 17.095 167.875 17.385 167.920 ;
        RECT 18.920 167.860 19.240 167.920 ;
        RECT 28.120 167.860 28.440 167.920 ;
        RECT 31.430 167.765 31.570 167.920 ;
        RECT 32.735 167.920 34.420 168.060 ;
        RECT 32.735 167.875 33.025 167.920 ;
        RECT 34.100 167.860 34.420 167.920 ;
        RECT 35.480 168.060 35.800 168.120 ;
        RECT 44.680 168.060 45.000 168.120 ;
        RECT 35.480 167.920 45.000 168.060 ;
        RECT 35.480 167.860 35.800 167.920 ;
        RECT 44.680 167.860 45.000 167.920 ;
        RECT 48.360 168.060 48.680 168.120 ;
        RECT 49.295 168.060 49.585 168.105 ;
        RECT 48.360 167.920 49.585 168.060 ;
        RECT 48.360 167.860 48.680 167.920 ;
        RECT 49.295 167.875 49.585 167.920 ;
        RECT 49.740 168.060 50.060 168.120 ;
        RECT 51.135 168.060 51.425 168.105 ;
        RECT 49.740 167.920 51.425 168.060 ;
        RECT 49.740 167.860 50.060 167.920 ;
        RECT 51.135 167.875 51.425 167.920 ;
        RECT 52.040 168.060 52.360 168.120 ;
        RECT 60.335 168.060 60.625 168.105 ;
        RECT 52.040 167.920 60.625 168.060 ;
        RECT 52.040 167.860 52.360 167.920 ;
        RECT 60.335 167.875 60.625 167.920 ;
        RECT 69.060 168.060 69.380 168.120 ;
        RECT 69.535 168.060 69.825 168.105 ;
        RECT 69.060 167.920 69.825 168.060 ;
        RECT 69.060 167.860 69.380 167.920 ;
        RECT 69.535 167.875 69.825 167.920 ;
        RECT 69.980 167.860 70.300 168.120 ;
        RECT 72.295 168.060 72.585 168.105 ;
        RECT 73.200 168.060 73.520 168.120 ;
        RECT 72.295 167.920 73.520 168.060 ;
        RECT 72.295 167.875 72.585 167.920 ;
        RECT 73.200 167.860 73.520 167.920 ;
        RECT 75.500 167.860 75.820 168.120 ;
        RECT 76.880 167.860 77.200 168.120 ;
        RECT 77.815 168.060 78.105 168.105 ;
        RECT 80.100 168.060 80.420 168.120 ;
        RECT 77.815 167.920 80.420 168.060 ;
        RECT 77.815 167.875 78.105 167.920 ;
        RECT 80.100 167.860 80.420 167.920 ;
        RECT 104.480 168.060 104.800 168.120 ;
        RECT 106.795 168.060 107.085 168.105 ;
        RECT 110.920 168.060 111.240 168.120 ;
        RECT 116.900 168.060 117.220 168.120 ;
        RECT 104.480 167.920 117.220 168.060 ;
        RECT 104.480 167.860 104.800 167.920 ;
        RECT 106.795 167.875 107.085 167.920 ;
        RECT 110.920 167.860 111.240 167.920 ;
        RECT 116.900 167.860 117.220 167.920 ;
        RECT 123.800 168.060 124.120 168.120 ;
        RECT 124.275 168.060 124.565 168.105 ;
        RECT 123.800 167.920 124.565 168.060 ;
        RECT 123.800 167.860 124.120 167.920 ;
        RECT 124.275 167.875 124.565 167.920 ;
        RECT 133.460 167.860 133.780 168.120 ;
        RECT 134.840 167.860 135.160 168.120 ;
        RECT 29.515 167.720 29.805 167.765 ;
        RECT 30.895 167.720 31.185 167.765 ;
        RECT 21.540 167.580 24.210 167.720 ;
        RECT 19.840 167.380 20.160 167.440 ;
        RECT 21.540 167.380 21.680 167.580 ;
        RECT 19.840 167.240 21.680 167.380 ;
        RECT 22.600 167.425 22.920 167.440 ;
        RECT 24.070 167.425 24.210 167.580 ;
        RECT 29.515 167.580 31.185 167.720 ;
        RECT 29.515 167.535 29.805 167.580 ;
        RECT 30.895 167.535 31.185 167.580 ;
        RECT 31.355 167.535 31.645 167.765 ;
        RECT 36.400 167.720 36.720 167.780 ;
        RECT 40.080 167.720 40.400 167.780 ;
        RECT 31.890 167.580 36.720 167.720 ;
        RECT 22.600 167.380 22.950 167.425 ;
        RECT 22.600 167.240 23.115 167.380 ;
        RECT 19.840 167.180 20.160 167.240 ;
        RECT 22.600 167.195 22.950 167.240 ;
        RECT 23.995 167.195 24.285 167.425 ;
        RECT 22.600 167.180 22.920 167.195 ;
        RECT 27.660 167.180 27.980 167.440 ;
        RECT 28.120 167.380 28.440 167.440 ;
        RECT 28.120 167.240 28.635 167.380 ;
        RECT 28.120 167.180 28.440 167.240 ;
        RECT 29.960 167.180 30.280 167.440 ;
        RECT 31.890 167.425 32.030 167.580 ;
        RECT 36.400 167.520 36.720 167.580 ;
        RECT 36.950 167.580 40.400 167.720 ;
        RECT 31.815 167.195 32.105 167.425 ;
        RECT 35.480 167.380 35.770 167.425 ;
        RECT 36.950 167.380 37.090 167.580 ;
        RECT 40.080 167.520 40.400 167.580 ;
        RECT 44.220 167.720 44.540 167.780 ;
        RECT 47.440 167.720 47.760 167.780 ;
        RECT 49.830 167.720 49.970 167.860 ;
        RECT 59.400 167.765 59.720 167.780 ;
        RECT 44.220 167.580 49.970 167.720 ;
        RECT 44.220 167.520 44.540 167.580 ;
        RECT 35.480 167.240 37.090 167.380 ;
        RECT 35.480 167.195 35.770 167.240 ;
        RECT 37.320 167.180 37.640 167.440 ;
        RECT 37.780 167.180 38.100 167.440 ;
        RECT 42.380 167.180 42.700 167.440 ;
        RECT 43.760 167.180 44.080 167.440 ;
        RECT 46.150 167.425 46.290 167.580 ;
        RECT 47.440 167.520 47.760 167.580 ;
        RECT 59.290 167.535 59.720 167.765 ;
        RECT 59.400 167.520 59.720 167.535 ;
        RECT 59.860 167.520 60.180 167.780 ;
        RECT 70.070 167.720 70.210 167.860 ;
        RECT 75.040 167.720 75.360 167.780 ;
        RECT 70.070 167.580 75.360 167.720 ;
        RECT 45.155 167.195 45.445 167.425 ;
        RECT 46.075 167.195 46.365 167.425 ;
        RECT 19.405 167.040 19.695 167.085 ;
        RECT 21.925 167.040 22.215 167.085 ;
        RECT 23.115 167.040 23.405 167.085 ;
        RECT 19.405 166.900 23.405 167.040 ;
        RECT 19.405 166.855 19.695 166.900 ;
        RECT 21.925 166.855 22.215 166.900 ;
        RECT 23.115 166.855 23.405 166.900 ;
        RECT 41.475 167.040 41.765 167.085 ;
        RECT 42.840 167.040 43.160 167.100 ;
        RECT 41.475 166.900 43.160 167.040 ;
        RECT 41.475 166.855 41.765 166.900 ;
        RECT 42.840 166.840 43.160 166.900 ;
        RECT 43.300 167.040 43.620 167.100 ;
        RECT 45.230 167.040 45.370 167.195 ;
        RECT 46.980 167.180 47.300 167.440 ;
        RECT 49.880 167.380 50.170 167.425 ;
        RECT 50.660 167.380 50.980 167.440 ;
        RECT 49.880 167.240 50.980 167.380 ;
        RECT 49.880 167.195 50.170 167.240 ;
        RECT 50.660 167.180 50.980 167.240 ;
        RECT 56.755 167.380 57.045 167.425 ;
        RECT 69.060 167.380 69.380 167.440 ;
        RECT 69.995 167.380 70.285 167.425 ;
        RECT 56.755 167.240 59.170 167.380 ;
        RECT 56.755 167.195 57.045 167.240 ;
        RECT 43.300 166.900 45.370 167.040 ;
        RECT 46.520 167.040 46.840 167.100 ;
        RECT 47.455 167.040 47.745 167.085 ;
        RECT 46.520 166.900 47.745 167.040 ;
        RECT 43.300 166.840 43.620 166.900 ;
        RECT 46.520 166.840 46.840 166.900 ;
        RECT 47.455 166.855 47.745 166.900 ;
        RECT 48.820 166.840 49.140 167.100 ;
        RECT 53.445 167.040 53.735 167.085 ;
        RECT 55.965 167.040 56.255 167.085 ;
        RECT 57.155 167.040 57.445 167.085 ;
        RECT 53.445 166.900 57.445 167.040 ;
        RECT 53.445 166.855 53.735 166.900 ;
        RECT 55.965 166.855 56.255 166.900 ;
        RECT 57.155 166.855 57.445 166.900 ;
        RECT 58.035 167.040 58.325 167.085 ;
        RECT 58.480 167.040 58.800 167.100 ;
        RECT 58.035 166.900 58.800 167.040 ;
        RECT 58.035 166.855 58.325 166.900 ;
        RECT 58.480 166.840 58.800 166.900 ;
        RECT 19.840 166.700 20.130 166.745 ;
        RECT 21.410 166.700 21.700 166.745 ;
        RECT 23.510 166.700 23.800 166.745 ;
        RECT 19.840 166.560 23.800 166.700 ;
        RECT 19.840 166.515 20.130 166.560 ;
        RECT 21.410 166.515 21.700 166.560 ;
        RECT 23.510 166.515 23.800 166.560 ;
        RECT 44.235 166.700 44.525 166.745 ;
        RECT 48.910 166.700 49.050 166.840 ;
        RECT 44.235 166.560 49.050 166.700 ;
        RECT 50.675 166.700 50.965 166.745 ;
        RECT 53.880 166.700 54.170 166.745 ;
        RECT 55.450 166.700 55.740 166.745 ;
        RECT 57.550 166.700 57.840 166.745 ;
        RECT 59.030 166.700 59.170 167.240 ;
        RECT 69.060 167.240 70.285 167.380 ;
        RECT 69.060 167.180 69.380 167.240 ;
        RECT 69.995 167.195 70.285 167.240 ;
        RECT 71.375 167.195 71.665 167.425 ;
        RECT 60.320 167.040 60.640 167.100 ;
        RECT 61.715 167.040 62.005 167.085 ;
        RECT 60.320 166.900 62.005 167.040 ;
        RECT 60.320 166.840 60.640 166.900 ;
        RECT 61.715 166.855 62.005 166.900 ;
        RECT 67.235 167.040 67.525 167.085 ;
        RECT 69.520 167.040 69.840 167.100 ;
        RECT 67.235 166.900 69.840 167.040 ;
        RECT 67.235 166.855 67.525 166.900 ;
        RECT 69.520 166.840 69.840 166.900 ;
        RECT 70.900 166.840 71.220 167.100 ;
        RECT 71.450 167.040 71.590 167.195 ;
        RECT 72.740 167.180 73.060 167.440 ;
        RECT 73.290 167.425 73.430 167.580 ;
        RECT 75.040 167.520 75.360 167.580 ;
        RECT 85.620 167.765 85.940 167.780 ;
        RECT 85.620 167.720 85.970 167.765 ;
        RECT 97.750 167.720 98.040 167.765 ;
        RECT 99.435 167.720 99.725 167.765 ;
        RECT 109.095 167.720 109.385 167.765 ;
        RECT 123.355 167.720 123.645 167.765 ;
        RECT 127.910 167.720 128.200 167.765 ;
        RECT 129.780 167.720 130.100 167.780 ;
        RECT 85.620 167.580 86.135 167.720 ;
        RECT 97.750 167.580 99.725 167.720 ;
        RECT 85.620 167.535 85.970 167.580 ;
        RECT 97.750 167.535 98.040 167.580 ;
        RECT 99.435 167.535 99.725 167.580 ;
        RECT 101.810 167.580 118.050 167.720 ;
        RECT 85.620 167.520 85.940 167.535 ;
        RECT 73.215 167.195 73.505 167.425 ;
        RECT 73.660 167.380 73.980 167.440 ;
        RECT 74.135 167.380 74.425 167.425 ;
        RECT 73.660 167.240 74.425 167.380 ;
        RECT 73.660 167.180 73.980 167.240 ;
        RECT 74.135 167.195 74.425 167.240 ;
        RECT 74.595 167.380 74.885 167.425 ;
        RECT 77.800 167.380 78.120 167.440 ;
        RECT 74.595 167.240 78.120 167.380 ;
        RECT 74.595 167.195 74.885 167.240 ;
        RECT 77.800 167.180 78.120 167.240 ;
        RECT 79.640 167.180 79.960 167.440 ;
        RECT 86.540 167.380 86.860 167.440 ;
        RECT 87.015 167.380 87.305 167.425 ;
        RECT 86.540 167.240 87.305 167.380 ;
        RECT 86.540 167.180 86.860 167.240 ;
        RECT 87.015 167.195 87.305 167.240 ;
        RECT 98.500 167.380 98.820 167.440 ;
        RECT 98.975 167.380 99.265 167.425 ;
        RECT 98.500 167.240 99.265 167.380 ;
        RECT 98.500 167.180 98.820 167.240 ;
        RECT 98.975 167.195 99.265 167.240 ;
        RECT 100.355 167.195 100.645 167.425 ;
        RECT 75.960 167.040 76.280 167.100 ;
        RECT 71.450 166.900 76.280 167.040 ;
        RECT 75.960 166.840 76.280 166.900 ;
        RECT 82.425 167.040 82.715 167.085 ;
        RECT 84.945 167.040 85.235 167.085 ;
        RECT 86.135 167.040 86.425 167.085 ;
        RECT 82.425 166.900 86.425 167.040 ;
        RECT 82.425 166.855 82.715 166.900 ;
        RECT 84.945 166.855 85.235 166.900 ;
        RECT 86.135 166.855 86.425 166.900 ;
        RECT 94.385 167.040 94.675 167.085 ;
        RECT 96.905 167.040 97.195 167.085 ;
        RECT 98.095 167.040 98.385 167.085 ;
        RECT 94.385 166.900 98.385 167.040 ;
        RECT 100.430 167.040 100.570 167.195 ;
        RECT 100.800 167.180 101.120 167.440 ;
        RECT 101.810 167.085 101.950 167.580 ;
        RECT 109.095 167.535 109.385 167.580 ;
        RECT 102.195 167.380 102.485 167.425 ;
        RECT 103.100 167.380 103.420 167.440 ;
        RECT 102.195 167.240 103.420 167.380 ;
        RECT 102.195 167.195 102.485 167.240 ;
        RECT 103.100 167.180 103.420 167.240 ;
        RECT 105.860 167.180 106.180 167.440 ;
        RECT 107.240 167.380 107.560 167.440 ;
        RECT 108.175 167.380 108.465 167.425 ;
        RECT 107.240 167.240 108.465 167.380 ;
        RECT 107.240 167.180 107.560 167.240 ;
        RECT 108.175 167.195 108.465 167.240 ;
        RECT 108.620 167.180 108.940 167.440 ;
        RECT 109.555 167.195 109.845 167.425 ;
        RECT 110.015 167.195 110.305 167.425 ;
        RECT 100.430 166.900 101.030 167.040 ;
        RECT 94.385 166.855 94.675 166.900 ;
        RECT 96.905 166.855 97.195 166.900 ;
        RECT 98.095 166.855 98.385 166.900 ;
        RECT 50.675 166.560 53.650 166.700 ;
        RECT 44.235 166.515 44.525 166.560 ;
        RECT 50.675 166.515 50.965 166.560 ;
        RECT 34.575 166.360 34.865 166.405 ;
        RECT 45.140 166.360 45.460 166.420 ;
        RECT 34.575 166.220 45.460 166.360 ;
        RECT 34.575 166.175 34.865 166.220 ;
        RECT 45.140 166.160 45.460 166.220 ;
        RECT 46.535 166.360 46.825 166.405 ;
        RECT 50.200 166.360 50.520 166.420 ;
        RECT 46.535 166.220 50.520 166.360 ;
        RECT 53.510 166.360 53.650 166.560 ;
        RECT 53.880 166.560 57.840 166.700 ;
        RECT 53.880 166.515 54.170 166.560 ;
        RECT 55.450 166.515 55.740 166.560 ;
        RECT 57.550 166.515 57.840 166.560 ;
        RECT 58.570 166.560 59.170 166.700 ;
        RECT 69.075 166.700 69.365 166.745 ;
        RECT 72.280 166.700 72.600 166.760 ;
        RECT 69.075 166.560 72.600 166.700 ;
        RECT 58.020 166.360 58.340 166.420 ;
        RECT 58.570 166.405 58.710 166.560 ;
        RECT 69.075 166.515 69.365 166.560 ;
        RECT 72.280 166.500 72.600 166.560 ;
        RECT 82.860 166.700 83.150 166.745 ;
        RECT 84.430 166.700 84.720 166.745 ;
        RECT 86.530 166.700 86.820 166.745 ;
        RECT 82.860 166.560 86.820 166.700 ;
        RECT 82.860 166.515 83.150 166.560 ;
        RECT 84.430 166.515 84.720 166.560 ;
        RECT 86.530 166.515 86.820 166.560 ;
        RECT 94.820 166.700 95.110 166.745 ;
        RECT 96.390 166.700 96.680 166.745 ;
        RECT 98.490 166.700 98.780 166.745 ;
        RECT 94.820 166.560 98.780 166.700 ;
        RECT 94.820 166.515 95.110 166.560 ;
        RECT 96.390 166.515 96.680 166.560 ;
        RECT 98.490 166.515 98.780 166.560 ;
        RECT 53.510 166.220 58.340 166.360 ;
        RECT 46.535 166.175 46.825 166.220 ;
        RECT 50.200 166.160 50.520 166.220 ;
        RECT 58.020 166.160 58.340 166.220 ;
        RECT 58.495 166.175 58.785 166.405 ;
        RECT 67.220 166.360 67.540 166.420 ;
        RECT 69.995 166.360 70.285 166.405 ;
        RECT 67.220 166.220 70.285 166.360 ;
        RECT 67.220 166.160 67.540 166.220 ;
        RECT 69.995 166.175 70.285 166.220 ;
        RECT 70.440 166.360 70.760 166.420 ;
        RECT 77.815 166.360 78.105 166.405 ;
        RECT 70.440 166.220 78.105 166.360 ;
        RECT 70.440 166.160 70.760 166.220 ;
        RECT 77.815 166.175 78.105 166.220 ;
        RECT 92.060 166.160 92.380 166.420 ;
        RECT 100.890 166.360 101.030 166.900 ;
        RECT 101.735 166.855 102.025 167.085 ;
        RECT 104.940 167.040 105.260 167.100 ;
        RECT 107.715 167.040 108.005 167.085 ;
        RECT 108.710 167.040 108.850 167.180 ;
        RECT 104.940 166.900 108.850 167.040 ;
        RECT 109.080 167.040 109.400 167.100 ;
        RECT 109.630 167.040 109.770 167.195 ;
        RECT 109.080 166.900 109.770 167.040 ;
        RECT 110.090 167.040 110.230 167.195 ;
        RECT 110.460 167.180 110.780 167.440 ;
        RECT 110.935 167.195 111.225 167.425 ;
        RECT 111.010 167.040 111.150 167.195 ;
        RECT 111.380 167.180 111.700 167.440 ;
        RECT 112.300 167.180 112.620 167.440 ;
        RECT 115.060 167.380 115.380 167.440 ;
        RECT 115.535 167.380 115.825 167.425 ;
        RECT 113.310 167.240 115.825 167.380 ;
        RECT 111.855 167.040 112.145 167.085 ;
        RECT 113.310 167.040 113.450 167.240 ;
        RECT 115.060 167.180 115.380 167.240 ;
        RECT 115.535 167.195 115.825 167.240 ;
        RECT 115.980 167.180 116.300 167.440 ;
        RECT 116.900 167.180 117.220 167.440 ;
        RECT 117.375 167.195 117.665 167.425 ;
        RECT 110.090 166.900 110.690 167.040 ;
        RECT 111.010 166.900 113.450 167.040 ;
        RECT 104.940 166.840 105.260 166.900 ;
        RECT 107.715 166.855 108.005 166.900 ;
        RECT 109.080 166.840 109.400 166.900 ;
        RECT 108.160 166.700 108.480 166.760 ;
        RECT 110.550 166.700 110.690 166.900 ;
        RECT 111.855 166.855 112.145 166.900 ;
        RECT 113.680 166.840 114.000 167.100 ;
        RECT 117.450 167.040 117.590 167.195 ;
        RECT 116.990 166.900 117.590 167.040 ;
        RECT 117.910 167.040 118.050 167.580 ;
        RECT 123.355 167.580 126.790 167.720 ;
        RECT 123.355 167.535 123.645 167.580 ;
        RECT 126.650 167.440 126.790 167.580 ;
        RECT 127.910 167.580 130.100 167.720 ;
        RECT 127.910 167.535 128.200 167.580 ;
        RECT 129.780 167.520 130.100 167.580 ;
        RECT 119.200 167.180 119.520 167.440 ;
        RECT 121.500 167.380 121.820 167.440 ;
        RECT 124.275 167.380 124.565 167.425 ;
        RECT 121.500 167.240 124.565 167.380 ;
        RECT 121.500 167.180 121.820 167.240 ;
        RECT 124.275 167.195 124.565 167.240 ;
        RECT 125.195 167.195 125.485 167.425 ;
        RECT 125.270 167.040 125.410 167.195 ;
        RECT 126.560 167.180 126.880 167.440 ;
        RECT 133.935 167.380 134.225 167.425 ;
        RECT 134.380 167.380 134.700 167.440 ;
        RECT 133.935 167.240 134.700 167.380 ;
        RECT 133.935 167.195 134.225 167.240 ;
        RECT 134.380 167.180 134.700 167.240 ;
        RECT 135.760 167.180 136.080 167.440 ;
        RECT 117.910 166.900 125.410 167.040 ;
        RECT 127.455 167.040 127.745 167.085 ;
        RECT 128.645 167.040 128.935 167.085 ;
        RECT 131.165 167.040 131.455 167.085 ;
        RECT 127.455 166.900 131.455 167.040 ;
        RECT 108.160 166.560 114.370 166.700 ;
        RECT 108.160 166.500 108.480 166.560 ;
        RECT 114.230 166.420 114.370 166.560 ;
        RECT 114.600 166.500 114.920 166.760 ;
        RECT 116.990 166.700 117.130 166.900 ;
        RECT 127.455 166.855 127.745 166.900 ;
        RECT 128.645 166.855 128.935 166.900 ;
        RECT 131.165 166.855 131.455 166.900 ;
        RECT 117.360 166.700 117.680 166.760 ;
        RECT 121.500 166.700 121.820 166.760 ;
        RECT 116.990 166.560 121.820 166.700 ;
        RECT 117.360 166.500 117.680 166.560 ;
        RECT 121.500 166.500 121.820 166.560 ;
        RECT 127.060 166.700 127.350 166.745 ;
        RECT 129.160 166.700 129.450 166.745 ;
        RECT 130.730 166.700 131.020 166.745 ;
        RECT 127.060 166.560 131.020 166.700 ;
        RECT 127.060 166.515 127.350 166.560 ;
        RECT 129.160 166.515 129.450 166.560 ;
        RECT 130.730 166.515 131.020 166.560 ;
        RECT 110.000 166.360 110.320 166.420 ;
        RECT 100.890 166.220 110.320 166.360 ;
        RECT 110.000 166.160 110.320 166.220 ;
        RECT 114.140 166.360 114.460 166.420 ;
        RECT 115.980 166.360 116.300 166.420 ;
        RECT 116.915 166.360 117.205 166.405 ;
        RECT 114.140 166.220 117.205 166.360 ;
        RECT 114.140 166.160 114.460 166.220 ;
        RECT 115.980 166.160 116.300 166.220 ;
        RECT 116.915 166.175 117.205 166.220 ;
        RECT 118.280 166.360 118.600 166.420 ;
        RECT 118.755 166.360 119.045 166.405 ;
        RECT 118.280 166.220 119.045 166.360 ;
        RECT 118.280 166.160 118.600 166.220 ;
        RECT 118.755 166.175 119.045 166.220 ;
        RECT 136.680 166.160 137.000 166.420 ;
        RECT 13.330 165.540 138.910 166.020 ;
        RECT 21.680 165.340 22.000 165.400 ;
        RECT 22.615 165.340 22.905 165.385 ;
        RECT 27.660 165.340 27.980 165.400 ;
        RECT 21.680 165.200 27.980 165.340 ;
        RECT 21.680 165.140 22.000 165.200 ;
        RECT 22.615 165.155 22.905 165.200 ;
        RECT 27.660 165.140 27.980 165.200 ;
        RECT 34.560 165.340 34.880 165.400 ;
        RECT 35.035 165.340 35.325 165.385 ;
        RECT 41.920 165.340 42.240 165.400 ;
        RECT 34.560 165.200 35.325 165.340 ;
        RECT 34.560 165.140 34.880 165.200 ;
        RECT 35.035 165.155 35.325 165.200 ;
        RECT 35.555 165.200 42.240 165.340 ;
        RECT 16.200 165.000 16.490 165.045 ;
        RECT 18.300 165.000 18.590 165.045 ;
        RECT 19.870 165.000 20.160 165.045 ;
        RECT 16.200 164.860 20.160 165.000 ;
        RECT 16.200 164.815 16.490 164.860 ;
        RECT 18.300 164.815 18.590 164.860 ;
        RECT 19.870 164.815 20.160 164.860 ;
        RECT 28.580 165.000 28.900 165.060 ;
        RECT 35.555 165.000 35.695 165.200 ;
        RECT 41.920 165.140 42.240 165.200 ;
        RECT 42.380 165.340 42.700 165.400 ;
        RECT 45.155 165.340 45.445 165.385 ;
        RECT 42.380 165.200 45.445 165.340 ;
        RECT 42.380 165.140 42.700 165.200 ;
        RECT 45.155 165.155 45.445 165.200 ;
        RECT 51.135 165.340 51.425 165.385 ;
        RECT 56.180 165.340 56.500 165.400 ;
        RECT 51.135 165.200 56.500 165.340 ;
        RECT 51.135 165.155 51.425 165.200 ;
        RECT 56.180 165.140 56.500 165.200 ;
        RECT 69.995 165.340 70.285 165.385 ;
        RECT 70.440 165.340 70.760 165.400 ;
        RECT 69.995 165.200 70.760 165.340 ;
        RECT 69.995 165.155 70.285 165.200 ;
        RECT 70.440 165.140 70.760 165.200 ;
        RECT 70.900 165.140 71.220 165.400 ;
        RECT 73.675 165.340 73.965 165.385 ;
        RECT 74.580 165.340 74.900 165.400 ;
        RECT 73.675 165.200 74.900 165.340 ;
        RECT 73.675 165.155 73.965 165.200 ;
        RECT 74.580 165.140 74.900 165.200 ;
        RECT 78.260 165.140 78.580 165.400 ;
        RECT 83.780 165.340 84.100 165.400 ;
        RECT 83.780 165.200 88.150 165.340 ;
        RECT 83.780 165.140 84.100 165.200 ;
        RECT 28.580 164.860 35.695 165.000 ;
        RECT 39.635 165.000 39.925 165.045 ;
        RECT 43.760 165.000 44.080 165.060 ;
        RECT 39.635 164.860 44.080 165.000 ;
        RECT 28.580 164.800 28.900 164.860 ;
        RECT 39.635 164.815 39.925 164.860 ;
        RECT 43.760 164.800 44.080 164.860 ;
        RECT 46.520 165.000 46.840 165.060 ;
        RECT 46.520 164.860 48.130 165.000 ;
        RECT 46.520 164.800 46.840 164.860 ;
        RECT 16.595 164.660 16.885 164.705 ;
        RECT 17.785 164.660 18.075 164.705 ;
        RECT 20.305 164.660 20.595 164.705 ;
        RECT 39.160 164.660 39.480 164.720 ;
        RECT 43.315 164.660 43.605 164.705 ;
        RECT 44.680 164.660 45.000 164.720 ;
        RECT 47.990 164.705 48.130 164.860 ;
        RECT 52.500 164.800 52.820 165.060 ;
        RECT 55.260 165.000 55.550 165.045 ;
        RECT 56.830 165.000 57.120 165.045 ;
        RECT 58.930 165.000 59.220 165.045 ;
        RECT 55.260 164.860 59.220 165.000 ;
        RECT 55.260 164.815 55.550 164.860 ;
        RECT 56.830 164.815 57.120 164.860 ;
        RECT 58.930 164.815 59.220 164.860 ;
        RECT 68.140 164.800 68.460 165.060 ;
        RECT 16.595 164.520 20.595 164.660 ;
        RECT 16.595 164.475 16.885 164.520 ;
        RECT 17.785 164.475 18.075 164.520 ;
        RECT 20.305 164.475 20.595 164.520 ;
        RECT 36.030 164.520 42.150 164.660 ;
        RECT 15.715 164.320 16.005 164.365 ;
        RECT 19.380 164.320 19.700 164.380 ;
        RECT 15.715 164.180 19.700 164.320 ;
        RECT 15.715 164.135 16.005 164.180 ;
        RECT 19.380 164.120 19.700 164.180 ;
        RECT 27.660 164.320 27.980 164.380 ;
        RECT 36.030 164.365 36.170 164.520 ;
        RECT 39.160 164.460 39.480 164.520 ;
        RECT 27.660 164.180 29.270 164.320 ;
        RECT 27.660 164.120 27.980 164.180 ;
        RECT 17.050 163.980 17.340 164.025 ;
        RECT 17.540 163.980 17.860 164.040 ;
        RECT 17.050 163.840 17.860 163.980 ;
        RECT 17.050 163.795 17.340 163.840 ;
        RECT 17.540 163.780 17.860 163.840 ;
        RECT 28.580 163.780 28.900 164.040 ;
        RECT 29.130 163.980 29.270 164.180 ;
        RECT 35.955 164.135 36.245 164.365 ;
        RECT 36.860 164.120 37.180 164.380 ;
        RECT 37.335 164.135 37.625 164.365 ;
        RECT 37.410 163.980 37.550 164.135 ;
        RECT 40.540 164.120 40.860 164.380 ;
        RECT 41.015 164.320 41.305 164.365 ;
        RECT 42.010 164.320 42.150 164.520 ;
        RECT 43.315 164.520 46.165 164.660 ;
        RECT 43.315 164.475 43.605 164.520 ;
        RECT 44.680 164.460 45.000 164.520 ;
        RECT 42.855 164.320 43.145 164.365 ;
        RECT 41.015 164.180 41.690 164.320 ;
        RECT 42.010 164.180 43.145 164.320 ;
        RECT 41.015 164.135 41.305 164.180 ;
        RECT 29.130 163.840 37.550 163.980 ;
        RECT 28.135 163.640 28.425 163.685 ;
        RECT 29.960 163.640 30.280 163.700 ;
        RECT 28.135 163.500 30.280 163.640 ;
        RECT 41.550 163.640 41.690 164.180 ;
        RECT 42.855 164.135 43.145 164.180 ;
        RECT 43.760 164.120 44.080 164.380 ;
        RECT 44.220 164.120 44.540 164.380 ;
        RECT 46.025 164.365 46.165 164.520 ;
        RECT 47.915 164.475 48.205 164.705 ;
        RECT 49.280 164.660 49.600 164.720 ;
        RECT 49.755 164.660 50.045 164.705 ;
        RECT 49.280 164.520 50.045 164.660 ;
        RECT 49.280 164.460 49.600 164.520 ;
        RECT 49.755 164.475 50.045 164.520 ;
        RECT 50.340 164.660 50.630 164.705 ;
        RECT 51.580 164.660 51.900 164.720 ;
        RECT 50.340 164.520 51.900 164.660 ;
        RECT 50.340 164.475 50.630 164.520 ;
        RECT 51.580 164.460 51.900 164.520 ;
        RECT 54.825 164.660 55.115 164.705 ;
        RECT 57.345 164.660 57.635 164.705 ;
        RECT 58.535 164.660 58.825 164.705 ;
        RECT 54.825 164.520 58.825 164.660 ;
        RECT 70.530 164.660 70.670 165.140 ;
        RECT 73.215 164.815 73.505 165.045 ;
        RECT 71.375 164.660 71.665 164.705 ;
        RECT 70.530 164.520 71.665 164.660 ;
        RECT 54.825 164.475 55.115 164.520 ;
        RECT 57.345 164.475 57.635 164.520 ;
        RECT 58.535 164.475 58.825 164.520 ;
        RECT 71.375 164.475 71.665 164.520 ;
        RECT 45.735 164.180 46.165 164.365 ;
        RECT 46.535 164.320 46.825 164.365 ;
        RECT 47.440 164.320 47.760 164.380 ;
        RECT 46.535 164.180 47.760 164.320 ;
        RECT 45.735 164.135 46.025 164.180 ;
        RECT 46.535 164.135 46.825 164.180 ;
        RECT 47.440 164.120 47.760 164.180 ;
        RECT 58.020 164.365 58.340 164.380 ;
        RECT 58.020 164.320 58.370 164.365 ;
        RECT 58.940 164.320 59.260 164.380 ;
        RECT 59.415 164.320 59.705 164.365 ;
        RECT 66.775 164.320 67.065 164.365 ;
        RECT 58.020 164.180 58.535 164.320 ;
        RECT 58.940 164.180 59.705 164.320 ;
        RECT 58.020 164.135 58.370 164.180 ;
        RECT 58.020 164.120 58.340 164.135 ;
        RECT 58.940 164.120 59.260 164.180 ;
        RECT 59.415 164.135 59.705 164.180 ;
        RECT 62.710 164.180 67.065 164.320 ;
        RECT 41.935 163.980 42.225 164.025 ;
        RECT 49.295 163.980 49.585 164.025 ;
        RECT 51.120 163.980 51.440 164.040 ;
        RECT 41.935 163.840 45.830 163.980 ;
        RECT 41.935 163.795 42.225 163.840 ;
        RECT 45.690 163.700 45.830 163.840 ;
        RECT 49.295 163.840 51.440 163.980 ;
        RECT 59.490 163.980 59.630 164.135 ;
        RECT 62.710 164.040 62.850 164.180 ;
        RECT 66.775 164.135 67.065 164.180 ;
        RECT 60.795 163.980 61.085 164.025 ;
        RECT 62.620 163.980 62.940 164.040 ;
        RECT 59.490 163.840 62.940 163.980 ;
        RECT 49.295 163.795 49.585 163.840 ;
        RECT 51.120 163.780 51.440 163.840 ;
        RECT 60.795 163.795 61.085 163.840 ;
        RECT 62.620 163.780 62.940 163.840 ;
        RECT 63.080 163.780 63.400 164.040 ;
        RECT 73.290 163.980 73.430 164.815 ;
        RECT 74.595 164.660 74.885 164.705 ;
        RECT 78.350 164.660 78.490 165.140 ;
        RECT 81.020 165.000 81.310 165.045 ;
        RECT 82.590 165.000 82.880 165.045 ;
        RECT 84.690 165.000 84.980 165.045 ;
        RECT 81.020 164.860 84.980 165.000 ;
        RECT 88.010 165.000 88.150 165.200 ;
        RECT 97.120 165.140 97.440 165.400 ;
        RECT 104.480 165.140 104.800 165.400 ;
        RECT 106.780 165.340 107.100 165.400 ;
        RECT 110.460 165.340 110.780 165.400 ;
        RECT 106.780 165.200 110.780 165.340 ;
        RECT 106.780 165.140 107.100 165.200 ;
        RECT 110.460 165.140 110.780 165.200 ;
        RECT 112.760 165.340 113.080 165.400 ;
        RECT 114.140 165.340 114.460 165.400 ;
        RECT 112.760 165.200 114.460 165.340 ;
        RECT 112.760 165.140 113.080 165.200 ;
        RECT 114.140 165.140 114.460 165.200 ;
        RECT 115.535 165.340 115.825 165.385 ;
        RECT 125.640 165.340 125.960 165.400 ;
        RECT 115.535 165.200 125.960 165.340 ;
        RECT 115.535 165.155 115.825 165.200 ;
        RECT 125.640 165.140 125.960 165.200 ;
        RECT 93.900 165.000 94.220 165.060 ;
        RECT 119.200 165.000 119.520 165.060 ;
        RECT 88.010 164.860 88.610 165.000 ;
        RECT 81.020 164.815 81.310 164.860 ;
        RECT 82.590 164.815 82.880 164.860 ;
        RECT 84.690 164.815 84.980 164.860 ;
        RECT 88.470 164.720 88.610 164.860 ;
        RECT 92.610 164.860 119.520 165.000 ;
        RECT 74.595 164.520 78.490 164.660 ;
        RECT 80.585 164.660 80.875 164.705 ;
        RECT 83.105 164.660 83.395 164.705 ;
        RECT 84.295 164.660 84.585 164.705 ;
        RECT 87.935 164.660 88.225 164.705 ;
        RECT 80.585 164.520 84.585 164.660 ;
        RECT 74.595 164.475 74.885 164.520 ;
        RECT 80.585 164.475 80.875 164.520 ;
        RECT 83.105 164.475 83.395 164.520 ;
        RECT 84.295 164.475 84.585 164.520 ;
        RECT 84.790 164.520 88.225 164.660 ;
        RECT 77.355 164.320 77.645 164.365 ;
        RECT 84.790 164.320 84.930 164.520 ;
        RECT 87.935 164.475 88.225 164.520 ;
        RECT 88.380 164.460 88.700 164.720 ;
        RECT 77.355 164.180 84.930 164.320 ;
        RECT 77.355 164.135 77.645 164.180 ;
        RECT 85.160 164.120 85.480 164.380 ;
        RECT 90.680 164.320 91.000 164.380 ;
        RECT 92.075 164.320 92.365 164.365 ;
        RECT 92.610 164.320 92.750 164.860 ;
        RECT 93.900 164.800 94.220 164.860 ;
        RECT 119.200 164.800 119.520 164.860 ;
        RECT 99.420 164.460 99.740 164.720 ;
        RECT 99.895 164.475 100.185 164.705 ;
        RECT 90.680 164.180 92.750 164.320 ;
        RECT 94.360 164.320 94.680 164.380 ;
        RECT 97.120 164.320 97.440 164.380 ;
        RECT 99.970 164.320 100.110 164.475 ;
        RECT 105.400 164.460 105.720 164.720 ;
        RECT 112.300 164.660 112.620 164.720 ;
        RECT 113.695 164.660 113.985 164.705 ;
        RECT 115.980 164.660 116.300 164.720 ;
        RECT 112.300 164.520 113.985 164.660 ;
        RECT 112.300 164.460 112.620 164.520 ;
        RECT 113.695 164.475 113.985 164.520 ;
        RECT 114.230 164.520 116.300 164.660 ;
        RECT 94.360 164.180 100.110 164.320 ;
        RECT 104.020 164.320 104.340 164.380 ;
        RECT 106.335 164.320 106.625 164.365 ;
        RECT 104.020 164.180 111.610 164.320 ;
        RECT 90.680 164.120 91.000 164.180 ;
        RECT 92.075 164.135 92.365 164.180 ;
        RECT 94.360 164.120 94.680 164.180 ;
        RECT 97.120 164.120 97.440 164.180 ;
        RECT 104.020 164.120 104.340 164.180 ;
        RECT 106.335 164.135 106.625 164.180 ;
        RECT 80.560 163.980 80.880 164.040 ;
        RECT 73.290 163.840 80.880 163.980 ;
        RECT 80.560 163.780 80.880 163.840 ;
        RECT 83.950 163.980 84.240 164.025 ;
        RECT 83.950 163.840 85.850 163.980 ;
        RECT 83.950 163.795 84.240 163.840 ;
        RECT 43.760 163.640 44.080 163.700 ;
        RECT 41.550 163.500 44.080 163.640 ;
        RECT 28.135 163.455 28.425 163.500 ;
        RECT 29.960 163.440 30.280 163.500 ;
        RECT 43.760 163.440 44.080 163.500 ;
        RECT 45.600 163.440 45.920 163.700 ;
        RECT 46.060 163.440 46.380 163.700 ;
        RECT 69.980 163.440 70.300 163.700 ;
        RECT 85.710 163.685 85.850 163.840 ;
        RECT 95.740 163.780 96.060 164.040 ;
        RECT 85.635 163.455 85.925 163.685 ;
        RECT 87.460 163.440 87.780 163.700 ;
        RECT 98.960 163.440 99.280 163.700 ;
        RECT 105.415 163.640 105.705 163.685 ;
        RECT 106.320 163.640 106.640 163.700 ;
        RECT 105.415 163.500 106.640 163.640 ;
        RECT 111.470 163.640 111.610 164.180 ;
        RECT 111.855 164.135 112.145 164.365 ;
        RECT 111.930 163.980 112.070 164.135 ;
        RECT 112.760 164.120 113.080 164.380 ;
        RECT 113.235 164.330 113.525 164.365 ;
        RECT 114.230 164.330 114.370 164.520 ;
        RECT 115.980 164.460 116.300 164.520 ;
        RECT 129.320 164.660 129.640 164.720 ;
        RECT 132.555 164.660 132.845 164.705 ;
        RECT 129.320 164.520 132.845 164.660 ;
        RECT 129.320 164.460 129.640 164.520 ;
        RECT 132.555 164.475 132.845 164.520 ;
        RECT 113.235 164.190 114.370 164.330 ;
        RECT 114.615 164.320 114.905 164.365 ;
        RECT 115.520 164.320 115.840 164.380 ;
        RECT 113.235 164.135 113.525 164.190 ;
        RECT 114.615 164.180 115.840 164.320 ;
        RECT 114.615 164.135 114.905 164.180 ;
        RECT 115.520 164.120 115.840 164.180 ;
        RECT 116.440 164.320 116.760 164.380 ;
        RECT 116.915 164.320 117.205 164.365 ;
        RECT 116.440 164.180 117.205 164.320 ;
        RECT 116.440 164.120 116.760 164.180 ;
        RECT 116.915 164.135 117.205 164.180 ;
        RECT 117.360 164.120 117.680 164.380 ;
        RECT 119.215 164.320 119.505 164.365 ;
        RECT 126.560 164.320 126.880 164.380 ;
        RECT 119.215 164.180 126.880 164.320 ;
        RECT 119.215 164.135 119.505 164.180 ;
        RECT 126.560 164.120 126.880 164.180 ;
        RECT 133.460 164.320 133.780 164.380 ;
        RECT 136.695 164.320 136.985 164.365 ;
        RECT 133.460 164.180 136.985 164.320 ;
        RECT 133.460 164.120 133.780 164.180 ;
        RECT 136.695 164.135 136.985 164.180 ;
        RECT 113.680 163.980 114.000 164.040 ;
        RECT 111.930 163.840 114.000 163.980 ;
        RECT 113.680 163.780 114.000 163.840 ;
        RECT 114.140 163.980 114.460 164.040 ;
        RECT 115.995 163.980 116.285 164.025 ;
        RECT 117.450 163.980 117.590 164.120 ;
        RECT 114.140 163.840 116.285 163.980 ;
        RECT 114.140 163.780 114.460 163.840 ;
        RECT 115.995 163.795 116.285 163.840 ;
        RECT 116.530 163.840 117.590 163.980 ;
        RECT 131.635 163.980 131.925 164.025 ;
        RECT 133.935 163.980 134.225 164.025 ;
        RECT 131.635 163.840 134.225 163.980 ;
        RECT 116.530 163.640 116.670 163.840 ;
        RECT 131.635 163.795 131.925 163.840 ;
        RECT 133.935 163.795 134.225 163.840 ;
        RECT 111.470 163.500 116.670 163.640 ;
        RECT 105.415 163.455 105.705 163.500 ;
        RECT 106.320 163.440 106.640 163.500 ;
        RECT 117.360 163.440 117.680 163.700 ;
        RECT 127.940 163.640 128.260 163.700 ;
        RECT 129.795 163.640 130.085 163.685 ;
        RECT 127.940 163.500 130.085 163.640 ;
        RECT 127.940 163.440 128.260 163.500 ;
        RECT 129.795 163.455 130.085 163.500 ;
        RECT 130.240 163.640 130.560 163.700 ;
        RECT 132.095 163.640 132.385 163.685 ;
        RECT 130.240 163.500 132.385 163.640 ;
        RECT 130.240 163.440 130.560 163.500 ;
        RECT 132.095 163.455 132.385 163.500 ;
        RECT 13.330 162.820 138.910 163.300 ;
        RECT 26.740 162.620 27.060 162.680 ;
        RECT 23.610 162.480 27.060 162.620 ;
        RECT 23.610 161.985 23.750 162.480 ;
        RECT 26.740 162.420 27.060 162.480 ;
        RECT 30.880 162.420 31.200 162.680 ;
        RECT 44.235 162.435 44.525 162.665 ;
        RECT 49.295 162.620 49.585 162.665 ;
        RECT 50.660 162.620 50.980 162.680 ;
        RECT 49.295 162.480 50.980 162.620 ;
        RECT 49.295 162.435 49.585 162.480 ;
        RECT 44.310 162.280 44.450 162.435 ;
        RECT 50.660 162.420 50.980 162.480 ;
        RECT 63.080 162.620 63.400 162.680 ;
        RECT 81.480 162.620 81.800 162.680 ;
        RECT 90.680 162.620 91.000 162.680 ;
        RECT 113.220 162.620 113.540 162.680 ;
        RECT 63.080 162.480 91.000 162.620 ;
        RECT 63.080 162.420 63.400 162.480 ;
        RECT 81.480 162.420 81.800 162.480 ;
        RECT 90.680 162.420 91.000 162.480 ;
        RECT 105.950 162.480 113.540 162.620 ;
        RECT 44.695 162.280 44.985 162.325 ;
        RECT 92.075 162.280 92.365 162.325 ;
        RECT 92.520 162.280 92.840 162.340 ;
        RECT 95.740 162.280 96.060 162.340 ;
        RECT 24.070 162.140 30.040 162.280 ;
        RECT 44.310 162.140 44.985 162.280 ;
        RECT 23.535 161.755 23.825 161.985 ;
        RECT 24.070 161.645 24.210 162.140 ;
        RECT 29.900 162.000 30.040 162.140 ;
        RECT 44.695 162.095 44.985 162.140 ;
        RECT 45.230 162.140 46.290 162.280 ;
        RECT 26.740 161.940 27.060 162.000 ;
        RECT 29.900 161.985 30.280 162.000 ;
        RECT 29.055 161.940 29.345 161.985 ;
        RECT 26.740 161.800 29.345 161.940 ;
        RECT 26.740 161.740 27.060 161.800 ;
        RECT 29.055 161.755 29.345 161.800 ;
        RECT 29.825 161.940 30.280 161.985 ;
        RECT 39.160 161.940 39.480 162.000 ;
        RECT 29.825 161.800 39.480 161.940 ;
        RECT 29.825 161.755 30.280 161.800 ;
        RECT 23.995 161.415 24.285 161.645 ;
        RECT 25.375 161.600 25.665 161.645 ;
        RECT 27.200 161.600 27.520 161.660 ;
        RECT 25.375 161.460 27.520 161.600 ;
        RECT 29.130 161.600 29.270 161.755 ;
        RECT 29.960 161.740 30.280 161.755 ;
        RECT 39.160 161.740 39.480 161.800 ;
        RECT 39.620 161.740 39.940 162.000 ;
        RECT 42.395 161.940 42.685 161.985 ;
        RECT 43.300 161.940 43.620 162.000 ;
        RECT 42.395 161.800 43.620 161.940 ;
        RECT 42.395 161.755 42.685 161.800 ;
        RECT 43.300 161.740 43.620 161.800 ;
        RECT 43.760 161.940 44.080 162.000 ;
        RECT 45.230 161.940 45.370 162.140 ;
        RECT 43.760 161.800 45.370 161.940 ;
        RECT 43.760 161.740 44.080 161.800 ;
        RECT 45.600 161.740 45.920 162.000 ;
        RECT 46.150 161.985 46.290 162.140 ;
        RECT 87.090 162.140 96.060 162.280 ;
        RECT 46.075 161.940 46.365 161.985 ;
        RECT 51.135 161.940 51.425 161.985 ;
        RECT 52.500 161.940 52.820 162.000 ;
        RECT 66.760 161.985 67.080 162.000 ;
        RECT 46.075 161.800 52.820 161.940 ;
        RECT 46.075 161.755 46.365 161.800 ;
        RECT 51.135 161.755 51.425 161.800 ;
        RECT 52.500 161.740 52.820 161.800 ;
        RECT 66.730 161.755 67.080 161.985 ;
        RECT 66.760 161.740 67.080 161.755 ;
        RECT 72.280 161.940 72.600 162.000 ;
        RECT 75.515 161.940 75.805 161.985 ;
        RECT 72.280 161.800 75.805 161.940 ;
        RECT 72.280 161.740 72.600 161.800 ;
        RECT 75.515 161.755 75.805 161.800 ;
        RECT 83.895 161.940 84.185 161.985 ;
        RECT 85.160 161.940 85.480 162.000 ;
        RECT 87.090 161.940 87.230 162.140 ;
        RECT 92.075 162.095 92.365 162.140 ;
        RECT 92.520 162.080 92.840 162.140 ;
        RECT 95.740 162.080 96.060 162.140 ;
        RECT 98.975 162.280 99.265 162.325 ;
        RECT 99.880 162.280 100.200 162.340 ;
        RECT 98.975 162.140 100.200 162.280 ;
        RECT 98.975 162.095 99.265 162.140 ;
        RECT 99.880 162.080 100.200 162.140 ;
        RECT 103.575 162.280 103.865 162.325 ;
        RECT 104.940 162.280 105.260 162.340 ;
        RECT 103.575 162.140 105.260 162.280 ;
        RECT 103.575 162.095 103.865 162.140 ;
        RECT 104.940 162.080 105.260 162.140 ;
        RECT 83.895 161.800 84.930 161.940 ;
        RECT 83.895 161.755 84.185 161.800 ;
        RECT 38.700 161.600 39.020 161.660 ;
        RECT 39.710 161.600 39.850 161.740 ;
        RECT 29.130 161.460 39.850 161.600 ;
        RECT 42.855 161.600 43.145 161.645 ;
        RECT 47.440 161.600 47.760 161.660 ;
        RECT 42.855 161.460 47.760 161.600 ;
        RECT 25.375 161.415 25.665 161.460 ;
        RECT 27.200 161.400 27.520 161.460 ;
        RECT 38.700 161.400 39.020 161.460 ;
        RECT 42.855 161.415 43.145 161.460 ;
        RECT 47.440 161.400 47.760 161.460 ;
        RECT 50.200 161.600 50.520 161.660 ;
        RECT 50.675 161.600 50.965 161.645 ;
        RECT 50.200 161.460 50.965 161.600 ;
        RECT 50.200 161.400 50.520 161.460 ;
        RECT 50.675 161.415 50.965 161.460 ;
        RECT 62.620 161.600 62.940 161.660 ;
        RECT 65.395 161.600 65.685 161.645 ;
        RECT 62.620 161.460 65.685 161.600 ;
        RECT 62.620 161.400 62.940 161.460 ;
        RECT 65.395 161.415 65.685 161.460 ;
        RECT 66.275 161.600 66.565 161.645 ;
        RECT 67.465 161.600 67.755 161.645 ;
        RECT 69.985 161.600 70.275 161.645 ;
        RECT 66.275 161.460 70.275 161.600 ;
        RECT 66.275 161.415 66.565 161.460 ;
        RECT 67.465 161.415 67.755 161.460 ;
        RECT 69.985 161.415 70.275 161.460 ;
        RECT 80.585 161.600 80.875 161.645 ;
        RECT 83.105 161.600 83.395 161.645 ;
        RECT 84.295 161.600 84.585 161.645 ;
        RECT 80.585 161.460 84.585 161.600 ;
        RECT 84.790 161.600 84.930 161.800 ;
        RECT 85.160 161.800 87.230 161.940 ;
        RECT 85.160 161.740 85.480 161.800 ;
        RECT 87.475 161.755 87.765 161.985 ;
        RECT 84.790 161.460 85.850 161.600 ;
        RECT 80.585 161.415 80.875 161.460 ;
        RECT 83.105 161.415 83.395 161.460 ;
        RECT 84.295 161.415 84.585 161.460 ;
        RECT 37.320 161.260 37.640 161.320 ;
        RECT 85.710 161.305 85.850 161.460 ;
        RECT 46.995 161.260 47.285 161.305 ;
        RECT 37.320 161.120 47.285 161.260 ;
        RECT 37.320 161.060 37.640 161.120 ;
        RECT 46.995 161.075 47.285 161.120 ;
        RECT 65.880 161.260 66.170 161.305 ;
        RECT 67.980 161.260 68.270 161.305 ;
        RECT 69.550 161.260 69.840 161.305 ;
        RECT 72.755 161.260 73.045 161.305 ;
        RECT 65.880 161.120 69.840 161.260 ;
        RECT 65.880 161.075 66.170 161.120 ;
        RECT 67.980 161.075 68.270 161.120 ;
        RECT 69.550 161.075 69.840 161.120 ;
        RECT 71.450 161.120 73.045 161.260 ;
        RECT 40.095 160.920 40.385 160.965 ;
        RECT 40.540 160.920 40.860 160.980 ;
        RECT 41.920 160.920 42.240 160.980 ;
        RECT 40.095 160.780 42.240 160.920 ;
        RECT 40.095 160.735 40.385 160.780 ;
        RECT 40.540 160.720 40.860 160.780 ;
        RECT 41.920 160.720 42.240 160.780 ;
        RECT 46.060 160.720 46.380 160.980 ;
        RECT 69.060 160.920 69.380 160.980 ;
        RECT 71.450 160.920 71.590 161.120 ;
        RECT 72.755 161.075 73.045 161.120 ;
        RECT 81.020 161.260 81.310 161.305 ;
        RECT 82.590 161.260 82.880 161.305 ;
        RECT 84.690 161.260 84.980 161.305 ;
        RECT 81.020 161.120 84.980 161.260 ;
        RECT 81.020 161.075 81.310 161.120 ;
        RECT 82.590 161.075 82.880 161.120 ;
        RECT 84.690 161.075 84.980 161.120 ;
        RECT 85.635 161.075 85.925 161.305 ;
        RECT 87.550 161.260 87.690 161.755 ;
        RECT 87.920 161.740 88.240 162.000 ;
        RECT 97.120 161.940 97.440 162.000 ;
        RECT 103.115 161.940 103.405 161.985 ;
        RECT 105.415 161.940 105.705 161.985 ;
        RECT 97.120 161.800 100.110 161.940 ;
        RECT 97.120 161.740 97.440 161.800 ;
        RECT 88.380 161.400 88.700 161.660 ;
        RECT 99.420 161.400 99.740 161.660 ;
        RECT 99.970 161.645 100.110 161.800 ;
        RECT 103.115 161.800 105.705 161.940 ;
        RECT 103.115 161.755 103.405 161.800 ;
        RECT 105.415 161.755 105.705 161.800 ;
        RECT 99.895 161.415 100.185 161.645 ;
        RECT 104.035 161.600 104.325 161.645 ;
        RECT 105.950 161.600 106.090 162.480 ;
        RECT 113.220 162.420 113.540 162.480 ;
        RECT 114.600 162.620 114.920 162.680 ;
        RECT 118.280 162.620 118.600 162.680 ;
        RECT 114.600 162.480 118.600 162.620 ;
        RECT 114.600 162.420 114.920 162.480 ;
        RECT 118.280 162.420 118.600 162.480 ;
        RECT 118.755 162.620 119.045 162.665 ;
        RECT 119.660 162.620 119.980 162.680 ;
        RECT 118.755 162.480 119.980 162.620 ;
        RECT 118.755 162.435 119.045 162.480 ;
        RECT 119.660 162.420 119.980 162.480 ;
        RECT 133.460 162.420 133.780 162.680 ;
        RECT 134.855 162.620 135.145 162.665 ;
        RECT 135.760 162.620 136.080 162.680 ;
        RECT 134.855 162.480 136.080 162.620 ;
        RECT 134.855 162.435 135.145 162.480 ;
        RECT 135.760 162.420 136.080 162.480 ;
        RECT 106.320 162.280 106.640 162.340 ;
        RECT 110.015 162.280 110.305 162.325 ;
        RECT 106.320 162.140 110.305 162.280 ;
        RECT 106.320 162.080 106.640 162.140 ;
        RECT 110.015 162.095 110.305 162.140 ;
        RECT 110.475 162.280 110.765 162.325 ;
        RECT 110.475 162.140 114.830 162.280 ;
        RECT 110.475 162.095 110.765 162.140 ;
        RECT 109.080 161.740 109.400 162.000 ;
        RECT 110.920 161.740 111.240 162.000 ;
        RECT 111.380 161.940 111.700 162.000 ;
        RECT 112.300 161.940 112.620 162.000 ;
        RECT 113.695 161.940 113.985 161.985 ;
        RECT 111.380 161.800 113.985 161.940 ;
        RECT 111.380 161.740 111.700 161.800 ;
        RECT 112.300 161.740 112.620 161.800 ;
        RECT 113.695 161.755 113.985 161.800 ;
        RECT 114.140 161.940 114.460 162.000 ;
        RECT 114.690 161.940 114.830 162.140 ;
        RECT 119.200 162.080 119.520 162.340 ;
        RECT 114.140 161.800 114.830 161.940 ;
        RECT 115.980 161.940 116.300 162.000 ;
        RECT 116.915 161.940 117.205 161.985 ;
        RECT 115.980 161.800 117.205 161.940 ;
        RECT 114.140 161.740 114.460 161.800 ;
        RECT 115.980 161.740 116.300 161.800 ;
        RECT 116.915 161.755 117.205 161.800 ;
        RECT 117.820 161.740 118.140 162.000 ;
        RECT 124.260 161.740 124.580 162.000 ;
        RECT 125.195 161.755 125.485 161.985 ;
        RECT 104.035 161.460 106.090 161.600 ;
        RECT 104.035 161.415 104.325 161.460 ;
        RECT 108.175 161.415 108.465 161.645 ;
        RECT 97.135 161.260 97.425 161.305 ;
        RECT 87.550 161.120 97.425 161.260 ;
        RECT 97.135 161.075 97.425 161.120 ;
        RECT 100.340 161.260 100.660 161.320 ;
        RECT 108.250 161.260 108.390 161.415 ;
        RECT 113.220 161.400 113.540 161.660 ;
        RECT 114.600 161.400 114.920 161.660 ;
        RECT 122.880 161.400 123.200 161.660 ;
        RECT 100.340 161.120 108.390 161.260 ;
        RECT 110.460 161.260 110.780 161.320 ;
        RECT 118.740 161.260 119.060 161.320 ;
        RECT 125.270 161.260 125.410 161.755 ;
        RECT 126.560 161.740 126.880 162.000 ;
        RECT 127.940 161.985 128.260 162.000 ;
        RECT 127.910 161.940 128.260 161.985 ;
        RECT 127.745 161.800 128.260 161.940 ;
        RECT 133.550 161.940 133.690 162.420 ;
        RECT 133.935 161.940 134.225 161.985 ;
        RECT 133.550 161.800 134.225 161.940 ;
        RECT 127.910 161.755 128.260 161.800 ;
        RECT 133.935 161.755 134.225 161.800 ;
        RECT 135.775 161.755 136.065 161.985 ;
        RECT 127.940 161.740 128.260 161.755 ;
        RECT 127.455 161.600 127.745 161.645 ;
        RECT 128.645 161.600 128.935 161.645 ;
        RECT 131.165 161.600 131.455 161.645 ;
        RECT 127.455 161.460 131.455 161.600 ;
        RECT 127.455 161.415 127.745 161.460 ;
        RECT 128.645 161.415 128.935 161.460 ;
        RECT 131.165 161.415 131.455 161.460 ;
        RECT 131.620 161.600 131.940 161.660 ;
        RECT 135.850 161.600 135.990 161.755 ;
        RECT 131.620 161.460 135.990 161.600 ;
        RECT 131.620 161.400 131.940 161.460 ;
        RECT 110.460 161.120 125.410 161.260 ;
        RECT 127.060 161.260 127.350 161.305 ;
        RECT 129.160 161.260 129.450 161.305 ;
        RECT 130.730 161.260 131.020 161.305 ;
        RECT 127.060 161.120 131.020 161.260 ;
        RECT 100.340 161.060 100.660 161.120 ;
        RECT 110.460 161.060 110.780 161.120 ;
        RECT 118.740 161.060 119.060 161.120 ;
        RECT 127.060 161.075 127.350 161.120 ;
        RECT 129.160 161.075 129.450 161.120 ;
        RECT 130.730 161.075 131.020 161.120 ;
        RECT 136.680 161.060 137.000 161.320 ;
        RECT 69.060 160.780 71.590 160.920 ;
        RECT 69.060 160.720 69.380 160.780 ;
        RECT 72.280 160.720 72.600 160.980 ;
        RECT 78.275 160.920 78.565 160.965 ;
        RECT 80.560 160.920 80.880 160.980 ;
        RECT 78.275 160.780 80.880 160.920 ;
        RECT 78.275 160.735 78.565 160.780 ;
        RECT 80.560 160.720 80.880 160.780 ;
        RECT 101.260 160.720 101.580 160.980 ;
        RECT 111.840 160.720 112.160 160.980 ;
        RECT 112.300 160.720 112.620 160.980 ;
        RECT 116.900 160.920 117.220 160.980 ;
        RECT 117.835 160.920 118.125 160.965 ;
        RECT 120.120 160.920 120.440 160.980 ;
        RECT 124.260 160.920 124.580 160.980 ;
        RECT 116.900 160.780 124.580 160.920 ;
        RECT 116.900 160.720 117.220 160.780 ;
        RECT 117.835 160.735 118.125 160.780 ;
        RECT 120.120 160.720 120.440 160.780 ;
        RECT 124.260 160.720 124.580 160.780 ;
        RECT 125.640 160.920 125.960 160.980 ;
        RECT 126.115 160.920 126.405 160.965 ;
        RECT 125.640 160.780 126.405 160.920 ;
        RECT 125.640 160.720 125.960 160.780 ;
        RECT 126.115 160.735 126.405 160.780 ;
        RECT 13.330 160.100 138.910 160.580 ;
        RECT 66.760 159.700 67.080 159.960 ;
        RECT 87.460 159.900 87.780 159.960 ;
        RECT 88.855 159.900 89.145 159.945 ;
        RECT 87.460 159.760 89.145 159.900 ;
        RECT 87.460 159.700 87.780 159.760 ;
        RECT 88.855 159.715 89.145 159.760 ;
        RECT 99.435 159.900 99.725 159.945 ;
        RECT 100.340 159.900 100.660 159.960 ;
        RECT 99.435 159.760 100.660 159.900 ;
        RECT 99.435 159.715 99.725 159.760 ;
        RECT 100.340 159.700 100.660 159.760 ;
        RECT 107.255 159.900 107.545 159.945 ;
        RECT 109.080 159.900 109.400 159.960 ;
        RECT 107.255 159.760 109.400 159.900 ;
        RECT 107.255 159.715 107.545 159.760 ;
        RECT 109.080 159.700 109.400 159.760 ;
        RECT 35.940 159.560 36.260 159.620 ;
        RECT 41.000 159.560 41.320 159.620 ;
        RECT 35.940 159.420 41.320 159.560 ;
        RECT 35.940 159.360 36.260 159.420 ;
        RECT 41.000 159.360 41.320 159.420 ;
        RECT 93.020 159.560 93.310 159.605 ;
        RECT 95.120 159.560 95.410 159.605 ;
        RECT 96.690 159.560 96.980 159.605 ;
        RECT 93.020 159.420 96.980 159.560 ;
        RECT 93.020 159.375 93.310 159.420 ;
        RECT 95.120 159.375 95.410 159.420 ;
        RECT 96.690 159.375 96.980 159.420 ;
        RECT 118.280 159.560 118.600 159.620 ;
        RECT 130.280 159.560 130.570 159.605 ;
        RECT 132.380 159.560 132.670 159.605 ;
        RECT 133.950 159.560 134.240 159.605 ;
        RECT 118.280 159.420 125.870 159.560 ;
        RECT 118.280 159.360 118.600 159.420 ;
        RECT 35.035 159.220 35.325 159.265 ;
        RECT 40.095 159.220 40.385 159.265 ;
        RECT 35.035 159.080 40.385 159.220 ;
        RECT 35.035 159.035 35.325 159.080 ;
        RECT 40.095 159.035 40.385 159.080 ;
        RECT 69.060 159.020 69.380 159.280 ;
        RECT 69.535 159.035 69.825 159.265 ;
        RECT 69.980 159.220 70.300 159.280 ;
        RECT 75.055 159.220 75.345 159.265 ;
        RECT 69.980 159.080 75.345 159.220 ;
        RECT 38.700 158.680 39.020 158.940 ;
        RECT 39.620 158.680 39.940 158.940 ;
        RECT 69.610 158.880 69.750 159.035 ;
        RECT 69.980 159.020 70.300 159.080 ;
        RECT 75.055 159.035 75.345 159.080 ;
        RECT 75.960 159.220 76.280 159.280 ;
        RECT 83.780 159.220 84.100 159.280 ;
        RECT 75.960 159.080 84.100 159.220 ;
        RECT 75.960 159.020 76.280 159.080 ;
        RECT 83.780 159.020 84.100 159.080 ;
        RECT 84.240 159.220 84.560 159.280 ;
        RECT 85.635 159.220 85.925 159.265 ;
        RECT 84.240 159.080 85.925 159.220 ;
        RECT 84.240 159.020 84.560 159.080 ;
        RECT 85.635 159.035 85.925 159.080 ;
        RECT 86.555 159.220 86.845 159.265 ;
        RECT 92.060 159.220 92.380 159.280 ;
        RECT 86.555 159.080 92.380 159.220 ;
        RECT 86.555 159.035 86.845 159.080 ;
        RECT 92.060 159.020 92.380 159.080 ;
        RECT 92.520 159.020 92.840 159.280 ;
        RECT 93.415 159.220 93.705 159.265 ;
        RECT 94.605 159.220 94.895 159.265 ;
        RECT 97.125 159.220 97.415 159.265 ;
        RECT 93.415 159.080 97.415 159.220 ;
        RECT 93.415 159.035 93.705 159.080 ;
        RECT 94.605 159.035 94.895 159.080 ;
        RECT 97.125 159.035 97.415 159.080 ;
        RECT 99.420 159.220 99.740 159.280 ;
        RECT 104.035 159.220 104.325 159.265 ;
        RECT 99.420 159.080 104.325 159.220 ;
        RECT 99.420 159.020 99.740 159.080 ;
        RECT 104.035 159.035 104.325 159.080 ;
        RECT 109.095 159.220 109.385 159.265 ;
        RECT 112.300 159.220 112.620 159.280 ;
        RECT 125.730 159.265 125.870 159.420 ;
        RECT 130.280 159.420 134.240 159.560 ;
        RECT 130.280 159.375 130.570 159.420 ;
        RECT 132.380 159.375 132.670 159.420 ;
        RECT 133.950 159.375 134.240 159.420 ;
        RECT 109.095 159.080 112.620 159.220 ;
        RECT 109.095 159.035 109.385 159.080 ;
        RECT 112.300 159.020 112.620 159.080 ;
        RECT 116.070 159.080 117.590 159.220 ;
        RECT 76.050 158.880 76.190 159.020 ;
        RECT 69.610 158.740 76.190 158.880 ;
        RECT 93.870 158.880 94.160 158.925 ;
        RECT 101.260 158.880 101.580 158.940 ;
        RECT 93.870 158.740 101.580 158.880 ;
        RECT 93.870 158.695 94.160 158.740 ;
        RECT 101.260 158.680 101.580 158.740 ;
        RECT 107.700 158.680 108.020 158.940 ;
        RECT 108.175 158.880 108.465 158.925 ;
        RECT 109.540 158.880 109.860 158.940 ;
        RECT 108.175 158.740 109.860 158.880 ;
        RECT 108.175 158.695 108.465 158.740 ;
        RECT 109.540 158.680 109.860 158.740 ;
        RECT 110.460 158.680 110.780 158.940 ;
        RECT 111.855 158.695 112.145 158.925 ;
        RECT 115.075 158.880 115.365 158.925 ;
        RECT 116.070 158.880 116.210 159.080 ;
        RECT 115.075 158.740 116.210 158.880 ;
        RECT 115.075 158.695 115.365 158.740 ;
        RECT 116.455 158.695 116.745 158.925 ;
        RECT 68.615 158.540 68.905 158.585 ;
        RECT 72.740 158.540 73.060 158.600 ;
        RECT 103.560 158.540 103.880 158.600 ;
        RECT 68.615 158.400 69.980 158.540 ;
        RECT 68.615 158.355 68.905 158.400 ;
        RECT 15.700 158.200 16.020 158.260 ;
        RECT 65.840 158.200 66.160 158.260 ;
        RECT 15.700 158.060 66.160 158.200 ;
        RECT 69.840 158.200 69.980 158.400 ;
        RECT 72.740 158.400 103.880 158.540 ;
        RECT 72.740 158.340 73.060 158.400 ;
        RECT 103.560 158.340 103.880 158.400 ;
        RECT 106.320 158.540 106.640 158.600 ;
        RECT 109.095 158.540 109.385 158.585 ;
        RECT 106.320 158.400 109.385 158.540 ;
        RECT 111.930 158.540 112.070 158.695 ;
        RECT 112.300 158.540 112.620 158.600 ;
        RECT 111.930 158.400 112.620 158.540 ;
        RECT 106.320 158.340 106.640 158.400 ;
        RECT 109.095 158.355 109.385 158.400 ;
        RECT 112.300 158.340 112.620 158.400 ;
        RECT 114.140 158.540 114.460 158.600 ;
        RECT 116.530 158.540 116.670 158.695 ;
        RECT 116.900 158.680 117.220 158.940 ;
        RECT 117.450 158.880 117.590 159.080 ;
        RECT 125.655 159.035 125.945 159.265 ;
        RECT 130.675 159.220 130.965 159.265 ;
        RECT 131.865 159.220 132.155 159.265 ;
        RECT 134.385 159.220 134.675 159.265 ;
        RECT 130.675 159.080 134.675 159.220 ;
        RECT 130.675 159.035 130.965 159.080 ;
        RECT 131.865 159.035 132.155 159.080 ;
        RECT 134.385 159.035 134.675 159.080 ;
        RECT 118.295 158.880 118.585 158.925 ;
        RECT 122.880 158.880 123.200 158.940 ;
        RECT 129.795 158.880 130.085 158.925 ;
        RECT 117.450 158.740 118.585 158.880 ;
        RECT 118.295 158.695 118.585 158.740 ;
        RECT 119.290 158.740 130.085 158.880 ;
        RECT 114.140 158.400 116.670 158.540 ;
        RECT 114.140 158.340 114.460 158.400 ;
        RECT 117.360 158.340 117.680 158.600 ;
        RECT 119.290 158.585 119.430 158.740 ;
        RECT 122.880 158.680 123.200 158.740 ;
        RECT 129.795 158.695 130.085 158.740 ;
        RECT 119.215 158.355 119.505 158.585 ;
        RECT 131.020 158.540 131.310 158.585 ;
        RECT 128.950 158.400 131.310 158.540 ;
        RECT 71.820 158.200 72.140 158.260 ;
        RECT 69.840 158.060 72.140 158.200 ;
        RECT 15.700 158.000 16.020 158.060 ;
        RECT 65.840 158.000 66.160 158.060 ;
        RECT 71.820 158.000 72.140 158.060 ;
        RECT 72.280 158.000 72.600 158.260 ;
        RECT 87.000 158.000 87.320 158.260 ;
        RECT 110.475 158.200 110.765 158.245 ;
        RECT 113.220 158.200 113.540 158.260 ;
        RECT 110.475 158.060 113.540 158.200 ;
        RECT 110.475 158.015 110.765 158.060 ;
        RECT 113.220 158.000 113.540 158.060 ;
        RECT 115.520 158.000 115.840 158.260 ;
        RECT 116.440 158.200 116.760 158.260 ;
        RECT 119.290 158.200 119.430 158.355 ;
        RECT 116.440 158.060 119.430 158.200 ;
        RECT 116.440 158.000 116.760 158.060 ;
        RECT 126.560 158.000 126.880 158.260 ;
        RECT 127.020 158.000 127.340 158.260 ;
        RECT 128.950 158.245 129.090 158.400 ;
        RECT 131.020 158.355 131.310 158.400 ;
        RECT 128.875 158.015 129.165 158.245 ;
        RECT 135.300 158.200 135.620 158.260 ;
        RECT 136.695 158.200 136.985 158.245 ;
        RECT 135.300 158.060 136.985 158.200 ;
        RECT 135.300 158.000 135.620 158.060 ;
        RECT 136.695 158.015 136.985 158.060 ;
        RECT 13.330 157.380 138.910 157.860 ;
        RECT 15.700 156.980 16.020 157.240 ;
        RECT 29.975 157.180 30.265 157.225 ;
        RECT 30.880 157.180 31.200 157.240 ;
        RECT 29.975 157.040 31.200 157.180 ;
        RECT 29.975 156.995 30.265 157.040 ;
        RECT 30.880 156.980 31.200 157.040 ;
        RECT 36.860 157.180 37.180 157.240 ;
        RECT 38.255 157.180 38.545 157.225 ;
        RECT 36.860 157.040 38.545 157.180 ;
        RECT 36.860 156.980 37.180 157.040 ;
        RECT 38.255 156.995 38.545 157.040 ;
        RECT 69.980 157.180 70.300 157.240 ;
        RECT 72.295 157.180 72.585 157.225 ;
        RECT 69.980 157.040 72.585 157.180 ;
        RECT 69.980 156.980 70.300 157.040 ;
        RECT 72.295 156.995 72.585 157.040 ;
        RECT 99.420 156.980 99.740 157.240 ;
        RECT 111.840 157.180 112.160 157.240 ;
        RECT 102.730 157.040 112.160 157.180 ;
        RECT 16.620 156.840 16.940 156.900 ;
        RECT 35.480 156.840 35.800 156.900 ;
        RECT 35.955 156.840 36.245 156.885 ;
        RECT 38.700 156.840 39.020 156.900 ;
        RECT 40.555 156.840 40.845 156.885 ;
        RECT 16.620 156.700 35.250 156.840 ;
        RECT 16.620 156.640 16.940 156.700 ;
        RECT 12.020 156.500 12.340 156.560 ;
        RECT 14.795 156.500 15.085 156.545 ;
        RECT 12.020 156.360 15.085 156.500 ;
        RECT 12.020 156.300 12.340 156.360 ;
        RECT 14.795 156.315 15.085 156.360 ;
        RECT 19.380 156.300 19.700 156.560 ;
        RECT 19.840 156.500 20.160 156.560 ;
        RECT 20.675 156.500 20.965 156.545 ;
        RECT 19.840 156.360 20.965 156.500 ;
        RECT 19.840 156.300 20.160 156.360 ;
        RECT 20.675 156.315 20.965 156.360 ;
        RECT 27.200 156.500 27.520 156.560 ;
        RECT 27.675 156.500 27.965 156.545 ;
        RECT 27.200 156.360 27.965 156.500 ;
        RECT 27.200 156.300 27.520 156.360 ;
        RECT 27.675 156.315 27.965 156.360 ;
        RECT 30.270 156.500 30.560 156.545 ;
        RECT 31.800 156.500 32.120 156.560 ;
        RECT 30.270 156.360 32.120 156.500 ;
        RECT 30.270 156.315 30.560 156.360 ;
        RECT 31.800 156.300 32.120 156.360 ;
        RECT 20.275 156.160 20.565 156.205 ;
        RECT 21.465 156.160 21.755 156.205 ;
        RECT 23.985 156.160 24.275 156.205 ;
        RECT 20.275 156.020 24.275 156.160 ;
        RECT 20.275 155.975 20.565 156.020 ;
        RECT 21.465 155.975 21.755 156.020 ;
        RECT 23.985 155.975 24.275 156.020 ;
        RECT 19.880 155.820 20.170 155.865 ;
        RECT 21.980 155.820 22.270 155.865 ;
        RECT 23.550 155.820 23.840 155.865 ;
        RECT 19.880 155.680 23.840 155.820 ;
        RECT 19.880 155.635 20.170 155.680 ;
        RECT 21.980 155.635 22.270 155.680 ;
        RECT 23.550 155.635 23.840 155.680 ;
        RECT 26.295 155.480 26.585 155.525 ;
        RECT 28.120 155.480 28.440 155.540 ;
        RECT 26.295 155.340 28.440 155.480 ;
        RECT 26.295 155.295 26.585 155.340 ;
        RECT 28.120 155.280 28.440 155.340 ;
        RECT 30.895 155.480 31.185 155.525 ;
        RECT 31.340 155.480 31.660 155.540 ;
        RECT 30.895 155.340 31.660 155.480 ;
        RECT 35.110 155.480 35.250 156.700 ;
        RECT 35.480 156.700 40.845 156.840 ;
        RECT 35.480 156.640 35.800 156.700 ;
        RECT 35.955 156.655 36.245 156.700 ;
        RECT 38.700 156.640 39.020 156.700 ;
        RECT 40.555 156.655 40.845 156.700 ;
        RECT 66.300 156.840 66.620 156.900 ;
        RECT 93.870 156.840 94.160 156.885 ;
        RECT 102.730 156.840 102.870 157.040 ;
        RECT 111.840 156.980 112.160 157.040 ;
        RECT 121.975 157.180 122.265 157.225 ;
        RECT 126.560 157.180 126.880 157.240 ;
        RECT 121.975 157.040 126.880 157.180 ;
        RECT 121.975 156.995 122.265 157.040 ;
        RECT 126.560 156.980 126.880 157.040 ;
        RECT 127.020 157.180 127.340 157.240 ;
        RECT 132.095 157.180 132.385 157.225 ;
        RECT 127.020 157.040 132.385 157.180 ;
        RECT 127.020 156.980 127.340 157.040 ;
        RECT 132.095 156.995 132.385 157.040 ;
        RECT 120.135 156.840 120.425 156.885 ;
        RECT 122.880 156.840 123.200 156.900 ;
        RECT 123.355 156.840 123.645 156.885 ;
        RECT 66.300 156.700 79.870 156.840 ;
        RECT 66.300 156.640 66.620 156.700 ;
        RECT 39.620 156.500 39.940 156.560 ;
        RECT 37.410 156.360 39.940 156.500 ;
        RECT 37.410 155.880 37.550 156.360 ;
        RECT 39.620 156.300 39.940 156.360 ;
        RECT 66.730 156.500 67.020 156.545 ;
        RECT 68.140 156.500 68.460 156.560 ;
        RECT 66.730 156.360 68.460 156.500 ;
        RECT 66.730 156.315 67.020 156.360 ;
        RECT 68.140 156.300 68.460 156.360 ;
        RECT 74.580 156.300 74.900 156.560 ;
        RECT 79.730 156.545 79.870 156.700 ;
        RECT 93.870 156.700 102.870 156.840 ;
        RECT 107.790 156.700 116.210 156.840 ;
        RECT 93.870 156.655 94.160 156.700 ;
        RECT 75.055 156.500 75.345 156.545 ;
        RECT 76.895 156.500 77.185 156.545 ;
        RECT 75.055 156.360 77.185 156.500 ;
        RECT 75.055 156.315 75.345 156.360 ;
        RECT 76.895 156.315 77.185 156.360 ;
        RECT 79.655 156.315 79.945 156.545 ;
        RECT 92.520 156.300 92.840 156.560 ;
        RECT 106.320 156.545 106.640 156.560 ;
        RECT 107.790 156.545 107.930 156.700 ;
        RECT 106.320 156.500 106.670 156.545 ;
        RECT 106.320 156.360 106.835 156.500 ;
        RECT 106.320 156.315 106.670 156.360 ;
        RECT 107.715 156.315 108.005 156.545 ;
        RECT 112.300 156.500 112.620 156.560 ;
        RECT 109.170 156.360 112.620 156.500 ;
        RECT 106.320 156.300 106.640 156.315 ;
        RECT 62.620 156.160 62.940 156.220 ;
        RECT 65.395 156.160 65.685 156.205 ;
        RECT 62.620 156.020 65.685 156.160 ;
        RECT 62.620 155.960 62.940 156.020 ;
        RECT 65.395 155.975 65.685 156.020 ;
        RECT 66.275 156.160 66.565 156.205 ;
        RECT 67.465 156.160 67.755 156.205 ;
        RECT 69.985 156.160 70.275 156.205 ;
        RECT 66.275 156.020 70.275 156.160 ;
        RECT 66.275 155.975 66.565 156.020 ;
        RECT 67.465 155.975 67.755 156.020 ;
        RECT 69.985 155.975 70.275 156.020 ;
        RECT 75.960 155.960 76.280 156.220 ;
        RECT 93.415 156.160 93.705 156.205 ;
        RECT 94.605 156.160 94.895 156.205 ;
        RECT 97.125 156.160 97.415 156.205 ;
        RECT 93.415 156.020 97.415 156.160 ;
        RECT 93.415 155.975 93.705 156.020 ;
        RECT 94.605 155.975 94.895 156.020 ;
        RECT 97.125 155.975 97.415 156.020 ;
        RECT 103.125 156.160 103.415 156.205 ;
        RECT 105.645 156.160 105.935 156.205 ;
        RECT 106.835 156.160 107.125 156.205 ;
        RECT 103.125 156.020 107.125 156.160 ;
        RECT 103.125 155.975 103.415 156.020 ;
        RECT 105.645 155.975 105.935 156.020 ;
        RECT 106.835 155.975 107.125 156.020 ;
        RECT 37.320 155.620 37.640 155.880 ;
        RECT 65.880 155.820 66.170 155.865 ;
        RECT 67.980 155.820 68.270 155.865 ;
        RECT 69.550 155.820 69.840 155.865 ;
        RECT 72.755 155.820 73.045 155.865 ;
        RECT 40.170 155.680 65.610 155.820 ;
        RECT 40.170 155.480 40.310 155.680 ;
        RECT 35.110 155.340 40.310 155.480 ;
        RECT 40.540 155.480 40.860 155.540 ;
        RECT 41.475 155.480 41.765 155.525 ;
        RECT 40.540 155.340 41.765 155.480 ;
        RECT 65.470 155.480 65.610 155.680 ;
        RECT 65.880 155.680 69.840 155.820 ;
        RECT 65.880 155.635 66.170 155.680 ;
        RECT 67.980 155.635 68.270 155.680 ;
        RECT 69.550 155.635 69.840 155.680 ;
        RECT 71.450 155.680 73.045 155.820 ;
        RECT 66.760 155.480 67.080 155.540 ;
        RECT 65.470 155.340 67.080 155.480 ;
        RECT 30.895 155.295 31.185 155.340 ;
        RECT 31.340 155.280 31.660 155.340 ;
        RECT 40.540 155.280 40.860 155.340 ;
        RECT 41.475 155.295 41.765 155.340 ;
        RECT 66.760 155.280 67.080 155.340 ;
        RECT 69.060 155.480 69.380 155.540 ;
        RECT 71.450 155.480 71.590 155.680 ;
        RECT 72.755 155.635 73.045 155.680 ;
        RECT 93.020 155.820 93.310 155.865 ;
        RECT 95.120 155.820 95.410 155.865 ;
        RECT 96.690 155.820 96.980 155.865 ;
        RECT 93.020 155.680 96.980 155.820 ;
        RECT 93.020 155.635 93.310 155.680 ;
        RECT 95.120 155.635 95.410 155.680 ;
        RECT 96.690 155.635 96.980 155.680 ;
        RECT 103.560 155.820 103.850 155.865 ;
        RECT 105.130 155.820 105.420 155.865 ;
        RECT 107.230 155.820 107.520 155.865 ;
        RECT 103.560 155.680 107.520 155.820 ;
        RECT 103.560 155.635 103.850 155.680 ;
        RECT 105.130 155.635 105.420 155.680 ;
        RECT 107.230 155.635 107.520 155.680 ;
        RECT 109.170 155.540 109.310 156.360 ;
        RECT 112.300 156.300 112.620 156.360 ;
        RECT 114.715 156.500 115.005 156.545 ;
        RECT 115.520 156.500 115.840 156.560 ;
        RECT 114.715 156.360 115.840 156.500 ;
        RECT 114.715 156.315 115.005 156.360 ;
        RECT 115.520 156.300 115.840 156.360 ;
        RECT 116.070 156.205 116.210 156.700 ;
        RECT 120.135 156.700 126.790 156.840 ;
        RECT 120.135 156.655 120.425 156.700 ;
        RECT 122.880 156.640 123.200 156.700 ;
        RECT 123.355 156.655 123.645 156.700 ;
        RECT 116.915 156.315 117.205 156.545 ;
        RECT 111.405 156.160 111.695 156.205 ;
        RECT 113.925 156.160 114.215 156.205 ;
        RECT 115.115 156.160 115.405 156.205 ;
        RECT 111.405 156.020 115.405 156.160 ;
        RECT 111.405 155.975 111.695 156.020 ;
        RECT 113.925 155.975 114.215 156.020 ;
        RECT 115.115 155.975 115.405 156.020 ;
        RECT 115.995 156.160 116.285 156.205 ;
        RECT 116.440 156.160 116.760 156.220 ;
        RECT 115.995 156.020 116.760 156.160 ;
        RECT 115.995 155.975 116.285 156.020 ;
        RECT 116.440 155.960 116.760 156.020 ;
        RECT 111.840 155.820 112.130 155.865 ;
        RECT 113.410 155.820 113.700 155.865 ;
        RECT 115.510 155.820 115.800 155.865 ;
        RECT 111.840 155.680 115.800 155.820 ;
        RECT 111.840 155.635 112.130 155.680 ;
        RECT 113.410 155.635 113.700 155.680 ;
        RECT 115.510 155.635 115.800 155.680 ;
        RECT 69.060 155.340 71.590 155.480 ;
        RECT 84.240 155.480 84.560 155.540 ;
        RECT 97.120 155.480 97.440 155.540 ;
        RECT 84.240 155.340 97.440 155.480 ;
        RECT 69.060 155.280 69.380 155.340 ;
        RECT 84.240 155.280 84.560 155.340 ;
        RECT 97.120 155.280 97.440 155.340 ;
        RECT 100.815 155.480 101.105 155.525 ;
        RECT 101.260 155.480 101.580 155.540 ;
        RECT 100.815 155.340 101.580 155.480 ;
        RECT 100.815 155.295 101.105 155.340 ;
        RECT 101.260 155.280 101.580 155.340 ;
        RECT 109.080 155.280 109.400 155.540 ;
        RECT 109.540 155.480 109.860 155.540 ;
        RECT 116.990 155.480 117.130 156.315 ;
        RECT 117.820 156.300 118.140 156.560 ;
        RECT 118.280 156.500 118.600 156.560 ;
        RECT 119.215 156.500 119.505 156.545 ;
        RECT 118.280 156.360 119.505 156.500 ;
        RECT 118.280 156.300 118.600 156.360 ;
        RECT 119.215 156.315 119.505 156.360 ;
        RECT 120.580 156.300 120.900 156.560 ;
        RECT 121.040 156.300 121.360 156.560 ;
        RECT 122.435 156.315 122.725 156.545 ;
        RECT 117.375 156.160 117.665 156.205 ;
        RECT 122.510 156.160 122.650 156.315 ;
        RECT 123.800 156.300 124.120 156.560 ;
        RECT 124.275 156.315 124.565 156.545 ;
        RECT 124.350 156.160 124.490 156.315 ;
        RECT 125.640 156.300 125.960 156.560 ;
        RECT 126.650 156.545 126.790 156.700 ;
        RECT 126.575 156.315 126.865 156.545 ;
        RECT 127.020 156.300 127.340 156.560 ;
        RECT 127.495 156.315 127.785 156.545 ;
        RECT 130.715 156.500 131.005 156.545 ;
        RECT 135.300 156.500 135.620 156.560 ;
        RECT 130.715 156.360 135.620 156.500 ;
        RECT 130.715 156.315 131.005 156.360 ;
        RECT 127.570 156.160 127.710 156.315 ;
        RECT 135.300 156.300 135.620 156.360 ;
        RECT 135.775 156.500 136.065 156.545 ;
        RECT 136.220 156.500 136.540 156.560 ;
        RECT 135.775 156.360 136.540 156.500 ;
        RECT 135.775 156.315 136.065 156.360 ;
        RECT 136.220 156.300 136.540 156.360 ;
        RECT 117.375 156.020 122.650 156.160 ;
        RECT 123.890 156.020 127.710 156.160 ;
        RECT 117.375 155.975 117.665 156.020 ;
        RECT 121.040 155.820 121.360 155.880 ;
        RECT 123.340 155.820 123.660 155.880 ;
        RECT 123.890 155.820 124.030 156.020 ;
        RECT 121.040 155.680 124.030 155.820 ;
        RECT 128.415 155.820 128.705 155.865 ;
        RECT 130.240 155.820 130.560 155.880 ;
        RECT 128.415 155.680 130.560 155.820 ;
        RECT 121.040 155.620 121.360 155.680 ;
        RECT 123.340 155.620 123.660 155.680 ;
        RECT 128.415 155.635 128.705 155.680 ;
        RECT 130.240 155.620 130.560 155.680 ;
        RECT 131.620 155.620 131.940 155.880 ;
        RECT 109.540 155.340 117.130 155.480 ;
        RECT 125.195 155.480 125.485 155.525 ;
        RECT 130.700 155.480 131.020 155.540 ;
        RECT 125.195 155.340 131.020 155.480 ;
        RECT 109.540 155.280 109.860 155.340 ;
        RECT 125.195 155.295 125.485 155.340 ;
        RECT 130.700 155.280 131.020 155.340 ;
        RECT 136.680 155.280 137.000 155.540 ;
        RECT 13.330 154.660 138.910 155.140 ;
        RECT 15.715 154.460 16.005 154.505 ;
        RECT 16.620 154.460 16.940 154.520 ;
        RECT 15.715 154.320 16.940 154.460 ;
        RECT 15.715 154.275 16.005 154.320 ;
        RECT 16.620 154.260 16.940 154.320 ;
        RECT 19.840 154.260 20.160 154.520 ;
        RECT 20.760 154.260 21.080 154.520 ;
        RECT 41.460 154.460 41.780 154.520 ;
        RECT 42.395 154.460 42.685 154.505 ;
        RECT 41.460 154.320 42.685 154.460 ;
        RECT 41.460 154.260 41.780 154.320 ;
        RECT 42.395 154.275 42.685 154.320 ;
        RECT 62.635 154.460 62.925 154.505 ;
        RECT 66.300 154.460 66.620 154.520 ;
        RECT 62.635 154.320 66.620 154.460 ;
        RECT 62.635 154.275 62.925 154.320 ;
        RECT 66.300 154.260 66.620 154.320 ;
        RECT 68.140 154.460 68.460 154.520 ;
        RECT 69.995 154.460 70.285 154.505 ;
        RECT 68.140 154.320 70.285 154.460 ;
        RECT 68.140 154.260 68.460 154.320 ;
        RECT 69.995 154.275 70.285 154.320 ;
        RECT 74.580 154.460 74.900 154.520 ;
        RECT 98.975 154.460 99.265 154.505 ;
        RECT 74.580 154.320 99.265 154.460 ;
        RECT 74.580 154.260 74.900 154.320 ;
        RECT 98.975 154.275 99.265 154.320 ;
        RECT 108.635 154.460 108.925 154.505 ;
        RECT 114.600 154.460 114.920 154.520 ;
        RECT 108.635 154.320 114.920 154.460 ;
        RECT 108.635 154.275 108.925 154.320 ;
        RECT 114.600 154.260 114.920 154.320 ;
        RECT 119.215 154.460 119.505 154.505 ;
        RECT 126.560 154.460 126.880 154.520 ;
        RECT 119.215 154.320 126.880 154.460 ;
        RECT 119.215 154.275 119.505 154.320 ;
        RECT 126.560 154.260 126.880 154.320 ;
        RECT 136.695 154.460 136.985 154.505 ;
        RECT 138.060 154.460 138.380 154.520 ;
        RECT 136.695 154.320 138.380 154.460 ;
        RECT 136.695 154.275 136.985 154.320 ;
        RECT 138.060 154.260 138.380 154.320 ;
        RECT 65.380 154.120 65.670 154.165 ;
        RECT 66.950 154.120 67.240 154.165 ;
        RECT 69.050 154.120 69.340 154.165 ;
        RECT 65.380 153.980 69.340 154.120 ;
        RECT 65.380 153.935 65.670 153.980 ;
        RECT 66.950 153.935 67.240 153.980 ;
        RECT 69.050 153.935 69.340 153.980 ;
        RECT 71.820 154.120 72.140 154.180 ;
        RECT 94.835 154.120 95.125 154.165 ;
        RECT 100.340 154.120 100.660 154.180 ;
        RECT 71.820 153.980 95.125 154.120 ;
        RECT 71.820 153.920 72.140 153.980 ;
        RECT 94.835 153.935 95.125 153.980 ;
        RECT 97.210 153.980 100.660 154.120 ;
        RECT 23.980 153.780 24.300 153.840 ;
        RECT 21.540 153.640 24.300 153.780 ;
        RECT 18.475 153.255 18.765 153.485 ;
        RECT 19.395 153.440 19.685 153.485 ;
        RECT 21.540 153.440 21.680 153.640 ;
        RECT 23.980 153.580 24.300 153.640 ;
        RECT 24.440 153.780 24.760 153.840 ;
        RECT 37.320 153.780 37.640 153.840 ;
        RECT 64.945 153.780 65.235 153.825 ;
        RECT 67.465 153.780 67.755 153.825 ;
        RECT 68.655 153.780 68.945 153.825 ;
        RECT 24.440 153.640 29.730 153.780 ;
        RECT 24.440 153.580 24.760 153.640 ;
        RECT 19.395 153.300 21.680 153.440 ;
        RECT 19.395 153.255 19.685 153.300 ;
        RECT 15.240 152.900 15.560 153.160 ;
        RECT 18.550 152.760 18.690 153.255 ;
        RECT 22.140 153.240 22.460 153.500 ;
        RECT 23.075 153.440 23.365 153.485 ;
        RECT 25.820 153.440 26.140 153.500 ;
        RECT 23.075 153.300 26.140 153.440 ;
        RECT 23.075 153.255 23.365 153.300 ;
        RECT 25.820 153.240 26.140 153.300 ;
        RECT 28.120 153.240 28.440 153.500 ;
        RECT 18.935 153.100 19.225 153.145 ;
        RECT 20.615 153.100 20.905 153.145 ;
        RECT 18.935 152.960 20.905 153.100 ;
        RECT 18.935 152.915 19.225 152.960 ;
        RECT 20.615 152.915 20.905 152.960 ;
        RECT 21.220 153.100 21.540 153.160 ;
        RECT 21.695 153.100 21.985 153.145 ;
        RECT 21.220 152.960 21.985 153.100 ;
        RECT 21.220 152.900 21.540 152.960 ;
        RECT 21.695 152.915 21.985 152.960 ;
        RECT 24.440 152.900 24.760 153.160 ;
        RECT 25.375 153.100 25.665 153.145 ;
        RECT 27.660 153.100 27.980 153.160 ;
        RECT 29.590 153.145 29.730 153.640 ;
        RECT 36.025 153.640 37.640 153.780 ;
        RECT 36.025 153.485 36.165 153.640 ;
        RECT 37.320 153.580 37.640 153.640 ;
        RECT 55.350 153.640 59.170 153.780 ;
        RECT 35.950 153.255 36.240 153.485 ;
        RECT 36.400 153.240 36.720 153.500 ;
        RECT 40.540 153.240 40.860 153.500 ;
        RECT 41.475 153.440 41.765 153.485 ;
        RECT 44.680 153.440 45.000 153.500 ;
        RECT 41.475 153.300 45.000 153.440 ;
        RECT 41.475 153.255 41.765 153.300 ;
        RECT 25.375 152.960 27.980 153.100 ;
        RECT 25.375 152.915 25.665 152.960 ;
        RECT 27.660 152.900 27.980 152.960 ;
        RECT 29.515 153.100 29.805 153.145 ;
        RECT 36.490 153.100 36.630 153.240 ;
        RECT 29.515 152.960 36.630 153.100 ;
        RECT 29.515 152.915 29.805 152.960 ;
        RECT 41.550 152.820 41.690 153.255 ;
        RECT 44.680 153.240 45.000 153.300 ;
        RECT 50.660 153.440 50.980 153.500 ;
        RECT 55.350 153.485 55.490 153.640 ;
        RECT 59.030 153.485 59.170 153.640 ;
        RECT 64.945 153.640 68.945 153.780 ;
        RECT 64.945 153.595 65.235 153.640 ;
        RECT 67.465 153.595 67.755 153.640 ;
        RECT 68.655 153.595 68.945 153.640 ;
        RECT 72.280 153.580 72.600 153.840 ;
        RECT 73.215 153.780 73.505 153.825 ;
        RECT 75.960 153.780 76.280 153.840 ;
        RECT 82.875 153.780 83.165 153.825 ;
        RECT 84.240 153.780 84.560 153.840 ;
        RECT 73.215 153.640 76.280 153.780 ;
        RECT 73.215 153.595 73.505 153.640 ;
        RECT 75.960 153.580 76.280 153.640 ;
        RECT 82.030 153.640 84.560 153.780 ;
        RECT 55.275 153.440 55.565 153.485 ;
        RECT 58.035 153.440 58.325 153.485 ;
        RECT 50.660 153.300 55.565 153.440 ;
        RECT 50.660 153.240 50.980 153.300 ;
        RECT 55.275 153.255 55.565 153.300 ;
        RECT 57.190 153.300 58.325 153.440 ;
        RECT 52.960 153.100 53.280 153.160 ;
        RECT 54.355 153.100 54.645 153.145 ;
        RECT 52.960 152.960 54.645 153.100 ;
        RECT 52.960 152.900 53.280 152.960 ;
        RECT 54.355 152.915 54.645 152.960 ;
        RECT 55.720 153.100 56.040 153.160 ;
        RECT 57.190 153.145 57.330 153.300 ;
        RECT 58.035 153.255 58.325 153.300 ;
        RECT 58.955 153.255 59.245 153.485 ;
        RECT 68.255 153.440 68.545 153.485 ;
        RECT 69.060 153.440 69.380 153.500 ;
        RECT 68.255 153.300 69.380 153.440 ;
        RECT 68.255 153.255 68.545 153.300 ;
        RECT 69.060 153.240 69.380 153.300 ;
        RECT 69.520 153.240 69.840 153.500 ;
        RECT 73.660 153.440 73.980 153.500 ;
        RECT 82.030 153.440 82.170 153.640 ;
        RECT 82.875 153.595 83.165 153.640 ;
        RECT 84.240 153.580 84.560 153.640 ;
        RECT 84.700 153.580 85.020 153.840 ;
        RECT 97.210 153.825 97.350 153.980 ;
        RECT 100.340 153.920 100.660 153.980 ;
        RECT 109.540 154.120 109.860 154.180 ;
        RECT 110.935 154.120 111.225 154.165 ;
        RECT 120.135 154.120 120.425 154.165 ;
        RECT 121.040 154.120 121.360 154.180 ;
        RECT 109.540 153.980 111.225 154.120 ;
        RECT 109.540 153.920 109.860 153.980 ;
        RECT 110.935 153.935 111.225 153.980 ;
        RECT 116.070 153.980 121.360 154.120 ;
        RECT 97.135 153.595 97.425 153.825 ;
        RECT 97.580 153.780 97.900 153.840 ;
        RECT 116.070 153.825 116.210 153.980 ;
        RECT 120.135 153.935 120.425 153.980 ;
        RECT 121.040 153.920 121.360 153.980 ;
        RECT 122.460 154.120 122.750 154.165 ;
        RECT 124.560 154.120 124.850 154.165 ;
        RECT 126.130 154.120 126.420 154.165 ;
        RECT 122.460 153.980 126.420 154.120 ;
        RECT 122.460 153.935 122.750 153.980 ;
        RECT 124.560 153.935 124.850 153.980 ;
        RECT 126.130 153.935 126.420 153.980 ;
        RECT 128.875 154.120 129.165 154.165 ;
        RECT 128.875 153.980 132.770 154.120 ;
        RECT 128.875 153.935 129.165 153.980 ;
        RECT 132.630 153.840 132.770 153.980 ;
        RECT 101.735 153.780 102.025 153.825 ;
        RECT 97.580 153.640 102.025 153.780 ;
        RECT 97.580 153.580 97.900 153.640 ;
        RECT 101.735 153.595 102.025 153.640 ;
        RECT 115.995 153.595 116.285 153.825 ;
        RECT 116.440 153.780 116.760 153.840 ;
        RECT 121.500 153.780 121.820 153.840 ;
        RECT 121.975 153.780 122.265 153.825 ;
        RECT 116.440 153.640 122.265 153.780 ;
        RECT 116.440 153.580 116.760 153.640 ;
        RECT 121.500 153.580 121.820 153.640 ;
        RECT 121.975 153.595 122.265 153.640 ;
        RECT 122.855 153.780 123.145 153.825 ;
        RECT 124.045 153.780 124.335 153.825 ;
        RECT 126.565 153.780 126.855 153.825 ;
        RECT 122.855 153.640 126.855 153.780 ;
        RECT 122.855 153.595 123.145 153.640 ;
        RECT 124.045 153.595 124.335 153.640 ;
        RECT 126.565 153.595 126.855 153.640 ;
        RECT 132.540 153.580 132.860 153.840 ;
        RECT 73.660 153.300 82.170 153.440 ;
        RECT 82.415 153.440 82.705 153.485 ;
        RECT 101.260 153.440 101.580 153.500 ;
        RECT 104.495 153.440 104.785 153.485 ;
        RECT 82.415 153.300 101.030 153.440 ;
        RECT 73.660 153.240 73.980 153.300 ;
        RECT 82.415 153.255 82.705 153.300 ;
        RECT 57.115 153.100 57.405 153.145 ;
        RECT 55.720 152.960 57.405 153.100 ;
        RECT 55.720 152.900 56.040 152.960 ;
        RECT 57.115 152.915 57.405 152.960 ;
        RECT 71.835 153.100 72.125 153.145 ;
        RECT 71.835 152.960 75.730 153.100 ;
        RECT 71.835 152.915 72.125 152.960 ;
        RECT 22.600 152.760 22.920 152.820 ;
        RECT 18.550 152.620 22.920 152.760 ;
        RECT 22.600 152.560 22.920 152.620 ;
        RECT 23.520 152.560 23.840 152.820 ;
        RECT 26.740 152.560 27.060 152.820 ;
        RECT 28.595 152.760 28.885 152.805 ;
        RECT 31.800 152.760 32.120 152.820 ;
        RECT 28.595 152.620 32.120 152.760 ;
        RECT 28.595 152.575 28.885 152.620 ;
        RECT 31.800 152.560 32.120 152.620 ;
        RECT 34.560 152.560 34.880 152.820 ;
        RECT 40.095 152.760 40.385 152.805 ;
        RECT 41.460 152.760 41.780 152.820 ;
        RECT 40.095 152.620 41.780 152.760 ;
        RECT 40.095 152.575 40.385 152.620 ;
        RECT 41.460 152.560 41.780 152.620 ;
        RECT 52.500 152.760 52.820 152.820 ;
        RECT 56.655 152.760 56.945 152.805 ;
        RECT 52.500 152.620 56.945 152.760 ;
        RECT 52.500 152.560 52.820 152.620 ;
        RECT 56.655 152.575 56.945 152.620 ;
        RECT 58.940 152.560 59.260 152.820 ;
        RECT 74.580 152.560 74.900 152.820 ;
        RECT 75.590 152.760 75.730 152.960 ;
        RECT 75.960 152.900 76.280 153.160 ;
        RECT 96.675 153.100 96.965 153.145 ;
        RECT 100.340 153.100 100.660 153.160 ;
        RECT 96.675 152.960 100.660 153.100 ;
        RECT 100.890 153.100 101.030 153.300 ;
        RECT 101.260 153.300 104.785 153.440 ;
        RECT 101.260 153.240 101.580 153.300 ;
        RECT 104.495 153.255 104.785 153.300 ;
        RECT 107.715 153.440 108.005 153.485 ;
        RECT 108.175 153.440 108.465 153.485 ;
        RECT 107.715 153.300 108.465 153.440 ;
        RECT 107.715 153.255 108.005 153.300 ;
        RECT 108.175 153.255 108.465 153.300 ;
        RECT 108.620 153.440 108.940 153.500 ;
        RECT 110.475 153.440 110.765 153.485 ;
        RECT 108.620 153.300 110.765 153.440 ;
        RECT 108.620 153.240 108.940 153.300 ;
        RECT 110.475 153.255 110.765 153.300 ;
        RECT 111.380 153.240 111.700 153.500 ;
        RECT 117.360 153.240 117.680 153.500 ;
        RECT 121.040 153.440 121.360 153.500 ;
        RECT 126.100 153.440 126.420 153.500 ;
        RECT 121.040 153.300 126.420 153.440 ;
        RECT 121.040 153.240 121.360 153.300 ;
        RECT 126.100 153.240 126.420 153.300 ;
        RECT 133.920 153.240 134.240 153.500 ;
        RECT 135.775 153.255 136.065 153.485 ;
        RECT 109.080 153.100 109.400 153.160 ;
        RECT 100.890 152.960 109.400 153.100 ;
        RECT 96.675 152.915 96.965 152.960 ;
        RECT 100.340 152.900 100.660 152.960 ;
        RECT 109.080 152.900 109.400 152.960 ;
        RECT 123.310 153.100 123.600 153.145 ;
        RECT 124.260 153.100 124.580 153.160 ;
        RECT 123.310 152.960 124.580 153.100 ;
        RECT 123.310 152.915 123.600 152.960 ;
        RECT 124.260 152.900 124.580 152.960 ;
        RECT 124.720 153.100 125.040 153.160 ;
        RECT 135.850 153.100 135.990 153.255 ;
        RECT 124.720 152.960 135.990 153.100 ;
        RECT 124.720 152.900 125.040 152.960 ;
        RECT 80.115 152.760 80.405 152.805 ;
        RECT 75.590 152.620 80.405 152.760 ;
        RECT 80.115 152.575 80.405 152.620 ;
        RECT 81.940 152.560 82.260 152.820 ;
        RECT 87.460 152.560 87.780 152.820 ;
        RECT 100.800 152.560 101.120 152.820 ;
        RECT 112.760 152.760 113.080 152.820 ;
        RECT 116.915 152.760 117.205 152.805 ;
        RECT 112.760 152.620 117.205 152.760 ;
        RECT 112.760 152.560 113.080 152.620 ;
        RECT 116.915 152.575 117.205 152.620 ;
        RECT 129.320 152.760 129.640 152.820 ;
        RECT 129.795 152.760 130.085 152.805 ;
        RECT 129.320 152.620 130.085 152.760 ;
        RECT 129.320 152.560 129.640 152.620 ;
        RECT 129.795 152.575 130.085 152.620 ;
        RECT 134.840 152.560 135.160 152.820 ;
        RECT 13.330 151.940 138.910 152.420 ;
        RECT 21.695 151.740 21.985 151.785 ;
        RECT 23.520 151.740 23.840 151.800 ;
        RECT 21.695 151.600 23.840 151.740 ;
        RECT 21.695 151.555 21.985 151.600 ;
        RECT 23.520 151.540 23.840 151.600 ;
        RECT 27.660 151.740 27.980 151.800 ;
        RECT 29.975 151.740 30.265 151.785 ;
        RECT 35.480 151.740 35.800 151.800 ;
        RECT 27.660 151.600 30.265 151.740 ;
        RECT 27.660 151.540 27.980 151.600 ;
        RECT 29.975 151.555 30.265 151.600 ;
        RECT 32.810 151.600 35.800 151.740 ;
        RECT 17.555 151.215 17.845 151.445 ;
        RECT 22.615 151.400 22.905 151.445 ;
        RECT 24.300 151.400 24.590 151.445 ;
        RECT 22.615 151.260 24.590 151.400 ;
        RECT 30.050 151.400 30.190 151.555 ;
        RECT 30.050 151.260 31.110 151.400 ;
        RECT 22.615 151.215 22.905 151.260 ;
        RECT 24.300 151.215 24.590 151.260 ;
        RECT 17.630 151.060 17.770 151.215 ;
        RECT 20.760 151.060 21.080 151.120 ;
        RECT 17.630 150.920 21.080 151.060 ;
        RECT 20.760 150.860 21.080 150.920 ;
        RECT 21.235 151.060 21.525 151.105 ;
        RECT 22.140 151.060 22.460 151.120 ;
        RECT 23.520 151.060 23.840 151.120 ;
        RECT 21.235 150.920 23.840 151.060 ;
        RECT 21.235 150.875 21.525 150.920 ;
        RECT 22.140 150.860 22.460 150.920 ;
        RECT 23.520 150.860 23.840 150.920 ;
        RECT 28.580 151.060 28.900 151.120 ;
        RECT 30.435 151.060 30.725 151.105 ;
        RECT 28.580 150.920 30.725 151.060 ;
        RECT 28.580 150.860 28.900 150.920 ;
        RECT 30.435 150.875 30.725 150.920 ;
        RECT 17.630 150.580 20.070 150.720 ;
        RECT 16.635 150.040 16.925 150.085 ;
        RECT 17.080 150.040 17.400 150.100 ;
        RECT 17.630 150.085 17.770 150.580 ;
        RECT 19.930 150.425 20.070 150.580 ;
        RECT 23.060 150.520 23.380 150.780 ;
        RECT 23.955 150.720 24.245 150.765 ;
        RECT 25.145 150.720 25.435 150.765 ;
        RECT 27.665 150.720 27.955 150.765 ;
        RECT 23.955 150.580 27.955 150.720 ;
        RECT 30.970 150.720 31.110 151.260 ;
        RECT 32.810 151.105 32.950 151.600 ;
        RECT 35.480 151.540 35.800 151.600 ;
        RECT 69.075 151.740 69.365 151.785 ;
        RECT 74.120 151.740 74.440 151.800 ;
        RECT 69.075 151.600 74.440 151.740 ;
        RECT 69.075 151.555 69.365 151.600 ;
        RECT 74.120 151.540 74.440 151.600 ;
        RECT 74.580 151.740 74.900 151.800 ;
        RECT 85.635 151.740 85.925 151.785 ;
        RECT 87.460 151.740 87.780 151.800 ;
        RECT 74.580 151.600 85.390 151.740 ;
        RECT 74.580 151.540 74.900 151.600 ;
        RECT 33.195 151.400 33.485 151.445 ;
        RECT 34.560 151.400 34.880 151.460 ;
        RECT 35.035 151.400 35.325 151.445 ;
        RECT 33.195 151.260 34.330 151.400 ;
        RECT 33.195 151.215 33.485 151.260 ;
        RECT 34.190 151.105 34.330 151.260 ;
        RECT 34.560 151.260 35.325 151.400 ;
        RECT 34.560 151.200 34.880 151.260 ;
        RECT 35.035 151.215 35.325 151.260 ;
        RECT 36.860 151.400 37.180 151.460 ;
        RECT 39.635 151.400 39.925 151.445 ;
        RECT 62.620 151.400 62.940 151.460 ;
        RECT 69.520 151.400 69.840 151.460 ;
        RECT 36.860 151.260 39.925 151.400 ;
        RECT 36.860 151.200 37.180 151.260 ;
        RECT 39.635 151.215 39.925 151.260 ;
        RECT 57.650 151.260 76.190 151.400 ;
        RECT 32.735 150.875 33.025 151.105 ;
        RECT 33.655 150.875 33.945 151.105 ;
        RECT 34.115 150.875 34.405 151.105 ;
        RECT 35.495 150.875 35.785 151.105 ;
        RECT 35.955 151.060 36.245 151.105 ;
        RECT 37.780 151.060 38.100 151.120 ;
        RECT 41.000 151.060 41.320 151.120 ;
        RECT 35.955 150.920 41.320 151.060 ;
        RECT 35.955 150.875 36.245 150.920 ;
        RECT 33.730 150.720 33.870 150.875 ;
        RECT 35.570 150.720 35.710 150.875 ;
        RECT 37.780 150.860 38.100 150.920 ;
        RECT 41.000 150.860 41.320 150.920 ;
        RECT 41.475 151.060 41.765 151.105 ;
        RECT 46.060 151.060 46.380 151.120 ;
        RECT 53.420 151.060 53.740 151.120 ;
        RECT 41.475 150.920 53.740 151.060 ;
        RECT 41.475 150.875 41.765 150.920 ;
        RECT 46.060 150.860 46.380 150.920 ;
        RECT 30.970 150.580 35.710 150.720 ;
        RECT 36.400 150.720 36.720 150.780 ;
        RECT 40.555 150.720 40.845 150.765 ;
        RECT 36.400 150.580 40.845 150.720 ;
        RECT 23.955 150.535 24.245 150.580 ;
        RECT 25.145 150.535 25.435 150.580 ;
        RECT 27.665 150.535 27.955 150.580 ;
        RECT 36.400 150.520 36.720 150.580 ;
        RECT 40.555 150.535 40.845 150.580 ;
        RECT 19.395 150.195 19.685 150.425 ;
        RECT 19.855 150.380 20.145 150.425 ;
        RECT 21.220 150.380 21.540 150.440 ;
        RECT 19.855 150.240 21.540 150.380 ;
        RECT 19.855 150.195 20.145 150.240 ;
        RECT 16.635 149.900 17.400 150.040 ;
        RECT 16.635 149.855 16.925 149.900 ;
        RECT 17.080 149.840 17.400 149.900 ;
        RECT 17.555 149.855 17.845 150.085 ;
        RECT 19.470 150.040 19.610 150.195 ;
        RECT 21.220 150.180 21.540 150.240 ;
        RECT 23.560 150.380 23.850 150.425 ;
        RECT 25.660 150.380 25.950 150.425 ;
        RECT 27.230 150.380 27.520 150.425 ;
        RECT 23.560 150.240 27.520 150.380 ;
        RECT 23.560 150.195 23.850 150.240 ;
        RECT 25.660 150.195 25.950 150.240 ;
        RECT 27.230 150.195 27.520 150.240 ;
        RECT 41.000 150.180 41.320 150.440 ;
        RECT 50.290 150.425 50.430 150.920 ;
        RECT 53.420 150.860 53.740 150.920 ;
        RECT 53.880 151.060 54.200 151.120 ;
        RECT 55.780 151.060 56.070 151.105 ;
        RECT 53.880 150.920 56.070 151.060 ;
        RECT 53.880 150.860 54.200 150.920 ;
        RECT 55.780 150.875 56.070 150.920 ;
        RECT 56.640 151.060 56.960 151.120 ;
        RECT 57.650 151.105 57.790 151.260 ;
        RECT 62.620 151.200 62.940 151.260 ;
        RECT 69.520 151.200 69.840 151.260 ;
        RECT 58.940 151.105 59.260 151.120 ;
        RECT 57.115 151.060 57.405 151.105 ;
        RECT 57.575 151.060 57.865 151.105 ;
        RECT 58.910 151.060 59.260 151.105 ;
        RECT 56.640 150.920 57.865 151.060 ;
        RECT 58.745 150.920 59.260 151.060 ;
        RECT 56.640 150.860 56.960 150.920 ;
        RECT 57.115 150.875 57.405 150.920 ;
        RECT 57.575 150.875 57.865 150.920 ;
        RECT 58.910 150.875 59.260 150.920 ;
        RECT 58.940 150.860 59.260 150.875 ;
        RECT 65.840 150.860 66.160 151.120 ;
        RECT 66.760 150.860 67.080 151.120 ;
        RECT 68.615 151.060 68.905 151.105 ;
        RECT 73.200 151.060 73.520 151.120 ;
        RECT 68.615 150.920 73.520 151.060 ;
        RECT 68.615 150.875 68.905 150.920 ;
        RECT 73.200 150.860 73.520 150.920 ;
        RECT 74.580 151.105 74.900 151.120 ;
        RECT 76.050 151.105 76.190 151.260 ;
        RECT 77.800 151.105 78.120 151.120 ;
        RECT 74.580 151.060 74.930 151.105 ;
        RECT 75.975 151.060 76.265 151.105 ;
        RECT 76.435 151.060 76.725 151.105 ;
        RECT 74.580 150.920 75.095 151.060 ;
        RECT 75.975 150.920 76.725 151.060 ;
        RECT 74.580 150.875 74.930 150.920 ;
        RECT 75.975 150.875 76.265 150.920 ;
        RECT 76.435 150.875 76.725 150.920 ;
        RECT 77.770 150.875 78.120 151.105 ;
        RECT 74.580 150.860 74.900 150.875 ;
        RECT 77.800 150.860 78.120 150.875 ;
        RECT 52.525 150.720 52.815 150.765 ;
        RECT 55.045 150.720 55.335 150.765 ;
        RECT 56.235 150.720 56.525 150.765 ;
        RECT 52.525 150.580 56.525 150.720 ;
        RECT 52.525 150.535 52.815 150.580 ;
        RECT 55.045 150.535 55.335 150.580 ;
        RECT 56.235 150.535 56.525 150.580 ;
        RECT 58.455 150.720 58.745 150.765 ;
        RECT 59.645 150.720 59.935 150.765 ;
        RECT 62.165 150.720 62.455 150.765 ;
        RECT 58.455 150.580 62.455 150.720 ;
        RECT 58.455 150.535 58.745 150.580 ;
        RECT 59.645 150.535 59.935 150.580 ;
        RECT 62.165 150.535 62.455 150.580 ;
        RECT 71.385 150.720 71.675 150.765 ;
        RECT 73.905 150.720 74.195 150.765 ;
        RECT 75.095 150.720 75.385 150.765 ;
        RECT 71.385 150.580 75.385 150.720 ;
        RECT 71.385 150.535 71.675 150.580 ;
        RECT 73.905 150.535 74.195 150.580 ;
        RECT 75.095 150.535 75.385 150.580 ;
        RECT 77.315 150.720 77.605 150.765 ;
        RECT 78.505 150.720 78.795 150.765 ;
        RECT 81.025 150.720 81.315 150.765 ;
        RECT 77.315 150.580 81.315 150.720 ;
        RECT 77.315 150.535 77.605 150.580 ;
        RECT 78.505 150.535 78.795 150.580 ;
        RECT 81.025 150.535 81.315 150.580 ;
        RECT 83.780 150.520 84.100 150.780 ;
        RECT 85.250 150.720 85.390 151.600 ;
        RECT 85.635 151.600 87.780 151.740 ;
        RECT 85.635 151.555 85.925 151.600 ;
        RECT 87.460 151.540 87.780 151.600 ;
        RECT 117.820 151.740 118.140 151.800 ;
        RECT 117.820 151.600 118.970 151.740 ;
        RECT 117.820 151.540 118.140 151.600 ;
        RECT 86.095 151.400 86.385 151.445 ;
        RECT 86.540 151.400 86.860 151.460 ;
        RECT 86.095 151.260 86.860 151.400 ;
        RECT 86.095 151.215 86.385 151.260 ;
        RECT 86.540 151.200 86.860 151.260 ;
        RECT 93.440 151.400 93.760 151.460 ;
        RECT 93.440 151.260 98.270 151.400 ;
        RECT 93.440 151.200 93.760 151.260 ;
        RECT 98.130 151.105 98.270 151.260 ;
        RECT 118.280 151.200 118.600 151.460 ;
        RECT 92.995 151.060 93.285 151.105 ;
        RECT 95.295 151.060 95.585 151.105 ;
        RECT 92.995 150.920 95.585 151.060 ;
        RECT 92.995 150.875 93.285 150.920 ;
        RECT 95.295 150.875 95.585 150.920 ;
        RECT 98.055 150.875 98.345 151.105 ;
        RECT 115.060 151.060 115.380 151.120 ;
        RECT 118.830 151.105 118.970 151.600 ;
        RECT 124.260 151.540 124.580 151.800 ;
        RECT 126.115 151.740 126.405 151.785 ;
        RECT 129.320 151.740 129.640 151.800 ;
        RECT 126.115 151.600 129.640 151.740 ;
        RECT 126.115 151.555 126.405 151.600 ;
        RECT 129.320 151.540 129.640 151.600 ;
        RECT 133.475 151.740 133.765 151.785 ;
        RECT 133.920 151.740 134.240 151.800 ;
        RECT 133.475 151.600 134.240 151.740 ;
        RECT 133.475 151.555 133.765 151.600 ;
        RECT 133.920 151.540 134.240 151.600 ;
        RECT 126.560 151.200 126.880 151.460 ;
        RECT 117.835 151.060 118.125 151.105 ;
        RECT 115.060 150.920 118.125 151.060 ;
        RECT 115.060 150.860 115.380 150.920 ;
        RECT 117.835 150.875 118.125 150.920 ;
        RECT 118.755 150.875 119.045 151.105 ;
        RECT 132.540 150.860 132.860 151.120 ;
        RECT 86.555 150.720 86.845 150.765 ;
        RECT 85.250 150.580 86.845 150.720 ;
        RECT 86.555 150.535 86.845 150.580 ;
        RECT 91.600 150.720 91.920 150.780 ;
        RECT 93.455 150.720 93.745 150.765 ;
        RECT 91.600 150.580 93.745 150.720 ;
        RECT 50.215 150.195 50.505 150.425 ;
        RECT 52.960 150.380 53.250 150.425 ;
        RECT 54.530 150.380 54.820 150.425 ;
        RECT 56.630 150.380 56.920 150.425 ;
        RECT 52.960 150.240 56.920 150.380 ;
        RECT 52.960 150.195 53.250 150.240 ;
        RECT 54.530 150.195 54.820 150.240 ;
        RECT 56.630 150.195 56.920 150.240 ;
        RECT 58.060 150.380 58.350 150.425 ;
        RECT 60.160 150.380 60.450 150.425 ;
        RECT 61.730 150.380 62.020 150.425 ;
        RECT 58.060 150.240 62.020 150.380 ;
        RECT 58.060 150.195 58.350 150.240 ;
        RECT 60.160 150.195 60.450 150.240 ;
        RECT 61.730 150.195 62.020 150.240 ;
        RECT 71.820 150.380 72.110 150.425 ;
        RECT 73.390 150.380 73.680 150.425 ;
        RECT 75.490 150.380 75.780 150.425 ;
        RECT 71.820 150.240 75.780 150.380 ;
        RECT 71.820 150.195 72.110 150.240 ;
        RECT 73.390 150.195 73.680 150.240 ;
        RECT 75.490 150.195 75.780 150.240 ;
        RECT 76.920 150.380 77.210 150.425 ;
        RECT 79.020 150.380 79.310 150.425 ;
        RECT 80.590 150.380 80.880 150.425 ;
        RECT 76.920 150.240 80.880 150.380 ;
        RECT 83.870 150.380 84.010 150.520 ;
        RECT 85.620 150.380 85.940 150.440 ;
        RECT 83.870 150.240 85.940 150.380 ;
        RECT 86.630 150.380 86.770 150.535 ;
        RECT 91.600 150.520 91.920 150.580 ;
        RECT 93.455 150.535 93.745 150.580 ;
        RECT 93.915 150.535 94.205 150.765 ;
        RECT 110.000 150.720 110.320 150.780 ;
        RECT 110.000 150.580 122.650 150.720 ;
        RECT 93.990 150.380 94.130 150.535 ;
        RECT 110.000 150.520 110.320 150.580 ;
        RECT 86.630 150.240 94.130 150.380 ;
        RECT 94.360 150.380 94.680 150.440 ;
        RECT 121.040 150.380 121.360 150.440 ;
        RECT 94.360 150.240 121.360 150.380 ;
        RECT 122.510 150.380 122.650 150.580 ;
        RECT 127.035 150.535 127.325 150.765 ;
        RECT 127.110 150.380 127.250 150.535 ;
        RECT 122.510 150.240 127.250 150.380 ;
        RECT 76.920 150.195 77.210 150.240 ;
        RECT 79.020 150.195 79.310 150.240 ;
        RECT 80.590 150.195 80.880 150.240 ;
        RECT 85.620 150.180 85.940 150.240 ;
        RECT 94.360 150.180 94.680 150.240 ;
        RECT 121.040 150.180 121.360 150.240 ;
        RECT 22.140 150.040 22.460 150.100 ;
        RECT 24.440 150.040 24.760 150.100 ;
        RECT 19.470 149.900 24.760 150.040 ;
        RECT 22.140 149.840 22.460 149.900 ;
        RECT 24.440 149.840 24.760 149.900 ;
        RECT 26.280 150.040 26.600 150.100 ;
        RECT 30.895 150.040 31.185 150.085 ;
        RECT 26.280 149.900 31.185 150.040 ;
        RECT 26.280 149.840 26.600 149.900 ;
        RECT 30.895 149.855 31.185 149.900 ;
        RECT 32.720 150.040 33.040 150.100 ;
        RECT 35.940 150.040 36.260 150.100 ;
        RECT 32.720 149.900 36.260 150.040 ;
        RECT 32.720 149.840 33.040 149.900 ;
        RECT 35.940 149.840 36.260 149.900 ;
        RECT 36.875 150.040 37.165 150.085 ;
        RECT 38.240 150.040 38.560 150.100 ;
        RECT 36.875 149.900 38.560 150.040 ;
        RECT 36.875 149.855 37.165 149.900 ;
        RECT 38.240 149.840 38.560 149.900 ;
        RECT 40.540 149.840 40.860 150.100 ;
        RECT 64.460 149.840 64.780 150.100 ;
        RECT 77.340 150.040 77.660 150.100 ;
        RECT 81.940 150.040 82.260 150.100 ;
        RECT 83.335 150.040 83.625 150.085 ;
        RECT 77.340 149.900 83.625 150.040 ;
        RECT 77.340 149.840 77.660 149.900 ;
        RECT 81.940 149.840 82.260 149.900 ;
        RECT 83.335 149.855 83.625 149.900 ;
        RECT 83.795 150.040 84.085 150.085 ;
        RECT 84.700 150.040 85.020 150.100 ;
        RECT 83.795 149.900 85.020 150.040 ;
        RECT 83.795 149.855 84.085 149.900 ;
        RECT 84.700 149.840 85.020 149.900 ;
        RECT 91.140 149.840 91.460 150.100 ;
        RECT 116.440 150.040 116.760 150.100 ;
        RECT 132.080 150.040 132.400 150.100 ;
        RECT 116.440 149.900 132.400 150.040 ;
        RECT 116.440 149.840 116.760 149.900 ;
        RECT 132.080 149.840 132.400 149.900 ;
        RECT 13.330 149.220 138.910 149.700 ;
        RECT 23.535 148.835 23.825 149.065 ;
        RECT 17.120 148.680 17.410 148.725 ;
        RECT 19.220 148.680 19.510 148.725 ;
        RECT 20.790 148.680 21.080 148.725 ;
        RECT 17.120 148.540 21.080 148.680 ;
        RECT 23.610 148.680 23.750 148.835 ;
        RECT 23.980 148.820 24.300 149.080 ;
        RECT 24.900 149.020 25.220 149.080 ;
        RECT 26.280 149.020 26.600 149.080 ;
        RECT 24.900 148.880 26.600 149.020 ;
        RECT 24.900 148.820 25.220 148.880 ;
        RECT 26.280 148.820 26.600 148.880 ;
        RECT 29.975 149.020 30.265 149.065 ;
        RECT 31.800 149.020 32.120 149.080 ;
        RECT 33.180 149.020 33.500 149.080 ;
        RECT 35.955 149.020 36.245 149.065 ;
        RECT 29.975 148.880 33.500 149.020 ;
        RECT 29.975 148.835 30.265 148.880 ;
        RECT 24.440 148.680 24.760 148.740 ;
        RECT 30.050 148.680 30.190 148.835 ;
        RECT 31.800 148.820 32.120 148.880 ;
        RECT 33.180 148.820 33.500 148.880 ;
        RECT 33.730 148.880 36.245 149.020 ;
        RECT 23.610 148.540 30.190 148.680 ;
        RECT 17.120 148.495 17.410 148.540 ;
        RECT 19.220 148.495 19.510 148.540 ;
        RECT 20.790 148.495 21.080 148.540 ;
        RECT 24.440 148.480 24.760 148.540 ;
        RECT 30.895 148.495 31.185 148.725 ;
        RECT 17.515 148.340 17.805 148.385 ;
        RECT 18.705 148.340 18.995 148.385 ;
        RECT 21.225 148.340 21.515 148.385 ;
        RECT 17.515 148.200 21.515 148.340 ;
        RECT 17.515 148.155 17.805 148.200 ;
        RECT 18.705 148.155 18.995 148.200 ;
        RECT 21.225 148.155 21.515 148.200 ;
        RECT 23.520 148.340 23.840 148.400 ;
        RECT 27.215 148.340 27.505 148.385 ;
        RECT 30.970 148.340 31.110 148.495 ;
        RECT 33.730 148.340 33.870 148.880 ;
        RECT 35.955 148.835 36.245 148.880 ;
        RECT 48.360 149.020 48.680 149.080 ;
        RECT 50.675 149.020 50.965 149.065 ;
        RECT 55.720 149.020 56.040 149.080 ;
        RECT 48.360 148.880 56.040 149.020 ;
        RECT 48.360 148.820 48.680 148.880 ;
        RECT 50.675 148.835 50.965 148.880 ;
        RECT 55.720 148.820 56.040 148.880 ;
        RECT 65.395 149.020 65.685 149.065 ;
        RECT 65.840 149.020 66.160 149.080 ;
        RECT 65.395 148.880 66.160 149.020 ;
        RECT 65.395 148.835 65.685 148.880 ;
        RECT 65.840 148.820 66.160 148.880 ;
        RECT 66.315 149.020 66.605 149.065 ;
        RECT 94.360 149.020 94.680 149.080 ;
        RECT 66.315 148.880 94.680 149.020 ;
        RECT 66.315 148.835 66.605 148.880 ;
        RECT 94.360 148.820 94.680 148.880 ;
        RECT 100.800 149.020 101.120 149.080 ;
        RECT 101.735 149.020 102.025 149.065 ;
        RECT 100.800 148.880 102.025 149.020 ;
        RECT 100.800 148.820 101.120 148.880 ;
        RECT 101.735 148.835 102.025 148.880 ;
        RECT 109.080 149.020 109.400 149.080 ;
        RECT 118.740 149.020 119.060 149.080 ;
        RECT 121.960 149.020 122.280 149.080 ;
        RECT 109.080 148.880 122.280 149.020 ;
        RECT 34.100 148.680 34.420 148.740 ;
        RECT 37.795 148.680 38.085 148.725 ;
        RECT 34.100 148.540 38.085 148.680 ;
        RECT 34.100 148.480 34.420 148.540 ;
        RECT 37.795 148.495 38.085 148.540 ;
        RECT 51.595 148.495 51.885 148.725 ;
        RECT 53.000 148.680 53.290 148.725 ;
        RECT 55.100 148.680 55.390 148.725 ;
        RECT 56.670 148.680 56.960 148.725 ;
        RECT 53.000 148.540 56.960 148.680 ;
        RECT 65.930 148.680 66.070 148.820 ;
        RECT 67.680 148.680 68.000 148.740 ;
        RECT 65.930 148.540 68.000 148.680 ;
        RECT 53.000 148.495 53.290 148.540 ;
        RECT 55.100 148.495 55.390 148.540 ;
        RECT 56.670 148.495 56.960 148.540 ;
        RECT 23.520 148.200 27.505 148.340 ;
        RECT 23.520 148.140 23.840 148.200 ;
        RECT 15.700 148.000 16.020 148.060 ;
        RECT 16.635 148.000 16.925 148.045 ;
        RECT 23.060 148.000 23.380 148.060 ;
        RECT 24.990 148.045 25.130 148.200 ;
        RECT 27.215 148.155 27.505 148.200 ;
        RECT 29.590 148.200 30.650 148.340 ;
        RECT 30.970 148.200 32.490 148.340 ;
        RECT 15.700 147.860 23.380 148.000 ;
        RECT 15.700 147.800 16.020 147.860 ;
        RECT 16.635 147.815 16.925 147.860 ;
        RECT 23.060 147.800 23.380 147.860 ;
        RECT 24.915 147.815 25.205 148.045 ;
        RECT 25.820 147.800 26.140 148.060 ;
        RECT 26.280 148.000 26.600 148.060 ;
        RECT 26.755 148.000 27.045 148.045 ;
        RECT 26.280 147.860 27.045 148.000 ;
        RECT 26.280 147.800 26.600 147.860 ;
        RECT 26.755 147.815 27.045 147.860 ;
        RECT 27.660 147.800 27.980 148.060 ;
        RECT 28.120 147.800 28.440 148.060 ;
        RECT 17.970 147.660 18.260 147.705 ;
        RECT 18.460 147.660 18.780 147.720 ;
        RECT 17.970 147.520 18.780 147.660 ;
        RECT 25.910 147.660 26.050 147.800 ;
        RECT 29.590 147.660 29.730 148.200 ;
        RECT 29.975 147.815 30.265 148.045 ;
        RECT 25.910 147.520 29.730 147.660 ;
        RECT 17.970 147.475 18.260 147.520 ;
        RECT 18.460 147.460 18.780 147.520 ;
        RECT 30.050 147.320 30.190 147.815 ;
        RECT 30.510 147.660 30.650 148.200 ;
        RECT 31.340 147.800 31.660 148.060 ;
        RECT 31.800 148.000 32.120 148.060 ;
        RECT 32.350 148.045 32.490 148.200 ;
        RECT 33.270 148.200 33.870 148.340 ;
        RECT 34.560 148.340 34.880 148.400 ;
        RECT 38.240 148.340 38.560 148.400 ;
        RECT 34.560 148.200 38.560 148.340 ;
        RECT 32.275 148.000 32.565 148.045 ;
        RECT 31.800 147.860 32.565 148.000 ;
        RECT 31.800 147.800 32.120 147.860 ;
        RECT 32.275 147.815 32.565 147.860 ;
        RECT 32.720 147.800 33.040 148.060 ;
        RECT 33.270 148.045 33.410 148.200 ;
        RECT 34.560 148.140 34.880 148.200 ;
        RECT 38.240 148.140 38.560 148.200 ;
        RECT 33.195 147.815 33.485 148.045 ;
        RECT 35.480 148.000 35.800 148.060 ;
        RECT 33.730 147.860 35.800 148.000 ;
        RECT 33.270 147.660 33.410 147.815 ;
        RECT 30.510 147.520 33.410 147.660 ;
        RECT 33.730 147.320 33.870 147.860 ;
        RECT 35.480 147.800 35.800 147.860 ;
        RECT 38.700 148.000 39.020 148.060 ;
        RECT 39.175 148.000 39.465 148.045 ;
        RECT 38.700 147.860 39.465 148.000 ;
        RECT 38.700 147.800 39.020 147.860 ;
        RECT 39.175 147.815 39.465 147.860 ;
        RECT 39.635 148.000 39.925 148.045 ;
        RECT 40.540 148.000 40.860 148.060 ;
        RECT 39.635 147.860 40.860 148.000 ;
        RECT 39.635 147.815 39.925 147.860 ;
        RECT 40.540 147.800 40.860 147.860 ;
        RECT 41.000 148.000 41.320 148.060 ;
        RECT 43.315 148.000 43.605 148.045 ;
        RECT 41.000 147.860 43.605 148.000 ;
        RECT 41.000 147.800 41.320 147.860 ;
        RECT 43.315 147.815 43.605 147.860 ;
        RECT 44.695 148.000 44.985 148.045 ;
        RECT 47.900 148.000 48.220 148.060 ;
        RECT 44.695 147.860 48.220 148.000 ;
        RECT 44.695 147.815 44.985 147.860 ;
        RECT 47.900 147.800 48.220 147.860 ;
        RECT 50.660 147.800 50.980 148.060 ;
        RECT 51.670 148.000 51.810 148.495 ;
        RECT 67.680 148.480 68.000 148.540 ;
        RECT 81.940 148.680 82.230 148.725 ;
        RECT 83.510 148.680 83.800 148.725 ;
        RECT 85.610 148.680 85.900 148.725 ;
        RECT 81.940 148.540 85.900 148.680 ;
        RECT 81.940 148.495 82.230 148.540 ;
        RECT 83.510 148.495 83.800 148.540 ;
        RECT 85.610 148.495 85.900 148.540 ;
        RECT 87.040 148.680 87.330 148.725 ;
        RECT 89.140 148.680 89.430 148.725 ;
        RECT 90.710 148.680 91.000 148.725 ;
        RECT 87.040 148.540 91.000 148.680 ;
        RECT 87.040 148.495 87.330 148.540 ;
        RECT 89.140 148.495 89.430 148.540 ;
        RECT 90.710 148.495 91.000 148.540 ;
        RECT 93.440 148.480 93.760 148.740 ;
        RECT 95.320 148.680 95.610 148.725 ;
        RECT 97.420 148.680 97.710 148.725 ;
        RECT 98.990 148.680 99.280 148.725 ;
        RECT 95.320 148.540 99.280 148.680 ;
        RECT 95.320 148.495 95.610 148.540 ;
        RECT 97.420 148.495 97.710 148.540 ;
        RECT 98.990 148.495 99.280 148.540 ;
        RECT 53.395 148.340 53.685 148.385 ;
        RECT 54.585 148.340 54.875 148.385 ;
        RECT 57.105 148.340 57.395 148.385 ;
        RECT 53.395 148.200 57.395 148.340 ;
        RECT 53.395 148.155 53.685 148.200 ;
        RECT 54.585 148.155 54.875 148.200 ;
        RECT 57.105 148.155 57.395 148.200 ;
        RECT 64.460 148.340 64.780 148.400 ;
        RECT 68.600 148.340 68.920 148.400 ;
        RECT 64.460 148.200 71.590 148.340 ;
        RECT 64.460 148.140 64.780 148.200 ;
        RECT 68.600 148.140 68.920 148.200 ;
        RECT 52.515 148.000 52.805 148.045 ;
        RECT 56.640 148.000 56.960 148.060 ;
        RECT 51.670 147.860 52.270 148.000 ;
        RECT 34.575 147.660 34.865 147.705 ;
        RECT 36.860 147.660 37.180 147.720 ;
        RECT 34.575 147.520 37.180 147.660 ;
        RECT 34.575 147.475 34.865 147.520 ;
        RECT 36.860 147.460 37.180 147.520 ;
        RECT 45.615 147.660 45.905 147.705 ;
        RECT 49.755 147.660 50.045 147.705 ;
        RECT 50.750 147.660 50.890 147.800 ;
        RECT 45.615 147.520 50.890 147.660 ;
        RECT 52.130 147.660 52.270 147.860 ;
        RECT 52.515 147.860 56.960 148.000 ;
        RECT 52.515 147.815 52.805 147.860 ;
        RECT 56.640 147.800 56.960 147.860 ;
        RECT 66.760 148.000 67.080 148.060 ;
        RECT 67.235 148.000 67.525 148.045 ;
        RECT 66.760 147.860 67.525 148.000 ;
        RECT 66.760 147.800 67.080 147.860 ;
        RECT 67.235 147.815 67.525 147.860 ;
        RECT 67.680 148.000 68.000 148.060 ;
        RECT 71.450 148.045 71.590 148.200 ;
        RECT 72.740 148.140 73.060 148.400 ;
        RECT 77.340 148.140 77.660 148.400 ;
        RECT 81.505 148.340 81.795 148.385 ;
        RECT 84.025 148.340 84.315 148.385 ;
        RECT 85.215 148.340 85.505 148.385 ;
        RECT 81.505 148.200 85.505 148.340 ;
        RECT 81.505 148.155 81.795 148.200 ;
        RECT 84.025 148.155 84.315 148.200 ;
        RECT 85.215 148.155 85.505 148.200 ;
        RECT 87.435 148.340 87.725 148.385 ;
        RECT 88.625 148.340 88.915 148.385 ;
        RECT 91.145 148.340 91.435 148.385 ;
        RECT 87.435 148.200 91.435 148.340 ;
        RECT 87.435 148.155 87.725 148.200 ;
        RECT 88.625 148.155 88.915 148.200 ;
        RECT 91.145 148.155 91.435 148.200 ;
        RECT 95.715 148.340 96.005 148.385 ;
        RECT 96.905 148.340 97.195 148.385 ;
        RECT 99.425 148.340 99.715 148.385 ;
        RECT 95.715 148.200 99.715 148.340 ;
        RECT 101.810 148.340 101.950 148.835 ;
        RECT 109.080 148.820 109.400 148.880 ;
        RECT 118.740 148.820 119.060 148.880 ;
        RECT 121.960 148.820 122.280 148.880 ;
        RECT 111.840 148.680 112.160 148.740 ;
        RECT 130.280 148.680 130.570 148.725 ;
        RECT 132.380 148.680 132.670 148.725 ;
        RECT 133.950 148.680 134.240 148.725 ;
        RECT 111.840 148.540 116.210 148.680 ;
        RECT 111.840 148.480 112.160 148.540 ;
        RECT 106.795 148.340 107.085 148.385 ;
        RECT 115.075 148.340 115.365 148.385 ;
        RECT 101.810 148.200 107.085 148.340 ;
        RECT 95.715 148.155 96.005 148.200 ;
        RECT 96.905 148.155 97.195 148.200 ;
        RECT 99.425 148.155 99.715 148.200 ;
        RECT 106.795 148.155 107.085 148.200 ;
        RECT 112.390 148.200 115.365 148.340 ;
        RECT 70.455 148.000 70.745 148.045 ;
        RECT 67.680 147.860 70.745 148.000 ;
        RECT 67.680 147.800 68.000 147.860 ;
        RECT 70.455 147.815 70.745 147.860 ;
        RECT 71.375 147.815 71.665 148.045 ;
        RECT 84.760 147.815 85.050 148.045 ;
        RECT 86.080 148.000 86.400 148.060 ;
        RECT 86.555 148.000 86.845 148.045 ;
        RECT 92.520 148.000 92.840 148.060 ;
        RECT 94.835 148.000 95.125 148.045 ;
        RECT 86.080 147.860 95.125 148.000 ;
        RECT 53.740 147.660 54.030 147.705 ;
        RECT 52.130 147.520 54.030 147.660 ;
        RECT 45.615 147.475 45.905 147.520 ;
        RECT 49.755 147.475 50.045 147.520 ;
        RECT 53.740 147.475 54.030 147.520 ;
        RECT 64.475 147.660 64.765 147.705 ;
        RECT 66.850 147.660 66.990 147.800 ;
        RECT 64.475 147.520 66.990 147.660 ;
        RECT 70.900 147.660 71.220 147.720 ;
        RECT 83.780 147.660 84.100 147.720 ;
        RECT 70.900 147.520 84.100 147.660 ;
        RECT 64.475 147.475 64.765 147.520 ;
        RECT 70.900 147.460 71.220 147.520 ;
        RECT 83.780 147.460 84.100 147.520 ;
        RECT 84.835 147.380 84.975 147.815 ;
        RECT 86.080 147.800 86.400 147.860 ;
        RECT 86.555 147.815 86.845 147.860 ;
        RECT 92.520 147.800 92.840 147.860 ;
        RECT 94.835 147.815 95.125 147.860 ;
        RECT 100.340 148.000 100.660 148.060 ;
        RECT 112.390 148.045 112.530 148.200 ;
        RECT 115.075 148.155 115.365 148.200 ;
        RECT 110.475 148.000 110.765 148.045 ;
        RECT 100.340 147.860 110.765 148.000 ;
        RECT 100.340 147.800 100.660 147.860 ;
        RECT 110.475 147.815 110.765 147.860 ;
        RECT 111.395 147.815 111.685 148.045 ;
        RECT 112.315 147.815 112.605 148.045 ;
        RECT 112.775 147.815 113.065 148.045 ;
        RECT 87.890 147.660 88.180 147.705 ;
        RECT 91.140 147.660 91.460 147.720 ;
        RECT 87.890 147.520 91.460 147.660 ;
        RECT 87.890 147.475 88.180 147.520 ;
        RECT 91.140 147.460 91.460 147.520 ;
        RECT 96.170 147.660 96.460 147.705 ;
        RECT 100.800 147.660 101.120 147.720 ;
        RECT 96.170 147.520 101.120 147.660 ;
        RECT 96.170 147.475 96.460 147.520 ;
        RECT 100.800 147.460 101.120 147.520 ;
        RECT 110.000 147.660 110.320 147.720 ;
        RECT 111.470 147.660 111.610 147.815 ;
        RECT 110.000 147.520 111.610 147.660 ;
        RECT 110.000 147.460 110.320 147.520 ;
        RECT 30.050 147.180 33.870 147.320 ;
        RECT 35.020 147.120 35.340 147.380 ;
        RECT 35.940 147.120 36.260 147.380 ;
        RECT 39.635 147.320 39.925 147.365 ;
        RECT 40.080 147.320 40.400 147.380 ;
        RECT 39.635 147.180 40.400 147.320 ;
        RECT 39.635 147.135 39.925 147.180 ;
        RECT 40.080 147.120 40.400 147.180 ;
        RECT 43.775 147.320 44.065 147.365 ;
        RECT 45.140 147.320 45.460 147.380 ;
        RECT 43.775 147.180 45.460 147.320 ;
        RECT 43.775 147.135 44.065 147.180 ;
        RECT 45.140 147.120 45.460 147.180 ;
        RECT 50.805 147.320 51.095 147.365 ;
        RECT 54.340 147.320 54.660 147.380 ;
        RECT 50.805 147.180 54.660 147.320 ;
        RECT 50.805 147.135 51.095 147.180 ;
        RECT 54.340 147.120 54.660 147.180 ;
        RECT 55.720 147.320 56.040 147.380 ;
        RECT 59.415 147.320 59.705 147.365 ;
        RECT 55.720 147.180 59.705 147.320 ;
        RECT 55.720 147.120 56.040 147.180 ;
        RECT 59.415 147.135 59.705 147.180 ;
        RECT 65.525 147.320 65.815 147.365 ;
        RECT 69.520 147.320 69.840 147.380 ;
        RECT 65.525 147.180 69.840 147.320 ;
        RECT 65.525 147.135 65.815 147.180 ;
        RECT 69.520 147.120 69.840 147.180 ;
        RECT 74.135 147.320 74.425 147.365 ;
        RECT 75.500 147.320 75.820 147.380 ;
        RECT 74.135 147.180 75.820 147.320 ;
        RECT 74.135 147.135 74.425 147.180 ;
        RECT 75.500 147.120 75.820 147.180 ;
        RECT 79.195 147.320 79.485 147.365 ;
        RECT 84.240 147.320 84.560 147.380 ;
        RECT 79.195 147.180 84.560 147.320 ;
        RECT 79.195 147.135 79.485 147.180 ;
        RECT 84.240 147.120 84.560 147.180 ;
        RECT 84.700 147.120 85.020 147.380 ;
        RECT 102.640 147.320 102.960 147.380 ;
        RECT 104.035 147.320 104.325 147.365 ;
        RECT 102.640 147.180 104.325 147.320 ;
        RECT 102.640 147.120 102.960 147.180 ;
        RECT 104.035 147.135 104.325 147.180 ;
        RECT 106.780 147.320 107.100 147.380 ;
        RECT 107.715 147.320 108.005 147.365 ;
        RECT 106.780 147.180 108.005 147.320 ;
        RECT 106.780 147.120 107.100 147.180 ;
        RECT 107.715 147.135 108.005 147.180 ;
        RECT 111.380 147.320 111.700 147.380 ;
        RECT 112.850 147.320 112.990 147.815 ;
        RECT 113.220 147.800 113.540 148.060 ;
        RECT 116.070 148.045 116.210 148.540 ;
        RECT 130.280 148.540 134.240 148.680 ;
        RECT 130.280 148.495 130.570 148.540 ;
        RECT 132.380 148.495 132.670 148.540 ;
        RECT 133.950 148.495 134.240 148.540 ;
        RECT 130.675 148.340 130.965 148.385 ;
        RECT 131.865 148.340 132.155 148.385 ;
        RECT 134.385 148.340 134.675 148.385 ;
        RECT 130.675 148.200 134.675 148.340 ;
        RECT 130.675 148.155 130.965 148.200 ;
        RECT 131.865 148.155 132.155 148.200 ;
        RECT 134.385 148.155 134.675 148.200 ;
        RECT 115.995 148.000 116.285 148.045 ;
        RECT 124.720 148.000 125.040 148.060 ;
        RECT 115.995 147.860 125.040 148.000 ;
        RECT 115.995 147.815 116.285 147.860 ;
        RECT 124.720 147.800 125.040 147.860 ;
        RECT 129.780 147.800 130.100 148.060 ;
        RECT 113.310 147.660 113.450 147.800 ;
        RECT 113.310 147.520 116.670 147.660 ;
        RECT 111.380 147.180 112.990 147.320 ;
        RECT 111.380 147.120 111.700 147.180 ;
        RECT 114.600 147.120 114.920 147.380 ;
        RECT 116.530 147.320 116.670 147.520 ;
        RECT 116.900 147.460 117.220 147.720 ;
        RECT 129.320 147.660 129.640 147.720 ;
        RECT 131.020 147.660 131.310 147.705 ;
        RECT 129.320 147.520 131.310 147.660 ;
        RECT 129.320 147.460 129.640 147.520 ;
        RECT 131.020 147.475 131.310 147.520 ;
        RECT 123.800 147.320 124.120 147.380 ;
        RECT 127.940 147.320 128.260 147.380 ;
        RECT 116.530 147.180 128.260 147.320 ;
        RECT 123.800 147.120 124.120 147.180 ;
        RECT 127.940 147.120 128.260 147.180 ;
        RECT 136.220 147.320 136.540 147.380 ;
        RECT 136.695 147.320 136.985 147.365 ;
        RECT 136.220 147.180 136.985 147.320 ;
        RECT 136.220 147.120 136.540 147.180 ;
        RECT 136.695 147.135 136.985 147.180 ;
        RECT 13.330 146.500 138.910 146.980 ;
        RECT 8.340 146.300 8.660 146.360 ;
        RECT 8.340 146.160 74.350 146.300 ;
        RECT 8.340 146.100 8.660 146.160 ;
        RECT 23.535 145.960 23.825 146.005 ;
        RECT 34.100 145.960 34.420 146.020 ;
        RECT 36.415 145.960 36.705 146.005 ;
        RECT 39.160 145.960 39.480 146.020 ;
        RECT 39.635 145.960 39.925 146.005 ;
        RECT 23.535 145.820 24.670 145.960 ;
        RECT 23.535 145.775 23.825 145.820 ;
        RECT 15.700 145.420 16.020 145.680 ;
        RECT 17.080 145.665 17.400 145.680 ;
        RECT 17.050 145.620 17.400 145.665 ;
        RECT 16.885 145.480 17.400 145.620 ;
        RECT 17.050 145.435 17.400 145.480 ;
        RECT 17.080 145.420 17.400 145.435 ;
        RECT 22.600 145.620 22.920 145.680 ;
        RECT 23.075 145.620 23.365 145.665 ;
        RECT 22.600 145.480 23.365 145.620 ;
        RECT 22.600 145.420 22.920 145.480 ;
        RECT 23.075 145.435 23.365 145.480 ;
        RECT 23.980 145.420 24.300 145.680 ;
        RECT 24.530 145.665 24.670 145.820 ;
        RECT 34.100 145.820 35.250 145.960 ;
        RECT 34.100 145.760 34.420 145.820 ;
        RECT 24.455 145.435 24.745 145.665 ;
        RECT 25.375 145.620 25.665 145.665 ;
        RECT 26.740 145.620 27.060 145.680 ;
        RECT 25.375 145.480 27.060 145.620 ;
        RECT 25.375 145.435 25.665 145.480 ;
        RECT 16.595 145.280 16.885 145.325 ;
        RECT 17.785 145.280 18.075 145.325 ;
        RECT 20.305 145.280 20.595 145.325 ;
        RECT 16.595 145.140 20.595 145.280 ;
        RECT 16.595 145.095 16.885 145.140 ;
        RECT 17.785 145.095 18.075 145.140 ;
        RECT 20.305 145.095 20.595 145.140 ;
        RECT 22.140 145.280 22.460 145.340 ;
        RECT 23.520 145.280 23.840 145.340 ;
        RECT 25.450 145.280 25.590 145.435 ;
        RECT 26.740 145.420 27.060 145.480 ;
        RECT 31.800 145.620 32.120 145.680 ;
        RECT 32.275 145.620 32.565 145.665 ;
        RECT 31.800 145.480 32.565 145.620 ;
        RECT 31.800 145.420 32.120 145.480 ;
        RECT 32.275 145.435 32.565 145.480 ;
        RECT 33.655 145.435 33.945 145.665 ;
        RECT 22.140 145.140 22.830 145.280 ;
        RECT 22.140 145.080 22.460 145.140 ;
        RECT 22.690 144.985 22.830 145.140 ;
        RECT 23.520 145.140 25.590 145.280 ;
        RECT 23.520 145.080 23.840 145.140 ;
        RECT 16.200 144.940 16.490 144.985 ;
        RECT 18.300 144.940 18.590 144.985 ;
        RECT 19.870 144.940 20.160 144.985 ;
        RECT 16.200 144.800 20.160 144.940 ;
        RECT 16.200 144.755 16.490 144.800 ;
        RECT 18.300 144.755 18.590 144.800 ;
        RECT 19.870 144.755 20.160 144.800 ;
        RECT 22.615 144.755 22.905 144.985 ;
        RECT 24.440 144.400 24.760 144.660 ;
        RECT 32.720 144.400 33.040 144.660 ;
        RECT 33.730 144.600 33.870 145.435 ;
        RECT 34.560 145.420 34.880 145.680 ;
        RECT 35.110 145.665 35.250 145.820 ;
        RECT 36.415 145.820 39.925 145.960 ;
        RECT 36.415 145.775 36.705 145.820 ;
        RECT 39.160 145.760 39.480 145.820 ;
        RECT 39.635 145.775 39.925 145.820 ;
        RECT 40.080 145.960 40.400 146.020 ;
        RECT 40.635 145.960 40.925 146.005 ;
        RECT 40.080 145.820 40.925 145.960 ;
        RECT 40.080 145.760 40.400 145.820 ;
        RECT 40.635 145.775 40.925 145.820 ;
        RECT 41.090 145.820 46.750 145.960 ;
        RECT 35.035 145.435 35.325 145.665 ;
        RECT 35.480 145.420 35.800 145.680 ;
        RECT 36.860 145.420 37.180 145.680 ;
        RECT 37.335 145.435 37.625 145.665 ;
        RECT 37.780 145.620 38.100 145.680 ;
        RECT 41.090 145.620 41.230 145.820 ;
        RECT 46.610 145.680 46.750 145.820 ;
        RECT 47.900 145.760 48.220 146.020 ;
        RECT 49.280 145.760 49.600 146.020 ;
        RECT 51.580 145.960 51.900 146.020 ;
        RECT 50.750 145.820 51.900 145.960 ;
        RECT 43.315 145.620 43.605 145.665 ;
        RECT 37.780 145.480 41.230 145.620 ;
        RECT 41.550 145.480 43.605 145.620 ;
        RECT 34.115 145.280 34.405 145.325 ;
        RECT 37.410 145.280 37.550 145.435 ;
        RECT 37.780 145.420 38.100 145.480 ;
        RECT 41.000 145.280 41.320 145.340 ;
        RECT 34.115 145.140 37.550 145.280 ;
        RECT 38.330 145.140 41.320 145.280 ;
        RECT 34.115 145.095 34.405 145.140 ;
        RECT 34.560 144.940 34.880 145.000 ;
        RECT 35.940 144.940 36.260 145.000 ;
        RECT 37.780 144.940 38.100 145.000 ;
        RECT 38.330 144.985 38.470 145.140 ;
        RECT 41.000 145.080 41.320 145.140 ;
        RECT 41.550 144.985 41.690 145.480 ;
        RECT 43.315 145.435 43.605 145.480 ;
        RECT 44.695 145.620 44.985 145.665 ;
        RECT 45.140 145.620 45.460 145.680 ;
        RECT 44.695 145.480 45.460 145.620 ;
        RECT 44.695 145.435 44.985 145.480 ;
        RECT 45.140 145.420 45.460 145.480 ;
        RECT 46.060 145.420 46.380 145.680 ;
        RECT 46.520 145.620 46.840 145.680 ;
        RECT 46.520 145.480 49.050 145.620 ;
        RECT 49.290 145.545 49.580 145.760 ;
        RECT 50.750 145.665 50.890 145.820 ;
        RECT 51.580 145.760 51.900 145.820 ;
        RECT 54.800 145.760 55.120 146.020 ;
        RECT 55.260 145.960 55.580 146.020 ;
        RECT 55.815 145.960 56.105 146.005 ;
        RECT 57.575 145.960 57.865 146.005 ;
        RECT 55.260 145.820 56.105 145.960 ;
        RECT 55.260 145.760 55.580 145.820 ;
        RECT 55.815 145.775 56.105 145.820 ;
        RECT 56.270 145.820 57.865 145.960 ;
        RECT 46.520 145.420 46.840 145.480 ;
        RECT 47.900 145.080 48.220 145.340 ;
        RECT 34.560 144.800 36.260 144.940 ;
        RECT 34.560 144.740 34.880 144.800 ;
        RECT 35.940 144.740 36.260 144.800 ;
        RECT 36.490 144.800 38.100 144.940 ;
        RECT 36.490 144.600 36.630 144.800 ;
        RECT 37.780 144.740 38.100 144.800 ;
        RECT 38.255 144.755 38.545 144.985 ;
        RECT 41.475 144.755 41.765 144.985 ;
        RECT 44.220 144.940 44.540 145.000 ;
        RECT 48.360 144.940 48.680 145.000 ;
        RECT 44.220 144.800 48.680 144.940 ;
        RECT 48.910 144.940 49.050 145.480 ;
        RECT 49.755 145.425 50.045 145.655 ;
        RECT 50.675 145.435 50.965 145.665 ;
        RECT 51.165 145.435 51.455 145.665 ;
        RECT 49.830 145.280 49.970 145.425 ;
        RECT 50.200 145.280 50.520 145.340 ;
        RECT 49.830 145.140 50.520 145.280 ;
        RECT 50.200 145.080 50.520 145.140 ;
        RECT 50.750 144.940 50.890 145.435 ;
        RECT 51.240 145.280 51.380 145.435 ;
        RECT 52.040 145.420 52.360 145.680 ;
        RECT 52.515 145.620 52.805 145.665 ;
        RECT 52.515 145.435 52.810 145.620 ;
        RECT 52.975 145.610 53.265 145.665 ;
        RECT 53.420 145.610 53.740 145.680 ;
        RECT 52.975 145.470 53.740 145.610 ;
        RECT 52.975 145.435 53.265 145.470 ;
        RECT 51.240 145.140 51.395 145.280 ;
        RECT 48.910 144.800 50.890 144.940 ;
        RECT 44.220 144.740 44.540 144.800 ;
        RECT 48.360 144.740 48.680 144.800 ;
        RECT 33.730 144.460 36.630 144.600 ;
        RECT 36.860 144.600 37.180 144.660 ;
        RECT 40.555 144.600 40.845 144.645 ;
        RECT 36.860 144.460 40.845 144.600 ;
        RECT 36.860 144.400 37.180 144.460 ;
        RECT 40.555 144.415 40.845 144.460 ;
        RECT 46.980 144.600 47.300 144.660 ;
        RECT 48.835 144.600 49.125 144.645 ;
        RECT 46.980 144.460 49.125 144.600 ;
        RECT 46.980 144.400 47.300 144.460 ;
        RECT 48.835 144.415 49.125 144.460 ;
        RECT 49.280 144.600 49.600 144.660 ;
        RECT 50.215 144.600 50.505 144.645 ;
        RECT 49.280 144.460 50.505 144.600 ;
        RECT 51.255 144.600 51.395 145.140 ;
        RECT 52.670 145.240 52.810 145.435 ;
        RECT 53.420 145.420 53.740 145.470 ;
        RECT 54.340 145.620 54.660 145.680 ;
        RECT 56.270 145.620 56.410 145.820 ;
        RECT 57.575 145.775 57.865 145.820 ;
        RECT 68.600 145.760 68.920 146.020 ;
        RECT 74.210 146.005 74.350 146.160 ;
        RECT 81.480 146.100 81.800 146.360 ;
        RECT 87.000 146.300 87.320 146.360 ;
        RECT 88.840 146.300 89.160 146.360 ;
        RECT 90.235 146.300 90.525 146.345 ;
        RECT 87.000 146.160 90.525 146.300 ;
        RECT 87.000 146.100 87.320 146.160 ;
        RECT 88.840 146.100 89.160 146.160 ;
        RECT 90.235 146.115 90.525 146.160 ;
        RECT 100.340 146.100 100.660 146.360 ;
        RECT 100.800 146.100 101.120 146.360 ;
        RECT 102.640 146.100 102.960 146.360 ;
        RECT 104.955 146.115 105.245 146.345 ;
        RECT 84.700 146.005 85.020 146.020 ;
        RECT 69.995 145.775 70.285 146.005 ;
        RECT 71.075 145.960 71.365 146.005 ;
        RECT 72.755 145.960 73.045 146.005 ;
        RECT 71.075 145.820 73.045 145.960 ;
        RECT 71.075 145.775 71.365 145.820 ;
        RECT 72.755 145.775 73.045 145.820 ;
        RECT 74.135 145.775 74.425 146.005 ;
        RECT 84.560 145.775 85.020 146.005 ;
        RECT 94.790 145.960 95.080 146.005 ;
        RECT 105.030 145.960 105.170 146.115 ;
        RECT 106.780 146.100 107.100 146.360 ;
        RECT 108.160 146.300 108.480 146.360 ;
        RECT 113.220 146.300 113.540 146.360 ;
        RECT 108.160 146.160 113.540 146.300 ;
        RECT 108.160 146.100 108.480 146.160 ;
        RECT 113.220 146.100 113.540 146.160 ;
        RECT 114.600 146.300 114.920 146.360 ;
        RECT 123.815 146.300 124.105 146.345 ;
        RECT 124.720 146.300 125.040 146.360 ;
        RECT 114.600 146.160 118.280 146.300 ;
        RECT 114.600 146.100 114.920 146.160 ;
        RECT 118.140 146.005 118.280 146.160 ;
        RECT 123.815 146.160 125.040 146.300 ;
        RECT 123.815 146.115 124.105 146.160 ;
        RECT 124.720 146.100 125.040 146.160 ;
        RECT 129.320 146.100 129.640 146.360 ;
        RECT 134.840 146.100 135.160 146.360 ;
        RECT 136.680 146.100 137.000 146.360 ;
        RECT 94.790 145.820 105.170 145.960 ;
        RECT 109.170 145.820 112.530 145.960 ;
        RECT 94.790 145.775 95.080 145.820 ;
        RECT 54.340 145.480 56.410 145.620 ;
        RECT 54.340 145.420 54.660 145.480 ;
        RECT 57.115 145.435 57.405 145.665 ;
        RECT 57.190 145.280 57.330 145.435 ;
        RECT 58.020 145.420 58.340 145.680 ;
        RECT 66.760 145.420 67.080 145.680 ;
        RECT 70.070 145.620 70.210 145.775 ;
        RECT 84.700 145.760 85.020 145.775 ;
        RECT 71.820 145.620 72.140 145.680 ;
        RECT 70.070 145.480 72.140 145.620 ;
        RECT 71.820 145.420 72.140 145.480 ;
        RECT 73.200 145.420 73.520 145.680 ;
        RECT 83.320 145.420 83.640 145.680 ;
        RECT 92.060 145.620 92.380 145.680 ;
        RECT 83.870 145.480 92.380 145.620 ;
        RECT 70.900 145.280 71.220 145.340 ;
        RECT 75.960 145.280 76.280 145.340 ;
        RECT 83.870 145.280 84.010 145.480 ;
        RECT 92.060 145.420 92.380 145.480 ;
        RECT 92.520 145.620 92.840 145.680 ;
        RECT 93.455 145.620 93.745 145.665 ;
        RECT 92.520 145.480 93.745 145.620 ;
        RECT 92.520 145.420 92.840 145.480 ;
        RECT 93.455 145.435 93.745 145.480 ;
        RECT 103.115 145.620 103.405 145.665 ;
        RECT 105.400 145.620 105.720 145.680 ;
        RECT 103.115 145.480 105.720 145.620 ;
        RECT 103.115 145.435 103.405 145.480 ;
        RECT 105.400 145.420 105.720 145.480 ;
        RECT 107.255 145.620 107.545 145.665 ;
        RECT 108.620 145.620 108.940 145.680 ;
        RECT 109.170 145.665 109.310 145.820 ;
        RECT 112.390 145.680 112.530 145.820 ;
        RECT 118.140 145.775 118.430 146.005 ;
        RECT 126.560 145.960 126.880 146.020 ;
        RECT 130.240 145.960 130.560 146.020 ;
        RECT 126.560 145.820 127.710 145.960 ;
        RECT 126.560 145.760 126.880 145.820 ;
        RECT 107.255 145.480 108.940 145.620 ;
        RECT 107.255 145.435 107.545 145.480 ;
        RECT 108.620 145.420 108.940 145.480 ;
        RECT 109.095 145.435 109.385 145.665 ;
        RECT 109.540 145.620 109.860 145.680 ;
        RECT 110.375 145.620 110.665 145.665 ;
        RECT 109.540 145.480 110.665 145.620 ;
        RECT 109.540 145.420 109.860 145.480 ;
        RECT 110.375 145.435 110.665 145.480 ;
        RECT 112.300 145.620 112.620 145.680 ;
        RECT 115.980 145.620 116.300 145.680 ;
        RECT 116.915 145.620 117.205 145.665 ;
        RECT 112.300 145.480 117.205 145.620 ;
        RECT 112.300 145.420 112.620 145.480 ;
        RECT 115.980 145.420 116.300 145.480 ;
        RECT 116.915 145.435 117.205 145.480 ;
        RECT 117.360 145.420 117.680 145.680 ;
        RECT 127.570 145.665 127.710 145.820 ;
        RECT 128.030 145.820 130.560 145.960 ;
        RECT 128.030 145.680 128.170 145.820 ;
        RECT 130.240 145.760 130.560 145.820 ;
        RECT 130.715 145.960 131.005 146.005 ;
        RECT 136.220 145.960 136.540 146.020 ;
        RECT 130.715 145.820 136.540 145.960 ;
        RECT 130.715 145.775 131.005 145.820 ;
        RECT 136.220 145.760 136.540 145.820 ;
        RECT 126.115 145.435 126.405 145.665 ;
        RECT 127.035 145.435 127.325 145.665 ;
        RECT 127.495 145.435 127.785 145.665 ;
        RECT 53.815 145.240 57.330 145.280 ;
        RECT 52.670 145.140 57.330 145.240 ;
        RECT 69.610 145.140 71.220 145.280 ;
        RECT 52.670 145.100 53.955 145.140 ;
        RECT 56.730 144.985 56.870 145.140 ;
        RECT 69.610 144.985 69.750 145.140 ;
        RECT 70.900 145.080 71.220 145.140 ;
        RECT 71.910 145.140 84.010 145.280 ;
        RECT 84.215 145.280 84.505 145.325 ;
        RECT 85.405 145.280 85.695 145.325 ;
        RECT 87.925 145.280 88.215 145.325 ;
        RECT 84.215 145.140 88.215 145.280 ;
        RECT 71.910 144.985 72.050 145.140 ;
        RECT 75.960 145.080 76.280 145.140 ;
        RECT 84.215 145.095 84.505 145.140 ;
        RECT 85.405 145.095 85.695 145.140 ;
        RECT 87.925 145.095 88.215 145.140 ;
        RECT 94.335 145.280 94.625 145.325 ;
        RECT 95.525 145.280 95.815 145.325 ;
        RECT 98.045 145.280 98.335 145.325 ;
        RECT 94.335 145.140 98.335 145.280 ;
        RECT 94.335 145.095 94.625 145.140 ;
        RECT 95.525 145.095 95.815 145.140 ;
        RECT 98.045 145.095 98.335 145.140 ;
        RECT 103.575 145.095 103.865 145.325 ;
        RECT 107.715 145.095 108.005 145.325 ;
        RECT 109.975 145.280 110.265 145.325 ;
        RECT 111.165 145.280 111.455 145.325 ;
        RECT 113.685 145.280 113.975 145.325 ;
        RECT 117.450 145.280 117.590 145.420 ;
        RECT 109.975 145.140 113.975 145.280 ;
        RECT 109.975 145.095 110.265 145.140 ;
        RECT 111.165 145.095 111.455 145.140 ;
        RECT 113.685 145.095 113.975 145.140 ;
        RECT 114.690 145.140 117.590 145.280 ;
        RECT 117.795 145.280 118.085 145.325 ;
        RECT 118.985 145.280 119.275 145.325 ;
        RECT 121.505 145.280 121.795 145.325 ;
        RECT 117.795 145.140 121.795 145.280 ;
        RECT 56.655 144.940 56.945 144.985 ;
        RECT 56.655 144.800 57.055 144.940 ;
        RECT 56.655 144.755 56.945 144.800 ;
        RECT 69.535 144.755 69.825 144.985 ;
        RECT 71.835 144.755 72.125 144.985 ;
        RECT 83.820 144.940 84.110 144.985 ;
        RECT 85.920 144.940 86.210 144.985 ;
        RECT 87.490 144.940 87.780 144.985 ;
        RECT 83.820 144.800 87.780 144.940 ;
        RECT 83.820 144.755 84.110 144.800 ;
        RECT 85.920 144.755 86.210 144.800 ;
        RECT 87.490 144.755 87.780 144.800 ;
        RECT 93.940 144.940 94.230 144.985 ;
        RECT 96.040 144.940 96.330 144.985 ;
        RECT 97.610 144.940 97.900 144.985 ;
        RECT 93.940 144.800 97.900 144.940 ;
        RECT 93.940 144.755 94.230 144.800 ;
        RECT 96.040 144.755 96.330 144.800 ;
        RECT 97.610 144.755 97.900 144.800 ;
        RECT 99.420 144.940 99.740 145.000 ;
        RECT 103.650 144.940 103.790 145.095 ;
        RECT 107.790 144.940 107.930 145.095 ;
        RECT 99.420 144.800 107.930 144.940 ;
        RECT 109.580 144.940 109.870 144.985 ;
        RECT 111.680 144.940 111.970 144.985 ;
        RECT 113.250 144.940 113.540 144.985 ;
        RECT 109.580 144.800 113.540 144.940 ;
        RECT 99.420 144.740 99.740 144.800 ;
        RECT 109.580 144.755 109.870 144.800 ;
        RECT 111.680 144.755 111.970 144.800 ;
        RECT 113.250 144.755 113.540 144.800 ;
        RECT 52.960 144.600 53.280 144.660 ;
        RECT 51.255 144.460 53.280 144.600 ;
        RECT 49.280 144.400 49.600 144.460 ;
        RECT 50.215 144.415 50.505 144.460 ;
        RECT 52.960 144.400 53.280 144.460 ;
        RECT 53.880 144.600 54.200 144.660 ;
        RECT 54.355 144.600 54.645 144.645 ;
        RECT 53.880 144.460 54.645 144.600 ;
        RECT 53.880 144.400 54.200 144.460 ;
        RECT 54.355 144.415 54.645 144.460 ;
        RECT 55.720 144.400 56.040 144.660 ;
        RECT 67.220 144.600 67.540 144.660 ;
        RECT 68.140 144.600 68.460 144.660 ;
        RECT 68.615 144.600 68.905 144.645 ;
        RECT 67.220 144.460 68.905 144.600 ;
        RECT 67.220 144.400 67.540 144.460 ;
        RECT 68.140 144.400 68.460 144.460 ;
        RECT 68.615 144.415 68.905 144.460 ;
        RECT 69.980 144.600 70.300 144.660 ;
        RECT 70.915 144.600 71.205 144.645 ;
        RECT 69.980 144.460 71.205 144.600 ;
        RECT 69.980 144.400 70.300 144.460 ;
        RECT 70.915 144.415 71.205 144.460 ;
        RECT 110.000 144.600 110.320 144.660 ;
        RECT 114.690 144.600 114.830 145.140 ;
        RECT 117.795 145.095 118.085 145.140 ;
        RECT 118.985 145.095 119.275 145.140 ;
        RECT 121.505 145.095 121.795 145.140 ;
        RECT 115.060 144.940 115.380 145.000 ;
        RECT 115.995 144.940 116.285 144.985 ;
        RECT 116.440 144.940 116.760 145.000 ;
        RECT 115.060 144.800 116.760 144.940 ;
        RECT 115.060 144.740 115.380 144.800 ;
        RECT 115.995 144.755 116.285 144.800 ;
        RECT 116.440 144.740 116.760 144.800 ;
        RECT 117.400 144.940 117.690 144.985 ;
        RECT 119.500 144.940 119.790 144.985 ;
        RECT 121.070 144.940 121.360 144.985 ;
        RECT 126.190 144.940 126.330 145.435 ;
        RECT 127.110 145.280 127.250 145.435 ;
        RECT 127.940 145.420 128.260 145.680 ;
        RECT 128.400 145.620 128.720 145.680 ;
        RECT 129.795 145.620 130.085 145.665 ;
        RECT 128.400 145.480 130.085 145.620 ;
        RECT 128.400 145.420 128.720 145.480 ;
        RECT 129.795 145.435 130.085 145.480 ;
        RECT 133.920 145.420 134.240 145.680 ;
        RECT 135.775 145.435 136.065 145.665 ;
        RECT 131.635 145.280 131.925 145.325 ;
        RECT 127.110 145.140 131.925 145.280 ;
        RECT 131.635 145.095 131.925 145.140 ;
        RECT 117.400 144.800 121.360 144.940 ;
        RECT 117.400 144.755 117.690 144.800 ;
        RECT 119.500 144.755 119.790 144.800 ;
        RECT 121.070 144.755 121.360 144.800 ;
        RECT 122.050 144.800 126.330 144.940 ;
        RECT 110.000 144.460 114.830 144.600 ;
        RECT 115.520 144.600 115.840 144.660 ;
        RECT 122.050 144.600 122.190 144.800 ;
        RECT 115.520 144.460 122.190 144.600 ;
        RECT 122.420 144.600 122.740 144.660 ;
        RECT 135.850 144.600 135.990 145.435 ;
        RECT 122.420 144.460 135.990 144.600 ;
        RECT 110.000 144.400 110.320 144.460 ;
        RECT 115.520 144.400 115.840 144.460 ;
        RECT 122.420 144.400 122.740 144.460 ;
        RECT 13.330 143.780 138.910 144.260 ;
        RECT 18.460 143.380 18.780 143.640 ;
        RECT 19.395 143.580 19.685 143.625 ;
        RECT 20.760 143.580 21.080 143.640 ;
        RECT 19.395 143.440 21.080 143.580 ;
        RECT 19.395 143.395 19.685 143.440 ;
        RECT 20.760 143.380 21.080 143.440 ;
        RECT 33.655 143.580 33.945 143.625 ;
        RECT 34.100 143.580 34.420 143.640 ;
        RECT 33.655 143.440 34.420 143.580 ;
        RECT 33.655 143.395 33.945 143.440 ;
        RECT 34.100 143.380 34.420 143.440 ;
        RECT 39.160 143.380 39.480 143.640 ;
        RECT 42.840 143.580 43.160 143.640 ;
        RECT 43.315 143.580 43.605 143.625 ;
        RECT 42.840 143.440 43.605 143.580 ;
        RECT 42.840 143.380 43.160 143.440 ;
        RECT 43.315 143.395 43.605 143.440 ;
        RECT 45.140 143.380 45.460 143.640 ;
        RECT 47.900 143.580 48.220 143.640 ;
        RECT 48.835 143.580 49.125 143.625 ;
        RECT 47.900 143.440 49.125 143.580 ;
        RECT 47.900 143.380 48.220 143.440 ;
        RECT 48.835 143.395 49.125 143.440 ;
        RECT 51.135 143.580 51.425 143.625 ;
        RECT 51.580 143.580 51.900 143.640 ;
        RECT 51.135 143.440 51.900 143.580 ;
        RECT 51.135 143.395 51.425 143.440 ;
        RECT 51.580 143.380 51.900 143.440 ;
        RECT 53.895 143.580 54.185 143.625 ;
        RECT 58.020 143.580 58.340 143.640 ;
        RECT 53.895 143.440 58.340 143.580 ;
        RECT 53.895 143.395 54.185 143.440 ;
        RECT 58.020 143.380 58.340 143.440 ;
        RECT 77.355 143.580 77.645 143.625 ;
        RECT 77.800 143.580 78.120 143.640 ;
        RECT 77.355 143.440 78.120 143.580 ;
        RECT 77.355 143.395 77.645 143.440 ;
        RECT 77.800 143.380 78.120 143.440 ;
        RECT 84.700 143.580 85.020 143.640 ;
        RECT 85.635 143.580 85.925 143.625 ;
        RECT 84.700 143.440 85.925 143.580 ;
        RECT 84.700 143.380 85.020 143.440 ;
        RECT 85.635 143.395 85.925 143.440 ;
        RECT 98.960 143.580 99.280 143.640 ;
        RECT 100.355 143.580 100.645 143.625 ;
        RECT 98.960 143.440 100.645 143.580 ;
        RECT 98.960 143.380 99.280 143.440 ;
        RECT 100.355 143.395 100.645 143.440 ;
        RECT 108.635 143.580 108.925 143.625 ;
        RECT 109.540 143.580 109.860 143.640 ;
        RECT 108.635 143.440 109.860 143.580 ;
        RECT 108.635 143.395 108.925 143.440 ;
        RECT 35.020 143.040 35.340 143.300 ;
        RECT 35.495 143.240 35.785 143.285 ;
        RECT 38.700 143.240 39.020 143.300 ;
        RECT 35.495 143.100 39.020 143.240 ;
        RECT 35.495 143.055 35.785 143.100 ;
        RECT 38.700 143.040 39.020 143.100 ;
        RECT 42.395 143.240 42.685 143.285 ;
        RECT 93.940 143.240 94.230 143.285 ;
        RECT 96.040 143.240 96.330 143.285 ;
        RECT 97.610 143.240 97.900 143.285 ;
        RECT 42.395 143.100 49.970 143.240 ;
        RECT 42.395 143.055 42.685 143.100 ;
        RECT 45.950 142.900 46.240 142.945 ;
        RECT 49.280 142.900 49.600 142.960 ;
        RECT 36.030 142.760 38.470 142.900 ;
        RECT 36.030 142.620 36.170 142.760 ;
        RECT 32.720 142.560 33.040 142.620 ;
        RECT 34.575 142.560 34.865 142.605 ;
        RECT 32.720 142.420 34.865 142.560 ;
        RECT 32.720 142.360 33.040 142.420 ;
        RECT 34.575 142.375 34.865 142.420 ;
        RECT 35.940 142.360 36.260 142.620 ;
        RECT 36.400 142.560 36.720 142.620 ;
        RECT 38.330 142.605 38.470 142.760 ;
        RECT 45.950 142.760 49.600 142.900 ;
        RECT 45.950 142.715 46.240 142.760 ;
        RECT 49.280 142.700 49.600 142.760 ;
        RECT 36.875 142.560 37.165 142.605 ;
        RECT 37.335 142.560 37.625 142.605 ;
        RECT 36.400 142.420 37.625 142.560 ;
        RECT 36.400 142.360 36.720 142.420 ;
        RECT 36.875 142.375 37.165 142.420 ;
        RECT 37.335 142.375 37.625 142.420 ;
        RECT 38.255 142.375 38.545 142.605 ;
        RECT 41.920 142.560 42.240 142.620 ;
        RECT 43.315 142.560 43.605 142.605 ;
        RECT 41.920 142.420 43.605 142.560 ;
        RECT 41.920 142.360 42.240 142.420 ;
        RECT 43.315 142.375 43.605 142.420 ;
        RECT 43.775 142.375 44.065 142.605 ;
        RECT 45.140 142.560 45.460 142.620 ;
        RECT 46.535 142.560 46.825 142.605 ;
        RECT 45.140 142.420 46.825 142.560 ;
        RECT 20.315 142.220 20.605 142.265 ;
        RECT 21.220 142.220 21.540 142.280 ;
        RECT 20.315 142.080 21.540 142.220 ;
        RECT 20.315 142.035 20.605 142.080 ;
        RECT 21.220 142.020 21.540 142.080 ;
        RECT 19.315 141.880 19.605 141.925 ;
        RECT 24.440 141.880 24.760 141.940 ;
        RECT 19.315 141.740 24.760 141.880 ;
        RECT 43.850 141.880 43.990 142.375 ;
        RECT 45.140 142.360 45.460 142.420 ;
        RECT 46.535 142.375 46.825 142.420 ;
        RECT 46.980 142.360 47.300 142.620 ;
        RECT 48.360 142.560 48.680 142.620 ;
        RECT 49.830 142.605 49.970 143.100 ;
        RECT 93.940 143.100 97.900 143.240 ;
        RECT 93.940 143.055 94.230 143.100 ;
        RECT 96.040 143.055 96.330 143.100 ;
        RECT 97.610 143.055 97.900 143.100 ;
        RECT 53.420 142.900 53.740 142.960 ;
        RECT 51.670 142.760 53.740 142.900 ;
        RECT 51.670 142.605 51.810 142.760 ;
        RECT 53.420 142.700 53.740 142.760 ;
        RECT 74.580 142.900 74.900 142.960 ;
        RECT 82.415 142.900 82.705 142.945 ;
        RECT 74.580 142.760 82.705 142.900 ;
        RECT 74.580 142.700 74.900 142.760 ;
        RECT 82.415 142.715 82.705 142.760 ;
        RECT 47.530 142.420 48.680 142.560 ;
        RECT 44.695 142.220 44.985 142.265 ;
        RECT 47.530 142.220 47.670 142.420 ;
        RECT 48.360 142.360 48.680 142.420 ;
        RECT 49.755 142.375 50.045 142.605 ;
        RECT 50.215 142.375 50.505 142.605 ;
        RECT 51.595 142.375 51.885 142.605 ;
        RECT 52.515 142.560 52.805 142.605 ;
        RECT 55.260 142.560 55.580 142.620 ;
        RECT 52.515 142.420 55.580 142.560 ;
        RECT 52.515 142.375 52.805 142.420 ;
        RECT 44.695 142.080 47.670 142.220 ;
        RECT 48.820 142.220 49.140 142.280 ;
        RECT 50.290 142.220 50.430 142.375 ;
        RECT 55.260 142.360 55.580 142.420 ;
        RECT 69.075 142.375 69.365 142.605 ;
        RECT 48.820 142.080 50.430 142.220 ;
        RECT 51.120 142.220 51.440 142.280 ;
        RECT 53.895 142.220 54.185 142.265 ;
        RECT 55.720 142.220 56.040 142.280 ;
        RECT 51.120 142.080 56.040 142.220 ;
        RECT 69.150 142.220 69.290 142.375 ;
        RECT 69.980 142.360 70.300 142.620 ;
        RECT 75.500 142.360 75.820 142.620 ;
        RECT 82.490 142.560 82.630 142.715 ;
        RECT 88.840 142.700 89.160 142.960 ;
        RECT 92.520 142.900 92.840 142.960 ;
        RECT 93.455 142.900 93.745 142.945 ;
        RECT 92.520 142.760 93.745 142.900 ;
        RECT 92.520 142.700 92.840 142.760 ;
        RECT 93.455 142.715 93.745 142.760 ;
        RECT 94.335 142.900 94.625 142.945 ;
        RECT 95.525 142.900 95.815 142.945 ;
        RECT 98.045 142.900 98.335 142.945 ;
        RECT 94.335 142.760 98.335 142.900 ;
        RECT 100.430 142.900 100.570 143.395 ;
        RECT 109.540 143.380 109.860 143.440 ;
        RECT 111.840 143.380 112.160 143.640 ;
        RECT 113.220 143.580 113.540 143.640 ;
        RECT 115.520 143.580 115.840 143.640 ;
        RECT 113.220 143.440 115.840 143.580 ;
        RECT 113.220 143.380 113.540 143.440 ;
        RECT 115.520 143.380 115.840 143.440 ;
        RECT 117.360 143.580 117.680 143.640 ;
        RECT 117.360 143.440 118.280 143.580 ;
        RECT 117.360 143.380 117.680 143.440 ;
        RECT 107.240 143.240 107.560 143.300 ;
        RECT 111.930 143.240 112.070 143.380 ;
        RECT 107.240 143.100 112.070 143.240 ;
        RECT 112.800 143.240 113.090 143.285 ;
        RECT 114.900 143.240 115.190 143.285 ;
        RECT 116.470 143.240 116.760 143.285 ;
        RECT 112.800 143.100 116.760 143.240 ;
        RECT 107.240 143.040 107.560 143.100 ;
        RECT 112.800 143.055 113.090 143.100 ;
        RECT 114.900 143.055 115.190 143.100 ;
        RECT 116.470 143.055 116.760 143.100 ;
        RECT 106.795 142.900 107.085 142.945 ;
        RECT 100.430 142.760 107.085 142.900 ;
        RECT 94.335 142.715 94.625 142.760 ;
        RECT 95.525 142.715 95.815 142.760 ;
        RECT 98.045 142.715 98.335 142.760 ;
        RECT 106.795 142.715 107.085 142.760 ;
        RECT 112.300 142.700 112.620 142.960 ;
        RECT 113.195 142.900 113.485 142.945 ;
        RECT 114.385 142.900 114.675 142.945 ;
        RECT 116.905 142.900 117.195 142.945 ;
        RECT 113.195 142.760 117.195 142.900 ;
        RECT 113.195 142.715 113.485 142.760 ;
        RECT 114.385 142.715 114.675 142.760 ;
        RECT 116.905 142.715 117.195 142.760 ;
        RECT 98.960 142.560 99.280 142.620 ;
        RECT 82.490 142.420 99.280 142.560 ;
        RECT 98.960 142.360 99.280 142.420 ;
        RECT 109.080 142.560 109.400 142.620 ;
        RECT 110.015 142.560 110.305 142.605 ;
        RECT 109.080 142.420 110.305 142.560 ;
        RECT 109.080 142.360 109.400 142.420 ;
        RECT 110.015 142.375 110.305 142.420 ;
        RECT 110.460 142.360 110.780 142.620 ;
        RECT 110.935 142.375 111.225 142.605 ;
        RECT 111.855 142.560 112.145 142.605 ;
        RECT 115.520 142.560 115.840 142.620 ;
        RECT 111.855 142.420 115.840 142.560 ;
        RECT 118.140 142.560 118.280 143.440 ;
        RECT 123.800 143.240 124.120 143.300 ;
        RECT 128.400 143.240 128.720 143.300 ;
        RECT 123.800 143.100 128.720 143.240 ;
        RECT 123.800 143.040 124.120 143.100 ;
        RECT 128.400 143.040 128.720 143.100 ;
        RECT 130.280 143.240 130.570 143.285 ;
        RECT 132.380 143.240 132.670 143.285 ;
        RECT 133.950 143.240 134.240 143.285 ;
        RECT 130.280 143.100 134.240 143.240 ;
        RECT 130.280 143.055 130.570 143.100 ;
        RECT 132.380 143.055 132.670 143.100 ;
        RECT 133.950 143.055 134.240 143.100 ;
        RECT 125.195 142.900 125.485 142.945 ;
        RECT 130.675 142.900 130.965 142.945 ;
        RECT 131.865 142.900 132.155 142.945 ;
        RECT 134.385 142.900 134.675 142.945 ;
        RECT 125.195 142.760 126.790 142.900 ;
        RECT 125.195 142.715 125.485 142.760 ;
        RECT 124.720 142.560 125.040 142.620 ;
        RECT 126.650 142.605 126.790 142.760 ;
        RECT 130.675 142.760 134.675 142.900 ;
        RECT 130.675 142.715 130.965 142.760 ;
        RECT 131.865 142.715 132.155 142.760 ;
        RECT 134.385 142.715 134.675 142.760 ;
        RECT 125.655 142.560 125.945 142.605 ;
        RECT 118.140 142.420 125.945 142.560 ;
        RECT 111.855 142.375 112.145 142.420 ;
        RECT 72.740 142.220 73.060 142.280 ;
        RECT 69.150 142.080 73.060 142.220 ;
        RECT 44.695 142.035 44.985 142.080 ;
        RECT 48.820 142.020 49.140 142.080 ;
        RECT 51.120 142.020 51.440 142.080 ;
        RECT 53.895 142.035 54.185 142.080 ;
        RECT 55.720 142.020 56.040 142.080 ;
        RECT 72.740 142.020 73.060 142.080 ;
        RECT 75.055 142.220 75.345 142.265 ;
        RECT 79.180 142.220 79.500 142.280 ;
        RECT 75.055 142.080 79.500 142.220 ;
        RECT 75.055 142.035 75.345 142.080 ;
        RECT 79.180 142.020 79.500 142.080 ;
        RECT 83.335 142.220 83.625 142.265 ;
        RECT 84.240 142.220 84.560 142.280 ;
        RECT 83.335 142.080 84.560 142.220 ;
        RECT 83.335 142.035 83.625 142.080 ;
        RECT 84.240 142.020 84.560 142.080 ;
        RECT 94.790 142.220 95.080 142.265 ;
        RECT 97.120 142.220 97.440 142.280 ;
        RECT 94.790 142.080 97.440 142.220 ;
        RECT 94.790 142.035 95.080 142.080 ;
        RECT 97.120 142.020 97.440 142.080 ;
        RECT 47.900 141.880 48.220 141.940 ;
        RECT 50.200 141.880 50.520 141.940 ;
        RECT 52.975 141.880 53.265 141.925 ;
        RECT 54.340 141.880 54.660 141.940 ;
        RECT 43.850 141.740 54.660 141.880 ;
        RECT 19.315 141.695 19.605 141.740 ;
        RECT 24.440 141.680 24.760 141.740 ;
        RECT 47.900 141.680 48.220 141.740 ;
        RECT 50.200 141.680 50.520 141.740 ;
        RECT 52.975 141.695 53.265 141.740 ;
        RECT 54.340 141.680 54.660 141.740 ;
        RECT 68.140 141.680 68.460 141.940 ;
        RECT 83.795 141.880 84.085 141.925 ;
        RECT 86.095 141.880 86.385 141.925 ;
        RECT 83.795 141.740 86.385 141.880 ;
        RECT 83.795 141.695 84.085 141.740 ;
        RECT 86.095 141.695 86.385 141.740 ;
        RECT 104.020 141.680 104.340 141.940 ;
        RECT 111.010 141.880 111.150 142.375 ;
        RECT 115.520 142.360 115.840 142.420 ;
        RECT 124.720 142.360 125.040 142.420 ;
        RECT 125.655 142.375 125.945 142.420 ;
        RECT 126.575 142.375 126.865 142.605 ;
        RECT 127.035 142.375 127.325 142.605 ;
        RECT 113.680 142.265 114.000 142.280 ;
        RECT 113.650 142.035 114.000 142.265 ;
        RECT 113.680 142.020 114.000 142.035 ;
        RECT 116.900 142.220 117.220 142.280 ;
        RECT 119.675 142.220 119.965 142.265 ;
        RECT 116.900 142.080 119.965 142.220 ;
        RECT 116.900 142.020 117.220 142.080 ;
        RECT 119.675 142.035 119.965 142.080 ;
        RECT 120.595 142.220 120.885 142.265 ;
        RECT 122.420 142.220 122.740 142.280 ;
        RECT 120.595 142.080 122.740 142.220 ;
        RECT 120.595 142.035 120.885 142.080 ;
        RECT 114.140 141.880 114.460 141.940 ;
        RECT 111.010 141.740 114.460 141.880 ;
        RECT 114.140 141.680 114.460 141.740 ;
        RECT 118.280 141.880 118.600 141.940 ;
        RECT 119.215 141.880 119.505 141.925 ;
        RECT 120.670 141.880 120.810 142.035 ;
        RECT 122.420 142.020 122.740 142.080 ;
        RECT 123.355 142.220 123.645 142.265 ;
        RECT 123.800 142.220 124.120 142.280 ;
        RECT 123.355 142.080 124.120 142.220 ;
        RECT 123.355 142.035 123.645 142.080 ;
        RECT 123.800 142.020 124.120 142.080 ;
        RECT 124.275 142.035 124.565 142.265 ;
        RECT 126.100 142.220 126.420 142.280 ;
        RECT 127.110 142.220 127.250 142.375 ;
        RECT 127.480 142.360 127.800 142.620 ;
        RECT 127.940 142.560 128.260 142.620 ;
        RECT 129.780 142.560 130.100 142.620 ;
        RECT 127.940 142.420 130.100 142.560 ;
        RECT 127.940 142.360 128.260 142.420 ;
        RECT 129.780 142.360 130.100 142.420 ;
        RECT 126.100 142.080 127.250 142.220 ;
        RECT 127.570 142.220 127.710 142.360 ;
        RECT 128.400 142.220 128.720 142.280 ;
        RECT 127.570 142.080 128.720 142.220 ;
        RECT 118.280 141.740 120.810 141.880 ;
        RECT 118.280 141.680 118.600 141.740 ;
        RECT 119.215 141.695 119.505 141.740 ;
        RECT 121.500 141.680 121.820 141.940 ;
        RECT 124.350 141.880 124.490 142.035 ;
        RECT 126.100 142.020 126.420 142.080 ;
        RECT 128.400 142.020 128.720 142.080 ;
        RECT 128.875 142.220 129.165 142.265 ;
        RECT 131.020 142.220 131.310 142.265 ;
        RECT 128.875 142.080 131.310 142.220 ;
        RECT 128.875 142.035 129.165 142.080 ;
        RECT 131.020 142.035 131.310 142.080 ;
        RECT 127.480 141.880 127.800 141.940 ;
        RECT 135.760 141.880 136.080 141.940 ;
        RECT 136.695 141.880 136.985 141.925 ;
        RECT 124.350 141.740 136.985 141.880 ;
        RECT 127.480 141.680 127.800 141.740 ;
        RECT 135.760 141.680 136.080 141.740 ;
        RECT 136.695 141.695 136.985 141.740 ;
        RECT 13.330 141.060 138.910 141.540 ;
        RECT 33.195 140.860 33.485 140.905 ;
        RECT 38.700 140.860 39.020 140.920 ;
        RECT 33.195 140.720 39.020 140.860 ;
        RECT 33.195 140.675 33.485 140.720 ;
        RECT 38.700 140.660 39.020 140.720 ;
        RECT 46.980 140.860 47.300 140.920 ;
        RECT 47.915 140.860 48.205 140.905 ;
        RECT 46.980 140.720 48.205 140.860 ;
        RECT 46.980 140.660 47.300 140.720 ;
        RECT 47.915 140.675 48.205 140.720 ;
        RECT 48.360 140.660 48.680 140.920 ;
        RECT 49.740 140.860 50.060 140.920 ;
        RECT 51.120 140.860 51.440 140.920 ;
        RECT 49.370 140.720 51.440 140.860 ;
        RECT 35.495 140.520 35.785 140.565 ;
        RECT 36.860 140.520 37.180 140.580 ;
        RECT 35.495 140.380 37.180 140.520 ;
        RECT 35.495 140.335 35.785 140.380 ;
        RECT 36.860 140.320 37.180 140.380 ;
        RECT 46.075 140.520 46.365 140.565 ;
        RECT 46.520 140.520 46.840 140.580 ;
        RECT 49.370 140.565 49.510 140.720 ;
        RECT 49.740 140.660 50.060 140.720 ;
        RECT 51.120 140.660 51.440 140.720 ;
        RECT 53.435 140.675 53.725 140.905 ;
        RECT 46.075 140.380 46.840 140.520 ;
        RECT 46.075 140.335 46.365 140.380 ;
        RECT 46.520 140.320 46.840 140.380 ;
        RECT 49.295 140.335 49.585 140.565 ;
        RECT 50.660 140.520 50.980 140.580 ;
        RECT 52.500 140.565 52.820 140.580 ;
        RECT 51.595 140.520 51.885 140.565 ;
        RECT 50.660 140.380 51.885 140.520 ;
        RECT 50.660 140.320 50.980 140.380 ;
        RECT 51.595 140.335 51.885 140.380 ;
        RECT 52.500 140.335 52.885 140.565 ;
        RECT 53.510 140.520 53.650 140.675 ;
        RECT 97.120 140.660 97.440 140.920 ;
        RECT 98.975 140.860 99.265 140.905 ;
        RECT 104.020 140.860 104.340 140.920 ;
        RECT 98.975 140.720 104.340 140.860 ;
        RECT 98.975 140.675 99.265 140.720 ;
        RECT 104.020 140.660 104.340 140.720 ;
        RECT 105.400 140.660 105.720 140.920 ;
        RECT 113.680 140.660 114.000 140.920 ;
        RECT 114.140 140.660 114.460 140.920 ;
        RECT 128.400 140.860 128.720 140.920 ;
        RECT 124.810 140.720 128.720 140.860 ;
        RECT 59.460 140.520 59.750 140.565 ;
        RECT 121.500 140.520 121.820 140.580 ;
        RECT 53.510 140.380 59.750 140.520 ;
        RECT 59.460 140.335 59.750 140.380 ;
        RECT 107.790 140.380 111.150 140.520 ;
        RECT 52.500 140.320 52.820 140.335 ;
        RECT 22.140 139.980 22.460 140.240 ;
        RECT 23.075 140.180 23.365 140.225 ;
        RECT 30.880 140.180 31.200 140.240 ;
        RECT 23.075 140.040 31.200 140.180 ;
        RECT 23.075 139.995 23.365 140.040 ;
        RECT 30.880 139.980 31.200 140.040 ;
        RECT 34.575 139.995 34.865 140.225 ;
        RECT 31.800 139.840 32.120 139.900 ;
        RECT 33.195 139.840 33.485 139.885 ;
        RECT 31.800 139.700 33.485 139.840 ;
        RECT 34.650 139.840 34.790 139.995 ;
        RECT 35.020 139.980 35.340 140.240 ;
        RECT 36.400 139.980 36.720 140.240 ;
        RECT 46.995 140.180 47.285 140.225 ;
        RECT 47.900 140.180 48.220 140.240 ;
        RECT 46.995 140.040 48.220 140.180 ;
        RECT 46.995 139.995 47.285 140.040 ;
        RECT 47.900 139.980 48.220 140.040 ;
        RECT 50.200 139.980 50.520 140.240 ;
        RECT 67.650 140.180 67.940 140.225 ;
        RECT 72.280 140.180 72.600 140.240 ;
        RECT 67.650 140.040 72.600 140.180 ;
        RECT 67.650 139.995 67.940 140.040 ;
        RECT 72.280 139.980 72.600 140.040 ;
        RECT 99.435 140.180 99.725 140.225 ;
        RECT 105.860 140.180 106.180 140.240 ;
        RECT 99.435 140.040 106.180 140.180 ;
        RECT 99.435 139.995 99.725 140.040 ;
        RECT 105.860 139.980 106.180 140.040 ;
        RECT 106.320 139.980 106.640 140.240 ;
        RECT 106.795 140.180 107.085 140.225 ;
        RECT 107.240 140.180 107.560 140.240 ;
        RECT 107.790 140.225 107.930 140.380 ;
        RECT 106.795 140.040 107.560 140.180 ;
        RECT 106.795 139.995 107.085 140.040 ;
        RECT 107.240 139.980 107.560 140.040 ;
        RECT 107.715 139.995 108.005 140.225 ;
        RECT 108.175 139.995 108.465 140.225 ;
        RECT 110.000 140.180 110.320 140.240 ;
        RECT 110.475 140.180 110.765 140.225 ;
        RECT 110.000 140.040 110.765 140.180 ;
        RECT 41.920 139.840 42.240 139.900 ;
        RECT 34.650 139.700 42.240 139.840 ;
        RECT 31.800 139.640 32.120 139.700 ;
        RECT 33.195 139.655 33.485 139.700 ;
        RECT 41.920 139.640 42.240 139.700 ;
        RECT 56.205 139.840 56.495 139.885 ;
        RECT 58.725 139.840 59.015 139.885 ;
        RECT 59.915 139.840 60.205 139.885 ;
        RECT 56.205 139.700 60.205 139.840 ;
        RECT 56.205 139.655 56.495 139.700 ;
        RECT 58.725 139.655 59.015 139.700 ;
        RECT 59.915 139.655 60.205 139.700 ;
        RECT 60.795 139.840 61.085 139.885 ;
        RECT 62.620 139.840 62.940 139.900 ;
        RECT 66.315 139.840 66.605 139.885 ;
        RECT 60.795 139.700 66.605 139.840 ;
        RECT 60.795 139.655 61.085 139.700 ;
        RECT 62.620 139.640 62.940 139.700 ;
        RECT 66.315 139.655 66.605 139.700 ;
        RECT 67.195 139.840 67.485 139.885 ;
        RECT 68.385 139.840 68.675 139.885 ;
        RECT 70.905 139.840 71.195 139.885 ;
        RECT 67.195 139.700 71.195 139.840 ;
        RECT 67.195 139.655 67.485 139.700 ;
        RECT 68.385 139.655 68.675 139.700 ;
        RECT 70.905 139.655 71.195 139.700 ;
        RECT 98.960 139.840 99.280 139.900 ;
        RECT 99.895 139.840 100.185 139.885 ;
        RECT 103.100 139.840 103.420 139.900 ;
        RECT 98.960 139.700 103.420 139.840 ;
        RECT 98.960 139.640 99.280 139.700 ;
        RECT 99.895 139.655 100.185 139.700 ;
        RECT 103.100 139.640 103.420 139.700 ;
        RECT 105.400 139.840 105.720 139.900 ;
        RECT 108.250 139.840 108.390 139.995 ;
        RECT 110.000 139.980 110.320 140.040 ;
        RECT 110.475 139.995 110.765 140.040 ;
        RECT 105.400 139.700 108.390 139.840 ;
        RECT 105.400 139.640 105.720 139.700 ;
        RECT 35.480 139.500 35.800 139.560 ;
        RECT 36.415 139.500 36.705 139.545 ;
        RECT 35.480 139.360 36.705 139.500 ;
        RECT 35.480 139.300 35.800 139.360 ;
        RECT 36.415 139.315 36.705 139.360 ;
        RECT 56.640 139.500 56.930 139.545 ;
        RECT 58.210 139.500 58.500 139.545 ;
        RECT 60.310 139.500 60.600 139.545 ;
        RECT 56.640 139.360 60.600 139.500 ;
        RECT 56.640 139.315 56.930 139.360 ;
        RECT 58.210 139.315 58.500 139.360 ;
        RECT 60.310 139.315 60.600 139.360 ;
        RECT 66.800 139.500 67.090 139.545 ;
        RECT 68.900 139.500 69.190 139.545 ;
        RECT 70.470 139.500 70.760 139.545 ;
        RECT 66.800 139.360 70.760 139.500 ;
        RECT 111.010 139.500 111.150 140.380 ;
        RECT 111.470 140.380 121.820 140.520 ;
        RECT 111.470 140.225 111.610 140.380 ;
        RECT 121.500 140.320 121.820 140.380 ;
        RECT 111.395 139.995 111.685 140.225 ;
        RECT 111.840 139.980 112.160 140.240 ;
        RECT 112.315 140.180 112.605 140.225 ;
        RECT 113.680 140.180 114.000 140.240 ;
        RECT 112.315 140.040 114.000 140.180 ;
        RECT 112.315 139.995 112.605 140.040 ;
        RECT 113.680 139.980 114.000 140.040 ;
        RECT 115.060 139.980 115.380 140.240 ;
        RECT 115.980 139.980 116.300 140.240 ;
        RECT 124.810 140.180 124.950 140.720 ;
        RECT 128.400 140.660 128.720 140.720 ;
        RECT 136.680 140.660 137.000 140.920 ;
        RECT 125.180 140.520 125.500 140.580 ;
        RECT 126.575 140.520 126.865 140.565 ;
        RECT 125.180 140.380 126.865 140.520 ;
        RECT 125.180 140.320 125.500 140.380 ;
        RECT 126.575 140.335 126.865 140.380 ;
        RECT 116.530 140.040 124.950 140.180 ;
        RECT 113.770 139.840 113.910 139.980 ;
        RECT 116.530 139.840 116.670 140.040 ;
        RECT 125.640 139.980 125.960 140.240 ;
        RECT 126.100 139.980 126.420 140.240 ;
        RECT 127.480 139.980 127.800 140.240 ;
        RECT 127.940 139.980 128.260 140.240 ;
        RECT 129.290 140.180 129.580 140.225 ;
        RECT 133.000 140.180 133.320 140.240 ;
        RECT 129.290 140.040 133.320 140.180 ;
        RECT 129.290 139.995 129.580 140.040 ;
        RECT 133.000 139.980 133.320 140.040 ;
        RECT 135.760 140.225 136.080 140.240 ;
        RECT 135.760 140.180 136.095 140.225 ;
        RECT 135.760 140.040 136.275 140.180 ;
        RECT 135.760 139.995 136.095 140.040 ;
        RECT 135.760 139.980 136.080 139.995 ;
        RECT 113.770 139.700 116.670 139.840 ;
        RECT 117.820 139.840 118.140 139.900 ;
        RECT 126.560 139.840 126.880 139.900 ;
        RECT 117.820 139.700 126.880 139.840 ;
        RECT 117.820 139.640 118.140 139.700 ;
        RECT 126.560 139.640 126.880 139.700 ;
        RECT 128.835 139.840 129.125 139.885 ;
        RECT 130.025 139.840 130.315 139.885 ;
        RECT 132.545 139.840 132.835 139.885 ;
        RECT 128.835 139.700 132.835 139.840 ;
        RECT 128.835 139.655 129.125 139.700 ;
        RECT 130.025 139.655 130.315 139.700 ;
        RECT 132.545 139.655 132.835 139.700 ;
        RECT 128.440 139.500 128.730 139.545 ;
        RECT 130.540 139.500 130.830 139.545 ;
        RECT 132.110 139.500 132.400 139.545 ;
        RECT 111.010 139.360 125.870 139.500 ;
        RECT 66.800 139.315 67.090 139.360 ;
        RECT 68.900 139.315 69.190 139.360 ;
        RECT 70.470 139.315 70.760 139.360 ;
        RECT 23.075 139.160 23.365 139.205 ;
        RECT 24.900 139.160 25.220 139.220 ;
        RECT 23.075 139.020 25.220 139.160 ;
        RECT 23.075 138.975 23.365 139.020 ;
        RECT 24.900 138.960 25.220 139.020 ;
        RECT 31.340 139.160 31.660 139.220 ;
        RECT 34.115 139.160 34.405 139.205 ;
        RECT 31.340 139.020 34.405 139.160 ;
        RECT 31.340 138.960 31.660 139.020 ;
        RECT 34.115 138.975 34.405 139.020 ;
        RECT 44.220 139.160 44.540 139.220 ;
        RECT 52.515 139.160 52.805 139.205 ;
        RECT 44.220 139.020 52.805 139.160 ;
        RECT 44.220 138.960 44.540 139.020 ;
        RECT 52.515 138.975 52.805 139.020 ;
        RECT 53.895 139.160 54.185 139.205 ;
        RECT 54.340 139.160 54.660 139.220 ;
        RECT 53.895 139.020 54.660 139.160 ;
        RECT 53.895 138.975 54.185 139.020 ;
        RECT 54.340 138.960 54.660 139.020 ;
        RECT 73.215 139.160 73.505 139.205 ;
        RECT 74.120 139.160 74.440 139.220 ;
        RECT 73.215 139.020 74.440 139.160 ;
        RECT 73.215 138.975 73.505 139.020 ;
        RECT 74.120 138.960 74.440 139.020 ;
        RECT 111.380 139.160 111.700 139.220 ;
        RECT 124.735 139.160 125.025 139.205 ;
        RECT 111.380 139.020 125.025 139.160 ;
        RECT 125.730 139.160 125.870 139.360 ;
        RECT 128.440 139.360 132.400 139.500 ;
        RECT 128.440 139.315 128.730 139.360 ;
        RECT 130.540 139.315 130.830 139.360 ;
        RECT 132.110 139.315 132.400 139.360 ;
        RECT 133.460 139.160 133.780 139.220 ;
        RECT 125.730 139.020 133.780 139.160 ;
        RECT 111.380 138.960 111.700 139.020 ;
        RECT 124.735 138.975 125.025 139.020 ;
        RECT 133.460 138.960 133.780 139.020 ;
        RECT 134.840 138.960 135.160 139.220 ;
        RECT 13.330 138.340 138.910 138.820 ;
        RECT 20.760 138.140 21.080 138.200 ;
        RECT 24.915 138.140 25.205 138.185 ;
        RECT 33.655 138.140 33.945 138.185 ;
        RECT 35.940 138.140 36.260 138.200 ;
        RECT 20.760 138.000 33.410 138.140 ;
        RECT 20.760 137.940 21.080 138.000 ;
        RECT 24.915 137.955 25.205 138.000 ;
        RECT 25.820 137.800 26.140 137.860 ;
        RECT 33.270 137.800 33.410 138.000 ;
        RECT 33.655 138.000 36.260 138.140 ;
        RECT 33.655 137.955 33.945 138.000 ;
        RECT 35.940 137.940 36.260 138.000 ;
        RECT 52.500 137.940 52.820 138.200 ;
        RECT 105.860 138.140 106.180 138.200 ;
        RECT 107.255 138.140 107.545 138.185 ;
        RECT 105.860 138.000 107.545 138.140 ;
        RECT 105.860 137.940 106.180 138.000 ;
        RECT 107.255 137.955 107.545 138.000 ;
        RECT 108.620 138.140 108.940 138.200 ;
        RECT 110.475 138.140 110.765 138.185 ;
        RECT 125.640 138.140 125.960 138.200 ;
        RECT 131.620 138.140 131.940 138.200 ;
        RECT 108.620 138.000 110.765 138.140 ;
        RECT 108.620 137.940 108.940 138.000 ;
        RECT 110.475 137.955 110.765 138.000 ;
        RECT 118.830 138.000 131.940 138.140 ;
        RECT 64.960 137.800 65.250 137.845 ;
        RECT 67.060 137.800 67.350 137.845 ;
        RECT 68.630 137.800 68.920 137.845 ;
        RECT 72.295 137.800 72.585 137.845 ;
        RECT 25.820 137.660 27.890 137.800 ;
        RECT 33.270 137.660 36.170 137.800 ;
        RECT 25.820 137.600 26.140 137.660 ;
        RECT 22.140 137.460 22.460 137.520 ;
        RECT 22.140 137.320 26.970 137.460 ;
        RECT 22.140 137.260 22.460 137.320 ;
        RECT 26.830 137.165 26.970 137.320 ;
        RECT 27.750 137.165 27.890 137.660 ;
        RECT 36.030 137.520 36.170 137.660 ;
        RECT 64.960 137.660 68.920 137.800 ;
        RECT 64.960 137.615 65.250 137.660 ;
        RECT 67.060 137.615 67.350 137.660 ;
        RECT 68.630 137.615 68.920 137.660 ;
        RECT 69.840 137.660 72.585 137.800 ;
        RECT 35.940 137.260 36.260 137.520 ;
        RECT 43.760 137.460 44.080 137.520 ;
        RECT 52.960 137.460 53.280 137.520 ;
        RECT 43.760 137.320 53.280 137.460 ;
        RECT 43.760 137.260 44.080 137.320 ;
        RECT 52.960 137.260 53.280 137.320 ;
        RECT 53.895 137.460 54.185 137.505 ;
        RECT 55.260 137.460 55.580 137.520 ;
        RECT 53.895 137.320 55.580 137.460 ;
        RECT 53.895 137.275 54.185 137.320 ;
        RECT 19.395 137.120 19.685 137.165 ;
        RECT 21.695 137.120 21.985 137.165 ;
        RECT 19.395 136.980 21.985 137.120 ;
        RECT 19.395 136.935 19.685 136.980 ;
        RECT 21.695 136.935 21.985 136.980 ;
        RECT 22.230 136.980 26.050 137.120 ;
        RECT 14.780 136.780 15.100 136.840 ;
        RECT 21.220 136.780 21.540 136.840 ;
        RECT 22.230 136.780 22.370 136.980 ;
        RECT 14.780 136.640 20.990 136.780 ;
        RECT 14.780 136.580 15.100 136.640 ;
        RECT 17.540 136.440 17.860 136.500 ;
        RECT 18.475 136.440 18.765 136.485 ;
        RECT 17.540 136.300 18.765 136.440 ;
        RECT 17.540 136.240 17.860 136.300 ;
        RECT 18.475 136.255 18.765 136.300 ;
        RECT 19.840 136.240 20.160 136.500 ;
        RECT 20.300 136.240 20.620 136.500 ;
        RECT 20.850 136.440 20.990 136.640 ;
        RECT 21.220 136.640 22.370 136.780 ;
        RECT 21.220 136.580 21.540 136.640 ;
        RECT 22.600 136.580 22.920 136.840 ;
        RECT 23.520 136.780 23.840 136.840 ;
        RECT 24.900 136.825 25.220 136.840 ;
        RECT 25.910 136.825 26.050 136.980 ;
        RECT 26.755 136.935 27.045 137.165 ;
        RECT 27.675 137.120 27.965 137.165 ;
        RECT 29.960 137.120 30.280 137.180 ;
        RECT 27.675 136.980 30.280 137.120 ;
        RECT 27.675 136.935 27.965 136.980 ;
        RECT 29.960 136.920 30.280 136.980 ;
        RECT 35.020 136.920 35.340 137.180 ;
        RECT 49.280 136.920 49.600 137.180 ;
        RECT 50.200 136.920 50.520 137.180 ;
        RECT 50.675 136.935 50.965 137.165 ;
        RECT 51.580 137.120 51.900 137.180 ;
        RECT 53.970 137.120 54.110 137.275 ;
        RECT 55.260 137.260 55.580 137.320 ;
        RECT 62.620 137.460 62.940 137.520 ;
        RECT 64.475 137.460 64.765 137.505 ;
        RECT 62.620 137.320 64.765 137.460 ;
        RECT 62.620 137.260 62.940 137.320 ;
        RECT 64.475 137.275 64.765 137.320 ;
        RECT 65.355 137.460 65.645 137.505 ;
        RECT 66.545 137.460 66.835 137.505 ;
        RECT 69.065 137.460 69.355 137.505 ;
        RECT 65.355 137.320 69.355 137.460 ;
        RECT 65.355 137.275 65.645 137.320 ;
        RECT 66.545 137.275 66.835 137.320 ;
        RECT 69.065 137.275 69.355 137.320 ;
        RECT 51.580 136.980 54.110 137.120 ;
        RECT 23.520 136.640 24.670 136.780 ;
        RECT 23.520 136.580 23.840 136.640 ;
        RECT 23.610 136.440 23.750 136.580 ;
        RECT 20.850 136.300 23.750 136.440 ;
        RECT 23.980 136.240 24.300 136.500 ;
        RECT 24.530 136.440 24.670 136.640 ;
        RECT 24.810 136.595 25.220 136.825 ;
        RECT 25.835 136.780 26.125 136.825 ;
        RECT 33.655 136.780 33.945 136.825 ;
        RECT 34.100 136.780 34.420 136.840 ;
        RECT 25.835 136.640 26.970 136.780 ;
        RECT 25.835 136.595 26.125 136.640 ;
        RECT 24.900 136.580 25.220 136.595 ;
        RECT 26.830 136.500 26.970 136.640 ;
        RECT 33.655 136.640 34.420 136.780 ;
        RECT 33.655 136.595 33.945 136.640 ;
        RECT 34.100 136.580 34.420 136.640 ;
        RECT 49.755 136.780 50.045 136.825 ;
        RECT 50.750 136.780 50.890 136.935 ;
        RECT 51.580 136.920 51.900 136.980 ;
        RECT 54.340 136.920 54.660 137.180 ;
        RECT 65.810 137.120 66.100 137.165 ;
        RECT 69.840 137.120 69.980 137.660 ;
        RECT 72.295 137.615 72.585 137.660 ;
        RECT 78.760 137.800 79.050 137.845 ;
        RECT 80.860 137.800 81.150 137.845 ;
        RECT 82.430 137.800 82.720 137.845 ;
        RECT 111.380 137.800 111.700 137.860 ;
        RECT 115.060 137.800 115.380 137.860 ;
        RECT 78.760 137.660 82.720 137.800 ;
        RECT 78.760 137.615 79.050 137.660 ;
        RECT 80.860 137.615 81.150 137.660 ;
        RECT 82.430 137.615 82.720 137.660 ;
        RECT 110.090 137.660 111.700 137.800 ;
        RECT 73.200 137.460 73.520 137.520 ;
        RECT 75.055 137.460 75.345 137.505 ;
        RECT 73.200 137.320 75.345 137.460 ;
        RECT 73.200 137.260 73.520 137.320 ;
        RECT 75.055 137.275 75.345 137.320 ;
        RECT 79.155 137.460 79.445 137.505 ;
        RECT 80.345 137.460 80.635 137.505 ;
        RECT 82.865 137.460 83.155 137.505 ;
        RECT 79.155 137.320 83.155 137.460 ;
        RECT 79.155 137.275 79.445 137.320 ;
        RECT 80.345 137.275 80.635 137.320 ;
        RECT 82.865 137.275 83.155 137.320 ;
        RECT 88.855 137.275 89.145 137.505 ;
        RECT 92.060 137.460 92.380 137.520 ;
        RECT 97.135 137.460 97.425 137.505 ;
        RECT 106.780 137.460 107.100 137.520 ;
        RECT 109.080 137.460 109.400 137.520 ;
        RECT 92.060 137.320 107.100 137.460 ;
        RECT 65.810 136.980 69.980 137.120 ;
        RECT 74.135 137.120 74.425 137.165 ;
        RECT 74.580 137.120 74.900 137.180 ;
        RECT 74.135 136.980 74.900 137.120 ;
        RECT 65.810 136.935 66.100 136.980 ;
        RECT 74.135 136.935 74.425 136.980 ;
        RECT 49.755 136.640 50.890 136.780 ;
        RECT 49.755 136.595 50.045 136.640 ;
        RECT 26.280 136.440 26.600 136.500 ;
        RECT 24.530 136.300 26.600 136.440 ;
        RECT 26.280 136.240 26.600 136.300 ;
        RECT 26.740 136.240 27.060 136.500 ;
        RECT 27.215 136.440 27.505 136.485 ;
        RECT 28.120 136.440 28.440 136.500 ;
        RECT 27.215 136.300 28.440 136.440 ;
        RECT 27.215 136.255 27.505 136.300 ;
        RECT 28.120 136.240 28.440 136.300 ;
        RECT 34.560 136.440 34.880 136.500 ;
        RECT 36.860 136.440 37.180 136.500 ;
        RECT 41.460 136.440 41.780 136.500 ;
        RECT 34.560 136.300 41.780 136.440 ;
        RECT 34.560 136.240 34.880 136.300 ;
        RECT 36.860 136.240 37.180 136.300 ;
        RECT 41.460 136.240 41.780 136.300 ;
        RECT 51.120 136.240 51.440 136.500 ;
        RECT 71.375 136.440 71.665 136.485 ;
        RECT 74.210 136.440 74.350 136.935 ;
        RECT 74.580 136.920 74.900 136.980 ;
        RECT 78.275 137.120 78.565 137.165 ;
        RECT 81.480 137.120 81.800 137.180 ;
        RECT 78.275 136.980 81.800 137.120 ;
        RECT 78.275 136.935 78.565 136.980 ;
        RECT 81.480 136.920 81.800 136.980 ;
        RECT 81.940 137.120 82.260 137.180 ;
        RECT 88.930 137.120 89.070 137.275 ;
        RECT 92.060 137.260 92.380 137.320 ;
        RECT 97.135 137.275 97.425 137.320 ;
        RECT 106.780 137.260 107.100 137.320 ;
        RECT 108.250 137.320 109.400 137.460 ;
        RECT 81.940 136.980 89.070 137.120 ;
        RECT 81.940 136.920 82.260 136.980 ;
        RECT 101.735 136.935 102.025 137.165 ;
        RECT 106.320 137.120 106.640 137.180 ;
        RECT 108.250 137.165 108.390 137.320 ;
        RECT 109.080 137.260 109.400 137.320 ;
        RECT 108.175 137.120 108.465 137.165 ;
        RECT 106.320 136.980 108.465 137.120 ;
        RECT 79.610 136.780 79.900 136.825 ;
        RECT 80.560 136.780 80.880 136.840 ;
        RECT 79.610 136.640 80.880 136.780 ;
        RECT 79.610 136.595 79.900 136.640 ;
        RECT 80.560 136.580 80.880 136.640 ;
        RECT 96.215 136.780 96.505 136.825 ;
        RECT 98.515 136.780 98.805 136.825 ;
        RECT 96.215 136.640 98.805 136.780 ;
        RECT 96.215 136.595 96.505 136.640 ;
        RECT 98.515 136.595 98.805 136.640 ;
        RECT 71.375 136.300 74.350 136.440 ;
        RECT 74.595 136.440 74.885 136.485 ;
        RECT 78.720 136.440 79.040 136.500 ;
        RECT 74.595 136.300 79.040 136.440 ;
        RECT 71.375 136.255 71.665 136.300 ;
        RECT 74.595 136.255 74.885 136.300 ;
        RECT 78.720 136.240 79.040 136.300 ;
        RECT 80.100 136.440 80.420 136.500 ;
        RECT 85.175 136.440 85.465 136.485 ;
        RECT 80.100 136.300 85.465 136.440 ;
        RECT 80.100 136.240 80.420 136.300 ;
        RECT 85.175 136.255 85.465 136.300 ;
        RECT 85.620 136.440 85.940 136.500 ;
        RECT 86.095 136.440 86.385 136.485 ;
        RECT 85.620 136.300 86.385 136.440 ;
        RECT 85.620 136.240 85.940 136.300 ;
        RECT 86.095 136.255 86.385 136.300 ;
        RECT 87.920 136.240 88.240 136.500 ;
        RECT 88.395 136.440 88.685 136.485 ;
        RECT 90.680 136.440 91.000 136.500 ;
        RECT 88.395 136.300 91.000 136.440 ;
        RECT 88.395 136.255 88.685 136.300 ;
        RECT 90.680 136.240 91.000 136.300 ;
        RECT 94.360 136.240 94.680 136.500 ;
        RECT 96.660 136.240 96.980 136.500 ;
        RECT 101.810 136.440 101.950 136.935 ;
        RECT 106.320 136.920 106.640 136.980 ;
        RECT 108.175 136.935 108.465 136.980 ;
        RECT 108.635 136.935 108.925 137.165 ;
        RECT 108.710 136.780 108.850 136.935 ;
        RECT 109.540 136.920 109.860 137.180 ;
        RECT 110.090 137.165 110.230 137.660 ;
        RECT 111.380 137.600 111.700 137.660 ;
        RECT 111.930 137.660 115.380 137.800 ;
        RECT 110.015 136.935 110.305 137.165 ;
        RECT 110.460 137.120 110.780 137.180 ;
        RECT 111.930 137.165 112.070 137.660 ;
        RECT 115.060 137.600 115.380 137.660 ;
        RECT 117.835 137.615 118.125 137.845 ;
        RECT 117.910 137.460 118.050 137.615 ;
        RECT 112.850 137.320 118.050 137.460 ;
        RECT 112.850 137.165 112.990 137.320 ;
        RECT 111.395 137.120 111.685 137.165 ;
        RECT 110.460 136.980 111.685 137.120 ;
        RECT 110.460 136.920 110.780 136.980 ;
        RECT 111.395 136.935 111.685 136.980 ;
        RECT 111.855 136.935 112.145 137.165 ;
        RECT 112.775 136.935 113.065 137.165 ;
        RECT 113.220 136.920 113.540 137.180 ;
        RECT 114.600 136.920 114.920 137.180 ;
        RECT 115.535 137.120 115.825 137.165 ;
        RECT 116.900 137.120 117.220 137.180 ;
        RECT 118.830 137.165 118.970 138.000 ;
        RECT 125.640 137.940 125.960 138.000 ;
        RECT 131.620 137.940 131.940 138.000 ;
        RECT 133.000 137.940 133.320 138.200 ;
        RECT 133.460 137.940 133.780 138.200 ;
        RECT 125.180 137.800 125.500 137.860 ;
        RECT 129.780 137.800 130.100 137.860 ;
        RECT 125.180 137.660 135.530 137.800 ;
        RECT 125.180 137.600 125.500 137.660 ;
        RECT 129.780 137.600 130.100 137.660 ;
        RECT 125.270 137.460 125.410 137.600 ;
        RECT 119.750 137.320 125.410 137.460 ;
        RECT 127.020 137.460 127.340 137.520 ;
        RECT 129.320 137.460 129.640 137.520 ;
        RECT 127.020 137.320 129.640 137.460 ;
        RECT 119.750 137.165 119.890 137.320 ;
        RECT 127.020 137.260 127.340 137.320 ;
        RECT 129.320 137.260 129.640 137.320 ;
        RECT 130.240 137.460 130.560 137.520 ;
        RECT 130.240 137.320 131.850 137.460 ;
        RECT 130.240 137.260 130.560 137.320 ;
        RECT 115.535 136.980 117.220 137.120 ;
        RECT 115.535 136.935 115.825 136.980 ;
        RECT 116.900 136.920 117.220 136.980 ;
        RECT 118.755 136.935 119.045 137.165 ;
        RECT 119.675 136.935 119.965 137.165 ;
        RECT 120.595 137.120 120.885 137.165 ;
        RECT 121.040 137.120 121.360 137.180 ;
        RECT 120.595 136.980 121.360 137.120 ;
        RECT 120.595 136.935 120.885 136.980 ;
        RECT 121.040 136.920 121.360 136.980 ;
        RECT 124.720 137.120 125.040 137.180 ;
        RECT 129.795 137.120 130.085 137.165 ;
        RECT 124.720 136.980 130.085 137.120 ;
        RECT 124.720 136.920 125.040 136.980 ;
        RECT 129.795 136.935 130.085 136.980 ;
        RECT 130.715 136.935 131.005 137.165 ;
        RECT 108.710 136.640 114.370 136.780 ;
        RECT 104.480 136.440 104.800 136.500 ;
        RECT 108.620 136.440 108.940 136.500 ;
        RECT 101.810 136.300 108.940 136.440 ;
        RECT 104.480 136.240 104.800 136.300 ;
        RECT 108.620 136.240 108.940 136.300 ;
        RECT 110.000 136.440 110.320 136.500 ;
        RECT 113.695 136.440 113.985 136.485 ;
        RECT 110.000 136.300 113.985 136.440 ;
        RECT 114.230 136.440 114.370 136.640 ;
        RECT 119.215 136.595 119.505 136.825 ;
        RECT 122.420 136.780 122.740 136.840 ;
        RECT 127.035 136.780 127.325 136.825 ;
        RECT 122.420 136.640 127.325 136.780 ;
        RECT 118.280 136.440 118.600 136.500 ;
        RECT 114.230 136.300 118.600 136.440 ;
        RECT 119.290 136.440 119.430 136.595 ;
        RECT 122.420 136.580 122.740 136.640 ;
        RECT 127.035 136.595 127.325 136.640 ;
        RECT 127.955 136.595 128.245 136.825 ;
        RECT 128.875 136.780 129.165 136.825 ;
        RECT 130.790 136.780 130.930 136.935 ;
        RECT 131.160 136.920 131.480 137.180 ;
        RECT 131.710 137.165 131.850 137.320 ;
        RECT 131.635 136.935 131.925 137.165 ;
        RECT 132.080 137.120 132.400 137.180 ;
        RECT 135.390 137.165 135.530 137.660 ;
        RECT 134.395 137.120 134.685 137.165 ;
        RECT 132.080 136.980 134.685 137.120 ;
        RECT 132.080 136.920 132.400 136.980 ;
        RECT 134.395 136.935 134.685 136.980 ;
        RECT 135.315 136.935 135.605 137.165 ;
        RECT 136.220 136.920 136.540 137.180 ;
        RECT 128.875 136.640 130.930 136.780 ;
        RECT 128.875 136.595 129.165 136.640 ;
        RECT 123.800 136.440 124.120 136.500 ;
        RECT 119.290 136.300 124.120 136.440 ;
        RECT 128.030 136.440 128.170 136.595 ;
        RECT 134.840 136.580 135.160 136.840 ;
        RECT 134.930 136.440 135.070 136.580 ;
        RECT 135.760 136.440 136.080 136.500 ;
        RECT 128.030 136.300 136.080 136.440 ;
        RECT 110.000 136.240 110.320 136.300 ;
        RECT 113.695 136.255 113.985 136.300 ;
        RECT 118.280 136.240 118.600 136.300 ;
        RECT 123.800 136.240 124.120 136.300 ;
        RECT 135.760 136.240 136.080 136.300 ;
        RECT 13.330 135.620 138.910 136.100 ;
        RECT 15.715 135.420 16.005 135.465 ;
        RECT 19.840 135.420 20.160 135.480 ;
        RECT 15.715 135.280 20.160 135.420 ;
        RECT 15.715 135.235 16.005 135.280 ;
        RECT 19.840 135.220 20.160 135.280 ;
        RECT 22.140 135.420 22.460 135.480 ;
        RECT 23.535 135.420 23.825 135.465 ;
        RECT 22.140 135.280 23.825 135.420 ;
        RECT 22.140 135.220 22.460 135.280 ;
        RECT 23.535 135.235 23.825 135.280 ;
        RECT 24.375 135.420 24.665 135.465 ;
        RECT 26.280 135.420 26.600 135.480 ;
        RECT 27.660 135.420 27.980 135.480 ;
        RECT 24.375 135.280 27.980 135.420 ;
        RECT 24.375 135.235 24.665 135.280 ;
        RECT 26.280 135.220 26.600 135.280 ;
        RECT 27.660 135.220 27.980 135.280 ;
        RECT 29.515 135.420 29.805 135.465 ;
        RECT 31.800 135.420 32.120 135.480 ;
        RECT 29.515 135.280 32.120 135.420 ;
        RECT 29.515 135.235 29.805 135.280 ;
        RECT 23.060 135.080 23.380 135.140 ;
        RECT 16.250 134.940 23.380 135.080 ;
        RECT 14.780 134.540 15.100 134.800 ;
        RECT 16.250 134.785 16.390 134.940 ;
        RECT 23.060 134.880 23.380 134.940 ;
        RECT 24.900 135.080 25.220 135.140 ;
        RECT 25.375 135.080 25.665 135.125 ;
        RECT 27.200 135.080 27.520 135.140 ;
        RECT 29.590 135.080 29.730 135.235 ;
        RECT 31.800 135.220 32.120 135.280 ;
        RECT 33.195 135.420 33.485 135.465 ;
        RECT 34.100 135.420 34.420 135.480 ;
        RECT 33.195 135.280 34.420 135.420 ;
        RECT 33.195 135.235 33.485 135.280 ;
        RECT 34.100 135.220 34.420 135.280 ;
        RECT 36.400 135.220 36.720 135.480 ;
        RECT 46.995 135.420 47.285 135.465 ;
        RECT 49.295 135.420 49.585 135.465 ;
        RECT 50.200 135.420 50.520 135.480 ;
        RECT 46.995 135.280 50.520 135.420 ;
        RECT 46.995 135.235 47.285 135.280 ;
        RECT 49.295 135.235 49.585 135.280 ;
        RECT 50.200 135.220 50.520 135.280 ;
        RECT 69.980 135.420 70.300 135.480 ;
        RECT 72.295 135.420 72.585 135.465 ;
        RECT 69.980 135.280 72.585 135.420 ;
        RECT 69.980 135.220 70.300 135.280 ;
        RECT 72.295 135.235 72.585 135.280 ;
        RECT 24.900 134.940 26.970 135.080 ;
        RECT 24.900 134.880 25.220 134.940 ;
        RECT 25.375 134.895 25.665 134.940 ;
        RECT 17.540 134.785 17.860 134.800 ;
        RECT 26.830 134.785 26.970 134.940 ;
        RECT 27.200 134.940 29.730 135.080 ;
        RECT 29.960 135.080 30.280 135.140 ;
        RECT 48.835 135.080 49.125 135.125 ;
        RECT 51.580 135.080 51.900 135.140 ;
        RECT 29.960 134.940 32.490 135.080 ;
        RECT 27.200 134.880 27.520 134.940 ;
        RECT 29.960 134.880 30.280 134.940 ;
        RECT 15.715 134.555 16.005 134.785 ;
        RECT 16.175 134.555 16.465 134.785 ;
        RECT 17.510 134.740 17.860 134.785 ;
        RECT 17.345 134.600 17.860 134.740 ;
        RECT 17.510 134.555 17.860 134.600 ;
        RECT 26.755 134.555 27.045 134.785 ;
        RECT 27.660 134.740 27.980 134.800 ;
        RECT 29.055 134.740 29.345 134.785 ;
        RECT 27.660 134.600 29.345 134.740 ;
        RECT 15.790 134.400 15.930 134.555 ;
        RECT 17.540 134.540 17.860 134.555 ;
        RECT 17.055 134.400 17.345 134.445 ;
        RECT 18.245 134.400 18.535 134.445 ;
        RECT 20.765 134.400 21.055 134.445 ;
        RECT 15.790 134.260 16.390 134.400 ;
        RECT 16.250 133.720 16.390 134.260 ;
        RECT 17.055 134.260 21.055 134.400 ;
        RECT 26.830 134.400 26.970 134.555 ;
        RECT 27.660 134.540 27.980 134.600 ;
        RECT 29.055 134.555 29.345 134.600 ;
        RECT 30.435 134.740 30.725 134.785 ;
        RECT 31.340 134.740 31.660 134.800 ;
        RECT 32.350 134.785 32.490 134.940 ;
        RECT 48.835 134.940 51.900 135.080 ;
        RECT 72.370 135.080 72.510 135.235 ;
        RECT 73.200 135.220 73.520 135.480 ;
        RECT 80.560 135.420 80.880 135.480 ;
        RECT 81.035 135.420 81.325 135.465 ;
        RECT 80.560 135.280 81.325 135.420 ;
        RECT 80.560 135.220 80.880 135.280 ;
        RECT 81.035 135.235 81.325 135.280 ;
        RECT 99.895 135.420 100.185 135.465 ;
        RECT 104.480 135.420 104.800 135.480 ;
        RECT 99.895 135.280 104.800 135.420 ;
        RECT 99.895 135.235 100.185 135.280 ;
        RECT 104.480 135.220 104.800 135.280 ;
        RECT 112.775 135.420 113.065 135.465 ;
        RECT 114.600 135.420 114.920 135.480 ;
        RECT 112.775 135.280 114.920 135.420 ;
        RECT 112.775 135.235 113.065 135.280 ;
        RECT 114.600 135.220 114.920 135.280 ;
        RECT 136.680 135.220 137.000 135.480 ;
        RECT 72.370 134.940 75.730 135.080 ;
        RECT 48.835 134.895 49.125 134.940 ;
        RECT 51.580 134.880 51.900 134.940 ;
        RECT 30.435 134.600 31.660 134.740 ;
        RECT 30.435 134.555 30.725 134.600 ;
        RECT 30.510 134.400 30.650 134.555 ;
        RECT 31.340 134.540 31.660 134.600 ;
        RECT 32.275 134.555 32.565 134.785 ;
        RECT 26.830 134.260 30.650 134.400 ;
        RECT 30.895 134.400 31.185 134.445 ;
        RECT 31.800 134.400 32.120 134.460 ;
        RECT 30.895 134.260 32.120 134.400 ;
        RECT 17.055 134.215 17.345 134.260 ;
        RECT 18.245 134.215 18.535 134.260 ;
        RECT 20.765 134.215 21.055 134.260 ;
        RECT 30.895 134.215 31.185 134.260 ;
        RECT 31.800 134.200 32.120 134.260 ;
        RECT 16.660 134.060 16.950 134.105 ;
        RECT 18.760 134.060 19.050 134.105 ;
        RECT 20.330 134.060 20.620 134.105 ;
        RECT 16.660 133.920 20.620 134.060 ;
        RECT 16.660 133.875 16.950 133.920 ;
        RECT 18.760 133.875 19.050 133.920 ;
        RECT 20.330 133.875 20.620 133.920 ;
        RECT 25.820 133.860 26.140 134.120 ;
        RECT 28.595 134.060 28.885 134.105 ;
        RECT 31.340 134.060 31.660 134.120 ;
        RECT 28.595 133.920 31.660 134.060 ;
        RECT 32.350 134.060 32.490 134.555 ;
        RECT 33.640 134.540 33.960 134.800 ;
        RECT 34.100 134.740 34.420 134.800 ;
        RECT 35.035 134.740 35.325 134.785 ;
        RECT 34.100 134.600 35.325 134.740 ;
        RECT 34.100 134.540 34.420 134.600 ;
        RECT 35.035 134.555 35.325 134.600 ;
        RECT 35.495 134.555 35.785 134.785 ;
        RECT 41.460 134.740 41.780 134.800 ;
        RECT 46.980 134.740 47.300 134.800 ;
        RECT 47.455 134.740 47.745 134.785 ;
        RECT 41.460 134.600 47.745 134.740 ;
        RECT 34.560 134.400 34.880 134.460 ;
        RECT 35.570 134.400 35.710 134.555 ;
        RECT 41.460 134.540 41.780 134.600 ;
        RECT 46.980 134.540 47.300 134.600 ;
        RECT 47.455 134.555 47.745 134.600 ;
        RECT 47.900 134.540 48.220 134.800 ;
        RECT 52.040 134.740 52.360 134.800 ;
        RECT 54.860 134.740 55.150 134.785 ;
        RECT 52.040 134.600 55.150 134.740 ;
        RECT 52.040 134.540 52.360 134.600 ;
        RECT 54.860 134.555 55.150 134.600 ;
        RECT 56.195 134.740 56.485 134.785 ;
        RECT 62.620 134.740 62.940 134.800 ;
        RECT 66.760 134.785 67.080 134.800 ;
        RECT 65.395 134.740 65.685 134.785 ;
        RECT 56.195 134.600 65.685 134.740 ;
        RECT 56.195 134.555 56.485 134.600 ;
        RECT 62.620 134.540 62.940 134.600 ;
        RECT 65.395 134.555 65.685 134.600 ;
        RECT 66.730 134.555 67.080 134.785 ;
        RECT 66.760 134.540 67.080 134.555 ;
        RECT 72.740 134.540 73.060 134.800 ;
        RECT 73.750 134.785 73.890 134.940 ;
        RECT 73.675 134.555 73.965 134.785 ;
        RECT 74.120 134.540 74.440 134.800 ;
        RECT 34.560 134.260 35.710 134.400 ;
        RECT 46.060 134.400 46.380 134.460 ;
        RECT 48.820 134.400 49.140 134.460 ;
        RECT 46.060 134.260 49.140 134.400 ;
        RECT 34.560 134.200 34.880 134.260 ;
        RECT 46.060 134.200 46.380 134.260 ;
        RECT 48.820 134.200 49.140 134.260 ;
        RECT 51.605 134.400 51.895 134.445 ;
        RECT 54.125 134.400 54.415 134.445 ;
        RECT 55.315 134.400 55.605 134.445 ;
        RECT 51.605 134.260 55.605 134.400 ;
        RECT 51.605 134.215 51.895 134.260 ;
        RECT 54.125 134.215 54.415 134.260 ;
        RECT 55.315 134.215 55.605 134.260 ;
        RECT 66.275 134.400 66.565 134.445 ;
        RECT 67.465 134.400 67.755 134.445 ;
        RECT 69.985 134.400 70.275 134.445 ;
        RECT 66.275 134.260 70.275 134.400 ;
        RECT 72.830 134.400 72.970 134.540 ;
        RECT 72.830 134.260 73.890 134.400 ;
        RECT 66.275 134.215 66.565 134.260 ;
        RECT 67.465 134.215 67.755 134.260 ;
        RECT 69.985 134.215 70.275 134.260 ;
        RECT 73.750 134.120 73.890 134.260 ;
        RECT 34.115 134.060 34.405 134.105 ;
        RECT 32.350 133.920 34.405 134.060 ;
        RECT 28.595 133.875 28.885 133.920 ;
        RECT 31.340 133.860 31.660 133.920 ;
        RECT 34.115 133.875 34.405 133.920 ;
        RECT 52.040 134.060 52.330 134.105 ;
        RECT 53.610 134.060 53.900 134.105 ;
        RECT 55.710 134.060 56.000 134.105 ;
        RECT 52.040 133.920 56.000 134.060 ;
        RECT 52.040 133.875 52.330 133.920 ;
        RECT 53.610 133.875 53.900 133.920 ;
        RECT 55.710 133.875 56.000 133.920 ;
        RECT 65.880 134.060 66.170 134.105 ;
        RECT 67.980 134.060 68.270 134.105 ;
        RECT 69.550 134.060 69.840 134.105 ;
        RECT 65.880 133.920 69.840 134.060 ;
        RECT 65.880 133.875 66.170 133.920 ;
        RECT 67.980 133.875 68.270 133.920 ;
        RECT 69.550 133.875 69.840 133.920 ;
        RECT 73.660 133.860 73.980 134.120 ;
        RECT 22.600 133.720 22.920 133.780 ;
        RECT 23.075 133.720 23.365 133.765 ;
        RECT 24.455 133.720 24.745 133.765 ;
        RECT 27.200 133.720 27.520 133.780 ;
        RECT 16.250 133.580 27.520 133.720 ;
        RECT 22.600 133.520 22.920 133.580 ;
        RECT 23.075 133.535 23.365 133.580 ;
        RECT 24.455 133.535 24.745 133.580 ;
        RECT 27.200 133.520 27.520 133.580 ;
        RECT 30.435 133.720 30.725 133.765 ;
        RECT 30.880 133.720 31.200 133.780 ;
        RECT 30.435 133.580 31.200 133.720 ;
        RECT 30.435 133.535 30.725 133.580 ;
        RECT 30.880 133.520 31.200 133.580 ;
        RECT 31.800 133.720 32.120 133.780 ;
        RECT 35.940 133.720 36.260 133.780 ;
        RECT 52.500 133.720 52.820 133.780 ;
        RECT 31.800 133.580 52.820 133.720 ;
        RECT 75.590 133.720 75.730 134.940 ;
        RECT 75.960 134.880 76.280 135.140 ;
        RECT 94.360 135.125 94.680 135.140 ;
        RECT 94.330 135.080 94.680 135.125 ;
        RECT 112.300 135.080 112.620 135.140 ;
        RECT 126.100 135.080 126.420 135.140 ;
        RECT 130.700 135.080 131.020 135.140 ;
        RECT 81.570 134.940 93.210 135.080 ;
        RECT 94.165 134.940 94.680 135.080 ;
        RECT 81.570 134.800 81.710 134.940 ;
        RECT 93.070 134.800 93.210 134.940 ;
        RECT 94.330 134.895 94.680 134.940 ;
        RECT 94.360 134.880 94.680 134.895 ;
        RECT 105.950 134.940 117.130 135.080 ;
        RECT 77.340 134.740 77.660 134.800 ;
        RECT 79.195 134.740 79.485 134.785 ;
        RECT 80.100 134.740 80.420 134.800 ;
        RECT 77.340 134.600 80.420 134.740 ;
        RECT 77.340 134.540 77.660 134.600 ;
        RECT 79.195 134.555 79.485 134.600 ;
        RECT 80.100 134.540 80.420 134.600 ;
        RECT 81.480 134.540 81.800 134.800 ;
        RECT 82.830 134.740 83.120 134.785 ;
        RECT 85.620 134.740 85.940 134.800 ;
        RECT 82.830 134.600 85.940 134.740 ;
        RECT 82.830 134.555 83.120 134.600 ;
        RECT 85.620 134.540 85.940 134.600 ;
        RECT 92.980 134.540 93.300 134.800 ;
        RECT 102.195 134.740 102.485 134.785 ;
        RECT 104.020 134.740 104.340 134.800 ;
        RECT 105.950 134.785 106.090 134.940 ;
        RECT 112.300 134.880 112.620 134.940 ;
        RECT 107.240 134.785 107.560 134.800 ;
        RECT 102.195 134.600 104.340 134.740 ;
        RECT 102.195 134.555 102.485 134.600 ;
        RECT 104.020 134.540 104.340 134.600 ;
        RECT 105.875 134.555 106.165 134.785 ;
        RECT 107.210 134.555 107.560 134.785 ;
        RECT 107.240 134.540 107.560 134.555 ;
        RECT 108.620 134.740 108.940 134.800 ;
        RECT 116.990 134.785 117.130 134.940 ;
        RECT 126.100 134.940 131.850 135.080 ;
        RECT 126.100 134.880 126.420 134.940 ;
        RECT 130.700 134.880 131.020 134.940 ;
        RECT 113.695 134.740 113.985 134.785 ;
        RECT 108.620 134.600 113.985 134.740 ;
        RECT 108.620 134.540 108.940 134.600 ;
        RECT 113.695 134.555 113.985 134.600 ;
        RECT 116.915 134.555 117.205 134.785 ;
        RECT 117.360 134.740 117.680 134.800 ;
        RECT 128.400 134.785 128.720 134.800 ;
        RECT 118.195 134.740 118.485 134.785 ;
        RECT 117.360 134.600 118.485 134.740 ;
        RECT 117.360 134.540 117.680 134.600 ;
        RECT 118.195 134.555 118.485 134.600 ;
        RECT 128.370 134.555 128.720 134.785 ;
        RECT 131.710 134.740 131.850 134.940 ;
        RECT 131.710 134.600 132.310 134.740 ;
        RECT 128.400 134.540 128.720 134.555 ;
        RECT 77.815 134.215 78.105 134.445 ;
        RECT 78.720 134.400 79.040 134.460 ;
        RECT 82.375 134.400 82.665 134.445 ;
        RECT 83.565 134.400 83.855 134.445 ;
        RECT 86.085 134.400 86.375 134.445 ;
        RECT 78.720 134.260 81.710 134.400 ;
        RECT 76.895 134.060 77.185 134.105 ;
        RECT 77.890 134.060 78.030 134.215 ;
        RECT 78.720 134.200 79.040 134.260 ;
        RECT 76.895 133.920 78.030 134.060 ;
        RECT 76.895 133.875 77.185 133.920 ;
        RECT 75.975 133.720 76.265 133.765 ;
        RECT 78.720 133.720 79.040 133.780 ;
        RECT 75.590 133.580 79.040 133.720 ;
        RECT 81.570 133.720 81.710 134.260 ;
        RECT 82.375 134.260 86.375 134.400 ;
        RECT 82.375 134.215 82.665 134.260 ;
        RECT 83.565 134.215 83.855 134.260 ;
        RECT 86.085 134.215 86.375 134.260 ;
        RECT 93.875 134.400 94.165 134.445 ;
        RECT 95.065 134.400 95.355 134.445 ;
        RECT 97.585 134.400 97.875 134.445 ;
        RECT 93.875 134.260 97.875 134.400 ;
        RECT 93.875 134.215 94.165 134.260 ;
        RECT 95.065 134.215 95.355 134.260 ;
        RECT 97.585 134.215 97.875 134.260 ;
        RECT 102.640 134.200 102.960 134.460 ;
        RECT 103.100 134.200 103.420 134.460 ;
        RECT 106.755 134.400 107.045 134.445 ;
        RECT 107.945 134.400 108.235 134.445 ;
        RECT 110.465 134.400 110.755 134.445 ;
        RECT 106.755 134.260 110.755 134.400 ;
        RECT 106.755 134.215 107.045 134.260 ;
        RECT 107.945 134.215 108.235 134.260 ;
        RECT 110.465 134.215 110.755 134.260 ;
        RECT 117.795 134.400 118.085 134.445 ;
        RECT 118.985 134.400 119.275 134.445 ;
        RECT 121.505 134.400 121.795 134.445 ;
        RECT 117.795 134.260 121.795 134.400 ;
        RECT 117.795 134.215 118.085 134.260 ;
        RECT 118.985 134.215 119.275 134.260 ;
        RECT 121.505 134.215 121.795 134.260 ;
        RECT 127.020 134.200 127.340 134.460 ;
        RECT 127.915 134.400 128.205 134.445 ;
        RECT 129.105 134.400 129.395 134.445 ;
        RECT 131.625 134.400 131.915 134.445 ;
        RECT 127.915 134.260 131.915 134.400 ;
        RECT 127.915 134.215 128.205 134.260 ;
        RECT 129.105 134.215 129.395 134.260 ;
        RECT 131.625 134.215 131.915 134.260 ;
        RECT 81.980 134.060 82.270 134.105 ;
        RECT 84.080 134.060 84.370 134.105 ;
        RECT 85.650 134.060 85.940 134.105 ;
        RECT 81.980 133.920 85.940 134.060 ;
        RECT 81.980 133.875 82.270 133.920 ;
        RECT 84.080 133.875 84.370 133.920 ;
        RECT 85.650 133.875 85.940 133.920 ;
        RECT 93.480 134.060 93.770 134.105 ;
        RECT 95.580 134.060 95.870 134.105 ;
        RECT 97.150 134.060 97.440 134.105 ;
        RECT 93.480 133.920 97.440 134.060 ;
        RECT 93.480 133.875 93.770 133.920 ;
        RECT 95.580 133.875 95.870 133.920 ;
        RECT 97.150 133.875 97.440 133.920 ;
        RECT 106.360 134.060 106.650 134.105 ;
        RECT 108.460 134.060 108.750 134.105 ;
        RECT 110.030 134.060 110.320 134.105 ;
        RECT 106.360 133.920 110.320 134.060 ;
        RECT 106.360 133.875 106.650 133.920 ;
        RECT 108.460 133.875 108.750 133.920 ;
        RECT 110.030 133.875 110.320 133.920 ;
        RECT 111.380 134.060 111.700 134.120 ;
        RECT 116.900 134.060 117.220 134.120 ;
        RECT 111.380 133.920 117.220 134.060 ;
        RECT 111.380 133.860 111.700 133.920 ;
        RECT 116.900 133.860 117.220 133.920 ;
        RECT 117.400 134.060 117.690 134.105 ;
        RECT 119.500 134.060 119.790 134.105 ;
        RECT 121.070 134.060 121.360 134.105 ;
        RECT 126.100 134.060 126.420 134.120 ;
        RECT 117.400 133.920 121.360 134.060 ;
        RECT 117.400 133.875 117.690 133.920 ;
        RECT 119.500 133.875 119.790 133.920 ;
        RECT 121.070 133.875 121.360 133.920 ;
        RECT 121.590 133.920 126.420 134.060 ;
        RECT 86.080 133.720 86.400 133.780 ;
        RECT 87.920 133.720 88.240 133.780 ;
        RECT 81.570 133.580 88.240 133.720 ;
        RECT 31.800 133.520 32.120 133.580 ;
        RECT 35.940 133.520 36.260 133.580 ;
        RECT 52.500 133.520 52.820 133.580 ;
        RECT 75.975 133.535 76.265 133.580 ;
        RECT 78.720 133.520 79.040 133.580 ;
        RECT 86.080 133.520 86.400 133.580 ;
        RECT 87.920 133.520 88.240 133.580 ;
        RECT 88.395 133.720 88.685 133.765 ;
        RECT 90.680 133.720 91.000 133.780 ;
        RECT 94.820 133.720 95.140 133.780 ;
        RECT 88.395 133.580 95.140 133.720 ;
        RECT 88.395 133.535 88.685 133.580 ;
        RECT 90.680 133.520 91.000 133.580 ;
        RECT 94.820 133.520 95.140 133.580 ;
        RECT 100.340 133.520 100.660 133.780 ;
        RECT 110.460 133.720 110.780 133.780 ;
        RECT 114.155 133.720 114.445 133.765 ;
        RECT 110.460 133.580 114.445 133.720 ;
        RECT 110.460 133.520 110.780 133.580 ;
        RECT 114.155 133.535 114.445 133.580 ;
        RECT 118.280 133.720 118.600 133.780 ;
        RECT 121.590 133.720 121.730 133.920 ;
        RECT 126.100 133.860 126.420 133.920 ;
        RECT 127.520 134.060 127.810 134.105 ;
        RECT 129.620 134.060 129.910 134.105 ;
        RECT 131.190 134.060 131.480 134.105 ;
        RECT 127.520 133.920 131.480 134.060 ;
        RECT 132.170 134.060 132.310 134.600 ;
        RECT 135.760 134.540 136.080 134.800 ;
        RECT 133.935 134.060 134.225 134.105 ;
        RECT 135.760 134.060 136.080 134.120 ;
        RECT 132.170 133.920 136.080 134.060 ;
        RECT 127.520 133.875 127.810 133.920 ;
        RECT 129.620 133.875 129.910 133.920 ;
        RECT 131.190 133.875 131.480 133.920 ;
        RECT 133.935 133.875 134.225 133.920 ;
        RECT 135.760 133.860 136.080 133.920 ;
        RECT 118.280 133.580 121.730 133.720 ;
        RECT 123.800 133.720 124.120 133.780 ;
        RECT 134.380 133.720 134.700 133.780 ;
        RECT 123.800 133.580 134.700 133.720 ;
        RECT 118.280 133.520 118.600 133.580 ;
        RECT 123.800 133.520 124.120 133.580 ;
        RECT 134.380 133.520 134.700 133.580 ;
        RECT 13.330 132.900 138.910 133.380 ;
        RECT 24.900 132.500 25.220 132.760 ;
        RECT 27.675 132.700 27.965 132.745 ;
        RECT 31.800 132.700 32.120 132.760 ;
        RECT 27.675 132.560 32.120 132.700 ;
        RECT 27.675 132.515 27.965 132.560 ;
        RECT 31.800 132.500 32.120 132.560 ;
        RECT 34.115 132.700 34.405 132.745 ;
        RECT 35.480 132.700 35.800 132.760 ;
        RECT 34.115 132.560 35.800 132.700 ;
        RECT 34.115 132.515 34.405 132.560 ;
        RECT 35.480 132.500 35.800 132.560 ;
        RECT 41.460 132.500 41.780 132.760 ;
        RECT 44.220 132.700 44.540 132.760 ;
        RECT 44.695 132.700 44.985 132.745 ;
        RECT 42.470 132.560 43.990 132.700 ;
        RECT 18.500 132.360 18.790 132.405 ;
        RECT 20.600 132.360 20.890 132.405 ;
        RECT 22.170 132.360 22.460 132.405 ;
        RECT 18.500 132.220 22.460 132.360 ;
        RECT 18.500 132.175 18.790 132.220 ;
        RECT 20.600 132.175 20.890 132.220 ;
        RECT 22.170 132.175 22.460 132.220 ;
        RECT 35.060 132.360 35.350 132.405 ;
        RECT 37.160 132.360 37.450 132.405 ;
        RECT 38.730 132.360 39.020 132.405 ;
        RECT 35.060 132.220 39.020 132.360 ;
        RECT 35.060 132.175 35.350 132.220 ;
        RECT 37.160 132.175 37.450 132.220 ;
        RECT 38.730 132.175 39.020 132.220 ;
        RECT 18.895 132.020 19.185 132.065 ;
        RECT 20.085 132.020 20.375 132.065 ;
        RECT 22.605 132.020 22.895 132.065 ;
        RECT 29.515 132.020 29.805 132.065 ;
        RECT 31.340 132.020 31.660 132.080 ;
        RECT 32.735 132.020 33.025 132.065 ;
        RECT 35.455 132.020 35.745 132.065 ;
        RECT 36.645 132.020 36.935 132.065 ;
        RECT 39.165 132.020 39.455 132.065 ;
        RECT 18.895 131.880 22.895 132.020 ;
        RECT 18.895 131.835 19.185 131.880 ;
        RECT 20.085 131.835 20.375 131.880 ;
        RECT 22.605 131.835 22.895 131.880 ;
        RECT 28.210 131.880 29.805 132.020 ;
        RECT 18.015 131.680 18.305 131.725 ;
        RECT 23.060 131.680 23.380 131.740 ;
        RECT 18.015 131.540 23.380 131.680 ;
        RECT 18.015 131.495 18.305 131.540 ;
        RECT 23.060 131.480 23.380 131.540 ;
        RECT 19.350 131.340 19.640 131.385 ;
        RECT 23.980 131.340 24.300 131.400 ;
        RECT 19.350 131.200 24.300 131.340 ;
        RECT 19.350 131.155 19.640 131.200 ;
        RECT 23.980 131.140 24.300 131.200 ;
        RECT 26.740 131.140 27.060 131.400 ;
        RECT 27.780 131.340 28.070 131.385 ;
        RECT 28.210 131.340 28.350 131.880 ;
        RECT 29.515 131.835 29.805 131.880 ;
        RECT 30.050 131.880 35.250 132.020 ;
        RECT 29.040 131.480 29.360 131.740 ;
        RECT 30.050 131.725 30.190 131.880 ;
        RECT 31.340 131.820 31.660 131.880 ;
        RECT 32.735 131.835 33.025 131.880 ;
        RECT 29.975 131.495 30.265 131.725 ;
        RECT 32.275 131.680 32.565 131.725 ;
        RECT 34.100 131.680 34.420 131.740 ;
        RECT 32.275 131.540 34.420 131.680 ;
        RECT 32.275 131.495 32.565 131.540 ;
        RECT 34.100 131.480 34.420 131.540 ;
        RECT 34.575 131.495 34.865 131.725 ;
        RECT 35.110 131.680 35.250 131.880 ;
        RECT 35.455 131.880 39.455 132.020 ;
        RECT 35.455 131.835 35.745 131.880 ;
        RECT 36.645 131.835 36.935 131.880 ;
        RECT 39.165 131.835 39.455 131.880 ;
        RECT 41.935 131.680 42.225 131.725 ;
        RECT 42.470 131.680 42.610 132.560 ;
        RECT 43.315 132.175 43.605 132.405 ;
        RECT 35.110 131.540 42.610 131.680 ;
        RECT 43.390 131.680 43.530 132.175 ;
        RECT 43.850 132.020 43.990 132.560 ;
        RECT 44.220 132.560 44.985 132.700 ;
        RECT 44.220 132.500 44.540 132.560 ;
        RECT 44.695 132.515 44.985 132.560 ;
        RECT 46.980 132.500 47.300 132.760 ;
        RECT 47.915 132.700 48.205 132.745 ;
        RECT 49.280 132.700 49.600 132.760 ;
        RECT 47.915 132.560 49.600 132.700 ;
        RECT 47.915 132.515 48.205 132.560 ;
        RECT 49.280 132.500 49.600 132.560 ;
        RECT 50.675 132.515 50.965 132.745 ;
        RECT 51.595 132.700 51.885 132.745 ;
        RECT 52.040 132.700 52.360 132.760 ;
        RECT 51.595 132.560 52.360 132.700 ;
        RECT 51.595 132.515 51.885 132.560 ;
        RECT 45.615 132.360 45.905 132.405 ;
        RECT 50.200 132.360 50.520 132.420 ;
        RECT 45.615 132.220 50.520 132.360 ;
        RECT 50.750 132.360 50.890 132.515 ;
        RECT 52.040 132.500 52.360 132.560 ;
        RECT 66.760 132.700 67.080 132.760 ;
        RECT 67.695 132.700 67.985 132.745 ;
        RECT 66.760 132.560 67.985 132.700 ;
        RECT 66.760 132.500 67.080 132.560 ;
        RECT 67.695 132.515 67.985 132.560 ;
        RECT 72.280 132.500 72.600 132.760 ;
        RECT 78.720 132.700 79.040 132.760 ;
        RECT 79.195 132.700 79.485 132.745 ;
        RECT 78.720 132.560 79.485 132.700 ;
        RECT 78.720 132.500 79.040 132.560 ;
        RECT 79.195 132.515 79.485 132.560 ;
        RECT 81.495 132.700 81.785 132.745 ;
        RECT 81.940 132.700 82.260 132.760 ;
        RECT 81.495 132.560 82.260 132.700 ;
        RECT 81.495 132.515 81.785 132.560 ;
        RECT 52.500 132.360 52.820 132.420 ;
        RECT 73.200 132.360 73.520 132.420 ;
        RECT 50.750 132.220 52.820 132.360 ;
        RECT 45.615 132.175 45.905 132.220 ;
        RECT 50.200 132.160 50.520 132.220 ;
        RECT 52.500 132.160 52.820 132.220 ;
        RECT 69.840 132.220 73.520 132.360 ;
        RECT 79.270 132.360 79.410 132.515 ;
        RECT 81.940 132.500 82.260 132.560 ;
        RECT 82.830 132.515 83.120 132.745 ;
        RECT 99.880 132.700 100.200 132.760 ;
        RECT 101.275 132.700 101.565 132.745 ;
        RECT 99.880 132.560 101.565 132.700 ;
        RECT 82.400 132.360 82.720 132.420 ;
        RECT 82.905 132.360 83.045 132.515 ;
        RECT 99.880 132.500 100.200 132.560 ;
        RECT 101.275 132.515 101.565 132.560 ;
        RECT 79.270 132.220 83.045 132.360 ;
        RECT 84.740 132.360 85.030 132.405 ;
        RECT 86.840 132.360 87.130 132.405 ;
        RECT 88.410 132.360 88.700 132.405 ;
        RECT 84.740 132.220 88.700 132.360 ;
        RECT 47.900 132.020 48.220 132.080 ;
        RECT 50.660 132.020 50.980 132.080 ;
        RECT 43.850 131.880 48.220 132.020 ;
        RECT 47.900 131.820 48.220 131.880 ;
        RECT 49.830 131.880 50.980 132.020 ;
        RECT 48.375 131.680 48.665 131.725 ;
        RECT 43.390 131.540 48.665 131.680 ;
        RECT 41.935 131.495 42.225 131.540 ;
        RECT 48.375 131.495 48.665 131.540 ;
        RECT 27.780 131.200 28.350 131.340 ;
        RECT 29.500 131.340 29.820 131.400 ;
        RECT 34.650 131.340 34.790 131.495 ;
        RECT 48.820 131.480 49.140 131.740 ;
        RECT 49.280 131.480 49.600 131.740 ;
        RECT 29.500 131.200 34.790 131.340 ;
        RECT 35.910 131.340 36.200 131.385 ;
        RECT 36.400 131.340 36.720 131.400 ;
        RECT 35.910 131.200 36.720 131.340 ;
        RECT 27.780 131.155 28.070 131.200 ;
        RECT 29.500 131.140 29.820 131.200 ;
        RECT 35.910 131.155 36.200 131.200 ;
        RECT 36.400 131.140 36.720 131.200 ;
        RECT 41.460 131.340 41.780 131.400 ;
        RECT 42.395 131.340 42.685 131.385 ;
        RECT 41.460 131.200 42.685 131.340 ;
        RECT 41.460 131.140 41.780 131.200 ;
        RECT 42.395 131.155 42.685 131.200 ;
        RECT 43.315 131.155 43.605 131.385 ;
        RECT 28.580 130.800 28.900 131.060 ;
        RECT 43.390 131.000 43.530 131.155 ;
        RECT 43.760 131.140 44.080 131.400 ;
        RECT 44.680 131.385 45.000 131.400 ;
        RECT 44.680 131.155 45.065 131.385 ;
        RECT 44.680 131.140 45.000 131.155 ;
        RECT 46.060 131.140 46.380 131.400 ;
        RECT 49.830 131.385 49.970 131.880 ;
        RECT 50.660 131.820 50.980 131.880 ;
        RECT 68.615 131.680 68.905 131.725 ;
        RECT 69.840 131.680 69.980 132.220 ;
        RECT 73.200 132.160 73.520 132.220 ;
        RECT 82.400 132.160 82.720 132.220 ;
        RECT 84.740 132.175 85.030 132.220 ;
        RECT 86.840 132.175 87.130 132.220 ;
        RECT 88.410 132.175 88.700 132.220 ;
        RECT 94.860 132.360 95.150 132.405 ;
        RECT 96.960 132.360 97.250 132.405 ;
        RECT 98.530 132.360 98.820 132.405 ;
        RECT 94.860 132.220 98.820 132.360 ;
        RECT 94.860 132.175 95.150 132.220 ;
        RECT 96.960 132.175 97.250 132.220 ;
        RECT 98.530 132.175 98.820 132.220 ;
        RECT 74.120 132.020 74.440 132.080 ;
        RECT 80.115 132.020 80.405 132.065 ;
        RECT 70.990 131.880 80.405 132.020 ;
        RECT 70.990 131.740 71.130 131.880 ;
        RECT 74.120 131.820 74.440 131.880 ;
        RECT 80.115 131.835 80.405 131.880 ;
        RECT 81.480 132.020 81.800 132.080 ;
        RECT 84.255 132.020 84.545 132.065 ;
        RECT 81.480 131.880 84.545 132.020 ;
        RECT 68.615 131.540 69.980 131.680 ;
        RECT 68.615 131.495 68.905 131.540 ;
        RECT 70.900 131.480 71.220 131.740 ;
        RECT 71.835 131.680 72.125 131.725 ;
        RECT 73.215 131.680 73.505 131.725 ;
        RECT 71.835 131.540 73.505 131.680 ;
        RECT 71.835 131.495 72.125 131.540 ;
        RECT 73.215 131.495 73.505 131.540 ;
        RECT 73.660 131.480 73.980 131.740 ;
        RECT 75.960 131.680 76.280 131.740 ;
        RECT 78.735 131.680 79.025 131.725 ;
        RECT 74.210 131.540 79.025 131.680 ;
        RECT 51.120 131.385 51.440 131.400 ;
        RECT 49.755 131.155 50.045 131.385 ;
        RECT 50.835 131.155 51.440 131.385 ;
        RECT 51.120 131.140 51.440 131.155 ;
        RECT 68.140 131.340 68.460 131.400 ;
        RECT 69.535 131.340 69.825 131.385 ;
        RECT 68.140 131.200 69.825 131.340 ;
        RECT 68.140 131.140 68.460 131.200 ;
        RECT 69.535 131.155 69.825 131.200 ;
        RECT 69.980 131.140 70.300 131.400 ;
        RECT 46.150 131.000 46.290 131.140 ;
        RECT 43.390 130.860 46.290 131.000 ;
        RECT 47.125 131.000 47.415 131.045 ;
        RECT 47.900 131.000 48.220 131.060 ;
        RECT 47.125 130.860 48.220 131.000 ;
        RECT 70.070 131.000 70.210 131.140 ;
        RECT 74.210 131.000 74.350 131.540 ;
        RECT 75.960 131.480 76.280 131.540 ;
        RECT 78.735 131.495 79.025 131.540 ;
        RECT 80.190 131.340 80.330 131.835 ;
        RECT 81.480 131.820 81.800 131.880 ;
        RECT 84.255 131.835 84.545 131.880 ;
        RECT 85.135 132.020 85.425 132.065 ;
        RECT 86.325 132.020 86.615 132.065 ;
        RECT 88.845 132.020 89.135 132.065 ;
        RECT 85.135 131.880 89.135 132.020 ;
        RECT 85.135 131.835 85.425 131.880 ;
        RECT 86.325 131.835 86.615 131.880 ;
        RECT 88.845 131.835 89.135 131.880 ;
        RECT 92.980 132.020 93.300 132.080 ;
        RECT 94.375 132.020 94.665 132.065 ;
        RECT 92.980 131.880 94.665 132.020 ;
        RECT 92.980 131.820 93.300 131.880 ;
        RECT 94.375 131.835 94.665 131.880 ;
        RECT 95.255 132.020 95.545 132.065 ;
        RECT 96.445 132.020 96.735 132.065 ;
        RECT 98.965 132.020 99.255 132.065 ;
        RECT 95.255 131.880 99.255 132.020 ;
        RECT 101.350 132.020 101.490 132.515 ;
        RECT 104.020 132.500 104.340 132.760 ;
        RECT 107.240 132.700 107.560 132.760 ;
        RECT 107.715 132.700 108.005 132.745 ;
        RECT 107.240 132.560 108.005 132.700 ;
        RECT 107.240 132.500 107.560 132.560 ;
        RECT 107.715 132.515 108.005 132.560 ;
        RECT 116.455 132.700 116.745 132.745 ;
        RECT 117.360 132.700 117.680 132.760 ;
        RECT 116.455 132.560 117.680 132.700 ;
        RECT 116.455 132.515 116.745 132.560 ;
        RECT 117.360 132.500 117.680 132.560 ;
        RECT 122.420 132.700 122.740 132.760 ;
        RECT 122.420 132.560 132.770 132.700 ;
        RECT 122.420 132.500 122.740 132.560 ;
        RECT 102.640 132.360 102.960 132.420 ;
        RECT 111.395 132.360 111.685 132.405 ;
        RECT 118.740 132.360 119.060 132.420 ;
        RECT 102.640 132.220 107.930 132.360 ;
        RECT 102.640 132.160 102.960 132.220 ;
        RECT 106.795 132.020 107.085 132.065 ;
        RECT 101.350 131.880 107.085 132.020 ;
        RECT 107.790 132.020 107.930 132.220 ;
        RECT 109.630 132.220 111.685 132.360 ;
        RECT 109.630 132.020 109.770 132.220 ;
        RECT 111.395 132.175 111.685 132.220 ;
        RECT 118.140 132.220 119.060 132.360 ;
        RECT 107.790 131.880 109.770 132.020 ;
        RECT 110.460 132.020 110.780 132.080 ;
        RECT 114.600 132.020 114.920 132.080 ;
        RECT 118.140 132.020 118.280 132.220 ;
        RECT 118.740 132.160 119.060 132.220 ;
        RECT 125.640 132.360 125.960 132.420 ;
        RECT 132.095 132.360 132.385 132.405 ;
        RECT 125.640 132.220 132.385 132.360 ;
        RECT 125.640 132.160 125.960 132.220 ;
        RECT 132.095 132.175 132.385 132.220 ;
        RECT 120.135 132.020 120.425 132.065 ;
        RECT 123.800 132.020 124.120 132.080 ;
        RECT 110.460 131.880 112.530 132.020 ;
        RECT 95.255 131.835 95.545 131.880 ;
        RECT 96.445 131.835 96.735 131.880 ;
        RECT 98.965 131.835 99.255 131.880 ;
        RECT 106.795 131.835 107.085 131.880 ;
        RECT 110.460 131.820 110.780 131.880 ;
        RECT 95.710 131.680 96.000 131.725 ;
        RECT 100.340 131.680 100.660 131.740 ;
        RECT 95.710 131.540 100.660 131.680 ;
        RECT 95.710 131.495 96.000 131.540 ;
        RECT 100.340 131.480 100.660 131.540 ;
        RECT 109.080 131.480 109.400 131.740 ;
        RECT 109.555 131.495 109.845 131.725 ;
        RECT 80.560 131.340 80.880 131.400 ;
        RECT 81.955 131.340 82.245 131.385 ;
        RECT 80.190 131.200 82.245 131.340 ;
        RECT 80.560 131.140 80.880 131.200 ;
        RECT 81.955 131.155 82.245 131.200 ;
        RECT 84.700 131.340 85.020 131.400 ;
        RECT 85.480 131.340 85.770 131.385 ;
        RECT 84.700 131.200 85.770 131.340 ;
        RECT 84.700 131.140 85.020 131.200 ;
        RECT 85.480 131.155 85.770 131.200 ;
        RECT 94.820 131.340 95.140 131.400 ;
        RECT 109.630 131.340 109.770 131.495 ;
        RECT 110.000 131.480 110.320 131.740 ;
        RECT 112.390 131.725 112.530 131.880 ;
        RECT 112.850 131.880 114.920 132.020 ;
        RECT 112.850 131.725 112.990 131.880 ;
        RECT 114.600 131.820 114.920 131.880 ;
        RECT 117.910 131.880 118.280 132.020 ;
        RECT 118.830 131.880 120.425 132.020 ;
        RECT 110.935 131.495 111.225 131.725 ;
        RECT 112.315 131.495 112.605 131.725 ;
        RECT 112.775 131.495 113.065 131.725 ;
        RECT 111.010 131.340 111.150 131.495 ;
        RECT 113.680 131.480 114.000 131.740 ;
        RECT 114.155 131.680 114.445 131.725 ;
        RECT 115.060 131.680 115.380 131.740 ;
        RECT 114.155 131.540 115.380 131.680 ;
        RECT 114.155 131.495 114.445 131.540 ;
        RECT 115.060 131.480 115.380 131.540 ;
        RECT 115.520 131.680 115.840 131.740 ;
        RECT 117.910 131.725 118.050 131.880 ;
        RECT 117.835 131.680 118.125 131.725 ;
        RECT 115.520 131.540 118.125 131.680 ;
        RECT 115.520 131.480 115.840 131.540 ;
        RECT 117.835 131.495 118.125 131.540 ;
        RECT 118.280 131.480 118.600 131.740 ;
        RECT 118.830 131.725 118.970 131.880 ;
        RECT 120.135 131.835 120.425 131.880 ;
        RECT 121.130 131.880 124.120 132.020 ;
        RECT 118.755 131.495 119.045 131.725 ;
        RECT 119.660 131.480 119.980 131.740 ;
        RECT 121.130 131.725 121.270 131.880 ;
        RECT 123.800 131.820 124.120 131.880 ;
        RECT 124.720 132.020 125.040 132.080 ;
        RECT 126.100 132.020 126.420 132.080 ;
        RECT 124.720 131.880 125.870 132.020 ;
        RECT 124.720 131.820 125.040 131.880 ;
        RECT 125.730 131.725 125.870 131.880 ;
        RECT 126.100 131.880 127.250 132.020 ;
        RECT 126.100 131.820 126.420 131.880 ;
        RECT 127.110 131.725 127.250 131.880 ;
        RECT 128.875 131.835 129.165 132.065 ;
        RECT 132.630 132.020 132.770 132.560 ;
        RECT 136.680 132.500 137.000 132.760 ;
        RECT 131.710 131.880 134.150 132.020 ;
        RECT 121.055 131.495 121.345 131.725 ;
        RECT 125.655 131.495 125.945 131.725 ;
        RECT 126.575 131.495 126.865 131.725 ;
        RECT 127.035 131.495 127.325 131.725 ;
        RECT 116.900 131.340 117.220 131.400 ;
        RECT 94.820 131.200 110.690 131.340 ;
        RECT 111.010 131.200 117.220 131.340 ;
        RECT 94.820 131.140 95.140 131.200 ;
        RECT 70.070 130.860 74.350 131.000 ;
        RECT 82.400 131.000 82.720 131.060 ;
        RECT 82.955 131.000 83.245 131.045 ;
        RECT 82.400 130.860 83.245 131.000 ;
        RECT 47.125 130.815 47.415 130.860 ;
        RECT 47.900 130.800 48.220 130.860 ;
        RECT 82.400 130.800 82.720 130.860 ;
        RECT 82.955 130.815 83.245 130.860 ;
        RECT 83.795 131.000 84.085 131.045 ;
        RECT 87.460 131.000 87.780 131.060 ;
        RECT 83.795 130.860 87.780 131.000 ;
        RECT 83.795 130.815 84.085 130.860 ;
        RECT 87.460 130.800 87.780 130.860 ;
        RECT 91.155 131.000 91.445 131.045 ;
        RECT 93.440 131.000 93.760 131.060 ;
        RECT 91.155 130.860 93.760 131.000 ;
        RECT 110.550 131.000 110.690 131.200 ;
        RECT 112.850 131.060 112.990 131.200 ;
        RECT 116.900 131.140 117.220 131.200 ;
        RECT 121.975 131.340 122.265 131.385 ;
        RECT 122.420 131.340 122.740 131.400 ;
        RECT 121.975 131.200 122.740 131.340 ;
        RECT 126.650 131.340 126.790 131.495 ;
        RECT 127.480 131.480 127.800 131.740 ;
        RECT 128.400 131.680 128.720 131.740 ;
        RECT 128.950 131.680 129.090 131.835 ;
        RECT 131.710 131.725 131.850 131.880 ;
        RECT 128.400 131.540 129.090 131.680 ;
        RECT 128.400 131.480 128.720 131.540 ;
        RECT 131.635 131.495 131.925 131.725 ;
        RECT 129.795 131.340 130.085 131.385 ;
        RECT 126.650 131.200 130.085 131.340 ;
        RECT 121.975 131.155 122.265 131.200 ;
        RECT 122.420 131.140 122.740 131.200 ;
        RECT 129.795 131.155 130.085 131.200 ;
        RECT 130.700 131.140 131.020 131.400 ;
        RECT 132.080 131.340 132.400 131.400 ;
        RECT 134.010 131.385 134.150 131.880 ;
        RECT 134.380 131.680 134.700 131.740 ;
        RECT 135.775 131.680 136.065 131.725 ;
        RECT 134.380 131.540 136.065 131.680 ;
        RECT 134.380 131.480 134.700 131.540 ;
        RECT 135.775 131.495 136.065 131.540 ;
        RECT 133.015 131.340 133.305 131.385 ;
        RECT 132.080 131.200 133.305 131.340 ;
        RECT 132.080 131.140 132.400 131.200 ;
        RECT 133.015 131.155 133.305 131.200 ;
        RECT 133.935 131.155 134.225 131.385 ;
        RECT 110.920 131.000 111.240 131.060 ;
        RECT 110.550 130.860 111.240 131.000 ;
        RECT 91.155 130.815 91.445 130.860 ;
        RECT 93.440 130.800 93.760 130.860 ;
        RECT 110.920 130.800 111.240 130.860 ;
        RECT 112.760 130.800 113.080 131.060 ;
        RECT 13.330 130.180 138.910 130.660 ;
        RECT 22.155 129.980 22.445 130.025 ;
        RECT 25.820 129.980 26.140 130.040 ;
        RECT 22.155 129.840 26.140 129.980 ;
        RECT 22.155 129.795 22.445 129.840 ;
        RECT 25.820 129.780 26.140 129.840 ;
        RECT 26.740 129.980 27.060 130.040 ;
        RECT 35.035 129.980 35.325 130.025 ;
        RECT 36.400 129.980 36.720 130.040 ;
        RECT 26.740 129.840 30.485 129.980 ;
        RECT 26.740 129.780 27.060 129.840 ;
        RECT 23.060 129.640 23.380 129.700 ;
        RECT 29.500 129.640 29.820 129.700 ;
        RECT 23.060 129.500 29.820 129.640 ;
        RECT 23.060 129.440 23.380 129.500 ;
        RECT 27.775 129.300 28.065 129.345 ;
        RECT 28.580 129.300 28.900 129.360 ;
        RECT 29.130 129.345 29.270 129.500 ;
        RECT 29.500 129.440 29.820 129.500 ;
        RECT 27.775 129.160 28.900 129.300 ;
        RECT 27.775 129.115 28.065 129.160 ;
        RECT 28.580 129.100 28.900 129.160 ;
        RECT 29.055 129.115 29.345 129.345 ;
        RECT 30.345 129.300 30.485 129.840 ;
        RECT 35.035 129.840 36.720 129.980 ;
        RECT 35.035 129.795 35.325 129.840 ;
        RECT 36.400 129.780 36.720 129.840 ;
        RECT 43.775 129.980 44.065 130.025 ;
        RECT 45.140 129.980 45.460 130.040 ;
        RECT 43.775 129.840 45.460 129.980 ;
        RECT 43.775 129.795 44.065 129.840 ;
        RECT 45.140 129.780 45.460 129.840 ;
        RECT 45.615 129.980 45.905 130.025 ;
        RECT 46.060 129.980 46.380 130.040 ;
        RECT 45.615 129.840 46.380 129.980 ;
        RECT 45.615 129.795 45.905 129.840 ;
        RECT 35.480 129.685 35.800 129.700 ;
        RECT 35.480 129.455 36.085 129.685 ;
        RECT 36.875 129.640 37.165 129.685 ;
        RECT 43.300 129.640 43.620 129.700 ;
        RECT 36.875 129.500 43.620 129.640 ;
        RECT 36.875 129.455 37.165 129.500 ;
        RECT 35.480 129.440 35.800 129.455 ;
        RECT 36.950 129.300 37.090 129.455 ;
        RECT 43.300 129.440 43.620 129.500 ;
        RECT 30.345 129.160 37.090 129.300 ;
        RECT 41.935 129.300 42.225 129.345 ;
        RECT 45.690 129.300 45.830 129.795 ;
        RECT 46.060 129.780 46.380 129.840 ;
        RECT 65.855 129.980 66.145 130.025 ;
        RECT 69.520 129.980 69.840 130.040 ;
        RECT 65.855 129.840 69.840 129.980 ;
        RECT 65.855 129.795 66.145 129.840 ;
        RECT 69.520 129.780 69.840 129.840 ;
        RECT 70.915 129.980 71.205 130.025 ;
        RECT 73.660 129.980 73.980 130.040 ;
        RECT 70.915 129.840 73.980 129.980 ;
        RECT 70.915 129.795 71.205 129.840 ;
        RECT 73.660 129.780 73.980 129.840 ;
        RECT 79.655 129.980 79.945 130.025 ;
        RECT 82.400 129.980 82.720 130.040 ;
        RECT 79.655 129.840 82.720 129.980 ;
        RECT 79.655 129.795 79.945 129.840 ;
        RECT 82.400 129.780 82.720 129.840 ;
        RECT 84.700 129.780 85.020 130.040 ;
        RECT 90.220 129.980 90.540 130.040 ;
        RECT 108.160 129.980 108.480 130.040 ;
        RECT 115.520 129.980 115.840 130.040 ;
        RECT 119.200 129.980 119.520 130.040 ;
        RECT 121.040 129.980 121.360 130.040 ;
        RECT 90.220 129.840 108.480 129.980 ;
        RECT 90.220 129.780 90.540 129.840 ;
        RECT 108.160 129.780 108.480 129.840 ;
        RECT 114.690 129.840 115.840 129.980 ;
        RECT 50.200 129.640 50.520 129.700 ;
        RECT 51.180 129.640 51.470 129.685 ;
        RECT 62.620 129.640 62.940 129.700 ;
        RECT 81.020 129.640 81.340 129.700 ;
        RECT 91.140 129.640 91.460 129.700 ;
        RECT 114.690 129.640 114.830 129.840 ;
        RECT 115.520 129.780 115.840 129.840 ;
        RECT 117.910 129.840 121.360 129.980 ;
        RECT 117.910 129.685 118.050 129.840 ;
        RECT 119.200 129.780 119.520 129.840 ;
        RECT 121.040 129.780 121.360 129.840 ;
        RECT 126.100 129.980 126.420 130.040 ;
        RECT 131.160 129.980 131.480 130.040 ;
        RECT 126.100 129.840 131.480 129.980 ;
        RECT 126.100 129.780 126.420 129.840 ;
        RECT 131.160 129.780 131.480 129.840 ;
        RECT 136.680 129.780 137.000 130.040 ;
        RECT 116.915 129.640 117.205 129.685 ;
        RECT 50.200 129.500 51.470 129.640 ;
        RECT 50.200 129.440 50.520 129.500 ;
        RECT 51.180 129.455 51.470 129.500 ;
        RECT 52.590 129.500 62.940 129.640 ;
        RECT 52.590 129.345 52.730 129.500 ;
        RECT 62.620 129.440 62.940 129.500 ;
        RECT 63.170 129.500 91.460 129.640 ;
        RECT 41.935 129.160 45.830 129.300 ;
        RECT 41.935 129.115 42.225 129.160 ;
        RECT 52.515 129.115 52.805 129.345 ;
        RECT 56.180 129.300 56.500 129.360 ;
        RECT 58.955 129.300 59.245 129.345 ;
        RECT 63.170 129.300 63.310 129.500 ;
        RECT 81.020 129.440 81.340 129.500 ;
        RECT 91.140 129.440 91.460 129.500 ;
        RECT 93.530 129.500 114.830 129.640 ;
        RECT 115.150 129.500 117.205 129.640 ;
        RECT 93.530 129.360 93.670 129.500 ;
        RECT 56.180 129.160 63.310 129.300 ;
        RECT 64.000 129.300 64.320 129.360 ;
        RECT 65.395 129.300 65.685 129.345 ;
        RECT 64.000 129.160 65.685 129.300 ;
        RECT 56.180 129.100 56.500 129.160 ;
        RECT 58.955 129.115 59.245 129.160 ;
        RECT 64.000 129.100 64.320 129.160 ;
        RECT 65.395 129.115 65.685 129.160 ;
        RECT 66.315 129.115 66.605 129.345 ;
        RECT 68.155 129.115 68.445 129.345 ;
        RECT 24.465 128.960 24.755 129.005 ;
        RECT 26.985 128.960 27.275 129.005 ;
        RECT 28.175 128.960 28.465 129.005 ;
        RECT 24.465 128.820 28.465 128.960 ;
        RECT 24.465 128.775 24.755 128.820 ;
        RECT 26.985 128.775 27.275 128.820 ;
        RECT 28.175 128.775 28.465 128.820 ;
        RECT 41.460 128.760 41.780 129.020 ;
        RECT 47.925 128.960 48.215 129.005 ;
        RECT 50.445 128.960 50.735 129.005 ;
        RECT 51.635 128.960 51.925 129.005 ;
        RECT 47.925 128.820 51.925 128.960 ;
        RECT 47.925 128.775 48.215 128.820 ;
        RECT 50.445 128.775 50.735 128.820 ;
        RECT 51.635 128.775 51.925 128.820 ;
        RECT 24.900 128.620 25.190 128.665 ;
        RECT 26.470 128.620 26.760 128.665 ;
        RECT 28.570 128.620 28.860 128.665 ;
        RECT 24.900 128.480 28.860 128.620 ;
        RECT 24.900 128.435 25.190 128.480 ;
        RECT 26.470 128.435 26.760 128.480 ;
        RECT 28.570 128.435 28.860 128.480 ;
        RECT 48.360 128.620 48.650 128.665 ;
        RECT 49.930 128.620 50.220 128.665 ;
        RECT 52.030 128.620 52.320 128.665 ;
        RECT 48.360 128.480 52.320 128.620 ;
        RECT 66.390 128.620 66.530 129.115 ;
        RECT 68.230 128.960 68.370 129.115 ;
        RECT 69.060 129.100 69.380 129.360 ;
        RECT 69.980 129.100 70.300 129.360 ;
        RECT 70.900 129.100 71.220 129.360 ;
        RECT 79.195 129.115 79.485 129.345 ;
        RECT 76.420 128.960 76.740 129.020 ;
        RECT 79.270 128.960 79.410 129.115 ;
        RECT 80.560 129.100 80.880 129.360 ;
        RECT 81.940 129.100 82.260 129.360 ;
        RECT 86.555 129.300 86.845 129.345 ;
        RECT 93.440 129.300 93.760 129.360 ;
        RECT 86.555 129.160 93.760 129.300 ;
        RECT 86.555 129.115 86.845 129.160 ;
        RECT 93.440 129.100 93.760 129.160 ;
        RECT 99.435 129.300 99.725 129.345 ;
        RECT 102.640 129.300 102.960 129.360 ;
        RECT 114.230 129.345 114.370 129.500 ;
        RECT 115.150 129.345 115.290 129.500 ;
        RECT 116.915 129.455 117.205 129.500 ;
        RECT 117.835 129.455 118.125 129.685 ;
        RECT 118.755 129.640 119.045 129.685 ;
        RECT 124.260 129.640 124.580 129.700 ;
        RECT 118.755 129.500 124.580 129.640 ;
        RECT 118.755 129.455 119.045 129.500 ;
        RECT 124.260 129.440 124.580 129.500 ;
        RECT 99.435 129.160 102.960 129.300 ;
        RECT 99.435 129.115 99.725 129.160 ;
        RECT 102.640 129.100 102.960 129.160 ;
        RECT 114.155 129.115 114.445 129.345 ;
        RECT 114.615 129.115 114.905 129.345 ;
        RECT 115.075 129.115 115.365 129.345 ;
        RECT 115.995 129.300 116.285 129.345 ;
        RECT 119.660 129.300 119.980 129.360 ;
        RECT 124.720 129.300 125.040 129.360 ;
        RECT 115.995 129.160 118.280 129.300 ;
        RECT 115.995 129.115 116.285 129.160 ;
        RECT 68.230 128.820 79.410 128.960 ;
        RECT 76.420 128.760 76.740 128.820 ;
        RECT 68.140 128.620 68.460 128.680 ;
        RECT 66.390 128.480 68.460 128.620 ;
        RECT 48.360 128.435 48.650 128.480 ;
        RECT 49.930 128.435 50.220 128.480 ;
        RECT 52.030 128.435 52.320 128.480 ;
        RECT 68.140 128.420 68.460 128.480 ;
        RECT 35.940 128.080 36.260 128.340 ;
        RECT 68.600 128.080 68.920 128.340 ;
        RECT 79.270 128.280 79.410 128.820 ;
        RECT 86.080 128.960 86.400 129.020 ;
        RECT 87.015 128.960 87.305 129.005 ;
        RECT 86.080 128.820 87.305 128.960 ;
        RECT 86.080 128.760 86.400 128.820 ;
        RECT 87.015 128.775 87.305 128.820 ;
        RECT 87.460 128.760 87.780 129.020 ;
        RECT 99.880 128.760 100.200 129.020 ;
        RECT 100.815 128.960 101.105 129.005 ;
        RECT 103.100 128.960 103.420 129.020 ;
        RECT 100.815 128.820 103.420 128.960 ;
        RECT 114.690 128.960 114.830 129.115 ;
        RECT 117.360 128.960 117.680 129.020 ;
        RECT 114.690 128.820 117.680 128.960 ;
        RECT 118.140 128.960 118.280 129.160 ;
        RECT 119.660 129.160 125.040 129.300 ;
        RECT 119.660 129.100 119.980 129.160 ;
        RECT 124.720 129.100 125.040 129.160 ;
        RECT 125.640 129.100 125.960 129.360 ;
        RECT 126.190 129.345 126.330 129.780 ;
        RECT 127.955 129.640 128.245 129.685 ;
        RECT 129.640 129.640 129.930 129.685 ;
        RECT 127.955 129.500 129.930 129.640 ;
        RECT 127.955 129.455 128.245 129.500 ;
        RECT 129.640 129.455 129.930 129.500 ;
        RECT 126.115 129.115 126.405 129.345 ;
        RECT 126.560 129.300 126.880 129.360 ;
        RECT 128.860 129.300 129.180 129.360 ;
        RECT 135.775 129.300 136.065 129.345 ;
        RECT 126.560 129.160 129.180 129.300 ;
        RECT 126.560 129.100 126.880 129.160 ;
        RECT 128.860 129.100 129.180 129.160 ;
        RECT 135.390 129.160 136.065 129.300 ;
        RECT 119.750 128.960 119.890 129.100 ;
        RECT 128.415 128.960 128.705 129.005 ;
        RECT 118.140 128.820 119.890 128.960 ;
        RECT 127.110 128.820 128.705 128.960 ;
        RECT 100.815 128.775 101.105 128.820 ;
        RECT 103.100 128.760 103.420 128.820 ;
        RECT 117.360 128.760 117.680 128.820 ;
        RECT 127.110 128.680 127.250 128.820 ;
        RECT 128.415 128.775 128.705 128.820 ;
        RECT 129.295 128.960 129.585 129.005 ;
        RECT 130.485 128.960 130.775 129.005 ;
        RECT 133.005 128.960 133.295 129.005 ;
        RECT 129.295 128.820 133.295 128.960 ;
        RECT 129.295 128.775 129.585 128.820 ;
        RECT 130.485 128.775 130.775 128.820 ;
        RECT 133.005 128.775 133.295 128.820 ;
        RECT 107.700 128.620 108.020 128.680 ;
        RECT 109.080 128.620 109.400 128.680 ;
        RECT 126.560 128.620 126.880 128.680 ;
        RECT 107.700 128.480 126.880 128.620 ;
        RECT 107.700 128.420 108.020 128.480 ;
        RECT 109.080 128.420 109.400 128.480 ;
        RECT 126.560 128.420 126.880 128.480 ;
        RECT 127.020 128.420 127.340 128.680 ;
        RECT 128.900 128.620 129.190 128.665 ;
        RECT 131.000 128.620 131.290 128.665 ;
        RECT 132.570 128.620 132.860 128.665 ;
        RECT 128.900 128.480 132.860 128.620 ;
        RECT 128.900 128.435 129.190 128.480 ;
        RECT 131.000 128.435 131.290 128.480 ;
        RECT 132.570 128.435 132.860 128.480 ;
        RECT 81.035 128.280 81.325 128.325 ;
        RECT 79.270 128.140 81.325 128.280 ;
        RECT 81.035 128.095 81.325 128.140 ;
        RECT 83.335 128.280 83.625 128.325 ;
        RECT 89.760 128.280 90.080 128.340 ;
        RECT 83.335 128.140 90.080 128.280 ;
        RECT 83.335 128.095 83.625 128.140 ;
        RECT 89.760 128.080 90.080 128.140 ;
        RECT 97.120 128.280 97.440 128.340 ;
        RECT 97.595 128.280 97.885 128.325 ;
        RECT 97.120 128.140 97.885 128.280 ;
        RECT 97.120 128.080 97.440 128.140 ;
        RECT 97.595 128.095 97.885 128.140 ;
        RECT 112.760 128.080 113.080 128.340 ;
        RECT 132.080 128.280 132.400 128.340 ;
        RECT 135.390 128.325 135.530 129.160 ;
        RECT 135.775 129.115 136.065 129.160 ;
        RECT 135.315 128.280 135.605 128.325 ;
        RECT 132.080 128.140 135.605 128.280 ;
        RECT 132.080 128.080 132.400 128.140 ;
        RECT 135.315 128.095 135.605 128.140 ;
        RECT 13.330 127.460 138.910 127.940 ;
        RECT 69.060 127.260 69.380 127.320 ;
        RECT 71.375 127.260 71.665 127.305 ;
        RECT 69.060 127.120 71.665 127.260 ;
        RECT 69.060 127.060 69.380 127.120 ;
        RECT 71.375 127.075 71.665 127.120 ;
        RECT 75.975 127.260 76.265 127.305 ;
        RECT 78.720 127.260 79.040 127.320 ;
        RECT 75.975 127.120 79.040 127.260 ;
        RECT 75.975 127.075 76.265 127.120 ;
        RECT 78.720 127.060 79.040 127.120 ;
        RECT 80.560 127.260 80.880 127.320 ;
        RECT 81.495 127.260 81.785 127.305 ;
        RECT 80.560 127.120 81.785 127.260 ;
        RECT 80.560 127.060 80.880 127.120 ;
        RECT 81.495 127.075 81.785 127.120 ;
        RECT 102.640 127.060 102.960 127.320 ;
        RECT 115.520 127.260 115.840 127.320 ;
        RECT 129.795 127.260 130.085 127.305 ;
        RECT 115.520 127.120 130.085 127.260 ;
        RECT 115.520 127.060 115.840 127.120 ;
        RECT 129.795 127.075 130.085 127.120 ;
        RECT 136.680 127.060 137.000 127.320 ;
        RECT 64.000 126.580 64.320 126.640 ;
        RECT 57.190 126.440 64.320 126.580 ;
        RECT 78.810 126.580 78.950 127.060 ;
        RECT 83.795 126.920 84.085 126.965 ;
        RECT 96.240 126.920 96.530 126.965 ;
        RECT 98.340 126.920 98.630 126.965 ;
        RECT 99.910 126.920 100.200 126.965 ;
        RECT 83.795 126.780 87.690 126.920 ;
        RECT 83.795 126.735 84.085 126.780 ;
        RECT 87.550 126.625 87.690 126.780 ;
        RECT 96.240 126.780 100.200 126.920 ;
        RECT 96.240 126.735 96.530 126.780 ;
        RECT 98.340 126.735 98.630 126.780 ;
        RECT 99.910 126.735 100.200 126.780 ;
        RECT 112.800 126.920 113.090 126.965 ;
        RECT 114.900 126.920 115.190 126.965 ;
        RECT 116.470 126.920 116.760 126.965 ;
        RECT 112.800 126.780 116.760 126.920 ;
        RECT 112.800 126.735 113.090 126.780 ;
        RECT 114.900 126.735 115.190 126.780 ;
        RECT 116.470 126.735 116.760 126.780 ;
        RECT 119.200 126.720 119.520 126.980 ;
        RECT 78.810 126.440 81.250 126.580 ;
        RECT 23.060 126.240 23.380 126.300 ;
        RECT 25.835 126.240 26.125 126.285 ;
        RECT 27.215 126.240 27.505 126.285 ;
        RECT 23.060 126.100 27.505 126.240 ;
        RECT 23.060 126.040 23.380 126.100 ;
        RECT 25.835 126.055 26.125 126.100 ;
        RECT 27.215 126.055 27.505 126.100 ;
        RECT 31.340 126.240 31.660 126.300 ;
        RECT 57.190 126.285 57.330 126.440 ;
        RECT 64.000 126.380 64.320 126.440 ;
        RECT 31.340 126.100 39.850 126.240 ;
        RECT 31.340 126.040 31.660 126.100 ;
        RECT 39.710 125.560 39.850 126.100 ;
        RECT 56.195 126.055 56.485 126.285 ;
        RECT 57.115 126.055 57.405 126.285 ;
        RECT 59.875 126.240 60.165 126.285 ;
        RECT 62.620 126.240 62.940 126.300 ;
        RECT 59.875 126.100 62.940 126.240 ;
        RECT 59.875 126.055 60.165 126.100 ;
        RECT 56.270 125.900 56.410 126.055 ;
        RECT 62.620 126.040 62.940 126.100 ;
        RECT 74.580 126.040 74.900 126.300 ;
        RECT 76.420 126.240 76.740 126.300 ;
        RECT 78.275 126.240 78.565 126.285 ;
        RECT 76.420 126.100 78.565 126.240 ;
        RECT 76.420 126.040 76.740 126.100 ;
        RECT 78.275 126.055 78.565 126.100 ;
        RECT 79.195 126.240 79.485 126.285 ;
        RECT 80.560 126.240 80.880 126.300 ;
        RECT 81.110 126.285 81.250 126.440 ;
        RECT 87.475 126.395 87.765 126.625 ;
        RECT 96.635 126.580 96.925 126.625 ;
        RECT 97.825 126.580 98.115 126.625 ;
        RECT 100.345 126.580 100.635 126.625 ;
        RECT 96.635 126.440 100.635 126.580 ;
        RECT 96.635 126.395 96.925 126.440 ;
        RECT 97.825 126.395 98.115 126.440 ;
        RECT 100.345 126.395 100.635 126.440 ;
        RECT 106.780 126.380 107.100 126.640 ;
        RECT 112.300 126.380 112.620 126.640 ;
        RECT 113.195 126.580 113.485 126.625 ;
        RECT 114.385 126.580 114.675 126.625 ;
        RECT 116.905 126.580 117.195 126.625 ;
        RECT 131.620 126.580 131.940 126.640 ;
        RECT 113.195 126.440 117.195 126.580 ;
        RECT 113.195 126.395 113.485 126.440 ;
        RECT 114.385 126.395 114.675 126.440 ;
        RECT 116.905 126.395 117.195 126.440 ;
        RECT 130.790 126.440 131.940 126.580 ;
        RECT 79.195 126.100 80.880 126.240 ;
        RECT 79.195 126.055 79.485 126.100 ;
        RECT 63.080 125.900 63.400 125.960 ;
        RECT 56.270 125.760 63.400 125.900 ;
        RECT 63.080 125.700 63.400 125.760 ;
        RECT 69.980 125.900 70.300 125.960 ;
        RECT 75.815 125.900 76.105 125.945 ;
        RECT 69.980 125.760 76.105 125.900 ;
        RECT 69.980 125.700 70.300 125.760 ;
        RECT 75.815 125.715 76.105 125.760 ;
        RECT 56.180 125.560 56.500 125.620 ;
        RECT 39.710 125.420 56.500 125.560 ;
        RECT 56.180 125.360 56.500 125.420 ;
        RECT 56.655 125.560 56.945 125.605 ;
        RECT 57.560 125.560 57.880 125.620 ;
        RECT 56.655 125.420 57.880 125.560 ;
        RECT 56.655 125.375 56.945 125.420 ;
        RECT 57.560 125.360 57.880 125.420 ;
        RECT 75.040 125.360 75.360 125.620 ;
        RECT 76.510 125.560 76.650 126.040 ;
        RECT 76.895 125.900 77.185 125.945 ;
        RECT 79.270 125.900 79.410 126.055 ;
        RECT 80.560 126.040 80.880 126.100 ;
        RECT 81.035 126.055 81.325 126.285 ;
        RECT 82.415 126.055 82.705 126.285 ;
        RECT 82.490 125.900 82.630 126.055 ;
        RECT 95.740 126.040 96.060 126.300 ;
        RECT 97.120 126.285 97.440 126.300 ;
        RECT 97.090 126.240 97.440 126.285 ;
        RECT 96.925 126.100 97.440 126.240 ;
        RECT 97.090 126.055 97.440 126.100 ;
        RECT 97.120 126.040 97.440 126.055 ;
        RECT 99.880 126.240 100.200 126.300 ;
        RECT 101.720 126.240 102.040 126.300 ;
        RECT 99.880 126.100 108.850 126.240 ;
        RECT 99.880 126.040 100.200 126.100 ;
        RECT 101.720 126.040 102.040 126.100 ;
        RECT 76.895 125.760 79.410 125.900 ;
        RECT 79.730 125.760 82.630 125.900 ;
        RECT 83.780 125.900 84.100 125.960 ;
        RECT 86.080 125.900 86.400 125.960 ;
        RECT 86.555 125.900 86.845 125.945 ;
        RECT 83.780 125.760 86.845 125.900 ;
        RECT 76.895 125.715 77.185 125.760 ;
        RECT 79.730 125.560 79.870 125.760 ;
        RECT 83.780 125.700 84.100 125.760 ;
        RECT 86.080 125.700 86.400 125.760 ;
        RECT 86.555 125.715 86.845 125.760 ;
        RECT 95.280 125.900 95.600 125.960 ;
        RECT 105.875 125.900 106.165 125.945 ;
        RECT 108.175 125.900 108.465 125.945 ;
        RECT 95.280 125.760 104.710 125.900 ;
        RECT 95.280 125.700 95.600 125.760 ;
        RECT 76.510 125.420 79.870 125.560 ;
        RECT 80.115 125.560 80.405 125.605 ;
        RECT 81.020 125.560 81.340 125.620 ;
        RECT 80.115 125.420 81.340 125.560 ;
        RECT 80.115 125.375 80.405 125.420 ;
        RECT 81.020 125.360 81.340 125.420 ;
        RECT 84.700 125.360 85.020 125.620 ;
        RECT 87.015 125.560 87.305 125.605 ;
        RECT 90.220 125.560 90.540 125.620 ;
        RECT 87.015 125.420 90.540 125.560 ;
        RECT 87.015 125.375 87.305 125.420 ;
        RECT 90.220 125.360 90.540 125.420 ;
        RECT 104.020 125.360 104.340 125.620 ;
        RECT 104.570 125.560 104.710 125.760 ;
        RECT 105.875 125.760 108.465 125.900 ;
        RECT 108.710 125.900 108.850 126.100 ;
        RECT 110.920 126.040 111.240 126.300 ;
        RECT 112.760 126.240 113.080 126.300 ;
        RECT 113.595 126.240 113.885 126.285 ;
        RECT 112.760 126.100 113.885 126.240 ;
        RECT 112.760 126.040 113.080 126.100 ;
        RECT 113.595 126.055 113.885 126.100 ;
        RECT 127.940 126.240 128.260 126.300 ;
        RECT 130.790 126.285 130.930 126.440 ;
        RECT 131.620 126.380 131.940 126.440 ;
        RECT 130.715 126.240 131.005 126.285 ;
        RECT 127.940 126.100 131.005 126.240 ;
        RECT 127.940 126.040 128.260 126.100 ;
        RECT 130.715 126.055 131.005 126.100 ;
        RECT 131.175 126.240 131.465 126.285 ;
        RECT 132.080 126.240 132.400 126.300 ;
        RECT 131.175 126.100 132.400 126.240 ;
        RECT 131.175 126.055 131.465 126.100 ;
        RECT 132.080 126.040 132.400 126.100 ;
        RECT 132.555 126.240 132.845 126.285 ;
        RECT 133.460 126.240 133.780 126.300 ;
        RECT 132.555 126.100 133.780 126.240 ;
        RECT 132.555 126.055 132.845 126.100 ;
        RECT 133.460 126.040 133.780 126.100 ;
        RECT 133.935 126.055 134.225 126.285 ;
        RECT 120.120 125.900 120.440 125.960 ;
        RECT 127.480 125.900 127.800 125.960 ;
        RECT 108.710 125.760 127.800 125.900 ;
        RECT 105.875 125.715 106.165 125.760 ;
        RECT 108.175 125.715 108.465 125.760 ;
        RECT 120.120 125.700 120.440 125.760 ;
        RECT 127.480 125.700 127.800 125.760 ;
        RECT 129.780 125.900 130.100 125.960 ;
        RECT 131.635 125.900 131.925 125.945 ;
        RECT 129.780 125.760 131.925 125.900 ;
        RECT 129.780 125.700 130.100 125.760 ;
        RECT 131.635 125.715 131.925 125.760 ;
        RECT 106.335 125.560 106.625 125.605 ;
        RECT 114.140 125.560 114.460 125.620 ;
        RECT 104.570 125.420 114.460 125.560 ;
        RECT 106.335 125.375 106.625 125.420 ;
        RECT 114.140 125.360 114.460 125.420 ;
        RECT 125.180 125.560 125.500 125.620 ;
        RECT 134.010 125.560 134.150 126.055 ;
        RECT 135.760 126.040 136.080 126.300 ;
        RECT 125.180 125.420 134.150 125.560 ;
        RECT 125.180 125.360 125.500 125.420 ;
        RECT 134.840 125.360 135.160 125.620 ;
        RECT 13.330 124.740 138.910 125.220 ;
        RECT 105.875 124.355 106.165 124.585 ;
        RECT 118.295 124.540 118.585 124.585 ;
        RECT 119.660 124.540 119.980 124.600 ;
        RECT 118.295 124.400 119.980 124.540 ;
        RECT 118.295 124.355 118.585 124.400 ;
        RECT 16.620 124.200 16.940 124.260 ;
        RECT 24.295 124.200 24.585 124.245 ;
        RECT 16.620 124.060 24.585 124.200 ;
        RECT 16.620 124.000 16.940 124.060 ;
        RECT 24.295 124.015 24.585 124.060 ;
        RECT 25.375 124.015 25.665 124.245 ;
        RECT 66.730 124.200 67.020 124.245 ;
        RECT 68.600 124.200 68.920 124.260 ;
        RECT 57.650 124.060 62.850 124.200 ;
        RECT 20.760 123.520 21.080 123.580 ;
        RECT 25.450 123.520 25.590 124.015 ;
        RECT 57.650 123.905 57.790 124.060 ;
        RECT 62.710 123.920 62.850 124.060 ;
        RECT 66.730 124.060 68.920 124.200 ;
        RECT 66.730 124.015 67.020 124.060 ;
        RECT 68.600 124.000 68.920 124.060 ;
        RECT 80.115 124.200 80.405 124.245 ;
        RECT 83.320 124.200 83.640 124.260 ;
        RECT 80.115 124.060 83.640 124.200 ;
        RECT 80.115 124.015 80.405 124.060 ;
        RECT 83.320 124.000 83.640 124.060 ;
        RECT 84.210 124.200 84.500 124.245 ;
        RECT 84.700 124.200 85.020 124.260 ;
        RECT 84.210 124.060 85.020 124.200 ;
        RECT 84.210 124.015 84.500 124.060 ;
        RECT 84.700 124.000 85.020 124.060 ;
        RECT 89.760 124.200 90.080 124.260 ;
        RECT 97.090 124.200 97.380 124.245 ;
        RECT 104.020 124.200 104.340 124.260 ;
        RECT 89.760 124.060 94.130 124.200 ;
        RECT 89.760 124.000 90.080 124.060 ;
        RECT 58.940 123.905 59.260 123.920 ;
        RECT 28.135 123.675 28.425 123.905 ;
        RECT 57.575 123.675 57.865 123.905 ;
        RECT 58.910 123.860 59.260 123.905 ;
        RECT 58.745 123.720 59.260 123.860 ;
        RECT 58.910 123.675 59.260 123.720 ;
        RECT 20.760 123.380 25.590 123.520 ;
        RECT 20.760 123.320 21.080 123.380 ;
        RECT 22.600 123.180 22.920 123.240 ;
        RECT 28.210 123.180 28.350 123.675 ;
        RECT 58.940 123.660 59.260 123.675 ;
        RECT 62.620 123.860 62.940 123.920 ;
        RECT 65.395 123.860 65.685 123.905 ;
        RECT 62.620 123.720 65.685 123.860 ;
        RECT 62.620 123.660 62.940 123.720 ;
        RECT 65.395 123.675 65.685 123.720 ;
        RECT 81.480 123.860 81.800 123.920 ;
        RECT 82.875 123.860 83.165 123.905 ;
        RECT 81.480 123.720 83.165 123.860 ;
        RECT 83.410 123.860 83.550 124.000 ;
        RECT 92.995 123.860 93.285 123.905 ;
        RECT 83.410 123.720 93.285 123.860 ;
        RECT 81.480 123.660 81.800 123.720 ;
        RECT 82.875 123.675 83.165 123.720 ;
        RECT 92.995 123.675 93.285 123.720 ;
        RECT 54.355 123.520 54.645 123.565 ;
        RECT 55.720 123.520 56.040 123.580 ;
        RECT 54.355 123.380 56.040 123.520 ;
        RECT 54.355 123.335 54.645 123.380 ;
        RECT 55.720 123.320 56.040 123.380 ;
        RECT 58.455 123.520 58.745 123.565 ;
        RECT 59.645 123.520 59.935 123.565 ;
        RECT 62.165 123.520 62.455 123.565 ;
        RECT 58.455 123.380 62.455 123.520 ;
        RECT 58.455 123.335 58.745 123.380 ;
        RECT 59.645 123.335 59.935 123.380 ;
        RECT 62.165 123.335 62.455 123.380 ;
        RECT 66.275 123.520 66.565 123.565 ;
        RECT 67.465 123.520 67.755 123.565 ;
        RECT 69.985 123.520 70.275 123.565 ;
        RECT 72.755 123.520 73.045 123.565 ;
        RECT 66.275 123.380 70.275 123.520 ;
        RECT 66.275 123.335 66.565 123.380 ;
        RECT 67.465 123.335 67.755 123.380 ;
        RECT 69.985 123.335 70.275 123.380 ;
        RECT 72.370 123.380 73.045 123.520 ;
        RECT 32.260 123.180 32.580 123.240 ;
        RECT 22.600 123.040 32.580 123.180 ;
        RECT 22.600 122.980 22.920 123.040 ;
        RECT 32.260 122.980 32.580 123.040 ;
        RECT 58.060 123.180 58.350 123.225 ;
        RECT 60.160 123.180 60.450 123.225 ;
        RECT 61.730 123.180 62.020 123.225 ;
        RECT 58.060 123.040 62.020 123.180 ;
        RECT 58.060 122.995 58.350 123.040 ;
        RECT 60.160 122.995 60.450 123.040 ;
        RECT 61.730 122.995 62.020 123.040 ;
        RECT 65.880 123.180 66.170 123.225 ;
        RECT 67.980 123.180 68.270 123.225 ;
        RECT 69.550 123.180 69.840 123.225 ;
        RECT 65.880 123.040 69.840 123.180 ;
        RECT 65.880 122.995 66.170 123.040 ;
        RECT 67.980 122.995 68.270 123.040 ;
        RECT 69.550 122.995 69.840 123.040 ;
        RECT 72.370 122.900 72.510 123.380 ;
        RECT 72.755 123.335 73.045 123.380 ;
        RECT 80.560 123.320 80.880 123.580 ;
        RECT 81.020 123.320 81.340 123.580 ;
        RECT 83.755 123.520 84.045 123.565 ;
        RECT 84.945 123.520 85.235 123.565 ;
        RECT 87.465 123.520 87.755 123.565 ;
        RECT 90.220 123.520 90.540 123.580 ;
        RECT 93.990 123.565 94.130 124.060 ;
        RECT 97.090 124.060 104.340 124.200 ;
        RECT 105.950 124.200 106.090 124.355 ;
        RECT 119.660 124.340 119.980 124.400 ;
        RECT 108.160 124.200 108.480 124.260 ;
        RECT 105.950 124.060 108.480 124.200 ;
        RECT 97.090 124.015 97.380 124.060 ;
        RECT 104.020 124.000 104.340 124.060 ;
        RECT 108.160 124.000 108.480 124.060 ;
        RECT 102.640 123.860 102.960 123.920 ;
        RECT 104.495 123.860 104.785 123.905 ;
        RECT 102.640 123.720 104.785 123.860 ;
        RECT 102.640 123.660 102.960 123.720 ;
        RECT 104.495 123.675 104.785 123.720 ;
        RECT 106.335 123.860 106.625 123.905 ;
        RECT 108.620 123.860 108.940 123.920 ;
        RECT 106.335 123.720 108.940 123.860 ;
        RECT 106.335 123.675 106.625 123.720 ;
        RECT 108.620 123.660 108.940 123.720 ;
        RECT 117.360 123.660 117.680 123.920 ;
        RECT 119.750 123.860 119.890 124.340 ;
        RECT 126.575 124.200 126.865 124.245 ;
        RECT 128.260 124.200 128.550 124.245 ;
        RECT 126.575 124.060 128.550 124.200 ;
        RECT 126.575 124.015 126.865 124.060 ;
        RECT 128.260 124.015 128.550 124.060 ;
        RECT 123.355 123.860 123.645 123.905 ;
        RECT 119.750 123.720 123.645 123.860 ;
        RECT 123.355 123.675 123.645 123.720 ;
        RECT 124.260 123.660 124.580 123.920 ;
        RECT 124.735 123.675 125.025 123.905 ;
        RECT 125.195 123.860 125.485 123.905 ;
        RECT 126.100 123.860 126.420 123.920 ;
        RECT 125.195 123.720 126.420 123.860 ;
        RECT 125.195 123.675 125.485 123.720 ;
        RECT 83.755 123.380 87.755 123.520 ;
        RECT 83.755 123.335 84.045 123.380 ;
        RECT 84.945 123.335 85.235 123.380 ;
        RECT 87.465 123.335 87.755 123.380 ;
        RECT 89.850 123.380 90.540 123.520 ;
        RECT 89.850 123.225 89.990 123.380 ;
        RECT 90.220 123.320 90.540 123.380 ;
        RECT 93.455 123.335 93.745 123.565 ;
        RECT 93.915 123.335 94.205 123.565 ;
        RECT 83.360 123.180 83.650 123.225 ;
        RECT 85.460 123.180 85.750 123.225 ;
        RECT 87.030 123.180 87.320 123.225 ;
        RECT 83.360 123.040 87.320 123.180 ;
        RECT 83.360 122.995 83.650 123.040 ;
        RECT 85.460 122.995 85.750 123.040 ;
        RECT 87.030 122.995 87.320 123.040 ;
        RECT 89.775 122.995 90.065 123.225 ;
        RECT 90.680 123.180 91.000 123.240 ;
        RECT 93.530 123.180 93.670 123.335 ;
        RECT 95.740 123.320 96.060 123.580 ;
        RECT 96.635 123.520 96.925 123.565 ;
        RECT 97.825 123.520 98.115 123.565 ;
        RECT 100.345 123.520 100.635 123.565 ;
        RECT 96.635 123.380 100.635 123.520 ;
        RECT 96.635 123.335 96.925 123.380 ;
        RECT 97.825 123.335 98.115 123.380 ;
        RECT 100.345 123.335 100.635 123.380 ;
        RECT 104.035 123.520 104.325 123.565 ;
        RECT 110.920 123.520 111.240 123.580 ;
        RECT 104.035 123.380 111.240 123.520 ;
        RECT 104.035 123.335 104.325 123.380 ;
        RECT 96.240 123.180 96.530 123.225 ;
        RECT 98.340 123.180 98.630 123.225 ;
        RECT 99.910 123.180 100.200 123.225 ;
        RECT 90.680 123.040 94.130 123.180 ;
        RECT 90.680 122.980 91.000 123.040 ;
        RECT 21.680 122.840 22.000 122.900 ;
        RECT 23.535 122.840 23.825 122.885 ;
        RECT 21.680 122.700 23.825 122.840 ;
        RECT 21.680 122.640 22.000 122.700 ;
        RECT 23.535 122.655 23.825 122.700 ;
        RECT 24.440 122.640 24.760 122.900 ;
        RECT 24.900 122.840 25.220 122.900 ;
        RECT 31.800 122.840 32.120 122.900 ;
        RECT 40.540 122.840 40.860 122.900 ;
        RECT 24.900 122.700 40.860 122.840 ;
        RECT 24.900 122.640 25.220 122.700 ;
        RECT 31.800 122.640 32.120 122.700 ;
        RECT 40.540 122.640 40.860 122.700 ;
        RECT 57.115 122.840 57.405 122.885 ;
        RECT 63.080 122.840 63.400 122.900 ;
        RECT 57.115 122.700 63.400 122.840 ;
        RECT 57.115 122.655 57.405 122.700 ;
        RECT 63.080 122.640 63.400 122.700 ;
        RECT 64.475 122.840 64.765 122.885 ;
        RECT 68.600 122.840 68.920 122.900 ;
        RECT 64.475 122.700 68.920 122.840 ;
        RECT 64.475 122.655 64.765 122.700 ;
        RECT 68.600 122.640 68.920 122.700 ;
        RECT 72.280 122.640 72.600 122.900 ;
        RECT 75.975 122.840 76.265 122.885 ;
        RECT 76.420 122.840 76.740 122.900 ;
        RECT 75.975 122.700 76.740 122.840 ;
        RECT 75.975 122.655 76.265 122.700 ;
        RECT 76.420 122.640 76.740 122.700 ;
        RECT 78.260 122.640 78.580 122.900 ;
        RECT 90.220 122.840 90.540 122.900 ;
        RECT 91.155 122.840 91.445 122.885 ;
        RECT 90.220 122.700 91.445 122.840 ;
        RECT 93.990 122.840 94.130 123.040 ;
        RECT 96.240 123.040 100.200 123.180 ;
        RECT 96.240 122.995 96.530 123.040 ;
        RECT 98.340 122.995 98.630 123.040 ;
        RECT 99.910 122.995 100.200 123.040 ;
        RECT 102.655 123.180 102.945 123.225 ;
        RECT 104.110 123.180 104.250 123.335 ;
        RECT 110.920 123.320 111.240 123.380 ;
        RECT 117.820 123.520 118.140 123.580 ;
        RECT 124.810 123.520 124.950 123.675 ;
        RECT 126.100 123.660 126.420 123.720 ;
        RECT 127.020 123.660 127.340 123.920 ;
        RECT 117.820 123.380 124.950 123.520 ;
        RECT 127.915 123.520 128.205 123.565 ;
        RECT 129.105 123.520 129.395 123.565 ;
        RECT 131.625 123.520 131.915 123.565 ;
        RECT 127.915 123.380 131.915 123.520 ;
        RECT 117.820 123.320 118.140 123.380 ;
        RECT 127.915 123.335 128.205 123.380 ;
        RECT 129.105 123.335 129.395 123.380 ;
        RECT 131.625 123.335 131.915 123.380 ;
        RECT 104.480 123.180 104.800 123.240 ;
        RECT 102.655 123.040 104.800 123.180 ;
        RECT 102.655 122.995 102.945 123.040 ;
        RECT 104.480 122.980 104.800 123.040 ;
        RECT 127.520 123.180 127.810 123.225 ;
        RECT 129.620 123.180 129.910 123.225 ;
        RECT 131.190 123.180 131.480 123.225 ;
        RECT 127.520 123.040 131.480 123.180 ;
        RECT 127.520 122.995 127.810 123.040 ;
        RECT 129.620 122.995 129.910 123.040 ;
        RECT 131.190 122.995 131.480 123.040 ;
        RECT 96.660 122.840 96.980 122.900 ;
        RECT 107.700 122.840 108.020 122.900 ;
        RECT 93.990 122.700 108.020 122.840 ;
        RECT 90.220 122.640 90.540 122.700 ;
        RECT 91.155 122.655 91.445 122.700 ;
        RECT 96.660 122.640 96.980 122.700 ;
        RECT 107.700 122.640 108.020 122.700 ;
        RECT 110.000 122.840 110.320 122.900 ;
        RECT 111.840 122.840 112.160 122.900 ;
        RECT 110.000 122.700 112.160 122.840 ;
        RECT 110.000 122.640 110.320 122.700 ;
        RECT 111.840 122.640 112.160 122.700 ;
        RECT 133.920 122.640 134.240 122.900 ;
        RECT 13.330 122.020 138.910 122.500 ;
        RECT 16.175 121.820 16.465 121.865 ;
        RECT 17.540 121.820 17.860 121.880 ;
        RECT 25.360 121.820 25.680 121.880 ;
        RECT 35.020 121.820 35.340 121.880 ;
        RECT 40.080 121.820 40.400 121.880 ;
        RECT 57.560 121.820 57.880 121.880 ;
        RECT 72.280 121.820 72.600 121.880 ;
        RECT 74.135 121.820 74.425 121.865 ;
        RECT 16.175 121.680 34.790 121.820 ;
        RECT 16.175 121.635 16.465 121.680 ;
        RECT 17.540 121.620 17.860 121.680 ;
        RECT 18.920 121.480 19.210 121.525 ;
        RECT 20.490 121.480 20.780 121.525 ;
        RECT 22.590 121.480 22.880 121.525 ;
        RECT 18.920 121.340 22.880 121.480 ;
        RECT 18.920 121.295 19.210 121.340 ;
        RECT 20.490 121.295 20.780 121.340 ;
        RECT 22.590 121.295 22.880 121.340 ;
        RECT 18.485 121.140 18.775 121.185 ;
        RECT 21.005 121.140 21.295 121.185 ;
        RECT 22.195 121.140 22.485 121.185 ;
        RECT 18.485 121.000 22.485 121.140 ;
        RECT 18.485 120.955 18.775 121.000 ;
        RECT 21.005 120.955 21.295 121.000 ;
        RECT 22.195 120.955 22.485 121.000 ;
        RECT 21.680 120.845 22.000 120.860 ;
        RECT 21.680 120.800 22.030 120.845 ;
        RECT 22.600 120.800 22.920 120.860 ;
        RECT 23.610 120.845 23.750 121.680 ;
        RECT 25.360 121.620 25.680 121.680 ;
        RECT 25.820 121.480 26.140 121.540 ;
        RECT 25.820 121.340 34.330 121.480 ;
        RECT 25.820 121.280 26.140 121.340 ;
        RECT 23.075 120.800 23.365 120.845 ;
        RECT 21.680 120.660 22.195 120.800 ;
        RECT 22.600 120.660 23.365 120.800 ;
        RECT 21.680 120.615 22.030 120.660 ;
        RECT 21.680 120.600 22.000 120.615 ;
        RECT 22.600 120.600 22.920 120.660 ;
        RECT 23.075 120.615 23.365 120.660 ;
        RECT 23.535 120.615 23.825 120.845 ;
        RECT 24.915 120.615 25.205 120.845 ;
        RECT 28.135 120.800 28.425 120.845 ;
        RECT 31.340 120.800 31.660 120.860 ;
        RECT 34.190 120.845 34.330 121.340 ;
        RECT 34.650 121.140 34.790 121.680 ;
        RECT 35.020 121.680 40.400 121.820 ;
        RECT 35.020 121.620 35.340 121.680 ;
        RECT 40.080 121.620 40.400 121.680 ;
        RECT 52.590 121.680 57.880 121.820 ;
        RECT 37.320 121.280 37.640 121.540 ;
        RECT 37.795 121.295 38.085 121.525 ;
        RECT 38.700 121.480 39.020 121.540 ;
        RECT 41.015 121.480 41.305 121.525 ;
        RECT 38.700 121.340 41.305 121.480 ;
        RECT 37.410 121.140 37.550 121.280 ;
        RECT 34.650 121.000 37.550 121.140 ;
        RECT 37.870 121.140 38.010 121.295 ;
        RECT 38.700 121.280 39.020 121.340 ;
        RECT 41.015 121.295 41.305 121.340 ;
        RECT 43.760 121.480 44.080 121.540 ;
        RECT 47.440 121.480 47.760 121.540 ;
        RECT 43.760 121.340 47.760 121.480 ;
        RECT 43.760 121.280 44.080 121.340 ;
        RECT 47.440 121.280 47.760 121.340 ;
        RECT 40.540 121.140 40.860 121.200 ;
        RECT 41.475 121.140 41.765 121.185 ;
        RECT 37.870 121.000 42.615 121.140 ;
        RECT 34.650 120.845 34.790 121.000 ;
        RECT 40.540 120.940 40.860 121.000 ;
        RECT 41.475 120.955 41.765 121.000 ;
        RECT 28.135 120.660 31.660 120.800 ;
        RECT 28.135 120.615 28.425 120.660 ;
        RECT 24.990 120.460 25.130 120.615 ;
        RECT 31.340 120.600 31.660 120.660 ;
        RECT 34.115 120.615 34.405 120.845 ;
        RECT 34.575 120.615 34.865 120.845 ;
        RECT 35.020 120.600 35.340 120.860 ;
        RECT 36.400 120.800 36.720 120.860 ;
        RECT 36.400 120.660 39.850 120.800 ;
        RECT 36.400 120.600 36.720 120.660 ;
        RECT 30.880 120.460 31.200 120.520 ;
        RECT 24.990 120.320 31.200 120.460 ;
        RECT 30.880 120.260 31.200 120.320 ;
        RECT 32.260 120.260 32.580 120.520 ;
        RECT 33.195 120.460 33.485 120.505 ;
        RECT 35.480 120.460 35.800 120.520 ;
        RECT 33.195 120.320 35.800 120.460 ;
        RECT 33.195 120.275 33.485 120.320 ;
        RECT 35.480 120.260 35.800 120.320 ;
        RECT 35.940 120.260 36.260 120.520 ;
        RECT 37.320 120.460 37.640 120.520 ;
        RECT 39.175 120.460 39.465 120.505 ;
        RECT 37.320 120.320 39.465 120.460 ;
        RECT 39.710 120.460 39.850 120.660 ;
        RECT 40.080 120.600 40.400 120.860 ;
        RECT 41.920 120.800 42.240 120.860 ;
        RECT 42.475 120.845 42.615 121.000 ;
        RECT 52.590 120.845 52.730 121.680 ;
        RECT 57.560 121.620 57.880 121.680 ;
        RECT 69.840 121.680 74.425 121.820 ;
        RECT 53.895 121.295 54.185 121.525 ;
        RECT 54.840 121.480 55.130 121.525 ;
        RECT 56.940 121.480 57.230 121.525 ;
        RECT 58.510 121.480 58.800 121.525 ;
        RECT 54.840 121.340 58.800 121.480 ;
        RECT 54.840 121.295 55.130 121.340 ;
        RECT 56.940 121.295 57.230 121.340 ;
        RECT 58.510 121.295 58.800 121.340 ;
        RECT 53.970 121.140 54.110 121.295 ;
        RECT 55.235 121.140 55.525 121.185 ;
        RECT 56.425 121.140 56.715 121.185 ;
        RECT 58.945 121.140 59.235 121.185 ;
        RECT 53.970 121.000 55.030 121.140 ;
        RECT 40.630 120.660 42.240 120.800 ;
        RECT 40.630 120.460 40.770 120.660 ;
        RECT 41.920 120.600 42.240 120.660 ;
        RECT 42.400 120.615 42.690 120.845 ;
        RECT 52.515 120.615 52.805 120.845 ;
        RECT 54.340 120.600 54.660 120.860 ;
        RECT 39.710 120.320 40.770 120.460 ;
        RECT 53.895 120.460 54.185 120.505 ;
        RECT 54.890 120.460 55.030 121.000 ;
        RECT 55.235 121.000 59.235 121.140 ;
        RECT 55.235 120.955 55.525 121.000 ;
        RECT 56.425 120.955 56.715 121.000 ;
        RECT 58.945 120.955 59.235 121.000 ;
        RECT 68.600 120.940 68.920 121.200 ;
        RECT 69.200 121.140 69.490 121.185 ;
        RECT 69.840 121.140 69.980 121.680 ;
        RECT 72.280 121.620 72.600 121.680 ;
        RECT 74.135 121.635 74.425 121.680 ;
        RECT 75.960 121.620 76.280 121.880 ;
        RECT 90.680 121.620 91.000 121.880 ;
        RECT 102.640 121.820 102.960 121.880 ;
        RECT 104.955 121.820 105.245 121.865 ;
        RECT 120.595 121.820 120.885 121.865 ;
        RECT 102.640 121.680 105.245 121.820 ;
        RECT 102.640 121.620 102.960 121.680 ;
        RECT 104.955 121.635 105.245 121.680 ;
        RECT 111.930 121.680 120.885 121.820 ;
        RECT 84.280 121.480 84.570 121.525 ;
        RECT 86.380 121.480 86.670 121.525 ;
        RECT 87.950 121.480 88.240 121.525 ;
        RECT 84.280 121.340 88.240 121.480 ;
        RECT 84.280 121.295 84.570 121.340 ;
        RECT 86.380 121.295 86.670 121.340 ;
        RECT 87.950 121.295 88.240 121.340 ;
        RECT 69.200 121.000 69.980 121.140 ;
        RECT 73.675 121.140 73.965 121.185 ;
        RECT 81.480 121.140 81.800 121.200 ;
        RECT 83.795 121.140 84.085 121.185 ;
        RECT 73.675 121.000 79.410 121.140 ;
        RECT 69.200 120.955 69.490 121.000 ;
        RECT 73.675 120.955 73.965 121.000 ;
        RECT 65.380 120.800 65.700 120.860 ;
        RECT 66.775 120.800 67.065 120.845 ;
        RECT 65.380 120.660 67.065 120.800 ;
        RECT 68.690 120.800 68.830 120.940 ;
        RECT 73.750 120.800 73.890 120.955 ;
        RECT 68.690 120.660 73.890 120.800 ;
        RECT 65.380 120.600 65.700 120.660 ;
        RECT 66.775 120.615 67.065 120.660 ;
        RECT 74.135 120.615 74.425 120.845 ;
        RECT 75.055 120.800 75.345 120.845 ;
        RECT 75.960 120.800 76.280 120.860 ;
        RECT 75.055 120.660 76.280 120.800 ;
        RECT 75.055 120.615 75.345 120.660 ;
        RECT 55.580 120.460 55.870 120.505 ;
        RECT 53.895 120.320 54.570 120.460 ;
        RECT 54.890 120.320 55.870 120.460 ;
        RECT 37.320 120.260 37.640 120.320 ;
        RECT 39.175 120.275 39.465 120.320 ;
        RECT 53.895 120.275 54.185 120.320 ;
        RECT 23.995 120.120 24.285 120.165 ;
        RECT 24.900 120.120 25.220 120.180 ;
        RECT 23.995 119.980 25.220 120.120 ;
        RECT 23.995 119.935 24.285 119.980 ;
        RECT 24.900 119.920 25.220 119.980 ;
        RECT 25.835 120.120 26.125 120.165 ;
        RECT 31.340 120.120 31.660 120.180 ;
        RECT 25.835 119.980 31.660 120.120 ;
        RECT 25.835 119.935 26.125 119.980 ;
        RECT 31.340 119.920 31.660 119.980 ;
        RECT 36.400 120.120 36.720 120.180 ;
        RECT 38.715 120.120 39.005 120.165 ;
        RECT 41.460 120.120 41.780 120.180 ;
        RECT 36.400 119.980 41.780 120.120 ;
        RECT 36.400 119.920 36.720 119.980 ;
        RECT 38.715 119.935 39.005 119.980 ;
        RECT 41.460 119.920 41.780 119.980 ;
        RECT 52.960 119.920 53.280 120.180 ;
        RECT 54.430 120.120 54.570 120.320 ;
        RECT 55.580 120.275 55.870 120.320 ;
        RECT 60.320 120.460 60.640 120.520 ;
        RECT 61.715 120.460 62.005 120.505 ;
        RECT 60.320 120.320 62.005 120.460 ;
        RECT 60.320 120.260 60.640 120.320 ;
        RECT 61.715 120.275 62.005 120.320 ;
        RECT 68.155 120.460 68.445 120.505 ;
        RECT 74.210 120.460 74.350 120.615 ;
        RECT 75.960 120.600 76.280 120.660 ;
        RECT 76.880 120.800 77.200 120.860 ;
        RECT 79.270 120.845 79.410 121.000 ;
        RECT 81.480 121.000 84.085 121.140 ;
        RECT 81.480 120.940 81.800 121.000 ;
        RECT 83.795 120.955 84.085 121.000 ;
        RECT 84.675 121.140 84.965 121.185 ;
        RECT 85.865 121.140 86.155 121.185 ;
        RECT 88.385 121.140 88.675 121.185 ;
        RECT 84.675 121.000 88.675 121.140 ;
        RECT 84.675 120.955 84.965 121.000 ;
        RECT 85.865 120.955 86.155 121.000 ;
        RECT 88.385 120.955 88.675 121.000 ;
        RECT 96.200 121.140 96.520 121.200 ;
        RECT 105.860 121.140 106.180 121.200 ;
        RECT 110.460 121.140 110.780 121.200 ;
        RECT 96.200 121.000 110.780 121.140 ;
        RECT 96.200 120.940 96.520 121.000 ;
        RECT 105.860 120.940 106.180 121.000 ;
        RECT 110.460 120.940 110.780 121.000 ;
        RECT 78.275 120.800 78.565 120.845 ;
        RECT 76.880 120.660 78.565 120.800 ;
        RECT 76.880 120.600 77.200 120.660 ;
        RECT 78.275 120.615 78.565 120.660 ;
        RECT 79.195 120.615 79.485 120.845 ;
        RECT 85.130 120.800 85.420 120.845 ;
        RECT 90.220 120.800 90.540 120.860 ;
        RECT 85.130 120.660 90.540 120.800 ;
        RECT 85.130 120.615 85.420 120.660 ;
        RECT 90.220 120.600 90.540 120.660 ;
        RECT 102.655 120.800 102.945 120.845 ;
        RECT 104.480 120.800 104.800 120.860 ;
        RECT 110.000 120.800 110.320 120.860 ;
        RECT 110.935 120.800 111.225 120.845 ;
        RECT 102.655 120.660 105.170 120.800 ;
        RECT 102.655 120.615 102.945 120.660 ;
        RECT 104.480 120.600 104.800 120.660 ;
        RECT 75.500 120.460 75.820 120.520 ;
        RECT 78.735 120.460 79.025 120.505 ;
        RECT 68.155 120.320 72.510 120.460 ;
        RECT 74.210 120.320 79.025 120.460 ;
        RECT 68.155 120.275 68.445 120.320 ;
        RECT 58.940 120.120 59.260 120.180 ;
        RECT 54.430 119.980 59.260 120.120 ;
        RECT 58.940 119.920 59.260 119.980 ;
        RECT 61.255 120.120 61.545 120.165 ;
        RECT 64.000 120.120 64.320 120.180 ;
        RECT 61.255 119.980 64.320 120.120 ;
        RECT 61.255 119.935 61.545 119.980 ;
        RECT 64.000 119.920 64.320 119.980 ;
        RECT 64.460 120.120 64.780 120.180 ;
        RECT 69.520 120.120 69.840 120.180 ;
        RECT 64.460 119.980 69.840 120.120 ;
        RECT 64.460 119.920 64.780 119.980 ;
        RECT 69.520 119.920 69.840 119.980 ;
        RECT 69.980 119.920 70.300 120.180 ;
        RECT 70.440 119.920 70.760 120.180 ;
        RECT 72.370 120.120 72.510 120.320 ;
        RECT 75.500 120.260 75.820 120.320 ;
        RECT 78.735 120.275 79.025 120.320 ;
        RECT 101.260 120.460 101.580 120.520 ;
        RECT 105.030 120.505 105.170 120.660 ;
        RECT 110.000 120.660 111.225 120.800 ;
        RECT 110.000 120.600 110.320 120.660 ;
        RECT 110.935 120.615 111.225 120.660 ;
        RECT 111.380 120.600 111.700 120.860 ;
        RECT 111.930 120.845 112.070 121.680 ;
        RECT 120.595 121.635 120.885 121.680 ;
        RECT 124.260 121.820 124.580 121.880 ;
        RECT 131.635 121.820 131.925 121.865 ;
        RECT 124.260 121.680 131.925 121.820 ;
        RECT 124.260 121.620 124.580 121.680 ;
        RECT 131.635 121.635 131.925 121.680 ;
        RECT 113.720 121.480 114.010 121.525 ;
        RECT 115.820 121.480 116.110 121.525 ;
        RECT 117.390 121.480 117.680 121.525 ;
        RECT 113.720 121.340 117.680 121.480 ;
        RECT 113.720 121.295 114.010 121.340 ;
        RECT 115.820 121.295 116.110 121.340 ;
        RECT 117.390 121.295 117.680 121.340 ;
        RECT 118.280 121.480 118.600 121.540 ;
        RECT 120.135 121.480 120.425 121.525 ;
        RECT 121.960 121.480 122.280 121.540 ;
        RECT 129.780 121.480 130.100 121.540 ;
        RECT 118.280 121.340 121.730 121.480 ;
        RECT 118.280 121.280 118.600 121.340 ;
        RECT 120.135 121.295 120.425 121.340 ;
        RECT 112.300 121.140 112.620 121.200 ;
        RECT 113.235 121.140 113.525 121.185 ;
        RECT 112.300 121.000 113.525 121.140 ;
        RECT 112.300 120.940 112.620 121.000 ;
        RECT 113.235 120.955 113.525 121.000 ;
        RECT 114.115 121.140 114.405 121.185 ;
        RECT 115.305 121.140 115.595 121.185 ;
        RECT 117.825 121.140 118.115 121.185 ;
        RECT 114.115 121.000 118.115 121.140 ;
        RECT 114.115 120.955 114.405 121.000 ;
        RECT 115.305 120.955 115.595 121.000 ;
        RECT 117.825 120.955 118.115 121.000 ;
        RECT 111.855 120.615 112.145 120.845 ;
        RECT 112.775 120.800 113.065 120.845 ;
        RECT 119.660 120.800 119.980 120.860 ;
        RECT 121.590 120.845 121.730 121.340 ;
        RECT 121.960 121.340 130.100 121.480 ;
        RECT 121.960 121.280 122.280 121.340 ;
        RECT 129.780 121.280 130.100 121.340 ;
        RECT 124.720 121.140 125.040 121.200 ;
        RECT 133.920 121.140 134.240 121.200 ;
        RECT 124.720 121.000 129.505 121.140 ;
        RECT 124.720 120.940 125.040 121.000 ;
        RECT 112.775 120.660 119.980 120.800 ;
        RECT 112.775 120.615 113.065 120.660 ;
        RECT 119.660 120.600 119.980 120.660 ;
        RECT 121.515 120.800 121.805 120.845 ;
        RECT 125.180 120.800 125.500 120.860 ;
        RECT 121.515 120.660 125.500 120.800 ;
        RECT 129.365 120.800 129.505 121.000 ;
        RECT 130.790 121.000 134.240 121.140 ;
        RECT 130.790 120.845 130.930 121.000 ;
        RECT 133.920 120.940 134.240 121.000 ;
        RECT 129.795 120.800 130.085 120.845 ;
        RECT 129.365 120.660 130.085 120.800 ;
        RECT 121.515 120.615 121.805 120.660 ;
        RECT 125.180 120.600 125.500 120.660 ;
        RECT 129.795 120.615 130.085 120.660 ;
        RECT 130.715 120.615 131.005 120.845 ;
        RECT 131.250 120.660 134.150 120.800 ;
        RECT 104.035 120.460 104.325 120.505 ;
        RECT 101.260 120.320 104.325 120.460 ;
        RECT 101.260 120.260 101.580 120.320 ;
        RECT 104.035 120.275 104.325 120.320 ;
        RECT 104.955 120.275 105.245 120.505 ;
        RECT 109.555 120.460 109.845 120.505 ;
        RECT 114.460 120.460 114.750 120.505 ;
        RECT 109.555 120.320 114.750 120.460 ;
        RECT 109.555 120.275 109.845 120.320 ;
        RECT 114.460 120.275 114.750 120.320 ;
        RECT 122.420 120.260 122.740 120.520 ;
        RECT 131.250 120.460 131.390 120.660 ;
        RECT 126.190 120.320 131.390 120.460 ;
        RECT 74.120 120.120 74.440 120.180 ;
        RECT 72.370 119.980 74.440 120.120 ;
        RECT 74.120 119.920 74.440 119.980 ;
        RECT 102.195 120.120 102.485 120.165 ;
        RECT 103.100 120.120 103.420 120.180 ;
        RECT 102.195 119.980 103.420 120.120 ;
        RECT 102.195 119.935 102.485 119.980 ;
        RECT 103.100 119.920 103.420 119.980 ;
        RECT 105.875 120.120 106.165 120.165 ;
        RECT 115.520 120.120 115.840 120.180 ;
        RECT 105.875 119.980 115.840 120.120 ;
        RECT 122.510 120.120 122.650 120.260 ;
        RECT 126.190 120.120 126.330 120.320 ;
        RECT 133.000 120.260 133.320 120.520 ;
        RECT 134.010 120.505 134.150 120.660 ;
        RECT 135.760 120.600 136.080 120.860 ;
        RECT 133.935 120.460 134.225 120.505 ;
        RECT 134.380 120.460 134.700 120.520 ;
        RECT 133.935 120.320 134.700 120.460 ;
        RECT 133.935 120.275 134.225 120.320 ;
        RECT 134.380 120.260 134.700 120.320 ;
        RECT 122.510 119.980 126.330 120.120 ;
        RECT 130.240 120.120 130.560 120.180 ;
        RECT 132.095 120.120 132.385 120.165 ;
        RECT 130.240 119.980 132.385 120.120 ;
        RECT 105.875 119.935 106.165 119.980 ;
        RECT 115.520 119.920 115.840 119.980 ;
        RECT 130.240 119.920 130.560 119.980 ;
        RECT 132.095 119.935 132.385 119.980 ;
        RECT 136.680 119.920 137.000 120.180 ;
        RECT 13.330 119.300 138.910 119.780 ;
        RECT 16.620 118.900 16.940 119.160 ;
        RECT 20.760 118.900 21.080 119.160 ;
        RECT 21.695 119.100 21.985 119.145 ;
        RECT 31.355 119.100 31.645 119.145 ;
        RECT 36.860 119.100 37.180 119.160 ;
        RECT 21.695 118.960 23.750 119.100 ;
        RECT 21.695 118.915 21.985 118.960 ;
        RECT 17.540 118.560 17.860 118.820 ;
        RECT 18.475 118.760 18.765 118.805 ;
        RECT 23.060 118.760 23.380 118.820 ;
        RECT 18.475 118.620 23.380 118.760 ;
        RECT 18.475 118.575 18.765 118.620 ;
        RECT 23.060 118.560 23.380 118.620 ;
        RECT 22.600 118.420 22.920 118.480 ;
        RECT 23.610 118.465 23.750 118.960 ;
        RECT 31.355 118.960 37.180 119.100 ;
        RECT 31.355 118.915 31.645 118.960 ;
        RECT 36.860 118.900 37.180 118.960 ;
        RECT 38.700 118.900 39.020 119.160 ;
        RECT 51.580 119.100 51.900 119.160 ;
        RECT 48.450 118.960 51.900 119.100 ;
        RECT 23.980 118.760 24.300 118.820 ;
        RECT 25.820 118.760 26.140 118.820 ;
        RECT 23.980 118.620 26.140 118.760 ;
        RECT 23.980 118.560 24.300 118.620 ;
        RECT 25.820 118.560 26.140 118.620 ;
        RECT 30.420 118.560 30.740 118.820 ;
        RECT 34.100 118.760 34.420 118.820 ;
        RECT 34.100 118.620 38.470 118.760 ;
        RECT 34.100 118.560 34.420 118.620 ;
        RECT 22.230 118.280 22.920 118.420 ;
        RECT 18.935 118.080 19.225 118.125 ;
        RECT 21.680 118.080 22.000 118.140 ;
        RECT 22.230 118.125 22.370 118.280 ;
        RECT 22.600 118.220 22.920 118.280 ;
        RECT 23.490 118.235 23.780 118.465 ;
        RECT 29.515 118.420 29.805 118.465 ;
        RECT 27.290 118.280 29.805 118.420 ;
        RECT 18.935 117.940 22.000 118.080 ;
        RECT 18.935 117.895 19.225 117.940 ;
        RECT 21.680 117.880 22.000 117.940 ;
        RECT 22.155 117.895 22.445 118.125 ;
        RECT 23.035 118.080 23.325 118.125 ;
        RECT 24.225 118.080 24.515 118.125 ;
        RECT 26.745 118.080 27.035 118.125 ;
        RECT 23.035 117.940 27.035 118.080 ;
        RECT 23.035 117.895 23.325 117.940 ;
        RECT 24.225 117.895 24.515 117.940 ;
        RECT 26.745 117.895 27.035 117.940 ;
        RECT 22.230 117.740 22.370 117.895 ;
        RECT 20.390 117.600 22.370 117.740 ;
        RECT 22.640 117.740 22.930 117.785 ;
        RECT 24.740 117.740 25.030 117.785 ;
        RECT 26.310 117.740 26.600 117.785 ;
        RECT 22.640 117.600 26.600 117.740 ;
        RECT 17.540 117.400 17.860 117.460 ;
        RECT 20.390 117.400 20.530 117.600 ;
        RECT 22.640 117.555 22.930 117.600 ;
        RECT 24.740 117.555 25.030 117.600 ;
        RECT 26.310 117.555 26.600 117.600 ;
        RECT 17.540 117.260 20.530 117.400 ;
        RECT 20.775 117.400 21.065 117.445 ;
        RECT 23.520 117.400 23.840 117.460 ;
        RECT 20.775 117.260 23.840 117.400 ;
        RECT 17.540 117.200 17.860 117.260 ;
        RECT 20.775 117.215 21.065 117.260 ;
        RECT 23.520 117.200 23.840 117.260 ;
        RECT 23.980 117.400 24.300 117.460 ;
        RECT 26.740 117.400 27.060 117.460 ;
        RECT 27.290 117.400 27.430 118.280 ;
        RECT 29.515 118.235 29.805 118.280 ;
        RECT 31.800 118.220 32.120 118.480 ;
        RECT 33.150 118.420 33.440 118.465 ;
        RECT 35.940 118.420 36.260 118.480 ;
        RECT 33.150 118.280 36.260 118.420 ;
        RECT 33.150 118.235 33.440 118.280 ;
        RECT 35.940 118.220 36.260 118.280 ;
        RECT 32.695 118.080 32.985 118.125 ;
        RECT 33.885 118.080 34.175 118.125 ;
        RECT 36.405 118.080 36.695 118.125 ;
        RECT 32.695 117.940 36.695 118.080 ;
        RECT 32.695 117.895 32.985 117.940 ;
        RECT 33.885 117.895 34.175 117.940 ;
        RECT 36.405 117.895 36.695 117.940 ;
        RECT 32.300 117.740 32.590 117.785 ;
        RECT 34.400 117.740 34.690 117.785 ;
        RECT 35.970 117.740 36.260 117.785 ;
        RECT 32.300 117.600 36.260 117.740 ;
        RECT 38.330 117.740 38.470 118.620 ;
        RECT 38.790 118.420 38.930 118.900 ;
        RECT 44.680 118.760 45.000 118.820 ;
        RECT 48.450 118.805 48.590 118.960 ;
        RECT 51.580 118.900 51.900 118.960 ;
        RECT 52.960 119.100 53.280 119.160 ;
        RECT 52.960 118.960 64.230 119.100 ;
        RECT 52.960 118.900 53.280 118.960 ;
        RECT 47.455 118.760 47.745 118.805 ;
        RECT 44.680 118.620 47.745 118.760 ;
        RECT 44.680 118.560 45.000 118.620 ;
        RECT 47.455 118.575 47.745 118.620 ;
        RECT 48.375 118.575 48.665 118.805 ;
        RECT 48.910 118.620 50.890 118.760 ;
        RECT 48.910 118.465 49.050 118.620 ;
        RECT 40.555 118.420 40.845 118.465 ;
        RECT 42.395 118.420 42.685 118.465 ;
        RECT 38.790 118.280 42.685 118.420 ;
        RECT 40.555 118.235 40.845 118.280 ;
        RECT 42.395 118.235 42.685 118.280 ;
        RECT 43.315 118.235 43.605 118.465 ;
        RECT 46.995 118.235 47.285 118.465 ;
        RECT 48.835 118.235 49.125 118.465 ;
        RECT 50.115 118.420 50.405 118.465 ;
        RECT 49.370 118.280 50.405 118.420 ;
        RECT 50.750 118.420 50.890 118.620 ;
        RECT 56.180 118.560 56.500 118.820 ;
        RECT 64.090 118.760 64.230 118.960 ;
        RECT 64.460 118.900 64.780 119.160 ;
        RECT 65.380 119.100 65.700 119.160 ;
        RECT 71.360 119.100 71.680 119.160 ;
        RECT 76.880 119.100 77.200 119.160 ;
        RECT 65.380 118.960 71.680 119.100 ;
        RECT 65.380 118.900 65.700 118.960 ;
        RECT 71.360 118.900 71.680 118.960 ;
        RECT 76.510 118.960 77.200 119.100 ;
        RECT 68.140 118.760 68.460 118.820 ;
        RECT 72.755 118.760 73.045 118.805 ;
        RECT 76.510 118.760 76.650 118.960 ;
        RECT 76.880 118.900 77.200 118.960 ;
        RECT 100.355 118.915 100.645 119.145 ;
        RECT 106.795 119.100 107.085 119.145 ;
        RECT 109.080 119.100 109.400 119.160 ;
        RECT 106.795 118.960 109.400 119.100 ;
        RECT 106.795 118.915 107.085 118.960 ;
        RECT 78.720 118.760 79.040 118.820 ;
        RECT 81.480 118.760 81.800 118.820 ;
        RECT 87.935 118.760 88.225 118.805 ;
        RECT 94.835 118.760 95.125 118.805 ;
        RECT 95.740 118.760 96.060 118.820 ;
        RECT 64.090 118.620 73.045 118.760 ;
        RECT 68.140 118.560 68.460 118.620 ;
        RECT 72.755 118.575 73.045 118.620 ;
        RECT 74.670 118.620 76.650 118.760 ;
        RECT 76.970 118.620 96.060 118.760 ;
        RECT 54.340 118.420 54.660 118.480 ;
        RECT 65.395 118.420 65.685 118.465 ;
        RECT 50.750 118.280 65.685 118.420 ;
        RECT 41.920 117.880 42.240 118.140 ;
        RECT 43.390 117.740 43.530 118.235 ;
        RECT 47.070 118.080 47.210 118.235 ;
        RECT 47.900 118.080 48.220 118.140 ;
        RECT 49.370 118.080 49.510 118.280 ;
        RECT 50.115 118.235 50.405 118.280 ;
        RECT 54.340 118.220 54.660 118.280 ;
        RECT 60.410 118.140 60.550 118.280 ;
        RECT 65.395 118.235 65.685 118.280 ;
        RECT 65.840 118.420 66.160 118.480 ;
        RECT 66.675 118.420 66.965 118.465 ;
        RECT 73.675 118.420 73.965 118.465 ;
        RECT 65.840 118.280 66.965 118.420 ;
        RECT 65.840 118.220 66.160 118.280 ;
        RECT 66.675 118.235 66.965 118.280 ;
        RECT 72.370 118.280 73.965 118.420 ;
        RECT 47.070 117.940 48.220 118.080 ;
        RECT 47.900 117.880 48.220 117.940 ;
        RECT 48.450 117.940 49.510 118.080 ;
        RECT 49.715 118.080 50.005 118.125 ;
        RECT 50.905 118.080 51.195 118.125 ;
        RECT 53.425 118.080 53.715 118.125 ;
        RECT 49.715 117.940 53.715 118.080 ;
        RECT 48.450 117.785 48.590 117.940 ;
        RECT 49.715 117.895 50.005 117.940 ;
        RECT 50.905 117.895 51.195 117.940 ;
        RECT 53.425 117.895 53.715 117.940 ;
        RECT 60.320 117.880 60.640 118.140 ;
        RECT 61.715 118.080 62.005 118.125 ;
        RECT 64.000 118.080 64.320 118.140 ;
        RECT 61.715 117.940 64.320 118.080 ;
        RECT 61.715 117.895 62.005 117.940 ;
        RECT 64.000 117.880 64.320 117.940 ;
        RECT 66.275 118.080 66.565 118.125 ;
        RECT 67.465 118.080 67.755 118.125 ;
        RECT 69.985 118.080 70.275 118.125 ;
        RECT 66.275 117.940 70.275 118.080 ;
        RECT 66.275 117.895 66.565 117.940 ;
        RECT 67.465 117.895 67.755 117.940 ;
        RECT 69.985 117.895 70.275 117.940 ;
        RECT 38.330 117.600 43.530 117.740 ;
        RECT 32.300 117.555 32.590 117.600 ;
        RECT 34.400 117.555 34.690 117.600 ;
        RECT 35.970 117.555 36.260 117.600 ;
        RECT 48.375 117.555 48.665 117.785 ;
        RECT 49.320 117.740 49.610 117.785 ;
        RECT 51.420 117.740 51.710 117.785 ;
        RECT 52.990 117.740 53.280 117.785 ;
        RECT 49.320 117.600 53.280 117.740 ;
        RECT 49.320 117.555 49.610 117.600 ;
        RECT 51.420 117.555 51.710 117.600 ;
        RECT 52.990 117.555 53.280 117.600 ;
        RECT 55.720 117.540 56.040 117.800 ;
        RECT 58.940 117.740 59.260 117.800 ;
        RECT 65.880 117.740 66.170 117.785 ;
        RECT 67.980 117.740 68.270 117.785 ;
        RECT 69.550 117.740 69.840 117.785 ;
        RECT 58.940 117.600 65.150 117.740 ;
        RECT 58.940 117.540 59.260 117.600 ;
        RECT 23.980 117.260 27.430 117.400 ;
        RECT 29.055 117.400 29.345 117.445 ;
        RECT 30.880 117.400 31.200 117.460 ;
        RECT 35.020 117.400 35.340 117.460 ;
        RECT 29.055 117.260 35.340 117.400 ;
        RECT 23.980 117.200 24.300 117.260 ;
        RECT 26.740 117.200 27.060 117.260 ;
        RECT 29.055 117.215 29.345 117.260 ;
        RECT 30.880 117.200 31.200 117.260 ;
        RECT 35.020 117.200 35.340 117.260 ;
        RECT 39.620 117.200 39.940 117.460 ;
        RECT 40.080 117.400 40.400 117.460 ;
        RECT 41.475 117.400 41.765 117.445 ;
        RECT 41.920 117.400 42.240 117.460 ;
        RECT 40.080 117.260 42.240 117.400 ;
        RECT 40.080 117.200 40.400 117.260 ;
        RECT 41.475 117.215 41.765 117.260 ;
        RECT 41.920 117.200 42.240 117.260 ;
        RECT 44.220 117.200 44.540 117.460 ;
        RECT 65.010 117.400 65.150 117.600 ;
        RECT 65.880 117.600 69.840 117.740 ;
        RECT 65.880 117.555 66.170 117.600 ;
        RECT 67.980 117.555 68.270 117.600 ;
        RECT 69.550 117.555 69.840 117.600 ;
        RECT 66.760 117.400 67.080 117.460 ;
        RECT 65.010 117.260 67.080 117.400 ;
        RECT 66.760 117.200 67.080 117.260 ;
        RECT 68.600 117.400 68.920 117.460 ;
        RECT 69.980 117.400 70.300 117.460 ;
        RECT 68.600 117.260 70.300 117.400 ;
        RECT 68.600 117.200 68.920 117.260 ;
        RECT 69.980 117.200 70.300 117.260 ;
        RECT 71.360 117.400 71.680 117.460 ;
        RECT 72.370 117.445 72.510 118.280 ;
        RECT 73.675 118.235 73.965 118.280 ;
        RECT 74.120 118.420 74.440 118.480 ;
        RECT 74.670 118.465 74.810 118.620 ;
        RECT 74.595 118.420 74.885 118.465 ;
        RECT 74.120 118.280 74.885 118.420 ;
        RECT 73.750 118.080 73.890 118.235 ;
        RECT 74.120 118.220 74.440 118.280 ;
        RECT 74.595 118.235 74.885 118.280 ;
        RECT 75.055 118.235 75.345 118.465 ;
        RECT 75.130 118.080 75.270 118.235 ;
        RECT 75.500 118.220 75.820 118.480 ;
        RECT 76.970 118.465 77.110 118.620 ;
        RECT 78.720 118.560 79.040 118.620 ;
        RECT 81.480 118.560 81.800 118.620 ;
        RECT 87.935 118.575 88.225 118.620 ;
        RECT 94.835 118.575 95.125 118.620 ;
        RECT 95.740 118.560 96.060 118.620 ;
        RECT 96.675 118.760 96.965 118.805 ;
        RECT 97.120 118.760 97.440 118.820 ;
        RECT 99.880 118.760 100.200 118.820 ;
        RECT 96.675 118.620 100.200 118.760 ;
        RECT 96.675 118.575 96.965 118.620 ;
        RECT 97.120 118.560 97.440 118.620 ;
        RECT 99.880 118.560 100.200 118.620 ;
        RECT 78.260 118.465 78.580 118.480 ;
        RECT 76.895 118.235 77.185 118.465 ;
        RECT 78.230 118.420 78.580 118.465 ;
        RECT 78.065 118.280 78.580 118.420 ;
        RECT 78.230 118.235 78.580 118.280 ;
        RECT 78.260 118.220 78.580 118.235 ;
        RECT 80.560 118.420 80.880 118.480 ;
        RECT 80.560 118.280 84.010 118.420 ;
        RECT 80.560 118.220 80.880 118.280 ;
        RECT 75.960 118.080 76.280 118.140 ;
        RECT 73.750 117.940 76.280 118.080 ;
        RECT 75.960 117.880 76.280 117.940 ;
        RECT 76.420 117.880 76.740 118.140 ;
        RECT 77.775 118.080 78.065 118.125 ;
        RECT 78.965 118.080 79.255 118.125 ;
        RECT 81.485 118.080 81.775 118.125 ;
        RECT 77.775 117.940 81.775 118.080 ;
        RECT 77.775 117.895 78.065 117.940 ;
        RECT 78.965 117.895 79.255 117.940 ;
        RECT 81.485 117.895 81.775 117.940 ;
        RECT 83.870 118.080 84.010 118.280 ;
        RECT 91.140 118.220 91.460 118.480 ;
        RECT 92.060 118.420 92.380 118.480 ;
        RECT 96.200 118.420 96.520 118.480 ;
        RECT 92.060 118.280 96.520 118.420 ;
        RECT 100.430 118.420 100.570 118.915 ;
        RECT 109.080 118.900 109.400 118.960 ;
        RECT 111.380 119.100 111.700 119.160 ;
        RECT 112.760 119.100 113.080 119.160 ;
        RECT 111.380 118.960 113.080 119.100 ;
        RECT 111.380 118.900 111.700 118.960 ;
        RECT 112.760 118.900 113.080 118.960 ;
        RECT 118.740 119.100 119.060 119.160 ;
        RECT 122.880 119.100 123.200 119.160 ;
        RECT 124.720 119.100 125.040 119.160 ;
        RECT 118.740 118.960 125.040 119.100 ;
        RECT 118.740 118.900 119.060 118.960 ;
        RECT 122.880 118.900 123.200 118.960 ;
        RECT 124.720 118.900 125.040 118.960 ;
        RECT 126.575 119.100 126.865 119.145 ;
        RECT 126.575 118.960 127.710 119.100 ;
        RECT 126.575 118.915 126.865 118.960 ;
        RECT 101.260 118.560 101.580 118.820 ;
        RECT 112.300 118.760 112.620 118.820 ;
        RECT 120.595 118.760 120.885 118.805 ;
        RECT 127.570 118.760 127.710 118.960 ;
        RECT 128.260 118.760 128.550 118.805 ;
        RECT 136.235 118.760 136.525 118.805 ;
        RECT 112.300 118.620 127.250 118.760 ;
        RECT 127.570 118.620 128.550 118.760 ;
        RECT 112.300 118.560 112.620 118.620 ;
        RECT 120.595 118.575 120.885 118.620 ;
        RECT 127.110 118.480 127.250 118.620 ;
        RECT 128.260 118.575 128.550 118.620 ;
        RECT 130.330 118.620 136.525 118.760 ;
        RECT 103.100 118.420 103.420 118.480 ;
        RECT 100.430 118.280 103.420 118.420 ;
        RECT 92.060 118.220 92.380 118.280 ;
        RECT 96.200 118.220 96.520 118.280 ;
        RECT 103.100 118.220 103.420 118.280 ;
        RECT 105.860 118.220 106.180 118.480 ;
        RECT 108.160 118.220 108.480 118.480 ;
        RECT 109.095 118.420 109.385 118.465 ;
        RECT 109.095 118.280 114.370 118.420 ;
        RECT 109.095 118.235 109.385 118.280 ;
        RECT 99.880 118.080 100.200 118.140 ;
        RECT 102.640 118.080 102.960 118.140 ;
        RECT 83.870 117.940 100.200 118.080 ;
        RECT 74.580 117.740 74.900 117.800 ;
        RECT 83.870 117.785 84.010 117.940 ;
        RECT 99.880 117.880 100.200 117.940 ;
        RECT 100.430 117.940 102.960 118.080 ;
        RECT 114.230 118.080 114.370 118.280 ;
        RECT 114.600 118.220 114.920 118.480 ;
        RECT 115.520 118.420 115.840 118.480 ;
        RECT 117.835 118.420 118.125 118.465 ;
        RECT 115.520 118.280 118.125 118.420 ;
        RECT 115.520 118.220 115.840 118.280 ;
        RECT 117.835 118.235 118.125 118.280 ;
        RECT 118.280 118.220 118.600 118.480 ;
        RECT 118.755 118.235 119.045 118.465 ;
        RECT 118.830 118.080 118.970 118.235 ;
        RECT 119.660 118.220 119.980 118.480 ;
        RECT 123.340 118.220 123.660 118.480 ;
        RECT 124.275 118.235 124.565 118.465 ;
        RECT 121.960 118.080 122.280 118.140 ;
        RECT 114.230 117.940 122.280 118.080 ;
        RECT 124.350 118.080 124.490 118.235 ;
        RECT 124.720 118.220 125.040 118.480 ;
        RECT 125.195 118.420 125.485 118.465 ;
        RECT 126.560 118.420 126.880 118.480 ;
        RECT 125.195 118.280 126.880 118.420 ;
        RECT 125.195 118.235 125.485 118.280 ;
        RECT 126.560 118.220 126.880 118.280 ;
        RECT 127.020 118.220 127.340 118.480 ;
        RECT 130.330 118.420 130.470 118.620 ;
        RECT 136.235 118.575 136.525 118.620 ;
        RECT 127.570 118.280 130.470 118.420 ;
        RECT 127.570 118.080 127.710 118.280 ;
        RECT 134.380 118.220 134.700 118.480 ;
        RECT 135.315 118.420 135.605 118.465 ;
        RECT 135.760 118.420 136.080 118.480 ;
        RECT 135.315 118.280 136.080 118.420 ;
        RECT 135.315 118.235 135.605 118.280 ;
        RECT 124.350 117.940 127.710 118.080 ;
        RECT 127.915 118.080 128.205 118.125 ;
        RECT 129.105 118.080 129.395 118.125 ;
        RECT 131.625 118.080 131.915 118.125 ;
        RECT 135.390 118.080 135.530 118.235 ;
        RECT 135.760 118.220 136.080 118.280 ;
        RECT 127.915 117.940 131.915 118.080 ;
        RECT 77.380 117.740 77.670 117.785 ;
        RECT 79.480 117.740 79.770 117.785 ;
        RECT 81.050 117.740 81.340 117.785 ;
        RECT 74.580 117.600 76.190 117.740 ;
        RECT 74.580 117.540 74.900 117.600 ;
        RECT 76.050 117.445 76.190 117.600 ;
        RECT 77.380 117.600 81.340 117.740 ;
        RECT 77.380 117.555 77.670 117.600 ;
        RECT 79.480 117.555 79.770 117.600 ;
        RECT 81.050 117.555 81.340 117.600 ;
        RECT 83.795 117.555 84.085 117.785 ;
        RECT 96.660 117.740 96.980 117.800 ;
        RECT 99.435 117.740 99.725 117.785 ;
        RECT 96.660 117.600 99.725 117.740 ;
        RECT 96.660 117.540 96.980 117.600 ;
        RECT 99.435 117.555 99.725 117.600 ;
        RECT 100.430 117.445 100.570 117.940 ;
        RECT 102.640 117.880 102.960 117.940 ;
        RECT 121.960 117.880 122.280 117.940 ;
        RECT 127.915 117.895 128.205 117.940 ;
        RECT 129.105 117.895 129.395 117.940 ;
        RECT 131.625 117.895 131.915 117.940 ;
        RECT 134.010 117.940 135.530 118.080 ;
        RECT 112.760 117.740 113.080 117.800 ;
        RECT 115.535 117.740 115.825 117.785 ;
        RECT 125.180 117.740 125.500 117.800 ;
        RECT 112.760 117.600 125.500 117.740 ;
        RECT 112.760 117.540 113.080 117.600 ;
        RECT 115.535 117.555 115.825 117.600 ;
        RECT 125.180 117.540 125.500 117.600 ;
        RECT 127.520 117.740 127.810 117.785 ;
        RECT 129.620 117.740 129.910 117.785 ;
        RECT 131.190 117.740 131.480 117.785 ;
        RECT 127.520 117.600 131.480 117.740 ;
        RECT 127.520 117.555 127.810 117.600 ;
        RECT 129.620 117.555 129.910 117.600 ;
        RECT 131.190 117.555 131.480 117.600 ;
        RECT 132.080 117.740 132.400 117.800 ;
        RECT 134.010 117.785 134.150 117.940 ;
        RECT 133.935 117.740 134.225 117.785 ;
        RECT 132.080 117.600 134.225 117.740 ;
        RECT 132.080 117.540 132.400 117.600 ;
        RECT 133.935 117.555 134.225 117.600 ;
        RECT 72.295 117.400 72.585 117.445 ;
        RECT 71.360 117.260 72.585 117.400 ;
        RECT 71.360 117.200 71.680 117.260 ;
        RECT 72.295 117.215 72.585 117.260 ;
        RECT 75.975 117.215 76.265 117.445 ;
        RECT 100.355 117.215 100.645 117.445 ;
        RECT 102.190 117.400 102.485 117.475 ;
        RECT 104.950 117.400 105.245 117.475 ;
        RECT 102.190 117.260 105.245 117.400 ;
        RECT 102.190 117.205 102.485 117.260 ;
        RECT 104.950 117.205 105.245 117.260 ;
        RECT 111.380 117.400 111.700 117.460 ;
        RECT 116.915 117.400 117.205 117.445 ;
        RECT 111.380 117.260 117.205 117.400 ;
        RECT 111.380 117.200 111.700 117.260 ;
        RECT 116.915 117.215 117.205 117.260 ;
        RECT 13.330 116.580 138.910 117.060 ;
        RECT 19.855 116.380 20.145 116.425 ;
        RECT 21.680 116.380 22.000 116.440 ;
        RECT 19.855 116.240 22.000 116.380 ;
        RECT 19.855 116.195 20.145 116.240 ;
        RECT 21.680 116.180 22.000 116.240 ;
        RECT 23.520 116.180 23.840 116.440 ;
        RECT 35.940 116.180 36.260 116.440 ;
        RECT 36.860 116.180 37.180 116.440 ;
        RECT 44.680 116.380 45.000 116.440 ;
        RECT 46.075 116.380 46.365 116.425 ;
        RECT 44.680 116.240 46.365 116.380 ;
        RECT 44.680 116.180 45.000 116.240 ;
        RECT 46.075 116.195 46.365 116.240 ;
        RECT 65.380 116.380 65.700 116.440 ;
        RECT 66.315 116.380 66.605 116.425 ;
        RECT 65.380 116.240 66.605 116.380 ;
        RECT 65.380 116.180 65.700 116.240 ;
        RECT 66.315 116.195 66.605 116.240 ;
        RECT 66.760 116.380 67.080 116.440 ;
        RECT 67.695 116.380 67.985 116.425 ;
        RECT 66.760 116.240 67.985 116.380 ;
        RECT 66.760 116.180 67.080 116.240 ;
        RECT 67.695 116.195 67.985 116.240 ;
        RECT 68.615 116.195 68.905 116.425 ;
        RECT 83.780 116.380 84.100 116.440 ;
        RECT 76.970 116.240 84.100 116.380 ;
        RECT 22.615 116.040 22.905 116.085 ;
        RECT 24.440 116.040 24.760 116.100 ;
        RECT 35.480 116.040 35.800 116.100 ;
        RECT 38.240 116.040 38.560 116.100 ;
        RECT 38.715 116.040 39.005 116.085 ;
        RECT 22.615 115.900 24.760 116.040 ;
        RECT 22.615 115.855 22.905 115.900 ;
        RECT 24.440 115.840 24.760 115.900 ;
        RECT 28.670 115.900 35.250 116.040 ;
        RECT 22.230 115.560 26.050 115.700 ;
        RECT 22.230 115.405 22.370 115.560 ;
        RECT 25.910 115.420 26.050 115.560 ;
        RECT 21.695 115.360 21.985 115.405 ;
        RECT 22.155 115.360 22.445 115.405 ;
        RECT 21.695 115.220 22.445 115.360 ;
        RECT 21.695 115.175 21.985 115.220 ;
        RECT 22.155 115.175 22.445 115.220 ;
        RECT 23.075 115.175 23.365 115.405 ;
        RECT 24.455 115.175 24.745 115.405 ;
        RECT 19.855 115.020 20.145 115.065 ;
        RECT 20.760 115.020 21.080 115.080 ;
        RECT 19.855 114.880 21.080 115.020 ;
        RECT 19.855 114.835 20.145 114.880 ;
        RECT 20.760 114.820 21.080 114.880 ;
        RECT 18.935 114.680 19.225 114.725 ;
        RECT 19.380 114.680 19.700 114.740 ;
        RECT 18.935 114.540 19.700 114.680 ;
        RECT 23.150 114.680 23.290 115.175 ;
        RECT 24.530 115.020 24.670 115.175 ;
        RECT 25.360 115.160 25.680 115.420 ;
        RECT 25.820 115.160 26.140 115.420 ;
        RECT 27.200 115.160 27.520 115.420 ;
        RECT 27.675 115.175 27.965 115.405 ;
        RECT 27.750 115.020 27.890 115.175 ;
        RECT 28.120 115.160 28.440 115.420 ;
        RECT 28.670 115.405 28.810 115.900 ;
        RECT 29.515 115.700 29.805 115.745 ;
        RECT 33.655 115.700 33.945 115.745 ;
        RECT 29.515 115.560 33.945 115.700 ;
        RECT 35.110 115.700 35.250 115.900 ;
        RECT 35.480 115.900 39.005 116.040 ;
        RECT 35.480 115.840 35.800 115.900 ;
        RECT 38.240 115.840 38.560 115.900 ;
        RECT 38.715 115.855 39.005 115.900 ;
        RECT 45.155 115.855 45.445 116.085 ;
        RECT 52.515 116.040 52.805 116.085 ;
        RECT 48.910 115.900 52.805 116.040 ;
        RECT 36.400 115.700 36.720 115.760 ;
        RECT 35.110 115.560 36.720 115.700 ;
        RECT 29.515 115.515 29.805 115.560 ;
        RECT 33.655 115.515 33.945 115.560 ;
        RECT 36.400 115.500 36.720 115.560 ;
        RECT 36.860 115.700 37.180 115.760 ;
        RECT 45.230 115.700 45.370 115.855 ;
        RECT 48.910 115.745 49.050 115.900 ;
        RECT 52.515 115.855 52.805 115.900 ;
        RECT 55.260 116.040 55.550 116.085 ;
        RECT 56.830 116.040 57.120 116.085 ;
        RECT 58.930 116.040 59.220 116.085 ;
        RECT 55.260 115.900 59.220 116.040 ;
        RECT 55.260 115.855 55.550 115.900 ;
        RECT 56.830 115.855 57.120 115.900 ;
        RECT 58.930 115.855 59.220 115.900 ;
        RECT 63.080 116.040 63.400 116.100 ;
        RECT 68.690 116.040 68.830 116.195 ;
        RECT 63.080 115.900 68.830 116.040 ;
        RECT 63.080 115.840 63.400 115.900 ;
        RECT 36.860 115.560 45.370 115.700 ;
        RECT 47.915 115.700 48.205 115.745 ;
        RECT 48.835 115.700 49.125 115.745 ;
        RECT 47.915 115.560 49.125 115.700 ;
        RECT 36.860 115.500 37.180 115.560 ;
        RECT 47.915 115.515 48.205 115.560 ;
        RECT 48.835 115.515 49.125 115.560 ;
        RECT 54.825 115.700 55.115 115.745 ;
        RECT 57.345 115.700 57.635 115.745 ;
        RECT 58.535 115.700 58.825 115.745 ;
        RECT 54.825 115.560 58.825 115.700 ;
        RECT 54.825 115.515 55.115 115.560 ;
        RECT 57.345 115.515 57.635 115.560 ;
        RECT 58.535 115.515 58.825 115.560 ;
        RECT 59.860 115.700 60.180 115.760 ;
        RECT 62.620 115.700 62.940 115.760 ;
        RECT 63.555 115.700 63.845 115.745 ;
        RECT 59.860 115.560 63.845 115.700 ;
        RECT 59.860 115.500 60.180 115.560 ;
        RECT 62.620 115.500 62.940 115.560 ;
        RECT 63.555 115.515 63.845 115.560 ;
        RECT 66.300 115.700 66.620 115.760 ;
        RECT 70.440 115.700 70.760 115.760 ;
        RECT 66.300 115.560 70.760 115.700 ;
        RECT 66.300 115.500 66.620 115.560 ;
        RECT 70.440 115.500 70.760 115.560 ;
        RECT 73.215 115.700 73.505 115.745 ;
        RECT 74.120 115.700 74.440 115.760 ;
        RECT 73.215 115.560 74.440 115.700 ;
        RECT 73.215 115.515 73.505 115.560 ;
        RECT 28.595 115.175 28.885 115.405 ;
        RECT 31.340 115.360 31.660 115.420 ;
        RECT 31.815 115.360 32.105 115.405 ;
        RECT 31.340 115.220 32.105 115.360 ;
        RECT 31.340 115.160 31.660 115.220 ;
        RECT 31.815 115.175 32.105 115.220 ;
        RECT 32.735 115.175 33.025 115.405 ;
        RECT 33.195 115.360 33.485 115.405 ;
        RECT 34.100 115.360 34.420 115.420 ;
        RECT 33.195 115.220 34.420 115.360 ;
        RECT 33.195 115.175 33.485 115.220 ;
        RECT 29.500 115.020 29.820 115.080 ;
        RECT 24.530 114.880 26.050 115.020 ;
        RECT 27.750 114.880 29.820 115.020 ;
        RECT 32.810 115.020 32.950 115.175 ;
        RECT 34.100 115.160 34.420 115.220 ;
        RECT 34.575 115.360 34.865 115.405 ;
        RECT 37.320 115.360 37.640 115.420 ;
        RECT 34.575 115.220 37.640 115.360 ;
        RECT 34.575 115.175 34.865 115.220 ;
        RECT 37.320 115.160 37.640 115.220 ;
        RECT 40.540 115.160 40.860 115.420 ;
        RECT 41.000 115.360 41.320 115.420 ;
        RECT 41.000 115.220 41.515 115.360 ;
        RECT 41.000 115.160 41.320 115.220 ;
        RECT 42.380 115.160 42.700 115.420 ;
        RECT 43.085 115.360 43.375 115.405 ;
        RECT 43.760 115.360 44.080 115.420 ;
        RECT 43.085 115.220 44.080 115.360 ;
        RECT 43.085 115.175 43.375 115.220 ;
        RECT 43.760 115.160 44.080 115.220 ;
        RECT 59.415 115.360 59.705 115.405 ;
        RECT 60.320 115.360 60.640 115.420 ;
        RECT 59.415 115.220 60.640 115.360 ;
        RECT 59.415 115.175 59.705 115.220 ;
        RECT 60.320 115.160 60.640 115.220 ;
        RECT 62.175 115.175 62.465 115.405 ;
        RECT 63.095 115.175 63.385 115.405 ;
        RECT 64.000 115.360 64.320 115.420 ;
        RECT 66.775 115.360 67.065 115.405 ;
        RECT 64.000 115.220 67.065 115.360 ;
        RECT 39.620 115.020 39.940 115.080 ;
        RECT 32.810 114.880 39.940 115.020 ;
        RECT 25.360 114.680 25.680 114.740 ;
        RECT 23.150 114.540 25.680 114.680 ;
        RECT 25.910 114.680 26.050 114.880 ;
        RECT 29.500 114.820 29.820 114.880 ;
        RECT 39.620 114.820 39.940 114.880 ;
        RECT 41.935 114.835 42.225 115.065 ;
        RECT 53.420 115.020 53.740 115.080 ;
        RECT 42.930 114.880 53.740 115.020 ;
        RECT 30.880 114.680 31.200 114.740 ;
        RECT 25.910 114.540 31.200 114.680 ;
        RECT 18.935 114.495 19.225 114.540 ;
        RECT 19.380 114.480 19.700 114.540 ;
        RECT 25.360 114.480 25.680 114.540 ;
        RECT 30.880 114.480 31.200 114.540 ;
        RECT 35.480 114.480 35.800 114.740 ;
        RECT 36.860 114.480 37.180 114.740 ;
        RECT 42.010 114.680 42.150 114.835 ;
        RECT 42.930 114.680 43.070 114.880 ;
        RECT 53.420 114.820 53.740 114.880 ;
        RECT 58.190 115.020 58.480 115.065 ;
        RECT 61.255 115.020 61.545 115.065 ;
        RECT 58.190 114.880 61.545 115.020 ;
        RECT 58.190 114.835 58.480 114.880 ;
        RECT 61.255 114.835 61.545 114.880 ;
        RECT 42.010 114.540 43.070 114.680 ;
        RECT 43.300 114.680 43.620 114.740 ;
        RECT 43.775 114.680 44.065 114.725 ;
        RECT 43.300 114.540 44.065 114.680 ;
        RECT 43.300 114.480 43.620 114.540 ;
        RECT 43.775 114.495 44.065 114.540 ;
        RECT 46.075 114.680 46.365 114.725 ;
        RECT 47.900 114.680 48.220 114.740 ;
        RECT 46.075 114.540 48.220 114.680 ;
        RECT 46.075 114.495 46.365 114.540 ;
        RECT 47.900 114.480 48.220 114.540 ;
        RECT 51.580 114.680 51.900 114.740 ;
        RECT 62.250 114.680 62.390 115.175 ;
        RECT 62.620 115.020 62.940 115.080 ;
        RECT 63.170 115.020 63.310 115.175 ;
        RECT 64.000 115.160 64.320 115.220 ;
        RECT 66.775 115.175 67.065 115.220 ;
        RECT 67.235 115.360 67.525 115.405 ;
        RECT 70.900 115.360 71.220 115.420 ;
        RECT 73.290 115.360 73.430 115.515 ;
        RECT 74.120 115.500 74.440 115.560 ;
        RECT 74.595 115.700 74.885 115.745 ;
        RECT 75.040 115.700 75.360 115.760 ;
        RECT 74.595 115.560 75.360 115.700 ;
        RECT 74.595 115.515 74.885 115.560 ;
        RECT 75.040 115.500 75.360 115.560 ;
        RECT 76.970 115.360 77.110 116.240 ;
        RECT 83.780 116.180 84.100 116.240 ;
        RECT 94.820 116.180 95.140 116.440 ;
        RECT 104.020 116.380 104.340 116.440 ;
        RECT 104.495 116.380 104.785 116.425 ;
        RECT 112.300 116.380 112.620 116.440 ;
        RECT 104.020 116.240 112.620 116.380 ;
        RECT 104.020 116.180 104.340 116.240 ;
        RECT 104.495 116.195 104.785 116.240 ;
        RECT 112.300 116.180 112.620 116.240 ;
        RECT 77.355 115.855 77.645 116.085 ;
        RECT 78.760 116.040 79.050 116.085 ;
        RECT 80.860 116.040 81.150 116.085 ;
        RECT 82.430 116.040 82.720 116.085 ;
        RECT 78.760 115.900 82.720 116.040 ;
        RECT 78.760 115.855 79.050 115.900 ;
        RECT 80.860 115.855 81.150 115.900 ;
        RECT 82.430 115.855 82.720 115.900 ;
        RECT 98.040 116.040 98.360 116.100 ;
        RECT 110.920 116.040 111.240 116.100 ;
        RECT 98.040 115.900 111.240 116.040 ;
        RECT 67.235 115.220 73.430 115.360 ;
        RECT 75.130 115.220 77.110 115.360 ;
        RECT 67.235 115.175 67.525 115.220 ;
        RECT 70.900 115.160 71.220 115.220 ;
        RECT 68.140 115.065 68.460 115.080 ;
        RECT 68.140 115.020 68.745 115.065 ;
        RECT 62.620 114.880 68.895 115.020 ;
        RECT 62.620 114.820 62.940 114.880 ;
        RECT 68.140 114.835 68.745 114.880 ;
        RECT 68.140 114.820 68.460 114.835 ;
        RECT 69.520 114.820 69.840 115.080 ;
        RECT 70.440 115.020 70.760 115.080 ;
        RECT 75.130 115.065 75.270 115.220 ;
        RECT 75.055 115.020 75.345 115.065 ;
        RECT 70.440 114.880 75.345 115.020 ;
        RECT 77.430 115.020 77.570 115.855 ;
        RECT 98.040 115.840 98.360 115.900 ;
        RECT 110.920 115.840 111.240 115.900 ;
        RECT 111.880 116.040 112.170 116.085 ;
        RECT 113.980 116.040 114.270 116.085 ;
        RECT 115.550 116.040 115.840 116.085 ;
        RECT 111.880 115.900 115.840 116.040 ;
        RECT 111.880 115.855 112.170 115.900 ;
        RECT 113.980 115.855 114.270 115.900 ;
        RECT 115.550 115.855 115.840 115.900 ;
        RECT 130.280 116.040 130.570 116.085 ;
        RECT 132.380 116.040 132.670 116.085 ;
        RECT 133.950 116.040 134.240 116.085 ;
        RECT 130.280 115.900 134.240 116.040 ;
        RECT 130.280 115.855 130.570 115.900 ;
        RECT 132.380 115.855 132.670 115.900 ;
        RECT 133.950 115.855 134.240 115.900 ;
        RECT 79.155 115.700 79.445 115.745 ;
        RECT 80.345 115.700 80.635 115.745 ;
        RECT 82.865 115.700 83.155 115.745 ;
        RECT 79.155 115.560 83.155 115.700 ;
        RECT 79.155 115.515 79.445 115.560 ;
        RECT 80.345 115.515 80.635 115.560 ;
        RECT 82.865 115.515 83.155 115.560 ;
        RECT 92.980 115.700 93.300 115.760 ;
        RECT 108.160 115.700 108.480 115.760 ;
        RECT 92.980 115.560 102.410 115.700 ;
        RECT 92.980 115.500 93.300 115.560 ;
        RECT 78.275 115.360 78.565 115.405 ;
        RECT 78.720 115.360 79.040 115.420 ;
        RECT 78.275 115.220 79.040 115.360 ;
        RECT 78.275 115.175 78.565 115.220 ;
        RECT 78.720 115.160 79.040 115.220 ;
        RECT 95.295 115.360 95.585 115.405 ;
        RECT 97.120 115.360 97.440 115.420 ;
        RECT 102.270 115.405 102.410 115.560 ;
        RECT 104.110 115.560 108.480 115.700 ;
        RECT 104.110 115.405 104.250 115.560 ;
        RECT 108.160 115.500 108.480 115.560 ;
        RECT 112.275 115.700 112.565 115.745 ;
        RECT 113.465 115.700 113.755 115.745 ;
        RECT 115.985 115.700 116.275 115.745 ;
        RECT 127.480 115.700 127.800 115.760 ;
        RECT 129.795 115.700 130.085 115.745 ;
        RECT 112.275 115.560 116.275 115.700 ;
        RECT 112.275 115.515 112.565 115.560 ;
        RECT 113.465 115.515 113.755 115.560 ;
        RECT 115.985 115.515 116.275 115.560 ;
        RECT 122.510 115.560 130.085 115.700 ;
        RECT 95.295 115.220 97.440 115.360 ;
        RECT 95.295 115.175 95.585 115.220 ;
        RECT 97.120 115.160 97.440 115.220 ;
        RECT 97.595 115.360 97.885 115.405 ;
        RECT 98.975 115.360 99.265 115.405 ;
        RECT 97.595 115.220 99.265 115.360 ;
        RECT 97.595 115.175 97.885 115.220 ;
        RECT 98.975 115.175 99.265 115.220 ;
        RECT 101.735 115.175 102.025 115.405 ;
        RECT 102.195 115.360 102.485 115.405 ;
        RECT 104.035 115.360 104.325 115.405 ;
        RECT 102.195 115.220 104.325 115.360 ;
        RECT 102.195 115.175 102.485 115.220 ;
        RECT 104.035 115.175 104.325 115.220 ;
        RECT 105.415 115.175 105.705 115.405 ;
        RECT 111.395 115.360 111.685 115.405 ;
        RECT 111.840 115.360 112.160 115.420 ;
        RECT 122.510 115.405 122.650 115.560 ;
        RECT 127.480 115.500 127.800 115.560 ;
        RECT 129.795 115.515 130.085 115.560 ;
        RECT 130.675 115.700 130.965 115.745 ;
        RECT 131.865 115.700 132.155 115.745 ;
        RECT 134.385 115.700 134.675 115.745 ;
        RECT 130.675 115.560 134.675 115.700 ;
        RECT 130.675 115.515 130.965 115.560 ;
        RECT 131.865 115.515 132.155 115.560 ;
        RECT 134.385 115.515 134.675 115.560 ;
        RECT 122.435 115.360 122.725 115.405 ;
        RECT 111.395 115.220 122.725 115.360 ;
        RECT 111.395 115.175 111.685 115.220 ;
        RECT 79.500 115.020 79.790 115.065 ;
        RECT 77.430 114.880 79.790 115.020 ;
        RECT 70.440 114.820 70.760 114.880 ;
        RECT 75.055 114.835 75.345 114.880 ;
        RECT 79.500 114.835 79.790 114.880 ;
        RECT 85.620 115.020 85.940 115.080 ;
        RECT 88.395 115.020 88.685 115.065 ;
        RECT 85.620 114.880 88.685 115.020 ;
        RECT 85.620 114.820 85.940 114.880 ;
        RECT 88.395 114.835 88.685 114.880 ;
        RECT 96.215 115.020 96.505 115.065 ;
        RECT 97.670 115.020 97.810 115.175 ;
        RECT 96.215 114.880 97.810 115.020 ;
        RECT 99.435 115.020 99.725 115.065 ;
        RECT 101.810 115.020 101.950 115.175 ;
        RECT 105.490 115.020 105.630 115.175 ;
        RECT 111.840 115.160 112.160 115.220 ;
        RECT 122.435 115.175 122.725 115.220 ;
        RECT 123.340 115.360 123.660 115.420 ;
        RECT 123.815 115.360 124.105 115.405 ;
        RECT 123.340 115.220 124.105 115.360 ;
        RECT 123.340 115.160 123.660 115.220 ;
        RECT 123.815 115.175 124.105 115.220 ;
        RECT 124.735 115.175 125.025 115.405 ;
        RECT 112.760 115.065 113.080 115.080 ;
        RECT 99.435 114.880 105.630 115.020 ;
        RECT 96.215 114.835 96.505 114.880 ;
        RECT 99.435 114.835 99.725 114.880 ;
        RECT 51.580 114.540 62.390 114.680 ;
        RECT 64.920 114.680 65.240 114.740 ;
        RECT 65.395 114.680 65.685 114.725 ;
        RECT 64.920 114.540 65.685 114.680 ;
        RECT 51.580 114.480 51.900 114.540 ;
        RECT 64.920 114.480 65.240 114.540 ;
        RECT 65.395 114.495 65.685 114.540 ;
        RECT 69.980 114.480 70.300 114.740 ;
        RECT 75.515 114.680 75.805 114.725 ;
        RECT 85.175 114.680 85.465 114.725 ;
        RECT 87.000 114.680 87.320 114.740 ;
        RECT 75.515 114.540 87.320 114.680 ;
        RECT 75.515 114.495 75.805 114.540 ;
        RECT 85.175 114.495 85.465 114.540 ;
        RECT 87.000 114.480 87.320 114.540 ;
        RECT 90.680 114.680 91.000 114.740 ;
        RECT 96.290 114.680 96.430 114.835 ;
        RECT 90.680 114.540 96.430 114.680 ;
        RECT 90.680 114.480 91.000 114.540 ;
        RECT 103.100 114.480 103.420 114.740 ;
        RECT 105.490 114.680 105.630 114.880 ;
        RECT 112.730 114.835 113.080 115.065 ;
        RECT 112.760 114.820 113.080 114.835 ;
        RECT 116.900 115.020 117.220 115.080 ;
        RECT 118.755 115.020 119.045 115.065 ;
        RECT 116.900 114.880 119.045 115.020 ;
        RECT 124.810 115.020 124.950 115.175 ;
        RECT 125.180 115.160 125.500 115.420 ;
        RECT 125.655 115.360 125.945 115.405 ;
        RECT 126.560 115.360 126.880 115.420 ;
        RECT 130.240 115.360 130.560 115.420 ;
        RECT 125.655 115.220 126.880 115.360 ;
        RECT 125.655 115.175 125.945 115.220 ;
        RECT 126.560 115.160 126.880 115.220 ;
        RECT 127.110 115.220 130.560 115.360 ;
        RECT 127.110 115.020 127.250 115.220 ;
        RECT 130.240 115.160 130.560 115.220 ;
        RECT 124.810 114.880 127.250 115.020 ;
        RECT 127.940 115.020 128.260 115.080 ;
        RECT 131.020 115.020 131.310 115.065 ;
        RECT 127.940 114.880 131.310 115.020 ;
        RECT 116.900 114.820 117.220 114.880 ;
        RECT 118.755 114.835 119.045 114.880 ;
        RECT 127.940 114.820 128.260 114.880 ;
        RECT 131.020 114.835 131.310 114.880 ;
        RECT 114.140 114.680 114.460 114.740 ;
        RECT 105.490 114.540 114.460 114.680 ;
        RECT 114.140 114.480 114.460 114.540 ;
        RECT 118.280 114.680 118.600 114.740 ;
        RECT 119.660 114.680 119.980 114.740 ;
        RECT 118.280 114.540 119.980 114.680 ;
        RECT 118.280 114.480 118.600 114.540 ;
        RECT 119.660 114.480 119.980 114.540 ;
        RECT 127.020 114.480 127.340 114.740 ;
        RECT 136.220 114.680 136.540 114.740 ;
        RECT 136.695 114.680 136.985 114.725 ;
        RECT 136.220 114.540 136.985 114.680 ;
        RECT 136.220 114.480 136.540 114.540 ;
        RECT 136.695 114.495 136.985 114.540 ;
        RECT 13.330 113.860 138.910 114.340 ;
        RECT 26.740 113.660 27.060 113.720 ;
        RECT 27.215 113.660 27.505 113.705 ;
        RECT 26.740 113.520 27.505 113.660 ;
        RECT 26.740 113.460 27.060 113.520 ;
        RECT 27.215 113.475 27.505 113.520 ;
        RECT 29.500 113.460 29.820 113.720 ;
        RECT 30.880 113.460 31.200 113.720 ;
        RECT 41.000 113.660 41.320 113.720 ;
        RECT 41.000 113.520 44.450 113.660 ;
        RECT 41.000 113.460 41.320 113.520 ;
        RECT 25.820 113.320 26.140 113.380 ;
        RECT 27.975 113.320 28.265 113.365 ;
        RECT 25.820 113.180 28.265 113.320 ;
        RECT 25.820 113.120 26.140 113.180 ;
        RECT 27.975 113.135 28.265 113.180 ;
        RECT 29.055 113.320 29.345 113.365 ;
        RECT 30.970 113.320 31.110 113.460 ;
        RECT 29.055 113.180 31.110 113.320 ;
        RECT 35.480 113.320 35.800 113.380 ;
        RECT 44.310 113.320 44.450 113.520 ;
        RECT 44.680 113.460 45.000 113.720 ;
        RECT 47.900 113.460 48.220 113.720 ;
        RECT 53.420 113.460 53.740 113.720 ;
        RECT 61.255 113.660 61.545 113.705 ;
        RECT 65.840 113.660 66.160 113.720 ;
        RECT 61.255 113.520 66.160 113.660 ;
        RECT 61.255 113.475 61.545 113.520 ;
        RECT 65.840 113.460 66.160 113.520 ;
        RECT 68.615 113.660 68.905 113.705 ;
        RECT 90.680 113.660 91.000 113.720 ;
        RECT 68.615 113.520 91.000 113.660 ;
        RECT 68.615 113.475 68.905 113.520 ;
        RECT 90.680 113.460 91.000 113.520 ;
        RECT 91.155 113.660 91.445 113.705 ;
        RECT 91.600 113.660 91.920 113.720 ;
        RECT 91.155 113.520 91.920 113.660 ;
        RECT 91.155 113.475 91.445 113.520 ;
        RECT 91.600 113.460 91.920 113.520 ;
        RECT 103.100 113.660 103.420 113.720 ;
        RECT 111.855 113.660 112.145 113.705 ;
        RECT 112.760 113.660 113.080 113.720 ;
        RECT 117.820 113.660 118.140 113.720 ;
        RECT 129.320 113.660 129.640 113.720 ;
        RECT 103.100 113.520 107.930 113.660 ;
        RECT 103.100 113.460 103.420 113.520 ;
        RECT 52.515 113.320 52.805 113.365 ;
        RECT 69.980 113.320 70.300 113.380 ;
        RECT 85.620 113.320 85.940 113.380 ;
        RECT 35.480 113.180 42.610 113.320 ;
        RECT 44.310 113.180 46.290 113.320 ;
        RECT 29.055 113.135 29.345 113.180 ;
        RECT 35.480 113.120 35.800 113.180 ;
        RECT 19.380 113.025 19.700 113.040 ;
        RECT 19.350 112.980 19.700 113.025 ;
        RECT 19.185 112.840 19.700 112.980 ;
        RECT 19.350 112.795 19.700 112.840 ;
        RECT 30.435 112.980 30.725 113.025 ;
        RECT 30.880 112.980 31.200 113.040 ;
        RECT 30.435 112.840 31.200 112.980 ;
        RECT 30.435 112.795 30.725 112.840 ;
        RECT 19.380 112.780 19.700 112.795 ;
        RECT 30.880 112.780 31.200 112.840 ;
        RECT 41.935 112.795 42.225 113.025 ;
        RECT 42.470 112.980 42.610 113.180 ;
        RECT 42.760 112.980 43.050 113.025 ;
        RECT 42.470 112.840 43.050 112.980 ;
        RECT 42.760 112.795 43.050 112.840 ;
        RECT 17.540 112.640 17.860 112.700 ;
        RECT 18.015 112.640 18.305 112.685 ;
        RECT 17.540 112.500 18.305 112.640 ;
        RECT 17.540 112.440 17.860 112.500 ;
        RECT 18.015 112.455 18.305 112.500 ;
        RECT 18.895 112.640 19.185 112.685 ;
        RECT 20.085 112.640 20.375 112.685 ;
        RECT 22.605 112.640 22.895 112.685 ;
        RECT 18.895 112.500 22.895 112.640 ;
        RECT 18.895 112.455 19.185 112.500 ;
        RECT 20.085 112.455 20.375 112.500 ;
        RECT 22.605 112.455 22.895 112.500 ;
        RECT 24.900 112.640 25.220 112.700 ;
        RECT 31.355 112.640 31.645 112.685 ;
        RECT 24.900 112.500 31.645 112.640 ;
        RECT 24.900 112.440 25.220 112.500 ;
        RECT 31.355 112.455 31.645 112.500 ;
        RECT 18.500 112.300 18.790 112.345 ;
        RECT 20.600 112.300 20.890 112.345 ;
        RECT 22.170 112.300 22.460 112.345 ;
        RECT 18.500 112.160 22.460 112.300 ;
        RECT 18.500 112.115 18.790 112.160 ;
        RECT 20.600 112.115 20.890 112.160 ;
        RECT 22.170 112.115 22.460 112.160 ;
        RECT 23.980 111.960 24.300 112.020 ;
        RECT 24.915 111.960 25.205 112.005 ;
        RECT 23.980 111.820 25.205 111.960 ;
        RECT 23.980 111.760 24.300 111.820 ;
        RECT 24.915 111.775 25.205 111.820 ;
        RECT 25.360 111.960 25.680 112.020 ;
        RECT 28.135 111.960 28.425 112.005 ;
        RECT 25.360 111.820 28.425 111.960 ;
        RECT 42.010 111.960 42.150 112.795 ;
        RECT 43.300 112.780 43.620 113.040 ;
        RECT 43.775 112.980 44.065 113.025 ;
        RECT 44.220 112.980 44.540 113.040 ;
        RECT 46.150 113.025 46.290 113.180 ;
        RECT 47.070 113.180 52.805 113.320 ;
        RECT 47.070 113.040 47.210 113.180 ;
        RECT 52.515 113.135 52.805 113.180 ;
        RECT 62.710 113.180 70.300 113.320 ;
        RECT 43.775 112.840 44.540 112.980 ;
        RECT 43.775 112.795 44.065 112.840 ;
        RECT 44.220 112.780 44.540 112.840 ;
        RECT 44.695 112.980 44.985 113.025 ;
        RECT 45.155 112.980 45.445 113.025 ;
        RECT 44.695 112.840 45.445 112.980 ;
        RECT 44.695 112.795 44.985 112.840 ;
        RECT 45.155 112.795 45.445 112.840 ;
        RECT 46.075 112.795 46.365 113.025 ;
        RECT 46.150 112.640 46.290 112.795 ;
        RECT 46.980 112.780 47.300 113.040 ;
        RECT 47.440 112.780 47.760 113.040 ;
        RECT 48.360 112.980 48.680 113.040 ;
        RECT 48.835 112.980 49.125 113.025 ;
        RECT 48.360 112.840 49.125 112.980 ;
        RECT 48.360 112.780 48.680 112.840 ;
        RECT 48.835 112.795 49.125 112.840 ;
        RECT 50.200 112.980 50.520 113.040 ;
        RECT 51.135 112.980 51.425 113.025 ;
        RECT 50.200 112.840 51.425 112.980 ;
        RECT 50.200 112.780 50.520 112.840 ;
        RECT 51.135 112.795 51.425 112.840 ;
        RECT 51.595 112.795 51.885 113.025 ;
        RECT 49.295 112.640 49.585 112.685 ;
        RECT 46.150 112.500 49.585 112.640 ;
        RECT 49.295 112.455 49.585 112.500 ;
        RECT 47.440 112.300 47.760 112.360 ;
        RECT 51.670 112.300 51.810 112.795 ;
        RECT 59.860 112.780 60.180 113.040 ;
        RECT 60.335 112.980 60.625 113.025 ;
        RECT 62.160 112.980 62.480 113.040 ;
        RECT 62.710 113.025 62.850 113.180 ;
        RECT 69.980 113.120 70.300 113.180 ;
        RECT 83.410 113.180 85.940 113.320 ;
        RECT 60.335 112.840 62.480 112.980 ;
        RECT 60.335 112.795 60.625 112.840 ;
        RECT 62.160 112.780 62.480 112.840 ;
        RECT 62.635 112.795 62.925 113.025 ;
        RECT 65.380 112.780 65.700 113.040 ;
        RECT 66.300 112.780 66.620 113.040 ;
        RECT 71.360 112.780 71.680 113.040 ;
        RECT 83.410 113.025 83.550 113.180 ;
        RECT 85.620 113.120 85.940 113.180 ;
        RECT 101.260 113.320 101.580 113.380 ;
        RECT 105.875 113.320 106.165 113.365 ;
        RECT 101.260 113.180 104.250 113.320 ;
        RECT 101.260 113.120 101.580 113.180 ;
        RECT 104.110 113.040 104.250 113.180 ;
        RECT 104.570 113.180 106.165 113.320 ;
        RECT 84.700 113.025 85.020 113.040 ;
        RECT 83.335 112.795 83.625 113.025 ;
        RECT 84.670 112.795 85.020 113.025 ;
        RECT 84.700 112.780 85.020 112.795 ;
        RECT 92.060 112.780 92.380 113.040 ;
        RECT 92.520 112.780 92.840 113.040 ;
        RECT 93.455 112.795 93.745 113.025 ;
        RECT 93.915 112.795 94.205 113.025 ;
        RECT 61.255 112.455 61.545 112.685 ;
        RECT 63.095 112.640 63.385 112.685 ;
        RECT 67.220 112.640 67.540 112.700 ;
        RECT 67.695 112.640 67.985 112.685 ;
        RECT 63.095 112.500 66.070 112.640 ;
        RECT 63.095 112.455 63.385 112.500 ;
        RECT 47.440 112.160 51.810 112.300 ;
        RECT 47.440 112.100 47.760 112.160 ;
        RECT 50.200 111.960 50.520 112.020 ;
        RECT 42.010 111.820 50.520 111.960 ;
        RECT 25.360 111.760 25.680 111.820 ;
        RECT 28.135 111.775 28.425 111.820 ;
        RECT 50.200 111.760 50.520 111.820 ;
        RECT 50.675 111.960 50.965 112.005 ;
        RECT 51.670 111.960 51.810 112.160 ;
        RECT 50.675 111.820 51.810 111.960 ;
        RECT 61.330 111.960 61.470 112.455 ;
        RECT 65.930 112.360 66.070 112.500 ;
        RECT 67.220 112.500 67.985 112.640 ;
        RECT 67.220 112.440 67.540 112.500 ;
        RECT 67.695 112.455 67.985 112.500 ;
        RECT 68.140 112.640 68.460 112.700 ;
        RECT 69.535 112.640 69.825 112.685 ;
        RECT 68.140 112.500 69.825 112.640 ;
        RECT 68.140 112.440 68.460 112.500 ;
        RECT 69.535 112.455 69.825 112.500 ;
        RECT 69.980 112.440 70.300 112.700 ;
        RECT 70.915 112.640 71.205 112.685 ;
        RECT 75.040 112.640 75.360 112.700 ;
        RECT 70.915 112.500 75.360 112.640 ;
        RECT 70.915 112.455 71.205 112.500 ;
        RECT 75.040 112.440 75.360 112.500 ;
        RECT 84.215 112.640 84.505 112.685 ;
        RECT 85.405 112.640 85.695 112.685 ;
        RECT 87.925 112.640 88.215 112.685 ;
        RECT 84.215 112.500 88.215 112.640 ;
        RECT 84.215 112.455 84.505 112.500 ;
        RECT 85.405 112.455 85.695 112.500 ;
        RECT 87.925 112.455 88.215 112.500 ;
        RECT 64.460 112.100 64.780 112.360 ;
        RECT 65.840 112.100 66.160 112.360 ;
        RECT 70.455 112.300 70.745 112.345 ;
        RECT 67.310 112.160 70.745 112.300 ;
        RECT 67.310 111.960 67.450 112.160 ;
        RECT 70.455 112.115 70.745 112.160 ;
        RECT 83.820 112.300 84.110 112.345 ;
        RECT 85.920 112.300 86.210 112.345 ;
        RECT 87.490 112.300 87.780 112.345 ;
        RECT 83.820 112.160 87.780 112.300 ;
        RECT 93.530 112.300 93.670 112.795 ;
        RECT 93.990 112.640 94.130 112.795 ;
        RECT 103.560 112.780 103.880 113.040 ;
        RECT 104.020 112.780 104.340 113.040 ;
        RECT 104.570 113.025 104.710 113.180 ;
        RECT 105.875 113.135 106.165 113.180 ;
        RECT 104.495 112.795 104.785 113.025 ;
        RECT 104.940 112.980 105.260 113.040 ;
        RECT 105.415 112.980 105.705 113.025 ;
        RECT 104.940 112.840 105.705 112.980 ;
        RECT 104.940 112.780 105.260 112.840 ;
        RECT 105.415 112.795 105.705 112.840 ;
        RECT 106.780 112.780 107.100 113.040 ;
        RECT 107.790 113.025 107.930 113.520 ;
        RECT 111.855 113.520 113.080 113.660 ;
        RECT 111.855 113.475 112.145 113.520 ;
        RECT 112.760 113.460 113.080 113.520 ;
        RECT 113.770 113.520 118.140 113.660 ;
        RECT 110.000 113.320 110.320 113.380 ;
        RECT 110.000 113.180 113.450 113.320 ;
        RECT 110.000 113.120 110.320 113.180 ;
        RECT 111.930 113.040 112.070 113.180 ;
        RECT 107.715 112.980 108.005 113.025 ;
        RECT 109.555 112.980 109.845 113.025 ;
        RECT 107.715 112.840 109.845 112.980 ;
        RECT 107.715 112.795 108.005 112.840 ;
        RECT 109.555 112.795 109.845 112.840 ;
        RECT 93.990 112.500 108.390 112.640 ;
        RECT 107.700 112.300 108.020 112.360 ;
        RECT 93.530 112.160 108.020 112.300 ;
        RECT 83.820 112.115 84.110 112.160 ;
        RECT 85.920 112.115 86.210 112.160 ;
        RECT 87.490 112.115 87.780 112.160 ;
        RECT 107.700 112.100 108.020 112.160 ;
        RECT 61.330 111.820 67.450 111.960 ;
        RECT 50.675 111.775 50.965 111.820 ;
        RECT 67.680 111.760 68.000 112.020 ;
        RECT 90.235 111.960 90.525 112.005 ;
        RECT 92.520 111.960 92.840 112.020 ;
        RECT 90.235 111.820 92.840 111.960 ;
        RECT 90.235 111.775 90.525 111.820 ;
        RECT 92.520 111.760 92.840 111.820 ;
        RECT 102.195 111.960 102.485 112.005 ;
        RECT 104.480 111.960 104.800 112.020 ;
        RECT 102.195 111.820 104.800 111.960 ;
        RECT 108.250 111.960 108.390 112.500 ;
        RECT 109.630 112.300 109.770 112.795 ;
        RECT 110.460 112.780 110.780 113.040 ;
        RECT 111.840 112.780 112.160 113.040 ;
        RECT 113.310 113.025 113.450 113.180 ;
        RECT 113.770 113.025 113.910 113.520 ;
        RECT 117.820 113.460 118.140 113.520 ;
        RECT 125.730 113.520 129.640 113.660 ;
        RECT 116.900 113.120 117.220 113.380 ;
        RECT 124.260 113.320 124.580 113.380 ;
        RECT 125.730 113.320 125.870 113.520 ;
        RECT 129.320 113.460 129.640 113.520 ;
        RECT 133.000 113.660 133.320 113.720 ;
        RECT 134.395 113.660 134.685 113.705 ;
        RECT 135.760 113.660 136.080 113.720 ;
        RECT 133.000 113.520 136.080 113.660 ;
        RECT 133.000 113.460 133.320 113.520 ;
        RECT 134.395 113.475 134.685 113.520 ;
        RECT 135.760 113.460 136.080 113.520 ;
        RECT 136.695 113.660 136.985 113.705 ;
        RECT 138.520 113.660 138.840 113.720 ;
        RECT 136.695 113.520 138.840 113.660 ;
        RECT 136.695 113.475 136.985 113.520 ;
        RECT 138.520 113.460 138.840 113.520 ;
        RECT 124.260 113.180 125.870 113.320 ;
        RECT 124.260 113.120 124.580 113.180 ;
        RECT 113.235 112.795 113.525 113.025 ;
        RECT 113.695 112.795 113.985 113.025 ;
        RECT 114.155 112.795 114.445 113.025 ;
        RECT 115.060 112.980 115.380 113.040 ;
        RECT 123.815 112.980 124.105 113.025 ;
        RECT 115.060 112.840 124.105 112.980 ;
        RECT 112.760 112.640 113.080 112.700 ;
        RECT 113.770 112.640 113.910 112.795 ;
        RECT 112.760 112.500 113.910 112.640 ;
        RECT 114.230 112.640 114.370 112.795 ;
        RECT 115.060 112.780 115.380 112.840 ;
        RECT 123.815 112.795 124.105 112.840 ;
        RECT 124.735 112.795 125.025 113.025 ;
        RECT 120.120 112.640 120.440 112.700 ;
        RECT 114.230 112.500 120.440 112.640 ;
        RECT 112.760 112.440 113.080 112.500 ;
        RECT 120.120 112.440 120.440 112.500 ;
        RECT 121.040 112.440 121.360 112.700 ;
        RECT 118.740 112.300 119.060 112.360 ;
        RECT 109.630 112.160 119.060 112.300 ;
        RECT 124.810 112.300 124.950 112.795 ;
        RECT 125.180 112.780 125.500 113.040 ;
        RECT 125.730 113.025 125.870 113.180 ;
        RECT 127.020 113.320 127.340 113.380 ;
        RECT 128.720 113.320 129.010 113.365 ;
        RECT 127.020 113.180 129.010 113.320 ;
        RECT 127.020 113.120 127.340 113.180 ;
        RECT 128.720 113.135 129.010 113.180 ;
        RECT 125.655 112.795 125.945 113.025 ;
        RECT 127.480 112.780 127.800 113.040 ;
        RECT 127.940 112.780 128.260 113.040 ;
        RECT 131.160 112.980 131.480 113.040 ;
        RECT 135.775 112.980 136.065 113.025 ;
        RECT 136.220 112.980 136.540 113.040 ;
        RECT 131.160 112.840 136.540 112.980 ;
        RECT 131.160 112.780 131.480 112.840 ;
        RECT 135.775 112.795 136.065 112.840 ;
        RECT 136.220 112.780 136.540 112.840 ;
        RECT 127.035 112.640 127.325 112.685 ;
        RECT 128.030 112.640 128.170 112.780 ;
        RECT 127.035 112.500 128.170 112.640 ;
        RECT 128.375 112.640 128.665 112.685 ;
        RECT 129.565 112.640 129.855 112.685 ;
        RECT 132.085 112.640 132.375 112.685 ;
        RECT 128.375 112.500 132.375 112.640 ;
        RECT 127.035 112.455 127.325 112.500 ;
        RECT 128.375 112.455 128.665 112.500 ;
        RECT 129.565 112.455 129.855 112.500 ;
        RECT 132.085 112.455 132.375 112.500 ;
        RECT 125.180 112.300 125.500 112.360 ;
        RECT 124.810 112.160 125.500 112.300 ;
        RECT 118.740 112.100 119.060 112.160 ;
        RECT 125.180 112.100 125.500 112.160 ;
        RECT 127.980 112.300 128.270 112.345 ;
        RECT 130.080 112.300 130.370 112.345 ;
        RECT 131.650 112.300 131.940 112.345 ;
        RECT 127.980 112.160 131.940 112.300 ;
        RECT 127.980 112.115 128.270 112.160 ;
        RECT 130.080 112.115 130.370 112.160 ;
        RECT 131.650 112.115 131.940 112.160 ;
        RECT 110.920 111.960 111.240 112.020 ;
        RECT 108.250 111.820 111.240 111.960 ;
        RECT 102.195 111.775 102.485 111.820 ;
        RECT 104.480 111.760 104.800 111.820 ;
        RECT 110.920 111.760 111.240 111.820 ;
        RECT 111.395 111.960 111.685 112.005 ;
        RECT 112.300 111.960 112.620 112.020 ;
        RECT 111.395 111.820 112.620 111.960 ;
        RECT 111.395 111.775 111.685 111.820 ;
        RECT 112.300 111.760 112.620 111.820 ;
        RECT 13.330 111.140 138.910 111.620 ;
        RECT 44.695 110.940 44.985 110.985 ;
        RECT 46.980 110.940 47.300 111.000 ;
        RECT 61.715 110.940 62.005 110.985 ;
        RECT 64.920 110.940 65.240 111.000 ;
        RECT 67.680 110.940 68.000 111.000 ;
        RECT 44.695 110.800 51.810 110.940 ;
        RECT 44.695 110.755 44.985 110.800 ;
        RECT 46.980 110.740 47.300 110.800 ;
        RECT 18.040 110.600 18.330 110.645 ;
        RECT 20.140 110.600 20.430 110.645 ;
        RECT 21.710 110.600 22.000 110.645 ;
        RECT 18.040 110.460 22.000 110.600 ;
        RECT 18.040 110.415 18.330 110.460 ;
        RECT 20.140 110.415 20.430 110.460 ;
        RECT 21.710 110.415 22.000 110.460 ;
        RECT 47.440 110.600 47.730 110.645 ;
        RECT 49.010 110.600 49.300 110.645 ;
        RECT 51.110 110.600 51.400 110.645 ;
        RECT 47.440 110.460 51.400 110.600 ;
        RECT 47.440 110.415 47.730 110.460 ;
        RECT 49.010 110.415 49.300 110.460 ;
        RECT 51.110 110.415 51.400 110.460 ;
        RECT 17.540 110.060 17.860 110.320 ;
        RECT 18.435 110.260 18.725 110.305 ;
        RECT 19.625 110.260 19.915 110.305 ;
        RECT 22.145 110.260 22.435 110.305 ;
        RECT 18.435 110.120 22.435 110.260 ;
        RECT 18.435 110.075 18.725 110.120 ;
        RECT 19.625 110.075 19.915 110.120 ;
        RECT 22.145 110.075 22.435 110.120 ;
        RECT 25.820 110.260 26.140 110.320 ;
        RECT 29.515 110.260 29.805 110.305 ;
        RECT 25.820 110.120 29.805 110.260 ;
        RECT 25.820 110.060 26.140 110.120 ;
        RECT 29.515 110.075 29.805 110.120 ;
        RECT 47.005 110.260 47.295 110.305 ;
        RECT 49.525 110.260 49.815 110.305 ;
        RECT 50.715 110.260 51.005 110.305 ;
        RECT 47.005 110.120 51.005 110.260 ;
        RECT 51.670 110.260 51.810 110.800 ;
        RECT 61.715 110.800 68.000 110.940 ;
        RECT 61.715 110.755 62.005 110.800 ;
        RECT 64.920 110.740 65.240 110.800 ;
        RECT 67.680 110.740 68.000 110.800 ;
        RECT 69.995 110.940 70.285 110.985 ;
        RECT 70.900 110.940 71.220 111.000 ;
        RECT 69.995 110.800 71.220 110.940 ;
        RECT 69.995 110.755 70.285 110.800 ;
        RECT 70.900 110.740 71.220 110.800 ;
        RECT 79.180 110.940 79.500 111.000 ;
        RECT 82.415 110.940 82.705 110.985 ;
        RECT 79.180 110.800 82.705 110.940 ;
        RECT 79.180 110.740 79.500 110.800 ;
        RECT 82.415 110.755 82.705 110.800 ;
        RECT 88.380 110.940 88.700 111.000 ;
        RECT 103.560 110.940 103.880 111.000 ;
        RECT 104.940 110.940 105.260 111.000 ;
        RECT 88.380 110.800 103.880 110.940 ;
        RECT 88.380 110.740 88.700 110.800 ;
        RECT 103.560 110.740 103.880 110.800 ;
        RECT 104.110 110.800 111.610 110.940 ;
        RECT 63.080 110.600 63.400 110.660 ;
        RECT 62.250 110.460 63.400 110.600 ;
        RECT 52.515 110.260 52.805 110.305 ;
        RECT 51.670 110.120 52.805 110.260 ;
        RECT 47.005 110.075 47.295 110.120 ;
        RECT 49.525 110.075 49.815 110.120 ;
        RECT 50.715 110.075 51.005 110.120 ;
        RECT 52.515 110.075 52.805 110.120 ;
        RECT 23.980 109.920 24.300 109.980 ;
        RECT 27.200 109.920 27.520 109.980 ;
        RECT 27.675 109.920 27.965 109.965 ;
        RECT 23.980 109.780 27.965 109.920 ;
        RECT 23.980 109.720 24.300 109.780 ;
        RECT 27.200 109.720 27.520 109.780 ;
        RECT 27.675 109.735 27.965 109.780 ;
        RECT 28.580 109.920 28.900 109.980 ;
        RECT 30.880 109.920 31.200 109.980 ;
        RECT 28.580 109.780 31.200 109.920 ;
        RECT 28.580 109.720 28.900 109.780 ;
        RECT 30.880 109.720 31.200 109.780 ;
        RECT 36.860 109.920 37.180 109.980 ;
        RECT 43.315 109.920 43.605 109.965 ;
        RECT 36.860 109.780 43.605 109.920 ;
        RECT 36.860 109.720 37.180 109.780 ;
        RECT 43.315 109.735 43.605 109.780 ;
        RECT 51.580 109.720 51.900 109.980 ;
        RECT 55.735 109.920 56.025 109.965 ;
        RECT 56.195 109.920 56.485 109.965 ;
        RECT 55.735 109.780 56.485 109.920 ;
        RECT 55.735 109.735 56.025 109.780 ;
        RECT 56.195 109.735 56.485 109.780 ;
        RECT 61.255 109.920 61.545 109.965 ;
        RECT 62.250 109.920 62.390 110.460 ;
        RECT 63.080 110.400 63.400 110.460 ;
        RECT 63.580 110.600 63.870 110.645 ;
        RECT 65.680 110.600 65.970 110.645 ;
        RECT 67.250 110.600 67.540 110.645 ;
        RECT 97.595 110.600 97.885 110.645 ;
        RECT 100.800 110.600 101.120 110.660 ;
        RECT 63.580 110.460 67.540 110.600 ;
        RECT 63.580 110.415 63.870 110.460 ;
        RECT 65.680 110.415 65.970 110.460 ;
        RECT 67.250 110.415 67.540 110.460 ;
        RECT 82.950 110.460 92.750 110.600 ;
        RECT 62.620 110.060 62.940 110.320 ;
        RECT 63.170 110.260 63.310 110.400 ;
        RECT 63.975 110.260 64.265 110.305 ;
        RECT 65.165 110.260 65.455 110.305 ;
        RECT 67.685 110.260 67.975 110.305 ;
        RECT 63.170 110.120 63.770 110.260 ;
        RECT 61.255 109.780 62.390 109.920 ;
        RECT 61.255 109.735 61.545 109.780 ;
        RECT 63.095 109.735 63.385 109.965 ;
        RECT 18.890 109.580 19.180 109.625 ;
        RECT 19.380 109.580 19.700 109.640 ;
        RECT 18.890 109.440 19.700 109.580 ;
        RECT 18.890 109.395 19.180 109.440 ;
        RECT 19.380 109.380 19.700 109.440 ;
        RECT 23.520 109.580 23.840 109.640 ;
        RECT 26.755 109.580 27.045 109.625 ;
        RECT 28.135 109.580 28.425 109.625 ;
        RECT 23.520 109.440 27.045 109.580 ;
        RECT 23.520 109.380 23.840 109.440 ;
        RECT 26.755 109.395 27.045 109.440 ;
        RECT 27.290 109.440 28.425 109.580 ;
        RECT 18.460 109.240 18.780 109.300 ;
        RECT 24.455 109.240 24.745 109.285 ;
        RECT 26.280 109.240 26.600 109.300 ;
        RECT 27.290 109.240 27.430 109.440 ;
        RECT 28.135 109.395 28.425 109.440 ;
        RECT 50.370 109.580 50.660 109.625 ;
        RECT 52.040 109.580 52.360 109.640 ;
        RECT 50.370 109.440 52.360 109.580 ;
        RECT 50.370 109.395 50.660 109.440 ;
        RECT 52.040 109.380 52.360 109.440 ;
        RECT 60.320 109.580 60.640 109.640 ;
        RECT 63.170 109.580 63.310 109.735 ;
        RECT 60.320 109.440 63.310 109.580 ;
        RECT 63.630 109.580 63.770 110.120 ;
        RECT 63.975 110.120 67.975 110.260 ;
        RECT 63.975 110.075 64.265 110.120 ;
        RECT 65.165 110.075 65.455 110.120 ;
        RECT 67.685 110.075 67.975 110.120 ;
        RECT 64.460 109.965 64.780 109.980 ;
        RECT 64.430 109.920 64.780 109.965 ;
        RECT 64.265 109.780 64.780 109.920 ;
        RECT 64.430 109.735 64.780 109.780 ;
        RECT 64.460 109.720 64.780 109.735 ;
        RECT 76.880 109.920 77.200 109.980 ;
        RECT 78.275 109.920 78.565 109.965 ;
        RECT 81.020 109.920 81.340 109.980 ;
        RECT 82.950 109.920 83.090 110.460 ;
        RECT 92.060 110.260 92.380 110.320 ;
        RECT 83.410 110.120 92.380 110.260 ;
        RECT 92.610 110.260 92.750 110.460 ;
        RECT 97.595 110.460 101.120 110.600 ;
        RECT 97.595 110.415 97.885 110.460 ;
        RECT 100.800 110.400 101.120 110.460 ;
        RECT 102.180 110.260 102.500 110.320 ;
        RECT 104.110 110.260 104.250 110.800 ;
        RECT 104.940 110.740 105.260 110.800 ;
        RECT 104.520 110.600 104.810 110.645 ;
        RECT 106.620 110.600 106.910 110.645 ;
        RECT 108.190 110.600 108.480 110.645 ;
        RECT 104.520 110.460 108.480 110.600 ;
        RECT 104.520 110.415 104.810 110.460 ;
        RECT 106.620 110.415 106.910 110.460 ;
        RECT 108.190 110.415 108.480 110.460 ;
        RECT 92.610 110.120 93.670 110.260 ;
        RECT 83.410 109.980 83.550 110.120 ;
        RECT 92.060 110.060 92.380 110.120 ;
        RECT 76.880 109.780 83.090 109.920 ;
        RECT 76.880 109.720 77.200 109.780 ;
        RECT 78.275 109.735 78.565 109.780 ;
        RECT 81.020 109.720 81.340 109.780 ;
        RECT 83.320 109.720 83.640 109.980 ;
        RECT 83.795 109.735 84.085 109.965 ;
        RECT 84.715 109.735 85.005 109.965 ;
        RECT 67.220 109.580 67.540 109.640 ;
        RECT 63.630 109.440 67.540 109.580 ;
        RECT 60.320 109.380 60.640 109.440 ;
        RECT 67.220 109.380 67.540 109.440 ;
        RECT 79.180 109.580 79.500 109.640 ;
        RECT 83.870 109.580 84.010 109.735 ;
        RECT 79.180 109.440 84.010 109.580 ;
        RECT 79.180 109.380 79.500 109.440 ;
        RECT 18.460 109.100 27.430 109.240 ;
        RECT 30.880 109.240 31.200 109.300 ;
        RECT 43.775 109.240 44.065 109.285 ;
        RECT 46.520 109.240 46.840 109.300 ;
        RECT 30.880 109.100 46.840 109.240 ;
        RECT 18.460 109.040 18.780 109.100 ;
        RECT 24.455 109.055 24.745 109.100 ;
        RECT 26.280 109.040 26.600 109.100 ;
        RECT 30.880 109.040 31.200 109.100 ;
        RECT 43.775 109.055 44.065 109.100 ;
        RECT 46.520 109.040 46.840 109.100 ;
        RECT 48.360 109.240 48.680 109.300 ;
        RECT 56.655 109.240 56.945 109.285 ;
        RECT 48.360 109.100 56.945 109.240 ;
        RECT 48.360 109.040 48.680 109.100 ;
        RECT 56.655 109.055 56.945 109.100 ;
        RECT 62.635 109.240 62.925 109.285 ;
        RECT 64.460 109.240 64.780 109.300 ;
        RECT 62.635 109.100 64.780 109.240 ;
        RECT 62.635 109.055 62.925 109.100 ;
        RECT 64.460 109.040 64.780 109.100 ;
        RECT 80.115 109.240 80.405 109.285 ;
        RECT 80.560 109.240 80.880 109.300 ;
        RECT 80.115 109.100 80.880 109.240 ;
        RECT 84.790 109.240 84.930 109.735 ;
        RECT 85.160 109.720 85.480 109.980 ;
        RECT 91.140 109.720 91.460 109.980 ;
        RECT 93.530 109.965 93.670 110.120 ;
        RECT 99.925 110.120 104.250 110.260 ;
        RECT 104.915 110.260 105.205 110.305 ;
        RECT 106.105 110.260 106.395 110.305 ;
        RECT 108.625 110.260 108.915 110.305 ;
        RECT 104.915 110.120 108.915 110.260 ;
        RECT 93.455 109.920 93.745 109.965 ;
        RECT 98.040 109.920 98.360 109.980 ;
        RECT 99.925 109.965 100.065 110.120 ;
        RECT 102.180 110.060 102.500 110.120 ;
        RECT 104.915 110.075 105.205 110.120 ;
        RECT 106.105 110.075 106.395 110.120 ;
        RECT 108.625 110.075 108.915 110.120 ;
        RECT 111.470 110.260 111.610 110.800 ;
        RECT 115.520 110.740 115.840 111.000 ;
        RECT 128.860 110.940 129.180 111.000 ;
        RECT 130.700 110.940 131.020 111.000 ;
        RECT 119.750 110.800 131.020 110.940 ;
        RECT 115.060 110.260 115.380 110.320 ;
        RECT 111.470 110.120 115.380 110.260 ;
        RECT 115.610 110.260 115.750 110.740 ;
        RECT 119.750 110.260 119.890 110.800 ;
        RECT 128.860 110.740 129.180 110.800 ;
        RECT 130.700 110.740 131.020 110.800 ;
        RECT 131.160 110.600 131.480 110.660 ;
        RECT 126.190 110.460 131.480 110.600 ;
        RECT 115.610 110.120 119.890 110.260 ;
        RECT 93.455 109.780 98.360 109.920 ;
        RECT 93.455 109.735 93.745 109.780 ;
        RECT 98.040 109.720 98.360 109.780 ;
        RECT 99.835 109.735 100.125 109.965 ;
        RECT 100.800 109.720 101.120 109.980 ;
        RECT 101.260 109.720 101.580 109.980 ;
        RECT 101.720 109.720 102.040 109.980 ;
        RECT 103.560 109.920 103.880 109.980 ;
        RECT 111.470 109.965 111.610 110.120 ;
        RECT 115.060 110.060 115.380 110.120 ;
        RECT 104.035 109.920 104.325 109.965 ;
        RECT 103.560 109.780 104.325 109.920 ;
        RECT 103.560 109.720 103.880 109.780 ;
        RECT 104.035 109.735 104.325 109.780 ;
        RECT 111.395 109.735 111.685 109.965 ;
        RECT 112.300 109.720 112.620 109.980 ;
        RECT 112.760 109.720 113.080 109.980 ;
        RECT 113.235 109.735 113.525 109.965 ;
        RECT 114.140 109.920 114.460 109.980 ;
        RECT 119.750 109.965 119.890 110.120 ;
        RECT 120.120 110.260 120.440 110.320 ;
        RECT 121.055 110.260 121.345 110.305 ;
        RECT 120.120 110.120 121.345 110.260 ;
        RECT 120.120 110.060 120.440 110.120 ;
        RECT 121.055 110.075 121.345 110.120 ;
        RECT 125.180 110.060 125.500 110.320 ;
        RECT 118.755 109.920 119.045 109.965 ;
        RECT 114.140 109.780 119.045 109.920 ;
        RECT 85.620 109.580 85.940 109.640 ;
        RECT 87.015 109.580 87.305 109.625 ;
        RECT 85.620 109.440 87.305 109.580 ;
        RECT 85.620 109.380 85.940 109.440 ;
        RECT 87.015 109.395 87.305 109.440 ;
        RECT 92.060 109.580 92.380 109.640 ;
        RECT 92.535 109.580 92.825 109.625 ;
        RECT 92.060 109.440 92.825 109.580 ;
        RECT 92.060 109.380 92.380 109.440 ;
        RECT 92.535 109.395 92.825 109.440 ;
        RECT 98.515 109.395 98.805 109.625 ;
        RECT 99.435 109.580 99.725 109.625 ;
        RECT 102.640 109.580 102.960 109.640 ;
        RECT 99.435 109.440 102.960 109.580 ;
        RECT 99.435 109.395 99.725 109.440 ;
        RECT 87.460 109.240 87.780 109.300 ;
        RECT 84.790 109.100 87.780 109.240 ;
        RECT 80.115 109.055 80.405 109.100 ;
        RECT 80.560 109.040 80.880 109.100 ;
        RECT 87.460 109.040 87.780 109.100 ;
        RECT 87.920 109.240 88.240 109.300 ;
        RECT 91.615 109.240 91.905 109.285 ;
        RECT 87.920 109.100 91.905 109.240 ;
        RECT 87.920 109.040 88.240 109.100 ;
        RECT 91.615 109.055 91.905 109.100 ;
        RECT 97.580 109.240 97.900 109.300 ;
        RECT 98.590 109.240 98.730 109.395 ;
        RECT 102.640 109.380 102.960 109.440 ;
        RECT 103.115 109.580 103.405 109.625 ;
        RECT 105.260 109.580 105.550 109.625 ;
        RECT 103.115 109.440 105.550 109.580 ;
        RECT 113.310 109.580 113.450 109.735 ;
        RECT 114.140 109.720 114.460 109.780 ;
        RECT 118.755 109.735 119.045 109.780 ;
        RECT 119.675 109.735 119.965 109.965 ;
        RECT 120.595 109.920 120.885 109.965 ;
        RECT 122.420 109.920 122.740 109.980 ;
        RECT 126.190 109.965 126.330 110.460 ;
        RECT 131.160 110.400 131.480 110.460 ;
        RECT 120.595 109.780 125.870 109.920 ;
        RECT 120.595 109.735 120.885 109.780 ;
        RECT 122.420 109.720 122.740 109.780 ;
        RECT 116.440 109.580 116.760 109.640 ;
        RECT 113.310 109.440 116.760 109.580 ;
        RECT 103.115 109.395 103.405 109.440 ;
        RECT 105.260 109.395 105.550 109.440 ;
        RECT 116.440 109.380 116.760 109.440 ;
        RECT 118.280 109.580 118.600 109.640 ;
        RECT 121.975 109.580 122.265 109.625 ;
        RECT 118.280 109.440 122.265 109.580 ;
        RECT 118.280 109.380 118.600 109.440 ;
        RECT 121.975 109.395 122.265 109.440 ;
        RECT 110.935 109.240 111.225 109.285 ;
        RECT 111.380 109.240 111.700 109.300 ;
        RECT 97.580 109.100 111.700 109.240 ;
        RECT 97.580 109.040 97.900 109.100 ;
        RECT 110.935 109.055 111.225 109.100 ;
        RECT 111.380 109.040 111.700 109.100 ;
        RECT 114.600 109.040 114.920 109.300 ;
        RECT 122.050 109.240 122.190 109.395 ;
        RECT 122.880 109.380 123.200 109.640 ;
        RECT 125.730 109.580 125.870 109.780 ;
        RECT 126.115 109.735 126.405 109.965 ;
        RECT 130.700 109.720 131.020 109.980 ;
        RECT 131.160 109.720 131.480 109.980 ;
        RECT 132.540 109.720 132.860 109.980 ;
        RECT 133.935 109.735 134.225 109.965 ;
        RECT 127.035 109.580 127.325 109.625 ;
        RECT 125.730 109.440 127.325 109.580 ;
        RECT 127.035 109.395 127.325 109.440 ;
        RECT 127.570 109.440 130.470 109.580 ;
        RECT 127.570 109.240 127.710 109.440 ;
        RECT 122.050 109.100 127.710 109.240 ;
        RECT 129.780 109.040 130.100 109.300 ;
        RECT 130.330 109.240 130.470 109.440 ;
        RECT 131.620 109.380 131.940 109.640 ;
        RECT 134.010 109.240 134.150 109.735 ;
        RECT 135.760 109.720 136.080 109.980 ;
        RECT 130.330 109.100 134.150 109.240 ;
        RECT 134.840 109.040 135.160 109.300 ;
        RECT 136.680 109.040 137.000 109.300 ;
        RECT 13.330 108.420 138.910 108.900 ;
        RECT 18.935 108.035 19.225 108.265 ;
        RECT 18.460 107.680 18.780 107.940 ;
        RECT 19.010 107.880 19.150 108.035 ;
        RECT 19.380 108.020 19.700 108.280 ;
        RECT 21.680 108.020 22.000 108.280 ;
        RECT 27.215 108.220 27.505 108.265 ;
        RECT 28.120 108.220 28.440 108.280 ;
        RECT 22.690 108.080 28.440 108.220 ;
        RECT 20.155 107.880 20.445 107.925 ;
        RECT 19.010 107.740 20.445 107.880 ;
        RECT 20.155 107.695 20.445 107.740 ;
        RECT 21.235 107.880 21.525 107.925 ;
        RECT 22.690 107.880 22.830 108.080 ;
        RECT 27.215 108.035 27.505 108.080 ;
        RECT 28.120 108.020 28.440 108.080 ;
        RECT 37.795 108.220 38.085 108.265 ;
        RECT 40.080 108.220 40.400 108.280 ;
        RECT 37.795 108.080 40.400 108.220 ;
        RECT 37.795 108.035 38.085 108.080 ;
        RECT 40.080 108.020 40.400 108.080 ;
        RECT 40.540 108.020 40.860 108.280 ;
        RECT 48.360 108.020 48.680 108.280 ;
        RECT 52.040 108.220 52.360 108.280 ;
        RECT 52.515 108.220 52.805 108.265 ;
        RECT 62.620 108.220 62.940 108.280 ;
        RECT 78.720 108.220 79.040 108.280 ;
        RECT 52.040 108.080 52.805 108.220 ;
        RECT 52.040 108.020 52.360 108.080 ;
        RECT 52.515 108.035 52.805 108.080 ;
        RECT 62.250 108.080 79.040 108.220 ;
        RECT 30.880 107.880 31.200 107.940 ;
        RECT 33.655 107.880 33.945 107.925 ;
        RECT 21.235 107.740 22.830 107.880 ;
        RECT 23.150 107.740 26.510 107.880 ;
        RECT 21.235 107.695 21.525 107.740 ;
        RECT 17.555 107.355 17.845 107.585 ;
        RECT 18.935 107.540 19.225 107.585 ;
        RECT 20.760 107.540 21.080 107.600 ;
        RECT 23.150 107.585 23.290 107.740 ;
        RECT 26.370 107.600 26.510 107.740 ;
        RECT 30.880 107.740 33.945 107.880 ;
        RECT 30.880 107.680 31.200 107.740 ;
        RECT 33.655 107.695 33.945 107.740 ;
        RECT 34.100 107.880 34.420 107.940 ;
        RECT 34.655 107.880 34.945 107.925 ;
        RECT 40.630 107.880 40.770 108.020 ;
        RECT 47.440 107.880 47.760 107.940 ;
        RECT 34.100 107.740 34.945 107.880 ;
        RECT 34.100 107.680 34.420 107.740 ;
        RECT 34.655 107.695 34.945 107.740 ;
        RECT 36.950 107.740 40.770 107.880 ;
        RECT 44.770 107.740 47.760 107.880 ;
        RECT 18.935 107.400 21.080 107.540 ;
        RECT 18.935 107.355 19.225 107.400 ;
        RECT 17.630 107.200 17.770 107.355 ;
        RECT 20.760 107.340 21.080 107.400 ;
        RECT 23.075 107.355 23.365 107.585 ;
        RECT 23.520 107.340 23.840 107.600 ;
        RECT 23.980 107.340 24.300 107.600 ;
        RECT 24.900 107.340 25.220 107.600 ;
        RECT 25.375 107.355 25.665 107.585 ;
        RECT 22.615 107.200 22.905 107.245 ;
        RECT 17.630 107.060 22.905 107.200 ;
        RECT 23.610 107.200 23.750 107.340 ;
        RECT 25.450 107.200 25.590 107.355 ;
        RECT 26.280 107.340 26.600 107.600 ;
        RECT 36.950 107.585 37.090 107.740 ;
        RECT 36.875 107.355 37.165 107.585 ;
        RECT 38.240 107.340 38.560 107.600 ;
        RECT 39.635 107.540 39.925 107.585 ;
        RECT 40.080 107.540 40.400 107.600 ;
        RECT 44.770 107.585 44.910 107.740 ;
        RECT 47.440 107.680 47.760 107.740 ;
        RECT 49.280 107.880 49.600 107.940 ;
        RECT 52.975 107.880 53.265 107.925 ;
        RECT 49.280 107.740 53.265 107.880 ;
        RECT 49.280 107.680 49.600 107.740 ;
        RECT 52.975 107.695 53.265 107.740 ;
        RECT 54.815 107.880 55.105 107.925 ;
        RECT 56.035 107.880 56.325 107.925 ;
        RECT 54.815 107.740 56.325 107.880 ;
        RECT 54.815 107.695 55.105 107.740 ;
        RECT 56.035 107.695 56.325 107.740 ;
        RECT 57.115 107.695 57.405 107.925 ;
        RECT 39.635 107.400 40.400 107.540 ;
        RECT 39.635 107.355 39.925 107.400 ;
        RECT 40.080 107.340 40.400 107.400 ;
        RECT 40.555 107.355 40.845 107.585 ;
        RECT 44.695 107.355 44.985 107.585 ;
        RECT 23.610 107.060 25.590 107.200 ;
        RECT 38.330 107.200 38.470 107.340 ;
        RECT 40.630 107.200 40.770 107.355 ;
        RECT 45.140 107.340 45.460 107.600 ;
        RECT 46.520 107.340 46.840 107.600 ;
        RECT 48.835 107.540 49.125 107.585 ;
        RECT 49.740 107.540 50.060 107.600 ;
        RECT 48.835 107.400 50.060 107.540 ;
        RECT 48.835 107.355 49.125 107.400 ;
        RECT 49.740 107.340 50.060 107.400 ;
        RECT 50.200 107.540 50.520 107.600 ;
        RECT 52.500 107.540 52.820 107.600 ;
        RECT 53.895 107.540 54.185 107.585 ;
        RECT 50.200 107.400 54.185 107.540 ;
        RECT 50.200 107.340 50.520 107.400 ;
        RECT 52.500 107.340 52.820 107.400 ;
        RECT 53.895 107.355 54.185 107.400 ;
        RECT 54.340 107.540 54.660 107.600 ;
        RECT 57.190 107.540 57.330 107.695 ;
        RECT 62.250 107.585 62.390 108.080 ;
        RECT 62.620 108.020 62.940 108.080 ;
        RECT 78.720 108.020 79.040 108.080 ;
        RECT 84.700 108.220 85.020 108.280 ;
        RECT 85.635 108.220 85.925 108.265 ;
        RECT 84.700 108.080 85.925 108.220 ;
        RECT 84.700 108.020 85.020 108.080 ;
        RECT 85.635 108.035 85.925 108.080 ;
        RECT 87.460 108.220 87.780 108.280 ;
        RECT 91.155 108.220 91.445 108.265 ;
        RECT 129.780 108.220 130.100 108.280 ;
        RECT 87.460 108.080 91.445 108.220 ;
        RECT 87.460 108.020 87.780 108.080 ;
        RECT 91.155 108.035 91.445 108.080 ;
        RECT 101.810 108.080 130.100 108.220 ;
        RECT 63.095 107.880 63.385 107.925 ;
        RECT 68.140 107.880 68.460 107.940 ;
        RECT 85.160 107.880 85.480 107.940 ;
        RECT 101.810 107.880 101.950 108.080 ;
        RECT 129.780 108.020 130.100 108.080 ;
        RECT 104.480 107.925 104.800 107.940 ;
        RECT 104.450 107.880 104.800 107.925 ;
        RECT 125.655 107.880 125.945 107.925 ;
        RECT 127.340 107.880 127.630 107.925 ;
        RECT 63.095 107.740 68.460 107.880 ;
        RECT 63.095 107.695 63.385 107.740 ;
        RECT 68.140 107.680 68.460 107.740 ;
        RECT 74.210 107.740 78.950 107.880 ;
        RECT 54.340 107.400 57.330 107.540 ;
        RECT 54.340 107.340 54.660 107.400 ;
        RECT 62.175 107.355 62.465 107.585 ;
        RECT 62.620 107.340 62.940 107.600 ;
        RECT 74.210 107.585 74.350 107.740 ;
        RECT 63.785 107.540 64.075 107.585 ;
        RECT 66.775 107.540 67.065 107.585 ;
        RECT 63.785 107.400 67.065 107.540 ;
        RECT 63.785 107.355 64.075 107.400 ;
        RECT 66.775 107.355 67.065 107.400 ;
        RECT 74.135 107.355 74.425 107.585 ;
        RECT 75.470 107.540 75.760 107.585 ;
        RECT 78.260 107.540 78.580 107.600 ;
        RECT 75.470 107.400 78.580 107.540 ;
        RECT 78.810 107.540 78.950 107.740 ;
        RECT 85.160 107.740 101.950 107.880 ;
        RECT 104.285 107.740 104.800 107.880 ;
        RECT 85.160 107.680 85.480 107.740 ;
        RECT 104.450 107.695 104.800 107.740 ;
        RECT 104.480 107.680 104.800 107.695 ;
        RECT 118.140 107.740 124.950 107.880 ;
        RECT 85.620 107.540 85.940 107.600 ;
        RECT 78.810 107.400 85.940 107.540 ;
        RECT 75.470 107.355 75.760 107.400 ;
        RECT 78.260 107.340 78.580 107.400 ;
        RECT 85.620 107.340 85.940 107.400 ;
        RECT 87.000 107.340 87.320 107.600 ;
        RECT 87.460 107.340 87.780 107.600 ;
        RECT 87.920 107.340 88.240 107.600 ;
        RECT 88.855 107.355 89.145 107.585 ;
        RECT 91.600 107.540 91.920 107.600 ;
        RECT 92.075 107.540 92.365 107.585 ;
        RECT 91.600 107.400 92.365 107.540 ;
        RECT 38.330 107.060 40.770 107.200 ;
        RECT 47.455 107.200 47.745 107.245 ;
        RECT 49.295 107.200 49.585 107.245 ;
        RECT 47.455 107.060 49.585 107.200 ;
        RECT 20.850 106.580 20.990 107.060 ;
        RECT 22.615 107.015 22.905 107.060 ;
        RECT 47.455 107.015 47.745 107.060 ;
        RECT 49.295 107.015 49.585 107.060 ;
        RECT 22.690 106.860 22.830 107.015 ;
        RECT 64.460 107.000 64.780 107.260 ;
        RECT 67.680 107.200 68.000 107.260 ;
        RECT 69.535 107.200 69.825 107.245 ;
        RECT 67.680 107.060 69.825 107.200 ;
        RECT 67.680 107.000 68.000 107.060 ;
        RECT 69.535 107.015 69.825 107.060 ;
        RECT 75.015 107.200 75.305 107.245 ;
        RECT 76.205 107.200 76.495 107.245 ;
        RECT 78.725 107.200 79.015 107.245 ;
        RECT 75.015 107.060 79.015 107.200 ;
        RECT 75.015 107.015 75.305 107.060 ;
        RECT 76.205 107.015 76.495 107.060 ;
        RECT 78.725 107.015 79.015 107.060 ;
        RECT 81.480 107.200 81.800 107.260 ;
        RECT 88.930 107.200 89.070 107.355 ;
        RECT 91.600 107.340 91.920 107.400 ;
        RECT 92.075 107.355 92.365 107.400 ;
        RECT 92.520 107.340 92.840 107.600 ;
        RECT 92.980 107.340 93.300 107.600 ;
        RECT 93.915 107.540 94.205 107.585 ;
        RECT 106.780 107.540 107.100 107.600 ;
        RECT 93.915 107.400 107.100 107.540 ;
        RECT 93.915 107.355 94.205 107.400 ;
        RECT 106.780 107.340 107.100 107.400 ;
        RECT 114.140 107.340 114.460 107.600 ;
        RECT 114.615 107.355 114.905 107.585 ;
        RECT 115.060 107.540 115.380 107.600 ;
        RECT 116.440 107.540 116.760 107.600 ;
        RECT 118.140 107.540 118.280 107.740 ;
        RECT 115.060 107.400 118.280 107.540 ;
        RECT 122.435 107.540 122.725 107.585 ;
        RECT 122.880 107.540 123.200 107.600 ;
        RECT 122.435 107.400 123.200 107.540 ;
        RECT 89.760 107.200 90.080 107.260 ;
        RECT 93.070 107.200 93.210 107.340 ;
        RECT 81.480 107.060 90.080 107.200 ;
        RECT 81.480 107.000 81.800 107.060 ;
        RECT 89.760 107.000 90.080 107.060 ;
        RECT 92.610 107.060 93.210 107.200 ;
        RECT 24.900 106.860 25.220 106.920 ;
        RECT 28.580 106.860 28.900 106.920 ;
        RECT 40.095 106.860 40.385 106.905 ;
        RECT 22.690 106.720 28.900 106.860 ;
        RECT 24.900 106.660 25.220 106.720 ;
        RECT 28.580 106.660 28.900 106.720 ;
        RECT 34.650 106.720 40.385 106.860 ;
        RECT 20.300 106.320 20.620 106.580 ;
        RECT 20.760 106.320 21.080 106.580 ;
        RECT 34.650 106.565 34.790 106.720 ;
        RECT 40.095 106.675 40.385 106.720 ;
        RECT 49.740 106.860 50.060 106.920 ;
        RECT 74.620 106.860 74.910 106.905 ;
        RECT 76.720 106.860 77.010 106.905 ;
        RECT 78.290 106.860 78.580 106.905 ;
        RECT 49.740 106.720 56.410 106.860 ;
        RECT 49.740 106.660 50.060 106.720 ;
        RECT 34.575 106.335 34.865 106.565 ;
        RECT 35.480 106.320 35.800 106.580 ;
        RECT 35.955 106.520 36.245 106.565 ;
        RECT 36.400 106.520 36.720 106.580 ;
        RECT 35.955 106.380 36.720 106.520 ;
        RECT 35.955 106.335 36.245 106.380 ;
        RECT 36.400 106.320 36.720 106.380 ;
        RECT 46.075 106.520 46.365 106.565 ;
        RECT 49.280 106.520 49.600 106.580 ;
        RECT 46.075 106.380 49.600 106.520 ;
        RECT 46.075 106.335 46.365 106.380 ;
        RECT 49.280 106.320 49.600 106.380 ;
        RECT 55.260 106.320 55.580 106.580 ;
        RECT 56.270 106.565 56.410 106.720 ;
        RECT 74.620 106.720 78.580 106.860 ;
        RECT 74.620 106.675 74.910 106.720 ;
        RECT 76.720 106.675 77.010 106.720 ;
        RECT 78.290 106.675 78.580 106.720 ;
        RECT 80.100 106.860 80.420 106.920 ;
        RECT 88.840 106.860 89.160 106.920 ;
        RECT 92.610 106.860 92.750 107.060 ;
        RECT 103.100 107.000 103.420 107.260 ;
        RECT 103.995 107.200 104.285 107.245 ;
        RECT 105.185 107.200 105.475 107.245 ;
        RECT 107.705 107.200 107.995 107.245 ;
        RECT 103.995 107.060 107.995 107.200 ;
        RECT 103.995 107.015 104.285 107.060 ;
        RECT 105.185 107.015 105.475 107.060 ;
        RECT 107.705 107.015 107.995 107.060 ;
        RECT 109.080 107.200 109.400 107.260 ;
        RECT 114.690 107.200 114.830 107.355 ;
        RECT 115.060 107.340 115.380 107.400 ;
        RECT 116.440 107.340 116.760 107.400 ;
        RECT 122.435 107.355 122.725 107.400 ;
        RECT 122.880 107.340 123.200 107.400 ;
        RECT 123.340 107.340 123.660 107.600 ;
        RECT 123.800 107.340 124.120 107.600 ;
        RECT 124.260 107.340 124.580 107.600 ;
        RECT 124.810 107.540 124.950 107.740 ;
        RECT 125.655 107.740 127.630 107.880 ;
        RECT 125.655 107.695 125.945 107.740 ;
        RECT 127.340 107.695 127.630 107.740 ;
        RECT 134.855 107.880 135.145 107.925 ;
        RECT 135.760 107.880 136.080 107.940 ;
        RECT 134.855 107.740 136.080 107.880 ;
        RECT 134.855 107.695 135.145 107.740 ;
        RECT 135.760 107.680 136.080 107.740 ;
        RECT 126.560 107.540 126.880 107.600 ;
        RECT 124.810 107.400 126.880 107.540 ;
        RECT 126.560 107.340 126.880 107.400 ;
        RECT 131.160 107.540 131.480 107.600 ;
        RECT 134.395 107.540 134.685 107.585 ;
        RECT 131.160 107.400 134.685 107.540 ;
        RECT 131.160 107.340 131.480 107.400 ;
        RECT 134.395 107.355 134.685 107.400 ;
        RECT 135.315 107.355 135.605 107.585 ;
        RECT 136.235 107.355 136.525 107.585 ;
        RECT 120.580 107.200 120.900 107.260 ;
        RECT 109.080 107.060 120.900 107.200 ;
        RECT 109.080 107.000 109.400 107.060 ;
        RECT 120.580 107.000 120.900 107.060 ;
        RECT 121.040 107.200 121.360 107.260 ;
        RECT 126.115 107.200 126.405 107.245 ;
        RECT 121.040 107.060 126.405 107.200 ;
        RECT 121.040 107.000 121.360 107.060 ;
        RECT 126.115 107.015 126.405 107.060 ;
        RECT 126.995 107.200 127.285 107.245 ;
        RECT 128.185 107.200 128.475 107.245 ;
        RECT 130.705 107.200 130.995 107.245 ;
        RECT 126.995 107.060 130.995 107.200 ;
        RECT 126.995 107.015 127.285 107.060 ;
        RECT 128.185 107.015 128.475 107.060 ;
        RECT 130.705 107.015 130.995 107.060 ;
        RECT 131.620 107.200 131.940 107.260 ;
        RECT 135.390 107.200 135.530 107.355 ;
        RECT 131.620 107.060 135.530 107.200 ;
        RECT 131.620 107.000 131.940 107.060 ;
        RECT 80.100 106.720 87.690 106.860 ;
        RECT 80.100 106.660 80.420 106.720 ;
        RECT 87.550 106.580 87.690 106.720 ;
        RECT 88.840 106.720 92.750 106.860 ;
        RECT 103.600 106.860 103.890 106.905 ;
        RECT 105.700 106.860 105.990 106.905 ;
        RECT 107.270 106.860 107.560 106.905 ;
        RECT 103.600 106.720 107.560 106.860 ;
        RECT 88.840 106.660 89.160 106.720 ;
        RECT 103.600 106.675 103.890 106.720 ;
        RECT 105.700 106.675 105.990 106.720 ;
        RECT 107.270 106.675 107.560 106.720 ;
        RECT 110.460 106.860 110.780 106.920 ;
        RECT 116.440 106.860 116.760 106.920 ;
        RECT 110.460 106.720 116.760 106.860 ;
        RECT 110.460 106.660 110.780 106.720 ;
        RECT 116.440 106.660 116.760 106.720 ;
        RECT 126.600 106.860 126.890 106.905 ;
        RECT 128.700 106.860 128.990 106.905 ;
        RECT 130.270 106.860 130.560 106.905 ;
        RECT 126.600 106.720 130.560 106.860 ;
        RECT 126.600 106.675 126.890 106.720 ;
        RECT 128.700 106.675 128.990 106.720 ;
        RECT 130.270 106.675 130.560 106.720 ;
        RECT 132.540 106.860 132.860 106.920 ;
        RECT 134.380 106.860 134.700 106.920 ;
        RECT 136.310 106.860 136.450 107.355 ;
        RECT 132.540 106.720 134.150 106.860 ;
        RECT 132.540 106.660 132.860 106.720 ;
        RECT 56.195 106.335 56.485 106.565 ;
        RECT 61.255 106.520 61.545 106.565 ;
        RECT 61.700 106.520 62.020 106.580 ;
        RECT 61.255 106.380 62.020 106.520 ;
        RECT 61.255 106.335 61.545 106.380 ;
        RECT 61.700 106.320 62.020 106.380 ;
        RECT 77.340 106.520 77.660 106.580 ;
        RECT 79.180 106.520 79.500 106.580 ;
        RECT 81.035 106.520 81.325 106.565 ;
        RECT 77.340 106.380 81.325 106.520 ;
        RECT 77.340 106.320 77.660 106.380 ;
        RECT 79.180 106.320 79.500 106.380 ;
        RECT 81.035 106.335 81.325 106.380 ;
        RECT 87.460 106.520 87.780 106.580 ;
        RECT 94.820 106.520 95.140 106.580 ;
        RECT 87.460 106.380 95.140 106.520 ;
        RECT 87.460 106.320 87.780 106.380 ;
        RECT 94.820 106.320 95.140 106.380 ;
        RECT 106.780 106.520 107.100 106.580 ;
        RECT 110.015 106.520 110.305 106.565 ;
        RECT 112.300 106.520 112.620 106.580 ;
        RECT 106.780 106.380 112.620 106.520 ;
        RECT 106.780 106.320 107.100 106.380 ;
        RECT 110.015 106.335 110.305 106.380 ;
        RECT 112.300 106.320 112.620 106.380 ;
        RECT 115.520 106.320 115.840 106.580 ;
        RECT 127.940 106.520 128.260 106.580 ;
        RECT 133.090 106.565 133.230 106.720 ;
        RECT 133.015 106.520 133.305 106.565 ;
        RECT 127.940 106.380 133.305 106.520 ;
        RECT 127.940 106.320 128.260 106.380 ;
        RECT 133.015 106.335 133.305 106.380 ;
        RECT 133.460 106.320 133.780 106.580 ;
        RECT 134.010 106.520 134.150 106.720 ;
        RECT 134.380 106.720 136.450 106.860 ;
        RECT 134.380 106.660 134.700 106.720 ;
        RECT 135.760 106.520 136.080 106.580 ;
        RECT 134.010 106.380 136.080 106.520 ;
        RECT 135.760 106.320 136.080 106.380 ;
        RECT 13.330 105.700 138.910 106.180 ;
        RECT 20.300 105.500 20.620 105.560 ;
        RECT 29.960 105.500 30.280 105.560 ;
        RECT 20.300 105.360 30.280 105.500 ;
        RECT 20.300 105.300 20.620 105.360 ;
        RECT 29.960 105.300 30.280 105.360 ;
        RECT 31.815 105.500 32.105 105.545 ;
        RECT 34.100 105.500 34.420 105.560 ;
        RECT 31.815 105.360 34.420 105.500 ;
        RECT 31.815 105.315 32.105 105.360 ;
        RECT 34.100 105.300 34.420 105.360 ;
        RECT 35.480 105.500 35.800 105.560 ;
        RECT 35.480 105.360 41.690 105.500 ;
        RECT 35.480 105.300 35.800 105.360 ;
        RECT 34.600 105.160 34.890 105.205 ;
        RECT 36.700 105.160 36.990 105.205 ;
        RECT 38.270 105.160 38.560 105.205 ;
        RECT 34.600 105.020 38.560 105.160 ;
        RECT 34.600 104.975 34.890 105.020 ;
        RECT 36.700 104.975 36.990 105.020 ;
        RECT 38.270 104.975 38.560 105.020 ;
        RECT 40.540 105.160 40.860 105.220 ;
        RECT 41.015 105.160 41.305 105.205 ;
        RECT 40.540 105.020 41.305 105.160 ;
        RECT 40.540 104.960 40.860 105.020 ;
        RECT 41.015 104.975 41.305 105.020 ;
        RECT 34.995 104.820 35.285 104.865 ;
        RECT 36.185 104.820 36.475 104.865 ;
        RECT 38.705 104.820 38.995 104.865 ;
        RECT 34.995 104.680 38.995 104.820 ;
        RECT 34.995 104.635 35.285 104.680 ;
        RECT 36.185 104.635 36.475 104.680 ;
        RECT 38.705 104.635 38.995 104.680 ;
        RECT 21.220 104.480 21.540 104.540 ;
        RECT 23.075 104.480 23.365 104.525 ;
        RECT 23.520 104.480 23.840 104.540 ;
        RECT 21.220 104.340 23.840 104.480 ;
        RECT 21.220 104.280 21.540 104.340 ;
        RECT 23.075 104.295 23.365 104.340 ;
        RECT 23.520 104.280 23.840 104.340 ;
        RECT 34.100 104.280 34.420 104.540 ;
        RECT 38.240 104.480 38.560 104.540 ;
        RECT 35.110 104.340 38.560 104.480 ;
        RECT 41.550 104.480 41.690 105.360 ;
        RECT 50.660 105.300 50.980 105.560 ;
        RECT 52.500 105.300 52.820 105.560 ;
        RECT 78.260 105.300 78.580 105.560 ;
        RECT 82.415 105.500 82.705 105.545 ;
        RECT 84.240 105.500 84.560 105.560 ;
        RECT 82.415 105.360 84.560 105.500 ;
        RECT 82.415 105.315 82.705 105.360 ;
        RECT 84.240 105.300 84.560 105.360 ;
        RECT 87.000 105.500 87.320 105.560 ;
        RECT 99.420 105.500 99.740 105.560 ;
        RECT 87.000 105.360 99.740 105.500 ;
        RECT 87.000 105.300 87.320 105.360 ;
        RECT 99.420 105.300 99.740 105.360 ;
        RECT 116.440 105.500 116.760 105.560 ;
        RECT 118.280 105.500 118.600 105.560 ;
        RECT 116.440 105.360 118.600 105.500 ;
        RECT 116.440 105.300 116.760 105.360 ;
        RECT 118.280 105.300 118.600 105.360 ;
        RECT 123.340 105.500 123.660 105.560 ;
        RECT 127.035 105.500 127.325 105.545 ;
        RECT 123.340 105.360 127.325 105.500 ;
        RECT 123.340 105.300 123.660 105.360 ;
        RECT 127.035 105.315 127.325 105.360 ;
        RECT 127.480 105.500 127.800 105.560 ;
        RECT 134.380 105.500 134.700 105.560 ;
        RECT 127.480 105.360 134.700 105.500 ;
        RECT 127.480 105.300 127.800 105.360 ;
        RECT 134.380 105.300 134.700 105.360 ;
        RECT 136.680 105.300 137.000 105.560 ;
        RECT 44.220 105.160 44.510 105.205 ;
        RECT 45.790 105.160 46.080 105.205 ;
        RECT 47.890 105.160 48.180 105.205 ;
        RECT 44.220 105.020 48.180 105.160 ;
        RECT 44.220 104.975 44.510 105.020 ;
        RECT 45.790 104.975 46.080 105.020 ;
        RECT 47.890 104.975 48.180 105.020 ;
        RECT 48.835 105.160 49.125 105.205 ;
        RECT 49.280 105.160 49.600 105.220 ;
        RECT 48.835 105.020 49.600 105.160 ;
        RECT 48.835 104.975 49.125 105.020 ;
        RECT 49.280 104.960 49.600 105.020 ;
        RECT 55.260 105.160 55.550 105.205 ;
        RECT 56.830 105.160 57.120 105.205 ;
        RECT 58.930 105.160 59.220 105.205 ;
        RECT 55.260 105.020 59.220 105.160 ;
        RECT 55.260 104.975 55.550 105.020 ;
        RECT 56.830 104.975 57.120 105.020 ;
        RECT 58.930 104.975 59.220 105.020 ;
        RECT 60.820 105.160 61.110 105.205 ;
        RECT 62.920 105.160 63.210 105.205 ;
        RECT 64.490 105.160 64.780 105.205 ;
        RECT 60.820 105.020 64.780 105.160 ;
        RECT 60.820 104.975 61.110 105.020 ;
        RECT 62.920 104.975 63.210 105.020 ;
        RECT 64.490 104.975 64.780 105.020 ;
        RECT 76.880 104.960 77.200 105.220 ;
        RECT 78.720 105.160 79.040 105.220 ;
        RECT 81.480 105.160 81.800 105.220 ;
        RECT 78.720 105.020 81.800 105.160 ;
        RECT 78.720 104.960 79.040 105.020 ;
        RECT 81.480 104.960 81.800 105.020 ;
        RECT 86.120 105.160 86.410 105.205 ;
        RECT 88.220 105.160 88.510 105.205 ;
        RECT 89.790 105.160 90.080 105.205 ;
        RECT 86.120 105.020 90.080 105.160 ;
        RECT 86.120 104.975 86.410 105.020 ;
        RECT 88.220 104.975 88.510 105.020 ;
        RECT 89.790 104.975 90.080 105.020 ;
        RECT 92.520 105.160 92.840 105.220 ;
        RECT 93.900 105.160 94.220 105.220 ;
        RECT 92.520 105.020 94.220 105.160 ;
        RECT 92.520 104.960 92.840 105.020 ;
        RECT 93.900 104.960 94.220 105.020 ;
        RECT 96.200 104.960 96.520 105.220 ;
        RECT 104.480 105.160 104.800 105.220 ;
        RECT 110.460 105.160 110.780 105.220 ;
        RECT 104.480 105.020 110.780 105.160 ;
        RECT 104.480 104.960 104.800 105.020 ;
        RECT 110.460 104.960 110.780 105.020 ;
        RECT 111.880 105.160 112.170 105.205 ;
        RECT 113.980 105.160 114.270 105.205 ;
        RECT 115.550 105.160 115.840 105.205 ;
        RECT 111.880 105.020 115.840 105.160 ;
        RECT 111.880 104.975 112.170 105.020 ;
        RECT 113.980 104.975 114.270 105.020 ;
        RECT 115.550 104.975 115.840 105.020 ;
        RECT 126.560 105.160 126.880 105.220 ;
        RECT 134.855 105.160 135.145 105.205 ;
        RECT 126.560 105.020 135.145 105.160 ;
        RECT 126.560 104.960 126.880 105.020 ;
        RECT 134.855 104.975 135.145 105.020 ;
        RECT 43.785 104.820 44.075 104.865 ;
        RECT 46.305 104.820 46.595 104.865 ;
        RECT 47.495 104.820 47.785 104.865 ;
        RECT 43.785 104.680 47.785 104.820 ;
        RECT 43.785 104.635 44.075 104.680 ;
        RECT 46.305 104.635 46.595 104.680 ;
        RECT 47.495 104.635 47.785 104.680 ;
        RECT 48.375 104.820 48.665 104.865 ;
        RECT 51.580 104.820 51.900 104.880 ;
        RECT 48.375 104.680 51.900 104.820 ;
        RECT 48.375 104.635 48.665 104.680 ;
        RECT 51.580 104.620 51.900 104.680 ;
        RECT 54.825 104.820 55.115 104.865 ;
        RECT 57.345 104.820 57.635 104.865 ;
        RECT 58.535 104.820 58.825 104.865 ;
        RECT 54.825 104.680 58.825 104.820 ;
        RECT 54.825 104.635 55.115 104.680 ;
        RECT 57.345 104.635 57.635 104.680 ;
        RECT 58.535 104.635 58.825 104.680 ;
        RECT 61.215 104.820 61.505 104.865 ;
        RECT 62.405 104.820 62.695 104.865 ;
        RECT 64.925 104.820 65.215 104.865 ;
        RECT 61.215 104.680 65.215 104.820 ;
        RECT 61.215 104.635 61.505 104.680 ;
        RECT 62.405 104.635 62.695 104.680 ;
        RECT 64.925 104.635 65.215 104.680 ;
        RECT 47.040 104.480 47.330 104.525 ;
        RECT 41.550 104.340 47.330 104.480 ;
        RECT 51.670 104.480 51.810 104.620 ;
        RECT 59.415 104.480 59.705 104.525 ;
        RECT 60.320 104.480 60.640 104.540 ;
        RECT 61.700 104.525 62.020 104.540 ;
        RECT 61.670 104.480 62.020 104.525 ;
        RECT 51.670 104.340 60.640 104.480 ;
        RECT 61.505 104.340 62.020 104.480 ;
        RECT 76.970 104.480 77.110 104.960 ;
        RECT 77.800 104.820 78.120 104.880 ;
        RECT 77.800 104.680 84.470 104.820 ;
        RECT 77.800 104.620 78.120 104.680 ;
        RECT 79.730 104.525 79.870 104.680 ;
        RECT 77.355 104.480 77.645 104.525 ;
        RECT 76.970 104.340 77.645 104.480 ;
        RECT 20.760 104.140 21.080 104.200 ;
        RECT 22.155 104.140 22.445 104.185 ;
        RECT 20.760 104.000 22.445 104.140 ;
        RECT 20.760 103.940 21.080 104.000 ;
        RECT 22.155 103.955 22.445 104.000 ;
        RECT 32.735 103.955 33.025 104.185 ;
        RECT 33.655 104.140 33.945 104.185 ;
        RECT 35.110 104.140 35.250 104.340 ;
        RECT 38.240 104.280 38.560 104.340 ;
        RECT 47.040 104.295 47.330 104.340 ;
        RECT 59.415 104.295 59.705 104.340 ;
        RECT 60.320 104.280 60.640 104.340 ;
        RECT 61.670 104.295 62.020 104.340 ;
        RECT 77.355 104.295 77.645 104.340 ;
        RECT 79.655 104.295 79.945 104.525 ;
        RECT 61.700 104.280 62.020 104.295 ;
        RECT 80.100 104.280 80.420 104.540 ;
        RECT 80.560 104.280 80.880 104.540 ;
        RECT 81.480 104.280 81.800 104.540 ;
        RECT 83.320 104.280 83.640 104.540 ;
        RECT 83.795 104.295 84.085 104.525 ;
        RECT 35.480 104.185 35.800 104.200 ;
        RECT 33.655 104.000 35.250 104.140 ;
        RECT 33.655 103.955 33.945 104.000 ;
        RECT 35.450 103.955 35.800 104.185 ;
        RECT 23.980 103.600 24.300 103.860 ;
        RECT 32.810 103.800 32.950 103.955 ;
        RECT 35.480 103.940 35.800 103.955 ;
        RECT 46.520 104.140 46.840 104.200 ;
        RECT 50.675 104.140 50.965 104.185 ;
        RECT 54.340 104.140 54.660 104.200 ;
        RECT 46.520 104.000 54.660 104.140 ;
        RECT 46.520 103.940 46.840 104.000 ;
        RECT 50.675 103.955 50.965 104.000 ;
        RECT 54.340 103.940 54.660 104.000 ;
        RECT 55.260 104.140 55.580 104.200 ;
        RECT 58.080 104.140 58.370 104.185 ;
        RECT 55.260 104.000 58.370 104.140 ;
        RECT 55.260 103.940 55.580 104.000 ;
        RECT 58.080 103.955 58.370 104.000 ;
        RECT 76.435 104.140 76.725 104.185 ;
        RECT 76.880 104.140 77.200 104.200 ;
        RECT 76.435 104.000 77.200 104.140 ;
        RECT 76.435 103.955 76.725 104.000 ;
        RECT 76.880 103.940 77.200 104.000 ;
        RECT 78.260 104.140 78.580 104.200 ;
        RECT 83.870 104.140 84.010 104.295 ;
        RECT 78.260 104.000 84.010 104.140 ;
        RECT 78.260 103.940 78.580 104.000 ;
        RECT 40.080 103.800 40.400 103.860 ;
        RECT 41.000 103.800 41.320 103.860 ;
        RECT 41.475 103.800 41.765 103.845 ;
        RECT 32.810 103.660 41.765 103.800 ;
        RECT 40.080 103.600 40.400 103.660 ;
        RECT 41.000 103.600 41.320 103.660 ;
        RECT 41.475 103.615 41.765 103.660 ;
        RECT 51.120 103.800 51.440 103.860 ;
        RECT 51.595 103.800 51.885 103.845 ;
        RECT 51.120 103.660 51.885 103.800 ;
        RECT 51.120 103.600 51.440 103.660 ;
        RECT 51.595 103.615 51.885 103.660 ;
        RECT 67.235 103.800 67.525 103.845 ;
        RECT 67.680 103.800 68.000 103.860 ;
        RECT 67.235 103.660 68.000 103.800 ;
        RECT 67.235 103.615 67.525 103.660 ;
        RECT 67.680 103.600 68.000 103.660 ;
        RECT 75.515 103.800 75.805 103.845 ;
        RECT 80.560 103.800 80.880 103.860 ;
        RECT 75.515 103.660 80.880 103.800 ;
        RECT 84.330 103.800 84.470 104.680 ;
        RECT 85.620 104.620 85.940 104.880 ;
        RECT 86.515 104.820 86.805 104.865 ;
        RECT 87.705 104.820 87.995 104.865 ;
        RECT 90.225 104.820 90.515 104.865 ;
        RECT 86.515 104.680 90.515 104.820 ;
        RECT 86.515 104.635 86.805 104.680 ;
        RECT 87.705 104.635 87.995 104.680 ;
        RECT 90.225 104.635 90.515 104.680 ;
        RECT 91.600 104.820 91.920 104.880 ;
        RECT 96.660 104.820 96.980 104.880 ;
        RECT 103.100 104.820 103.420 104.880 ;
        RECT 112.275 104.820 112.565 104.865 ;
        RECT 113.465 104.820 113.755 104.865 ;
        RECT 115.985 104.820 116.275 104.865 ;
        RECT 91.600 104.680 99.190 104.820 ;
        RECT 91.600 104.620 91.920 104.680 ;
        RECT 84.700 104.280 85.020 104.540 ;
        RECT 85.175 104.480 85.465 104.525 ;
        RECT 86.080 104.480 86.400 104.540 ;
        RECT 96.290 104.525 96.430 104.680 ;
        RECT 96.660 104.620 96.980 104.680 ;
        RECT 99.050 104.540 99.190 104.680 ;
        RECT 103.100 104.680 111.610 104.820 ;
        RECT 103.100 104.620 103.420 104.680 ;
        RECT 85.175 104.340 86.400 104.480 ;
        RECT 85.175 104.295 85.465 104.340 ;
        RECT 86.080 104.280 86.400 104.340 ;
        RECT 96.215 104.295 96.505 104.525 ;
        RECT 97.135 104.480 97.425 104.525 ;
        RECT 97.135 104.340 98.730 104.480 ;
        RECT 97.135 104.295 97.425 104.340 ;
        RECT 87.000 104.185 87.320 104.200 ;
        RECT 86.970 103.955 87.320 104.185 ;
        RECT 87.000 103.940 87.320 103.955 ;
        RECT 93.900 103.940 94.220 104.200 ;
        RECT 94.820 104.140 95.140 104.200 ;
        RECT 98.055 104.140 98.345 104.185 ;
        RECT 94.820 104.000 98.345 104.140 ;
        RECT 98.590 104.140 98.730 104.340 ;
        RECT 98.960 104.280 99.280 104.540 ;
        RECT 99.895 104.295 100.185 104.525 ;
        RECT 99.970 104.140 100.110 104.295 ;
        RECT 109.080 104.280 109.400 104.540 ;
        RECT 111.470 104.525 111.610 104.680 ;
        RECT 112.275 104.680 116.275 104.820 ;
        RECT 112.275 104.635 112.565 104.680 ;
        RECT 113.465 104.635 113.755 104.680 ;
        RECT 115.985 104.635 116.275 104.680 ;
        RECT 129.870 104.680 133.230 104.820 ;
        RECT 110.475 104.295 110.765 104.525 ;
        RECT 111.395 104.480 111.685 104.525 ;
        RECT 118.740 104.480 119.060 104.540 ;
        RECT 121.040 104.480 121.360 104.540 ;
        RECT 126.575 104.480 126.865 104.525 ;
        RECT 111.395 104.340 121.360 104.480 ;
        RECT 111.395 104.295 111.685 104.340 ;
        RECT 110.550 104.140 110.690 104.295 ;
        RECT 118.740 104.280 119.060 104.340 ;
        RECT 121.040 104.280 121.360 104.340 ;
        RECT 125.270 104.340 128.630 104.480 ;
        RECT 98.590 104.000 110.690 104.140 ;
        RECT 94.820 103.940 95.140 104.000 ;
        RECT 98.055 103.955 98.345 104.000 ;
        RECT 88.380 103.800 88.700 103.860 ;
        RECT 84.330 103.660 88.700 103.800 ;
        RECT 75.515 103.615 75.805 103.660 ;
        RECT 80.560 103.600 80.880 103.660 ;
        RECT 88.380 103.600 88.700 103.660 ;
        RECT 92.980 103.600 93.300 103.860 ;
        RECT 110.550 103.800 110.690 104.000 ;
        RECT 110.935 104.140 111.225 104.185 ;
        RECT 111.840 104.140 112.160 104.200 ;
        RECT 110.935 104.000 112.160 104.140 ;
        RECT 110.935 103.955 111.225 104.000 ;
        RECT 111.840 103.940 112.160 104.000 ;
        RECT 112.730 104.140 113.020 104.185 ;
        RECT 114.600 104.140 114.920 104.200 ;
        RECT 112.730 104.000 114.920 104.140 ;
        RECT 112.730 103.955 113.020 104.000 ;
        RECT 114.600 103.940 114.920 104.000 ;
        RECT 115.520 104.140 115.840 104.200 ;
        RECT 125.270 104.140 125.410 104.340 ;
        RECT 126.575 104.295 126.865 104.340 ;
        RECT 115.520 104.000 125.410 104.140 ;
        RECT 125.655 104.140 125.945 104.185 ;
        RECT 127.480 104.140 127.800 104.200 ;
        RECT 125.655 104.000 127.800 104.140 ;
        RECT 115.520 103.940 115.840 104.000 ;
        RECT 125.655 103.955 125.945 104.000 ;
        RECT 127.480 103.940 127.800 104.000 ;
        RECT 127.940 103.940 128.260 104.200 ;
        RECT 128.490 104.140 128.630 104.340 ;
        RECT 128.875 104.140 129.165 104.185 ;
        RECT 129.870 104.140 130.010 104.680 ;
        RECT 130.700 104.280 131.020 104.540 ;
        RECT 131.175 104.480 131.465 104.525 ;
        RECT 132.080 104.480 132.400 104.540 ;
        RECT 133.090 104.525 133.230 104.680 ;
        RECT 131.175 104.340 132.400 104.480 ;
        RECT 131.175 104.295 131.465 104.340 ;
        RECT 132.080 104.280 132.400 104.340 ;
        RECT 132.555 104.295 132.845 104.525 ;
        RECT 133.015 104.295 133.305 104.525 ;
        RECT 128.490 104.000 130.010 104.140 ;
        RECT 128.875 103.955 129.165 104.000 ;
        RECT 131.620 103.940 131.940 104.200 ;
        RECT 132.630 104.140 132.770 104.295 ;
        RECT 135.760 104.280 136.080 104.540 ;
        RECT 133.935 104.140 134.225 104.185 ;
        RECT 135.300 104.140 135.620 104.200 ;
        RECT 132.630 104.000 135.620 104.140 ;
        RECT 133.935 103.955 134.225 104.000 ;
        RECT 135.300 103.940 135.620 104.000 ;
        RECT 114.140 103.800 114.460 103.860 ;
        RECT 110.550 103.660 114.460 103.800 ;
        RECT 114.140 103.600 114.460 103.660 ;
        RECT 118.280 103.800 118.600 103.860 ;
        RECT 124.260 103.800 124.580 103.860 ;
        RECT 118.280 103.660 124.580 103.800 ;
        RECT 118.280 103.600 118.600 103.660 ;
        RECT 124.260 103.600 124.580 103.660 ;
        RECT 124.735 103.800 125.025 103.845 ;
        RECT 125.180 103.800 125.500 103.860 ;
        RECT 124.735 103.660 125.500 103.800 ;
        RECT 124.735 103.615 125.025 103.660 ;
        RECT 125.180 103.600 125.500 103.660 ;
        RECT 126.100 103.800 126.420 103.860 ;
        RECT 129.795 103.800 130.085 103.845 ;
        RECT 126.100 103.660 130.085 103.800 ;
        RECT 126.100 103.600 126.420 103.660 ;
        RECT 129.795 103.615 130.085 103.660 ;
        RECT 13.330 102.980 138.910 103.460 ;
        RECT 17.540 102.580 17.860 102.840 ;
        RECT 23.980 102.780 24.300 102.840 ;
        RECT 29.845 102.780 30.135 102.825 ;
        RECT 23.980 102.640 30.135 102.780 ;
        RECT 23.980 102.580 24.300 102.640 ;
        RECT 29.845 102.595 30.135 102.640 ;
        RECT 35.480 102.580 35.800 102.840 ;
        RECT 36.415 102.780 36.705 102.825 ;
        RECT 36.860 102.780 37.180 102.840 ;
        RECT 36.415 102.640 37.180 102.780 ;
        RECT 36.415 102.595 36.705 102.640 ;
        RECT 36.860 102.580 37.180 102.640 ;
        RECT 38.240 102.780 38.560 102.840 ;
        RECT 40.635 102.780 40.925 102.825 ;
        RECT 38.240 102.640 40.925 102.780 ;
        RECT 38.240 102.580 38.560 102.640 ;
        RECT 40.635 102.595 40.925 102.640 ;
        RECT 41.475 102.595 41.765 102.825 ;
        RECT 46.995 102.780 47.285 102.825 ;
        RECT 50.660 102.780 50.980 102.840 ;
        RECT 80.100 102.780 80.420 102.840 ;
        RECT 46.995 102.640 50.980 102.780 ;
        RECT 46.995 102.595 47.285 102.640 ;
        RECT 17.630 102.440 17.770 102.580 ;
        RECT 17.630 102.300 28.810 102.440 ;
        RECT 17.555 101.915 17.845 102.145 ;
        RECT 18.475 102.100 18.765 102.145 ;
        RECT 21.220 102.100 21.540 102.160 ;
        RECT 28.670 102.145 28.810 102.300 ;
        RECT 30.880 102.240 31.200 102.500 ;
        RECT 39.635 102.440 39.925 102.485 ;
        RECT 40.080 102.440 40.400 102.500 ;
        RECT 39.635 102.300 40.400 102.440 ;
        RECT 39.635 102.255 39.925 102.300 ;
        RECT 40.080 102.240 40.400 102.300 ;
        RECT 41.550 102.440 41.690 102.595 ;
        RECT 50.660 102.580 50.980 102.640 ;
        RECT 76.050 102.640 80.420 102.780 ;
        RECT 45.140 102.440 45.460 102.500 ;
        RECT 41.550 102.300 45.460 102.440 ;
        RECT 18.475 101.960 21.540 102.100 ;
        RECT 18.475 101.915 18.765 101.960 ;
        RECT 17.630 101.760 17.770 101.915 ;
        RECT 21.220 101.900 21.540 101.960 ;
        RECT 27.315 102.100 27.605 102.145 ;
        RECT 28.595 102.100 28.885 102.145 ;
        RECT 34.100 102.100 34.420 102.160 ;
        RECT 27.315 101.960 28.350 102.100 ;
        RECT 27.315 101.915 27.605 101.960 ;
        RECT 24.005 101.760 24.295 101.805 ;
        RECT 26.525 101.760 26.815 101.805 ;
        RECT 27.715 101.760 28.005 101.805 ;
        RECT 17.630 101.620 20.990 101.760 ;
        RECT 20.850 101.480 20.990 101.620 ;
        RECT 24.005 101.620 28.005 101.760 ;
        RECT 28.210 101.760 28.350 101.960 ;
        RECT 28.595 101.960 34.420 102.100 ;
        RECT 28.595 101.915 28.885 101.960 ;
        RECT 34.100 101.900 34.420 101.960 ;
        RECT 38.255 102.100 38.545 102.145 ;
        RECT 41.550 102.100 41.690 102.300 ;
        RECT 45.140 102.240 45.460 102.300 ;
        RECT 46.075 102.440 46.365 102.485 ;
        RECT 47.440 102.440 47.760 102.500 ;
        RECT 46.075 102.300 47.760 102.440 ;
        RECT 46.075 102.255 46.365 102.300 ;
        RECT 47.440 102.240 47.760 102.300 ;
        RECT 51.580 102.440 51.900 102.500 ;
        RECT 51.580 102.300 54.570 102.440 ;
        RECT 51.580 102.240 51.900 102.300 ;
        RECT 38.255 101.960 41.690 102.100 ;
        RECT 51.120 102.100 51.440 102.160 ;
        RECT 54.430 102.145 54.570 102.300 ;
        RECT 53.020 102.100 53.310 102.145 ;
        RECT 51.120 101.960 53.310 102.100 ;
        RECT 38.255 101.915 38.545 101.960 ;
        RECT 51.120 101.900 51.440 101.960 ;
        RECT 53.020 101.915 53.310 101.960 ;
        RECT 54.355 101.915 54.645 102.145 ;
        RECT 73.660 102.100 73.980 102.160 ;
        RECT 76.050 102.145 76.190 102.640 ;
        RECT 80.100 102.580 80.420 102.640 ;
        RECT 86.555 102.780 86.845 102.825 ;
        RECT 87.000 102.780 87.320 102.840 ;
        RECT 86.555 102.640 87.320 102.780 ;
        RECT 86.555 102.595 86.845 102.640 ;
        RECT 87.000 102.580 87.320 102.640 ;
        RECT 104.940 102.780 105.260 102.840 ;
        RECT 105.415 102.780 105.705 102.825 ;
        RECT 112.760 102.780 113.080 102.840 ;
        RECT 114.140 102.780 114.460 102.840 ;
        RECT 118.280 102.780 118.600 102.840 ;
        RECT 104.940 102.640 110.230 102.780 ;
        RECT 104.940 102.580 105.260 102.640 ;
        RECT 105.415 102.595 105.705 102.640 ;
        RECT 77.815 102.440 78.105 102.485 ;
        RECT 76.510 102.300 78.105 102.440 ;
        RECT 76.510 102.145 76.650 102.300 ;
        RECT 77.815 102.255 78.105 102.300 ;
        RECT 79.655 102.440 79.945 102.485 ;
        RECT 81.020 102.440 81.340 102.500 ;
        RECT 79.655 102.300 81.340 102.440 ;
        RECT 79.655 102.255 79.945 102.300 ;
        RECT 81.020 102.240 81.340 102.300 ;
        RECT 82.875 102.440 83.165 102.485 ;
        RECT 92.980 102.440 93.300 102.500 ;
        RECT 82.875 102.300 86.770 102.440 ;
        RECT 82.875 102.255 83.165 102.300 ;
        RECT 86.630 102.160 86.770 102.300 ;
        RECT 88.930 102.300 93.300 102.440 ;
        RECT 75.515 102.100 75.805 102.145 ;
        RECT 73.660 101.960 75.805 102.100 ;
        RECT 73.660 101.900 73.980 101.960 ;
        RECT 75.515 101.915 75.805 101.960 ;
        RECT 75.975 101.915 76.265 102.145 ;
        RECT 76.435 101.915 76.725 102.145 ;
        RECT 77.355 101.915 77.645 102.145 ;
        RECT 78.260 102.100 78.580 102.160 ;
        RECT 78.735 102.100 79.025 102.145 ;
        RECT 78.260 101.960 79.025 102.100 ;
        RECT 49.765 101.760 50.055 101.805 ;
        RECT 52.285 101.760 52.575 101.805 ;
        RECT 53.475 101.760 53.765 101.805 ;
        RECT 28.210 101.620 29.270 101.760 ;
        RECT 24.005 101.575 24.295 101.620 ;
        RECT 26.525 101.575 26.815 101.620 ;
        RECT 27.715 101.575 28.005 101.620 ;
        RECT 18.015 101.420 18.305 101.465 ;
        RECT 19.855 101.420 20.145 101.465 ;
        RECT 20.300 101.420 20.620 101.480 ;
        RECT 18.015 101.280 19.610 101.420 ;
        RECT 18.015 101.235 18.305 101.280 ;
        RECT 18.920 100.880 19.240 101.140 ;
        RECT 19.470 101.080 19.610 101.280 ;
        RECT 19.855 101.280 20.620 101.420 ;
        RECT 19.855 101.235 20.145 101.280 ;
        RECT 20.300 101.220 20.620 101.280 ;
        RECT 20.760 101.420 21.080 101.480 ;
        RECT 29.130 101.465 29.270 101.620 ;
        RECT 49.765 101.620 53.765 101.760 ;
        RECT 75.590 101.760 75.730 101.915 ;
        RECT 75.590 101.620 76.190 101.760 ;
        RECT 49.765 101.575 50.055 101.620 ;
        RECT 52.285 101.575 52.575 101.620 ;
        RECT 53.475 101.575 53.765 101.620 ;
        RECT 21.695 101.420 21.985 101.465 ;
        RECT 20.760 101.280 21.985 101.420 ;
        RECT 20.760 101.220 21.080 101.280 ;
        RECT 21.695 101.235 21.985 101.280 ;
        RECT 24.440 101.420 24.730 101.465 ;
        RECT 26.010 101.420 26.300 101.465 ;
        RECT 28.110 101.420 28.400 101.465 ;
        RECT 24.440 101.280 28.400 101.420 ;
        RECT 24.440 101.235 24.730 101.280 ;
        RECT 26.010 101.235 26.300 101.280 ;
        RECT 28.110 101.235 28.400 101.280 ;
        RECT 29.055 101.235 29.345 101.465 ;
        RECT 30.880 101.420 31.200 101.480 ;
        RECT 29.590 101.280 31.200 101.420 ;
        RECT 29.590 101.080 29.730 101.280 ;
        RECT 30.880 101.220 31.200 101.280 ;
        RECT 47.440 101.220 47.760 101.480 ;
        RECT 50.200 101.420 50.490 101.465 ;
        RECT 51.770 101.420 52.060 101.465 ;
        RECT 53.870 101.420 54.160 101.465 ;
        RECT 50.200 101.280 54.160 101.420 ;
        RECT 50.200 101.235 50.490 101.280 ;
        RECT 51.770 101.235 52.060 101.280 ;
        RECT 53.870 101.235 54.160 101.280 ;
        RECT 19.470 100.940 29.730 101.080 ;
        RECT 29.960 100.880 30.280 101.140 ;
        RECT 36.400 100.880 36.720 101.140 ;
        RECT 40.555 101.080 40.845 101.125 ;
        RECT 41.000 101.080 41.320 101.140 ;
        RECT 40.555 100.940 41.320 101.080 ;
        RECT 40.555 100.895 40.845 100.940 ;
        RECT 41.000 100.880 41.320 100.940 ;
        RECT 74.120 100.880 74.440 101.140 ;
        RECT 76.050 101.080 76.190 101.620 ;
        RECT 77.430 101.420 77.570 101.915 ;
        RECT 78.260 101.900 78.580 101.960 ;
        RECT 78.735 101.915 79.025 101.960 ;
        RECT 83.320 102.100 83.640 102.160 ;
        RECT 83.795 102.100 84.085 102.145 ;
        RECT 83.320 101.960 84.085 102.100 ;
        RECT 83.320 101.900 83.640 101.960 ;
        RECT 83.795 101.915 84.085 101.960 ;
        RECT 84.255 101.915 84.545 102.145 ;
        RECT 81.020 101.760 81.340 101.820 ;
        RECT 84.330 101.760 84.470 101.915 ;
        RECT 85.160 101.900 85.480 102.160 ;
        RECT 85.635 102.100 85.925 102.145 ;
        RECT 85.635 101.960 86.310 102.100 ;
        RECT 85.635 101.915 85.925 101.960 ;
        RECT 81.020 101.620 84.470 101.760 ;
        RECT 81.020 101.560 81.340 101.620 ;
        RECT 78.720 101.420 79.040 101.480 ;
        RECT 77.430 101.280 79.040 101.420 ;
        RECT 78.720 101.220 79.040 101.280 ;
        RECT 84.700 101.080 85.020 101.140 ;
        RECT 76.050 100.940 85.020 101.080 ;
        RECT 86.170 101.080 86.310 101.960 ;
        RECT 86.540 101.900 86.860 102.160 ;
        RECT 87.920 101.900 88.240 102.160 ;
        RECT 88.930 102.145 89.070 102.300 ;
        RECT 92.980 102.240 93.300 102.300 ;
        RECT 98.960 102.440 99.280 102.500 ;
        RECT 109.555 102.440 109.845 102.485 ;
        RECT 98.960 102.300 109.845 102.440 ;
        RECT 98.960 102.240 99.280 102.300 ;
        RECT 109.555 102.255 109.845 102.300 ;
        RECT 88.395 101.915 88.685 102.145 ;
        RECT 88.855 101.915 89.145 102.145 ;
        RECT 87.000 101.760 87.320 101.820 ;
        RECT 88.470 101.760 88.610 101.915 ;
        RECT 89.760 101.900 90.080 102.160 ;
        RECT 98.040 102.100 98.360 102.160 ;
        RECT 99.795 102.100 100.085 102.145 ;
        RECT 98.040 101.960 100.085 102.100 ;
        RECT 98.040 101.900 98.360 101.960 ;
        RECT 99.795 101.915 100.085 101.960 ;
        RECT 108.620 101.900 108.940 102.160 ;
        RECT 109.080 101.900 109.400 102.160 ;
        RECT 87.000 101.620 88.610 101.760 ;
        RECT 87.000 101.560 87.320 101.620 ;
        RECT 98.500 101.560 98.820 101.820 ;
        RECT 99.395 101.760 99.685 101.805 ;
        RECT 100.585 101.760 100.875 101.805 ;
        RECT 103.105 101.760 103.395 101.805 ;
        RECT 99.395 101.620 103.395 101.760 ;
        RECT 99.395 101.575 99.685 101.620 ;
        RECT 100.585 101.575 100.875 101.620 ;
        RECT 103.105 101.575 103.395 101.620 ;
        RECT 99.000 101.420 99.290 101.465 ;
        RECT 101.100 101.420 101.390 101.465 ;
        RECT 102.670 101.420 102.960 101.465 ;
        RECT 109.630 101.420 109.770 102.255 ;
        RECT 110.090 102.160 110.230 102.640 ;
        RECT 112.760 102.640 114.460 102.780 ;
        RECT 112.760 102.580 113.080 102.640 ;
        RECT 114.140 102.580 114.460 102.640 ;
        RECT 114.690 102.640 118.600 102.780 ;
        RECT 111.840 102.440 112.160 102.500 ;
        RECT 114.690 102.440 114.830 102.640 ;
        RECT 118.280 102.580 118.600 102.640 ;
        RECT 127.955 102.780 128.245 102.825 ;
        RECT 134.380 102.780 134.700 102.840 ;
        RECT 135.315 102.780 135.605 102.825 ;
        RECT 127.955 102.640 129.090 102.780 ;
        RECT 127.955 102.595 128.245 102.640 ;
        RECT 118.740 102.440 119.060 102.500 ;
        RECT 124.260 102.440 124.580 102.500 ;
        RECT 128.950 102.440 129.090 102.640 ;
        RECT 134.380 102.640 135.605 102.780 ;
        RECT 134.380 102.580 134.700 102.640 ;
        RECT 135.315 102.595 135.605 102.640 ;
        RECT 129.640 102.440 129.930 102.485 ;
        RECT 111.840 102.300 114.830 102.440 ;
        RECT 111.840 102.240 112.160 102.300 ;
        RECT 110.000 102.100 110.320 102.160 ;
        RECT 110.475 102.100 110.765 102.145 ;
        RECT 110.000 101.960 110.765 102.100 ;
        RECT 110.000 101.900 110.320 101.960 ;
        RECT 110.475 101.915 110.765 101.960 ;
        RECT 114.140 101.900 114.460 102.160 ;
        RECT 114.690 102.145 114.830 102.300 ;
        RECT 116.990 102.300 128.630 102.440 ;
        RECT 128.950 102.300 129.930 102.440 ;
        RECT 114.615 101.915 114.905 102.145 ;
        RECT 115.060 101.900 115.380 102.160 ;
        RECT 115.995 102.100 116.285 102.145 ;
        RECT 116.440 102.100 116.760 102.160 ;
        RECT 116.990 102.145 117.130 102.300 ;
        RECT 118.740 102.240 119.060 102.300 ;
        RECT 124.260 102.240 124.580 102.300 ;
        RECT 115.995 101.960 116.760 102.100 ;
        RECT 115.995 101.915 116.285 101.960 ;
        RECT 116.440 101.900 116.760 101.960 ;
        RECT 116.915 101.915 117.205 102.145 ;
        RECT 118.195 102.100 118.485 102.145 ;
        RECT 117.450 101.960 118.485 102.100 ;
        RECT 112.775 101.760 113.065 101.805 ;
        RECT 117.450 101.760 117.590 101.960 ;
        RECT 118.195 101.915 118.485 101.960 ;
        RECT 122.880 102.100 123.200 102.160 ;
        RECT 124.735 102.100 125.025 102.145 ;
        RECT 122.880 101.960 125.025 102.100 ;
        RECT 122.880 101.900 123.200 101.960 ;
        RECT 124.735 101.915 125.025 101.960 ;
        RECT 125.180 102.100 125.500 102.160 ;
        RECT 125.655 102.100 125.945 102.145 ;
        RECT 125.180 101.960 125.945 102.100 ;
        RECT 125.180 101.900 125.500 101.960 ;
        RECT 125.655 101.915 125.945 101.960 ;
        RECT 126.115 101.915 126.405 102.145 ;
        RECT 126.575 102.100 126.865 102.145 ;
        RECT 127.020 102.100 127.340 102.160 ;
        RECT 128.490 102.145 128.630 102.300 ;
        RECT 129.640 102.255 129.930 102.300 ;
        RECT 126.575 101.960 127.340 102.100 ;
        RECT 126.575 101.915 126.865 101.960 ;
        RECT 112.775 101.620 117.590 101.760 ;
        RECT 117.795 101.760 118.085 101.805 ;
        RECT 118.985 101.760 119.275 101.805 ;
        RECT 121.505 101.760 121.795 101.805 ;
        RECT 117.795 101.620 121.795 101.760 ;
        RECT 112.775 101.575 113.065 101.620 ;
        RECT 117.795 101.575 118.085 101.620 ;
        RECT 118.985 101.575 119.275 101.620 ;
        RECT 121.505 101.575 121.795 101.620 ;
        RECT 123.800 101.760 124.120 101.820 ;
        RECT 126.190 101.760 126.330 101.915 ;
        RECT 127.020 101.900 127.340 101.960 ;
        RECT 128.415 101.915 128.705 102.145 ;
        RECT 135.390 102.100 135.530 102.595 ;
        RECT 136.680 102.580 137.000 102.840 ;
        RECT 135.775 102.100 136.065 102.145 ;
        RECT 135.390 101.960 136.065 102.100 ;
        RECT 135.775 101.915 136.065 101.960 ;
        RECT 129.295 101.760 129.585 101.805 ;
        RECT 130.485 101.760 130.775 101.805 ;
        RECT 133.005 101.760 133.295 101.805 ;
        RECT 123.800 101.620 127.250 101.760 ;
        RECT 123.800 101.560 124.120 101.620 ;
        RECT 127.110 101.480 127.250 101.620 ;
        RECT 129.295 101.620 133.295 101.760 ;
        RECT 129.295 101.575 129.585 101.620 ;
        RECT 130.485 101.575 130.775 101.620 ;
        RECT 133.005 101.575 133.295 101.620 ;
        RECT 110.460 101.420 110.780 101.480 ;
        RECT 99.000 101.280 102.960 101.420 ;
        RECT 99.000 101.235 99.290 101.280 ;
        RECT 101.100 101.235 101.390 101.280 ;
        RECT 102.670 101.235 102.960 101.280 ;
        RECT 107.330 101.280 108.390 101.420 ;
        RECT 109.630 101.280 110.780 101.420 ;
        RECT 107.330 101.080 107.470 101.280 ;
        RECT 86.170 100.940 107.470 101.080 ;
        RECT 84.700 100.880 85.020 100.940 ;
        RECT 107.700 100.880 108.020 101.140 ;
        RECT 108.250 101.080 108.390 101.280 ;
        RECT 110.460 101.220 110.780 101.280 ;
        RECT 117.400 101.420 117.690 101.465 ;
        RECT 119.500 101.420 119.790 101.465 ;
        RECT 121.070 101.420 121.360 101.465 ;
        RECT 126.100 101.420 126.420 101.480 ;
        RECT 117.400 101.280 121.360 101.420 ;
        RECT 117.400 101.235 117.690 101.280 ;
        RECT 119.500 101.235 119.790 101.280 ;
        RECT 121.070 101.235 121.360 101.280 ;
        RECT 123.430 101.280 126.420 101.420 ;
        RECT 123.430 101.080 123.570 101.280 ;
        RECT 126.100 101.220 126.420 101.280 ;
        RECT 127.020 101.220 127.340 101.480 ;
        RECT 128.900 101.420 129.190 101.465 ;
        RECT 131.000 101.420 131.290 101.465 ;
        RECT 132.570 101.420 132.860 101.465 ;
        RECT 128.900 101.280 132.860 101.420 ;
        RECT 128.900 101.235 129.190 101.280 ;
        RECT 131.000 101.235 131.290 101.280 ;
        RECT 132.570 101.235 132.860 101.280 ;
        RECT 108.250 100.940 123.570 101.080 ;
        RECT 123.800 100.880 124.120 101.140 ;
        RECT 13.330 100.260 138.910 100.740 ;
        RECT 21.680 100.060 22.000 100.120 ;
        RECT 25.375 100.060 25.665 100.105 ;
        RECT 21.680 99.920 25.665 100.060 ;
        RECT 21.680 99.860 22.000 99.920 ;
        RECT 25.375 99.875 25.665 99.920 ;
        RECT 49.295 100.060 49.585 100.105 ;
        RECT 49.740 100.060 50.060 100.120 ;
        RECT 49.295 99.920 50.060 100.060 ;
        RECT 49.295 99.875 49.585 99.920 ;
        RECT 49.740 99.860 50.060 99.920 ;
        RECT 76.880 100.060 77.200 100.120 ;
        RECT 81.020 100.060 81.340 100.120 ;
        RECT 76.880 99.920 81.340 100.060 ;
        RECT 76.880 99.860 77.200 99.920 ;
        RECT 81.020 99.860 81.340 99.920 ;
        RECT 81.480 100.060 81.800 100.120 ;
        RECT 83.335 100.060 83.625 100.105 ;
        RECT 81.480 99.920 83.625 100.060 ;
        RECT 81.480 99.860 81.800 99.920 ;
        RECT 83.335 99.875 83.625 99.920 ;
        RECT 85.160 100.060 85.480 100.120 ;
        RECT 87.015 100.060 87.305 100.105 ;
        RECT 85.160 99.920 87.305 100.060 ;
        RECT 85.160 99.860 85.480 99.920 ;
        RECT 87.015 99.875 87.305 99.920 ;
        RECT 98.040 99.860 98.360 100.120 ;
        RECT 102.180 99.860 102.500 100.120 ;
        RECT 112.760 100.060 113.080 100.120 ;
        RECT 102.730 99.920 113.080 100.060 ;
        RECT 18.960 99.720 19.250 99.765 ;
        RECT 21.060 99.720 21.350 99.765 ;
        RECT 22.630 99.720 22.920 99.765 ;
        RECT 18.960 99.580 22.920 99.720 ;
        RECT 18.960 99.535 19.250 99.580 ;
        RECT 21.060 99.535 21.350 99.580 ;
        RECT 22.630 99.535 22.920 99.580 ;
        RECT 70.940 99.720 71.230 99.765 ;
        RECT 73.040 99.720 73.330 99.765 ;
        RECT 74.610 99.720 74.900 99.765 ;
        RECT 99.420 99.720 99.740 99.780 ;
        RECT 102.730 99.720 102.870 99.920 ;
        RECT 112.760 99.860 113.080 99.920 ;
        RECT 115.060 100.060 115.380 100.120 ;
        RECT 115.995 100.060 116.285 100.105 ;
        RECT 115.060 99.920 116.285 100.060 ;
        RECT 115.060 99.860 115.380 99.920 ;
        RECT 115.995 99.875 116.285 99.920 ;
        RECT 116.440 100.060 116.760 100.120 ;
        RECT 117.375 100.060 117.665 100.105 ;
        RECT 116.440 99.920 117.665 100.060 ;
        RECT 116.440 99.860 116.760 99.920 ;
        RECT 117.375 99.875 117.665 99.920 ;
        RECT 135.300 100.060 135.620 100.120 ;
        RECT 136.695 100.060 136.985 100.105 ;
        RECT 135.300 99.920 136.985 100.060 ;
        RECT 135.300 99.860 135.620 99.920 ;
        RECT 136.695 99.875 136.985 99.920 ;
        RECT 116.900 99.720 117.220 99.780 ;
        RECT 70.940 99.580 74.900 99.720 ;
        RECT 70.940 99.535 71.230 99.580 ;
        RECT 73.040 99.535 73.330 99.580 ;
        RECT 74.610 99.535 74.900 99.580 ;
        RECT 99.050 99.580 102.870 99.720 ;
        RECT 104.570 99.580 117.220 99.720 ;
        RECT 17.540 99.380 17.860 99.440 ;
        RECT 18.475 99.380 18.765 99.425 ;
        RECT 17.540 99.240 18.765 99.380 ;
        RECT 17.540 99.180 17.860 99.240 ;
        RECT 18.475 99.195 18.765 99.240 ;
        RECT 19.355 99.380 19.645 99.425 ;
        RECT 20.545 99.380 20.835 99.425 ;
        RECT 23.065 99.380 23.355 99.425 ;
        RECT 50.200 99.380 50.520 99.440 ;
        RECT 19.355 99.240 23.355 99.380 ;
        RECT 19.355 99.195 19.645 99.240 ;
        RECT 20.545 99.195 20.835 99.240 ;
        RECT 23.065 99.195 23.355 99.240 ;
        RECT 48.910 99.240 50.520 99.380 ;
        RECT 18.920 99.040 19.240 99.100 ;
        RECT 48.910 99.085 49.050 99.240 ;
        RECT 50.200 99.180 50.520 99.240 ;
        RECT 71.335 99.380 71.625 99.425 ;
        RECT 72.525 99.380 72.815 99.425 ;
        RECT 75.045 99.380 75.335 99.425 ;
        RECT 91.600 99.380 91.920 99.440 ;
        RECT 71.335 99.240 75.335 99.380 ;
        RECT 71.335 99.195 71.625 99.240 ;
        RECT 72.525 99.195 72.815 99.240 ;
        RECT 75.045 99.195 75.335 99.240 ;
        RECT 88.010 99.240 91.920 99.380 ;
        RECT 88.010 99.100 88.150 99.240 ;
        RECT 91.600 99.180 91.920 99.240 ;
        RECT 19.755 99.040 20.045 99.085 ;
        RECT 18.920 98.900 20.045 99.040 ;
        RECT 18.920 98.840 19.240 98.900 ;
        RECT 19.755 98.855 20.045 98.900 ;
        RECT 48.835 98.855 49.125 99.085 ;
        RECT 49.280 99.040 49.600 99.100 ;
        RECT 49.755 99.040 50.045 99.085 ;
        RECT 49.280 98.900 50.045 99.040 ;
        RECT 49.280 98.840 49.600 98.900 ;
        RECT 49.755 98.855 50.045 98.900 ;
        RECT 70.440 98.840 70.760 99.100 ;
        RECT 71.790 99.040 72.080 99.085 ;
        RECT 74.120 99.040 74.440 99.100 ;
        RECT 71.790 98.900 74.440 99.040 ;
        RECT 71.790 98.855 72.080 98.900 ;
        RECT 74.120 98.840 74.440 98.900 ;
        RECT 79.640 98.840 79.960 99.100 ;
        RECT 80.100 98.840 80.420 99.100 ;
        RECT 80.560 98.840 80.880 99.100 ;
        RECT 81.480 98.840 81.800 99.100 ;
        RECT 82.415 98.855 82.705 99.085 ;
        RECT 82.490 98.700 82.630 98.855 ;
        RECT 87.920 98.840 88.240 99.100 ;
        RECT 89.775 99.040 90.065 99.085 ;
        RECT 97.580 99.040 97.900 99.100 ;
        RECT 89.775 98.900 97.900 99.040 ;
        RECT 99.050 99.040 99.190 99.580 ;
        RECT 99.420 99.520 99.740 99.580 ;
        RECT 99.335 99.040 99.625 99.085 ;
        RECT 99.050 98.900 99.625 99.040 ;
        RECT 89.775 98.855 90.065 98.900 ;
        RECT 97.580 98.840 97.900 98.900 ;
        RECT 99.335 98.855 99.625 98.900 ;
        RECT 99.895 98.855 100.185 99.085 ;
        RECT 100.355 98.855 100.645 99.085 ;
        RECT 101.275 99.040 101.565 99.085 ;
        RECT 102.180 99.040 102.500 99.100 ;
        RECT 101.275 98.900 102.500 99.040 ;
        RECT 101.275 98.855 101.565 98.900 ;
        RECT 71.910 98.560 82.630 98.700 ;
        RECT 71.910 98.420 72.050 98.560 ;
        RECT 71.820 98.160 72.140 98.420 ;
        RECT 77.355 98.360 77.645 98.405 ;
        RECT 77.800 98.360 78.120 98.420 ;
        RECT 77.355 98.220 78.120 98.360 ;
        RECT 77.355 98.175 77.645 98.220 ;
        RECT 77.800 98.160 78.120 98.220 ;
        RECT 78.260 98.160 78.580 98.420 ;
        RECT 82.490 98.360 82.630 98.560 ;
        RECT 88.380 98.500 88.700 98.760 ;
        RECT 88.840 98.500 89.160 98.760 ;
        RECT 96.200 98.700 96.520 98.760 ;
        RECT 99.970 98.700 100.110 98.855 ;
        RECT 96.200 98.560 100.110 98.700 ;
        RECT 100.430 98.700 100.570 98.855 ;
        RECT 102.180 98.840 102.500 98.900 ;
        RECT 102.640 99.040 102.960 99.100 ;
        RECT 103.115 99.040 103.405 99.085 ;
        RECT 104.570 99.040 104.710 99.580 ;
        RECT 116.900 99.520 117.220 99.580 ;
        RECT 130.280 99.720 130.570 99.765 ;
        RECT 132.380 99.720 132.670 99.765 ;
        RECT 133.950 99.720 134.240 99.765 ;
        RECT 130.280 99.580 134.240 99.720 ;
        RECT 130.280 99.535 130.570 99.580 ;
        RECT 132.380 99.535 132.670 99.580 ;
        RECT 133.950 99.535 134.240 99.580 ;
        RECT 123.800 99.380 124.120 99.440 ;
        RECT 115.150 99.240 124.120 99.380 ;
        RECT 102.640 98.900 104.710 99.040 ;
        RECT 102.640 98.840 102.960 98.900 ;
        RECT 103.115 98.855 103.405 98.900 ;
        RECT 104.940 98.840 105.260 99.100 ;
        RECT 109.080 99.040 109.400 99.100 ;
        RECT 115.150 99.085 115.290 99.240 ;
        RECT 123.800 99.180 124.120 99.240 ;
        RECT 124.260 99.380 124.580 99.440 ;
        RECT 129.795 99.380 130.085 99.425 ;
        RECT 124.260 99.240 130.085 99.380 ;
        RECT 124.260 99.180 124.580 99.240 ;
        RECT 129.795 99.195 130.085 99.240 ;
        RECT 130.675 99.380 130.965 99.425 ;
        RECT 131.865 99.380 132.155 99.425 ;
        RECT 134.385 99.380 134.675 99.425 ;
        RECT 130.675 99.240 134.675 99.380 ;
        RECT 130.675 99.195 130.965 99.240 ;
        RECT 131.865 99.195 132.155 99.240 ;
        RECT 134.385 99.195 134.675 99.240 ;
        RECT 115.075 99.040 115.365 99.085 ;
        RECT 109.080 98.900 115.365 99.040 ;
        RECT 109.080 98.840 109.400 98.900 ;
        RECT 115.075 98.855 115.365 98.900 ;
        RECT 115.980 99.040 116.300 99.100 ;
        RECT 116.455 99.040 116.745 99.085 ;
        RECT 115.980 98.900 116.745 99.040 ;
        RECT 115.980 98.840 116.300 98.900 ;
        RECT 116.455 98.855 116.745 98.900 ;
        RECT 122.880 99.040 123.200 99.100 ;
        RECT 125.655 99.040 125.945 99.085 ;
        RECT 122.880 98.900 125.945 99.040 ;
        RECT 122.880 98.840 123.200 98.900 ;
        RECT 104.035 98.700 104.325 98.745 ;
        RECT 100.430 98.560 104.325 98.700 ;
        RECT 96.200 98.500 96.520 98.560 ;
        RECT 92.980 98.360 93.300 98.420 ;
        RECT 82.490 98.220 93.300 98.360 ;
        RECT 99.970 98.360 100.110 98.560 ;
        RECT 104.035 98.515 104.325 98.560 ;
        RECT 105.400 98.700 105.720 98.760 ;
        RECT 105.875 98.700 106.165 98.745 ;
        RECT 105.400 98.560 106.165 98.700 ;
        RECT 105.400 98.500 105.720 98.560 ;
        RECT 105.875 98.515 106.165 98.560 ;
        RECT 114.155 98.700 114.445 98.745 ;
        RECT 115.520 98.700 115.840 98.760 ;
        RECT 114.155 98.560 115.840 98.700 ;
        RECT 114.155 98.515 114.445 98.560 ;
        RECT 115.520 98.500 115.840 98.560 ;
        RECT 104.940 98.360 105.260 98.420 ;
        RECT 99.970 98.220 105.260 98.360 ;
        RECT 92.980 98.160 93.300 98.220 ;
        RECT 104.940 98.160 105.260 98.220 ;
        RECT 116.440 98.360 116.760 98.420 ;
        RECT 122.970 98.360 123.110 98.840 ;
        RECT 124.350 98.760 124.490 98.900 ;
        RECT 125.655 98.855 125.945 98.900 ;
        RECT 126.560 98.840 126.880 99.100 ;
        RECT 127.020 98.840 127.340 99.100 ;
        RECT 127.495 99.040 127.785 99.085 ;
        RECT 128.400 99.040 128.720 99.100 ;
        RECT 127.495 98.900 128.720 99.040 ;
        RECT 129.870 99.040 130.010 99.195 ;
        RECT 129.870 98.900 132.310 99.040 ;
        RECT 127.495 98.855 127.785 98.900 ;
        RECT 128.400 98.840 128.720 98.900 ;
        RECT 124.260 98.500 124.580 98.760 ;
        RECT 116.440 98.220 123.110 98.360 ;
        RECT 123.340 98.360 123.660 98.420 ;
        RECT 127.110 98.360 127.250 98.840 ;
        RECT 132.170 98.760 132.310 98.900 ;
        RECT 128.875 98.700 129.165 98.745 ;
        RECT 131.020 98.700 131.310 98.745 ;
        RECT 128.875 98.560 131.310 98.700 ;
        RECT 128.875 98.515 129.165 98.560 ;
        RECT 131.020 98.515 131.310 98.560 ;
        RECT 132.080 98.500 132.400 98.760 ;
        RECT 131.620 98.360 131.940 98.420 ;
        RECT 123.340 98.220 131.940 98.360 ;
        RECT 116.440 98.160 116.760 98.220 ;
        RECT 123.340 98.160 123.660 98.220 ;
        RECT 131.620 98.160 131.940 98.220 ;
        RECT 13.330 97.540 138.910 98.020 ;
        RECT 81.480 97.140 81.800 97.400 ;
        RECT 94.820 97.340 95.140 97.400 ;
        RECT 91.230 97.200 95.140 97.340 ;
        RECT 81.570 97.000 81.710 97.140 ;
        RECT 91.230 97.045 91.370 97.200 ;
        RECT 94.820 97.140 95.140 97.200 ;
        RECT 105.860 97.140 106.180 97.400 ;
        RECT 108.620 97.340 108.940 97.400 ;
        RECT 115.520 97.340 115.840 97.400 ;
        RECT 108.620 97.200 111.150 97.340 ;
        RECT 108.620 97.140 108.940 97.200 ;
        RECT 81.570 96.860 90.450 97.000 ;
        RECT 72.250 96.660 72.540 96.705 ;
        RECT 78.260 96.660 78.580 96.720 ;
        RECT 72.250 96.520 78.580 96.660 ;
        RECT 72.250 96.475 72.540 96.520 ;
        RECT 78.260 96.460 78.580 96.520 ;
        RECT 79.640 96.660 79.960 96.720 ;
        RECT 82.950 96.705 83.090 96.860 ;
        RECT 81.035 96.660 81.325 96.705 ;
        RECT 79.640 96.520 81.325 96.660 ;
        RECT 79.640 96.460 79.960 96.520 ;
        RECT 81.035 96.475 81.325 96.520 ;
        RECT 81.495 96.475 81.785 96.705 ;
        RECT 81.955 96.475 82.245 96.705 ;
        RECT 82.875 96.475 83.165 96.705 ;
        RECT 70.440 96.320 70.760 96.380 ;
        RECT 70.915 96.320 71.205 96.365 ;
        RECT 70.440 96.180 71.205 96.320 ;
        RECT 70.440 96.120 70.760 96.180 ;
        RECT 70.915 96.135 71.205 96.180 ;
        RECT 71.795 96.320 72.085 96.365 ;
        RECT 72.985 96.320 73.275 96.365 ;
        RECT 75.505 96.320 75.795 96.365 ;
        RECT 71.795 96.180 75.795 96.320 ;
        RECT 71.795 96.135 72.085 96.180 ;
        RECT 72.985 96.135 73.275 96.180 ;
        RECT 75.505 96.135 75.795 96.180 ;
        RECT 70.990 95.640 71.130 96.135 ;
        RECT 71.400 95.980 71.690 96.025 ;
        RECT 73.500 95.980 73.790 96.025 ;
        RECT 75.070 95.980 75.360 96.025 ;
        RECT 71.400 95.840 75.360 95.980 ;
        RECT 81.570 95.980 81.710 96.475 ;
        RECT 82.030 96.320 82.170 96.475 ;
        RECT 84.700 96.460 85.020 96.720 ;
        RECT 85.175 96.475 85.465 96.705 ;
        RECT 84.240 96.320 84.560 96.380 ;
        RECT 82.030 96.180 84.560 96.320 ;
        RECT 84.240 96.120 84.560 96.180 ;
        RECT 85.250 96.320 85.390 96.475 ;
        RECT 85.620 96.460 85.940 96.720 ;
        RECT 86.630 96.705 86.770 96.860 ;
        RECT 86.555 96.475 86.845 96.705 ;
        RECT 87.000 96.460 87.320 96.720 ;
        RECT 87.920 96.460 88.240 96.720 ;
        RECT 88.395 96.475 88.685 96.705 ;
        RECT 87.090 96.320 87.230 96.460 ;
        RECT 85.250 96.180 87.230 96.320 ;
        RECT 87.460 96.320 87.780 96.380 ;
        RECT 88.470 96.320 88.610 96.475 ;
        RECT 88.840 96.460 89.160 96.720 ;
        RECT 89.760 96.460 90.080 96.720 ;
        RECT 87.460 96.180 88.610 96.320 ;
        RECT 90.310 96.320 90.450 96.860 ;
        RECT 91.155 96.815 91.445 97.045 ;
        RECT 91.600 97.000 91.920 97.060 ;
        RECT 92.995 97.000 93.285 97.045 ;
        RECT 91.600 96.860 93.285 97.000 ;
        RECT 91.600 96.800 91.920 96.860 ;
        RECT 92.995 96.815 93.285 96.860 ;
        RECT 102.180 97.000 102.500 97.060 ;
        RECT 106.780 97.000 107.100 97.060 ;
        RECT 102.180 96.860 109.310 97.000 ;
        RECT 102.180 96.800 102.500 96.860 ;
        RECT 106.780 96.800 107.100 96.860 ;
        RECT 92.075 96.660 92.365 96.705 ;
        RECT 92.520 96.660 92.840 96.720 ;
        RECT 92.075 96.520 92.840 96.660 ;
        RECT 92.075 96.475 92.365 96.520 ;
        RECT 92.520 96.460 92.840 96.520 ;
        RECT 93.455 96.475 93.745 96.705 ;
        RECT 93.530 96.320 93.670 96.475 ;
        RECT 94.360 96.460 94.680 96.720 ;
        RECT 94.835 96.475 95.125 96.705 ;
        RECT 90.310 96.180 93.670 96.320 ;
        RECT 94.910 96.320 95.050 96.475 ;
        RECT 95.280 96.460 95.600 96.720 ;
        RECT 98.500 96.460 98.820 96.720 ;
        RECT 99.850 96.660 100.140 96.705 ;
        RECT 104.020 96.660 104.340 96.720 ;
        RECT 107.255 96.660 107.545 96.705 ;
        RECT 99.850 96.520 104.340 96.660 ;
        RECT 99.850 96.475 100.140 96.520 ;
        RECT 104.020 96.460 104.340 96.520 ;
        RECT 104.570 96.520 107.545 96.660 ;
        RECT 96.200 96.320 96.520 96.380 ;
        RECT 94.910 96.180 96.520 96.320 ;
        RECT 85.250 95.980 85.390 96.180 ;
        RECT 87.460 96.120 87.780 96.180 ;
        RECT 81.570 95.840 85.390 95.980 ;
        RECT 71.400 95.795 71.690 95.840 ;
        RECT 73.500 95.795 73.790 95.840 ;
        RECT 75.070 95.795 75.360 95.840 ;
        RECT 76.420 95.640 76.740 95.700 ;
        RECT 70.990 95.500 76.740 95.640 ;
        RECT 76.420 95.440 76.740 95.500 ;
        RECT 76.880 95.640 77.200 95.700 ;
        RECT 77.815 95.640 78.105 95.685 ;
        RECT 76.880 95.500 78.105 95.640 ;
        RECT 76.880 95.440 77.200 95.500 ;
        RECT 77.815 95.455 78.105 95.500 ;
        RECT 79.640 95.440 79.960 95.700 ;
        RECT 83.320 95.440 83.640 95.700 ;
        RECT 85.250 95.640 85.390 95.840 ;
        RECT 86.080 95.980 86.400 96.040 ;
        RECT 87.015 95.980 87.305 96.025 ;
        RECT 90.680 95.980 91.000 96.040 ;
        RECT 94.910 95.980 95.050 96.180 ;
        RECT 96.200 96.120 96.520 96.180 ;
        RECT 99.395 96.320 99.685 96.365 ;
        RECT 100.585 96.320 100.875 96.365 ;
        RECT 103.105 96.320 103.395 96.365 ;
        RECT 99.395 96.180 103.395 96.320 ;
        RECT 99.395 96.135 99.685 96.180 ;
        RECT 100.585 96.135 100.875 96.180 ;
        RECT 103.105 96.135 103.395 96.180 ;
        RECT 99.000 95.980 99.290 96.025 ;
        RECT 101.100 95.980 101.390 96.025 ;
        RECT 102.670 95.980 102.960 96.025 ;
        RECT 86.080 95.840 87.305 95.980 ;
        RECT 86.080 95.780 86.400 95.840 ;
        RECT 87.015 95.795 87.305 95.840 ;
        RECT 89.850 95.840 95.050 95.980 ;
        RECT 96.290 95.840 98.730 95.980 ;
        RECT 89.850 95.640 89.990 95.840 ;
        RECT 90.680 95.780 91.000 95.840 ;
        RECT 85.250 95.500 89.990 95.640 ;
        RECT 90.220 95.640 90.540 95.700 ;
        RECT 96.290 95.640 96.430 95.840 ;
        RECT 90.220 95.500 96.430 95.640 ;
        RECT 90.220 95.440 90.540 95.500 ;
        RECT 96.660 95.440 96.980 95.700 ;
        RECT 98.590 95.640 98.730 95.840 ;
        RECT 99.000 95.840 102.960 95.980 ;
        RECT 99.000 95.795 99.290 95.840 ;
        RECT 101.100 95.795 101.390 95.840 ;
        RECT 102.670 95.795 102.960 95.840 ;
        RECT 104.570 95.640 104.710 96.520 ;
        RECT 107.255 96.475 107.545 96.520 ;
        RECT 107.715 96.475 108.005 96.705 ;
        RECT 104.940 96.320 105.260 96.380 ;
        RECT 107.790 96.320 107.930 96.475 ;
        RECT 108.160 96.460 108.480 96.720 ;
        RECT 109.170 96.705 109.310 96.860 ;
        RECT 110.460 96.800 110.780 97.060 ;
        RECT 111.010 97.000 111.150 97.200 ;
        RECT 114.230 97.200 115.840 97.340 ;
        RECT 114.230 97.045 114.370 97.200 ;
        RECT 115.520 97.140 115.840 97.200 ;
        RECT 118.280 97.340 118.600 97.400 ;
        RECT 120.580 97.340 120.900 97.400 ;
        RECT 122.880 97.340 123.200 97.400 ;
        RECT 118.280 97.200 123.200 97.340 ;
        RECT 118.280 97.140 118.600 97.200 ;
        RECT 120.580 97.140 120.900 97.200 ;
        RECT 122.880 97.140 123.200 97.200 ;
        RECT 123.340 97.140 123.660 97.400 ;
        RECT 111.010 96.860 111.610 97.000 ;
        RECT 109.095 96.475 109.385 96.705 ;
        RECT 109.555 96.475 109.845 96.705 ;
        RECT 104.940 96.180 107.930 96.320 ;
        RECT 104.940 96.120 105.260 96.180 ;
        RECT 105.415 95.980 105.705 96.025 ;
        RECT 106.320 95.980 106.640 96.040 ;
        RECT 109.630 95.980 109.770 96.475 ;
        RECT 110.000 96.460 110.320 96.720 ;
        RECT 111.470 96.705 111.610 96.860 ;
        RECT 114.155 96.815 114.445 97.045 ;
        RECT 115.060 97.000 115.380 97.060 ;
        RECT 123.430 97.000 123.570 97.140 ;
        RECT 125.640 97.000 125.960 97.060 ;
        RECT 115.060 96.860 123.570 97.000 ;
        RECT 123.890 96.860 125.960 97.000 ;
        RECT 115.060 96.800 115.380 96.860 ;
        RECT 110.935 96.475 111.225 96.705 ;
        RECT 111.395 96.660 111.685 96.705 ;
        RECT 114.600 96.660 114.920 96.720 ;
        RECT 111.395 96.520 114.920 96.660 ;
        RECT 111.395 96.475 111.685 96.520 ;
        RECT 110.090 96.040 110.230 96.460 ;
        RECT 110.460 96.320 110.780 96.380 ;
        RECT 111.010 96.320 111.150 96.475 ;
        RECT 114.600 96.460 114.920 96.520 ;
        RECT 116.440 96.660 116.760 96.720 ;
        RECT 116.915 96.660 117.205 96.705 ;
        RECT 117.835 96.660 118.125 96.705 ;
        RECT 116.440 96.520 117.205 96.660 ;
        RECT 116.440 96.460 116.760 96.520 ;
        RECT 116.915 96.475 117.205 96.520 ;
        RECT 117.450 96.520 118.125 96.660 ;
        RECT 115.995 96.320 116.285 96.365 ;
        RECT 117.450 96.320 117.590 96.520 ;
        RECT 117.835 96.475 118.125 96.520 ;
        RECT 118.280 96.460 118.600 96.720 ;
        RECT 118.755 96.475 119.045 96.705 ;
        RECT 121.960 96.660 122.280 96.720 ;
        RECT 122.435 96.660 122.725 96.705 ;
        RECT 121.960 96.520 122.725 96.660 ;
        RECT 110.460 96.180 111.150 96.320 ;
        RECT 111.930 96.180 115.290 96.320 ;
        RECT 110.460 96.120 110.780 96.180 ;
        RECT 105.415 95.840 109.770 95.980 ;
        RECT 105.415 95.795 105.705 95.840 ;
        RECT 106.320 95.780 106.640 95.840 ;
        RECT 110.000 95.780 110.320 96.040 ;
        RECT 111.930 95.640 112.070 96.180 ;
        RECT 115.150 95.980 115.290 96.180 ;
        RECT 115.995 96.180 117.590 96.320 ;
        RECT 115.995 96.135 116.285 96.180 ;
        RECT 118.830 95.980 118.970 96.475 ;
        RECT 121.960 96.460 122.280 96.520 ;
        RECT 122.435 96.475 122.725 96.520 ;
        RECT 122.880 96.460 123.200 96.720 ;
        RECT 123.355 96.660 123.645 96.705 ;
        RECT 123.890 96.660 124.030 96.860 ;
        RECT 125.640 96.800 125.960 96.860 ;
        RECT 130.330 96.860 132.770 97.000 ;
        RECT 123.355 96.520 124.030 96.660 ;
        RECT 123.355 96.475 123.645 96.520 ;
        RECT 124.260 96.460 124.580 96.720 ;
        RECT 130.330 96.660 130.470 96.860 ;
        RECT 124.810 96.520 130.470 96.660 ;
        RECT 130.815 96.660 131.105 96.705 ;
        RECT 131.620 96.660 131.940 96.720 ;
        RECT 130.815 96.520 131.940 96.660 ;
        RECT 119.200 96.320 119.520 96.380 ;
        RECT 124.810 96.320 124.950 96.520 ;
        RECT 130.815 96.475 131.105 96.520 ;
        RECT 131.620 96.460 131.940 96.520 ;
        RECT 132.080 96.460 132.400 96.720 ;
        RECT 132.630 96.660 132.770 96.860 ;
        RECT 133.935 96.660 134.225 96.705 ;
        RECT 132.630 96.520 134.225 96.660 ;
        RECT 133.935 96.475 134.225 96.520 ;
        RECT 135.300 96.660 135.620 96.720 ;
        RECT 135.775 96.660 136.065 96.705 ;
        RECT 135.300 96.520 136.065 96.660 ;
        RECT 135.300 96.460 135.620 96.520 ;
        RECT 135.775 96.475 136.065 96.520 ;
        RECT 119.200 96.180 124.950 96.320 ;
        RECT 127.505 96.320 127.795 96.365 ;
        RECT 130.025 96.320 130.315 96.365 ;
        RECT 131.215 96.320 131.505 96.365 ;
        RECT 127.505 96.180 131.505 96.320 ;
        RECT 119.200 96.120 119.520 96.180 ;
        RECT 127.505 96.135 127.795 96.180 ;
        RECT 130.025 96.135 130.315 96.180 ;
        RECT 131.215 96.135 131.505 96.180 ;
        RECT 115.150 95.840 118.970 95.980 ;
        RECT 127.940 95.980 128.230 96.025 ;
        RECT 129.510 95.980 129.800 96.025 ;
        RECT 131.610 95.980 131.900 96.025 ;
        RECT 127.940 95.840 131.900 95.980 ;
        RECT 127.940 95.795 128.230 95.840 ;
        RECT 129.510 95.795 129.800 95.840 ;
        RECT 131.610 95.795 131.900 95.840 ;
        RECT 134.840 95.780 135.160 96.040 ;
        RECT 136.680 95.780 137.000 96.040 ;
        RECT 98.590 95.500 112.070 95.640 ;
        RECT 112.315 95.640 112.605 95.685 ;
        RECT 113.680 95.640 114.000 95.700 ;
        RECT 112.315 95.500 114.000 95.640 ;
        RECT 112.315 95.455 112.605 95.500 ;
        RECT 113.680 95.440 114.000 95.500 ;
        RECT 120.120 95.440 120.440 95.700 ;
        RECT 121.055 95.640 121.345 95.685 ;
        RECT 122.420 95.640 122.740 95.700 ;
        RECT 121.055 95.500 122.740 95.640 ;
        RECT 121.055 95.455 121.345 95.500 ;
        RECT 122.420 95.440 122.740 95.500 ;
        RECT 123.340 95.640 123.660 95.700 ;
        RECT 125.195 95.640 125.485 95.685 ;
        RECT 123.340 95.500 125.485 95.640 ;
        RECT 123.340 95.440 123.660 95.500 ;
        RECT 125.195 95.455 125.485 95.500 ;
        RECT 13.330 94.820 138.910 95.300 ;
        RECT 85.175 94.620 85.465 94.665 ;
        RECT 88.380 94.620 88.700 94.680 ;
        RECT 85.175 94.480 88.700 94.620 ;
        RECT 85.175 94.435 85.465 94.480 ;
        RECT 88.380 94.420 88.700 94.480 ;
        RECT 90.220 94.620 90.540 94.680 ;
        RECT 90.220 94.480 101.030 94.620 ;
        RECT 90.220 94.420 90.540 94.480 ;
        RECT 78.760 94.280 79.050 94.325 ;
        RECT 80.860 94.280 81.150 94.325 ;
        RECT 82.430 94.280 82.720 94.325 ;
        RECT 78.760 94.140 82.720 94.280 ;
        RECT 78.760 94.095 79.050 94.140 ;
        RECT 80.860 94.095 81.150 94.140 ;
        RECT 82.430 94.095 82.720 94.140 ;
        RECT 87.500 94.280 87.790 94.325 ;
        RECT 89.600 94.280 89.890 94.325 ;
        RECT 91.170 94.280 91.460 94.325 ;
        RECT 87.500 94.140 91.460 94.280 ;
        RECT 87.500 94.095 87.790 94.140 ;
        RECT 89.600 94.095 89.890 94.140 ;
        RECT 91.170 94.095 91.460 94.140 ;
        RECT 94.860 94.280 95.150 94.325 ;
        RECT 96.960 94.280 97.250 94.325 ;
        RECT 98.530 94.280 98.820 94.325 ;
        RECT 94.860 94.140 98.820 94.280 ;
        RECT 94.860 94.095 95.150 94.140 ;
        RECT 96.960 94.095 97.250 94.140 ;
        RECT 98.530 94.095 98.820 94.140 ;
        RECT 79.155 93.940 79.445 93.985 ;
        RECT 80.345 93.940 80.635 93.985 ;
        RECT 82.865 93.940 83.155 93.985 ;
        RECT 79.155 93.800 83.155 93.940 ;
        RECT 79.155 93.755 79.445 93.800 ;
        RECT 80.345 93.755 80.635 93.800 ;
        RECT 82.865 93.755 83.155 93.800 ;
        RECT 87.895 93.940 88.185 93.985 ;
        RECT 89.085 93.940 89.375 93.985 ;
        RECT 91.605 93.940 91.895 93.985 ;
        RECT 87.895 93.800 91.895 93.940 ;
        RECT 87.895 93.755 88.185 93.800 ;
        RECT 89.085 93.755 89.375 93.800 ;
        RECT 91.605 93.755 91.895 93.800 ;
        RECT 95.255 93.940 95.545 93.985 ;
        RECT 96.445 93.940 96.735 93.985 ;
        RECT 98.965 93.940 99.255 93.985 ;
        RECT 95.255 93.800 99.255 93.940 ;
        RECT 100.890 93.940 101.030 94.480 ;
        RECT 102.640 94.420 102.960 94.680 ;
        RECT 104.020 94.420 104.340 94.680 ;
        RECT 123.340 94.620 123.660 94.680 ;
        RECT 108.710 94.480 123.660 94.620 ;
        RECT 101.260 94.280 101.580 94.340 ;
        RECT 101.260 94.140 107.470 94.280 ;
        RECT 101.260 94.080 101.580 94.140 ;
        RECT 104.480 93.940 104.800 94.000 ;
        RECT 100.890 93.800 104.800 93.940 ;
        RECT 95.255 93.755 95.545 93.800 ;
        RECT 96.445 93.755 96.735 93.800 ;
        RECT 98.965 93.755 99.255 93.800 ;
        RECT 104.480 93.740 104.800 93.800 ;
        RECT 104.940 93.940 105.260 94.000 ;
        RECT 104.940 93.800 106.090 93.940 ;
        RECT 104.940 93.740 105.260 93.800 ;
        RECT 76.420 93.600 76.740 93.660 ;
        RECT 78.275 93.600 78.565 93.645 ;
        RECT 85.160 93.600 85.480 93.660 ;
        RECT 87.015 93.600 87.305 93.645 ;
        RECT 94.375 93.600 94.665 93.645 ;
        RECT 98.500 93.600 98.820 93.660 ;
        RECT 105.950 93.645 106.090 93.800 ;
        RECT 106.780 93.740 107.100 94.000 ;
        RECT 107.330 93.940 107.470 94.140 ;
        RECT 108.710 93.940 108.850 94.480 ;
        RECT 123.340 94.420 123.660 94.480 ;
        RECT 125.640 94.620 125.960 94.680 ;
        RECT 126.115 94.620 126.405 94.665 ;
        RECT 125.640 94.480 126.405 94.620 ;
        RECT 125.640 94.420 125.960 94.480 ;
        RECT 126.115 94.435 126.405 94.480 ;
        RECT 131.620 94.620 131.940 94.680 ;
        RECT 133.015 94.620 133.305 94.665 ;
        RECT 131.620 94.480 133.305 94.620 ;
        RECT 131.620 94.420 131.940 94.480 ;
        RECT 133.015 94.435 133.305 94.480 ;
        RECT 114.140 94.280 114.430 94.325 ;
        RECT 115.710 94.280 116.000 94.325 ;
        RECT 117.810 94.280 118.100 94.325 ;
        RECT 114.140 94.140 118.100 94.280 ;
        RECT 114.140 94.095 114.430 94.140 ;
        RECT 115.710 94.095 116.000 94.140 ;
        RECT 117.810 94.095 118.100 94.140 ;
        RECT 119.240 94.280 119.530 94.325 ;
        RECT 121.340 94.280 121.630 94.325 ;
        RECT 122.910 94.280 123.200 94.325 ;
        RECT 119.240 94.140 123.200 94.280 ;
        RECT 119.240 94.095 119.530 94.140 ;
        RECT 121.340 94.095 121.630 94.140 ;
        RECT 122.910 94.095 123.200 94.140 ;
        RECT 124.720 94.280 125.040 94.340 ;
        RECT 124.720 94.140 135.990 94.280 ;
        RECT 124.720 94.080 125.040 94.140 ;
        RECT 113.705 93.940 113.995 93.985 ;
        RECT 116.225 93.940 116.515 93.985 ;
        RECT 117.415 93.940 117.705 93.985 ;
        RECT 107.330 93.800 107.930 93.940 ;
        RECT 108.710 93.800 109.310 93.940 ;
        RECT 105.415 93.600 105.705 93.645 ;
        RECT 76.420 93.460 98.820 93.600 ;
        RECT 76.420 93.400 76.740 93.460 ;
        RECT 78.275 93.415 78.565 93.460 ;
        RECT 85.160 93.400 85.480 93.460 ;
        RECT 87.015 93.415 87.305 93.460 ;
        RECT 94.375 93.415 94.665 93.460 ;
        RECT 98.500 93.400 98.820 93.460 ;
        RECT 104.570 93.460 105.705 93.600 ;
        RECT 104.570 93.320 104.710 93.460 ;
        RECT 105.415 93.415 105.705 93.460 ;
        RECT 105.875 93.415 106.165 93.645 ;
        RECT 106.320 93.400 106.640 93.660 ;
        RECT 106.870 93.585 107.010 93.740 ;
        RECT 107.790 93.645 107.930 93.800 ;
        RECT 107.255 93.585 107.545 93.645 ;
        RECT 106.870 93.445 107.545 93.585 ;
        RECT 107.255 93.415 107.545 93.445 ;
        RECT 107.715 93.415 108.005 93.645 ;
        RECT 108.620 93.400 108.940 93.660 ;
        RECT 109.170 93.645 109.310 93.800 ;
        RECT 113.705 93.800 117.705 93.940 ;
        RECT 113.705 93.755 113.995 93.800 ;
        RECT 116.225 93.755 116.515 93.800 ;
        RECT 117.415 93.755 117.705 93.800 ;
        RECT 118.295 93.940 118.585 93.985 ;
        RECT 118.740 93.940 119.060 94.000 ;
        RECT 118.295 93.800 119.060 93.940 ;
        RECT 118.295 93.755 118.585 93.800 ;
        RECT 118.740 93.740 119.060 93.800 ;
        RECT 119.635 93.940 119.925 93.985 ;
        RECT 120.825 93.940 121.115 93.985 ;
        RECT 123.345 93.940 123.635 93.985 ;
        RECT 119.635 93.800 123.635 93.940 ;
        RECT 119.635 93.755 119.925 93.800 ;
        RECT 120.825 93.755 121.115 93.800 ;
        RECT 123.345 93.755 123.635 93.800 ;
        RECT 125.180 93.940 125.500 94.000 ;
        RECT 125.180 93.800 131.850 93.940 ;
        RECT 125.180 93.740 125.500 93.800 ;
        RECT 109.095 93.415 109.385 93.645 ;
        RECT 109.675 93.600 109.965 93.645 ;
        RECT 109.630 93.415 109.965 93.600 ;
        RECT 110.460 93.600 110.780 93.660 ;
        RECT 115.520 93.600 115.840 93.660 ;
        RECT 120.120 93.645 120.440 93.660 ;
        RECT 120.090 93.600 120.440 93.645 ;
        RECT 127.955 93.600 128.245 93.645 ;
        RECT 128.400 93.600 128.720 93.660 ;
        RECT 110.460 93.460 114.370 93.600 ;
        RECT 79.640 93.305 79.960 93.320 ;
        RECT 79.610 93.260 79.960 93.305 ;
        RECT 79.445 93.120 79.960 93.260 ;
        RECT 79.610 93.075 79.960 93.120 ;
        RECT 88.350 93.260 88.640 93.305 ;
        RECT 91.140 93.260 91.460 93.320 ;
        RECT 88.350 93.120 91.460 93.260 ;
        RECT 88.350 93.075 88.640 93.120 ;
        RECT 79.640 93.060 79.960 93.075 ;
        RECT 91.140 93.060 91.460 93.120 ;
        RECT 95.710 93.260 96.000 93.305 ;
        RECT 96.660 93.260 96.980 93.320 ;
        RECT 95.710 93.120 96.980 93.260 ;
        RECT 95.710 93.075 96.000 93.120 ;
        RECT 96.660 93.060 96.980 93.120 ;
        RECT 101.720 93.260 102.040 93.320 ;
        RECT 102.195 93.260 102.485 93.305 ;
        RECT 101.720 93.120 102.485 93.260 ;
        RECT 101.720 93.060 102.040 93.120 ;
        RECT 102.195 93.075 102.485 93.120 ;
        RECT 104.480 93.060 104.800 93.320 ;
        RECT 109.630 93.260 109.770 93.415 ;
        RECT 110.460 93.400 110.780 93.460 ;
        RECT 109.170 93.120 109.770 93.260 ;
        RECT 109.170 92.980 109.310 93.120 ;
        RECT 92.520 92.920 92.840 92.980 ;
        RECT 93.915 92.920 94.205 92.965 ;
        RECT 96.200 92.920 96.520 92.980 ;
        RECT 104.940 92.920 105.260 92.980 ;
        RECT 92.520 92.780 105.260 92.920 ;
        RECT 92.520 92.720 92.840 92.780 ;
        RECT 93.915 92.735 94.205 92.780 ;
        RECT 96.200 92.720 96.520 92.780 ;
        RECT 104.940 92.720 105.260 92.780 ;
        RECT 109.080 92.720 109.400 92.980 ;
        RECT 109.540 92.920 109.860 92.980 ;
        RECT 110.475 92.920 110.765 92.965 ;
        RECT 109.540 92.780 110.765 92.920 ;
        RECT 109.540 92.720 109.860 92.780 ;
        RECT 110.475 92.735 110.765 92.780 ;
        RECT 111.395 92.920 111.685 92.965 ;
        RECT 113.680 92.920 114.000 92.980 ;
        RECT 111.395 92.780 114.000 92.920 ;
        RECT 114.230 92.920 114.370 93.460 ;
        RECT 115.520 93.460 118.280 93.600 ;
        RECT 119.925 93.460 120.440 93.600 ;
        RECT 115.520 93.400 115.840 93.460 ;
        RECT 116.900 93.305 117.220 93.320 ;
        RECT 116.900 93.075 117.250 93.305 ;
        RECT 118.140 93.260 118.280 93.460 ;
        RECT 120.090 93.415 120.440 93.460 ;
        RECT 120.120 93.400 120.440 93.415 ;
        RECT 124.810 93.460 128.720 93.600 ;
        RECT 124.810 93.260 124.950 93.460 ;
        RECT 127.955 93.415 128.245 93.460 ;
        RECT 128.400 93.400 128.720 93.460 ;
        RECT 129.795 93.415 130.085 93.645 ;
        RECT 130.240 93.600 130.560 93.660 ;
        RECT 130.715 93.600 131.005 93.645 ;
        RECT 130.240 93.460 131.005 93.600 ;
        RECT 118.140 93.120 124.950 93.260 ;
        RECT 125.180 93.260 125.500 93.320 ;
        RECT 125.180 93.120 126.790 93.260 ;
        RECT 116.900 93.060 117.220 93.075 ;
        RECT 125.180 93.060 125.500 93.120 ;
        RECT 121.960 92.920 122.280 92.980 ;
        RECT 114.230 92.780 122.280 92.920 ;
        RECT 111.395 92.735 111.685 92.780 ;
        RECT 113.680 92.720 114.000 92.780 ;
        RECT 121.960 92.720 122.280 92.780 ;
        RECT 122.880 92.920 123.200 92.980 ;
        RECT 125.655 92.920 125.945 92.965 ;
        RECT 122.880 92.780 125.945 92.920 ;
        RECT 126.650 92.920 126.790 93.120 ;
        RECT 127.020 93.060 127.340 93.320 ;
        RECT 129.870 92.920 130.010 93.415 ;
        RECT 130.240 93.400 130.560 93.460 ;
        RECT 130.715 93.415 131.005 93.460 ;
        RECT 131.160 93.400 131.480 93.660 ;
        RECT 131.710 93.645 131.850 93.800 ;
        RECT 135.850 93.645 135.990 94.140 ;
        RECT 131.635 93.415 131.925 93.645 ;
        RECT 135.775 93.415 136.065 93.645 ;
        RECT 126.650 92.780 130.010 92.920 ;
        RECT 122.880 92.720 123.200 92.780 ;
        RECT 125.655 92.735 125.945 92.780 ;
        RECT 136.680 92.720 137.000 92.980 ;
        RECT 13.330 92.100 138.910 92.580 ;
        RECT 83.795 91.900 84.085 91.945 ;
        RECT 85.620 91.900 85.940 91.960 ;
        RECT 83.795 91.760 85.940 91.900 ;
        RECT 83.795 91.715 84.085 91.760 ;
        RECT 85.620 91.700 85.940 91.760 ;
        RECT 91.140 91.700 91.460 91.960 ;
        RECT 91.600 91.900 91.920 91.960 ;
        RECT 94.360 91.900 94.680 91.960 ;
        RECT 95.295 91.900 95.585 91.945 ;
        RECT 105.860 91.900 106.180 91.960 ;
        RECT 91.600 91.760 93.670 91.900 ;
        RECT 91.600 91.700 91.920 91.760 ;
        RECT 77.770 91.560 78.060 91.605 ;
        RECT 83.320 91.560 83.640 91.620 ;
        RECT 77.770 91.420 83.640 91.560 ;
        RECT 77.770 91.375 78.060 91.420 ;
        RECT 83.320 91.360 83.640 91.420 ;
        RECT 84.240 91.560 84.560 91.620 ;
        RECT 86.095 91.560 86.385 91.605 ;
        RECT 84.240 91.420 86.385 91.560 ;
        RECT 84.240 91.360 84.560 91.420 ;
        RECT 86.095 91.375 86.385 91.420 ;
        RECT 87.015 91.560 87.305 91.605 ;
        RECT 88.380 91.560 88.700 91.620 ;
        RECT 87.015 91.420 88.700 91.560 ;
        RECT 87.015 91.375 87.305 91.420 ;
        RECT 88.380 91.360 88.700 91.420 ;
        RECT 90.680 91.560 91.000 91.620 ;
        RECT 90.680 91.420 93.210 91.560 ;
        RECT 90.680 91.360 91.000 91.420 ;
        RECT 76.420 91.020 76.740 91.280 ;
        RECT 84.770 91.220 85.060 91.265 ;
        RECT 85.635 91.220 85.925 91.265 ;
        RECT 87.935 91.220 88.225 91.265 ;
        RECT 84.770 91.080 85.345 91.220 ;
        RECT 84.770 91.035 85.060 91.080 ;
        RECT 77.315 90.880 77.605 90.925 ;
        RECT 78.505 90.880 78.795 90.925 ;
        RECT 81.025 90.880 81.315 90.925 ;
        RECT 77.315 90.740 81.315 90.880 ;
        RECT 77.315 90.695 77.605 90.740 ;
        RECT 78.505 90.695 78.795 90.740 ;
        RECT 81.025 90.695 81.315 90.740 ;
        RECT 85.205 90.880 85.345 91.080 ;
        RECT 85.635 91.080 88.225 91.220 ;
        RECT 85.635 91.035 85.925 91.080 ;
        RECT 87.935 91.035 88.225 91.080 ;
        RECT 87.460 90.880 87.780 90.940 ;
        RECT 85.205 90.740 87.780 90.880 ;
        RECT 88.010 90.880 88.150 91.035 ;
        RECT 92.520 91.020 92.840 91.280 ;
        RECT 93.070 91.265 93.210 91.420 ;
        RECT 93.530 91.265 93.670 91.760 ;
        RECT 94.360 91.760 95.585 91.900 ;
        RECT 94.360 91.700 94.680 91.760 ;
        RECT 95.295 91.715 95.585 91.760 ;
        RECT 104.110 91.760 106.180 91.900 ;
        RECT 96.215 91.560 96.505 91.605 ;
        RECT 99.420 91.560 99.740 91.620 ;
        RECT 101.260 91.560 101.580 91.620 ;
        RECT 96.215 91.420 101.580 91.560 ;
        RECT 96.215 91.375 96.505 91.420 ;
        RECT 99.420 91.360 99.740 91.420 ;
        RECT 101.260 91.360 101.580 91.420 ;
        RECT 103.270 91.560 103.560 91.605 ;
        RECT 104.110 91.560 104.250 91.760 ;
        RECT 105.860 91.700 106.180 91.760 ;
        RECT 106.780 91.700 107.100 91.960 ;
        RECT 107.240 91.900 107.560 91.960 ;
        RECT 109.095 91.900 109.385 91.945 ;
        RECT 107.240 91.760 109.385 91.900 ;
        RECT 107.240 91.700 107.560 91.760 ;
        RECT 109.095 91.715 109.385 91.760 ;
        RECT 109.540 91.900 109.860 91.960 ;
        RECT 113.220 91.900 113.540 91.960 ;
        RECT 115.075 91.900 115.365 91.945 ;
        RECT 109.540 91.760 112.070 91.900 ;
        RECT 109.540 91.700 109.860 91.760 ;
        RECT 103.270 91.420 104.250 91.560 ;
        RECT 109.170 91.420 110.230 91.560 ;
        RECT 103.270 91.375 103.560 91.420 ;
        RECT 109.170 91.280 109.310 91.420 ;
        RECT 92.995 91.035 93.285 91.265 ;
        RECT 93.455 91.035 93.745 91.265 ;
        RECT 94.360 91.020 94.680 91.280 ;
        RECT 94.820 91.220 95.140 91.280 ;
        RECT 97.120 91.220 97.440 91.280 ;
        RECT 101.720 91.220 102.040 91.280 ;
        RECT 94.820 91.080 97.440 91.220 ;
        RECT 94.820 91.020 95.140 91.080 ;
        RECT 97.120 91.020 97.440 91.080 ;
        RECT 99.510 91.080 102.040 91.220 ;
        RECT 94.910 90.880 95.050 91.020 ;
        RECT 88.010 90.740 95.050 90.880 ;
        RECT 76.920 90.540 77.210 90.585 ;
        RECT 79.020 90.540 79.310 90.585 ;
        RECT 80.590 90.540 80.880 90.585 ;
        RECT 76.920 90.400 80.880 90.540 ;
        RECT 76.920 90.355 77.210 90.400 ;
        RECT 79.020 90.355 79.310 90.400 ;
        RECT 80.590 90.355 80.880 90.400 ;
        RECT 83.335 90.540 83.625 90.585 ;
        RECT 83.780 90.540 84.100 90.600 ;
        RECT 85.205 90.540 85.345 90.740 ;
        RECT 87.460 90.680 87.780 90.740 ;
        RECT 83.335 90.400 85.345 90.540 ;
        RECT 92.980 90.540 93.300 90.600 ;
        RECT 94.360 90.540 94.680 90.600 ;
        RECT 99.510 90.540 99.650 91.080 ;
        RECT 101.720 91.020 102.040 91.080 ;
        RECT 104.955 91.220 105.245 91.265 ;
        RECT 105.400 91.220 105.720 91.280 ;
        RECT 104.955 91.080 105.720 91.220 ;
        RECT 104.955 91.035 105.245 91.080 ;
        RECT 105.400 91.020 105.720 91.080 ;
        RECT 105.875 91.220 106.165 91.265 ;
        RECT 106.320 91.220 106.640 91.280 ;
        RECT 105.875 91.080 106.640 91.220 ;
        RECT 105.875 91.035 106.165 91.080 ;
        RECT 106.320 91.020 106.640 91.080 ;
        RECT 109.080 91.020 109.400 91.280 ;
        RECT 110.090 91.265 110.230 91.420 ;
        RECT 110.920 91.360 111.240 91.620 ;
        RECT 111.930 91.265 112.070 91.760 ;
        RECT 113.220 91.760 115.365 91.900 ;
        RECT 113.220 91.700 113.540 91.760 ;
        RECT 115.075 91.715 115.365 91.760 ;
        RECT 116.900 91.700 117.220 91.960 ;
        RECT 118.740 91.900 119.060 91.960 ;
        RECT 118.140 91.760 119.060 91.900 ;
        RECT 112.760 91.560 113.080 91.620 ;
        RECT 118.140 91.560 118.280 91.760 ;
        RECT 118.740 91.700 119.060 91.760 ;
        RECT 120.120 91.900 120.440 91.960 ;
        RECT 124.260 91.900 124.580 91.960 ;
        RECT 120.120 91.760 124.580 91.900 ;
        RECT 120.120 91.700 120.440 91.760 ;
        RECT 124.260 91.700 124.580 91.760 ;
        RECT 127.020 91.900 127.340 91.960 ;
        RECT 127.955 91.900 128.245 91.945 ;
        RECT 127.020 91.760 128.245 91.900 ;
        RECT 127.020 91.700 127.340 91.760 ;
        RECT 127.955 91.715 128.245 91.760 ;
        RECT 130.240 91.700 130.560 91.960 ;
        RECT 122.420 91.605 122.740 91.620 ;
        RECT 122.390 91.560 122.740 91.605 ;
        RECT 112.760 91.420 121.270 91.560 ;
        RECT 122.225 91.420 122.740 91.560 ;
        RECT 112.760 91.360 113.080 91.420 ;
        RECT 109.895 91.080 110.230 91.265 ;
        RECT 109.895 91.035 110.185 91.080 ;
        RECT 110.475 91.035 110.765 91.265 ;
        RECT 111.855 91.035 112.145 91.265 ;
        RECT 99.905 90.880 100.195 90.925 ;
        RECT 102.425 90.880 102.715 90.925 ;
        RECT 103.615 90.880 103.905 90.925 ;
        RECT 99.905 90.740 103.905 90.880 ;
        RECT 99.905 90.695 100.195 90.740 ;
        RECT 102.425 90.695 102.715 90.740 ;
        RECT 103.615 90.695 103.905 90.740 ;
        RECT 104.495 90.695 104.785 90.925 ;
        RECT 108.620 90.880 108.940 90.940 ;
        RECT 110.550 90.880 110.690 91.035 ;
        RECT 112.300 91.020 112.620 91.280 ;
        RECT 113.220 91.020 113.540 91.280 ;
        RECT 113.680 91.020 114.000 91.280 ;
        RECT 114.155 91.220 114.445 91.265 ;
        RECT 114.600 91.220 114.920 91.280 ;
        RECT 114.155 91.080 114.920 91.220 ;
        RECT 114.155 91.035 114.445 91.080 ;
        RECT 114.600 91.020 114.920 91.080 ;
        RECT 118.280 91.020 118.600 91.280 ;
        RECT 118.755 91.035 119.045 91.265 ;
        RECT 108.620 90.740 110.690 90.880 ;
        RECT 118.830 90.880 118.970 91.035 ;
        RECT 119.200 91.020 119.520 91.280 ;
        RECT 120.120 91.020 120.440 91.280 ;
        RECT 121.130 91.265 121.270 91.420 ;
        RECT 122.390 91.375 122.740 91.420 ;
        RECT 122.420 91.360 122.740 91.375 ;
        RECT 123.340 91.360 123.660 91.620 ;
        RECT 128.400 91.360 128.720 91.620 ;
        RECT 121.055 91.035 121.345 91.265 ;
        RECT 123.430 91.220 123.570 91.360 ;
        RECT 129.335 91.220 129.625 91.265 ;
        RECT 132.080 91.220 132.400 91.280 ;
        RECT 123.430 91.080 132.400 91.220 ;
        RECT 129.335 91.035 129.625 91.080 ;
        RECT 132.080 91.020 132.400 91.080 ;
        RECT 133.920 91.220 134.240 91.280 ;
        RECT 135.775 91.220 136.065 91.265 ;
        RECT 133.920 91.080 136.065 91.220 ;
        RECT 133.920 91.020 134.240 91.080 ;
        RECT 135.775 91.035 136.065 91.080 ;
        RECT 120.580 90.880 120.900 90.940 ;
        RECT 118.830 90.740 120.900 90.880 ;
        RECT 92.980 90.400 99.650 90.540 ;
        RECT 100.340 90.540 100.630 90.585 ;
        RECT 101.910 90.540 102.200 90.585 ;
        RECT 104.010 90.540 104.300 90.585 ;
        RECT 100.340 90.400 104.300 90.540 ;
        RECT 104.570 90.540 104.710 90.695 ;
        RECT 108.620 90.680 108.940 90.740 ;
        RECT 120.580 90.680 120.900 90.740 ;
        RECT 121.935 90.880 122.225 90.925 ;
        RECT 123.125 90.880 123.415 90.925 ;
        RECT 125.645 90.880 125.935 90.925 ;
        RECT 121.935 90.740 125.935 90.880 ;
        RECT 121.935 90.695 122.225 90.740 ;
        RECT 123.125 90.695 123.415 90.740 ;
        RECT 125.645 90.695 125.935 90.740 ;
        RECT 121.540 90.540 121.830 90.585 ;
        RECT 123.640 90.540 123.930 90.585 ;
        RECT 125.210 90.540 125.500 90.585 ;
        RECT 104.570 90.400 111.610 90.540 ;
        RECT 83.335 90.355 83.625 90.400 ;
        RECT 83.780 90.340 84.100 90.400 ;
        RECT 92.980 90.340 93.300 90.400 ;
        RECT 94.360 90.340 94.680 90.400 ;
        RECT 100.340 90.355 100.630 90.400 ;
        RECT 101.910 90.355 102.200 90.400 ;
        RECT 104.010 90.355 104.300 90.400 ;
        RECT 97.595 90.200 97.885 90.245 ;
        RECT 100.800 90.200 101.120 90.260 ;
        RECT 97.595 90.060 101.120 90.200 ;
        RECT 97.595 90.015 97.885 90.060 ;
        RECT 100.800 90.000 101.120 90.060 ;
        RECT 104.480 90.200 104.800 90.260 ;
        RECT 107.240 90.200 107.560 90.260 ;
        RECT 110.460 90.200 110.780 90.260 ;
        RECT 104.480 90.060 110.780 90.200 ;
        RECT 111.470 90.200 111.610 90.400 ;
        RECT 121.540 90.400 125.500 90.540 ;
        RECT 121.540 90.355 121.830 90.400 ;
        RECT 123.640 90.355 123.930 90.400 ;
        RECT 125.210 90.355 125.500 90.400 ;
        RECT 112.760 90.200 113.080 90.260 ;
        RECT 111.470 90.060 113.080 90.200 ;
        RECT 104.480 90.000 104.800 90.060 ;
        RECT 107.240 90.000 107.560 90.060 ;
        RECT 110.460 90.000 110.780 90.060 ;
        RECT 112.760 90.000 113.080 90.060 ;
        RECT 113.220 90.200 113.540 90.260 ;
        RECT 115.520 90.200 115.840 90.260 ;
        RECT 113.220 90.060 115.840 90.200 ;
        RECT 113.220 90.000 113.540 90.060 ;
        RECT 115.520 90.000 115.840 90.060 ;
        RECT 136.680 90.000 137.000 90.260 ;
        RECT 13.330 89.380 138.910 89.860 ;
        RECT 59.860 89.180 60.180 89.240 ;
        RECT 60.795 89.180 61.085 89.225 ;
        RECT 59.860 89.040 61.085 89.180 ;
        RECT 59.860 88.980 60.180 89.040 ;
        RECT 60.795 88.995 61.085 89.040 ;
        RECT 100.800 89.180 101.120 89.240 ;
        RECT 114.140 89.180 114.460 89.240 ;
        RECT 117.835 89.180 118.125 89.225 ;
        RECT 100.800 89.040 105.630 89.180 ;
        RECT 100.800 88.980 101.120 89.040 ;
        RECT 101.260 88.840 101.580 88.900 ;
        RECT 104.495 88.840 104.785 88.885 ;
        RECT 101.260 88.700 104.785 88.840 ;
        RECT 101.260 88.640 101.580 88.700 ;
        RECT 104.495 88.655 104.785 88.700 ;
        RECT 70.900 88.300 71.220 88.560 ;
        RECT 97.580 88.500 97.900 88.560 ;
        RECT 104.940 88.500 105.260 88.560 ;
        RECT 97.580 88.360 105.260 88.500 ;
        RECT 97.580 88.300 97.900 88.360 ;
        RECT 59.400 88.160 59.720 88.220 ;
        RECT 59.875 88.160 60.165 88.205 ;
        RECT 59.400 88.020 60.165 88.160 ;
        RECT 59.400 87.960 59.720 88.020 ;
        RECT 59.875 87.975 60.165 88.020 ;
        RECT 67.680 87.960 68.000 88.220 ;
        RECT 69.060 88.160 69.380 88.220 ;
        RECT 69.535 88.160 69.825 88.205 ;
        RECT 69.060 88.020 69.825 88.160 ;
        RECT 69.060 87.960 69.380 88.020 ;
        RECT 69.535 87.975 69.825 88.020 ;
        RECT 75.515 88.160 75.805 88.205 ;
        RECT 76.880 88.160 77.200 88.220 ;
        RECT 75.515 88.020 77.200 88.160 ;
        RECT 75.515 87.975 75.805 88.020 ;
        RECT 76.880 87.960 77.200 88.020 ;
        RECT 77.340 87.960 77.660 88.220 ;
        RECT 77.800 88.160 78.120 88.220 ;
        RECT 80.575 88.160 80.865 88.205 ;
        RECT 77.800 88.020 80.865 88.160 ;
        RECT 77.800 87.960 78.120 88.020 ;
        RECT 80.575 87.975 80.865 88.020 ;
        RECT 83.780 87.960 84.100 88.220 ;
        RECT 87.015 88.160 87.305 88.205 ;
        RECT 88.380 88.160 88.700 88.220 ;
        RECT 87.015 88.020 88.700 88.160 ;
        RECT 87.015 87.975 87.305 88.020 ;
        RECT 88.380 87.960 88.700 88.020 ;
        RECT 90.235 88.160 90.525 88.205 ;
        RECT 92.060 88.160 92.380 88.220 ;
        RECT 90.235 88.020 92.380 88.160 ;
        RECT 90.235 87.975 90.525 88.020 ;
        RECT 92.060 87.960 92.380 88.020 ;
        RECT 93.455 88.160 93.745 88.205 ;
        RECT 93.900 88.160 94.220 88.220 ;
        RECT 93.455 88.020 94.220 88.160 ;
        RECT 93.455 87.975 93.745 88.020 ;
        RECT 93.900 87.960 94.220 88.020 ;
        RECT 96.660 87.960 96.980 88.220 ;
        RECT 99.420 87.960 99.740 88.220 ;
        RECT 99.970 88.205 100.110 88.360 ;
        RECT 104.940 88.300 105.260 88.360 ;
        RECT 105.490 88.500 105.630 89.040 ;
        RECT 114.140 89.040 118.125 89.180 ;
        RECT 114.140 88.980 114.460 89.040 ;
        RECT 117.835 88.995 118.125 89.040 ;
        RECT 109.540 88.640 109.860 88.900 ;
        RECT 115.535 88.840 115.825 88.885 ;
        RECT 119.200 88.840 119.520 88.900 ;
        RECT 115.535 88.700 119.520 88.840 ;
        RECT 115.535 88.655 115.825 88.700 ;
        RECT 119.200 88.640 119.520 88.700 ;
        RECT 119.675 88.655 119.965 88.885 ;
        RECT 109.630 88.500 109.770 88.640 ;
        RECT 105.490 88.360 109.770 88.500 ;
        RECT 112.300 88.500 112.620 88.560 ;
        RECT 119.750 88.500 119.890 88.655 ;
        RECT 112.300 88.360 117.130 88.500 ;
        RECT 99.895 88.160 100.185 88.205 ;
        RECT 99.895 88.020 100.295 88.160 ;
        RECT 99.895 87.975 100.185 88.020 ;
        RECT 100.800 87.960 101.120 88.220 ;
        RECT 105.490 88.205 105.630 88.360 ;
        RECT 112.300 88.300 112.620 88.360 ;
        RECT 105.415 87.975 105.705 88.205 ;
        RECT 106.320 88.160 106.640 88.220 ;
        RECT 107.255 88.160 107.545 88.205 ;
        RECT 106.320 88.020 107.545 88.160 ;
        RECT 106.320 87.960 106.640 88.020 ;
        RECT 107.255 87.975 107.545 88.020 ;
        RECT 109.555 88.160 109.845 88.205 ;
        RECT 110.000 88.160 110.320 88.220 ;
        RECT 109.555 88.020 110.320 88.160 ;
        RECT 109.555 87.975 109.845 88.020 ;
        RECT 110.000 87.960 110.320 88.020 ;
        RECT 111.380 87.960 111.700 88.220 ;
        RECT 113.220 88.160 113.540 88.220 ;
        RECT 116.990 88.205 117.130 88.360 ;
        RECT 118.140 88.360 119.890 88.500 ;
        RECT 113.695 88.160 113.985 88.205 ;
        RECT 113.220 88.020 113.985 88.160 ;
        RECT 113.220 87.960 113.540 88.020 ;
        RECT 113.695 87.975 113.985 88.020 ;
        RECT 116.915 87.975 117.205 88.205 ;
        RECT 117.360 88.160 117.680 88.220 ;
        RECT 118.140 88.160 118.280 88.360 ;
        RECT 117.360 88.020 118.280 88.160 ;
        RECT 117.360 87.960 117.680 88.020 ;
        RECT 118.755 87.975 119.045 88.205 ;
        RECT 122.435 88.160 122.725 88.205 ;
        RECT 122.880 88.160 123.200 88.220 ;
        RECT 122.435 88.020 123.200 88.160 ;
        RECT 122.435 87.975 122.725 88.020 ;
        RECT 101.735 87.820 102.025 87.865 ;
        RECT 108.160 87.820 108.480 87.880 ;
        RECT 114.615 87.820 114.905 87.865 ;
        RECT 118.830 87.820 118.970 87.975 ;
        RECT 122.880 87.960 123.200 88.020 ;
        RECT 123.800 88.160 124.120 88.220 ;
        RECT 124.275 88.160 124.565 88.205 ;
        RECT 123.800 88.020 124.565 88.160 ;
        RECT 123.800 87.960 124.120 88.020 ;
        RECT 124.275 87.975 124.565 88.020 ;
        RECT 127.020 88.160 127.340 88.220 ;
        RECT 127.495 88.160 127.785 88.205 ;
        RECT 127.020 88.020 127.785 88.160 ;
        RECT 127.020 87.960 127.340 88.020 ;
        RECT 127.495 87.975 127.785 88.020 ;
        RECT 132.080 87.960 132.400 88.220 ;
        RECT 101.735 87.680 108.480 87.820 ;
        RECT 101.735 87.635 102.025 87.680 ;
        RECT 108.160 87.620 108.480 87.680 ;
        RECT 113.770 87.680 118.970 87.820 ;
        RECT 113.770 87.540 113.910 87.680 ;
        RECT 114.615 87.635 114.905 87.680 ;
        RECT 65.840 87.480 66.160 87.540 ;
        RECT 66.775 87.480 67.065 87.525 ;
        RECT 65.840 87.340 67.065 87.480 ;
        RECT 65.840 87.280 66.160 87.340 ;
        RECT 66.775 87.295 67.065 87.340 ;
        RECT 72.280 87.480 72.600 87.540 ;
        RECT 74.595 87.480 74.885 87.525 ;
        RECT 72.280 87.340 74.885 87.480 ;
        RECT 72.280 87.280 72.600 87.340 ;
        RECT 74.595 87.295 74.885 87.340 ;
        RECT 75.500 87.480 75.820 87.540 ;
        RECT 76.435 87.480 76.725 87.525 ;
        RECT 75.500 87.340 76.725 87.480 ;
        RECT 75.500 87.280 75.820 87.340 ;
        RECT 76.435 87.295 76.725 87.340 ;
        RECT 78.720 87.480 79.040 87.540 ;
        RECT 79.655 87.480 79.945 87.525 ;
        RECT 78.720 87.340 79.945 87.480 ;
        RECT 78.720 87.280 79.040 87.340 ;
        RECT 79.655 87.295 79.945 87.340 ;
        RECT 81.940 87.480 82.260 87.540 ;
        RECT 82.875 87.480 83.165 87.525 ;
        RECT 81.940 87.340 83.165 87.480 ;
        RECT 81.940 87.280 82.260 87.340 ;
        RECT 82.875 87.295 83.165 87.340 ;
        RECT 85.160 87.480 85.480 87.540 ;
        RECT 86.095 87.480 86.385 87.525 ;
        RECT 85.160 87.340 86.385 87.480 ;
        RECT 85.160 87.280 85.480 87.340 ;
        RECT 86.095 87.295 86.385 87.340 ;
        RECT 88.380 87.480 88.700 87.540 ;
        RECT 89.315 87.480 89.605 87.525 ;
        RECT 88.380 87.340 89.605 87.480 ;
        RECT 88.380 87.280 88.700 87.340 ;
        RECT 89.315 87.295 89.605 87.340 ;
        RECT 91.600 87.480 91.920 87.540 ;
        RECT 92.535 87.480 92.825 87.525 ;
        RECT 91.600 87.340 92.825 87.480 ;
        RECT 91.600 87.280 91.920 87.340 ;
        RECT 92.535 87.295 92.825 87.340 ;
        RECT 94.820 87.480 95.140 87.540 ;
        RECT 95.755 87.480 96.045 87.525 ;
        RECT 94.820 87.340 96.045 87.480 ;
        RECT 94.820 87.280 95.140 87.340 ;
        RECT 95.755 87.295 96.045 87.340 ;
        RECT 98.040 87.480 98.360 87.540 ;
        RECT 98.515 87.480 98.805 87.525 ;
        RECT 98.040 87.340 98.805 87.480 ;
        RECT 98.040 87.280 98.360 87.340 ;
        RECT 98.515 87.295 98.805 87.340 ;
        RECT 104.940 87.480 105.260 87.540 ;
        RECT 106.335 87.480 106.625 87.525 ;
        RECT 104.940 87.340 106.625 87.480 ;
        RECT 104.940 87.280 105.260 87.340 ;
        RECT 106.335 87.295 106.625 87.340 ;
        RECT 107.700 87.480 108.020 87.540 ;
        RECT 108.635 87.480 108.925 87.525 ;
        RECT 107.700 87.340 108.925 87.480 ;
        RECT 107.700 87.280 108.020 87.340 ;
        RECT 108.635 87.295 108.925 87.340 ;
        RECT 110.920 87.480 111.240 87.540 ;
        RECT 112.315 87.480 112.605 87.525 ;
        RECT 110.920 87.340 112.605 87.480 ;
        RECT 110.920 87.280 111.240 87.340 ;
        RECT 112.315 87.295 112.605 87.340 ;
        RECT 113.680 87.280 114.000 87.540 ;
        RECT 120.580 87.480 120.900 87.540 ;
        RECT 121.515 87.480 121.805 87.525 ;
        RECT 120.580 87.340 121.805 87.480 ;
        RECT 120.580 87.280 120.900 87.340 ;
        RECT 121.515 87.295 121.805 87.340 ;
        RECT 123.800 87.480 124.120 87.540 ;
        RECT 125.195 87.480 125.485 87.525 ;
        RECT 123.800 87.340 125.485 87.480 ;
        RECT 123.800 87.280 124.120 87.340 ;
        RECT 125.195 87.295 125.485 87.340 ;
        RECT 127.020 87.480 127.340 87.540 ;
        RECT 128.415 87.480 128.705 87.525 ;
        RECT 127.020 87.340 128.705 87.480 ;
        RECT 127.020 87.280 127.340 87.340 ;
        RECT 128.415 87.295 128.705 87.340 ;
        RECT 130.240 87.480 130.560 87.540 ;
        RECT 131.175 87.480 131.465 87.525 ;
        RECT 130.240 87.340 131.465 87.480 ;
        RECT 130.240 87.280 130.560 87.340 ;
        RECT 131.175 87.295 131.465 87.340 ;
        RECT 13.330 86.660 138.910 87.140 ;
        RECT 12.920 51.400 48.800 51.880 ;
        RECT 21.745 51.200 22.035 51.245 ;
        RECT 26.790 51.200 27.110 51.260 ;
        RECT 21.745 51.060 27.110 51.200 ;
        RECT 21.745 51.015 22.035 51.060 ;
        RECT 26.790 51.000 27.110 51.060 ;
        RECT 32.325 51.200 32.615 51.245 ;
        RECT 33.230 51.200 33.550 51.260 ;
        RECT 32.325 51.060 33.550 51.200 ;
        RECT 32.325 51.015 32.615 51.060 ;
        RECT 33.230 51.000 33.550 51.060 ;
        RECT 39.670 51.200 39.990 51.260 ;
        RECT 40.605 51.200 40.895 51.245 ;
        RECT 39.670 51.060 40.895 51.200 ;
        RECT 39.670 51.000 39.990 51.060 ;
        RECT 40.605 51.015 40.895 51.060 ;
        RECT 24.045 50.860 24.335 50.905 ;
        RECT 31.390 50.860 31.710 50.920 ;
        RECT 38.290 50.860 38.610 50.920 ;
        RECT 24.045 50.720 31.710 50.860 ;
        RECT 24.045 50.675 24.335 50.720 ;
        RECT 31.390 50.660 31.710 50.720 ;
        RECT 32.860 50.720 38.610 50.860 ;
        RECT 27.265 50.520 27.555 50.565 ;
        RECT 20.900 50.380 27.555 50.520 ;
        RECT 18.510 50.180 18.830 50.240 ;
        RECT 20.900 50.225 21.040 50.380 ;
        RECT 27.265 50.335 27.555 50.380 ;
        RECT 20.825 50.180 21.115 50.225 ;
        RECT 18.510 50.040 21.115 50.180 ;
        RECT 18.510 49.980 18.830 50.040 ;
        RECT 20.825 49.995 21.115 50.040 ;
        RECT 23.110 49.980 23.430 50.240 ;
        RECT 23.570 49.980 23.890 50.240 ;
        RECT 24.505 50.180 24.795 50.225 ;
        RECT 32.860 50.180 33.000 50.720 ;
        RECT 38.290 50.660 38.610 50.720 ;
        RECT 24.505 50.040 33.000 50.180 ;
        RECT 33.245 50.180 33.535 50.225 ;
        RECT 33.690 50.180 34.010 50.240 ;
        RECT 33.245 50.040 34.010 50.180 ;
        RECT 24.505 49.995 24.795 50.040 ;
        RECT 33.245 49.995 33.535 50.040 ;
        RECT 33.690 49.980 34.010 50.040 ;
        RECT 36.450 50.180 36.770 50.240 ;
        RECT 37.385 50.180 37.675 50.225 ;
        RECT 36.450 50.040 37.675 50.180 ;
        RECT 36.450 49.980 36.770 50.040 ;
        RECT 37.385 49.995 37.675 50.040 ;
        RECT 41.510 49.980 41.830 50.240 ;
        RECT 44.270 49.980 44.590 50.240 ;
        RECT 45.650 49.980 45.970 50.240 ;
        RECT 47.030 49.980 47.350 50.240 ;
        RECT 25.410 49.300 25.730 49.560 ;
        RECT 30.470 49.300 30.790 49.560 ;
        RECT 34.150 49.500 34.470 49.560 ;
        RECT 36.925 49.500 37.215 49.545 ;
        RECT 34.150 49.360 37.215 49.500 ;
        RECT 34.150 49.300 34.470 49.360 ;
        RECT 36.925 49.315 37.215 49.360 ;
        RECT 40.130 49.500 40.450 49.560 ;
        RECT 43.365 49.500 43.655 49.545 ;
        RECT 40.130 49.360 43.655 49.500 ;
        RECT 40.130 49.300 40.450 49.360 ;
        RECT 43.365 49.315 43.655 49.360 ;
        RECT 43.810 49.500 44.130 49.560 ;
        RECT 44.745 49.500 45.035 49.545 ;
        RECT 43.810 49.360 45.035 49.500 ;
        RECT 43.810 49.300 44.130 49.360 ;
        RECT 44.745 49.315 45.035 49.360 ;
        RECT 46.125 49.500 46.415 49.545 ;
        RECT 46.570 49.500 46.890 49.560 ;
        RECT 46.125 49.360 46.890 49.500 ;
        RECT 46.125 49.315 46.415 49.360 ;
        RECT 46.570 49.300 46.890 49.360 ;
        RECT 12.920 48.680 48.800 49.160 ;
        RECT 18.510 48.280 18.830 48.540 ;
        RECT 23.110 48.480 23.430 48.540 ;
        RECT 32.785 48.480 33.075 48.525 ;
        RECT 33.690 48.480 34.010 48.540 ;
        RECT 23.110 48.340 28.400 48.480 ;
        RECT 23.110 48.280 23.430 48.340 ;
        RECT 25.410 48.140 25.730 48.200 ;
        RECT 27.110 48.140 27.400 48.185 ;
        RECT 25.410 48.000 27.400 48.140 ;
        RECT 28.260 48.140 28.400 48.340 ;
        RECT 32.785 48.340 34.010 48.480 ;
        RECT 32.785 48.295 33.075 48.340 ;
        RECT 33.690 48.280 34.010 48.340 ;
        RECT 33.245 48.140 33.535 48.185 ;
        RECT 28.260 48.000 33.535 48.140 ;
        RECT 25.410 47.940 25.730 48.000 ;
        RECT 27.110 47.955 27.400 48.000 ;
        RECT 33.245 47.955 33.535 48.000 ;
        RECT 34.150 47.940 34.470 48.200 ;
        RECT 24.145 47.800 24.435 47.845 ;
        RECT 26.330 47.800 26.650 47.860 ;
        RECT 24.145 47.660 26.650 47.800 ;
        RECT 24.145 47.615 24.435 47.660 ;
        RECT 26.330 47.600 26.650 47.660 ;
        RECT 35.070 47.600 35.390 47.860 ;
        RECT 35.545 47.615 35.835 47.845 ;
        RECT 36.450 47.800 36.770 47.860 ;
        RECT 37.385 47.800 37.675 47.845 ;
        RECT 36.450 47.660 37.675 47.800 ;
        RECT 20.835 47.460 21.125 47.505 ;
        RECT 23.355 47.460 23.645 47.505 ;
        RECT 24.545 47.460 24.835 47.505 ;
        RECT 20.835 47.320 24.835 47.460 ;
        RECT 20.835 47.275 21.125 47.320 ;
        RECT 23.355 47.275 23.645 47.320 ;
        RECT 24.545 47.275 24.835 47.320 ;
        RECT 25.425 47.460 25.715 47.505 ;
        RECT 25.885 47.460 26.175 47.505 ;
        RECT 25.425 47.320 26.175 47.460 ;
        RECT 25.425 47.275 25.715 47.320 ;
        RECT 25.885 47.275 26.175 47.320 ;
        RECT 26.765 47.460 27.055 47.505 ;
        RECT 27.955 47.460 28.245 47.505 ;
        RECT 30.475 47.460 30.765 47.505 ;
        RECT 26.765 47.320 30.765 47.460 ;
        RECT 26.765 47.275 27.055 47.320 ;
        RECT 27.955 47.275 28.245 47.320 ;
        RECT 30.475 47.275 30.765 47.320 ;
        RECT 31.850 47.460 32.170 47.520 ;
        RECT 35.620 47.460 35.760 47.615 ;
        RECT 36.450 47.600 36.770 47.660 ;
        RECT 37.385 47.615 37.675 47.660 ;
        RECT 38.290 47.800 38.610 47.860 ;
        RECT 40.145 47.800 40.435 47.845 ;
        RECT 38.290 47.660 40.435 47.800 ;
        RECT 38.290 47.600 38.610 47.660 ;
        RECT 40.145 47.615 40.435 47.660 ;
        RECT 41.050 47.600 41.370 47.860 ;
        RECT 41.525 47.800 41.815 47.845 ;
        RECT 44.270 47.800 44.590 47.860 ;
        RECT 41.525 47.660 44.590 47.800 ;
        RECT 41.525 47.615 41.815 47.660 ;
        RECT 44.270 47.600 44.590 47.660 ;
        RECT 47.030 47.600 47.350 47.860 ;
        RECT 31.850 47.320 35.760 47.460 ;
        RECT 35.990 47.460 36.310 47.520 ;
        RECT 38.380 47.460 38.520 47.600 ;
        RECT 35.990 47.320 38.520 47.460 ;
        RECT 21.270 47.120 21.560 47.165 ;
        RECT 22.840 47.120 23.130 47.165 ;
        RECT 24.940 47.120 25.230 47.165 ;
        RECT 21.270 46.980 25.230 47.120 ;
        RECT 21.270 46.935 21.560 46.980 ;
        RECT 22.840 46.935 23.130 46.980 ;
        RECT 24.940 46.935 25.230 46.980 ;
        RECT 24.030 46.780 24.350 46.840 ;
        RECT 25.960 46.780 26.100 47.275 ;
        RECT 31.850 47.260 32.170 47.320 ;
        RECT 35.990 47.260 36.310 47.320 ;
        RECT 42.445 47.275 42.735 47.505 ;
        RECT 26.370 47.120 26.660 47.165 ;
        RECT 28.470 47.120 28.760 47.165 ;
        RECT 30.040 47.120 30.330 47.165 ;
        RECT 26.370 46.980 30.330 47.120 ;
        RECT 26.370 46.935 26.660 46.980 ;
        RECT 28.470 46.935 28.760 46.980 ;
        RECT 30.040 46.935 30.330 46.980 ;
        RECT 30.930 47.120 31.250 47.180 ;
        RECT 36.465 47.120 36.755 47.165 ;
        RECT 30.930 46.980 36.755 47.120 ;
        RECT 30.930 46.920 31.250 46.980 ;
        RECT 36.465 46.935 36.755 46.980 ;
        RECT 37.845 47.120 38.135 47.165 ;
        RECT 40.605 47.120 40.895 47.165 ;
        RECT 37.845 46.980 40.895 47.120 ;
        RECT 37.845 46.935 38.135 46.980 ;
        RECT 40.605 46.935 40.895 46.980 ;
        RECT 41.510 47.120 41.830 47.180 ;
        RECT 42.520 47.120 42.660 47.275 ;
        RECT 41.510 46.980 42.660 47.120 ;
        RECT 44.730 47.120 45.050 47.180 ;
        RECT 46.125 47.120 46.415 47.165 ;
        RECT 44.730 46.980 46.415 47.120 ;
        RECT 41.510 46.920 41.830 46.980 ;
        RECT 44.730 46.920 45.050 46.980 ;
        RECT 46.125 46.935 46.415 46.980 ;
        RECT 34.610 46.780 34.930 46.840 ;
        RECT 24.030 46.640 34.930 46.780 ;
        RECT 24.030 46.580 24.350 46.640 ;
        RECT 34.610 46.580 34.930 46.640 ;
        RECT 37.370 46.780 37.690 46.840 ;
        RECT 39.225 46.780 39.515 46.825 ;
        RECT 37.370 46.640 39.515 46.780 ;
        RECT 37.370 46.580 37.690 46.640 ;
        RECT 39.225 46.595 39.515 46.640 ;
        RECT 43.350 46.780 43.670 46.840 ;
        RECT 45.665 46.780 45.955 46.825 ;
        RECT 43.350 46.640 45.955 46.780 ;
        RECT 43.350 46.580 43.670 46.640 ;
        RECT 45.665 46.595 45.955 46.640 ;
        RECT 12.920 45.960 48.800 46.440 ;
        RECT 26.330 45.560 26.650 45.820 ;
        RECT 31.390 45.760 31.710 45.820 ;
        RECT 33.705 45.760 33.995 45.805 ;
        RECT 36.450 45.760 36.770 45.820 ;
        RECT 31.390 45.620 33.995 45.760 ;
        RECT 31.390 45.560 31.710 45.620 ;
        RECT 33.705 45.575 33.995 45.620 ;
        RECT 34.700 45.620 39.900 45.760 ;
        RECT 14.870 45.420 15.160 45.465 ;
        RECT 16.970 45.420 17.260 45.465 ;
        RECT 18.540 45.420 18.830 45.465 ;
        RECT 34.700 45.420 34.840 45.620 ;
        RECT 36.450 45.560 36.770 45.620 ;
        RECT 14.870 45.280 18.830 45.420 ;
        RECT 14.870 45.235 15.160 45.280 ;
        RECT 16.970 45.235 17.260 45.280 ;
        RECT 18.540 45.235 18.830 45.280 ;
        RECT 29.640 45.280 34.840 45.420 ;
        RECT 35.110 45.420 35.400 45.465 ;
        RECT 37.210 45.420 37.500 45.465 ;
        RECT 38.780 45.420 39.070 45.465 ;
        RECT 35.110 45.280 39.070 45.420 ;
        RECT 29.640 45.125 29.780 45.280 ;
        RECT 35.110 45.235 35.400 45.280 ;
        RECT 37.210 45.235 37.500 45.280 ;
        RECT 38.780 45.235 39.070 45.280 ;
        RECT 15.265 45.080 15.555 45.125 ;
        RECT 16.455 45.080 16.745 45.125 ;
        RECT 18.975 45.080 19.265 45.125 ;
        RECT 15.265 44.940 19.265 45.080 ;
        RECT 15.265 44.895 15.555 44.940 ;
        RECT 16.455 44.895 16.745 44.940 ;
        RECT 18.975 44.895 19.265 44.940 ;
        RECT 29.565 44.895 29.855 45.125 ;
        RECT 34.610 44.880 34.930 45.140 ;
        RECT 35.505 45.080 35.795 45.125 ;
        RECT 36.695 45.080 36.985 45.125 ;
        RECT 39.215 45.080 39.505 45.125 ;
        RECT 35.505 44.940 39.505 45.080 ;
        RECT 35.505 44.895 35.795 44.940 ;
        RECT 36.695 44.895 36.985 44.940 ;
        RECT 39.215 44.895 39.505 44.940 ;
        RECT 14.385 44.740 14.675 44.785 ;
        RECT 24.030 44.740 24.350 44.800 ;
        RECT 14.385 44.600 24.350 44.740 ;
        RECT 14.385 44.555 14.675 44.600 ;
        RECT 24.030 44.540 24.350 44.600 ;
        RECT 24.505 44.555 24.795 44.785 ;
        RECT 28.185 44.740 28.475 44.785 ;
        RECT 30.470 44.740 30.790 44.800 ;
        RECT 28.185 44.600 30.790 44.740 ;
        RECT 28.185 44.555 28.475 44.600 ;
        RECT 15.720 44.400 16.010 44.445 ;
        RECT 16.210 44.400 16.530 44.460 ;
        RECT 24.580 44.400 24.720 44.555 ;
        RECT 30.470 44.540 30.790 44.600 ;
        RECT 30.930 44.540 31.250 44.800 ;
        RECT 31.850 44.740 32.170 44.800 ;
        RECT 33.690 44.740 34.010 44.800 ;
        RECT 31.850 44.600 34.010 44.740 ;
        RECT 31.850 44.540 32.170 44.600 ;
        RECT 33.690 44.540 34.010 44.600 ;
        RECT 34.150 44.740 34.470 44.800 ;
        RECT 35.070 44.740 35.390 44.800 ;
        RECT 34.150 44.600 35.390 44.740 ;
        RECT 34.150 44.540 34.470 44.600 ;
        RECT 35.070 44.540 35.390 44.600 ;
        RECT 35.960 44.740 36.250 44.785 ;
        RECT 37.370 44.740 37.690 44.800 ;
        RECT 35.960 44.600 37.690 44.740 ;
        RECT 39.760 44.740 39.900 45.620 ;
        RECT 41.510 45.560 41.830 45.820 ;
        RECT 44.270 45.560 44.590 45.820 ;
        RECT 42.445 44.740 42.735 44.785 ;
        RECT 39.760 44.600 42.735 44.740 ;
        RECT 35.960 44.555 36.250 44.600 ;
        RECT 37.370 44.540 37.690 44.600 ;
        RECT 42.445 44.555 42.735 44.600 ;
        RECT 43.350 44.540 43.670 44.800 ;
        RECT 44.730 44.540 45.050 44.800 ;
        RECT 47.030 44.540 47.350 44.800 ;
        RECT 15.720 44.260 16.530 44.400 ;
        RECT 15.720 44.215 16.010 44.260 ;
        RECT 16.210 44.200 16.530 44.260 ;
        RECT 21.360 44.260 24.720 44.400 ;
        RECT 28.645 44.400 28.935 44.445 ;
        RECT 36.450 44.400 36.770 44.460 ;
        RECT 28.645 44.260 36.770 44.400 ;
        RECT 21.360 44.120 21.500 44.260 ;
        RECT 28.645 44.215 28.935 44.260 ;
        RECT 36.450 44.200 36.770 44.260 ;
        RECT 21.270 43.860 21.590 44.120 ;
        RECT 21.730 43.860 22.050 44.120 ;
        RECT 30.470 44.060 30.790 44.120 ;
        RECT 32.785 44.060 33.075 44.105 ;
        RECT 30.470 43.920 33.075 44.060 ;
        RECT 30.470 43.860 30.790 43.920 ;
        RECT 32.785 43.875 33.075 43.920 ;
        RECT 45.650 43.860 45.970 44.120 ;
        RECT 46.110 43.860 46.430 44.120 ;
        RECT 12.920 43.240 48.800 43.720 ;
        RECT 13.910 43.040 14.230 43.100 ;
        RECT 14.845 43.040 15.135 43.085 ;
        RECT 13.910 42.900 15.135 43.040 ;
        RECT 13.910 42.840 14.230 42.900 ;
        RECT 14.845 42.855 15.135 42.900 ;
        RECT 16.210 42.840 16.530 43.100 ;
        RECT 18.065 43.040 18.355 43.085 ;
        RECT 21.730 43.040 22.050 43.100 ;
        RECT 18.065 42.900 22.050 43.040 ;
        RECT 18.065 42.855 18.355 42.900 ;
        RECT 21.730 42.840 22.050 42.900 ;
        RECT 24.030 43.040 24.350 43.100 ;
        RECT 26.330 43.040 26.650 43.100 ;
        RECT 24.030 42.900 26.650 43.040 ;
        RECT 24.030 42.840 24.350 42.900 ;
        RECT 26.330 42.840 26.650 42.900 ;
        RECT 27.250 43.040 27.570 43.100 ;
        RECT 30.930 43.040 31.250 43.100 ;
        RECT 43.810 43.040 44.130 43.100 ;
        RECT 27.250 42.900 31.250 43.040 ;
        RECT 27.250 42.840 27.570 42.900 ;
        RECT 30.930 42.840 31.250 42.900 ;
        RECT 37.460 42.900 44.130 43.040 ;
        RECT 35.990 42.500 36.310 42.760 ;
        RECT 15.765 42.360 16.055 42.405 ;
        RECT 21.270 42.360 21.590 42.420 ;
        RECT 15.765 42.220 21.590 42.360 ;
        RECT 15.765 42.175 16.055 42.220 ;
        RECT 21.270 42.160 21.590 42.220 ;
        RECT 30.485 42.360 30.775 42.405 ;
        RECT 30.930 42.360 31.250 42.420 ;
        RECT 37.460 42.405 37.600 42.900 ;
        RECT 43.810 42.840 44.130 42.900 ;
        RECT 46.110 42.840 46.430 43.100 ;
        RECT 39.225 42.700 39.515 42.745 ;
        RECT 40.590 42.700 40.910 42.760 ;
        RECT 39.225 42.560 40.910 42.700 ;
        RECT 39.225 42.515 39.515 42.560 ;
        RECT 40.590 42.500 40.910 42.560 ;
        RECT 41.050 42.700 41.370 42.760 ;
        RECT 46.200 42.700 46.340 42.840 ;
        RECT 41.050 42.560 46.340 42.700 ;
        RECT 41.050 42.500 41.370 42.560 ;
        RECT 30.485 42.220 31.250 42.360 ;
        RECT 30.485 42.175 30.775 42.220 ;
        RECT 30.930 42.160 31.250 42.220 ;
        RECT 37.385 42.175 37.675 42.405 ;
        RECT 40.130 42.160 40.450 42.420 ;
        RECT 42.520 42.405 42.660 42.560 ;
        RECT 41.525 42.175 41.815 42.405 ;
        RECT 42.445 42.175 42.735 42.405 ;
        RECT 18.525 41.835 18.815 42.065 ;
        RECT 19.445 42.020 19.735 42.065 ;
        RECT 19.890 42.020 20.210 42.080 ;
        RECT 19.445 41.880 20.210 42.020 ;
        RECT 19.445 41.835 19.735 41.880 ;
        RECT 16.670 41.680 16.990 41.740 ;
        RECT 18.600 41.680 18.740 41.835 ;
        RECT 19.890 41.820 20.210 41.880 ;
        RECT 34.165 42.020 34.455 42.065 ;
        RECT 34.610 42.020 34.930 42.080 ;
        RECT 34.165 41.880 34.930 42.020 ;
        RECT 34.165 41.835 34.455 41.880 ;
        RECT 34.610 41.820 34.930 41.880 ;
        RECT 36.925 42.020 37.215 42.065 ;
        RECT 40.220 42.020 40.360 42.160 ;
        RECT 36.925 41.880 40.360 42.020 ;
        RECT 41.600 42.020 41.740 42.175 ;
        RECT 43.810 42.160 44.130 42.420 ;
        RECT 45.190 42.160 45.510 42.420 ;
        RECT 46.125 42.360 46.415 42.405 ;
        RECT 46.570 42.360 46.890 42.420 ;
        RECT 46.125 42.220 46.890 42.360 ;
        RECT 46.125 42.175 46.415 42.220 ;
        RECT 46.570 42.160 46.890 42.220 ;
        RECT 42.905 42.020 43.195 42.065 ;
        RECT 41.600 41.880 43.195 42.020 ;
        RECT 36.925 41.835 37.215 41.880 ;
        RECT 42.905 41.835 43.195 41.880 ;
        RECT 36.450 41.680 36.770 41.740 ;
        RECT 41.050 41.680 41.370 41.740 ;
        RECT 16.670 41.540 36.770 41.680 ;
        RECT 16.670 41.480 16.990 41.540 ;
        RECT 36.450 41.480 36.770 41.540 ;
        RECT 37.460 41.540 41.370 41.680 ;
        RECT 30.945 41.340 31.235 41.385 ;
        RECT 31.390 41.340 31.710 41.400 ;
        RECT 37.460 41.385 37.600 41.540 ;
        RECT 41.050 41.480 41.370 41.540 ;
        RECT 30.945 41.200 31.710 41.340 ;
        RECT 30.945 41.155 31.235 41.200 ;
        RECT 31.390 41.140 31.710 41.200 ;
        RECT 37.385 41.155 37.675 41.385 ;
        RECT 38.290 41.140 38.610 41.400 ;
        RECT 12.920 40.520 48.800 41.000 ;
        RECT 27.250 40.320 27.570 40.380 ;
        RECT 18.600 40.180 27.570 40.320 ;
        RECT 16.670 39.440 16.990 39.700 ;
        RECT 17.605 39.640 17.895 39.685 ;
        RECT 18.600 39.640 18.740 40.180 ;
        RECT 27.250 40.120 27.570 40.180 ;
        RECT 33.245 40.320 33.535 40.365 ;
        RECT 33.690 40.320 34.010 40.380 ;
        RECT 33.245 40.180 34.010 40.320 ;
        RECT 33.245 40.135 33.535 40.180 ;
        RECT 33.690 40.120 34.010 40.180 ;
        RECT 43.365 40.320 43.655 40.365 ;
        RECT 45.190 40.320 45.510 40.380 ;
        RECT 43.365 40.180 45.510 40.320 ;
        RECT 43.365 40.135 43.655 40.180 ;
        RECT 45.190 40.120 45.510 40.180 ;
        RECT 19.010 39.980 19.300 40.025 ;
        RECT 21.110 39.980 21.400 40.025 ;
        RECT 22.680 39.980 22.970 40.025 ;
        RECT 19.010 39.840 22.970 39.980 ;
        RECT 19.010 39.795 19.300 39.840 ;
        RECT 21.110 39.795 21.400 39.840 ;
        RECT 22.680 39.795 22.970 39.840 ;
        RECT 25.425 39.795 25.715 40.025 ;
        RECT 26.830 39.980 27.120 40.025 ;
        RECT 28.930 39.980 29.220 40.025 ;
        RECT 30.500 39.980 30.790 40.025 ;
        RECT 26.830 39.840 30.790 39.980 ;
        RECT 26.830 39.795 27.120 39.840 ;
        RECT 28.930 39.795 29.220 39.840 ;
        RECT 30.500 39.795 30.790 39.840 ;
        RECT 17.605 39.500 18.740 39.640 ;
        RECT 19.405 39.640 19.695 39.685 ;
        RECT 20.595 39.640 20.885 39.685 ;
        RECT 23.115 39.640 23.405 39.685 ;
        RECT 19.405 39.500 23.405 39.640 ;
        RECT 17.605 39.455 17.895 39.500 ;
        RECT 19.405 39.455 19.695 39.500 ;
        RECT 20.595 39.455 20.885 39.500 ;
        RECT 23.115 39.455 23.405 39.500 ;
        RECT 18.525 39.300 18.815 39.345 ;
        RECT 21.270 39.300 21.590 39.360 ;
        RECT 24.030 39.300 24.350 39.360 ;
        RECT 18.525 39.160 24.350 39.300 ;
        RECT 25.500 39.300 25.640 39.795 ;
        RECT 35.070 39.780 35.390 40.040 ;
        RECT 41.970 39.980 42.290 40.040 ;
        RECT 46.570 39.980 46.890 40.040 ;
        RECT 39.760 39.840 46.890 39.980 ;
        RECT 26.330 39.440 26.650 39.700 ;
        RECT 39.760 39.685 39.900 39.840 ;
        RECT 41.970 39.780 42.290 39.840 ;
        RECT 46.570 39.780 46.890 39.840 ;
        RECT 27.225 39.640 27.515 39.685 ;
        RECT 28.415 39.640 28.705 39.685 ;
        RECT 30.935 39.640 31.225 39.685 ;
        RECT 27.225 39.500 31.225 39.640 ;
        RECT 27.225 39.455 27.515 39.500 ;
        RECT 28.415 39.455 28.705 39.500 ;
        RECT 30.935 39.455 31.225 39.500 ;
        RECT 39.685 39.455 39.975 39.685 ;
        RECT 40.145 39.640 40.435 39.685 ;
        RECT 42.890 39.640 43.210 39.700 ;
        RECT 40.145 39.500 43.210 39.640 ;
        RECT 40.145 39.455 40.435 39.500 ;
        RECT 42.890 39.440 43.210 39.500 ;
        RECT 34.610 39.300 34.930 39.360 ;
        RECT 25.500 39.160 35.760 39.300 ;
        RECT 18.525 39.115 18.815 39.160 ;
        RECT 21.270 39.100 21.590 39.160 ;
        RECT 24.030 39.100 24.350 39.160 ;
        RECT 34.610 39.100 34.930 39.160 ;
        RECT 35.620 39.020 35.760 39.160 ;
        RECT 39.225 39.115 39.515 39.345 ;
        RECT 40.605 39.115 40.895 39.345 ;
        RECT 41.050 39.300 41.370 39.360 ;
        RECT 41.525 39.300 41.815 39.345 ;
        RECT 41.050 39.160 41.815 39.300 ;
        RECT 19.890 39.005 20.210 39.020 ;
        RECT 19.860 38.960 20.210 39.005 ;
        RECT 27.680 38.960 27.970 39.005 ;
        RECT 34.150 38.960 34.470 39.020 ;
        RECT 19.455 38.820 27.480 38.960 ;
        RECT 19.860 38.775 20.210 38.820 ;
        RECT 19.890 38.760 20.210 38.775 ;
        RECT 14.370 38.420 14.690 38.680 ;
        RECT 16.225 38.620 16.515 38.665 ;
        RECT 18.970 38.620 19.290 38.680 ;
        RECT 16.225 38.480 19.290 38.620 ;
        RECT 27.340 38.620 27.480 38.820 ;
        RECT 27.680 38.820 34.470 38.960 ;
        RECT 27.680 38.775 27.970 38.820 ;
        RECT 34.150 38.760 34.470 38.820 ;
        RECT 35.530 38.960 35.850 39.020 ;
        RECT 36.925 38.960 37.215 39.005 ;
        RECT 35.530 38.820 37.215 38.960 ;
        RECT 39.300 38.960 39.440 39.115 ;
        RECT 40.680 38.960 40.820 39.115 ;
        RECT 41.050 39.100 41.370 39.160 ;
        RECT 41.525 39.115 41.815 39.160 ;
        RECT 42.445 39.300 42.735 39.345 ;
        RECT 43.810 39.300 44.130 39.360 ;
        RECT 42.445 39.160 44.130 39.300 ;
        RECT 42.445 39.115 42.735 39.160 ;
        RECT 43.810 39.100 44.130 39.160 ;
        RECT 44.270 39.100 44.590 39.360 ;
        RECT 45.650 39.100 45.970 39.360 ;
        RECT 46.110 39.300 46.430 39.360 ;
        RECT 46.585 39.300 46.875 39.345 ;
        RECT 46.110 39.160 46.875 39.300 ;
        RECT 46.110 39.100 46.430 39.160 ;
        RECT 46.585 39.115 46.875 39.160 ;
        RECT 41.985 38.960 42.275 39.005 ;
        RECT 39.300 38.820 39.900 38.960 ;
        RECT 40.680 38.820 42.275 38.960 ;
        RECT 35.530 38.760 35.850 38.820 ;
        RECT 36.925 38.775 37.215 38.820 ;
        RECT 33.690 38.620 34.010 38.680 ;
        RECT 34.625 38.620 34.915 38.665 ;
        RECT 27.340 38.480 34.915 38.620 ;
        RECT 16.225 38.435 16.515 38.480 ;
        RECT 18.970 38.420 19.290 38.480 ;
        RECT 33.690 38.420 34.010 38.480 ;
        RECT 34.625 38.435 34.915 38.480 ;
        RECT 38.305 38.620 38.595 38.665 ;
        RECT 39.210 38.620 39.530 38.680 ;
        RECT 38.305 38.480 39.530 38.620 ;
        RECT 39.760 38.620 39.900 38.820 ;
        RECT 41.985 38.775 42.275 38.820 ;
        RECT 44.360 38.620 44.500 39.100 ;
        RECT 39.760 38.480 44.500 38.620 ;
        RECT 38.305 38.435 38.595 38.480 ;
        RECT 39.210 38.420 39.530 38.480 ;
        RECT 12.920 37.800 48.800 38.280 ;
        RECT 34.150 37.400 34.470 37.660 ;
        RECT 36.450 37.600 36.770 37.660 ;
        RECT 41.065 37.600 41.355 37.645 ;
        RECT 36.450 37.460 41.355 37.600 ;
        RECT 36.450 37.400 36.770 37.460 ;
        RECT 41.065 37.415 41.355 37.460 ;
        RECT 46.125 37.415 46.415 37.645 ;
        RECT 14.370 37.260 14.690 37.320 ;
        RECT 19.950 37.260 20.240 37.305 ;
        RECT 14.370 37.120 20.240 37.260 ;
        RECT 14.370 37.060 14.690 37.120 ;
        RECT 19.950 37.075 20.240 37.120 ;
        RECT 24.950 37.060 25.270 37.320 ;
        RECT 46.200 37.260 46.340 37.415 ;
        RECT 44.820 37.120 46.340 37.260 ;
        RECT 44.820 36.980 44.960 37.120 ;
        RECT 21.270 36.720 21.590 36.980 ;
        RECT 39.210 36.720 39.530 36.980 ;
        RECT 40.130 36.720 40.450 36.980 ;
        RECT 44.730 36.720 45.050 36.980 ;
        RECT 45.665 36.920 45.955 36.965 ;
        RECT 46.110 36.920 46.430 36.980 ;
        RECT 45.665 36.780 46.430 36.920 ;
        RECT 45.665 36.735 45.955 36.780 ;
        RECT 46.110 36.720 46.430 36.780 ;
        RECT 47.030 36.720 47.350 36.980 ;
        RECT 16.695 36.580 16.985 36.625 ;
        RECT 19.215 36.580 19.505 36.625 ;
        RECT 20.405 36.580 20.695 36.625 ;
        RECT 16.695 36.440 20.695 36.580 ;
        RECT 16.695 36.395 16.985 36.440 ;
        RECT 19.215 36.395 19.505 36.440 ;
        RECT 20.405 36.395 20.695 36.440 ;
        RECT 31.390 36.580 31.710 36.640 ;
        RECT 36.925 36.580 37.215 36.625 ;
        RECT 31.390 36.440 37.215 36.580 ;
        RECT 31.390 36.380 31.710 36.440 ;
        RECT 36.925 36.395 37.215 36.440 ;
        RECT 17.130 36.240 17.420 36.285 ;
        RECT 18.700 36.240 18.990 36.285 ;
        RECT 20.800 36.240 21.090 36.285 ;
        RECT 17.130 36.100 21.090 36.240 ;
        RECT 17.130 36.055 17.420 36.100 ;
        RECT 18.700 36.055 18.990 36.100 ;
        RECT 20.800 36.055 21.090 36.100 ;
        RECT 14.370 35.700 14.690 35.960 ;
        RECT 30.930 35.900 31.250 35.960 ;
        RECT 31.405 35.900 31.695 35.945 ;
        RECT 30.930 35.760 31.695 35.900 ;
        RECT 30.930 35.700 31.250 35.760 ;
        RECT 31.405 35.715 31.695 35.760 ;
        RECT 35.990 35.900 36.310 35.960 ;
        RECT 39.225 35.900 39.515 35.945 ;
        RECT 35.990 35.760 39.515 35.900 ;
        RECT 35.990 35.700 36.310 35.760 ;
        RECT 39.225 35.715 39.515 35.760 ;
        RECT 42.430 35.900 42.750 35.960 ;
        RECT 45.665 35.900 45.955 35.945 ;
        RECT 42.430 35.760 45.955 35.900 ;
        RECT 42.430 35.700 42.750 35.760 ;
        RECT 45.665 35.715 45.955 35.760 ;
        RECT 12.920 35.080 48.800 35.560 ;
        RECT 18.970 34.680 19.290 34.940 ;
        RECT 27.250 34.680 27.570 34.940 ;
        RECT 27.710 34.880 28.030 34.940 ;
        RECT 29.565 34.880 29.855 34.925 ;
        RECT 27.710 34.740 29.855 34.880 ;
        RECT 27.710 34.680 28.030 34.740 ;
        RECT 29.565 34.695 29.855 34.740 ;
        RECT 38.290 34.680 38.610 34.940 ;
        RECT 45.650 34.880 45.970 34.940 ;
        RECT 46.585 34.880 46.875 34.925 ;
        RECT 45.650 34.740 46.875 34.880 ;
        RECT 45.650 34.680 45.970 34.740 ;
        RECT 46.585 34.695 46.875 34.740 ;
        RECT 28.645 34.540 28.935 34.585 ;
        RECT 31.850 34.540 32.170 34.600 ;
        RECT 35.990 34.540 36.310 34.600 ;
        RECT 28.645 34.400 32.170 34.540 ;
        RECT 28.645 34.355 28.935 34.400 ;
        RECT 14.370 34.200 14.690 34.260 ;
        RECT 15.765 34.200 16.055 34.245 ;
        RECT 28.720 34.200 28.860 34.355 ;
        RECT 31.850 34.340 32.170 34.400 ;
        RECT 34.700 34.400 36.310 34.540 ;
        RECT 14.370 34.060 16.055 34.200 ;
        RECT 14.370 34.000 14.690 34.060 ;
        RECT 15.765 34.015 16.055 34.060 ;
        RECT 27.340 34.060 28.860 34.200 ;
        RECT 29.105 34.200 29.395 34.245 ;
        RECT 34.700 34.200 34.840 34.400 ;
        RECT 35.990 34.340 36.310 34.400 ;
        RECT 44.270 34.340 44.590 34.600 ;
        RECT 29.105 34.060 34.840 34.200 ;
        RECT 22.190 33.660 22.510 33.920 ;
        RECT 27.340 33.905 27.480 34.060 ;
        RECT 29.105 34.015 29.395 34.060 ;
        RECT 35.070 34.000 35.390 34.260 ;
        RECT 44.360 34.200 44.500 34.340 ;
        RECT 37.920 34.060 44.500 34.200 ;
        RECT 26.345 33.675 26.635 33.905 ;
        RECT 27.265 33.675 27.555 33.905 ;
        RECT 26.420 33.520 26.560 33.675 ;
        RECT 27.710 33.660 28.030 33.920 ;
        RECT 30.025 33.860 30.315 33.905 ;
        RECT 30.470 33.860 30.790 33.920 ;
        RECT 30.025 33.720 30.790 33.860 ;
        RECT 30.025 33.675 30.315 33.720 ;
        RECT 30.470 33.660 30.790 33.720 ;
        RECT 31.390 33.660 31.710 33.920 ;
        RECT 37.920 33.905 38.060 34.060 ;
        RECT 37.845 33.675 38.135 33.905 ;
        RECT 38.765 33.860 39.055 33.905 ;
        RECT 40.605 33.860 40.895 33.905 ;
        RECT 41.050 33.860 41.370 33.920 ;
        RECT 41.600 33.905 41.740 34.060 ;
        RECT 38.765 33.720 41.370 33.860 ;
        RECT 38.765 33.675 39.055 33.720 ;
        RECT 40.605 33.675 40.895 33.720 ;
        RECT 41.050 33.660 41.370 33.720 ;
        RECT 41.525 33.675 41.815 33.905 ;
        RECT 41.970 33.660 42.290 33.920 ;
        RECT 43.365 33.675 43.655 33.905 ;
        RECT 31.865 33.520 32.155 33.565 ;
        RECT 26.420 33.380 32.155 33.520 ;
        RECT 31.865 33.335 32.155 33.380 ;
        RECT 40.145 33.520 40.435 33.565 ;
        RECT 42.430 33.520 42.750 33.580 ;
        RECT 43.440 33.520 43.580 33.675 ;
        RECT 44.270 33.660 44.590 33.920 ;
        RECT 44.730 33.860 45.050 33.920 ;
        RECT 45.665 33.860 45.955 33.905 ;
        RECT 44.730 33.720 45.955 33.860 ;
        RECT 44.730 33.660 45.050 33.720 ;
        RECT 45.665 33.675 45.955 33.720 ;
        RECT 45.190 33.520 45.510 33.580 ;
        RECT 40.145 33.380 42.750 33.520 ;
        RECT 40.145 33.335 40.435 33.380 ;
        RECT 42.430 33.320 42.750 33.380 ;
        RECT 42.980 33.380 45.510 33.520 ;
        RECT 19.430 32.980 19.750 33.240 ;
        RECT 36.925 33.180 37.215 33.225 ;
        RECT 37.830 33.180 38.150 33.240 ;
        RECT 36.925 33.040 38.150 33.180 ;
        RECT 36.925 32.995 37.215 33.040 ;
        RECT 37.830 32.980 38.150 33.040 ;
        RECT 40.590 33.180 40.910 33.240 ;
        RECT 42.980 33.225 43.120 33.380 ;
        RECT 45.190 33.320 45.510 33.380 ;
        RECT 41.065 33.180 41.355 33.225 ;
        RECT 40.590 33.040 41.355 33.180 ;
        RECT 40.590 32.980 40.910 33.040 ;
        RECT 41.065 32.995 41.355 33.040 ;
        RECT 42.905 32.995 43.195 33.225 ;
        RECT 12.920 32.360 48.800 32.840 ;
        RECT 13.910 32.160 14.230 32.220 ;
        RECT 14.845 32.160 15.135 32.205 ;
        RECT 13.910 32.020 15.135 32.160 ;
        RECT 13.910 31.960 14.230 32.020 ;
        RECT 14.845 31.975 15.135 32.020 ;
        RECT 18.525 32.160 18.815 32.205 ;
        RECT 19.430 32.160 19.750 32.220 ;
        RECT 18.525 32.020 19.750 32.160 ;
        RECT 18.525 31.975 18.815 32.020 ;
        RECT 19.430 31.960 19.750 32.020 ;
        RECT 27.710 32.160 28.030 32.220 ;
        RECT 34.610 32.160 34.930 32.220 ;
        RECT 27.710 32.020 34.930 32.160 ;
        RECT 27.710 31.960 28.030 32.020 ;
        RECT 34.610 31.960 34.930 32.020 ;
        RECT 44.270 32.160 44.590 32.220 ;
        RECT 46.585 32.160 46.875 32.205 ;
        RECT 44.270 32.020 46.875 32.160 ;
        RECT 44.270 31.960 44.590 32.020 ;
        RECT 46.585 31.975 46.875 32.020 ;
        RECT 22.160 31.820 22.450 31.865 ;
        RECT 25.870 31.820 26.190 31.880 ;
        RECT 27.250 31.820 27.570 31.880 ;
        RECT 42.430 31.820 42.750 31.880 ;
        RECT 22.160 31.680 27.570 31.820 ;
        RECT 22.160 31.635 22.450 31.680 ;
        RECT 25.870 31.620 26.190 31.680 ;
        RECT 27.250 31.620 27.570 31.680 ;
        RECT 40.220 31.680 42.750 31.820 ;
        RECT 14.370 31.480 14.690 31.540 ;
        RECT 15.765 31.480 16.055 31.525 ;
        RECT 14.370 31.340 16.055 31.480 ;
        RECT 14.370 31.280 14.690 31.340 ;
        RECT 15.765 31.295 16.055 31.340 ;
        RECT 30.025 31.480 30.315 31.525 ;
        RECT 32.325 31.480 32.615 31.525 ;
        RECT 30.025 31.340 32.615 31.480 ;
        RECT 30.025 31.295 30.315 31.340 ;
        RECT 32.325 31.295 32.615 31.340 ;
        RECT 38.290 31.480 38.610 31.540 ;
        RECT 40.220 31.525 40.360 31.680 ;
        RECT 42.430 31.620 42.750 31.680 ;
        RECT 39.685 31.480 39.975 31.525 ;
        RECT 38.290 31.340 39.975 31.480 ;
        RECT 38.290 31.280 38.610 31.340 ;
        RECT 39.685 31.295 39.975 31.340 ;
        RECT 40.145 31.295 40.435 31.525 ;
        RECT 40.590 31.280 40.910 31.540 ;
        RECT 43.365 31.480 43.655 31.525 ;
        RECT 43.810 31.480 44.130 31.540 ;
        RECT 43.365 31.340 44.130 31.480 ;
        RECT 43.365 31.295 43.655 31.340 ;
        RECT 43.810 31.280 44.130 31.340 ;
        RECT 44.270 31.280 44.590 31.540 ;
        RECT 45.665 31.480 45.955 31.525 ;
        RECT 46.110 31.480 46.430 31.540 ;
        RECT 45.665 31.340 46.430 31.480 ;
        RECT 45.665 31.295 45.955 31.340 ;
        RECT 46.110 31.280 46.430 31.340 ;
        RECT 18.985 31.140 19.275 31.185 ;
        RECT 19.430 31.140 19.750 31.200 ;
        RECT 18.985 31.000 19.750 31.140 ;
        RECT 18.985 30.955 19.275 31.000 ;
        RECT 19.430 30.940 19.750 31.000 ;
        RECT 19.890 30.940 20.210 31.200 ;
        RECT 20.825 30.955 21.115 31.185 ;
        RECT 21.705 31.140 21.995 31.185 ;
        RECT 22.895 31.140 23.185 31.185 ;
        RECT 25.415 31.140 25.705 31.185 ;
        RECT 21.705 31.000 25.705 31.140 ;
        RECT 21.705 30.955 21.995 31.000 ;
        RECT 22.895 30.955 23.185 31.000 ;
        RECT 25.415 30.955 25.705 31.000 ;
        RECT 30.485 30.955 30.775 31.185 ;
        RECT 31.405 31.140 31.695 31.185 ;
        RECT 33.690 31.140 34.010 31.200 ;
        RECT 31.405 31.000 34.010 31.140 ;
        RECT 31.405 30.955 31.695 31.000 ;
        RECT 14.370 30.800 14.690 30.860 ;
        RECT 20.900 30.800 21.040 30.955 ;
        RECT 14.370 30.660 21.040 30.800 ;
        RECT 21.310 30.800 21.600 30.845 ;
        RECT 23.410 30.800 23.700 30.845 ;
        RECT 24.980 30.800 25.270 30.845 ;
        RECT 21.310 30.660 25.270 30.800 ;
        RECT 14.370 30.600 14.690 30.660 ;
        RECT 21.310 30.615 21.600 30.660 ;
        RECT 23.410 30.615 23.700 30.660 ;
        RECT 24.980 30.615 25.270 30.660 ;
        RECT 27.250 30.800 27.570 30.860 ;
        RECT 28.185 30.800 28.475 30.845 ;
        RECT 27.250 30.660 28.475 30.800 ;
        RECT 30.560 30.800 30.700 30.955 ;
        RECT 33.690 30.940 34.010 31.000 ;
        RECT 34.150 31.140 34.470 31.200 ;
        RECT 35.085 31.140 35.375 31.185 ;
        RECT 34.150 31.000 35.375 31.140 ;
        RECT 34.150 30.940 34.470 31.000 ;
        RECT 35.085 30.955 35.375 31.000 ;
        RECT 41.065 31.140 41.355 31.185 ;
        RECT 44.730 31.140 45.050 31.200 ;
        RECT 41.065 31.000 45.050 31.140 ;
        RECT 41.065 30.955 41.355 31.000 ;
        RECT 44.730 30.940 45.050 31.000 ;
        RECT 35.990 30.800 36.310 30.860 ;
        RECT 41.985 30.800 42.275 30.845 ;
        RECT 30.560 30.660 42.275 30.800 ;
        RECT 27.250 30.600 27.570 30.660 ;
        RECT 28.185 30.615 28.475 30.660 ;
        RECT 35.990 30.600 36.310 30.660 ;
        RECT 41.985 30.615 42.275 30.660 ;
        RECT 16.670 30.260 16.990 30.520 ;
        RECT 12.920 29.640 48.800 30.120 ;
        RECT 21.285 29.440 21.575 29.485 ;
        RECT 22.190 29.440 22.510 29.500 ;
        RECT 21.285 29.300 22.510 29.440 ;
        RECT 21.285 29.255 21.575 29.300 ;
        RECT 22.190 29.240 22.510 29.300 ;
        RECT 36.005 29.440 36.295 29.485 ;
        RECT 36.910 29.440 37.230 29.500 ;
        RECT 36.005 29.300 37.230 29.440 ;
        RECT 36.005 29.255 36.295 29.300 ;
        RECT 36.910 29.240 37.230 29.300 ;
        RECT 42.890 29.440 43.210 29.500 ;
        RECT 43.825 29.440 44.115 29.485 ;
        RECT 42.890 29.300 44.115 29.440 ;
        RECT 42.890 29.240 43.210 29.300 ;
        RECT 43.825 29.255 44.115 29.300 ;
        RECT 14.870 29.100 15.160 29.145 ;
        RECT 16.970 29.100 17.260 29.145 ;
        RECT 18.540 29.100 18.830 29.145 ;
        RECT 14.870 28.960 18.830 29.100 ;
        RECT 14.870 28.915 15.160 28.960 ;
        RECT 16.970 28.915 17.260 28.960 ;
        RECT 18.540 28.915 18.830 28.960 ;
        RECT 26.830 29.100 27.120 29.145 ;
        RECT 28.930 29.100 29.220 29.145 ;
        RECT 30.500 29.100 30.790 29.145 ;
        RECT 26.830 28.960 30.790 29.100 ;
        RECT 26.830 28.915 27.120 28.960 ;
        RECT 28.930 28.915 29.220 28.960 ;
        RECT 30.500 28.915 30.790 28.960 ;
        RECT 35.530 28.900 35.850 29.160 ;
        RECT 14.370 28.560 14.690 28.820 ;
        RECT 15.265 28.760 15.555 28.805 ;
        RECT 16.455 28.760 16.745 28.805 ;
        RECT 18.975 28.760 19.265 28.805 ;
        RECT 15.265 28.620 19.265 28.760 ;
        RECT 15.265 28.575 15.555 28.620 ;
        RECT 16.455 28.575 16.745 28.620 ;
        RECT 18.975 28.575 19.265 28.620 ;
        RECT 27.225 28.760 27.515 28.805 ;
        RECT 28.415 28.760 28.705 28.805 ;
        RECT 30.935 28.760 31.225 28.805 ;
        RECT 27.225 28.620 31.225 28.760 ;
        RECT 27.225 28.575 27.515 28.620 ;
        RECT 28.415 28.575 28.705 28.620 ;
        RECT 30.935 28.575 31.225 28.620 ;
        RECT 33.705 28.760 33.995 28.805 ;
        RECT 34.610 28.760 34.930 28.820 ;
        RECT 33.705 28.620 34.930 28.760 ;
        RECT 33.705 28.575 33.995 28.620 ;
        RECT 34.610 28.560 34.930 28.620 ;
        RECT 42.430 28.760 42.750 28.820 ;
        RECT 42.430 28.620 46.340 28.760 ;
        RECT 42.430 28.560 42.750 28.620 ;
        RECT 14.460 28.420 14.600 28.560 ;
        RECT 21.270 28.420 21.590 28.480 ;
        RECT 26.345 28.420 26.635 28.465 ;
        RECT 14.460 28.280 26.635 28.420 ;
        RECT 21.270 28.220 21.590 28.280 ;
        RECT 26.345 28.235 26.635 28.280 ;
        RECT 27.680 28.235 27.970 28.465 ;
        RECT 15.720 28.080 16.010 28.125 ;
        RECT 16.670 28.080 16.990 28.140 ;
        RECT 15.720 27.940 16.990 28.080 ;
        RECT 15.720 27.895 16.010 27.940 ;
        RECT 16.670 27.880 16.990 27.940 ;
        RECT 26.420 27.740 26.560 28.235 ;
        RECT 27.250 28.080 27.570 28.140 ;
        RECT 27.800 28.080 27.940 28.235 ;
        RECT 40.130 28.220 40.450 28.480 ;
        RECT 42.890 28.420 43.210 28.480 ;
        RECT 44.745 28.420 45.035 28.465 ;
        RECT 42.890 28.280 45.035 28.420 ;
        RECT 42.890 28.220 43.210 28.280 ;
        RECT 44.745 28.235 45.035 28.280 ;
        RECT 45.190 28.220 45.510 28.480 ;
        RECT 45.650 28.220 45.970 28.480 ;
        RECT 46.200 28.465 46.340 28.620 ;
        RECT 46.125 28.235 46.415 28.465 ;
        RECT 27.250 27.940 27.940 28.080 ;
        RECT 27.250 27.880 27.570 27.940 ;
        RECT 31.390 27.740 31.710 27.800 ;
        RECT 26.420 27.600 31.710 27.740 ;
        RECT 31.390 27.540 31.710 27.600 ;
        RECT 33.245 27.740 33.535 27.785 ;
        RECT 34.150 27.740 34.470 27.800 ;
        RECT 33.245 27.600 34.470 27.740 ;
        RECT 33.245 27.555 33.535 27.600 ;
        RECT 34.150 27.540 34.470 27.600 ;
        RECT 41.050 27.740 41.370 27.800 ;
        RECT 43.365 27.740 43.655 27.785 ;
        RECT 41.050 27.600 43.655 27.740 ;
        RECT 41.050 27.540 41.370 27.600 ;
        RECT 43.365 27.555 43.655 27.600 ;
        RECT 12.920 26.920 48.800 27.400 ;
        RECT 41.050 26.520 41.370 26.780 ;
        RECT 44.730 26.520 45.050 26.780 ;
        RECT 35.990 26.380 36.310 26.440 ;
        RECT 31.020 26.240 36.310 26.380 ;
        RECT 15.765 26.040 16.055 26.085 ;
        RECT 22.190 26.040 22.510 26.100 ;
        RECT 15.765 25.900 22.510 26.040 ;
        RECT 15.765 25.855 16.055 25.900 ;
        RECT 22.190 25.840 22.510 25.900 ;
        RECT 24.965 26.040 25.255 26.085 ;
        RECT 27.265 26.040 27.555 26.085 ;
        RECT 24.965 25.900 27.555 26.040 ;
        RECT 24.965 25.855 25.255 25.900 ;
        RECT 27.265 25.855 27.555 25.900 ;
        RECT 14.370 25.700 14.690 25.760 ;
        RECT 17.145 25.700 17.435 25.745 ;
        RECT 14.370 25.560 17.435 25.700 ;
        RECT 14.370 25.500 14.690 25.560 ;
        RECT 17.145 25.515 17.435 25.560 ;
        RECT 21.730 25.500 22.050 25.760 ;
        RECT 25.870 25.500 26.190 25.760 ;
        RECT 26.805 25.700 27.095 25.745 ;
        RECT 31.020 25.700 31.160 26.240 ;
        RECT 35.990 26.180 36.310 26.240 ;
        RECT 45.190 26.380 45.510 26.440 ;
        RECT 47.045 26.380 47.335 26.425 ;
        RECT 45.190 26.240 47.335 26.380 ;
        RECT 45.190 26.180 45.510 26.240 ;
        RECT 47.045 26.195 47.335 26.240 ;
        RECT 31.390 25.840 31.710 26.100 ;
        RECT 32.740 26.040 33.030 26.085 ;
        RECT 36.910 26.040 37.230 26.100 ;
        RECT 32.740 25.900 36.680 26.040 ;
        RECT 32.740 25.855 33.030 25.900 ;
        RECT 26.805 25.560 31.160 25.700 ;
        RECT 32.285 25.700 32.575 25.745 ;
        RECT 33.475 25.700 33.765 25.745 ;
        RECT 35.995 25.700 36.285 25.745 ;
        RECT 32.285 25.560 36.285 25.700 ;
        RECT 26.805 25.515 27.095 25.560 ;
        RECT 32.285 25.515 32.575 25.560 ;
        RECT 33.475 25.515 33.765 25.560 ;
        RECT 35.995 25.515 36.285 25.560 ;
        RECT 13.910 25.360 14.230 25.420 ;
        RECT 14.845 25.360 15.135 25.405 ;
        RECT 13.910 25.220 15.135 25.360 ;
        RECT 13.910 25.160 14.230 25.220 ;
        RECT 14.845 25.175 15.135 25.220 ;
        RECT 19.430 25.360 19.750 25.420 ;
        RECT 31.890 25.360 32.180 25.405 ;
        RECT 33.990 25.360 34.280 25.405 ;
        RECT 35.560 25.360 35.850 25.405 ;
        RECT 19.430 25.220 31.620 25.360 ;
        RECT 19.430 25.160 19.750 25.220 ;
        RECT 18.970 25.020 19.290 25.080 ;
        RECT 20.365 25.020 20.655 25.065 ;
        RECT 18.970 24.880 20.655 25.020 ;
        RECT 18.970 24.820 19.290 24.880 ;
        RECT 20.365 24.835 20.655 24.880 ;
        RECT 29.105 25.020 29.395 25.065 ;
        RECT 30.470 25.020 30.790 25.080 ;
        RECT 29.105 24.880 30.790 25.020 ;
        RECT 31.480 25.020 31.620 25.220 ;
        RECT 31.890 25.220 35.850 25.360 ;
        RECT 36.540 25.360 36.680 25.900 ;
        RECT 36.910 25.900 42.200 26.040 ;
        RECT 36.910 25.840 37.230 25.900 ;
        RECT 37.830 25.700 38.150 25.760 ;
        RECT 42.060 25.745 42.200 25.900 ;
        RECT 43.350 25.840 43.670 26.100 ;
        RECT 44.730 26.040 45.050 26.100 ;
        RECT 45.665 26.040 45.955 26.085 ;
        RECT 44.730 25.900 45.955 26.040 ;
        RECT 44.730 25.840 45.050 25.900 ;
        RECT 45.665 25.855 45.955 25.900 ;
        RECT 41.525 25.700 41.815 25.745 ;
        RECT 37.830 25.560 41.815 25.700 ;
        RECT 37.830 25.500 38.150 25.560 ;
        RECT 41.525 25.515 41.815 25.560 ;
        RECT 41.985 25.515 42.275 25.745 ;
        RECT 42.890 25.700 43.210 25.760 ;
        RECT 46.110 25.700 46.430 25.760 ;
        RECT 42.890 25.560 46.430 25.700 ;
        RECT 42.890 25.500 43.210 25.560 ;
        RECT 46.110 25.500 46.430 25.560 ;
        RECT 39.225 25.360 39.515 25.405 ;
        RECT 36.540 25.220 39.515 25.360 ;
        RECT 31.890 25.175 32.180 25.220 ;
        RECT 33.990 25.175 34.280 25.220 ;
        RECT 35.560 25.175 35.850 25.220 ;
        RECT 39.225 25.175 39.515 25.220 ;
        RECT 44.285 25.360 44.575 25.405 ;
        RECT 47.030 25.360 47.350 25.420 ;
        RECT 44.285 25.220 47.350 25.360 ;
        RECT 44.285 25.175 44.575 25.220 ;
        RECT 47.030 25.160 47.350 25.220 ;
        RECT 37.830 25.020 38.150 25.080 ;
        RECT 31.480 24.880 38.150 25.020 ;
        RECT 29.105 24.835 29.395 24.880 ;
        RECT 30.470 24.820 30.790 24.880 ;
        RECT 37.830 24.820 38.150 24.880 ;
        RECT 38.305 25.020 38.595 25.065 ;
        RECT 40.130 25.020 40.450 25.080 ;
        RECT 38.305 24.880 40.450 25.020 ;
        RECT 38.305 24.835 38.595 24.880 ;
        RECT 40.130 24.820 40.450 24.880 ;
        RECT 43.810 25.020 44.130 25.080 ;
        RECT 45.665 25.020 45.955 25.065 ;
        RECT 43.810 24.880 45.955 25.020 ;
        RECT 43.810 24.820 44.130 24.880 ;
        RECT 45.665 24.835 45.955 24.880 ;
        RECT 12.920 24.200 48.800 24.680 ;
        RECT 14.370 23.800 14.690 24.060 ;
        RECT 31.390 24.000 31.710 24.060 ;
        RECT 32.785 24.000 33.075 24.045 ;
        RECT 31.390 23.860 33.075 24.000 ;
        RECT 31.390 23.800 31.710 23.860 ;
        RECT 32.785 23.815 33.075 23.860 ;
        RECT 40.605 24.000 40.895 24.045 ;
        RECT 42.890 24.000 43.210 24.060 ;
        RECT 40.605 23.860 43.210 24.000 ;
        RECT 40.605 23.815 40.895 23.860 ;
        RECT 42.890 23.800 43.210 23.860 ;
        RECT 43.825 24.000 44.115 24.045 ;
        RECT 44.270 24.000 44.590 24.060 ;
        RECT 43.825 23.860 44.590 24.000 ;
        RECT 43.825 23.815 44.115 23.860 ;
        RECT 44.270 23.800 44.590 23.860 ;
        RECT 17.130 23.660 17.420 23.705 ;
        RECT 18.700 23.660 18.990 23.705 ;
        RECT 20.800 23.660 21.090 23.705 ;
        RECT 17.130 23.520 21.090 23.660 ;
        RECT 17.130 23.475 17.420 23.520 ;
        RECT 18.700 23.475 18.990 23.520 ;
        RECT 20.800 23.475 21.090 23.520 ;
        RECT 37.845 23.660 38.135 23.705 ;
        RECT 43.350 23.660 43.670 23.720 ;
        RECT 37.845 23.520 43.670 23.660 ;
        RECT 37.845 23.475 38.135 23.520 ;
        RECT 43.350 23.460 43.670 23.520 ;
        RECT 16.695 23.320 16.985 23.365 ;
        RECT 19.215 23.320 19.505 23.365 ;
        RECT 20.405 23.320 20.695 23.365 ;
        RECT 16.695 23.180 20.695 23.320 ;
        RECT 16.695 23.135 16.985 23.180 ;
        RECT 19.215 23.135 19.505 23.180 ;
        RECT 20.405 23.135 20.695 23.180 ;
        RECT 21.270 23.120 21.590 23.380 ;
        RECT 46.570 23.320 46.890 23.380 ;
        RECT 37.000 23.180 46.890 23.320 ;
        RECT 26.345 22.980 26.635 23.025 ;
        RECT 30.930 22.980 31.250 23.040 ;
        RECT 37.000 23.025 37.140 23.180 ;
        RECT 46.570 23.120 46.890 23.180 ;
        RECT 26.345 22.840 31.250 22.980 ;
        RECT 26.345 22.795 26.635 22.840 ;
        RECT 30.930 22.780 31.250 22.840 ;
        RECT 36.925 22.795 37.215 23.025 ;
        RECT 38.290 22.780 38.610 23.040 ;
        RECT 39.670 22.780 39.990 23.040 ;
        RECT 41.050 22.780 41.370 23.040 ;
        RECT 42.445 22.795 42.735 23.025 ;
        RECT 43.365 22.980 43.655 23.025 ;
        RECT 43.810 22.980 44.130 23.040 ;
        RECT 43.365 22.840 44.130 22.980 ;
        RECT 43.365 22.795 43.655 22.840 ;
        RECT 17.130 22.640 17.450 22.700 ;
        RECT 19.950 22.640 20.240 22.685 ;
        RECT 42.520 22.640 42.660 22.795 ;
        RECT 43.810 22.780 44.130 22.840 ;
        RECT 44.730 22.780 45.050 23.040 ;
        RECT 46.110 22.780 46.430 23.040 ;
        RECT 47.030 22.780 47.350 23.040 ;
        RECT 44.820 22.640 44.960 22.780 ;
        RECT 17.130 22.500 20.240 22.640 ;
        RECT 17.130 22.440 17.450 22.500 ;
        RECT 19.950 22.455 20.240 22.500 ;
        RECT 39.300 22.500 44.960 22.640 ;
        RECT 39.300 22.345 39.440 22.500 ;
        RECT 39.225 22.115 39.515 22.345 ;
        RECT 41.985 22.300 42.275 22.345 ;
        RECT 42.430 22.300 42.750 22.360 ;
        RECT 41.985 22.160 42.750 22.300 ;
        RECT 41.985 22.115 42.275 22.160 ;
        RECT 42.430 22.100 42.750 22.160 ;
        RECT 42.890 22.100 43.210 22.360 ;
        RECT 12.920 21.480 48.800 21.960 ;
        RECT 17.130 21.080 17.450 21.340 ;
        RECT 18.970 21.080 19.290 21.340 ;
        RECT 19.430 21.080 19.750 21.340 ;
        RECT 21.730 21.280 22.050 21.340 ;
        RECT 24.030 21.280 24.350 21.340 ;
        RECT 26.345 21.280 26.635 21.325 ;
        RECT 21.730 21.140 26.635 21.280 ;
        RECT 21.730 21.080 22.050 21.140 ;
        RECT 24.030 21.080 24.350 21.140 ;
        RECT 26.345 21.095 26.635 21.140 ;
        RECT 30.470 21.080 30.790 21.340 ;
        RECT 35.990 21.080 36.310 21.340 ;
        RECT 45.650 21.280 45.970 21.340 ;
        RECT 46.125 21.280 46.415 21.325 ;
        RECT 45.650 21.140 46.415 21.280 ;
        RECT 45.650 21.080 45.970 21.140 ;
        RECT 46.125 21.095 46.415 21.140 ;
        RECT 14.370 20.600 14.690 20.660 ;
        RECT 15.765 20.600 16.055 20.645 ;
        RECT 14.370 20.460 16.055 20.600 ;
        RECT 30.560 20.600 30.700 21.080 ;
        RECT 31.390 20.940 31.710 21.000 ;
        RECT 31.390 20.800 33.460 20.940 ;
        RECT 31.390 20.740 31.710 20.800 ;
        RECT 33.320 20.645 33.460 20.800 ;
        RECT 31.910 20.600 32.200 20.645 ;
        RECT 30.560 20.460 32.200 20.600 ;
        RECT 14.370 20.400 14.690 20.460 ;
        RECT 15.765 20.415 16.055 20.460 ;
        RECT 31.910 20.415 32.200 20.460 ;
        RECT 33.245 20.415 33.535 20.645 ;
        RECT 35.545 20.600 35.835 20.645 ;
        RECT 39.225 20.600 39.515 20.645 ;
        RECT 35.545 20.460 39.515 20.600 ;
        RECT 35.545 20.415 35.835 20.460 ;
        RECT 39.225 20.415 39.515 20.460 ;
        RECT 42.890 20.600 43.210 20.660 ;
        RECT 45.205 20.600 45.495 20.645 ;
        RECT 42.890 20.460 45.495 20.600 ;
        RECT 42.890 20.400 43.210 20.460 ;
        RECT 45.205 20.415 45.495 20.460 ;
        RECT 20.365 20.260 20.655 20.305 ;
        RECT 25.870 20.260 26.190 20.320 ;
        RECT 20.365 20.120 26.190 20.260 ;
        RECT 20.365 20.075 20.655 20.120 ;
        RECT 25.870 20.060 26.190 20.120 ;
        RECT 28.655 20.260 28.945 20.305 ;
        RECT 31.175 20.260 31.465 20.305 ;
        RECT 32.365 20.260 32.655 20.305 ;
        RECT 28.655 20.120 32.655 20.260 ;
        RECT 28.655 20.075 28.945 20.120 ;
        RECT 31.175 20.075 31.465 20.120 ;
        RECT 32.365 20.075 32.655 20.120 ;
        RECT 36.910 20.060 37.230 20.320 ;
        RECT 37.370 20.260 37.690 20.320 ;
        RECT 41.985 20.260 42.275 20.305 ;
        RECT 37.370 20.120 42.275 20.260 ;
        RECT 37.370 20.060 37.690 20.120 ;
        RECT 41.985 20.075 42.275 20.120 ;
        RECT 42.430 20.260 42.750 20.320 ;
        RECT 43.825 20.260 44.115 20.305 ;
        RECT 42.430 20.120 44.115 20.260 ;
        RECT 42.430 20.060 42.750 20.120 ;
        RECT 43.825 20.075 44.115 20.120 ;
        RECT 44.285 20.260 44.575 20.305 ;
        RECT 47.030 20.260 47.350 20.320 ;
        RECT 44.285 20.120 47.350 20.260 ;
        RECT 44.285 20.075 44.575 20.120 ;
        RECT 47.030 20.060 47.350 20.120 ;
        RECT 11.610 19.920 11.930 19.980 ;
        RECT 14.845 19.920 15.135 19.965 ;
        RECT 11.610 19.780 15.135 19.920 ;
        RECT 11.610 19.720 11.930 19.780 ;
        RECT 14.845 19.735 15.135 19.780 ;
        RECT 29.090 19.920 29.380 19.965 ;
        RECT 30.660 19.920 30.950 19.965 ;
        RECT 32.760 19.920 33.050 19.965 ;
        RECT 29.090 19.780 33.050 19.920 ;
        RECT 29.090 19.735 29.380 19.780 ;
        RECT 30.660 19.735 30.950 19.780 ;
        RECT 32.760 19.735 33.050 19.780 ;
        RECT 31.390 19.580 31.710 19.640 ;
        RECT 33.705 19.580 33.995 19.625 ;
        RECT 31.390 19.440 33.995 19.580 ;
        RECT 31.390 19.380 31.710 19.440 ;
        RECT 33.705 19.395 33.995 19.440 ;
        RECT 12.920 18.760 48.800 19.240 ;
        RECT 34.150 18.560 34.470 18.620 ;
        RECT 28.260 18.420 34.470 18.560 ;
        RECT 24.030 17.340 24.350 17.600 ;
        RECT 28.260 17.585 28.400 18.420 ;
        RECT 34.150 18.360 34.470 18.420 ;
        RECT 41.985 18.560 42.275 18.605 ;
        RECT 43.810 18.560 44.130 18.620 ;
        RECT 41.985 18.420 44.130 18.560 ;
        RECT 41.985 18.375 42.275 18.420 ;
        RECT 43.810 18.360 44.130 18.420 ;
        RECT 46.110 18.560 46.430 18.620 ;
        RECT 46.585 18.560 46.875 18.605 ;
        RECT 46.110 18.420 46.875 18.560 ;
        RECT 46.110 18.360 46.430 18.420 ;
        RECT 46.585 18.375 46.875 18.420 ;
        RECT 29.130 18.220 29.420 18.265 ;
        RECT 31.230 18.220 31.520 18.265 ;
        RECT 32.800 18.220 33.090 18.265 ;
        RECT 29.130 18.080 33.090 18.220 ;
        RECT 29.130 18.035 29.420 18.080 ;
        RECT 31.230 18.035 31.520 18.080 ;
        RECT 32.800 18.035 33.090 18.080 ;
        RECT 35.545 18.220 35.835 18.265 ;
        RECT 37.370 18.220 37.690 18.280 ;
        RECT 35.545 18.080 37.690 18.220 ;
        RECT 35.545 18.035 35.835 18.080 ;
        RECT 37.370 18.020 37.690 18.080 ;
        RECT 43.350 18.220 43.670 18.280 ;
        RECT 45.665 18.220 45.955 18.265 ;
        RECT 43.350 18.080 45.955 18.220 ;
        RECT 43.350 18.020 43.670 18.080 ;
        RECT 45.665 18.035 45.955 18.080 ;
        RECT 29.525 17.880 29.815 17.925 ;
        RECT 30.715 17.880 31.005 17.925 ;
        RECT 33.235 17.880 33.525 17.925 ;
        RECT 29.525 17.740 33.525 17.880 ;
        RECT 29.525 17.695 29.815 17.740 ;
        RECT 30.715 17.695 31.005 17.740 ;
        RECT 33.235 17.695 33.525 17.740 ;
        RECT 42.430 17.880 42.750 17.940 ;
        RECT 44.285 17.880 44.575 17.925 ;
        RECT 42.430 17.740 44.575 17.880 ;
        RECT 42.430 17.680 42.750 17.740 ;
        RECT 44.285 17.695 44.575 17.740 ;
        RECT 28.185 17.355 28.475 17.585 ;
        RECT 28.645 17.540 28.935 17.585 ;
        RECT 29.090 17.540 29.410 17.600 ;
        RECT 28.645 17.400 29.410 17.540 ;
        RECT 28.645 17.355 28.935 17.400 ;
        RECT 29.090 17.340 29.410 17.400 ;
        RECT 37.370 17.340 37.690 17.600 ;
        RECT 40.130 17.340 40.450 17.600 ;
        RECT 42.890 17.340 43.210 17.600 ;
        RECT 29.980 17.200 30.270 17.245 ;
        RECT 31.390 17.200 31.710 17.260 ;
        RECT 29.980 17.060 31.710 17.200 ;
        RECT 29.980 17.015 30.270 17.060 ;
        RECT 31.390 17.000 31.710 17.060 ;
        RECT 33.780 17.060 36.680 17.200 ;
        RECT 33.780 16.920 33.920 17.060 ;
        RECT 24.965 16.860 25.255 16.905 ;
        RECT 26.790 16.860 27.110 16.920 ;
        RECT 24.965 16.720 27.110 16.860 ;
        RECT 24.965 16.675 25.255 16.720 ;
        RECT 26.790 16.660 27.110 16.720 ;
        RECT 27.265 16.860 27.555 16.905 ;
        RECT 29.550 16.860 29.870 16.920 ;
        RECT 27.265 16.720 29.870 16.860 ;
        RECT 27.265 16.675 27.555 16.720 ;
        RECT 29.550 16.660 29.870 16.720 ;
        RECT 33.690 16.660 34.010 16.920 ;
        RECT 36.540 16.905 36.680 17.060 ;
        RECT 36.465 16.675 36.755 16.905 ;
        RECT 39.670 16.860 39.990 16.920 ;
        RECT 41.065 16.860 41.355 16.905 ;
        RECT 39.670 16.720 41.355 16.860 ;
        RECT 39.670 16.660 39.990 16.720 ;
        RECT 41.065 16.675 41.355 16.720 ;
        RECT 12.920 16.040 48.800 16.520 ;
      LAYER met2 ;
        RECT 72.300 219.400 72.580 223.400 ;
        RECT 32.180 211.835 33.720 212.205 ;
        RECT 72.370 211.670 72.510 219.400 ;
        RECT 72.310 211.350 72.570 211.670 ;
        RECT 73.690 210.670 73.950 210.990 ;
        RECT 28.880 209.115 30.420 209.485 ;
        RECT 32.180 206.395 33.720 206.765 ;
        RECT 8.360 204.015 8.640 204.385 ;
        RECT 8.430 146.390 8.570 204.015 ;
        RECT 28.880 203.675 30.420 204.045 ;
        RECT 32.180 200.955 33.720 201.325 ;
        RECT 54.830 199.790 55.090 200.110 ;
        RECT 67.250 199.790 67.510 200.110 ;
        RECT 68.170 199.790 68.430 200.110 ;
        RECT 28.880 198.235 30.420 198.605 ;
        RECT 32.180 195.515 33.720 195.885 ;
        RECT 54.890 195.350 55.030 199.790 ;
        RECT 66.790 199.450 67.050 199.770 ;
        RECT 62.190 199.110 62.450 199.430 ;
        RECT 54.830 195.030 55.090 195.350 ;
        RECT 62.250 194.670 62.390 199.110 ;
        RECT 63.110 198.770 63.370 199.090 ;
        RECT 62.650 196.050 62.910 196.370 ;
        RECT 62.710 194.670 62.850 196.050 ;
        RECT 60.350 194.350 60.610 194.670 ;
        RECT 62.190 194.350 62.450 194.670 ;
        RECT 62.650 194.350 62.910 194.670 ;
        RECT 33.670 194.010 33.930 194.330 ;
        RECT 34.130 194.010 34.390 194.330 ;
        RECT 37.810 194.010 38.070 194.330 ;
        RECT 30.910 193.670 31.170 193.990 ;
        RECT 28.880 192.795 30.420 193.165 ;
        RECT 25.850 191.970 26.110 192.290 ;
        RECT 26.310 191.970 26.570 192.290 ;
        RECT 30.970 192.030 31.110 193.670 ;
        RECT 24.010 191.630 24.270 191.950 ;
        RECT 17.570 191.290 17.830 191.610 ;
        RECT 17.630 188.550 17.770 191.290 ;
        RECT 20.330 190.950 20.590 191.270 ;
        RECT 20.390 189.910 20.530 190.950 ;
        RECT 20.790 190.610 21.050 190.930 ;
        RECT 20.850 189.910 20.990 190.610 ;
        RECT 24.070 189.990 24.210 191.630 ;
        RECT 20.330 189.590 20.590 189.910 ;
        RECT 20.790 189.590 21.050 189.910 ;
        RECT 23.610 189.850 24.210 189.990 ;
        RECT 17.570 188.230 17.830 188.550 ;
        RECT 12.050 183.470 12.310 183.790 ;
        RECT 12.110 182.625 12.250 183.470 ;
        RECT 17.630 183.450 17.770 188.230 ;
        RECT 20.330 186.490 20.590 186.510 ;
        RECT 20.850 186.490 20.990 189.590 ;
        RECT 23.610 188.890 23.750 189.850 ;
        RECT 25.910 189.230 26.050 191.970 ;
        RECT 25.850 188.910 26.110 189.230 ;
        RECT 21.710 188.570 21.970 188.890 ;
        RECT 23.550 188.570 23.810 188.890 ;
        RECT 21.770 186.850 21.910 188.570 ;
        RECT 21.710 186.530 21.970 186.850 ;
        RECT 20.330 186.350 20.990 186.490 ;
        RECT 20.330 186.190 20.590 186.350 ;
        RECT 19.870 186.080 20.130 186.170 ;
        RECT 19.470 185.940 20.130 186.080 ;
        RECT 18.490 185.170 18.750 185.490 ;
        RECT 18.550 184.130 18.690 185.170 ;
        RECT 18.490 183.810 18.750 184.130 ;
        RECT 17.570 183.130 17.830 183.450 ;
        RECT 12.040 182.255 12.320 182.625 ;
        RECT 17.630 180.730 17.770 183.130 ;
        RECT 17.570 180.410 17.830 180.730 ;
        RECT 18.490 180.070 18.750 180.390 ;
        RECT 18.550 179.030 18.690 180.070 ;
        RECT 19.470 179.030 19.610 185.940 ;
        RECT 19.870 185.850 20.130 185.940 ;
        RECT 19.870 180.410 20.130 180.730 ;
        RECT 19.930 179.030 20.070 180.410 ;
        RECT 18.490 178.710 18.750 179.030 ;
        RECT 19.410 178.710 19.670 179.030 ;
        RECT 19.870 178.710 20.130 179.030 ;
        RECT 17.570 178.030 17.830 178.350 ;
        RECT 17.630 176.310 17.770 178.030 ;
        RECT 18.950 177.010 19.210 177.330 ;
        RECT 17.570 175.990 17.830 176.310 ;
        RECT 19.010 174.610 19.150 177.010 ;
        RECT 18.950 174.290 19.210 174.610 ;
        RECT 19.010 172.910 19.150 174.290 ;
        RECT 19.470 173.250 19.610 178.710 ;
        RECT 19.410 172.930 19.670 173.250 ;
        RECT 18.950 172.590 19.210 172.910 ;
        RECT 12.050 169.530 12.310 169.850 ;
        RECT 12.110 169.025 12.250 169.530 ;
        RECT 12.040 168.655 12.320 169.025 ;
        RECT 17.570 168.850 17.830 169.170 ;
        RECT 17.630 164.070 17.770 168.850 ;
        RECT 19.010 168.150 19.150 172.590 ;
        RECT 19.470 169.850 19.610 172.930 ;
        RECT 19.410 169.530 19.670 169.850 ;
        RECT 18.950 167.830 19.210 168.150 ;
        RECT 19.930 167.470 20.070 178.710 ;
        RECT 20.390 178.350 20.530 186.190 ;
        RECT 23.610 186.170 23.750 188.570 ;
        RECT 25.910 188.210 26.050 188.910 ;
        RECT 25.850 187.890 26.110 188.210 ;
        RECT 25.910 187.190 26.050 187.890 ;
        RECT 25.850 186.870 26.110 187.190 ;
        RECT 26.370 186.850 26.510 191.970 ;
        RECT 30.050 191.950 31.110 192.030 ;
        RECT 33.730 192.030 33.870 194.010 ;
        RECT 34.190 192.630 34.330 194.010 ;
        RECT 35.050 193.330 35.310 193.650 ;
        RECT 35.510 193.330 35.770 193.650 ;
        RECT 34.130 192.310 34.390 192.630 ;
        RECT 29.990 191.890 31.110 191.950 ;
        RECT 29.990 191.630 30.250 191.890 ;
        RECT 31.370 191.630 31.630 191.950 ;
        RECT 33.730 191.890 34.330 192.030 ;
        RECT 30.910 190.950 31.170 191.270 ;
        RECT 30.970 188.890 31.110 190.950 ;
        RECT 26.770 188.570 27.030 188.890 ;
        RECT 30.910 188.570 31.170 188.890 ;
        RECT 26.830 186.850 26.970 188.570 ;
        RECT 30.910 187.890 31.170 188.210 ;
        RECT 28.880 187.355 30.420 187.725 ;
        RECT 30.450 186.870 30.710 187.190 ;
        RECT 26.310 186.530 26.570 186.850 ;
        RECT 26.770 186.530 27.030 186.850 ;
        RECT 30.510 186.705 30.650 186.870 ;
        RECT 21.250 185.850 21.510 186.170 ;
        RECT 23.550 185.850 23.810 186.170 ;
        RECT 21.310 178.350 21.450 185.850 ;
        RECT 25.850 185.510 26.110 185.830 ;
        RECT 25.910 184.470 26.050 185.510 ;
        RECT 25.850 184.150 26.110 184.470 ;
        RECT 26.830 183.790 26.970 186.530 ;
        RECT 30.440 186.335 30.720 186.705 ;
        RECT 24.470 183.470 24.730 183.790 ;
        RECT 26.770 183.470 27.030 183.790 ;
        RECT 24.010 182.450 24.270 182.770 ;
        RECT 24.070 181.070 24.210 182.450 ;
        RECT 24.530 181.750 24.670 183.470 ;
        RECT 24.930 182.450 25.190 182.770 ;
        RECT 24.470 181.430 24.730 181.750 ;
        RECT 24.010 180.750 24.270 181.070 ;
        RECT 24.990 180.730 25.130 182.450 ;
        RECT 22.170 180.410 22.430 180.730 ;
        RECT 24.930 180.410 25.190 180.730 ;
        RECT 21.710 178.370 21.970 178.690 ;
        RECT 20.330 178.030 20.590 178.350 ;
        RECT 21.250 178.030 21.510 178.350 ;
        RECT 20.390 170.190 20.530 178.030 ;
        RECT 20.790 171.570 21.050 171.890 ;
        RECT 20.850 170.190 20.990 171.570 ;
        RECT 21.310 170.530 21.450 178.030 ;
        RECT 21.770 175.290 21.910 178.370 ;
        RECT 22.230 177.670 22.370 180.410 ;
        RECT 24.010 179.730 24.270 180.050 ;
        RECT 24.070 178.690 24.210 179.730 ;
        RECT 24.010 178.370 24.270 178.690 ;
        RECT 22.170 177.350 22.430 177.670 ;
        RECT 24.070 176.310 24.210 178.370 ;
        RECT 24.990 178.010 25.130 180.410 ;
        RECT 26.830 178.690 26.970 183.470 ;
        RECT 30.510 183.190 30.650 186.335 ;
        RECT 30.970 186.170 31.110 187.890 ;
        RECT 31.430 187.190 31.570 191.630 ;
        RECT 33.730 191.270 33.870 191.890 ;
        RECT 33.670 190.950 33.930 191.270 ;
        RECT 32.290 190.840 32.550 190.930 ;
        RECT 31.890 190.700 32.550 190.840 ;
        RECT 31.890 189.570 32.030 190.700 ;
        RECT 32.290 190.610 32.550 190.700 ;
        RECT 32.180 190.075 33.720 190.445 ;
        RECT 34.190 189.910 34.330 191.890 ;
        RECT 32.750 189.820 33.010 189.910 ;
        RECT 32.350 189.680 33.010 189.820 ;
        RECT 31.830 189.250 32.090 189.570 ;
        RECT 32.350 188.210 32.490 189.680 ;
        RECT 32.750 189.590 33.010 189.680 ;
        RECT 34.130 189.590 34.390 189.910 ;
        RECT 32.290 187.890 32.550 188.210 ;
        RECT 34.590 187.890 34.850 188.210 ;
        RECT 31.370 186.870 31.630 187.190 ;
        RECT 32.350 186.170 32.490 187.890 ;
        RECT 33.200 186.335 33.480 186.705 ;
        RECT 33.670 186.530 33.930 186.850 ;
        RECT 33.270 186.170 33.410 186.335 ;
        RECT 33.730 186.170 33.870 186.530 ;
        RECT 30.910 185.850 31.170 186.170 ;
        RECT 32.290 185.850 32.550 186.170 ;
        RECT 33.210 185.850 33.470 186.170 ;
        RECT 33.670 185.850 33.930 186.170 ;
        RECT 34.650 185.490 34.790 187.890 ;
        RECT 35.110 187.190 35.250 193.330 ;
        RECT 35.570 191.610 35.710 193.330 ;
        RECT 35.510 191.290 35.770 191.610 ;
        RECT 35.050 186.870 35.310 187.190 ;
        RECT 37.870 186.510 38.010 194.010 ;
        RECT 51.150 193.330 51.410 193.650 ;
        RECT 50.230 192.310 50.490 192.630 ;
        RECT 49.310 191.290 49.570 191.610 ;
        RECT 42.870 190.950 43.130 191.270 ;
        RECT 39.650 190.610 39.910 190.930 ;
        RECT 41.030 190.610 41.290 190.930 ;
        RECT 39.710 186.850 39.850 190.610 ;
        RECT 41.090 189.570 41.230 190.610 ;
        RECT 42.930 189.910 43.070 190.950 ;
        RECT 42.870 189.590 43.130 189.910 ;
        RECT 41.030 189.250 41.290 189.570 ;
        RECT 47.470 189.250 47.730 189.570 ;
        RECT 39.650 186.530 39.910 186.850 ;
        RECT 37.810 186.190 38.070 186.510 ;
        RECT 39.710 186.170 39.850 186.530 ;
        RECT 37.350 185.850 37.610 186.170 ;
        RECT 39.650 185.850 39.910 186.170 ;
        RECT 37.410 185.490 37.550 185.850 ;
        RECT 34.590 185.170 34.850 185.490 ;
        RECT 37.350 185.170 37.610 185.490 ;
        RECT 32.180 184.635 33.720 185.005 ;
        RECT 30.510 183.050 31.110 183.190 ;
        RECT 28.880 181.915 30.420 182.285 ;
        RECT 28.150 180.410 28.410 180.730 ;
        RECT 30.970 180.470 31.110 183.050 ;
        RECT 34.650 181.750 34.790 185.170 ;
        RECT 34.590 181.430 34.850 181.750 ;
        RECT 36.430 181.090 36.690 181.410 ;
        RECT 36.890 181.090 37.150 181.410 ;
        RECT 28.210 178.690 28.350 180.410 ;
        RECT 30.510 180.330 31.110 180.470 ;
        RECT 26.770 178.370 27.030 178.690 ;
        RECT 28.150 178.370 28.410 178.690 ;
        RECT 25.850 178.030 26.110 178.350 ;
        RECT 24.930 177.690 25.190 178.010 ;
        RECT 24.010 175.990 24.270 176.310 ;
        RECT 24.070 175.290 24.210 175.990 ;
        RECT 25.910 175.630 26.050 178.030 ;
        RECT 26.770 175.990 27.030 176.310 ;
        RECT 25.850 175.310 26.110 175.630 ;
        RECT 21.710 174.970 21.970 175.290 ;
        RECT 24.010 174.970 24.270 175.290 ;
        RECT 21.770 172.570 21.910 174.970 ;
        RECT 23.550 172.930 23.810 173.250 ;
        RECT 21.710 172.250 21.970 172.570 ;
        RECT 21.250 170.210 21.510 170.530 ;
        RECT 20.330 169.870 20.590 170.190 ;
        RECT 20.790 169.870 21.050 170.190 ;
        RECT 21.770 169.510 21.910 172.250 ;
        RECT 23.610 170.190 23.750 172.930 ;
        RECT 26.830 172.910 26.970 175.990 ;
        RECT 28.210 175.630 28.350 178.370 ;
        RECT 30.510 178.350 30.650 180.330 ;
        RECT 31.830 180.070 32.090 180.390 ;
        RECT 30.910 179.730 31.170 180.050 ;
        RECT 30.970 178.350 31.110 179.730 ;
        RECT 30.450 178.030 30.710 178.350 ;
        RECT 30.910 178.030 31.170 178.350 ;
        RECT 31.370 178.030 31.630 178.350 ;
        RECT 28.880 176.475 30.420 176.845 ;
        RECT 28.150 175.310 28.410 175.630 ;
        RECT 27.230 174.970 27.490 175.290 ;
        RECT 26.770 172.590 27.030 172.910 ;
        RECT 27.290 172.570 27.430 174.970 ;
        RECT 28.210 172.910 28.350 175.310 ;
        RECT 30.970 175.290 31.110 178.030 ;
        RECT 30.910 174.970 31.170 175.290 ;
        RECT 31.430 173.500 31.570 178.030 ;
        RECT 30.970 173.360 31.570 173.500 ;
        RECT 28.150 172.590 28.410 172.910 ;
        RECT 30.970 172.570 31.110 173.360 ;
        RECT 31.370 172.590 31.630 172.910 ;
        RECT 27.230 172.250 27.490 172.570 ;
        RECT 30.910 172.250 31.170 172.570 ;
        RECT 23.550 169.870 23.810 170.190 ;
        RECT 26.770 169.530 27.030 169.850 ;
        RECT 21.710 169.190 21.970 169.510 ;
        RECT 19.870 167.150 20.130 167.470 ;
        RECT 19.930 166.870 20.070 167.150 ;
        RECT 19.470 166.730 20.070 166.870 ;
        RECT 19.470 164.410 19.610 166.730 ;
        RECT 21.770 165.430 21.910 169.190 ;
        RECT 22.170 168.850 22.430 169.170 ;
        RECT 22.230 167.380 22.370 168.850 ;
        RECT 22.630 167.380 22.890 167.470 ;
        RECT 22.230 167.240 22.890 167.380 ;
        RECT 22.630 167.150 22.890 167.240 ;
        RECT 21.710 165.110 21.970 165.430 ;
        RECT 19.410 164.090 19.670 164.410 ;
        RECT 17.570 163.750 17.830 164.070 ;
        RECT 15.730 157.970 15.990 158.290 ;
        RECT 15.790 157.270 15.930 157.970 ;
        RECT 15.730 156.950 15.990 157.270 ;
        RECT 16.650 156.610 16.910 156.930 ;
        RECT 12.050 156.270 12.310 156.590 ;
        RECT 12.110 155.425 12.250 156.270 ;
        RECT 12.040 155.055 12.320 155.425 ;
        RECT 16.710 154.550 16.850 156.610 ;
        RECT 19.470 156.590 19.610 164.090 ;
        RECT 26.830 162.710 26.970 169.530 ;
        RECT 26.770 162.390 27.030 162.710 ;
        RECT 26.830 162.030 26.970 162.390 ;
        RECT 26.770 161.710 27.030 162.030 ;
        RECT 27.290 161.690 27.430 172.250 ;
        RECT 28.880 171.035 30.420 171.405 ;
        RECT 28.610 170.550 28.870 170.870 ;
        RECT 28.150 169.530 28.410 169.850 ;
        RECT 28.210 168.150 28.350 169.530 ;
        RECT 28.150 167.830 28.410 168.150 ;
        RECT 27.690 167.150 27.950 167.470 ;
        RECT 28.150 167.380 28.410 167.470 ;
        RECT 28.670 167.380 28.810 170.550 ;
        RECT 29.990 168.850 30.250 169.170 ;
        RECT 30.050 167.470 30.190 168.850 ;
        RECT 28.150 167.240 28.810 167.380 ;
        RECT 28.150 167.150 28.410 167.240 ;
        RECT 29.990 167.150 30.250 167.470 ;
        RECT 27.750 165.430 27.890 167.150 ;
        RECT 27.690 165.110 27.950 165.430 ;
        RECT 27.750 164.410 27.890 165.110 ;
        RECT 28.210 165.000 28.350 167.150 ;
        RECT 28.880 165.595 30.420 165.965 ;
        RECT 28.610 165.000 28.870 165.090 ;
        RECT 28.210 164.860 28.870 165.000 ;
        RECT 28.610 164.770 28.870 164.860 ;
        RECT 27.690 164.090 27.950 164.410 ;
        RECT 28.670 164.070 28.810 164.770 ;
        RECT 28.610 163.750 28.870 164.070 ;
        RECT 29.990 163.410 30.250 163.730 ;
        RECT 30.050 162.030 30.190 163.410 ;
        RECT 30.970 162.710 31.110 172.250 ;
        RECT 31.430 169.850 31.570 172.590 ;
        RECT 31.890 172.425 32.030 180.070 ;
        RECT 35.970 179.730 36.230 180.050 ;
        RECT 32.180 179.195 33.720 179.565 ;
        RECT 33.210 177.690 33.470 178.010 ;
        RECT 33.270 175.290 33.410 177.690 ;
        RECT 33.670 177.010 33.930 177.330 ;
        RECT 33.730 175.290 33.870 177.010 ;
        RECT 36.030 175.290 36.170 179.730 ;
        RECT 36.490 175.290 36.630 181.090 ;
        RECT 36.950 180.730 37.090 181.090 ;
        RECT 39.710 181.070 39.850 185.850 ;
        RECT 41.090 182.770 41.230 189.250 ;
        RECT 47.010 188.910 47.270 189.230 ;
        RECT 41.950 188.570 42.210 188.890 ;
        RECT 46.550 188.570 46.810 188.890 ;
        RECT 42.010 185.490 42.150 188.570 ;
        RECT 43.330 185.850 43.590 186.170 ;
        RECT 41.950 185.170 42.210 185.490 ;
        RECT 42.010 184.550 42.150 185.170 ;
        RECT 42.010 184.470 42.610 184.550 ;
        RECT 42.010 184.410 42.670 184.470 ;
        RECT 42.410 184.150 42.670 184.410 ;
        RECT 42.870 183.470 43.130 183.790 ;
        RECT 41.490 183.130 41.750 183.450 ;
        RECT 40.110 182.450 40.370 182.770 ;
        RECT 41.030 182.450 41.290 182.770 ;
        RECT 40.170 181.070 40.310 182.450 ;
        RECT 41.030 181.090 41.290 181.410 ;
        RECT 39.650 180.750 39.910 181.070 ;
        RECT 40.110 180.750 40.370 181.070 ;
        RECT 36.890 180.410 37.150 180.730 ;
        RECT 37.810 180.640 38.070 180.730 ;
        RECT 37.810 180.500 39.390 180.640 ;
        RECT 37.810 180.410 38.070 180.500 ;
        RECT 39.250 180.470 39.390 180.500 ;
        RECT 40.170 180.470 40.310 180.750 ;
        RECT 39.250 180.330 40.310 180.470 ;
        RECT 40.570 180.410 40.830 180.730 ;
        RECT 33.210 174.970 33.470 175.290 ;
        RECT 33.670 174.970 33.930 175.290 ;
        RECT 35.970 174.970 36.230 175.290 ;
        RECT 36.430 174.970 36.690 175.290 ;
        RECT 35.970 174.290 36.230 174.610 ;
        RECT 36.890 174.290 37.150 174.610 ;
        RECT 37.350 174.290 37.610 174.610 ;
        RECT 32.180 173.755 33.720 174.125 ;
        RECT 31.820 172.055 32.100 172.425 ;
        RECT 31.830 171.570 32.090 171.890 ;
        RECT 31.890 169.850 32.030 171.570 ;
        RECT 33.210 170.550 33.470 170.870 ;
        RECT 33.270 169.850 33.410 170.550 ;
        RECT 36.030 170.190 36.170 174.290 ;
        RECT 36.950 173.250 37.090 174.290 ;
        RECT 36.890 172.930 37.150 173.250 ;
        RECT 37.410 172.910 37.550 174.290 ;
        RECT 40.630 173.500 40.770 180.410 ;
        RECT 39.710 173.360 40.770 173.500 ;
        RECT 37.350 172.590 37.610 172.910 ;
        RECT 37.810 172.590 38.070 172.910 ;
        RECT 37.870 172.310 38.010 172.590 ;
        RECT 37.410 172.170 38.010 172.310 ;
        RECT 35.970 169.870 36.230 170.190 ;
        RECT 36.430 169.870 36.690 170.190 ;
        RECT 31.370 169.530 31.630 169.850 ;
        RECT 31.830 169.530 32.090 169.850 ;
        RECT 33.210 169.760 33.470 169.850 ;
        RECT 33.210 169.620 34.330 169.760 ;
        RECT 33.210 169.530 33.470 169.620 ;
        RECT 32.180 168.315 33.720 168.685 ;
        RECT 34.190 168.150 34.330 169.620 ;
        RECT 34.590 169.530 34.850 169.850 ;
        RECT 34.130 167.830 34.390 168.150 ;
        RECT 34.650 165.430 34.790 169.530 ;
        RECT 35.510 169.190 35.770 169.510 ;
        RECT 35.570 168.150 35.710 169.190 ;
        RECT 35.510 167.830 35.770 168.150 ;
        RECT 36.490 167.810 36.630 169.870 ;
        RECT 36.890 169.760 37.150 169.850 ;
        RECT 37.410 169.760 37.550 172.170 ;
        RECT 37.810 171.570 38.070 171.890 ;
        RECT 36.890 169.620 37.550 169.760 ;
        RECT 36.890 169.530 37.150 169.620 ;
        RECT 36.430 167.490 36.690 167.810 ;
        RECT 36.950 166.870 37.090 169.530 ;
        RECT 37.350 168.850 37.610 169.170 ;
        RECT 37.410 167.470 37.550 168.850 ;
        RECT 37.870 167.470 38.010 171.570 ;
        RECT 39.190 168.850 39.450 169.170 ;
        RECT 37.350 167.150 37.610 167.470 ;
        RECT 37.810 167.150 38.070 167.470 ;
        RECT 36.950 166.730 37.550 166.870 ;
        RECT 34.590 165.110 34.850 165.430 ;
        RECT 36.890 164.090 37.150 164.410 ;
        RECT 32.180 162.875 33.720 163.245 ;
        RECT 30.910 162.390 31.170 162.710 ;
        RECT 29.990 161.710 30.250 162.030 ;
        RECT 27.230 161.370 27.490 161.690 ;
        RECT 27.290 156.590 27.430 161.370 ;
        RECT 28.880 160.155 30.420 160.525 ;
        RECT 30.970 157.270 31.110 162.390 ;
        RECT 35.970 159.330 36.230 159.650 ;
        RECT 32.180 157.435 33.720 157.805 ;
        RECT 30.910 156.950 31.170 157.270 ;
        RECT 35.510 156.610 35.770 156.930 ;
        RECT 19.410 156.270 19.670 156.590 ;
        RECT 19.870 156.270 20.130 156.590 ;
        RECT 27.230 156.270 27.490 156.590 ;
        RECT 31.830 156.270 32.090 156.590 ;
        RECT 19.930 154.550 20.070 156.270 ;
        RECT 28.150 155.250 28.410 155.570 ;
        RECT 31.370 155.250 31.630 155.570 ;
        RECT 16.650 154.230 16.910 154.550 ;
        RECT 19.870 154.230 20.130 154.550 ;
        RECT 20.790 154.230 21.050 154.550 ;
        RECT 15.270 152.870 15.530 153.190 ;
        RECT 15.330 151.345 15.470 152.870 ;
        RECT 15.260 150.975 15.540 151.345 ;
        RECT 20.850 151.150 20.990 154.230 ;
        RECT 24.010 153.550 24.270 153.870 ;
        RECT 24.470 153.550 24.730 153.870 ;
        RECT 22.170 153.210 22.430 153.530 ;
        RECT 21.250 152.870 21.510 153.190 ;
        RECT 20.790 150.830 21.050 151.150 ;
        RECT 17.110 149.810 17.370 150.130 ;
        RECT 15.730 147.770 15.990 148.090 ;
        RECT 8.370 146.070 8.630 146.390 ;
        RECT 15.790 145.710 15.930 147.770 ;
        RECT 17.170 145.710 17.310 149.810 ;
        RECT 18.490 147.430 18.750 147.750 ;
        RECT 15.730 145.390 15.990 145.710 ;
        RECT 17.110 145.390 17.370 145.710 ;
        RECT 18.550 143.670 18.690 147.430 ;
        RECT 20.850 143.670 20.990 150.830 ;
        RECT 21.310 150.470 21.450 152.870 ;
        RECT 22.230 151.150 22.370 153.210 ;
        RECT 22.630 152.530 22.890 152.850 ;
        RECT 23.550 152.530 23.810 152.850 ;
        RECT 22.170 150.830 22.430 151.150 ;
        RECT 21.250 150.150 21.510 150.470 ;
        RECT 18.490 143.350 18.750 143.670 ;
        RECT 20.790 143.350 21.050 143.670 ;
        RECT 20.850 138.230 20.990 143.350 ;
        RECT 21.310 142.310 21.450 150.150 ;
        RECT 22.170 149.810 22.430 150.130 ;
        RECT 22.230 145.370 22.370 149.810 ;
        RECT 22.690 145.710 22.830 152.530 ;
        RECT 23.610 151.830 23.750 152.530 ;
        RECT 23.550 151.510 23.810 151.830 ;
        RECT 23.550 150.830 23.810 151.150 ;
        RECT 23.090 150.490 23.350 150.810 ;
        RECT 23.150 148.090 23.290 150.490 ;
        RECT 23.610 148.430 23.750 150.830 ;
        RECT 24.070 149.110 24.210 153.550 ;
        RECT 24.530 153.190 24.670 153.550 ;
        RECT 28.210 153.530 28.350 155.250 ;
        RECT 28.880 154.715 30.420 155.085 ;
        RECT 25.850 153.210 26.110 153.530 ;
        RECT 28.150 153.270 28.410 153.530 ;
        RECT 28.150 153.210 28.810 153.270 ;
        RECT 24.470 152.870 24.730 153.190 ;
        RECT 24.530 150.130 24.670 152.870 ;
        RECT 24.470 149.810 24.730 150.130 ;
        RECT 25.910 149.870 26.050 153.210 ;
        RECT 27.690 152.870 27.950 153.190 ;
        RECT 28.210 153.130 28.810 153.210 ;
        RECT 26.770 152.530 27.030 152.850 ;
        RECT 26.310 149.870 26.570 150.130 ;
        RECT 25.910 149.810 26.570 149.870 ;
        RECT 24.530 149.190 24.670 149.810 ;
        RECT 25.910 149.730 26.510 149.810 ;
        RECT 24.530 149.110 25.130 149.190 ;
        RECT 24.010 148.790 24.270 149.110 ;
        RECT 24.530 149.050 25.190 149.110 ;
        RECT 24.930 148.790 25.190 149.050 ;
        RECT 24.470 148.450 24.730 148.770 ;
        RECT 23.550 148.110 23.810 148.430 ;
        RECT 23.090 147.770 23.350 148.090 ;
        RECT 22.630 145.390 22.890 145.710 ;
        RECT 22.170 145.050 22.430 145.370 ;
        RECT 21.250 141.990 21.510 142.310 ;
        RECT 20.790 137.910 21.050 138.230 ;
        RECT 20.850 136.950 20.990 137.910 ;
        RECT 14.810 136.550 15.070 136.870 ;
        RECT 20.390 136.810 20.990 136.950 ;
        RECT 21.310 136.870 21.450 141.990 ;
        RECT 22.170 139.950 22.430 140.270 ;
        RECT 22.230 137.550 22.370 139.950 ;
        RECT 22.170 137.230 22.430 137.550 ;
        RECT 14.870 134.830 15.010 136.550 ;
        RECT 20.390 136.530 20.530 136.810 ;
        RECT 21.250 136.550 21.510 136.870 ;
        RECT 17.570 136.210 17.830 136.530 ;
        RECT 19.870 136.210 20.130 136.530 ;
        RECT 20.330 136.210 20.590 136.530 ;
        RECT 17.630 134.830 17.770 136.210 ;
        RECT 19.930 135.510 20.070 136.210 ;
        RECT 22.230 135.510 22.370 137.230 ;
        RECT 22.630 136.550 22.890 136.870 ;
        RECT 19.870 135.190 20.130 135.510 ;
        RECT 22.170 135.190 22.430 135.510 ;
        RECT 14.810 134.510 15.070 134.830 ;
        RECT 17.570 134.510 17.830 134.830 ;
        RECT 22.690 133.810 22.830 136.550 ;
        RECT 23.150 135.170 23.290 147.770 ;
        RECT 24.010 145.620 24.270 145.710 ;
        RECT 24.530 145.620 24.670 148.450 ;
        RECT 25.910 148.090 26.050 149.730 ;
        RECT 26.310 148.790 26.570 149.110 ;
        RECT 26.370 148.090 26.510 148.790 ;
        RECT 25.850 147.770 26.110 148.090 ;
        RECT 26.310 147.770 26.570 148.090 ;
        RECT 26.830 145.710 26.970 152.530 ;
        RECT 27.750 151.830 27.890 152.870 ;
        RECT 27.690 151.510 27.950 151.830 ;
        RECT 27.750 148.090 27.890 151.510 ;
        RECT 28.670 151.150 28.810 153.130 ;
        RECT 28.610 150.830 28.870 151.150 ;
        RECT 28.880 149.275 30.420 149.645 ;
        RECT 31.430 148.090 31.570 155.250 ;
        RECT 31.890 152.850 32.030 156.270 ;
        RECT 31.830 152.530 32.090 152.850 ;
        RECT 34.590 152.530 34.850 152.850 ;
        RECT 31.890 149.110 32.030 152.530 ;
        RECT 32.180 151.995 33.720 152.365 ;
        RECT 34.650 151.490 34.790 152.530 ;
        RECT 35.570 151.830 35.710 156.610 ;
        RECT 35.510 151.510 35.770 151.830 ;
        RECT 34.590 151.170 34.850 151.490 ;
        RECT 32.750 149.810 33.010 150.130 ;
        RECT 31.830 148.790 32.090 149.110 ;
        RECT 32.810 148.090 32.950 149.810 ;
        RECT 33.270 149.110 34.330 149.190 ;
        RECT 33.210 149.050 34.330 149.110 ;
        RECT 33.210 148.790 33.470 149.050 ;
        RECT 34.190 148.770 34.330 149.050 ;
        RECT 34.130 148.450 34.390 148.770 ;
        RECT 34.590 148.110 34.850 148.430 ;
        RECT 27.690 147.770 27.950 148.090 ;
        RECT 28.150 147.945 28.410 148.090 ;
        RECT 28.140 147.575 28.420 147.945 ;
        RECT 31.370 147.770 31.630 148.090 ;
        RECT 31.830 147.770 32.090 148.090 ;
        RECT 32.750 147.770 33.010 148.090 ;
        RECT 31.890 145.710 32.030 147.770 ;
        RECT 32.180 146.555 33.720 146.925 ;
        RECT 34.130 145.730 34.390 146.050 ;
        RECT 24.010 145.480 24.670 145.620 ;
        RECT 24.010 145.390 24.270 145.480 ;
        RECT 26.770 145.390 27.030 145.710 ;
        RECT 31.830 145.390 32.090 145.710 ;
        RECT 23.550 145.050 23.810 145.370 ;
        RECT 23.610 136.870 23.750 145.050 ;
        RECT 24.470 144.370 24.730 144.690 ;
        RECT 32.750 144.370 33.010 144.690 ;
        RECT 24.530 141.970 24.670 144.370 ;
        RECT 28.880 143.835 30.420 144.205 ;
        RECT 32.810 142.650 32.950 144.370 ;
        RECT 34.190 143.670 34.330 145.730 ;
        RECT 34.650 145.710 34.790 148.110 ;
        RECT 35.570 148.090 35.710 151.510 ;
        RECT 36.030 150.130 36.170 159.330 ;
        RECT 36.950 157.270 37.090 164.090 ;
        RECT 37.410 161.350 37.550 166.730 ;
        RECT 39.250 164.750 39.390 168.850 ;
        RECT 39.190 164.430 39.450 164.750 ;
        RECT 39.710 162.030 39.850 173.360 ;
        RECT 40.570 172.590 40.830 172.910 ;
        RECT 40.630 169.850 40.770 172.590 ;
        RECT 40.570 169.530 40.830 169.850 ;
        RECT 40.110 169.190 40.370 169.510 ;
        RECT 40.170 167.810 40.310 169.190 ;
        RECT 40.110 167.490 40.370 167.810 ;
        RECT 40.570 164.090 40.830 164.410 ;
        RECT 39.190 161.710 39.450 162.030 ;
        RECT 39.650 161.710 39.910 162.030 ;
        RECT 38.730 161.370 38.990 161.690 ;
        RECT 37.350 161.030 37.610 161.350 ;
        RECT 38.790 158.970 38.930 161.370 ;
        RECT 38.730 158.650 38.990 158.970 ;
        RECT 39.250 158.880 39.390 161.710 ;
        RECT 40.630 161.010 40.770 164.090 ;
        RECT 40.570 160.690 40.830 161.010 ;
        RECT 41.090 159.650 41.230 181.090 ;
        RECT 41.550 180.390 41.690 183.130 ;
        RECT 42.930 182.510 43.070 183.470 ;
        RECT 43.390 183.110 43.530 185.850 ;
        RECT 43.330 182.790 43.590 183.110 ;
        RECT 42.930 182.370 43.530 182.510 ;
        RECT 41.490 180.070 41.750 180.390 ;
        RECT 41.950 179.730 42.210 180.050 ;
        RECT 42.010 176.310 42.150 179.730 ;
        RECT 41.950 175.990 42.210 176.310 ;
        RECT 42.010 174.950 42.150 175.990 ;
        RECT 41.950 174.630 42.210 174.950 ;
        RECT 42.410 174.290 42.670 174.610 ;
        RECT 42.470 172.910 42.610 174.290 ;
        RECT 42.410 172.590 42.670 172.910 ;
        RECT 42.870 171.570 43.130 171.890 ;
        RECT 41.490 169.870 41.750 170.190 ;
        RECT 41.030 159.330 41.290 159.650 ;
        RECT 39.650 158.880 39.910 158.970 ;
        RECT 39.250 158.740 39.910 158.880 ;
        RECT 39.650 158.650 39.910 158.740 ;
        RECT 36.890 156.950 37.150 157.270 ;
        RECT 36.430 153.210 36.690 153.530 ;
        RECT 36.490 150.810 36.630 153.210 ;
        RECT 36.950 151.490 37.090 156.950 ;
        RECT 38.790 156.930 38.930 158.650 ;
        RECT 38.730 156.610 38.990 156.930 ;
        RECT 39.710 156.590 39.850 158.650 ;
        RECT 39.650 156.270 39.910 156.590 ;
        RECT 37.350 155.590 37.610 155.910 ;
        RECT 37.410 153.870 37.550 155.590 ;
        RECT 40.570 155.250 40.830 155.570 ;
        RECT 37.350 153.550 37.610 153.870 ;
        RECT 36.890 151.170 37.150 151.490 ;
        RECT 36.430 150.490 36.690 150.810 ;
        RECT 35.970 149.810 36.230 150.130 ;
        RECT 35.510 147.770 35.770 148.090 ;
        RECT 36.030 147.410 36.170 149.810 ;
        RECT 37.410 147.945 37.550 153.550 ;
        RECT 40.630 153.530 40.770 155.250 ;
        RECT 41.550 154.550 41.690 169.870 ;
        RECT 42.410 167.150 42.670 167.470 ;
        RECT 42.470 165.430 42.610 167.150 ;
        RECT 42.930 167.130 43.070 171.570 ;
        RECT 43.390 167.130 43.530 182.370 ;
        RECT 44.710 179.730 44.970 180.050 ;
        RECT 44.770 179.030 44.910 179.730 ;
        RECT 44.710 178.710 44.970 179.030 ;
        RECT 44.770 169.850 44.910 178.710 ;
        RECT 46.610 175.630 46.750 188.570 ;
        RECT 47.070 185.490 47.210 188.910 ;
        RECT 47.530 185.490 47.670 189.250 ;
        RECT 47.010 185.170 47.270 185.490 ;
        RECT 47.470 185.170 47.730 185.490 ;
        RECT 48.850 185.170 49.110 185.490 ;
        RECT 46.550 175.310 46.810 175.630 ;
        RECT 45.170 171.910 45.430 172.230 ;
        RECT 44.710 169.530 44.970 169.850 ;
        RECT 44.710 167.830 44.970 168.150 ;
        RECT 44.250 167.490 44.510 167.810 ;
        RECT 43.790 167.150 44.050 167.470 ;
        RECT 42.870 166.810 43.130 167.130 ;
        RECT 43.330 166.810 43.590 167.130 ;
        RECT 41.950 165.110 42.210 165.430 ;
        RECT 42.410 165.110 42.670 165.430 ;
        RECT 42.010 164.830 42.150 165.110 ;
        RECT 42.010 164.690 43.070 164.830 ;
        RECT 41.950 160.690 42.210 161.010 ;
        RECT 41.490 154.460 41.750 154.550 ;
        RECT 41.090 154.320 41.750 154.460 ;
        RECT 40.570 153.210 40.830 153.530 ;
        RECT 41.090 151.150 41.230 154.320 ;
        RECT 41.490 154.230 41.750 154.320 ;
        RECT 41.490 152.530 41.750 152.850 ;
        RECT 37.810 150.830 38.070 151.150 ;
        RECT 41.030 150.830 41.290 151.150 ;
        RECT 36.890 147.430 37.150 147.750 ;
        RECT 37.340 147.575 37.620 147.945 ;
        RECT 35.050 147.090 35.310 147.410 ;
        RECT 35.970 147.090 36.230 147.410 ;
        RECT 34.590 145.390 34.850 145.710 ;
        RECT 34.590 144.710 34.850 145.030 ;
        RECT 34.130 143.350 34.390 143.670 ;
        RECT 32.750 142.330 33.010 142.650 ;
        RECT 34.650 142.560 34.790 144.710 ;
        RECT 35.110 143.330 35.250 147.090 ;
        RECT 35.510 145.390 35.770 145.710 ;
        RECT 35.050 143.010 35.310 143.330 ;
        RECT 34.650 142.420 35.250 142.560 ;
        RECT 24.470 141.650 24.730 141.970 ;
        RECT 32.180 141.115 33.720 141.485 ;
        RECT 35.110 140.270 35.250 142.420 ;
        RECT 30.910 139.950 31.170 140.270 ;
        RECT 35.050 139.950 35.310 140.270 ;
        RECT 24.930 138.930 25.190 139.250 ;
        RECT 24.990 136.870 25.130 138.930 ;
        RECT 28.880 138.395 30.420 138.765 ;
        RECT 25.850 137.570 26.110 137.890 ;
        RECT 23.550 136.550 23.810 136.870 ;
        RECT 24.930 136.550 25.190 136.870 ;
        RECT 24.010 136.210 24.270 136.530 ;
        RECT 23.090 134.850 23.350 135.170 ;
        RECT 22.630 133.490 22.890 133.810 ;
        RECT 23.150 131.770 23.290 134.850 ;
        RECT 23.090 131.450 23.350 131.770 ;
        RECT 23.150 129.730 23.290 131.450 ;
        RECT 24.070 131.430 24.210 136.210 ;
        RECT 24.930 134.850 25.190 135.170 ;
        RECT 24.990 132.790 25.130 134.850 ;
        RECT 25.910 134.150 26.050 137.570 ;
        RECT 29.990 136.890 30.250 137.210 ;
        RECT 26.310 136.210 26.570 136.530 ;
        RECT 26.770 136.210 27.030 136.530 ;
        RECT 28.150 136.210 28.410 136.530 ;
        RECT 26.370 135.510 26.510 136.210 ;
        RECT 26.310 135.190 26.570 135.510 ;
        RECT 25.850 133.830 26.110 134.150 ;
        RECT 24.930 132.470 25.190 132.790 ;
        RECT 24.010 131.110 24.270 131.430 ;
        RECT 25.910 130.070 26.050 133.830 ;
        RECT 26.830 131.430 26.970 136.210 ;
        RECT 27.690 135.190 27.950 135.510 ;
        RECT 27.230 134.850 27.490 135.170 ;
        RECT 27.290 133.810 27.430 134.850 ;
        RECT 27.750 134.830 27.890 135.190 ;
        RECT 27.690 134.510 27.950 134.830 ;
        RECT 27.230 133.490 27.490 133.810 ;
        RECT 28.210 132.190 28.350 136.210 ;
        RECT 30.050 135.170 30.190 136.890 ;
        RECT 29.990 134.850 30.250 135.170 ;
        RECT 30.970 133.810 31.110 139.950 ;
        RECT 31.830 139.610 32.090 139.930 ;
        RECT 31.370 138.930 31.630 139.250 ;
        RECT 31.430 134.830 31.570 138.930 ;
        RECT 31.890 135.510 32.030 139.610 ;
        RECT 35.110 137.210 35.250 139.950 ;
        RECT 35.570 139.590 35.710 145.390 ;
        RECT 36.030 145.030 36.170 147.090 ;
        RECT 36.950 145.710 37.090 147.430 ;
        RECT 36.890 145.390 37.150 145.710 ;
        RECT 35.970 144.710 36.230 145.030 ;
        RECT 36.950 144.690 37.090 145.390 ;
        RECT 36.890 144.370 37.150 144.690 ;
        RECT 35.970 142.330 36.230 142.650 ;
        RECT 36.430 142.330 36.690 142.650 ;
        RECT 35.510 139.270 35.770 139.590 ;
        RECT 36.030 138.230 36.170 142.330 ;
        RECT 36.490 140.270 36.630 142.330 ;
        RECT 36.890 140.290 37.150 140.610 ;
        RECT 36.430 139.950 36.690 140.270 ;
        RECT 35.970 137.910 36.230 138.230 ;
        RECT 35.970 137.230 36.230 137.550 ;
        RECT 35.050 136.890 35.310 137.210 ;
        RECT 34.130 136.550 34.390 136.870 ;
        RECT 32.180 135.675 33.720 136.045 ;
        RECT 34.190 135.510 34.330 136.550 ;
        RECT 34.590 136.210 34.850 136.530 ;
        RECT 31.830 135.190 32.090 135.510 ;
        RECT 34.130 135.190 34.390 135.510 ;
        RECT 31.370 134.510 31.630 134.830 ;
        RECT 31.820 134.655 32.100 135.025 ;
        RECT 33.660 134.655 33.940 135.025 ;
        RECT 34.650 134.910 34.790 136.210 ;
        RECT 34.190 134.830 34.790 134.910 ;
        RECT 34.130 134.770 34.790 134.830 ;
        RECT 31.890 134.490 32.030 134.655 ;
        RECT 33.670 134.510 33.930 134.655 ;
        RECT 34.130 134.510 34.390 134.770 ;
        RECT 31.830 134.400 32.090 134.490 ;
        RECT 31.830 134.260 32.490 134.400 ;
        RECT 31.830 134.170 32.090 134.260 ;
        RECT 31.370 133.830 31.630 134.150 ;
        RECT 30.910 133.490 31.170 133.810 ;
        RECT 28.880 132.955 30.420 133.325 ;
        RECT 28.210 132.050 29.270 132.190 ;
        RECT 31.430 132.110 31.570 133.830 ;
        RECT 31.830 133.490 32.090 133.810 ;
        RECT 31.890 132.790 32.030 133.490 ;
        RECT 31.830 132.470 32.090 132.790 ;
        RECT 32.350 132.190 32.490 134.260 ;
        RECT 29.130 131.770 29.270 132.050 ;
        RECT 31.370 131.790 31.630 132.110 ;
        RECT 31.890 132.050 32.490 132.190 ;
        RECT 29.070 131.450 29.330 131.770 ;
        RECT 26.770 131.110 27.030 131.430 ;
        RECT 29.530 131.110 29.790 131.430 ;
        RECT 26.830 130.070 26.970 131.110 ;
        RECT 28.610 130.770 28.870 131.090 ;
        RECT 25.850 129.750 26.110 130.070 ;
        RECT 26.770 129.750 27.030 130.070 ;
        RECT 23.090 129.410 23.350 129.730 ;
        RECT 23.150 126.330 23.290 129.410 ;
        RECT 28.670 129.390 28.810 130.770 ;
        RECT 29.590 129.730 29.730 131.110 ;
        RECT 29.530 129.410 29.790 129.730 ;
        RECT 28.610 129.070 28.870 129.390 ;
        RECT 28.880 127.515 30.420 127.885 ;
        RECT 23.090 126.010 23.350 126.330 ;
        RECT 31.370 126.010 31.630 126.330 ;
        RECT 16.650 123.970 16.910 124.290 ;
        RECT 16.710 119.190 16.850 123.970 ;
        RECT 20.790 123.290 21.050 123.610 ;
        RECT 17.570 121.590 17.830 121.910 ;
        RECT 16.650 118.870 16.910 119.190 ;
        RECT 17.630 118.850 17.770 121.590 ;
        RECT 20.850 119.190 20.990 123.290 ;
        RECT 22.630 122.950 22.890 123.270 ;
        RECT 21.710 122.610 21.970 122.930 ;
        RECT 21.770 120.890 21.910 122.610 ;
        RECT 22.690 120.890 22.830 122.950 ;
        RECT 24.470 122.610 24.730 122.930 ;
        RECT 24.930 122.610 25.190 122.930 ;
        RECT 21.710 120.570 21.970 120.890 ;
        RECT 22.630 120.570 22.890 120.890 ;
        RECT 20.790 118.870 21.050 119.190 ;
        RECT 17.570 118.530 17.830 118.850 ;
        RECT 17.570 117.170 17.830 117.490 ;
        RECT 17.630 112.730 17.770 117.170 ;
        RECT 20.850 115.110 20.990 118.870 ;
        RECT 22.690 118.510 22.830 120.570 ;
        RECT 23.090 118.590 23.350 118.850 ;
        RECT 24.010 118.590 24.270 118.850 ;
        RECT 23.090 118.530 24.270 118.590 ;
        RECT 22.630 118.190 22.890 118.510 ;
        RECT 23.150 118.450 24.210 118.530 ;
        RECT 21.710 117.910 21.970 118.170 ;
        RECT 21.710 117.850 24.210 117.910 ;
        RECT 21.770 117.770 24.210 117.850 ;
        RECT 24.070 117.490 24.210 117.770 ;
        RECT 23.550 117.170 23.810 117.490 ;
        RECT 24.010 117.170 24.270 117.490 ;
        RECT 23.610 116.470 23.750 117.170 ;
        RECT 21.710 116.150 21.970 116.470 ;
        RECT 23.550 116.150 23.810 116.470 ;
        RECT 20.790 114.790 21.050 115.110 ;
        RECT 19.410 114.450 19.670 114.770 ;
        RECT 19.470 113.070 19.610 114.450 ;
        RECT 19.410 112.750 19.670 113.070 ;
        RECT 17.570 112.410 17.830 112.730 ;
        RECT 17.630 110.350 17.770 112.410 ;
        RECT 20.850 110.590 20.990 114.790 ;
        RECT 20.390 110.450 20.990 110.590 ;
        RECT 17.570 110.030 17.830 110.350 ;
        RECT 17.630 102.870 17.770 110.030 ;
        RECT 19.410 109.350 19.670 109.670 ;
        RECT 18.490 109.010 18.750 109.330 ;
        RECT 18.550 107.970 18.690 109.010 ;
        RECT 19.470 108.310 19.610 109.350 ;
        RECT 19.410 107.990 19.670 108.310 ;
        RECT 18.490 107.650 18.750 107.970 ;
        RECT 20.390 106.610 20.530 110.450 ;
        RECT 21.770 108.310 21.910 116.150 ;
        RECT 24.530 116.130 24.670 122.610 ;
        RECT 24.990 120.210 25.130 122.610 ;
        RECT 28.880 122.075 30.420 122.445 ;
        RECT 25.390 121.590 25.650 121.910 ;
        RECT 24.930 119.890 25.190 120.210 ;
        RECT 24.470 115.810 24.730 116.130 ;
        RECT 24.990 112.730 25.130 119.890 ;
        RECT 25.450 115.450 25.590 121.590 ;
        RECT 25.850 121.250 26.110 121.570 ;
        RECT 25.910 118.850 26.050 121.250 ;
        RECT 31.430 120.890 31.570 126.010 ;
        RECT 31.890 122.930 32.030 132.050 ;
        RECT 34.190 131.770 34.330 134.510 ;
        RECT 34.590 134.230 34.850 134.490 ;
        RECT 35.110 134.230 35.250 136.890 ;
        RECT 34.590 134.170 35.250 134.230 ;
        RECT 34.650 134.090 35.250 134.170 ;
        RECT 34.130 131.450 34.390 131.770 ;
        RECT 34.650 130.830 34.790 134.090 ;
        RECT 36.030 133.810 36.170 137.230 ;
        RECT 36.490 135.510 36.630 139.950 ;
        RECT 36.950 136.530 37.090 140.290 ;
        RECT 36.890 136.210 37.150 136.530 ;
        RECT 36.430 135.190 36.690 135.510 ;
        RECT 35.970 133.490 36.230 133.810 ;
        RECT 35.510 132.470 35.770 132.790 ;
        RECT 34.190 130.690 34.790 130.830 ;
        RECT 32.180 130.235 33.720 130.605 ;
        RECT 32.180 124.795 33.720 125.165 ;
        RECT 32.290 122.950 32.550 123.270 ;
        RECT 31.830 122.610 32.090 122.930 ;
        RECT 30.440 120.375 30.720 120.745 ;
        RECT 31.370 120.570 31.630 120.890 ;
        RECT 32.350 120.630 32.490 122.950 ;
        RECT 31.890 120.550 32.490 120.630 ;
        RECT 30.510 118.850 30.650 120.375 ;
        RECT 30.910 120.230 31.170 120.550 ;
        RECT 31.890 120.490 32.550 120.550 ;
        RECT 25.850 118.530 26.110 118.850 ;
        RECT 30.450 118.530 30.710 118.850 ;
        RECT 25.910 115.450 26.050 118.530 ;
        RECT 30.970 117.490 31.110 120.230 ;
        RECT 31.370 119.890 31.630 120.210 ;
        RECT 26.770 117.170 27.030 117.490 ;
        RECT 30.910 117.170 31.170 117.490 ;
        RECT 25.390 115.130 25.650 115.450 ;
        RECT 25.850 115.130 26.110 115.450 ;
        RECT 25.450 114.770 25.590 115.130 ;
        RECT 25.390 114.450 25.650 114.770 ;
        RECT 24.930 112.410 25.190 112.730 ;
        RECT 25.450 112.050 25.590 114.450 ;
        RECT 25.910 113.410 26.050 115.130 ;
        RECT 26.830 113.750 26.970 117.170 ;
        RECT 28.880 116.635 30.420 117.005 ;
        RECT 27.230 115.130 27.490 115.450 ;
        RECT 28.150 115.130 28.410 115.450 ;
        RECT 26.770 113.430 27.030 113.750 ;
        RECT 25.850 113.090 26.110 113.410 ;
        RECT 24.010 111.730 24.270 112.050 ;
        RECT 25.390 111.730 25.650 112.050 ;
        RECT 24.070 110.010 24.210 111.730 ;
        RECT 25.910 110.350 26.050 113.090 ;
        RECT 25.850 110.030 26.110 110.350 ;
        RECT 27.290 110.010 27.430 115.130 ;
        RECT 24.010 109.690 24.270 110.010 ;
        RECT 27.230 109.690 27.490 110.010 ;
        RECT 23.550 109.350 23.810 109.670 ;
        RECT 21.710 107.990 21.970 108.310 ;
        RECT 23.610 107.630 23.750 109.350 ;
        RECT 24.070 107.630 24.210 109.690 ;
        RECT 26.310 109.010 26.570 109.330 ;
        RECT 26.370 107.630 26.510 109.010 ;
        RECT 28.210 108.310 28.350 115.130 ;
        RECT 29.530 114.790 29.790 115.110 ;
        RECT 29.590 113.750 29.730 114.790 ;
        RECT 30.970 114.770 31.110 117.170 ;
        RECT 31.430 115.450 31.570 119.890 ;
        RECT 31.890 118.510 32.030 120.490 ;
        RECT 32.290 120.230 32.550 120.490 ;
        RECT 32.180 119.355 33.720 119.725 ;
        RECT 34.190 118.850 34.330 130.690 ;
        RECT 35.570 129.730 35.710 132.470 ;
        RECT 35.510 129.410 35.770 129.730 ;
        RECT 36.030 128.370 36.170 133.490 ;
        RECT 36.430 131.110 36.690 131.430 ;
        RECT 36.490 130.070 36.630 131.110 ;
        RECT 36.430 129.750 36.690 130.070 ;
        RECT 35.970 128.050 36.230 128.370 ;
        RECT 37.410 124.390 37.550 147.575 ;
        RECT 37.870 145.710 38.010 150.830 ;
        RECT 41.090 150.470 41.230 150.830 ;
        RECT 41.030 150.150 41.290 150.470 ;
        RECT 38.270 149.810 38.530 150.130 ;
        RECT 40.570 149.810 40.830 150.130 ;
        RECT 38.330 148.430 38.470 149.810 ;
        RECT 38.270 148.110 38.530 148.430 ;
        RECT 40.630 148.090 40.770 149.810 ;
        RECT 38.730 147.770 38.990 148.090 ;
        RECT 40.570 147.770 40.830 148.090 ;
        RECT 41.030 147.770 41.290 148.090 ;
        RECT 37.810 145.390 38.070 145.710 ;
        RECT 37.870 145.030 38.010 145.390 ;
        RECT 37.810 144.710 38.070 145.030 ;
        RECT 38.790 143.330 38.930 147.770 ;
        RECT 40.110 147.090 40.370 147.410 ;
        RECT 40.170 146.050 40.310 147.090 ;
        RECT 39.190 145.730 39.450 146.050 ;
        RECT 40.110 145.730 40.370 146.050 ;
        RECT 39.250 143.670 39.390 145.730 ;
        RECT 41.090 145.370 41.230 147.770 ;
        RECT 41.030 145.050 41.290 145.370 ;
        RECT 41.550 144.600 41.690 152.530 ;
        RECT 41.090 144.460 41.690 144.600 ;
        RECT 39.190 143.350 39.450 143.670 ;
        RECT 38.730 143.010 38.990 143.330 ;
        RECT 38.790 140.950 38.930 143.010 ;
        RECT 38.730 140.630 38.990 140.950 ;
        RECT 36.490 124.250 37.550 124.390 ;
        RECT 35.050 121.590 35.310 121.910 ;
        RECT 35.110 120.890 35.250 121.590 ;
        RECT 36.490 120.890 36.630 124.250 ;
        RECT 40.570 122.610 40.830 122.930 ;
        RECT 40.110 121.590 40.370 121.910 ;
        RECT 37.350 121.480 37.610 121.570 ;
        RECT 38.730 121.480 38.990 121.570 ;
        RECT 37.350 121.340 38.990 121.480 ;
        RECT 37.350 121.250 37.610 121.340 ;
        RECT 38.730 121.250 38.990 121.340 ;
        RECT 40.170 120.890 40.310 121.590 ;
        RECT 40.630 121.230 40.770 122.610 ;
        RECT 40.570 120.910 40.830 121.230 ;
        RECT 35.050 120.570 35.310 120.890 ;
        RECT 34.130 118.530 34.390 118.850 ;
        RECT 31.830 118.190 32.090 118.510 ;
        RECT 34.190 115.450 34.330 118.530 ;
        RECT 35.110 117.490 35.250 120.570 ;
        RECT 35.510 120.230 35.770 120.550 ;
        RECT 35.960 120.375 36.240 120.745 ;
        RECT 36.430 120.570 36.690 120.890 ;
        RECT 35.970 120.230 36.230 120.375 ;
        RECT 37.350 120.230 37.610 120.550 ;
        RECT 38.720 120.375 39.000 120.745 ;
        RECT 40.110 120.570 40.370 120.890 ;
        RECT 35.050 117.170 35.310 117.490 ;
        RECT 35.570 116.130 35.710 120.230 ;
        RECT 36.430 119.890 36.690 120.210 ;
        RECT 35.970 118.190 36.230 118.510 ;
        RECT 36.030 116.470 36.170 118.190 ;
        RECT 35.970 116.150 36.230 116.470 ;
        RECT 35.510 115.810 35.770 116.130 ;
        RECT 36.490 115.790 36.630 119.890 ;
        RECT 36.890 118.870 37.150 119.190 ;
        RECT 36.950 116.470 37.090 118.870 ;
        RECT 36.890 116.150 37.150 116.470 ;
        RECT 36.430 115.470 36.690 115.790 ;
        RECT 36.890 115.470 37.150 115.790 ;
        RECT 31.370 115.130 31.630 115.450 ;
        RECT 34.130 115.130 34.390 115.450 ;
        RECT 36.950 114.770 37.090 115.470 ;
        RECT 37.410 115.450 37.550 120.230 ;
        RECT 38.790 119.190 38.930 120.375 ;
        RECT 38.730 118.870 38.990 119.190 ;
        RECT 39.650 117.170 39.910 117.490 ;
        RECT 40.110 117.170 40.370 117.490 ;
        RECT 38.270 115.810 38.530 116.130 ;
        RECT 37.350 115.130 37.610 115.450 ;
        RECT 30.910 114.450 31.170 114.770 ;
        RECT 35.510 114.450 35.770 114.770 ;
        RECT 36.890 114.450 37.150 114.770 ;
        RECT 30.970 113.750 31.110 114.450 ;
        RECT 32.180 113.915 33.720 114.285 ;
        RECT 29.530 113.430 29.790 113.750 ;
        RECT 30.910 113.430 31.170 113.750 ;
        RECT 35.570 113.410 35.710 114.450 ;
        RECT 35.510 113.090 35.770 113.410 ;
        RECT 30.910 112.750 31.170 113.070 ;
        RECT 28.880 111.195 30.420 111.565 ;
        RECT 30.970 110.010 31.110 112.750 ;
        RECT 36.950 110.010 37.090 114.450 ;
        RECT 28.610 109.690 28.870 110.010 ;
        RECT 30.910 109.690 31.170 110.010 ;
        RECT 36.890 109.690 37.150 110.010 ;
        RECT 28.150 107.990 28.410 108.310 ;
        RECT 20.790 107.310 21.050 107.630 ;
        RECT 23.550 107.310 23.810 107.630 ;
        RECT 24.010 107.310 24.270 107.630 ;
        RECT 24.930 107.310 25.190 107.630 ;
        RECT 26.310 107.310 26.570 107.630 ;
        RECT 20.850 107.030 20.990 107.310 ;
        RECT 20.850 106.890 21.450 107.030 ;
        RECT 20.330 106.290 20.590 106.610 ;
        RECT 20.790 106.290 21.050 106.610 ;
        RECT 20.390 105.590 20.530 106.290 ;
        RECT 20.330 105.270 20.590 105.590 ;
        RECT 17.570 102.550 17.830 102.870 ;
        RECT 17.630 99.470 17.770 102.550 ;
        RECT 20.390 101.510 20.530 105.270 ;
        RECT 20.850 104.230 20.990 106.290 ;
        RECT 21.310 104.570 21.450 106.890 ;
        RECT 23.610 104.570 23.750 107.310 ;
        RECT 24.990 106.950 25.130 107.310 ;
        RECT 28.670 106.950 28.810 109.690 ;
        RECT 30.910 109.010 31.170 109.330 ;
        RECT 30.970 107.970 31.110 109.010 ;
        RECT 32.180 108.475 33.720 108.845 ;
        RECT 30.910 107.650 31.170 107.970 ;
        RECT 34.130 107.650 34.390 107.970 ;
        RECT 24.930 106.630 25.190 106.950 ;
        RECT 28.610 106.630 28.870 106.950 ;
        RECT 28.880 105.755 30.420 106.125 ;
        RECT 29.990 105.500 30.250 105.590 ;
        RECT 30.970 105.500 31.110 107.650 ;
        RECT 34.190 105.590 34.330 107.650 ;
        RECT 35.510 106.290 35.770 106.610 ;
        RECT 36.430 106.290 36.690 106.610 ;
        RECT 35.570 105.590 35.710 106.290 ;
        RECT 29.990 105.360 31.110 105.500 ;
        RECT 29.990 105.270 30.250 105.360 ;
        RECT 34.130 105.270 34.390 105.590 ;
        RECT 35.510 105.270 35.770 105.590 ;
        RECT 21.250 104.250 21.510 104.570 ;
        RECT 23.550 104.250 23.810 104.570 ;
        RECT 20.790 103.910 21.050 104.230 ;
        RECT 20.850 101.510 20.990 103.910 ;
        RECT 21.310 102.190 21.450 104.250 ;
        RECT 24.010 103.570 24.270 103.890 ;
        RECT 24.070 102.870 24.210 103.570 ;
        RECT 24.010 102.550 24.270 102.870 ;
        RECT 21.250 101.870 21.510 102.190 ;
        RECT 20.330 101.190 20.590 101.510 ;
        RECT 20.790 101.190 21.050 101.510 ;
        RECT 18.950 100.850 19.210 101.170 ;
        RECT 17.570 99.150 17.830 99.470 ;
        RECT 19.010 99.130 19.150 100.850 ;
        RECT 21.310 100.230 21.450 101.870 ;
        RECT 30.050 101.170 30.190 105.270 ;
        RECT 34.130 104.250 34.390 104.570 ;
        RECT 32.180 103.035 33.720 103.405 ;
        RECT 30.910 102.210 31.170 102.530 ;
        RECT 30.970 101.510 31.110 102.210 ;
        RECT 34.190 102.190 34.330 104.250 ;
        RECT 35.510 103.910 35.770 104.230 ;
        RECT 35.570 102.870 35.710 103.910 ;
        RECT 35.510 102.550 35.770 102.870 ;
        RECT 34.130 101.870 34.390 102.190 ;
        RECT 30.910 101.190 31.170 101.510 ;
        RECT 36.490 101.170 36.630 106.290 ;
        RECT 36.950 102.870 37.090 109.690 ;
        RECT 38.330 107.630 38.470 115.810 ;
        RECT 39.710 115.110 39.850 117.170 ;
        RECT 39.650 114.790 39.910 115.110 ;
        RECT 40.170 108.310 40.310 117.170 ;
        RECT 41.090 115.450 41.230 144.460 ;
        RECT 42.010 142.650 42.150 160.690 ;
        RECT 42.930 143.670 43.070 164.690 ;
        RECT 43.390 162.030 43.530 166.810 ;
        RECT 43.850 165.090 43.990 167.150 ;
        RECT 43.790 164.770 44.050 165.090 ;
        RECT 44.310 164.410 44.450 167.490 ;
        RECT 44.770 164.750 44.910 167.830 ;
        RECT 45.230 166.450 45.370 171.910 ;
        RECT 45.630 168.850 45.890 169.170 ;
        RECT 45.170 166.130 45.430 166.450 ;
        RECT 44.710 164.430 44.970 164.750 ;
        RECT 43.790 164.090 44.050 164.410 ;
        RECT 44.250 164.090 44.510 164.410 ;
        RECT 43.850 163.730 43.990 164.090 ;
        RECT 43.790 163.410 44.050 163.730 ;
        RECT 43.850 162.030 43.990 163.410 ;
        RECT 43.330 161.710 43.590 162.030 ;
        RECT 43.790 161.710 44.050 162.030 ;
        RECT 44.770 153.530 44.910 164.430 ;
        RECT 45.690 163.730 45.830 168.850 ;
        RECT 46.610 167.130 46.750 175.310 ;
        RECT 47.070 173.250 47.210 185.170 ;
        RECT 47.010 172.930 47.270 173.250 ;
        RECT 47.530 172.230 47.670 185.170 ;
        RECT 48.910 183.790 49.050 185.170 ;
        RECT 49.370 184.130 49.510 191.290 ;
        RECT 50.290 189.230 50.430 192.310 ;
        RECT 51.210 189.570 51.350 193.330 ;
        RECT 60.410 192.630 60.550 194.350 ;
        RECT 60.350 192.310 60.610 192.630 ;
        RECT 62.250 191.950 62.390 194.350 ;
        RECT 62.190 191.630 62.450 191.950 ;
        RECT 63.170 191.270 63.310 198.770 ;
        RECT 64.950 196.730 65.210 197.050 ;
        RECT 66.330 196.730 66.590 197.050 ;
        RECT 63.570 194.010 63.830 194.330 ;
        RECT 64.030 194.010 64.290 194.330 ;
        RECT 63.630 191.465 63.770 194.010 ;
        RECT 51.610 190.950 51.870 191.270 ;
        RECT 63.110 190.950 63.370 191.270 ;
        RECT 63.560 191.095 63.840 191.465 ;
        RECT 63.570 190.950 63.830 191.095 ;
        RECT 51.150 189.250 51.410 189.570 ;
        RECT 50.230 188.910 50.490 189.230 ;
        RECT 50.690 188.910 50.950 189.230 ;
        RECT 49.310 183.810 49.570 184.130 ;
        RECT 48.850 183.470 49.110 183.790 ;
        RECT 49.370 180.390 49.510 183.810 ;
        RECT 49.310 180.070 49.570 180.390 ;
        RECT 49.770 180.070 50.030 180.390 ;
        RECT 49.370 178.690 49.510 180.070 ;
        RECT 49.310 178.370 49.570 178.690 ;
        RECT 49.830 176.310 49.970 180.070 ;
        RECT 49.770 175.990 50.030 176.310 ;
        RECT 50.290 175.970 50.430 188.910 ;
        RECT 49.310 175.650 49.570 175.970 ;
        RECT 50.230 175.650 50.490 175.970 ;
        RECT 48.850 172.930 49.110 173.250 ;
        RECT 47.470 171.910 47.730 172.230 ;
        RECT 48.390 171.910 48.650 172.230 ;
        RECT 47.010 170.210 47.270 170.530 ;
        RECT 47.070 167.470 47.210 170.210 ;
        RECT 48.450 168.150 48.590 171.910 ;
        RECT 48.910 168.345 49.050 172.930 ;
        RECT 48.390 167.830 48.650 168.150 ;
        RECT 48.840 167.975 49.120 168.345 ;
        RECT 47.470 167.490 47.730 167.810 ;
        RECT 47.010 167.150 47.270 167.470 ;
        RECT 46.550 166.810 46.810 167.130 ;
        RECT 46.610 165.090 46.750 166.810 ;
        RECT 46.550 164.770 46.810 165.090 ;
        RECT 47.530 164.410 47.670 167.490 ;
        RECT 48.910 167.130 49.050 167.975 ;
        RECT 48.850 166.810 49.110 167.130 ;
        RECT 49.370 164.750 49.510 175.650 ;
        RECT 50.230 174.970 50.490 175.290 ;
        RECT 49.770 172.590 50.030 172.910 ;
        RECT 49.830 170.190 49.970 172.590 ;
        RECT 50.290 172.570 50.430 174.970 ;
        RECT 50.750 174.350 50.890 188.910 ;
        RECT 51.210 186.850 51.350 189.250 ;
        RECT 51.670 188.550 51.810 190.950 ;
        RECT 52.990 190.610 53.250 190.930 ;
        RECT 51.610 188.230 51.870 188.550 ;
        RECT 51.150 186.530 51.410 186.850 ;
        RECT 53.050 180.390 53.190 190.610 ;
        RECT 63.170 188.890 63.310 190.950 ;
        RECT 63.110 188.570 63.370 188.890 ;
        RECT 63.570 186.490 63.830 186.510 ;
        RECT 64.090 186.490 64.230 194.010 ;
        RECT 64.490 193.330 64.750 193.650 ;
        RECT 64.550 191.950 64.690 193.330 ;
        RECT 65.010 192.290 65.150 196.730 ;
        RECT 66.390 192.630 66.530 196.730 ;
        RECT 66.850 195.350 66.990 199.450 ;
        RECT 67.310 196.710 67.450 199.790 ;
        RECT 67.250 196.390 67.510 196.710 ;
        RECT 67.310 195.350 67.450 196.390 ;
        RECT 66.790 195.030 67.050 195.350 ;
        RECT 67.250 195.030 67.510 195.350 ;
        RECT 66.330 192.310 66.590 192.630 ;
        RECT 67.710 192.310 67.970 192.630 ;
        RECT 64.950 191.970 65.210 192.290 ;
        RECT 65.870 191.970 66.130 192.290 ;
        RECT 64.490 191.630 64.750 191.950 ;
        RECT 65.930 189.910 66.070 191.970 ;
        RECT 65.870 189.590 66.130 189.910 ;
        RECT 67.770 189.230 67.910 192.310 ;
        RECT 68.230 192.290 68.370 199.790 ;
        RECT 73.750 199.430 73.890 210.670 ;
        RECT 77.370 199.790 77.630 200.110 ;
        RECT 116.470 199.790 116.730 200.110 ;
        RECT 74.610 199.450 74.870 199.770 ;
        RECT 73.690 199.110 73.950 199.430 ;
        RECT 70.470 197.410 70.730 197.730 ;
        RECT 69.550 196.730 69.810 197.050 ;
        RECT 69.090 196.050 69.350 196.370 ;
        RECT 68.630 194.350 68.890 194.670 ;
        RECT 68.690 192.630 68.830 194.350 ;
        RECT 68.630 192.310 68.890 192.630 ;
        RECT 68.170 191.970 68.430 192.290 ;
        RECT 68.170 191.290 68.430 191.610 ;
        RECT 67.710 188.910 67.970 189.230 ;
        RECT 68.230 188.890 68.370 191.290 ;
        RECT 69.150 189.140 69.290 196.050 ;
        RECT 69.610 195.010 69.750 196.730 ;
        RECT 70.010 195.030 70.270 195.350 ;
        RECT 69.550 194.690 69.810 195.010 ;
        RECT 69.610 191.610 69.750 194.690 ;
        RECT 70.070 192.630 70.210 195.030 ;
        RECT 70.530 194.670 70.670 197.410 ;
        RECT 73.750 196.710 73.890 199.110 ;
        RECT 74.150 198.770 74.410 199.090 ;
        RECT 74.210 198.070 74.350 198.770 ;
        RECT 74.150 197.750 74.410 198.070 ;
        RECT 73.690 196.390 73.950 196.710 ;
        RECT 74.670 196.370 74.810 199.450 ;
        RECT 74.610 196.050 74.870 196.370 ;
        RECT 70.470 194.350 70.730 194.670 ;
        RECT 70.010 192.310 70.270 192.630 ;
        RECT 69.550 191.290 69.810 191.610 ;
        RECT 70.070 189.570 70.210 192.310 ;
        RECT 70.530 191.610 70.670 194.350 ;
        RECT 74.670 194.330 74.810 196.050 ;
        RECT 74.610 194.010 74.870 194.330 ;
        RECT 75.530 194.010 75.790 194.330 ;
        RECT 72.770 193.330 73.030 193.650 ;
        RECT 73.230 193.330 73.490 193.650 ;
        RECT 72.830 191.610 72.970 193.330 ;
        RECT 73.290 191.950 73.430 193.330 ;
        RECT 73.230 191.630 73.490 191.950 ;
        RECT 74.670 191.610 74.810 194.010 ;
        RECT 75.590 193.505 75.730 194.010 ;
        RECT 75.520 193.135 75.800 193.505 ;
        RECT 76.910 193.330 77.170 193.650 ;
        RECT 76.450 192.310 76.710 192.630 ;
        RECT 76.510 191.610 76.650 192.310 ;
        RECT 76.970 191.950 77.110 193.330 ;
        RECT 76.910 191.630 77.170 191.950 ;
        RECT 70.470 191.290 70.730 191.610 ;
        RECT 71.390 191.465 71.650 191.610 ;
        RECT 71.380 191.095 71.660 191.465 ;
        RECT 72.770 191.290 73.030 191.610 ;
        RECT 74.610 191.290 74.870 191.610 ;
        RECT 76.450 191.290 76.710 191.610 ;
        RECT 73.690 190.950 73.950 191.270 ;
        RECT 73.750 189.910 73.890 190.950 ;
        RECT 74.670 190.930 74.810 191.290 ;
        RECT 74.610 190.610 74.870 190.930 ;
        RECT 76.450 190.670 76.710 190.930 ;
        RECT 77.430 190.670 77.570 199.790 ;
        RECT 79.210 198.770 79.470 199.090 ;
        RECT 113.710 198.770 113.970 199.090 ;
        RECT 77.830 194.350 78.090 194.670 ;
        RECT 77.890 192.630 78.030 194.350 ;
        RECT 77.830 192.310 78.090 192.630 ;
        RECT 79.270 191.465 79.410 198.770 ;
        RECT 104.050 197.070 104.310 197.390 ;
        RECT 95.770 196.960 96.030 197.050 ;
        RECT 95.770 196.820 96.430 196.960 ;
        RECT 95.770 196.730 96.030 196.820 ;
        RECT 80.130 196.050 80.390 196.370 ;
        RECT 90.710 196.050 90.970 196.370 ;
        RECT 91.630 196.050 91.890 196.370 ;
        RECT 80.190 195.010 80.330 196.050 ;
        RECT 80.130 194.690 80.390 195.010 ;
        RECT 90.250 194.690 90.510 195.010 ;
        RECT 80.590 194.350 80.850 194.670 ;
        RECT 81.510 194.350 81.770 194.670 ;
        RECT 79.200 191.095 79.480 191.465 ;
        RECT 76.450 190.610 77.570 190.670 ;
        RECT 76.510 190.530 77.570 190.610 ;
        RECT 73.690 189.590 73.950 189.910 ;
        RECT 70.010 189.250 70.270 189.570 ;
        RECT 69.150 189.000 69.750 189.140 ;
        RECT 64.950 188.570 65.210 188.890 ;
        RECT 68.170 188.570 68.430 188.890 ;
        RECT 63.570 186.350 64.230 186.490 ;
        RECT 63.570 186.190 63.830 186.350 ;
        RECT 53.450 185.850 53.710 186.170 ;
        RECT 53.510 184.470 53.650 185.850 ;
        RECT 63.630 185.490 63.770 186.190 ;
        RECT 65.010 186.170 65.150 188.570 ;
        RECT 66.330 187.890 66.590 188.210 ;
        RECT 67.250 187.890 67.510 188.210 ;
        RECT 67.710 187.890 67.970 188.210 ;
        RECT 64.030 185.850 64.290 186.170 ;
        RECT 64.950 185.850 65.210 186.170 ;
        RECT 58.510 185.170 58.770 185.490 ;
        RECT 63.570 185.170 63.830 185.490 ;
        RECT 53.450 184.150 53.710 184.470 ;
        RECT 52.530 180.070 52.790 180.390 ;
        RECT 52.990 180.070 53.250 180.390 ;
        RECT 51.150 177.010 51.410 177.330 ;
        RECT 51.210 175.290 51.350 177.010 ;
        RECT 52.590 175.630 52.730 180.070 ;
        RECT 53.510 178.690 53.650 184.150 ;
        RECT 55.750 183.130 56.010 183.450 ;
        RECT 55.290 182.450 55.550 182.770 ;
        RECT 55.350 181.410 55.490 182.450 ;
        RECT 55.290 181.090 55.550 181.410 ;
        RECT 55.810 180.730 55.950 183.130 ;
        RECT 58.570 180.730 58.710 185.170 ;
        RECT 64.090 181.750 64.230 185.850 ;
        RECT 66.390 185.830 66.530 187.890 ;
        RECT 67.310 186.170 67.450 187.890 ;
        RECT 67.250 186.080 67.510 186.170 ;
        RECT 66.850 185.940 67.510 186.080 ;
        RECT 66.330 185.510 66.590 185.830 ;
        RECT 66.390 183.790 66.530 185.510 ;
        RECT 66.850 184.470 66.990 185.940 ;
        RECT 67.250 185.850 67.510 185.940 ;
        RECT 67.250 185.170 67.510 185.490 ;
        RECT 67.310 184.470 67.450 185.170 ;
        RECT 66.790 184.150 67.050 184.470 ;
        RECT 67.250 184.150 67.510 184.470 ;
        RECT 67.770 183.790 67.910 187.890 ;
        RECT 68.230 183.790 68.370 188.570 ;
        RECT 69.090 188.230 69.350 188.550 ;
        RECT 69.150 186.850 69.290 188.230 ;
        RECT 69.090 186.530 69.350 186.850 ;
        RECT 69.150 184.470 69.290 186.530 ;
        RECT 69.610 186.170 69.750 189.000 ;
        RECT 76.970 188.210 77.110 190.530 ;
        RECT 77.370 189.250 77.630 189.570 ;
        RECT 76.910 187.890 77.170 188.210 ;
        RECT 69.550 185.850 69.810 186.170 ;
        RECT 70.470 185.850 70.730 186.170 ;
        RECT 71.850 185.850 72.110 186.170 ;
        RECT 75.530 185.850 75.790 186.170 ;
        RECT 69.090 184.150 69.350 184.470 ;
        RECT 66.330 183.470 66.590 183.790 ;
        RECT 67.710 183.470 67.970 183.790 ;
        RECT 68.170 183.470 68.430 183.790 ;
        RECT 67.770 181.750 67.910 183.470 ;
        RECT 64.030 181.430 64.290 181.750 ;
        RECT 67.710 181.430 67.970 181.750 ;
        RECT 55.750 180.410 56.010 180.730 ;
        RECT 58.510 180.410 58.770 180.730 ;
        RECT 54.370 179.730 54.630 180.050 ;
        RECT 65.410 179.730 65.670 180.050 ;
        RECT 67.250 179.730 67.510 180.050 ;
        RECT 54.430 179.030 54.570 179.730 ;
        RECT 54.370 178.710 54.630 179.030 ;
        RECT 52.990 178.370 53.250 178.690 ;
        RECT 53.450 178.370 53.710 178.690 ;
        RECT 65.470 178.545 65.610 179.730 ;
        RECT 52.530 175.310 52.790 175.630 ;
        RECT 53.050 175.290 53.190 178.370 ;
        RECT 65.400 178.175 65.680 178.545 ;
        RECT 60.350 177.690 60.610 178.010 ;
        RECT 60.410 175.290 60.550 177.690 ;
        RECT 51.150 174.970 51.410 175.290 ;
        RECT 52.990 174.970 53.250 175.290 ;
        RECT 60.350 174.970 60.610 175.290 ;
        RECT 63.110 174.970 63.370 175.290 ;
        RECT 65.410 174.970 65.670 175.290 ;
        RECT 51.150 174.350 51.410 174.610 ;
        RECT 50.750 174.290 51.410 174.350 ;
        RECT 50.750 174.210 51.350 174.290 ;
        RECT 51.210 172.570 51.350 174.210 ;
        RECT 50.230 172.250 50.490 172.570 ;
        RECT 51.150 172.250 51.410 172.570 ;
        RECT 50.290 170.530 50.430 172.250 ;
        RECT 50.230 170.210 50.490 170.530 ;
        RECT 49.770 169.870 50.030 170.190 ;
        RECT 49.830 169.170 49.970 169.870 ;
        RECT 49.770 168.850 50.030 169.170 ;
        RECT 49.830 168.150 49.970 168.850 ;
        RECT 49.770 167.830 50.030 168.150 ;
        RECT 50.690 167.150 50.950 167.470 ;
        RECT 50.230 166.130 50.490 166.450 ;
        RECT 49.310 164.430 49.570 164.750 ;
        RECT 47.470 164.090 47.730 164.410 ;
        RECT 45.630 163.410 45.890 163.730 ;
        RECT 46.090 163.410 46.350 163.730 ;
        RECT 45.690 162.030 45.830 163.410 ;
        RECT 45.630 161.710 45.890 162.030 ;
        RECT 46.150 161.010 46.290 163.410 ;
        RECT 50.290 161.690 50.430 166.130 ;
        RECT 50.750 162.710 50.890 167.150 ;
        RECT 51.210 164.070 51.350 172.250 ;
        RECT 59.890 171.910 60.150 172.230 ;
        RECT 59.430 171.570 59.690 171.890 ;
        RECT 52.530 169.530 52.790 169.850 ;
        RECT 58.970 169.530 59.230 169.850 ;
        RECT 51.610 168.850 51.870 169.170 ;
        RECT 51.670 164.750 51.810 168.850 ;
        RECT 52.060 167.975 52.340 168.345 ;
        RECT 52.070 167.830 52.330 167.975 ;
        RECT 52.590 165.090 52.730 169.530 ;
        RECT 56.210 169.190 56.470 169.510 ;
        RECT 56.270 165.430 56.410 169.190 ;
        RECT 58.510 167.040 58.770 167.130 ;
        RECT 59.030 167.040 59.170 169.530 ;
        RECT 59.490 167.810 59.630 171.570 ;
        RECT 59.950 167.810 60.090 171.910 ;
        RECT 61.730 171.570 61.990 171.890 ;
        RECT 60.350 170.550 60.610 170.870 ;
        RECT 59.430 167.490 59.690 167.810 ;
        RECT 59.890 167.490 60.150 167.810 ;
        RECT 60.410 167.130 60.550 170.550 ;
        RECT 61.790 170.530 61.930 171.570 ;
        RECT 61.730 170.210 61.990 170.530 ;
        RECT 58.510 166.900 59.170 167.040 ;
        RECT 58.510 166.810 58.770 166.900 ;
        RECT 58.050 166.130 58.310 166.450 ;
        RECT 56.210 165.110 56.470 165.430 ;
        RECT 52.530 164.770 52.790 165.090 ;
        RECT 51.610 164.430 51.870 164.750 ;
        RECT 51.150 163.750 51.410 164.070 ;
        RECT 50.690 162.390 50.950 162.710 ;
        RECT 52.590 162.030 52.730 164.770 ;
        RECT 58.110 164.410 58.250 166.130 ;
        RECT 59.030 164.410 59.170 166.900 ;
        RECT 60.350 166.810 60.610 167.130 ;
        RECT 58.050 164.090 58.310 164.410 ;
        RECT 58.970 164.090 59.230 164.410 ;
        RECT 63.170 164.070 63.310 174.970 ;
        RECT 64.950 174.630 65.210 174.950 ;
        RECT 65.010 172.910 65.150 174.630 ;
        RECT 65.470 172.910 65.610 174.970 ;
        RECT 67.310 174.950 67.450 179.730 ;
        RECT 68.230 175.290 68.370 183.470 ;
        RECT 69.610 183.360 69.750 185.850 ;
        RECT 68.690 183.220 69.750 183.360 ;
        RECT 68.690 180.730 68.830 183.220 ;
        RECT 69.090 182.450 69.350 182.770 ;
        RECT 68.630 180.410 68.890 180.730 ;
        RECT 68.170 174.970 68.430 175.290 ;
        RECT 67.250 174.630 67.510 174.950 ;
        RECT 64.950 172.590 65.210 172.910 ;
        RECT 65.410 172.590 65.670 172.910 ;
        RECT 69.150 169.510 69.290 182.450 ;
        RECT 70.010 180.410 70.270 180.730 ;
        RECT 70.070 178.690 70.210 180.410 ;
        RECT 70.530 179.030 70.670 185.850 ;
        RECT 71.910 184.470 72.050 185.850 ;
        RECT 73.690 185.170 73.950 185.490 ;
        RECT 71.850 184.150 72.110 184.470 ;
        RECT 71.390 183.810 71.650 184.130 ;
        RECT 71.450 181.750 71.590 183.810 ;
        RECT 71.910 181.750 72.050 184.150 ;
        RECT 72.310 183.470 72.570 183.790 ;
        RECT 71.390 181.430 71.650 181.750 ;
        RECT 71.850 181.430 72.110 181.750 ;
        RECT 70.930 181.090 71.190 181.410 ;
        RECT 70.470 178.710 70.730 179.030 ;
        RECT 70.990 178.690 71.130 181.090 ;
        RECT 71.380 180.895 71.660 181.265 ;
        RECT 71.390 180.750 71.650 180.895 ;
        RECT 71.850 180.410 72.110 180.730 ;
        RECT 71.910 179.225 72.050 180.410 ;
        RECT 71.840 178.855 72.120 179.225 ;
        RECT 72.370 179.030 72.510 183.470 ;
        RECT 72.770 180.750 73.030 181.070 ;
        RECT 73.220 180.895 73.500 181.265 ;
        RECT 72.310 178.710 72.570 179.030 ;
        RECT 70.010 178.370 70.270 178.690 ;
        RECT 70.930 178.370 71.190 178.690 ;
        RECT 70.070 173.590 70.210 178.370 ;
        RECT 72.310 177.690 72.570 178.010 ;
        RECT 70.470 177.010 70.730 177.330 ;
        RECT 70.010 173.270 70.270 173.590 ;
        RECT 70.070 172.990 70.210 173.270 ;
        RECT 69.610 172.850 70.210 172.990 ;
        RECT 69.610 170.190 69.750 172.850 ;
        RECT 70.530 170.870 70.670 177.010 ;
        RECT 72.370 175.290 72.510 177.690 ;
        RECT 72.830 177.330 72.970 180.750 ;
        RECT 72.770 177.010 73.030 177.330 ;
        RECT 72.310 174.970 72.570 175.290 ;
        RECT 73.290 172.690 73.430 180.895 ;
        RECT 73.750 178.350 73.890 185.170 ;
        RECT 75.590 184.470 75.730 185.850 ;
        RECT 75.530 184.150 75.790 184.470 ;
        RECT 75.070 183.810 75.330 184.130 ;
        RECT 75.130 181.750 75.270 183.810 ;
        RECT 75.990 182.450 76.250 182.770 ;
        RECT 76.910 182.450 77.170 182.770 ;
        RECT 75.070 181.430 75.330 181.750 ;
        RECT 75.130 181.070 75.730 181.150 ;
        RECT 76.050 181.070 76.190 182.450 ;
        RECT 75.070 181.010 75.730 181.070 ;
        RECT 75.070 180.750 75.330 181.010 ;
        RECT 73.690 178.030 73.950 178.350 ;
        RECT 75.060 178.175 75.340 178.545 ;
        RECT 75.590 178.350 75.730 181.010 ;
        RECT 75.990 180.750 76.250 181.070 ;
        RECT 76.440 180.895 76.720 181.265 ;
        RECT 75.070 178.030 75.330 178.175 ;
        RECT 75.530 178.030 75.790 178.350 ;
        RECT 75.590 177.750 75.730 178.030 ;
        RECT 74.670 177.670 75.730 177.750 ;
        RECT 74.610 177.610 75.730 177.670 ;
        RECT 74.610 177.350 74.870 177.610 ;
        RECT 75.070 177.010 75.330 177.330 ;
        RECT 73.290 172.550 73.890 172.690 ;
        RECT 70.470 170.550 70.730 170.870 ;
        RECT 70.010 170.210 70.270 170.530 ;
        RECT 69.550 169.870 69.810 170.190 ;
        RECT 68.170 169.190 68.430 169.510 ;
        RECT 69.090 169.190 69.350 169.510 ;
        RECT 66.330 168.850 66.590 169.170 ;
        RECT 67.250 168.850 67.510 169.170 ;
        RECT 62.650 163.750 62.910 164.070 ;
        RECT 63.110 163.750 63.370 164.070 ;
        RECT 52.530 161.710 52.790 162.030 ;
        RECT 62.710 161.690 62.850 163.750 ;
        RECT 63.170 162.710 63.310 163.750 ;
        RECT 63.110 162.390 63.370 162.710 ;
        RECT 47.470 161.370 47.730 161.690 ;
        RECT 50.230 161.370 50.490 161.690 ;
        RECT 62.650 161.370 62.910 161.690 ;
        RECT 46.090 160.690 46.350 161.010 ;
        RECT 44.710 153.210 44.970 153.530 ;
        RECT 46.090 150.830 46.350 151.150 ;
        RECT 45.170 147.090 45.430 147.410 ;
        RECT 45.230 145.710 45.370 147.090 ;
        RECT 46.150 145.710 46.290 150.830 ;
        RECT 45.170 145.390 45.430 145.710 ;
        RECT 46.090 145.390 46.350 145.710 ;
        RECT 46.550 145.390 46.810 145.710 ;
        RECT 44.250 144.710 44.510 145.030 ;
        RECT 42.870 143.350 43.130 143.670 ;
        RECT 41.950 142.330 42.210 142.650 ;
        RECT 42.010 139.930 42.150 142.330 ;
        RECT 41.950 139.610 42.210 139.930 ;
        RECT 44.310 139.250 44.450 144.710 ;
        RECT 45.230 143.670 45.370 145.390 ;
        RECT 45.170 143.350 45.430 143.670 ;
        RECT 45.170 142.330 45.430 142.650 ;
        RECT 44.250 138.930 44.510 139.250 ;
        RECT 43.790 137.230 44.050 137.550 ;
        RECT 41.490 136.210 41.750 136.530 ;
        RECT 41.550 134.830 41.690 136.210 ;
        RECT 41.490 134.510 41.750 134.830 ;
        RECT 41.550 132.790 41.690 134.510 ;
        RECT 41.490 132.470 41.750 132.790 ;
        RECT 41.550 131.430 41.690 132.470 ;
        RECT 43.850 131.430 43.990 137.230 ;
        RECT 44.310 132.790 44.450 138.930 ;
        RECT 44.250 132.470 44.510 132.790 ;
        RECT 41.490 131.110 41.750 131.430 ;
        RECT 43.790 131.110 44.050 131.430 ;
        RECT 44.700 131.255 44.980 131.625 ;
        RECT 44.710 131.110 44.970 131.255 ;
        RECT 43.330 129.640 43.590 129.730 ;
        RECT 43.850 129.640 43.990 131.110 ;
        RECT 45.230 130.070 45.370 142.330 ;
        RECT 46.610 140.610 46.750 145.390 ;
        RECT 47.010 144.370 47.270 144.690 ;
        RECT 47.070 142.650 47.210 144.370 ;
        RECT 47.010 142.330 47.270 142.650 ;
        RECT 47.070 140.950 47.210 142.330 ;
        RECT 47.010 140.630 47.270 140.950 ;
        RECT 46.550 140.290 46.810 140.610 ;
        RECT 47.010 134.510 47.270 134.830 ;
        RECT 46.090 134.170 46.350 134.490 ;
        RECT 46.150 131.430 46.290 134.170 ;
        RECT 47.070 132.790 47.210 134.510 ;
        RECT 47.010 132.470 47.270 132.790 ;
        RECT 46.090 131.110 46.350 131.430 ;
        RECT 46.150 130.070 46.290 131.110 ;
        RECT 45.170 129.750 45.430 130.070 ;
        RECT 46.090 129.750 46.350 130.070 ;
        RECT 43.330 129.500 43.990 129.640 ;
        RECT 43.330 129.410 43.590 129.500 ;
        RECT 41.490 128.730 41.750 129.050 ;
        RECT 41.550 120.210 41.690 128.730 ;
        RECT 47.530 121.570 47.670 161.370 ;
        RECT 62.710 156.250 62.850 161.370 ;
        RECT 65.870 157.970 66.130 158.290 ;
        RECT 62.650 155.930 62.910 156.250 ;
        RECT 50.690 153.210 50.950 153.530 ;
        RECT 48.390 148.790 48.650 149.110 ;
        RECT 47.930 147.770 48.190 148.090 ;
        RECT 47.990 146.050 48.130 147.770 ;
        RECT 47.930 145.730 48.190 146.050 ;
        RECT 47.930 145.050 48.190 145.370 ;
        RECT 47.990 143.670 48.130 145.050 ;
        RECT 48.450 145.030 48.590 148.790 ;
        RECT 50.750 148.090 50.890 153.210 ;
        RECT 52.990 152.870 53.250 153.190 ;
        RECT 55.750 152.870 56.010 153.190 ;
        RECT 52.530 152.530 52.790 152.850 ;
        RECT 50.690 147.770 50.950 148.090 ;
        RECT 49.310 145.960 49.570 146.050 ;
        RECT 49.310 145.820 49.970 145.960 ;
        RECT 49.310 145.730 49.570 145.820 ;
        RECT 48.390 144.710 48.650 145.030 ;
        RECT 49.310 144.370 49.570 144.690 ;
        RECT 47.930 143.350 48.190 143.670 ;
        RECT 49.370 142.990 49.510 144.370 ;
        RECT 49.310 142.670 49.570 142.990 ;
        RECT 48.390 142.330 48.650 142.650 ;
        RECT 47.930 141.650 48.190 141.970 ;
        RECT 47.990 140.270 48.130 141.650 ;
        RECT 48.450 140.950 48.590 142.330 ;
        RECT 48.850 141.990 49.110 142.310 ;
        RECT 48.390 140.630 48.650 140.950 ;
        RECT 47.930 139.950 48.190 140.270 ;
        RECT 47.930 134.510 48.190 134.830 ;
        RECT 47.990 132.110 48.130 134.510 ;
        RECT 48.910 134.490 49.050 141.990 ;
        RECT 49.830 140.950 49.970 145.820 ;
        RECT 50.230 145.050 50.490 145.370 ;
        RECT 50.290 141.970 50.430 145.050 ;
        RECT 50.230 141.650 50.490 141.970 ;
        RECT 49.770 140.630 50.030 140.950 ;
        RECT 50.750 140.610 50.890 147.770 ;
        RECT 51.610 145.730 51.870 146.050 ;
        RECT 51.670 143.670 51.810 145.730 ;
        RECT 52.070 145.620 52.330 145.710 ;
        RECT 52.590 145.620 52.730 152.530 ;
        RECT 52.070 145.480 52.730 145.620 ;
        RECT 52.070 145.390 52.330 145.480 ;
        RECT 51.610 143.350 51.870 143.670 ;
        RECT 51.150 141.990 51.410 142.310 ;
        RECT 51.210 140.950 51.350 141.990 ;
        RECT 51.150 140.630 51.410 140.950 ;
        RECT 50.690 140.290 50.950 140.610 ;
        RECT 50.230 139.950 50.490 140.270 ;
        RECT 50.290 137.210 50.430 139.950 ;
        RECT 49.310 136.890 49.570 137.210 ;
        RECT 50.230 136.890 50.490 137.210 ;
        RECT 48.850 134.170 49.110 134.490 ;
        RECT 49.370 132.790 49.510 136.890 ;
        RECT 50.290 135.510 50.430 136.890 ;
        RECT 50.230 135.190 50.490 135.510 ;
        RECT 49.310 132.470 49.570 132.790 ;
        RECT 47.930 131.790 48.190 132.110 ;
        RECT 47.990 131.090 48.130 131.790 ;
        RECT 49.370 131.770 49.510 132.470 ;
        RECT 50.230 132.130 50.490 132.450 ;
        RECT 48.850 131.625 49.110 131.770 ;
        RECT 48.840 131.255 49.120 131.625 ;
        RECT 49.310 131.450 49.570 131.770 ;
        RECT 47.930 130.770 48.190 131.090 ;
        RECT 50.290 129.730 50.430 132.130 ;
        RECT 50.750 132.110 50.890 140.290 ;
        RECT 51.610 136.890 51.870 137.210 ;
        RECT 51.150 136.210 51.410 136.530 ;
        RECT 50.690 131.790 50.950 132.110 ;
        RECT 51.210 131.430 51.350 136.210 ;
        RECT 51.670 135.170 51.810 136.890 ;
        RECT 52.130 135.420 52.270 145.390 ;
        RECT 53.050 144.690 53.190 152.870 ;
        RECT 53.450 150.830 53.710 151.150 ;
        RECT 53.910 150.830 54.170 151.150 ;
        RECT 53.510 145.710 53.650 150.830 ;
        RECT 53.450 145.390 53.710 145.710 ;
        RECT 52.990 144.370 53.250 144.690 ;
        RECT 52.530 140.290 52.790 140.610 ;
        RECT 52.590 138.230 52.730 140.290 ;
        RECT 52.530 137.910 52.790 138.230 ;
        RECT 53.050 137.550 53.190 144.370 ;
        RECT 53.510 142.990 53.650 145.390 ;
        RECT 53.970 144.690 54.110 150.830 ;
        RECT 55.810 149.110 55.950 152.870 ;
        RECT 58.970 152.530 59.230 152.850 ;
        RECT 59.030 151.150 59.170 152.530 ;
        RECT 62.710 151.490 62.850 155.930 ;
        RECT 62.650 151.170 62.910 151.490 ;
        RECT 65.930 151.150 66.070 157.970 ;
        RECT 66.390 156.930 66.530 168.850 ;
        RECT 67.310 166.450 67.450 168.850 ;
        RECT 67.250 166.130 67.510 166.450 ;
        RECT 68.230 165.090 68.370 169.190 ;
        RECT 70.070 168.150 70.210 170.210 ;
        RECT 69.090 167.830 69.350 168.150 ;
        RECT 70.010 167.830 70.270 168.150 ;
        RECT 69.150 167.470 69.290 167.830 ;
        RECT 70.530 167.550 70.670 170.550 ;
        RECT 73.230 169.530 73.490 169.850 ;
        RECT 72.770 168.850 73.030 169.170 ;
        RECT 69.090 167.150 69.350 167.470 ;
        RECT 69.610 167.410 70.670 167.550 ;
        RECT 72.830 167.470 72.970 168.850 ;
        RECT 73.290 168.150 73.430 169.530 ;
        RECT 73.230 167.830 73.490 168.150 ;
        RECT 73.750 167.470 73.890 172.550 ;
        RECT 74.150 172.250 74.410 172.570 ;
        RECT 69.610 167.130 69.750 167.410 ;
        RECT 69.550 166.810 69.810 167.130 ;
        RECT 70.530 166.450 70.670 167.410 ;
        RECT 72.770 167.150 73.030 167.470 ;
        RECT 73.690 167.150 73.950 167.470 ;
        RECT 70.930 166.810 71.190 167.130 ;
        RECT 70.470 166.130 70.730 166.450 ;
        RECT 70.530 165.430 70.670 166.130 ;
        RECT 70.990 165.430 71.130 166.810 ;
        RECT 72.310 166.470 72.570 166.790 ;
        RECT 70.470 165.110 70.730 165.430 ;
        RECT 70.930 165.110 71.190 165.430 ;
        RECT 68.170 164.770 68.430 165.090 ;
        RECT 70.010 163.410 70.270 163.730 ;
        RECT 66.790 161.710 67.050 162.030 ;
        RECT 66.850 159.990 66.990 161.710 ;
        RECT 69.090 160.690 69.350 161.010 ;
        RECT 66.790 159.670 67.050 159.990 ;
        RECT 69.150 159.310 69.290 160.690 ;
        RECT 70.070 159.310 70.210 163.410 ;
        RECT 72.370 162.030 72.510 166.470 ;
        RECT 72.310 161.710 72.570 162.030 ;
        RECT 72.370 161.010 72.510 161.710 ;
        RECT 72.310 160.690 72.570 161.010 ;
        RECT 69.090 158.990 69.350 159.310 ;
        RECT 70.010 158.990 70.270 159.310 ;
        RECT 70.070 157.270 70.210 158.990 ;
        RECT 72.770 158.310 73.030 158.630 ;
        RECT 71.850 157.970 72.110 158.290 ;
        RECT 72.310 157.970 72.570 158.290 ;
        RECT 70.010 156.950 70.270 157.270 ;
        RECT 66.330 156.610 66.590 156.930 ;
        RECT 66.390 154.550 66.530 156.610 ;
        RECT 68.170 156.270 68.430 156.590 ;
        RECT 66.790 155.250 67.050 155.570 ;
        RECT 66.330 154.230 66.590 154.550 ;
        RECT 66.850 151.150 66.990 155.250 ;
        RECT 68.230 154.550 68.370 156.270 ;
        RECT 69.090 155.250 69.350 155.570 ;
        RECT 68.170 154.230 68.430 154.550 ;
        RECT 69.150 153.530 69.290 155.250 ;
        RECT 71.910 154.210 72.050 157.970 ;
        RECT 71.850 153.890 72.110 154.210 ;
        RECT 72.370 153.870 72.510 157.970 ;
        RECT 72.310 153.550 72.570 153.870 ;
        RECT 69.090 153.210 69.350 153.530 ;
        RECT 69.550 153.210 69.810 153.530 ;
        RECT 69.610 151.490 69.750 153.210 ;
        RECT 69.550 151.170 69.810 151.490 ;
        RECT 56.670 150.830 56.930 151.150 ;
        RECT 58.970 150.830 59.230 151.150 ;
        RECT 65.870 150.830 66.130 151.150 ;
        RECT 66.790 150.830 67.050 151.150 ;
        RECT 55.750 148.790 56.010 149.110 ;
        RECT 56.730 148.090 56.870 150.830 ;
        RECT 64.490 149.810 64.750 150.130 ;
        RECT 64.550 148.430 64.690 149.810 ;
        RECT 65.930 149.110 66.070 150.830 ;
        RECT 65.870 148.790 66.130 149.110 ;
        RECT 64.490 148.110 64.750 148.430 ;
        RECT 66.850 148.090 66.990 150.830 ;
        RECT 67.710 148.450 67.970 148.770 ;
        RECT 67.770 148.090 67.910 148.450 ;
        RECT 72.830 148.430 72.970 158.310 ;
        RECT 73.690 153.270 73.950 153.530 ;
        RECT 73.290 153.210 73.950 153.270 ;
        RECT 73.290 153.130 73.890 153.210 ;
        RECT 73.290 151.150 73.430 153.130 ;
        RECT 74.210 151.830 74.350 172.250 ;
        RECT 74.610 169.870 74.870 170.190 ;
        RECT 74.670 165.430 74.810 169.870 ;
        RECT 75.130 167.810 75.270 177.010 ;
        RECT 76.050 172.570 76.190 180.750 ;
        RECT 76.510 180.730 76.650 180.895 ;
        RECT 76.450 180.410 76.710 180.730 ;
        RECT 76.970 179.030 77.110 182.450 ;
        RECT 76.910 178.710 77.170 179.030 ;
        RECT 76.910 174.290 77.170 174.610 ;
        RECT 75.990 172.250 76.250 172.570 ;
        RECT 76.050 169.850 76.190 172.250 ;
        RECT 76.970 172.230 77.110 174.290 ;
        RECT 77.430 173.590 77.570 189.250 ;
        RECT 78.290 181.430 78.550 181.750 ;
        RECT 77.820 178.855 78.100 179.225 ;
        RECT 77.830 178.710 78.090 178.855 ;
        RECT 78.350 178.690 78.490 181.430 ;
        RECT 79.270 181.070 79.410 191.095 ;
        RECT 80.650 190.930 80.790 194.350 ;
        RECT 81.050 191.970 81.310 192.290 ;
        RECT 80.590 190.610 80.850 190.930 ;
        RECT 81.110 185.490 81.250 191.970 ;
        RECT 81.570 189.910 81.710 194.350 ;
        RECT 88.870 194.010 89.130 194.330 ;
        RECT 85.650 193.330 85.910 193.650 ;
        RECT 85.710 191.610 85.850 193.330 ;
        RECT 85.650 191.290 85.910 191.610 ;
        RECT 86.110 191.290 86.370 191.610 ;
        RECT 81.510 189.590 81.770 189.910 ;
        RECT 85.650 188.570 85.910 188.890 ;
        RECT 85.190 187.890 85.450 188.210 ;
        RECT 80.130 185.170 80.390 185.490 ;
        RECT 81.050 185.170 81.310 185.490 ;
        RECT 79.670 181.090 79.930 181.410 ;
        RECT 79.210 180.750 79.470 181.070 ;
        RECT 78.290 178.370 78.550 178.690 ;
        RECT 78.350 175.290 78.490 178.370 ;
        RECT 79.270 177.330 79.410 180.750 ;
        RECT 79.730 178.350 79.870 181.090 ;
        RECT 80.190 181.070 80.330 185.170 ;
        RECT 81.970 183.470 82.230 183.790 ;
        RECT 82.030 181.750 82.170 183.470 ;
        RECT 81.970 181.430 82.230 181.750 ;
        RECT 80.130 180.750 80.390 181.070 ;
        RECT 82.890 180.410 83.150 180.730 ;
        RECT 82.950 178.690 83.090 180.410 ;
        RECT 83.810 179.730 84.070 180.050 ;
        RECT 83.870 179.030 84.010 179.730 ;
        RECT 83.810 178.710 84.070 179.030 ;
        RECT 82.890 178.370 83.150 178.690 ;
        RECT 79.670 178.030 79.930 178.350 ;
        RECT 84.730 178.030 84.990 178.350 ;
        RECT 79.210 177.010 79.470 177.330 ;
        RECT 78.290 174.970 78.550 175.290 ;
        RECT 77.370 173.270 77.630 173.590 ;
        RECT 78.290 172.590 78.550 172.910 ;
        RECT 76.910 171.910 77.170 172.230 ;
        RECT 77.830 171.570 78.090 171.890 ;
        RECT 76.910 170.550 77.170 170.870 ;
        RECT 75.990 169.530 76.250 169.850 ;
        RECT 75.520 167.975 75.800 168.345 ;
        RECT 75.530 167.830 75.790 167.975 ;
        RECT 75.070 167.490 75.330 167.810 ;
        RECT 76.050 167.130 76.190 169.530 ;
        RECT 76.970 168.150 77.110 170.550 ;
        RECT 76.910 167.830 77.170 168.150 ;
        RECT 77.890 167.470 78.030 171.570 ;
        RECT 77.830 167.150 78.090 167.470 ;
        RECT 75.990 166.810 76.250 167.130 ;
        RECT 78.350 165.430 78.490 172.590 ;
        RECT 79.730 167.470 79.870 178.030 ;
        RECT 80.130 177.690 80.390 178.010 ;
        RECT 80.190 176.310 80.330 177.690 ;
        RECT 84.270 177.350 84.530 177.670 ;
        RECT 83.810 177.010 84.070 177.330 ;
        RECT 80.130 175.990 80.390 176.310 ;
        RECT 80.190 173.590 80.330 175.990 ;
        RECT 81.970 174.630 82.230 174.950 ;
        RECT 82.030 173.590 82.170 174.630 ;
        RECT 80.130 173.270 80.390 173.590 ;
        RECT 81.970 173.270 82.230 173.590 ;
        RECT 83.870 170.190 84.010 177.010 ;
        RECT 84.330 172.570 84.470 177.350 ;
        RECT 84.270 172.250 84.530 172.570 ;
        RECT 83.810 169.870 84.070 170.190 ;
        RECT 80.130 169.530 80.390 169.850 ;
        RECT 80.590 169.530 80.850 169.850 ;
        RECT 80.190 168.150 80.330 169.530 ;
        RECT 80.130 167.830 80.390 168.150 ;
        RECT 79.670 167.150 79.930 167.470 ;
        RECT 74.610 165.110 74.870 165.430 ;
        RECT 78.290 165.110 78.550 165.430 ;
        RECT 80.650 164.070 80.790 169.530 ;
        RECT 83.870 165.430 84.010 169.870 ;
        RECT 83.810 165.110 84.070 165.430 ;
        RECT 80.590 163.750 80.850 164.070 ;
        RECT 80.650 161.010 80.790 163.750 ;
        RECT 81.510 162.390 81.770 162.710 ;
        RECT 80.590 160.690 80.850 161.010 ;
        RECT 75.990 158.990 76.250 159.310 ;
        RECT 74.610 156.270 74.870 156.590 ;
        RECT 74.670 154.550 74.810 156.270 ;
        RECT 76.050 156.250 76.190 158.990 ;
        RECT 75.990 155.930 76.250 156.250 ;
        RECT 74.610 154.230 74.870 154.550 ;
        RECT 76.050 153.870 76.190 155.930 ;
        RECT 75.990 153.550 76.250 153.870 ;
        RECT 75.990 152.870 76.250 153.190 ;
        RECT 74.610 152.530 74.870 152.850 ;
        RECT 74.670 151.830 74.810 152.530 ;
        RECT 74.150 151.510 74.410 151.830 ;
        RECT 74.610 151.510 74.870 151.830 ;
        RECT 74.670 151.150 74.810 151.510 ;
        RECT 73.230 150.830 73.490 151.150 ;
        RECT 74.610 150.830 74.870 151.150 ;
        RECT 68.630 148.110 68.890 148.430 ;
        RECT 72.770 148.110 73.030 148.430 ;
        RECT 56.670 147.770 56.930 148.090 ;
        RECT 66.790 147.770 67.050 148.090 ;
        RECT 67.710 147.770 67.970 148.090 ;
        RECT 54.370 147.090 54.630 147.410 ;
        RECT 55.750 147.090 56.010 147.410 ;
        RECT 54.430 145.710 54.570 147.090 ;
        RECT 54.830 145.730 55.090 146.050 ;
        RECT 55.290 145.730 55.550 146.050 ;
        RECT 54.370 145.390 54.630 145.710 ;
        RECT 53.910 144.370 54.170 144.690 ;
        RECT 53.450 142.670 53.710 142.990 ;
        RECT 54.370 141.880 54.630 141.970 ;
        RECT 54.890 141.880 55.030 145.730 ;
        RECT 55.350 142.650 55.490 145.730 ;
        RECT 55.810 144.690 55.950 147.090 ;
        RECT 66.850 145.710 66.990 147.770 ;
        RECT 67.770 146.470 67.910 147.770 ;
        RECT 67.770 146.330 68.370 146.470 ;
        RECT 58.050 145.390 58.310 145.710 ;
        RECT 66.790 145.620 67.050 145.710 ;
        RECT 66.790 145.480 67.910 145.620 ;
        RECT 66.790 145.390 67.050 145.480 ;
        RECT 55.750 144.370 56.010 144.690 ;
        RECT 55.290 142.330 55.550 142.650 ;
        RECT 54.370 141.740 55.030 141.880 ;
        RECT 54.370 141.650 54.630 141.740 ;
        RECT 54.430 139.250 54.570 141.650 ;
        RECT 54.370 138.930 54.630 139.250 ;
        RECT 52.990 137.230 53.250 137.550 ;
        RECT 54.430 137.210 54.570 138.930 ;
        RECT 55.350 137.550 55.490 142.330 ;
        RECT 55.810 142.310 55.950 144.370 ;
        RECT 58.110 143.670 58.250 145.390 ;
        RECT 67.250 144.370 67.510 144.690 ;
        RECT 58.050 143.350 58.310 143.670 ;
        RECT 55.750 141.990 56.010 142.310 ;
        RECT 62.650 139.610 62.910 139.930 ;
        RECT 62.710 137.550 62.850 139.610 ;
        RECT 55.290 137.230 55.550 137.550 ;
        RECT 62.650 137.230 62.910 137.550 ;
        RECT 54.370 136.890 54.630 137.210 ;
        RECT 52.130 135.280 52.730 135.420 ;
        RECT 51.610 134.850 51.870 135.170 ;
        RECT 52.070 134.510 52.330 134.830 ;
        RECT 52.130 132.790 52.270 134.510 ;
        RECT 52.590 133.810 52.730 135.280 ;
        RECT 62.710 134.830 62.850 137.230 ;
        RECT 62.650 134.510 62.910 134.830 ;
        RECT 66.790 134.510 67.050 134.830 ;
        RECT 52.530 133.490 52.790 133.810 ;
        RECT 52.070 132.470 52.330 132.790 ;
        RECT 52.590 132.450 52.730 133.490 ;
        RECT 52.530 132.130 52.790 132.450 ;
        RECT 51.150 131.110 51.410 131.430 ;
        RECT 62.710 129.730 62.850 134.510 ;
        RECT 66.850 132.790 66.990 134.510 ;
        RECT 66.790 132.470 67.050 132.790 ;
        RECT 50.230 129.410 50.490 129.730 ;
        RECT 62.650 129.410 62.910 129.730 ;
        RECT 56.210 129.070 56.470 129.390 ;
        RECT 56.270 125.650 56.410 129.070 ;
        RECT 62.710 126.330 62.850 129.410 ;
        RECT 64.030 129.070 64.290 129.390 ;
        RECT 64.090 126.670 64.230 129.070 ;
        RECT 64.030 126.350 64.290 126.670 ;
        RECT 62.650 126.010 62.910 126.330 ;
        RECT 56.210 125.330 56.470 125.650 ;
        RECT 57.590 125.330 57.850 125.650 ;
        RECT 55.750 123.290 56.010 123.610 ;
        RECT 43.790 121.250 44.050 121.570 ;
        RECT 47.470 121.250 47.730 121.570 ;
        RECT 41.950 120.570 42.210 120.890 ;
        RECT 41.490 119.890 41.750 120.210 ;
        RECT 42.010 118.170 42.150 120.570 ;
        RECT 41.950 117.850 42.210 118.170 ;
        RECT 41.950 117.170 42.210 117.490 ;
        RECT 40.570 115.130 40.830 115.450 ;
        RECT 41.030 115.130 41.290 115.450 ;
        RECT 42.010 115.360 42.150 117.170 ;
        RECT 43.850 115.450 43.990 121.250 ;
        RECT 54.370 120.570 54.630 120.890 ;
        RECT 52.990 119.890 53.250 120.210 ;
        RECT 53.050 119.190 53.190 119.890 ;
        RECT 51.610 118.870 51.870 119.190 ;
        RECT 52.990 118.870 53.250 119.190 ;
        RECT 44.710 118.530 44.970 118.850 ;
        RECT 44.250 117.170 44.510 117.490 ;
        RECT 42.410 115.360 42.670 115.450 ;
        RECT 42.010 115.220 42.670 115.360 ;
        RECT 42.410 115.130 42.670 115.220 ;
        RECT 43.790 115.130 44.050 115.450 ;
        RECT 40.630 108.310 40.770 115.130 ;
        RECT 41.090 113.750 41.230 115.130 ;
        RECT 43.330 114.450 43.590 114.770 ;
        RECT 41.030 113.430 41.290 113.750 ;
        RECT 43.390 113.070 43.530 114.450 ;
        RECT 44.310 113.070 44.450 117.170 ;
        RECT 44.770 116.470 44.910 118.530 ;
        RECT 47.930 117.850 48.190 118.170 ;
        RECT 44.710 116.150 44.970 116.470 ;
        RECT 44.770 113.750 44.910 116.150 ;
        RECT 47.990 114.770 48.130 117.850 ;
        RECT 51.670 114.770 51.810 118.870 ;
        RECT 54.430 118.510 54.570 120.570 ;
        RECT 54.370 118.190 54.630 118.510 ;
        RECT 55.810 117.830 55.950 123.290 ;
        RECT 56.270 118.850 56.410 125.330 ;
        RECT 57.650 121.910 57.790 125.330 ;
        RECT 62.710 123.950 62.850 126.010 ;
        RECT 63.110 125.670 63.370 125.990 ;
        RECT 58.970 123.630 59.230 123.950 ;
        RECT 62.650 123.630 62.910 123.950 ;
        RECT 57.590 121.590 57.850 121.910 ;
        RECT 59.030 120.210 59.170 123.630 ;
        RECT 63.170 122.930 63.310 125.670 ;
        RECT 63.110 122.610 63.370 122.930 ;
        RECT 60.350 120.230 60.610 120.550 ;
        RECT 58.970 119.890 59.230 120.210 ;
        RECT 56.210 118.530 56.470 118.850 ;
        RECT 59.030 117.830 59.170 119.890 ;
        RECT 60.410 118.170 60.550 120.230 ;
        RECT 60.350 117.850 60.610 118.170 ;
        RECT 55.750 117.510 56.010 117.830 ;
        RECT 58.970 117.510 59.230 117.830 ;
        RECT 59.890 115.470 60.150 115.790 ;
        RECT 53.450 114.790 53.710 115.110 ;
        RECT 47.930 114.450 48.190 114.770 ;
        RECT 51.610 114.450 51.870 114.770 ;
        RECT 47.990 113.750 48.130 114.450 ;
        RECT 53.510 113.750 53.650 114.790 ;
        RECT 44.710 113.430 44.970 113.750 ;
        RECT 47.930 113.430 48.190 113.750 ;
        RECT 53.450 113.430 53.710 113.750 ;
        RECT 59.950 113.070 60.090 115.470 ;
        RECT 60.410 115.450 60.550 117.850 ;
        RECT 62.640 116.975 62.920 117.345 ;
        RECT 62.710 115.790 62.850 116.975 ;
        RECT 63.170 116.130 63.310 122.610 ;
        RECT 64.090 120.210 64.230 126.350 ;
        RECT 65.410 120.570 65.670 120.890 ;
        RECT 64.030 119.890 64.290 120.210 ;
        RECT 64.490 119.890 64.750 120.210 ;
        RECT 64.090 118.170 64.230 119.890 ;
        RECT 64.550 119.190 64.690 119.890 ;
        RECT 65.470 119.190 65.610 120.570 ;
        RECT 64.490 118.870 64.750 119.190 ;
        RECT 65.410 118.870 65.670 119.190 ;
        RECT 64.030 117.850 64.290 118.170 ;
        RECT 63.110 115.810 63.370 116.130 ;
        RECT 62.650 115.470 62.910 115.790 ;
        RECT 64.090 115.450 64.230 117.850 ;
        RECT 65.470 116.470 65.610 118.870 ;
        RECT 65.870 118.190 66.130 118.510 ;
        RECT 65.410 116.150 65.670 116.470 ;
        RECT 60.350 115.130 60.610 115.450 ;
        RECT 64.030 115.130 64.290 115.450 ;
        RECT 43.330 112.750 43.590 113.070 ;
        RECT 44.250 112.750 44.510 113.070 ;
        RECT 47.010 112.750 47.270 113.070 ;
        RECT 47.470 112.750 47.730 113.070 ;
        RECT 48.390 112.750 48.650 113.070 ;
        RECT 50.230 112.750 50.490 113.070 ;
        RECT 59.890 112.750 60.150 113.070 ;
        RECT 47.070 111.030 47.210 112.750 ;
        RECT 47.530 112.390 47.670 112.750 ;
        RECT 47.470 112.070 47.730 112.390 ;
        RECT 47.010 110.710 47.270 111.030 ;
        RECT 46.550 109.010 46.810 109.330 ;
        RECT 40.110 107.990 40.370 108.310 ;
        RECT 40.570 107.990 40.830 108.310 ;
        RECT 40.170 107.630 40.310 107.990 ;
        RECT 38.270 107.310 38.530 107.630 ;
        RECT 40.110 107.310 40.370 107.630 ;
        RECT 38.330 104.570 38.470 107.310 ;
        RECT 38.270 104.250 38.530 104.570 ;
        RECT 38.330 102.870 38.470 104.250 ;
        RECT 40.170 103.890 40.310 107.310 ;
        RECT 40.630 105.250 40.770 107.990 ;
        RECT 46.610 107.630 46.750 109.010 ;
        RECT 47.530 107.970 47.670 112.070 ;
        RECT 48.450 109.330 48.590 112.750 ;
        RECT 50.290 112.050 50.430 112.750 ;
        RECT 50.230 111.730 50.490 112.050 ;
        RECT 48.390 109.010 48.650 109.330 ;
        RECT 48.450 108.310 48.590 109.010 ;
        RECT 48.390 107.990 48.650 108.310 ;
        RECT 47.470 107.650 47.730 107.970 ;
        RECT 49.310 107.650 49.570 107.970 ;
        RECT 45.170 107.310 45.430 107.630 ;
        RECT 46.550 107.310 46.810 107.630 ;
        RECT 40.570 104.930 40.830 105.250 ;
        RECT 40.110 103.570 40.370 103.890 ;
        RECT 40.630 102.950 40.770 104.930 ;
        RECT 41.030 103.570 41.290 103.890 ;
        RECT 36.890 102.550 37.150 102.870 ;
        RECT 38.270 102.550 38.530 102.870 ;
        RECT 40.170 102.810 40.770 102.950 ;
        RECT 40.170 102.530 40.310 102.810 ;
        RECT 40.110 102.210 40.370 102.530 ;
        RECT 41.090 101.170 41.230 103.570 ;
        RECT 45.230 102.530 45.370 107.310 ;
        RECT 46.610 104.230 46.750 107.310 ;
        RECT 46.550 103.910 46.810 104.230 ;
        RECT 47.530 102.530 47.670 107.650 ;
        RECT 49.370 106.610 49.510 107.650 ;
        RECT 50.290 107.630 50.430 111.730 ;
        RECT 51.610 109.690 51.870 110.010 ;
        RECT 49.770 107.310 50.030 107.630 ;
        RECT 50.230 107.310 50.490 107.630 ;
        RECT 49.830 106.950 49.970 107.310 ;
        RECT 49.770 106.630 50.030 106.950 ;
        RECT 49.310 106.290 49.570 106.610 ;
        RECT 49.370 105.250 49.510 106.290 ;
        RECT 49.310 104.930 49.570 105.250 ;
        RECT 45.170 102.210 45.430 102.530 ;
        RECT 47.470 102.210 47.730 102.530 ;
        RECT 47.530 101.510 47.670 102.210 ;
        RECT 47.470 101.190 47.730 101.510 ;
        RECT 29.990 100.850 30.250 101.170 ;
        RECT 36.430 100.850 36.690 101.170 ;
        RECT 41.030 100.850 41.290 101.170 ;
        RECT 28.880 100.315 30.420 100.685 ;
        RECT 21.310 100.150 21.910 100.230 ;
        RECT 21.310 100.090 21.970 100.150 ;
        RECT 21.710 99.830 21.970 100.090 ;
        RECT 49.370 99.130 49.510 104.930 ;
        RECT 49.830 100.150 49.970 106.630 ;
        RECT 49.770 99.830 50.030 100.150 ;
        RECT 50.290 99.470 50.430 107.310 ;
        RECT 50.690 105.270 50.950 105.590 ;
        RECT 50.750 102.870 50.890 105.270 ;
        RECT 51.670 104.910 51.810 109.690 ;
        RECT 52.070 109.350 52.330 109.670 ;
        RECT 52.130 108.310 52.270 109.350 ;
        RECT 52.070 107.990 52.330 108.310 ;
        RECT 52.530 107.310 52.790 107.630 ;
        RECT 54.370 107.310 54.630 107.630 ;
        RECT 52.590 105.590 52.730 107.310 ;
        RECT 52.530 105.270 52.790 105.590 ;
        RECT 51.610 104.590 51.870 104.910 ;
        RECT 51.150 103.570 51.410 103.890 ;
        RECT 50.690 102.550 50.950 102.870 ;
        RECT 51.210 102.190 51.350 103.570 ;
        RECT 51.670 102.530 51.810 104.590 ;
        RECT 54.430 104.230 54.570 107.310 ;
        RECT 55.290 106.290 55.550 106.610 ;
        RECT 55.350 104.230 55.490 106.290 ;
        RECT 54.370 103.910 54.630 104.230 ;
        RECT 55.290 103.910 55.550 104.230 ;
        RECT 51.610 102.210 51.870 102.530 ;
        RECT 51.150 101.870 51.410 102.190 ;
        RECT 50.230 99.150 50.490 99.470 ;
        RECT 18.950 98.810 19.210 99.130 ;
        RECT 49.310 98.810 49.570 99.130 ;
        RECT 32.180 97.595 33.720 97.965 ;
        RECT 28.880 94.875 30.420 95.245 ;
        RECT 32.180 92.155 33.720 92.525 ;
        RECT 28.880 89.435 30.420 89.805 ;
        RECT 59.950 89.270 60.090 112.750 ;
        RECT 60.410 109.670 60.550 115.130 ;
        RECT 62.650 114.790 62.910 115.110 ;
        RECT 62.190 112.980 62.450 113.070 ;
        RECT 62.710 112.980 62.850 114.790 ;
        RECT 64.950 114.450 65.210 114.770 ;
        RECT 62.190 112.840 62.850 112.980 ;
        RECT 62.190 112.750 62.450 112.840 ;
        RECT 64.490 112.070 64.750 112.390 ;
        RECT 63.110 110.370 63.370 110.690 ;
        RECT 62.650 110.030 62.910 110.350 ;
        RECT 60.350 109.350 60.610 109.670 ;
        RECT 60.410 104.570 60.550 109.350 ;
        RECT 62.710 108.310 62.850 110.030 ;
        RECT 62.650 107.990 62.910 108.310 ;
        RECT 62.650 107.540 62.910 107.630 ;
        RECT 63.170 107.540 63.310 110.370 ;
        RECT 64.550 110.010 64.690 112.070 ;
        RECT 65.010 111.030 65.150 114.450 ;
        RECT 65.470 113.070 65.610 116.150 ;
        RECT 65.930 113.750 66.070 118.190 ;
        RECT 66.790 117.170 67.050 117.490 ;
        RECT 66.850 116.470 66.990 117.170 ;
        RECT 66.790 116.150 67.050 116.470 ;
        RECT 66.330 115.470 66.590 115.790 ;
        RECT 65.870 113.430 66.130 113.750 ;
        RECT 66.390 113.070 66.530 115.470 ;
        RECT 65.410 112.750 65.670 113.070 ;
        RECT 66.330 112.750 66.590 113.070 ;
        RECT 67.310 112.730 67.450 144.370 ;
        RECT 67.770 113.320 67.910 145.480 ;
        RECT 68.230 144.690 68.370 146.330 ;
        RECT 68.690 146.050 68.830 148.110 ;
        RECT 70.930 147.430 71.190 147.750 ;
        RECT 69.550 147.090 69.810 147.410 ;
        RECT 68.630 145.730 68.890 146.050 ;
        RECT 68.170 144.370 68.430 144.690 ;
        RECT 69.610 144.430 69.750 147.090 ;
        RECT 70.990 145.370 71.130 147.430 ;
        RECT 73.290 145.710 73.430 150.830 ;
        RECT 71.850 145.390 72.110 145.710 ;
        RECT 73.230 145.390 73.490 145.710 ;
        RECT 70.930 145.050 71.190 145.370 ;
        RECT 70.010 144.430 70.270 144.690 ;
        RECT 69.610 144.370 70.270 144.430 ;
        RECT 69.610 144.290 70.210 144.370 ;
        RECT 68.170 141.650 68.430 141.970 ;
        RECT 68.230 131.430 68.370 141.650 ;
        RECT 68.170 131.110 68.430 131.430 ;
        RECT 69.610 130.070 69.750 144.290 ;
        RECT 70.010 142.330 70.270 142.650 ;
        RECT 70.070 135.510 70.210 142.330 ;
        RECT 70.010 135.190 70.270 135.510 ;
        RECT 70.930 131.450 71.190 131.770 ;
        RECT 70.010 131.110 70.270 131.430 ;
        RECT 69.550 129.750 69.810 130.070 ;
        RECT 70.070 129.390 70.210 131.110 ;
        RECT 70.990 129.390 71.130 131.450 ;
        RECT 69.090 129.070 69.350 129.390 ;
        RECT 70.010 129.070 70.270 129.390 ;
        RECT 70.930 129.070 71.190 129.390 ;
        RECT 68.170 128.390 68.430 128.710 ;
        RECT 68.230 118.850 68.370 128.390 ;
        RECT 68.630 128.050 68.890 128.370 ;
        RECT 68.690 124.290 68.830 128.050 ;
        RECT 69.150 127.350 69.290 129.070 ;
        RECT 69.090 127.030 69.350 127.350 ;
        RECT 70.070 125.990 70.210 129.070 ;
        RECT 70.010 125.670 70.270 125.990 ;
        RECT 68.630 123.970 68.890 124.290 ;
        RECT 68.630 122.610 68.890 122.930 ;
        RECT 68.690 121.230 68.830 122.610 ;
        RECT 68.630 120.910 68.890 121.230 ;
        RECT 70.070 120.210 70.210 125.670 ;
        RECT 69.550 119.890 69.810 120.210 ;
        RECT 70.010 119.890 70.270 120.210 ;
        RECT 70.470 119.890 70.730 120.210 ;
        RECT 68.170 118.530 68.430 118.850 ;
        RECT 68.230 115.110 68.370 118.530 ;
        RECT 68.630 117.345 68.890 117.490 ;
        RECT 68.620 116.975 68.900 117.345 ;
        RECT 69.610 115.110 69.750 119.890 ;
        RECT 70.010 117.170 70.270 117.490 ;
        RECT 70.070 115.190 70.210 117.170 ;
        RECT 70.530 115.790 70.670 119.890 ;
        RECT 71.390 118.870 71.650 119.190 ;
        RECT 71.450 117.490 71.590 118.870 ;
        RECT 71.390 117.170 71.650 117.490 ;
        RECT 70.470 115.470 70.730 115.790 ;
        RECT 70.070 115.110 70.670 115.190 ;
        RECT 70.930 115.130 71.190 115.450 ;
        RECT 68.170 114.790 68.430 115.110 ;
        RECT 69.550 114.790 69.810 115.110 ;
        RECT 70.070 115.050 70.730 115.110 ;
        RECT 70.470 114.790 70.730 115.050 ;
        RECT 70.010 114.450 70.270 114.770 ;
        RECT 70.070 113.410 70.210 114.450 ;
        RECT 67.770 113.180 68.370 113.320 ;
        RECT 68.230 112.730 68.370 113.180 ;
        RECT 70.010 113.090 70.270 113.410 ;
        RECT 65.860 112.215 66.140 112.585 ;
        RECT 67.250 112.410 67.510 112.730 ;
        RECT 68.170 112.410 68.430 112.730 ;
        RECT 70.010 112.585 70.270 112.730 ;
        RECT 65.870 112.070 66.130 112.215 ;
        RECT 64.950 110.710 65.210 111.030 ;
        RECT 64.490 109.690 64.750 110.010 ;
        RECT 67.310 109.670 67.450 112.410 ;
        RECT 67.710 111.730 67.970 112.050 ;
        RECT 67.770 111.030 67.910 111.730 ;
        RECT 67.710 110.710 67.970 111.030 ;
        RECT 67.250 109.350 67.510 109.670 ;
        RECT 64.490 109.010 64.750 109.330 ;
        RECT 62.650 107.400 63.310 107.540 ;
        RECT 62.650 107.310 62.910 107.400 ;
        RECT 64.550 107.290 64.690 109.010 ;
        RECT 68.230 107.970 68.370 112.410 ;
        RECT 70.000 112.215 70.280 112.585 ;
        RECT 70.990 111.030 71.130 115.130 ;
        RECT 71.450 113.070 71.590 117.170 ;
        RECT 71.390 112.750 71.650 113.070 ;
        RECT 70.930 110.710 71.190 111.030 ;
        RECT 68.170 107.650 68.430 107.970 ;
        RECT 64.490 106.970 64.750 107.290 ;
        RECT 67.710 106.970 67.970 107.290 ;
        RECT 61.730 106.290 61.990 106.610 ;
        RECT 61.790 104.570 61.930 106.290 ;
        RECT 60.350 104.250 60.610 104.570 ;
        RECT 61.730 104.250 61.990 104.570 ;
        RECT 67.770 103.890 67.910 106.970 ;
        RECT 67.710 103.570 67.970 103.890 ;
        RECT 59.890 88.950 60.150 89.270 ;
        RECT 67.770 88.250 67.910 103.570 ;
        RECT 70.470 98.810 70.730 99.130 ;
        RECT 70.530 96.410 70.670 98.810 ;
        RECT 71.910 98.450 72.050 145.390 ;
        RECT 74.670 142.990 74.810 150.830 ;
        RECT 75.530 147.090 75.790 147.410 ;
        RECT 74.610 142.670 74.870 142.990 ;
        RECT 75.590 142.650 75.730 147.090 ;
        RECT 76.050 145.370 76.190 152.870 ;
        RECT 77.830 150.830 78.090 151.150 ;
        RECT 77.370 149.810 77.630 150.130 ;
        RECT 77.430 148.430 77.570 149.810 ;
        RECT 77.370 148.110 77.630 148.430 ;
        RECT 75.990 145.050 76.250 145.370 ;
        RECT 77.890 143.670 78.030 150.830 ;
        RECT 81.570 146.390 81.710 162.390 ;
        RECT 83.870 159.310 84.010 165.110 ;
        RECT 83.810 158.990 84.070 159.310 ;
        RECT 84.270 158.990 84.530 159.310 ;
        RECT 84.330 155.570 84.470 158.990 ;
        RECT 84.270 155.250 84.530 155.570 ;
        RECT 84.330 153.870 84.470 155.250 ;
        RECT 84.790 153.870 84.930 178.030 ;
        RECT 85.250 172.570 85.390 187.890 ;
        RECT 85.710 186.170 85.850 188.570 ;
        RECT 85.650 185.850 85.910 186.170 ;
        RECT 85.190 172.250 85.450 172.570 ;
        RECT 85.710 171.630 85.850 185.850 ;
        RECT 86.170 183.790 86.310 191.290 ;
        RECT 87.950 190.610 88.210 190.930 ;
        RECT 88.010 189.230 88.150 190.610 ;
        RECT 88.930 189.910 89.070 194.010 ;
        RECT 90.310 191.950 90.450 194.690 ;
        RECT 90.250 191.630 90.510 191.950 ;
        RECT 90.770 191.610 90.910 196.050 ;
        RECT 91.170 193.330 91.430 193.650 ;
        RECT 90.710 191.290 90.970 191.610 ;
        RECT 88.870 189.590 89.130 189.910 ;
        RECT 87.950 188.910 88.210 189.230 ;
        RECT 88.410 188.910 88.670 189.230 ;
        RECT 88.470 186.510 88.610 188.910 ;
        RECT 91.230 188.890 91.370 193.330 ;
        RECT 91.690 192.630 91.830 196.050 ;
        RECT 91.630 192.310 91.890 192.630 ;
        RECT 91.170 188.570 91.430 188.890 ;
        RECT 91.230 186.510 91.370 188.570 ;
        RECT 88.410 186.190 88.670 186.510 ;
        RECT 91.170 186.190 91.430 186.510 ;
        RECT 91.690 185.830 91.830 192.310 ;
        RECT 93.010 190.610 93.270 190.930 ;
        RECT 93.070 188.890 93.210 190.610 ;
        RECT 93.930 189.310 94.190 189.570 ;
        RECT 93.930 189.250 94.590 189.310 ;
        RECT 93.990 189.170 94.590 189.250 ;
        RECT 93.010 188.570 93.270 188.890 ;
        RECT 93.070 186.170 93.210 188.570 ;
        RECT 94.450 186.850 94.590 189.170 ;
        RECT 95.770 188.570 96.030 188.890 ;
        RECT 94.390 186.530 94.650 186.850 ;
        RECT 93.010 185.850 93.270 186.170 ;
        RECT 93.930 185.850 94.190 186.170 ;
        RECT 91.630 185.510 91.890 185.830 ;
        RECT 93.990 185.490 94.130 185.850 ;
        RECT 93.930 185.170 94.190 185.490 ;
        RECT 86.110 183.470 86.370 183.790 ;
        RECT 86.170 175.630 86.310 183.470 ;
        RECT 94.450 180.730 94.590 186.530 ;
        RECT 95.830 186.170 95.970 188.570 ;
        RECT 96.290 188.550 96.430 196.820 ;
        RECT 98.530 196.730 98.790 197.050 ;
        RECT 101.290 196.730 101.550 197.050 ;
        RECT 97.150 196.050 97.410 196.370 ;
        RECT 96.690 193.330 96.950 193.650 ;
        RECT 96.750 191.610 96.890 193.330 ;
        RECT 96.690 191.290 96.950 191.610 ;
        RECT 96.230 188.230 96.490 188.550 ;
        RECT 97.210 188.210 97.350 196.050 ;
        RECT 98.590 195.010 98.730 196.730 ;
        RECT 99.450 196.390 99.710 196.710 ;
        RECT 98.530 194.690 98.790 195.010 ;
        RECT 97.610 194.580 97.870 194.670 ;
        RECT 97.610 194.440 98.270 194.580 ;
        RECT 97.610 194.350 97.870 194.440 ;
        RECT 97.610 190.610 97.870 190.930 ;
        RECT 97.670 189.570 97.810 190.610 ;
        RECT 98.130 189.910 98.270 194.440 ;
        RECT 98.070 189.590 98.330 189.910 ;
        RECT 97.610 189.250 97.870 189.570 ;
        RECT 97.150 187.890 97.410 188.210 ;
        RECT 97.210 187.190 97.350 187.890 ;
        RECT 97.150 186.870 97.410 187.190 ;
        RECT 97.670 186.490 97.810 189.250 ;
        RECT 99.510 189.230 99.650 196.390 ;
        RECT 101.350 194.580 101.490 196.730 ;
        RECT 101.350 194.440 102.870 194.580 ;
        RECT 101.290 193.330 101.550 193.650 ;
        RECT 100.830 190.950 101.090 191.270 ;
        RECT 100.890 189.570 101.030 190.950 ;
        RECT 100.830 189.250 101.090 189.570 ;
        RECT 101.350 189.230 101.490 193.330 ;
        RECT 102.730 191.610 102.870 194.440 ;
        RECT 103.590 194.350 103.850 194.670 ;
        RECT 103.650 192.630 103.790 194.350 ;
        RECT 103.590 192.310 103.850 192.630 ;
        RECT 103.590 191.630 103.850 191.950 ;
        RECT 102.670 191.290 102.930 191.610 ;
        RECT 102.730 189.230 102.870 191.290 ;
        RECT 103.130 190.610 103.390 190.930 ;
        RECT 99.450 188.910 99.710 189.230 ;
        RECT 101.290 188.910 101.550 189.230 ;
        RECT 102.670 188.910 102.930 189.230 ;
        RECT 102.730 187.190 102.870 188.910 ;
        RECT 102.670 186.870 102.930 187.190 ;
        RECT 98.070 186.490 98.330 186.510 ;
        RECT 97.670 186.350 98.330 186.490 ;
        RECT 98.070 186.190 98.330 186.350 ;
        RECT 103.190 186.170 103.330 190.610 ;
        RECT 103.650 189.230 103.790 191.630 ;
        RECT 103.590 188.910 103.850 189.230 ;
        RECT 104.110 189.140 104.250 197.070 ;
        RECT 106.350 196.730 106.610 197.050 ;
        RECT 105.890 196.390 106.150 196.710 ;
        RECT 104.970 196.050 105.230 196.370 ;
        RECT 105.030 191.610 105.170 196.050 ;
        RECT 105.950 192.630 106.090 196.390 ;
        RECT 105.890 192.310 106.150 192.630 ;
        RECT 104.970 191.290 105.230 191.610 ;
        RECT 105.950 189.570 106.090 192.310 ;
        RECT 106.410 192.290 106.550 196.730 ;
        RECT 113.250 196.390 113.510 196.710 ;
        RECT 108.650 196.050 108.910 196.370 ;
        RECT 106.350 191.970 106.610 192.290 ;
        RECT 105.890 189.250 106.150 189.570 ;
        RECT 104.510 189.140 104.770 189.230 ;
        RECT 104.110 189.000 104.770 189.140 ;
        RECT 104.510 188.910 104.770 189.000 ;
        RECT 104.970 188.570 105.230 188.890 ;
        RECT 103.590 187.890 103.850 188.210 ;
        RECT 95.770 185.850 96.030 186.170 ;
        RECT 103.130 185.850 103.390 186.170 ;
        RECT 103.190 181.070 103.330 185.850 ;
        RECT 103.650 182.770 103.790 187.890 ;
        RECT 104.510 186.870 104.770 187.190 ;
        RECT 104.570 186.490 104.710 186.870 ;
        RECT 105.030 186.850 105.170 188.570 ;
        RECT 105.430 187.890 105.690 188.210 ;
        RECT 104.970 186.530 105.230 186.850 ;
        RECT 104.110 186.350 104.710 186.490 ;
        RECT 103.590 182.450 103.850 182.770 ;
        RECT 94.850 180.750 95.110 181.070 ;
        RECT 103.130 180.750 103.390 181.070 ;
        RECT 94.390 180.410 94.650 180.730 ;
        RECT 91.170 179.730 91.430 180.050 ;
        RECT 86.110 175.310 86.370 175.630 ;
        RECT 86.170 172.570 86.310 175.310 ;
        RECT 91.230 175.290 91.370 179.730 ;
        RECT 94.910 179.030 95.050 180.750 ;
        RECT 95.310 180.410 95.570 180.730 ;
        RECT 94.850 178.710 95.110 179.030 ;
        RECT 94.390 178.030 94.650 178.350 ;
        RECT 93.470 175.990 93.730 176.310 ;
        RECT 91.170 174.970 91.430 175.290 ;
        RECT 91.170 172.590 91.430 172.910 ;
        RECT 86.110 172.250 86.370 172.570 ;
        RECT 85.250 171.490 85.850 171.630 ;
        RECT 85.250 166.870 85.390 171.490 ;
        RECT 85.650 168.850 85.910 169.170 ;
        RECT 85.710 167.810 85.850 168.850 ;
        RECT 85.650 167.490 85.910 167.810 ;
        RECT 86.170 167.380 86.310 172.250 ;
        RECT 91.230 170.870 91.370 172.590 ;
        RECT 91.170 170.550 91.430 170.870 ;
        RECT 93.530 170.190 93.670 175.990 ;
        RECT 93.930 172.590 94.190 172.910 ;
        RECT 93.470 169.870 93.730 170.190 ;
        RECT 92.090 169.530 92.350 169.850 ;
        RECT 87.950 168.850 88.210 169.170 ;
        RECT 86.570 167.380 86.830 167.470 ;
        RECT 86.170 167.240 86.830 167.380 ;
        RECT 86.570 167.150 86.830 167.240 ;
        RECT 85.250 166.730 85.850 166.870 ;
        RECT 85.190 164.090 85.450 164.410 ;
        RECT 85.250 162.030 85.390 164.090 ;
        RECT 85.190 161.710 85.450 162.030 ;
        RECT 84.270 153.550 84.530 153.870 ;
        RECT 84.730 153.550 84.990 153.870 ;
        RECT 81.970 152.530 82.230 152.850 ;
        RECT 82.030 150.130 82.170 152.530 ;
        RECT 83.810 150.490 84.070 150.810 ;
        RECT 84.790 150.550 84.930 153.550 ;
        RECT 81.970 149.810 82.230 150.130 ;
        RECT 83.870 147.750 84.010 150.490 ;
        RECT 84.330 150.410 84.930 150.550 ;
        RECT 85.710 150.470 85.850 166.730 ;
        RECT 87.490 163.410 87.750 163.730 ;
        RECT 87.550 159.990 87.690 163.410 ;
        RECT 88.010 162.030 88.150 168.850 ;
        RECT 92.150 166.450 92.290 169.530 ;
        RECT 93.470 168.850 93.730 169.170 ;
        RECT 92.090 166.130 92.350 166.450 ;
        RECT 88.410 164.430 88.670 164.750 ;
        RECT 87.950 161.710 88.210 162.030 ;
        RECT 88.470 161.690 88.610 164.430 ;
        RECT 90.710 164.090 90.970 164.410 ;
        RECT 90.770 162.710 90.910 164.090 ;
        RECT 90.710 162.390 90.970 162.710 ;
        RECT 88.410 161.370 88.670 161.690 ;
        RECT 87.490 159.670 87.750 159.990 ;
        RECT 92.150 159.310 92.290 166.130 ;
        RECT 92.550 162.050 92.810 162.370 ;
        RECT 92.610 159.310 92.750 162.050 ;
        RECT 92.090 158.990 92.350 159.310 ;
        RECT 92.550 158.990 92.810 159.310 ;
        RECT 87.030 157.970 87.290 158.290 ;
        RECT 86.570 151.170 86.830 151.490 ;
        RECT 83.810 147.430 84.070 147.750 ;
        RECT 84.330 147.410 84.470 150.410 ;
        RECT 85.650 150.150 85.910 150.470 ;
        RECT 84.730 149.810 84.990 150.130 ;
        RECT 84.790 147.410 84.930 149.810 ;
        RECT 86.110 147.770 86.370 148.090 ;
        RECT 84.270 147.090 84.530 147.410 ;
        RECT 84.730 147.090 84.990 147.410 ;
        RECT 81.510 146.070 81.770 146.390 ;
        RECT 77.830 143.350 78.090 143.670 ;
        RECT 75.530 142.330 75.790 142.650 ;
        RECT 72.770 141.990 73.030 142.310 ;
        RECT 79.210 141.990 79.470 142.310 ;
        RECT 72.310 139.950 72.570 140.270 ;
        RECT 72.370 132.790 72.510 139.950 ;
        RECT 72.830 134.830 72.970 141.990 ;
        RECT 74.150 138.930 74.410 139.250 ;
        RECT 73.230 137.230 73.490 137.550 ;
        RECT 73.290 135.510 73.430 137.230 ;
        RECT 73.230 135.190 73.490 135.510 ;
        RECT 72.770 134.510 73.030 134.830 ;
        RECT 72.310 132.470 72.570 132.790 ;
        RECT 73.290 132.450 73.430 135.190 ;
        RECT 74.210 134.830 74.350 138.930 ;
        RECT 74.610 136.890 74.870 137.210 ;
        RECT 74.150 134.510 74.410 134.830 ;
        RECT 73.690 133.830 73.950 134.150 ;
        RECT 73.230 132.130 73.490 132.450 ;
        RECT 73.750 131.770 73.890 133.830 ;
        RECT 74.210 132.110 74.350 134.510 ;
        RECT 74.150 131.790 74.410 132.110 ;
        RECT 73.690 131.450 73.950 131.770 ;
        RECT 74.670 131.510 74.810 136.890 ;
        RECT 78.750 136.210 79.010 136.530 ;
        RECT 75.990 134.850 76.250 135.170 ;
        RECT 76.050 131.770 76.190 134.850 ;
        RECT 77.370 134.510 77.630 134.830 ;
        RECT 73.750 130.070 73.890 131.450 ;
        RECT 74.210 131.370 74.810 131.510 ;
        RECT 75.990 131.450 76.250 131.770 ;
        RECT 73.690 129.750 73.950 130.070 ;
        RECT 72.310 122.610 72.570 122.930 ;
        RECT 72.370 121.910 72.510 122.610 ;
        RECT 72.310 121.590 72.570 121.910 ;
        RECT 74.210 120.630 74.350 131.370 ;
        RECT 76.450 128.730 76.710 129.050 ;
        RECT 76.510 126.330 76.650 128.730 ;
        RECT 74.610 126.010 74.870 126.330 ;
        RECT 76.450 126.240 76.710 126.330 ;
        RECT 76.050 126.100 76.710 126.240 ;
        RECT 73.750 120.490 74.350 120.630 ;
        RECT 73.750 102.190 73.890 120.490 ;
        RECT 74.150 119.890 74.410 120.210 ;
        RECT 74.210 118.510 74.350 119.890 ;
        RECT 74.150 118.190 74.410 118.510 ;
        RECT 74.210 115.790 74.350 118.190 ;
        RECT 74.670 117.830 74.810 126.010 ;
        RECT 75.070 125.330 75.330 125.650 ;
        RECT 74.610 117.510 74.870 117.830 ;
        RECT 75.130 115.790 75.270 125.330 ;
        RECT 76.050 121.910 76.190 126.100 ;
        RECT 76.450 126.010 76.710 126.100 ;
        RECT 76.450 122.610 76.710 122.930 ;
        RECT 75.990 121.590 76.250 121.910 ;
        RECT 75.990 120.570 76.250 120.890 ;
        RECT 75.530 120.230 75.790 120.550 ;
        RECT 75.590 118.510 75.730 120.230 ;
        RECT 75.530 118.190 75.790 118.510 ;
        RECT 76.050 118.170 76.190 120.570 ;
        RECT 76.510 118.170 76.650 122.610 ;
        RECT 76.910 120.570 77.170 120.890 ;
        RECT 76.970 119.190 77.110 120.570 ;
        RECT 76.910 118.870 77.170 119.190 ;
        RECT 75.990 117.850 76.250 118.170 ;
        RECT 76.450 117.850 76.710 118.170 ;
        RECT 74.150 115.470 74.410 115.790 ;
        RECT 75.070 115.470 75.330 115.790 ;
        RECT 75.130 112.730 75.270 115.470 ;
        RECT 77.430 114.680 77.570 134.510 ;
        RECT 78.810 134.490 78.950 136.210 ;
        RECT 78.750 134.170 79.010 134.490 ;
        RECT 78.750 133.490 79.010 133.810 ;
        RECT 78.810 132.790 78.950 133.490 ;
        RECT 78.750 132.470 79.010 132.790 ;
        RECT 78.810 127.350 78.950 132.470 ;
        RECT 78.750 127.030 79.010 127.350 ;
        RECT 78.290 122.610 78.550 122.930 ;
        RECT 78.350 118.510 78.490 122.610 ;
        RECT 78.750 118.530 79.010 118.850 ;
        RECT 78.290 118.190 78.550 118.510 ;
        RECT 78.810 115.450 78.950 118.530 ;
        RECT 78.750 115.130 79.010 115.450 ;
        RECT 77.430 114.540 78.030 114.680 ;
        RECT 75.070 112.410 75.330 112.730 ;
        RECT 76.910 109.690 77.170 110.010 ;
        RECT 76.970 105.250 77.110 109.690 ;
        RECT 77.370 106.290 77.630 106.610 ;
        RECT 76.910 104.930 77.170 105.250 ;
        RECT 76.910 103.910 77.170 104.230 ;
        RECT 73.690 101.870 73.950 102.190 ;
        RECT 74.150 100.850 74.410 101.170 ;
        RECT 74.210 99.130 74.350 100.850 ;
        RECT 76.970 100.150 77.110 103.910 ;
        RECT 76.910 99.830 77.170 100.150 ;
        RECT 74.150 98.810 74.410 99.130 ;
        RECT 71.850 98.130 72.110 98.450 ;
        RECT 70.470 96.090 70.730 96.410 ;
        RECT 71.910 89.890 72.050 98.130 ;
        RECT 76.970 95.730 77.110 99.830 ;
        RECT 76.450 95.410 76.710 95.730 ;
        RECT 76.910 95.410 77.170 95.730 ;
        RECT 76.510 93.690 76.650 95.410 ;
        RECT 76.450 93.370 76.710 93.690 ;
        RECT 76.510 91.310 76.650 93.370 ;
        RECT 76.450 90.990 76.710 91.310 ;
        RECT 70.990 89.750 72.050 89.890 ;
        RECT 70.990 88.590 71.130 89.750 ;
        RECT 70.930 88.270 71.190 88.590 ;
        RECT 76.970 88.250 77.110 95.410 ;
        RECT 77.430 88.250 77.570 106.290 ;
        RECT 77.890 104.910 78.030 114.540 ;
        RECT 79.270 111.030 79.410 141.990 ;
        RECT 81.570 138.190 81.710 146.070 ;
        RECT 83.340 145.535 83.620 145.905 ;
        RECT 84.730 145.730 84.990 146.050 ;
        RECT 86.170 145.905 86.310 147.770 ;
        RECT 83.350 145.390 83.610 145.535 ;
        RECT 84.790 143.670 84.930 145.730 ;
        RECT 86.100 145.535 86.380 145.905 ;
        RECT 84.730 143.350 84.990 143.670 ;
        RECT 84.270 141.990 84.530 142.310 ;
        RECT 81.110 138.050 81.710 138.190 ;
        RECT 80.590 136.550 80.850 136.870 ;
        RECT 80.130 136.210 80.390 136.530 ;
        RECT 80.190 134.830 80.330 136.210 ;
        RECT 80.650 135.510 80.790 136.550 ;
        RECT 80.590 135.190 80.850 135.510 ;
        RECT 80.130 134.510 80.390 134.830 ;
        RECT 80.590 131.110 80.850 131.430 ;
        RECT 80.650 129.390 80.790 131.110 ;
        RECT 81.110 129.730 81.250 138.050 ;
        RECT 81.510 136.890 81.770 137.210 ;
        RECT 81.970 136.890 82.230 137.210 ;
        RECT 81.570 134.830 81.710 136.890 ;
        RECT 81.510 134.510 81.770 134.830 ;
        RECT 81.570 132.110 81.710 134.510 ;
        RECT 82.030 132.790 82.170 136.890 ;
        RECT 81.970 132.470 82.230 132.790 ;
        RECT 82.430 132.190 82.690 132.450 ;
        RECT 82.030 132.130 82.690 132.190 ;
        RECT 81.510 131.790 81.770 132.110 ;
        RECT 82.030 132.050 82.630 132.130 ;
        RECT 81.050 129.410 81.310 129.730 ;
        RECT 80.590 129.070 80.850 129.390 ;
        RECT 80.650 127.350 80.790 129.070 ;
        RECT 80.590 127.030 80.850 127.350 ;
        RECT 80.650 126.330 80.790 127.030 ;
        RECT 80.590 126.010 80.850 126.330 ;
        RECT 81.050 125.330 81.310 125.650 ;
        RECT 81.110 123.610 81.250 125.330 ;
        RECT 81.570 123.950 81.710 131.790 ;
        RECT 82.030 129.390 82.170 132.050 ;
        RECT 82.430 130.770 82.690 131.090 ;
        RECT 82.490 130.070 82.630 130.770 ;
        RECT 82.430 129.750 82.690 130.070 ;
        RECT 81.970 129.070 82.230 129.390 ;
        RECT 83.810 125.670 84.070 125.990 ;
        RECT 83.350 124.200 83.610 124.290 ;
        RECT 83.870 124.200 84.010 125.670 ;
        RECT 83.350 124.060 84.010 124.200 ;
        RECT 83.350 123.970 83.610 124.060 ;
        RECT 81.510 123.630 81.770 123.950 ;
        RECT 80.590 123.290 80.850 123.610 ;
        RECT 81.050 123.290 81.310 123.610 ;
        RECT 80.650 118.510 80.790 123.290 ;
        RECT 81.570 121.230 81.710 123.630 ;
        RECT 81.510 120.910 81.770 121.230 ;
        RECT 81.570 118.850 81.710 120.910 ;
        RECT 81.510 118.530 81.770 118.850 ;
        RECT 80.590 118.420 80.850 118.510 ;
        RECT 79.730 118.280 80.850 118.420 ;
        RECT 79.210 110.710 79.470 111.030 ;
        RECT 79.210 109.350 79.470 109.670 ;
        RECT 78.750 107.990 79.010 108.310 ;
        RECT 78.290 107.310 78.550 107.630 ;
        RECT 78.350 105.590 78.490 107.310 ;
        RECT 78.290 105.270 78.550 105.590 ;
        RECT 78.810 105.250 78.950 107.990 ;
        RECT 79.270 106.610 79.410 109.350 ;
        RECT 79.210 106.290 79.470 106.610 ;
        RECT 78.750 104.930 79.010 105.250 ;
        RECT 77.830 104.590 78.090 104.910 ;
        RECT 78.290 103.910 78.550 104.230 ;
        RECT 78.350 102.190 78.490 103.910 ;
        RECT 78.290 101.870 78.550 102.190 ;
        RECT 78.350 101.590 78.490 101.870 ;
        RECT 77.890 101.450 78.490 101.590 ;
        RECT 78.810 101.510 78.950 104.930 ;
        RECT 77.890 98.450 78.030 101.450 ;
        RECT 78.750 101.190 79.010 101.510 ;
        RECT 79.730 99.130 79.870 118.280 ;
        RECT 80.590 118.190 80.850 118.280 ;
        RECT 83.870 116.470 84.010 124.060 ;
        RECT 83.810 116.150 84.070 116.470 ;
        RECT 81.050 109.690 81.310 110.010 ;
        RECT 83.350 109.690 83.610 110.010 ;
        RECT 80.590 109.010 80.850 109.330 ;
        RECT 80.130 106.630 80.390 106.950 ;
        RECT 80.190 104.570 80.330 106.630 ;
        RECT 80.650 104.570 80.790 109.010 ;
        RECT 80.130 104.250 80.390 104.570 ;
        RECT 80.590 104.250 80.850 104.570 ;
        RECT 80.190 102.870 80.330 104.250 ;
        RECT 80.590 103.570 80.850 103.890 ;
        RECT 80.130 102.550 80.390 102.870 ;
        RECT 80.190 99.130 80.330 102.550 ;
        RECT 80.650 99.130 80.790 103.570 ;
        RECT 81.110 102.530 81.250 109.690 ;
        RECT 81.510 106.970 81.770 107.290 ;
        RECT 81.570 105.250 81.710 106.970 ;
        RECT 81.510 104.930 81.770 105.250 ;
        RECT 81.570 104.570 81.710 104.930 ;
        RECT 83.410 104.570 83.550 109.690 ;
        RECT 84.330 105.590 84.470 141.990 ;
        RECT 85.650 136.210 85.910 136.530 ;
        RECT 85.710 134.830 85.850 136.210 ;
        RECT 85.650 134.510 85.910 134.830 ;
        RECT 86.110 133.490 86.370 133.810 ;
        RECT 84.730 131.110 84.990 131.430 ;
        RECT 84.790 130.070 84.930 131.110 ;
        RECT 84.730 129.750 84.990 130.070 ;
        RECT 86.170 129.050 86.310 133.490 ;
        RECT 86.110 128.730 86.370 129.050 ;
        RECT 86.170 125.990 86.310 128.730 ;
        RECT 86.110 125.670 86.370 125.990 ;
        RECT 84.730 125.330 84.990 125.650 ;
        RECT 84.790 124.290 84.930 125.330 ;
        RECT 84.730 123.970 84.990 124.290 ;
        RECT 85.650 114.790 85.910 115.110 ;
        RECT 85.710 113.410 85.850 114.790 ;
        RECT 85.650 113.090 85.910 113.410 ;
        RECT 84.730 112.750 84.990 113.070 ;
        RECT 84.790 108.310 84.930 112.750 ;
        RECT 85.190 109.690 85.450 110.010 ;
        RECT 84.730 107.990 84.990 108.310 ;
        RECT 85.250 107.970 85.390 109.690 ;
        RECT 85.710 109.670 85.850 113.090 ;
        RECT 85.650 109.350 85.910 109.670 ;
        RECT 85.190 107.650 85.450 107.970 ;
        RECT 85.710 107.630 85.850 109.350 ;
        RECT 85.650 107.310 85.910 107.630 ;
        RECT 84.270 105.270 84.530 105.590 ;
        RECT 84.720 104.735 85.000 105.105 ;
        RECT 85.710 104.910 85.850 107.310 ;
        RECT 84.790 104.570 84.930 104.735 ;
        RECT 85.650 104.590 85.910 104.910 ;
        RECT 81.510 104.250 81.770 104.570 ;
        RECT 83.350 104.250 83.610 104.570 ;
        RECT 84.730 104.250 84.990 104.570 ;
        RECT 81.050 102.210 81.310 102.530 ;
        RECT 81.050 101.530 81.310 101.850 ;
        RECT 81.110 100.150 81.250 101.530 ;
        RECT 81.570 100.150 81.710 104.250 ;
        RECT 83.410 102.190 83.550 104.250 ;
        RECT 84.720 103.375 85.000 103.745 ;
        RECT 83.350 101.870 83.610 102.190 ;
        RECT 84.790 101.170 84.930 103.375 ;
        RECT 85.190 101.870 85.450 102.190 ;
        RECT 84.730 100.850 84.990 101.170 ;
        RECT 81.050 99.830 81.310 100.150 ;
        RECT 81.510 99.830 81.770 100.150 ;
        RECT 81.570 99.130 81.710 99.830 ;
        RECT 79.670 98.810 79.930 99.130 ;
        RECT 80.130 98.810 80.390 99.130 ;
        RECT 80.590 98.810 80.850 99.130 ;
        RECT 81.510 98.810 81.770 99.130 ;
        RECT 77.830 98.130 78.090 98.450 ;
        RECT 78.290 98.130 78.550 98.450 ;
        RECT 77.890 88.250 78.030 98.130 ;
        RECT 78.350 96.750 78.490 98.130 ;
        RECT 79.730 96.750 79.870 98.810 ;
        RECT 81.570 97.430 81.710 98.810 ;
        RECT 81.510 97.110 81.770 97.430 ;
        RECT 84.790 96.750 84.930 100.850 ;
        RECT 85.250 100.150 85.390 101.870 ;
        RECT 85.190 99.830 85.450 100.150 ;
        RECT 85.710 99.550 85.850 104.590 ;
        RECT 86.110 104.250 86.370 104.570 ;
        RECT 85.250 99.410 85.850 99.550 ;
        RECT 78.290 96.430 78.550 96.750 ;
        RECT 79.670 96.430 79.930 96.750 ;
        RECT 84.730 96.430 84.990 96.750 ;
        RECT 84.270 96.090 84.530 96.410 ;
        RECT 79.670 95.410 79.930 95.730 ;
        RECT 83.350 95.410 83.610 95.730 ;
        RECT 79.730 93.350 79.870 95.410 ;
        RECT 79.670 93.030 79.930 93.350 ;
        RECT 83.410 91.650 83.550 95.410 ;
        RECT 84.330 91.650 84.470 96.090 ;
        RECT 85.250 93.690 85.390 99.410 ;
        RECT 85.650 96.430 85.910 96.750 ;
        RECT 85.190 93.370 85.450 93.690 ;
        RECT 85.710 91.990 85.850 96.430 ;
        RECT 86.170 96.070 86.310 104.250 ;
        RECT 86.630 102.190 86.770 151.170 ;
        RECT 87.090 146.390 87.230 157.970 ;
        RECT 92.610 156.590 92.750 158.990 ;
        RECT 92.550 156.270 92.810 156.590 ;
        RECT 87.490 152.530 87.750 152.850 ;
        RECT 87.550 151.830 87.690 152.530 ;
        RECT 87.490 151.510 87.750 151.830 ;
        RECT 91.630 150.490 91.890 150.810 ;
        RECT 91.170 149.810 91.430 150.130 ;
        RECT 91.230 147.750 91.370 149.810 ;
        RECT 91.170 147.430 91.430 147.750 ;
        RECT 87.030 146.070 87.290 146.390 ;
        RECT 88.870 146.070 89.130 146.390 ;
        RECT 88.930 142.990 89.070 146.070 ;
        RECT 88.870 142.670 89.130 142.990 ;
        RECT 87.950 136.210 88.210 136.530 ;
        RECT 90.710 136.210 90.970 136.530 ;
        RECT 88.010 133.810 88.150 136.210 ;
        RECT 90.770 133.810 90.910 136.210 ;
        RECT 87.950 133.490 88.210 133.810 ;
        RECT 90.710 133.490 90.970 133.810 ;
        RECT 87.490 130.770 87.750 131.090 ;
        RECT 87.550 129.050 87.690 130.770 ;
        RECT 90.250 129.750 90.510 130.070 ;
        RECT 87.490 128.730 87.750 129.050 ;
        RECT 89.790 128.050 90.050 128.370 ;
        RECT 89.850 124.290 89.990 128.050 ;
        RECT 90.310 125.650 90.450 129.750 ;
        RECT 91.170 129.410 91.430 129.730 ;
        RECT 90.250 125.330 90.510 125.650 ;
        RECT 89.790 123.970 90.050 124.290 ;
        RECT 90.310 123.610 90.450 125.330 ;
        RECT 90.250 123.350 90.510 123.610 ;
        RECT 89.850 123.290 90.510 123.350 ;
        RECT 89.850 123.210 90.450 123.290 ;
        RECT 87.030 114.450 87.290 114.770 ;
        RECT 87.090 107.630 87.230 114.450 ;
        RECT 88.410 110.710 88.670 111.030 ;
        RECT 87.490 109.010 87.750 109.330 ;
        RECT 87.950 109.010 88.210 109.330 ;
        RECT 87.550 108.310 87.690 109.010 ;
        RECT 87.490 107.990 87.750 108.310 ;
        RECT 88.010 107.630 88.150 109.010 ;
        RECT 87.030 107.310 87.290 107.630 ;
        RECT 87.490 107.310 87.750 107.630 ;
        RECT 87.950 107.310 88.210 107.630 ;
        RECT 87.090 105.590 87.230 107.310 ;
        RECT 87.550 106.610 87.690 107.310 ;
        RECT 87.490 106.290 87.750 106.610 ;
        RECT 87.030 105.270 87.290 105.590 ;
        RECT 87.030 103.910 87.290 104.230 ;
        RECT 87.090 102.870 87.230 103.910 ;
        RECT 88.470 103.890 88.610 110.710 ;
        RECT 89.850 107.710 89.990 123.210 ;
        RECT 90.710 122.950 90.970 123.270 ;
        RECT 90.250 122.610 90.510 122.930 ;
        RECT 90.310 120.890 90.450 122.610 ;
        RECT 90.770 121.910 90.910 122.950 ;
        RECT 90.710 121.590 90.970 121.910 ;
        RECT 90.250 120.570 90.510 120.890 ;
        RECT 91.230 118.510 91.370 129.410 ;
        RECT 91.170 118.190 91.430 118.510 ;
        RECT 90.710 114.450 90.970 114.770 ;
        RECT 90.770 113.750 90.910 114.450 ;
        RECT 90.710 113.430 90.970 113.750 ;
        RECT 91.230 113.265 91.370 118.190 ;
        RECT 91.690 113.750 91.830 150.490 ;
        RECT 92.610 148.090 92.750 156.270 ;
        RECT 93.530 151.490 93.670 168.850 ;
        RECT 93.990 165.090 94.130 172.590 ;
        RECT 94.450 170.190 94.590 178.030 ;
        RECT 95.370 176.310 95.510 180.410 ;
        RECT 103.650 180.390 103.790 182.450 ;
        RECT 103.590 180.070 103.850 180.390 ;
        RECT 101.290 179.730 101.550 180.050 ;
        RECT 101.350 178.350 101.490 179.730 ;
        RECT 101.290 178.030 101.550 178.350 ;
        RECT 98.070 177.690 98.330 178.010 ;
        RECT 95.310 175.990 95.570 176.310 ;
        RECT 98.130 175.290 98.270 177.690 ;
        RECT 103.130 175.310 103.390 175.630 ;
        RECT 98.070 174.970 98.330 175.290 ;
        RECT 98.130 172.570 98.270 174.970 ;
        RECT 99.450 174.290 99.710 174.610 ;
        RECT 98.070 172.250 98.330 172.570 ;
        RECT 94.390 169.870 94.650 170.190 ;
        RECT 93.930 164.770 94.190 165.090 ;
        RECT 94.450 164.410 94.590 169.870 ;
        RECT 97.150 169.190 97.410 169.510 ;
        RECT 97.210 165.430 97.350 169.190 ;
        RECT 98.130 167.380 98.270 172.250 ;
        RECT 98.530 167.380 98.790 167.470 ;
        RECT 98.130 167.240 98.790 167.380 ;
        RECT 98.530 167.150 98.790 167.240 ;
        RECT 97.150 165.110 97.410 165.430 ;
        RECT 99.510 164.750 99.650 174.290 ;
        RECT 103.190 173.590 103.330 175.310 ;
        RECT 103.130 173.270 103.390 173.590 ;
        RECT 100.830 168.850 101.090 169.170 ;
        RECT 100.890 167.470 101.030 168.850 ;
        RECT 103.190 167.470 103.330 173.270 ;
        RECT 100.830 167.150 101.090 167.470 ;
        RECT 103.130 167.150 103.390 167.470 ;
        RECT 99.450 164.430 99.710 164.750 ;
        RECT 94.390 164.090 94.650 164.410 ;
        RECT 97.150 164.090 97.410 164.410 ;
        RECT 95.770 163.750 96.030 164.070 ;
        RECT 95.830 162.370 95.970 163.750 ;
        RECT 95.770 162.050 96.030 162.370 ;
        RECT 97.210 162.030 97.350 164.090 ;
        RECT 98.990 163.410 99.250 163.730 ;
        RECT 97.150 161.710 97.410 162.030 ;
        RECT 97.210 155.570 97.350 161.710 ;
        RECT 97.150 155.250 97.410 155.570 ;
        RECT 97.210 153.950 97.350 155.250 ;
        RECT 97.210 153.870 97.810 153.950 ;
        RECT 97.210 153.810 97.870 153.870 ;
        RECT 97.610 153.550 97.870 153.810 ;
        RECT 93.470 151.170 93.730 151.490 ;
        RECT 93.530 148.770 93.670 151.170 ;
        RECT 94.390 150.150 94.650 150.470 ;
        RECT 94.450 149.110 94.590 150.150 ;
        RECT 94.390 148.790 94.650 149.110 ;
        RECT 93.470 148.450 93.730 148.770 ;
        RECT 92.550 147.770 92.810 148.090 ;
        RECT 92.610 145.710 92.750 147.770 ;
        RECT 92.090 145.390 92.350 145.710 ;
        RECT 92.550 145.390 92.810 145.710 ;
        RECT 92.150 137.550 92.290 145.390 ;
        RECT 92.610 142.990 92.750 145.390 ;
        RECT 99.050 143.670 99.190 163.410 ;
        RECT 99.910 162.050 100.170 162.370 ;
        RECT 99.450 161.370 99.710 161.690 ;
        RECT 99.510 159.310 99.650 161.370 ;
        RECT 99.450 158.990 99.710 159.310 ;
        RECT 99.510 157.270 99.650 158.990 ;
        RECT 99.450 156.950 99.710 157.270 ;
        RECT 99.450 144.710 99.710 145.030 ;
        RECT 98.990 143.350 99.250 143.670 ;
        RECT 99.510 143.070 99.650 144.710 ;
        RECT 92.550 142.670 92.810 142.990 ;
        RECT 99.050 142.930 99.650 143.070 ;
        RECT 99.050 142.650 99.190 142.930 ;
        RECT 98.990 142.330 99.250 142.650 ;
        RECT 97.150 141.990 97.410 142.310 ;
        RECT 97.210 140.950 97.350 141.990 ;
        RECT 97.150 140.630 97.410 140.950 ;
        RECT 99.050 139.930 99.190 142.330 ;
        RECT 98.990 139.610 99.250 139.930 ;
        RECT 92.090 137.230 92.350 137.550 ;
        RECT 94.390 136.210 94.650 136.530 ;
        RECT 96.690 136.210 96.950 136.530 ;
        RECT 94.450 135.170 94.590 136.210 ;
        RECT 94.390 134.850 94.650 135.170 ;
        RECT 93.010 134.510 93.270 134.830 ;
        RECT 93.070 132.110 93.210 134.510 ;
        RECT 94.850 133.550 95.110 133.810 ;
        RECT 94.850 133.490 95.510 133.550 ;
        RECT 94.910 133.410 95.510 133.490 ;
        RECT 93.010 131.790 93.270 132.110 ;
        RECT 94.850 131.110 95.110 131.430 ;
        RECT 93.470 130.770 93.730 131.090 ;
        RECT 93.530 129.390 93.670 130.770 ;
        RECT 93.470 129.070 93.730 129.390 ;
        RECT 92.090 118.190 92.350 118.510 ;
        RECT 91.630 113.430 91.890 113.750 ;
        RECT 91.160 112.895 91.440 113.265 ;
        RECT 92.150 113.070 92.290 118.190 ;
        RECT 93.010 115.470 93.270 115.790 ;
        RECT 91.230 110.010 91.370 112.895 ;
        RECT 92.090 112.750 92.350 113.070 ;
        RECT 92.550 112.750 92.810 113.070 ;
        RECT 92.150 110.350 92.290 112.750 ;
        RECT 92.610 112.050 92.750 112.750 ;
        RECT 92.550 111.730 92.810 112.050 ;
        RECT 92.090 110.030 92.350 110.350 ;
        RECT 91.170 109.690 91.430 110.010 ;
        RECT 92.090 109.580 92.350 109.670 ;
        RECT 92.610 109.580 92.750 111.730 ;
        RECT 92.090 109.440 92.750 109.580 ;
        RECT 92.090 109.350 92.350 109.440 ;
        RECT 89.850 107.570 90.450 107.710 ;
        RECT 89.790 106.970 90.050 107.290 ;
        RECT 88.870 106.630 89.130 106.950 ;
        RECT 88.410 103.570 88.670 103.890 ;
        RECT 87.030 102.550 87.290 102.870 ;
        RECT 88.470 102.780 88.610 103.570 ;
        RECT 88.010 102.640 88.610 102.780 ;
        RECT 88.010 102.190 88.150 102.640 ;
        RECT 86.570 101.870 86.830 102.190 ;
        RECT 87.950 101.870 88.210 102.190 ;
        RECT 87.030 101.530 87.290 101.850 ;
        RECT 87.090 96.750 87.230 101.530 ;
        RECT 87.950 98.810 88.210 99.130 ;
        RECT 88.010 96.750 88.150 98.810 ;
        RECT 88.930 98.790 89.070 106.630 ;
        RECT 89.850 102.190 89.990 106.970 ;
        RECT 89.790 101.870 90.050 102.190 ;
        RECT 88.410 98.470 88.670 98.790 ;
        RECT 88.870 98.470 89.130 98.790 ;
        RECT 87.030 96.430 87.290 96.750 ;
        RECT 87.950 96.430 88.210 96.750 ;
        RECT 87.490 96.090 87.750 96.410 ;
        RECT 86.110 95.750 86.370 96.070 ;
        RECT 85.650 91.670 85.910 91.990 ;
        RECT 83.350 91.330 83.610 91.650 ;
        RECT 84.270 91.330 84.530 91.650 ;
        RECT 87.550 90.970 87.690 96.090 ;
        RECT 88.470 94.710 88.610 98.470 ;
        RECT 88.930 96.750 89.070 98.470 ;
        RECT 88.870 96.430 89.130 96.750 ;
        RECT 89.790 96.430 90.050 96.750 ;
        RECT 89.850 94.790 89.990 96.430 ;
        RECT 90.310 95.730 90.450 107.570 ;
        RECT 91.630 107.310 91.890 107.630 ;
        RECT 91.690 104.910 91.830 107.310 ;
        RECT 91.630 104.590 91.890 104.910 ;
        RECT 91.690 99.470 91.830 104.590 ;
        RECT 91.630 99.150 91.890 99.470 ;
        RECT 91.630 96.770 91.890 97.090 ;
        RECT 90.710 95.750 90.970 96.070 ;
        RECT 90.250 95.410 90.510 95.730 ;
        RECT 89.850 94.710 90.450 94.790 ;
        RECT 88.410 94.390 88.670 94.710 ;
        RECT 89.850 94.650 90.510 94.710 ;
        RECT 90.250 94.390 90.510 94.650 ;
        RECT 88.470 91.650 88.610 94.390 ;
        RECT 90.770 91.650 90.910 95.750 ;
        RECT 91.170 93.030 91.430 93.350 ;
        RECT 91.230 91.990 91.370 93.030 ;
        RECT 91.690 91.990 91.830 96.770 ;
        RECT 91.170 91.670 91.430 91.990 ;
        RECT 91.630 91.670 91.890 91.990 ;
        RECT 88.410 91.330 88.670 91.650 ;
        RECT 90.710 91.330 90.970 91.650 ;
        RECT 87.490 90.650 87.750 90.970 ;
        RECT 83.810 90.310 84.070 90.630 ;
        RECT 83.870 88.250 84.010 90.310 ;
        RECT 88.470 88.250 88.610 91.330 ;
        RECT 92.150 88.250 92.290 109.350 ;
        RECT 93.070 107.630 93.210 115.470 ;
        RECT 92.550 107.310 92.810 107.630 ;
        RECT 93.010 107.310 93.270 107.630 ;
        RECT 92.610 105.250 92.750 107.310 ;
        RECT 92.550 104.930 92.810 105.250 ;
        RECT 93.010 103.570 93.270 103.890 ;
        RECT 93.070 102.530 93.210 103.570 ;
        RECT 93.010 102.210 93.270 102.530 ;
        RECT 93.010 98.130 93.270 98.450 ;
        RECT 92.550 96.430 92.810 96.750 ;
        RECT 92.610 93.010 92.750 96.430 ;
        RECT 92.550 92.690 92.810 93.010 ;
        RECT 92.540 91.135 92.820 91.505 ;
        RECT 92.550 90.990 92.810 91.135 ;
        RECT 93.070 90.630 93.210 98.130 ;
        RECT 93.530 91.505 93.670 129.070 ;
        RECT 94.910 116.470 95.050 131.110 ;
        RECT 95.370 125.990 95.510 133.410 ;
        RECT 95.770 126.010 96.030 126.330 ;
        RECT 95.310 125.670 95.570 125.990 ;
        RECT 94.850 116.150 95.110 116.470 ;
        RECT 94.910 106.610 95.050 116.150 ;
        RECT 94.850 106.290 95.110 106.610 ;
        RECT 93.930 104.930 94.190 105.250 ;
        RECT 93.990 104.230 94.130 104.930 ;
        RECT 93.930 103.910 94.190 104.230 ;
        RECT 94.850 103.910 95.110 104.230 ;
        RECT 93.460 91.135 93.740 91.505 ;
        RECT 93.010 90.310 93.270 90.630 ;
        RECT 93.990 88.250 94.130 103.910 ;
        RECT 94.910 97.430 95.050 103.910 ;
        RECT 94.850 97.110 95.110 97.430 ;
        RECT 94.390 96.430 94.650 96.750 ;
        RECT 94.450 91.990 94.590 96.430 ;
        RECT 94.390 91.670 94.650 91.990 ;
        RECT 94.910 91.310 95.050 97.110 ;
        RECT 95.370 96.750 95.510 125.670 ;
        RECT 95.830 123.610 95.970 126.010 ;
        RECT 95.770 123.290 96.030 123.610 ;
        RECT 95.830 118.850 95.970 123.290 ;
        RECT 96.750 122.930 96.890 136.210 ;
        RECT 99.970 132.790 100.110 162.050 ;
        RECT 100.370 161.030 100.630 161.350 ;
        RECT 100.430 159.990 100.570 161.030 ;
        RECT 101.290 160.690 101.550 161.010 ;
        RECT 100.370 159.670 100.630 159.990 ;
        RECT 100.430 154.210 100.570 159.670 ;
        RECT 101.350 158.970 101.490 160.690 ;
        RECT 101.290 158.650 101.550 158.970 ;
        RECT 103.650 158.630 103.790 180.070 ;
        RECT 104.110 178.350 104.250 186.350 ;
        RECT 104.970 179.730 105.230 180.050 ;
        RECT 105.030 178.690 105.170 179.730 ;
        RECT 104.970 178.370 105.230 178.690 ;
        RECT 104.050 178.030 104.310 178.350 ;
        RECT 104.510 178.030 104.770 178.350 ;
        RECT 104.570 175.970 104.710 178.030 ;
        RECT 105.030 176.310 105.170 178.370 ;
        RECT 104.970 175.990 105.230 176.310 ;
        RECT 104.510 175.650 104.770 175.970 ;
        RECT 104.050 174.970 104.310 175.290 ;
        RECT 104.110 174.610 104.250 174.970 ;
        RECT 104.050 174.290 104.310 174.610 ;
        RECT 105.030 173.250 105.170 175.990 ;
        RECT 104.970 172.930 105.230 173.250 ;
        RECT 104.050 172.590 104.310 172.910 ;
        RECT 104.110 164.410 104.250 172.590 ;
        RECT 104.510 167.830 104.770 168.150 ;
        RECT 104.570 165.430 104.710 167.830 ;
        RECT 104.970 166.810 105.230 167.130 ;
        RECT 104.510 165.110 104.770 165.430 ;
        RECT 104.050 164.090 104.310 164.410 ;
        RECT 105.030 162.370 105.170 166.810 ;
        RECT 105.490 164.750 105.630 187.890 ;
        RECT 105.950 187.190 106.090 189.250 ;
        RECT 105.890 186.870 106.150 187.190 ;
        RECT 106.410 185.830 106.550 191.970 ;
        RECT 108.710 191.610 108.850 196.050 ;
        RECT 110.950 194.350 111.210 194.670 ;
        RECT 112.790 194.350 113.050 194.670 ;
        RECT 109.110 193.330 109.370 193.650 ;
        RECT 106.810 191.290 107.070 191.610 ;
        RECT 108.650 191.290 108.910 191.610 ;
        RECT 106.870 188.210 107.010 191.290 ;
        RECT 106.810 187.890 107.070 188.210 ;
        RECT 107.730 187.890 107.990 188.210 ;
        RECT 106.350 185.510 106.610 185.830 ;
        RECT 106.410 180.730 106.550 185.510 ;
        RECT 106.810 185.170 107.070 185.490 ;
        RECT 107.270 185.170 107.530 185.490 ;
        RECT 106.870 184.665 107.010 185.170 ;
        RECT 106.800 184.295 107.080 184.665 ;
        RECT 107.330 183.450 107.470 185.170 ;
        RECT 107.790 183.790 107.930 187.890 ;
        RECT 108.710 187.190 108.850 191.290 ;
        RECT 109.170 191.270 109.310 193.330 ;
        RECT 110.490 191.630 110.750 191.950 ;
        RECT 109.110 190.950 109.370 191.270 ;
        RECT 109.170 189.480 109.310 190.950 ;
        RECT 109.570 189.480 109.830 189.570 ;
        RECT 109.170 189.340 109.830 189.480 ;
        RECT 109.570 189.250 109.830 189.340 ;
        RECT 109.630 188.550 109.770 189.250 ;
        RECT 109.570 188.230 109.830 188.550 ;
        RECT 108.650 186.870 108.910 187.190 ;
        RECT 109.630 186.510 109.770 188.230 ;
        RECT 109.570 186.190 109.830 186.510 ;
        RECT 110.550 184.380 110.690 191.630 ;
        RECT 111.010 191.270 111.150 194.350 ;
        RECT 112.850 191.950 112.990 194.350 ;
        RECT 113.310 192.630 113.450 196.390 ;
        RECT 113.770 194.330 113.910 198.770 ;
        RECT 115.090 196.390 115.350 196.710 ;
        RECT 115.150 195.350 115.290 196.390 ;
        RECT 116.530 196.370 116.670 199.790 ;
        RECT 124.750 196.730 125.010 197.050 ;
        RECT 116.470 196.050 116.730 196.370 ;
        RECT 115.090 195.030 115.350 195.350 ;
        RECT 113.710 194.010 113.970 194.330 ;
        RECT 113.250 192.310 113.510 192.630 ;
        RECT 112.790 191.630 113.050 191.950 ;
        RECT 113.770 191.610 113.910 194.010 ;
        RECT 115.550 192.310 115.810 192.630 ;
        RECT 114.170 191.970 114.430 192.290 ;
        RECT 114.230 191.610 114.370 191.970 ;
        RECT 113.710 191.465 113.970 191.610 ;
        RECT 110.950 190.950 111.210 191.270 ;
        RECT 111.870 190.950 112.130 191.270 ;
        RECT 113.700 191.095 113.980 191.465 ;
        RECT 114.170 191.290 114.430 191.610 ;
        RECT 110.940 190.415 111.220 190.785 ;
        RECT 111.010 186.170 111.150 190.415 ;
        RECT 111.930 189.910 112.070 190.950 ;
        RECT 113.710 190.610 113.970 190.930 ;
        RECT 111.870 189.590 112.130 189.910 ;
        RECT 111.870 188.910 112.130 189.230 ;
        RECT 111.410 187.890 111.670 188.210 ;
        RECT 111.470 186.850 111.610 187.890 ;
        RECT 111.410 186.530 111.670 186.850 ;
        RECT 110.950 185.850 111.210 186.170 ;
        RECT 110.090 184.240 110.690 184.380 ;
        RECT 107.730 183.470 107.990 183.790 ;
        RECT 107.270 183.130 107.530 183.450 ;
        RECT 109.570 183.130 109.830 183.450 ;
        RECT 107.730 182.790 107.990 183.110 ;
        RECT 107.790 181.750 107.930 182.790 ;
        RECT 108.650 182.450 108.910 182.770 ;
        RECT 107.730 181.430 107.990 181.750 ;
        RECT 108.710 180.730 108.850 182.450 ;
        RECT 109.630 180.730 109.770 183.130 ;
        RECT 106.350 180.410 106.610 180.730 ;
        RECT 107.270 180.410 107.530 180.730 ;
        RECT 108.650 180.410 108.910 180.730 ;
        RECT 109.570 180.585 109.830 180.730 ;
        RECT 106.410 178.350 106.550 180.410 ;
        RECT 106.810 179.730 107.070 180.050 ;
        RECT 106.870 179.030 107.010 179.730 ;
        RECT 107.330 179.225 107.470 180.410 ;
        RECT 106.810 178.710 107.070 179.030 ;
        RECT 107.260 178.855 107.540 179.225 ;
        RECT 106.350 178.030 106.610 178.350 ;
        RECT 107.330 178.010 107.470 178.855 ;
        RECT 108.710 178.350 108.850 180.410 ;
        RECT 109.560 180.215 109.840 180.585 ;
        RECT 108.650 178.030 108.910 178.350 ;
        RECT 107.270 177.690 107.530 178.010 ;
        RECT 106.810 177.350 107.070 177.670 ;
        RECT 105.890 168.850 106.150 169.170 ;
        RECT 105.950 167.470 106.090 168.850 ;
        RECT 105.890 167.150 106.150 167.470 ;
        RECT 106.870 165.430 107.010 177.350 ;
        RECT 107.330 175.290 107.470 177.690 ;
        RECT 109.570 177.010 109.830 177.330 ;
        RECT 107.270 174.970 107.530 175.290 ;
        RECT 107.330 167.665 107.470 174.970 ;
        RECT 109.110 168.850 109.370 169.170 ;
        RECT 107.260 167.295 107.540 167.665 ;
        RECT 107.270 167.150 107.530 167.295 ;
        RECT 108.650 167.150 108.910 167.470 ;
        RECT 108.190 166.470 108.450 166.790 ;
        RECT 106.810 165.110 107.070 165.430 ;
        RECT 105.430 164.430 105.690 164.750 ;
        RECT 106.350 163.410 106.610 163.730 ;
        RECT 106.410 162.370 106.550 163.410 ;
        RECT 104.970 162.050 105.230 162.370 ;
        RECT 106.350 162.050 106.610 162.370 ;
        RECT 107.730 158.890 107.990 158.970 ;
        RECT 108.250 158.890 108.390 166.470 ;
        RECT 107.730 158.750 108.390 158.890 ;
        RECT 107.730 158.650 107.990 158.750 ;
        RECT 103.590 158.310 103.850 158.630 ;
        RECT 106.350 158.310 106.610 158.630 ;
        RECT 106.410 156.590 106.550 158.310 ;
        RECT 106.350 156.270 106.610 156.590 ;
        RECT 101.290 155.250 101.550 155.570 ;
        RECT 100.370 153.890 100.630 154.210 ;
        RECT 101.350 153.530 101.490 155.250 ;
        RECT 108.710 153.530 108.850 167.150 ;
        RECT 109.170 167.130 109.310 168.850 ;
        RECT 109.110 166.810 109.370 167.130 ;
        RECT 109.110 161.710 109.370 162.030 ;
        RECT 109.170 159.990 109.310 161.710 ;
        RECT 109.110 159.670 109.370 159.990 ;
        RECT 109.630 159.390 109.770 177.010 ;
        RECT 110.090 167.380 110.230 184.240 ;
        RECT 110.490 183.470 110.750 183.790 ;
        RECT 110.550 177.670 110.690 183.470 ;
        RECT 111.470 183.450 111.610 186.530 ;
        RECT 111.930 186.170 112.070 188.910 ;
        RECT 113.250 188.230 113.510 188.550 ;
        RECT 112.790 187.890 113.050 188.210 ;
        RECT 111.870 185.850 112.130 186.170 ;
        RECT 112.850 185.740 112.990 187.890 ;
        RECT 113.310 186.760 113.450 188.230 ;
        RECT 113.770 188.210 113.910 190.610 ;
        RECT 113.710 187.890 113.970 188.210 ;
        RECT 113.710 186.760 113.970 186.850 ;
        RECT 113.310 186.620 113.970 186.760 ;
        RECT 113.710 186.530 113.970 186.620 ;
        RECT 112.850 185.600 113.450 185.740 ;
        RECT 111.870 185.170 112.130 185.490 ;
        RECT 110.940 182.935 111.220 183.305 ;
        RECT 111.410 183.130 111.670 183.450 ;
        RECT 111.930 183.190 112.070 185.170 ;
        RECT 112.780 184.295 113.060 184.665 ;
        RECT 112.850 184.130 112.990 184.295 ;
        RECT 112.790 183.810 113.050 184.130 ;
        RECT 113.310 183.190 113.450 185.600 ;
        RECT 113.770 185.490 113.910 186.530 ;
        RECT 114.230 186.510 114.370 191.290 ;
        RECT 114.630 187.890 114.890 188.210 ;
        RECT 115.090 187.890 115.350 188.210 ;
        RECT 114.690 187.190 114.830 187.890 ;
        RECT 114.630 186.870 114.890 187.190 ;
        RECT 114.170 186.190 114.430 186.510 ;
        RECT 114.630 185.510 114.890 185.830 ;
        RECT 113.710 185.170 113.970 185.490 ;
        RECT 113.770 183.790 113.910 185.170 ;
        RECT 113.710 183.470 113.970 183.790 ;
        RECT 114.170 183.470 114.430 183.790 ;
        RECT 114.230 183.190 114.370 183.470 ;
        RECT 111.930 183.050 112.530 183.190 ;
        RECT 111.010 181.410 111.150 182.935 ;
        RECT 111.870 182.450 112.130 182.770 ;
        RECT 111.410 181.430 111.670 181.750 ;
        RECT 110.950 181.090 111.210 181.410 ;
        RECT 110.950 180.410 111.210 180.730 ;
        RECT 111.010 179.030 111.150 180.410 ;
        RECT 111.470 180.390 111.610 181.430 ;
        RECT 111.930 180.730 112.070 182.450 ;
        RECT 111.870 180.410 112.130 180.730 ;
        RECT 111.410 180.070 111.670 180.390 ;
        RECT 110.950 178.710 111.210 179.030 ;
        RECT 111.470 178.010 111.610 180.070 ;
        RECT 111.410 177.690 111.670 178.010 ;
        RECT 110.490 177.350 110.750 177.670 ;
        RECT 111.930 176.310 112.070 180.410 ;
        RECT 111.870 175.990 112.130 176.310 ;
        RECT 111.410 169.530 111.670 169.850 ;
        RECT 110.950 167.830 111.210 168.150 ;
        RECT 110.490 167.380 110.750 167.470 ;
        RECT 110.090 167.240 110.750 167.380 ;
        RECT 110.090 166.450 110.230 167.240 ;
        RECT 110.490 167.150 110.750 167.240 ;
        RECT 110.030 166.130 110.290 166.450 ;
        RECT 110.490 165.110 110.750 165.430 ;
        RECT 110.550 161.350 110.690 165.110 ;
        RECT 111.010 162.030 111.150 167.830 ;
        RECT 111.470 167.665 111.610 169.530 ;
        RECT 111.400 167.295 111.680 167.665 ;
        RECT 112.390 167.470 112.530 183.050 ;
        RECT 112.850 183.050 113.450 183.190 ;
        RECT 113.770 183.110 114.370 183.190 ;
        RECT 113.710 183.050 114.370 183.110 ;
        RECT 112.850 180.730 112.990 183.050 ;
        RECT 113.710 182.790 113.970 183.050 ;
        RECT 113.250 182.450 113.510 182.770 ;
        RECT 114.170 182.450 114.430 182.770 ;
        RECT 112.790 180.410 113.050 180.730 ;
        RECT 112.850 175.970 112.990 180.410 ;
        RECT 113.310 178.010 113.450 182.450 ;
        RECT 113.710 181.430 113.970 181.750 ;
        RECT 113.250 177.690 113.510 178.010 ;
        RECT 112.790 175.650 113.050 175.970 ;
        RECT 112.790 174.970 113.050 175.290 ;
        RECT 112.850 173.590 112.990 174.970 ;
        RECT 112.790 173.270 113.050 173.590 ;
        RECT 112.850 170.385 112.990 173.270 ;
        RECT 113.310 172.310 113.450 177.690 ;
        RECT 113.770 175.630 113.910 181.430 ;
        RECT 114.230 180.730 114.370 182.450 ;
        RECT 114.690 181.410 114.830 185.510 ;
        RECT 114.630 181.090 114.890 181.410 ;
        RECT 114.170 180.410 114.430 180.730 ;
        RECT 114.630 180.410 114.890 180.730 ;
        RECT 114.230 177.670 114.370 180.410 ;
        RECT 114.690 179.905 114.830 180.410 ;
        RECT 114.620 179.535 114.900 179.905 ;
        RECT 114.620 178.855 114.900 179.225 ;
        RECT 114.630 178.710 114.890 178.855 ;
        RECT 114.170 177.350 114.430 177.670 ;
        RECT 114.690 175.970 114.830 178.710 ;
        RECT 114.630 175.650 114.890 175.970 ;
        RECT 113.710 175.310 113.970 175.630 ;
        RECT 114.630 174.970 114.890 175.290 ;
        RECT 114.170 174.290 114.430 174.610 ;
        RECT 113.310 172.170 113.910 172.310 ;
        RECT 113.770 171.890 113.910 172.170 ;
        RECT 113.250 171.570 113.510 171.890 ;
        RECT 113.710 171.570 113.970 171.890 ;
        RECT 112.780 170.015 113.060 170.385 ;
        RECT 111.410 167.150 111.670 167.295 ;
        RECT 112.330 167.150 112.590 167.470 ;
        RECT 112.390 164.750 112.530 167.150 ;
        RECT 112.850 165.430 112.990 170.015 ;
        RECT 112.790 165.110 113.050 165.430 ;
        RECT 112.330 164.430 112.590 164.750 ;
        RECT 112.390 162.030 112.530 164.430 ;
        RECT 112.790 164.090 113.050 164.410 ;
        RECT 112.850 162.110 112.990 164.090 ;
        RECT 113.310 162.710 113.450 171.570 ;
        RECT 113.700 168.655 113.980 169.025 ;
        RECT 113.770 167.130 113.910 168.655 ;
        RECT 113.710 166.810 113.970 167.130 ;
        RECT 113.770 164.070 113.910 166.810 ;
        RECT 114.230 166.450 114.370 174.290 ;
        RECT 114.690 169.170 114.830 174.970 ;
        RECT 115.150 169.850 115.290 187.890 ;
        RECT 115.610 187.190 115.750 192.310 ;
        RECT 116.010 191.290 116.270 191.610 ;
        RECT 116.070 188.890 116.210 191.290 ;
        RECT 116.530 191.270 116.670 196.050 ;
        RECT 124.810 193.390 124.950 196.730 ;
        RECT 124.810 193.250 125.410 193.390 ;
        RECT 118.770 191.970 119.030 192.290 ;
        RECT 116.930 191.290 117.190 191.610 ;
        RECT 116.470 190.950 116.730 191.270 ;
        RECT 116.530 190.785 116.670 190.950 ;
        RECT 116.460 190.415 116.740 190.785 ;
        RECT 116.010 188.570 116.270 188.890 ;
        RECT 115.550 186.870 115.810 187.190 ;
        RECT 115.550 185.740 115.810 186.060 ;
        RECT 115.610 180.390 115.750 185.740 ;
        RECT 116.070 183.450 116.210 188.570 ;
        RECT 116.470 183.700 116.730 183.790 ;
        RECT 116.990 183.700 117.130 191.290 ;
        RECT 117.390 190.610 117.650 190.930 ;
        RECT 117.450 189.910 117.590 190.610 ;
        RECT 117.390 189.590 117.650 189.910 ;
        RECT 117.390 186.870 117.650 187.190 ;
        RECT 117.450 186.490 117.590 186.870 ;
        RECT 118.310 186.490 118.570 186.510 ;
        RECT 118.830 186.490 118.970 191.970 ;
        RECT 125.270 189.230 125.410 193.250 ;
        RECT 133.950 191.290 134.210 191.610 ;
        RECT 137.170 191.290 137.430 191.610 ;
        RECT 134.010 189.230 134.150 191.290 ;
        RECT 135.790 190.610 136.050 190.930 ;
        RECT 135.850 189.230 135.990 190.610 ;
        RECT 125.210 188.910 125.470 189.230 ;
        RECT 129.810 188.910 130.070 189.230 ;
        RECT 133.950 188.910 134.210 189.230 ;
        RECT 135.790 188.910 136.050 189.230 ;
        RECT 125.270 188.630 125.410 188.910 ;
        RECT 125.270 188.490 125.870 188.630 ;
        RECT 117.450 186.350 118.050 186.490 ;
        RECT 117.910 185.910 118.050 186.350 ;
        RECT 118.310 186.350 118.970 186.490 ;
        RECT 118.310 186.190 118.570 186.350 ;
        RECT 117.910 185.770 118.510 185.910 ;
        RECT 117.850 185.170 118.110 185.490 ;
        RECT 117.910 183.790 118.050 185.170 ;
        RECT 116.470 183.560 117.130 183.700 ;
        RECT 116.470 183.470 116.730 183.560 ;
        RECT 116.010 183.130 116.270 183.450 ;
        RECT 116.990 183.110 117.130 183.560 ;
        RECT 117.390 183.470 117.650 183.790 ;
        RECT 117.850 183.470 118.110 183.790 ;
        RECT 116.930 182.790 117.190 183.110 ;
        RECT 116.010 181.090 116.270 181.410 ;
        RECT 115.550 180.070 115.810 180.390 ;
        RECT 116.070 178.350 116.210 181.090 ;
        RECT 116.470 180.585 116.730 180.730 ;
        RECT 116.460 180.215 116.740 180.585 ;
        RECT 116.920 178.855 117.200 179.225 ;
        RECT 116.010 178.030 116.270 178.350 ;
        RECT 116.070 175.290 116.210 178.030 ;
        RECT 116.010 174.970 116.270 175.290 ;
        RECT 116.070 173.250 116.210 174.970 ;
        RECT 116.990 174.610 117.130 178.855 ;
        RECT 117.450 178.350 117.590 183.470 ;
        RECT 117.850 179.905 118.110 180.050 ;
        RECT 117.840 179.535 118.120 179.905 ;
        RECT 117.840 178.855 118.120 179.225 ;
        RECT 117.910 178.430 118.050 178.855 ;
        RECT 118.370 178.430 118.510 185.770 ;
        RECT 118.830 184.470 118.970 186.350 ;
        RECT 121.530 186.190 121.790 186.510 ;
        RECT 125.210 186.190 125.470 186.510 ;
        RECT 119.690 185.170 119.950 185.490 ;
        RECT 118.770 184.150 119.030 184.470 ;
        RECT 118.830 178.690 118.970 184.150 ;
        RECT 119.230 183.810 119.490 184.130 ;
        RECT 119.290 181.750 119.430 183.810 ;
        RECT 119.750 183.305 119.890 185.170 ;
        RECT 119.680 182.935 119.960 183.305 ;
        RECT 119.230 181.430 119.490 181.750 ;
        RECT 119.230 180.070 119.490 180.390 ;
        RECT 117.910 178.350 118.510 178.430 ;
        RECT 118.770 178.370 119.030 178.690 ;
        RECT 117.390 178.030 117.650 178.350 ;
        RECT 117.910 178.290 118.570 178.350 ;
        RECT 118.310 178.030 118.570 178.290 ;
        RECT 117.450 176.310 117.590 178.030 ;
        RECT 118.770 177.690 119.030 178.010 ;
        RECT 117.850 177.350 118.110 177.670 ;
        RECT 117.390 175.990 117.650 176.310 ;
        RECT 116.930 174.290 117.190 174.610 ;
        RECT 116.010 172.930 116.270 173.250 ;
        RECT 117.450 172.910 117.590 175.990 ;
        RECT 117.390 172.590 117.650 172.910 ;
        RECT 115.550 171.570 115.810 171.890 ;
        RECT 115.610 169.850 115.750 171.570 ;
        RECT 115.090 169.705 115.350 169.850 ;
        RECT 115.080 169.335 115.360 169.705 ;
        RECT 115.550 169.530 115.810 169.850 ;
        RECT 114.630 168.850 114.890 169.170 ;
        RECT 115.090 167.150 115.350 167.470 ;
        RECT 114.630 166.470 114.890 166.790 ;
        RECT 114.170 166.130 114.430 166.450 ;
        RECT 114.170 165.110 114.430 165.430 ;
        RECT 114.230 164.070 114.370 165.110 ;
        RECT 113.710 163.750 113.970 164.070 ;
        RECT 114.170 163.750 114.430 164.070 ;
        RECT 113.250 162.390 113.510 162.710 ;
        RECT 110.950 161.710 111.210 162.030 ;
        RECT 111.410 161.710 111.670 162.030 ;
        RECT 112.330 161.710 112.590 162.030 ;
        RECT 112.850 161.970 113.450 162.110 ;
        RECT 114.230 162.030 114.370 163.750 ;
        RECT 114.690 162.710 114.830 166.470 ;
        RECT 114.630 162.390 114.890 162.710 ;
        RECT 110.490 161.030 110.750 161.350 ;
        RECT 109.630 159.250 110.230 159.390 ;
        RECT 109.570 158.650 109.830 158.970 ;
        RECT 109.630 155.570 109.770 158.650 ;
        RECT 109.110 155.250 109.370 155.570 ;
        RECT 109.570 155.250 109.830 155.570 ;
        RECT 101.290 153.210 101.550 153.530 ;
        RECT 108.650 153.210 108.910 153.530 ;
        RECT 109.170 153.190 109.310 155.250 ;
        RECT 109.630 154.210 109.770 155.250 ;
        RECT 109.570 153.890 109.830 154.210 ;
        RECT 100.370 152.870 100.630 153.190 ;
        RECT 109.110 152.870 109.370 153.190 ;
        RECT 100.430 148.090 100.570 152.870 ;
        RECT 100.830 152.530 101.090 152.850 ;
        RECT 100.890 149.110 101.030 152.530 ;
        RECT 110.090 150.810 110.230 159.250 ;
        RECT 110.550 158.970 110.690 161.030 ;
        RECT 110.490 158.650 110.750 158.970 ;
        RECT 111.470 153.530 111.610 161.710 ;
        RECT 113.310 161.690 113.450 161.970 ;
        RECT 114.170 161.710 114.430 162.030 ;
        RECT 113.250 161.370 113.510 161.690 ;
        RECT 111.870 160.690 112.130 161.010 ;
        RECT 112.330 160.690 112.590 161.010 ;
        RECT 111.930 157.270 112.070 160.690 ;
        RECT 112.390 159.310 112.530 160.690 ;
        RECT 112.330 158.990 112.590 159.310 ;
        RECT 112.330 158.310 112.590 158.630 ;
        RECT 111.870 156.950 112.130 157.270 ;
        RECT 112.390 156.590 112.530 158.310 ;
        RECT 113.310 158.290 113.450 161.370 ;
        RECT 114.230 158.630 114.370 161.710 ;
        RECT 114.630 161.370 114.890 161.690 ;
        RECT 114.170 158.310 114.430 158.630 ;
        RECT 113.250 157.970 113.510 158.290 ;
        RECT 112.330 156.270 112.590 156.590 ;
        RECT 114.690 154.550 114.830 161.370 ;
        RECT 114.630 154.230 114.890 154.550 ;
        RECT 111.410 153.210 111.670 153.530 ;
        RECT 112.790 152.530 113.050 152.850 ;
        RECT 110.030 150.490 110.290 150.810 ;
        RECT 100.830 148.790 101.090 149.110 ;
        RECT 109.110 148.790 109.370 149.110 ;
        RECT 100.370 147.770 100.630 148.090 ;
        RECT 100.430 146.390 100.570 147.770 ;
        RECT 100.830 147.430 101.090 147.750 ;
        RECT 100.890 146.390 101.030 147.430 ;
        RECT 102.670 147.090 102.930 147.410 ;
        RECT 106.810 147.090 107.070 147.410 ;
        RECT 102.730 146.390 102.870 147.090 ;
        RECT 106.870 146.390 107.010 147.090 ;
        RECT 100.370 146.070 100.630 146.390 ;
        RECT 100.830 146.070 101.090 146.390 ;
        RECT 102.670 146.070 102.930 146.390 ;
        RECT 106.810 146.070 107.070 146.390 ;
        RECT 108.190 146.070 108.450 146.390 ;
        RECT 105.430 145.390 105.690 145.710 ;
        RECT 104.050 141.650 104.310 141.970 ;
        RECT 104.110 140.950 104.250 141.650 ;
        RECT 105.490 140.950 105.630 145.390 ;
        RECT 107.270 143.010 107.530 143.330 ;
        RECT 104.050 140.630 104.310 140.950 ;
        RECT 105.430 140.630 105.690 140.950 ;
        RECT 107.330 140.270 107.470 143.010 ;
        RECT 105.890 139.950 106.150 140.270 ;
        RECT 106.350 139.950 106.610 140.270 ;
        RECT 107.270 139.950 107.530 140.270 ;
        RECT 103.130 139.610 103.390 139.930 ;
        RECT 105.430 139.610 105.690 139.930 ;
        RECT 103.190 134.490 103.330 139.610 ;
        RECT 104.510 136.210 104.770 136.530 ;
        RECT 104.570 135.510 104.710 136.210 ;
        RECT 104.510 135.190 104.770 135.510 ;
        RECT 104.050 134.510 104.310 134.830 ;
        RECT 102.670 134.170 102.930 134.490 ;
        RECT 103.130 134.170 103.390 134.490 ;
        RECT 100.370 133.490 100.630 133.810 ;
        RECT 99.910 132.470 100.170 132.790 ;
        RECT 100.430 131.770 100.570 133.490 ;
        RECT 102.730 132.450 102.870 134.170 ;
        RECT 102.670 132.130 102.930 132.450 ;
        RECT 100.370 131.450 100.630 131.770 ;
        RECT 102.670 129.070 102.930 129.390 ;
        RECT 99.910 128.730 100.170 129.050 ;
        RECT 97.150 128.050 97.410 128.370 ;
        RECT 97.210 126.330 97.350 128.050 ;
        RECT 99.970 126.330 100.110 128.730 ;
        RECT 102.730 127.350 102.870 129.070 ;
        RECT 103.190 129.050 103.330 134.170 ;
        RECT 104.110 132.790 104.250 134.510 ;
        RECT 104.050 132.470 104.310 132.790 ;
        RECT 103.130 128.730 103.390 129.050 ;
        RECT 102.670 127.030 102.930 127.350 ;
        RECT 97.150 126.010 97.410 126.330 ;
        RECT 99.910 126.010 100.170 126.330 ;
        RECT 101.750 126.010 102.010 126.330 ;
        RECT 96.690 122.610 96.950 122.930 ;
        RECT 96.230 120.910 96.490 121.230 ;
        RECT 95.770 118.530 96.030 118.850 ;
        RECT 96.290 118.510 96.430 120.910 ;
        RECT 101.290 120.230 101.550 120.550 ;
        RECT 101.350 118.850 101.490 120.230 ;
        RECT 97.150 118.530 97.410 118.850 ;
        RECT 99.910 118.760 100.170 118.850 ;
        RECT 101.290 118.760 101.550 118.850 ;
        RECT 99.910 118.620 101.550 118.760 ;
        RECT 99.910 118.530 100.170 118.620 ;
        RECT 101.290 118.530 101.550 118.620 ;
        RECT 96.230 118.190 96.490 118.510 ;
        RECT 96.690 117.510 96.950 117.830 ;
        RECT 96.230 104.930 96.490 105.250 ;
        RECT 96.290 98.790 96.430 104.930 ;
        RECT 96.750 104.910 96.890 117.510 ;
        RECT 97.210 115.450 97.350 118.530 ;
        RECT 99.910 117.910 100.170 118.170 ;
        RECT 101.810 117.910 101.950 126.010 ;
        RECT 102.730 123.950 102.870 127.030 ;
        RECT 104.050 125.330 104.310 125.650 ;
        RECT 104.110 124.290 104.250 125.330 ;
        RECT 104.050 123.970 104.310 124.290 ;
        RECT 102.670 123.630 102.930 123.950 ;
        RECT 102.730 121.910 102.870 123.630 ;
        RECT 104.510 122.950 104.770 123.270 ;
        RECT 102.670 121.590 102.930 121.910 ;
        RECT 102.730 118.170 102.870 121.590 ;
        RECT 104.570 120.890 104.710 122.950 ;
        RECT 104.510 120.570 104.770 120.890 ;
        RECT 103.130 119.890 103.390 120.210 ;
        RECT 103.190 118.510 103.330 119.890 ;
        RECT 103.130 118.190 103.390 118.510 ;
        RECT 99.910 117.850 101.950 117.910 ;
        RECT 102.670 117.850 102.930 118.170 ;
        RECT 99.970 117.770 101.950 117.850 ;
        RECT 98.070 115.810 98.330 116.130 ;
        RECT 97.150 115.130 97.410 115.450 ;
        RECT 98.130 110.010 98.270 115.810 ;
        RECT 101.290 113.090 101.550 113.410 ;
        RECT 100.830 110.370 101.090 110.690 ;
        RECT 100.890 110.010 101.030 110.370 ;
        RECT 101.350 110.010 101.490 113.090 ;
        RECT 101.810 110.010 101.950 117.770 ;
        RECT 104.050 116.150 104.310 116.470 ;
        RECT 103.130 114.450 103.390 114.770 ;
        RECT 103.190 113.750 103.330 114.450 ;
        RECT 103.130 113.430 103.390 113.750 ;
        RECT 102.210 110.030 102.470 110.350 ;
        RECT 103.190 110.260 103.330 113.430 ;
        RECT 104.110 113.070 104.250 116.150 ;
        RECT 103.590 112.750 103.850 113.070 ;
        RECT 104.050 112.750 104.310 113.070 ;
        RECT 104.970 112.750 105.230 113.070 ;
        RECT 103.650 112.585 103.790 112.750 ;
        RECT 103.580 112.215 103.860 112.585 ;
        RECT 103.650 111.030 103.790 112.215 ;
        RECT 104.510 111.730 104.770 112.050 ;
        RECT 103.590 110.710 103.850 111.030 ;
        RECT 102.730 110.120 103.330 110.260 ;
        RECT 98.070 109.690 98.330 110.010 ;
        RECT 100.830 109.690 101.090 110.010 ;
        RECT 101.290 109.690 101.550 110.010 ;
        RECT 101.750 109.690 102.010 110.010 ;
        RECT 97.610 109.010 97.870 109.330 ;
        RECT 96.690 104.590 96.950 104.910 ;
        RECT 97.670 99.130 97.810 109.010 ;
        RECT 99.450 105.270 99.710 105.590 ;
        RECT 98.990 104.250 99.250 104.570 ;
        RECT 99.050 102.530 99.190 104.250 ;
        RECT 98.990 102.210 99.250 102.530 ;
        RECT 98.070 101.870 98.330 102.190 ;
        RECT 98.130 100.150 98.270 101.870 ;
        RECT 98.530 101.530 98.790 101.850 ;
        RECT 98.070 99.830 98.330 100.150 ;
        RECT 97.610 98.810 97.870 99.130 ;
        RECT 96.230 98.470 96.490 98.790 ;
        RECT 95.310 96.430 95.570 96.750 ;
        RECT 95.370 96.265 95.510 96.430 ;
        RECT 96.290 96.410 96.430 98.470 ;
        RECT 98.590 96.750 98.730 101.530 ;
        RECT 99.510 99.810 99.650 105.270 ;
        RECT 102.270 100.150 102.410 110.030 ;
        RECT 102.730 109.670 102.870 110.120 ;
        RECT 103.590 109.920 103.850 110.010 ;
        RECT 103.190 109.780 103.850 109.920 ;
        RECT 102.670 109.350 102.930 109.670 ;
        RECT 103.190 107.290 103.330 109.780 ;
        RECT 103.590 109.690 103.850 109.780 ;
        RECT 104.570 107.970 104.710 111.730 ;
        RECT 105.030 111.030 105.170 112.750 ;
        RECT 104.970 110.710 105.230 111.030 ;
        RECT 104.510 107.650 104.770 107.970 ;
        RECT 103.130 106.970 103.390 107.290 ;
        RECT 103.190 104.910 103.330 106.970 ;
        RECT 104.510 104.930 104.770 105.250 ;
        RECT 103.130 104.590 103.390 104.910 ;
        RECT 102.210 99.830 102.470 100.150 ;
        RECT 99.450 99.490 99.710 99.810 ;
        RECT 102.270 99.130 102.410 99.830 ;
        RECT 102.210 98.810 102.470 99.130 ;
        RECT 102.670 98.810 102.930 99.130 ;
        RECT 102.270 97.090 102.410 98.810 ;
        RECT 102.210 96.770 102.470 97.090 ;
        RECT 98.530 96.430 98.790 96.750 ;
        RECT 95.300 95.895 95.580 96.265 ;
        RECT 96.230 96.090 96.490 96.410 ;
        RECT 96.690 95.410 96.950 95.730 ;
        RECT 96.750 93.350 96.890 95.410 ;
        RECT 98.590 93.690 98.730 96.430 ;
        RECT 102.730 94.710 102.870 98.810 ;
        RECT 104.050 96.430 104.310 96.750 ;
        RECT 104.110 94.710 104.250 96.430 ;
        RECT 102.670 94.390 102.930 94.710 ;
        RECT 104.050 94.390 104.310 94.710 ;
        RECT 101.290 94.050 101.550 94.370 ;
        RECT 98.530 93.370 98.790 93.690 ;
        RECT 96.690 93.030 96.950 93.350 ;
        RECT 96.230 92.690 96.490 93.010 ;
        RECT 94.390 90.990 94.650 91.310 ;
        RECT 94.850 90.990 95.110 91.310 ;
        RECT 94.450 90.630 94.590 90.990 ;
        RECT 94.390 90.310 94.650 90.630 ;
        RECT 96.290 89.890 96.430 92.690 ;
        RECT 101.350 91.650 101.490 94.050 ;
        RECT 104.570 94.030 104.710 104.930 ;
        RECT 104.970 102.550 105.230 102.870 ;
        RECT 105.030 99.130 105.170 102.550 ;
        RECT 105.490 100.230 105.630 139.610 ;
        RECT 105.950 138.230 106.090 139.950 ;
        RECT 105.890 137.910 106.150 138.230 ;
        RECT 106.410 137.210 106.550 139.950 ;
        RECT 106.810 137.230 107.070 137.550 ;
        RECT 106.350 136.890 106.610 137.210 ;
        RECT 106.870 126.670 107.010 137.230 ;
        RECT 107.270 134.510 107.530 134.830 ;
        RECT 107.330 132.790 107.470 134.510 ;
        RECT 107.270 132.470 107.530 132.790 ;
        RECT 108.250 130.070 108.390 146.070 ;
        RECT 108.650 145.390 108.910 145.710 ;
        RECT 108.710 138.230 108.850 145.390 ;
        RECT 109.170 142.650 109.310 148.790 ;
        RECT 111.870 148.450 112.130 148.770 ;
        RECT 110.030 147.430 110.290 147.750 ;
        RECT 109.570 145.390 109.830 145.710 ;
        RECT 109.630 143.670 109.770 145.390 ;
        RECT 110.090 144.690 110.230 147.430 ;
        RECT 111.410 147.090 111.670 147.410 ;
        RECT 110.030 144.370 110.290 144.690 ;
        RECT 109.570 143.350 109.830 143.670 ;
        RECT 109.110 142.330 109.370 142.650 ;
        RECT 110.090 140.270 110.230 144.370 ;
        RECT 111.470 143.070 111.610 147.090 ;
        RECT 111.930 143.670 112.070 148.450 ;
        RECT 112.330 145.390 112.590 145.710 ;
        RECT 111.870 143.350 112.130 143.670 ;
        RECT 110.550 142.930 112.070 143.070 ;
        RECT 112.390 142.990 112.530 145.390 ;
        RECT 110.550 142.650 110.690 142.930 ;
        RECT 110.490 142.330 110.750 142.650 ;
        RECT 110.030 139.950 110.290 140.270 ;
        RECT 108.650 137.910 108.910 138.230 ;
        RECT 110.550 138.190 110.690 142.330 ;
        RECT 111.930 140.270 112.070 142.930 ;
        RECT 112.330 142.670 112.590 142.990 ;
        RECT 111.870 139.950 112.130 140.270 ;
        RECT 111.410 138.930 111.670 139.250 ;
        RECT 112.850 138.990 112.990 152.530 ;
        RECT 115.150 151.150 115.290 167.150 ;
        RECT 115.610 164.410 115.750 169.530 ;
        RECT 116.460 169.335 116.740 169.705 ;
        RECT 116.010 168.850 116.270 169.170 ;
        RECT 116.070 167.470 116.210 168.850 ;
        RECT 116.010 167.150 116.270 167.470 ;
        RECT 116.010 166.130 116.270 166.450 ;
        RECT 116.070 164.750 116.210 166.130 ;
        RECT 116.010 164.430 116.270 164.750 ;
        RECT 115.550 164.090 115.810 164.410 ;
        RECT 116.070 162.030 116.210 164.430 ;
        RECT 116.530 164.410 116.670 169.335 ;
        RECT 116.930 168.850 117.190 169.170 ;
        RECT 117.450 169.080 117.590 172.590 ;
        RECT 117.910 171.890 118.050 177.350 ;
        RECT 118.830 176.310 118.970 177.690 ;
        RECT 118.770 175.990 119.030 176.310 ;
        RECT 118.310 174.970 118.570 175.290 ;
        RECT 118.370 172.990 118.510 174.970 ;
        RECT 118.830 173.590 118.970 175.990 ;
        RECT 119.290 175.290 119.430 180.070 ;
        RECT 119.750 178.260 119.890 182.935 ;
        RECT 120.610 182.450 120.870 182.770 ;
        RECT 120.670 180.390 120.810 182.450 ;
        RECT 120.610 180.070 120.870 180.390 ;
        RECT 121.070 179.730 121.330 180.050 ;
        RECT 120.150 178.260 120.410 178.350 ;
        RECT 119.750 178.120 120.810 178.260 ;
        RECT 120.150 178.030 120.410 178.120 ;
        RECT 120.150 175.310 120.410 175.630 ;
        RECT 119.230 174.970 119.490 175.290 ;
        RECT 119.690 174.630 119.950 174.950 ;
        RECT 118.770 173.270 119.030 173.590 ;
        RECT 118.370 172.850 118.970 172.990 ;
        RECT 118.310 171.910 118.570 172.230 ;
        RECT 117.850 171.570 118.110 171.890 ;
        RECT 117.850 169.870 118.110 170.190 ;
        RECT 117.910 169.705 118.050 169.870 ;
        RECT 117.840 169.335 118.120 169.705 ;
        RECT 117.850 169.080 118.110 169.170 ;
        RECT 117.450 169.025 118.110 169.080 ;
        RECT 117.380 168.940 118.110 169.025 ;
        RECT 116.990 168.150 117.130 168.850 ;
        RECT 117.380 168.655 117.660 168.940 ;
        RECT 117.850 168.850 118.110 168.940 ;
        RECT 116.930 167.830 117.190 168.150 ;
        RECT 116.990 167.470 117.130 167.830 ;
        RECT 116.930 167.150 117.190 167.470 ;
        RECT 117.390 166.470 117.650 166.790 ;
        RECT 117.450 164.410 117.590 166.470 ;
        RECT 118.370 166.450 118.510 171.910 ;
        RECT 118.830 169.510 118.970 172.850 ;
        RECT 119.750 170.950 119.890 174.630 ;
        RECT 120.210 173.590 120.350 175.310 ;
        RECT 120.670 175.290 120.810 178.120 ;
        RECT 120.610 174.970 120.870 175.290 ;
        RECT 120.150 173.270 120.410 173.590 ;
        RECT 120.610 171.570 120.870 171.890 ;
        RECT 119.750 170.870 120.350 170.950 ;
        RECT 119.750 170.810 120.410 170.870 ;
        RECT 120.150 170.550 120.410 170.810 ;
        RECT 119.220 170.015 119.500 170.385 ;
        RECT 119.290 169.850 119.430 170.015 ;
        RECT 119.230 169.530 119.490 169.850 ;
        RECT 119.690 169.530 119.950 169.850 ;
        RECT 118.770 169.190 119.030 169.510 ;
        RECT 118.310 166.130 118.570 166.450 ;
        RECT 116.470 164.090 116.730 164.410 ;
        RECT 117.390 164.320 117.650 164.410 ;
        RECT 117.390 164.180 118.050 164.320 ;
        RECT 117.390 164.090 117.650 164.180 ;
        RECT 117.390 163.410 117.650 163.730 ;
        RECT 116.010 161.710 116.270 162.030 ;
        RECT 116.930 160.690 117.190 161.010 ;
        RECT 116.990 158.970 117.130 160.690 ;
        RECT 116.930 158.650 117.190 158.970 ;
        RECT 117.450 158.630 117.590 163.410 ;
        RECT 117.910 162.030 118.050 164.180 ;
        RECT 118.310 162.390 118.570 162.710 ;
        RECT 117.850 161.710 118.110 162.030 ;
        RECT 117.390 158.310 117.650 158.630 ;
        RECT 115.550 157.970 115.810 158.290 ;
        RECT 116.470 157.970 116.730 158.290 ;
        RECT 115.610 156.590 115.750 157.970 ;
        RECT 115.550 156.270 115.810 156.590 ;
        RECT 116.530 156.250 116.670 157.970 ;
        RECT 117.910 156.590 118.050 161.710 ;
        RECT 118.370 159.650 118.510 162.390 ;
        RECT 118.830 161.350 118.970 169.190 ;
        RECT 119.230 167.150 119.490 167.470 ;
        RECT 119.290 165.090 119.430 167.150 ;
        RECT 119.230 164.770 119.490 165.090 ;
        RECT 119.290 162.370 119.430 164.770 ;
        RECT 119.750 162.710 119.890 169.530 ;
        RECT 119.690 162.390 119.950 162.710 ;
        RECT 119.230 162.050 119.490 162.370 ;
        RECT 118.770 161.030 119.030 161.350 ;
        RECT 120.210 161.010 120.350 170.550 ;
        RECT 120.670 170.530 120.810 171.570 ;
        RECT 120.610 170.210 120.870 170.530 ;
        RECT 120.150 160.690 120.410 161.010 ;
        RECT 118.310 159.330 118.570 159.650 ;
        RECT 121.130 159.390 121.270 179.730 ;
        RECT 121.590 167.470 121.730 186.190 ;
        RECT 125.270 184.550 125.410 186.190 ;
        RECT 124.810 184.470 125.410 184.550 ;
        RECT 124.750 184.410 125.410 184.470 ;
        RECT 124.750 184.150 125.010 184.410 ;
        RECT 125.730 183.790 125.870 188.490 ;
        RECT 129.870 187.190 130.010 188.910 ;
        RECT 131.650 188.570 131.910 188.890 ;
        RECT 137.230 188.745 137.370 191.290 ;
        RECT 129.810 186.870 130.070 187.190 ;
        RECT 131.710 186.170 131.850 188.570 ;
        RECT 137.160 188.375 137.440 188.745 ;
        RECT 136.710 187.890 136.970 188.210 ;
        RECT 131.650 185.850 131.910 186.170 ;
        RECT 135.790 185.850 136.050 186.170 ;
        RECT 126.130 185.510 126.390 185.830 ;
        RECT 123.830 183.470 124.090 183.790 ;
        RECT 125.670 183.470 125.930 183.790 ;
        RECT 122.450 183.130 122.710 183.450 ;
        RECT 122.510 180.730 122.650 183.130 ;
        RECT 123.890 180.730 124.030 183.470 ;
        RECT 126.190 183.110 126.330 185.510 ;
        RECT 127.510 185.170 127.770 185.490 ;
        RECT 134.870 185.170 135.130 185.490 ;
        RECT 126.590 183.470 126.850 183.790 ;
        RECT 126.130 182.790 126.390 183.110 ;
        RECT 126.650 181.070 126.790 183.470 ;
        RECT 127.570 181.750 127.710 185.170 ;
        RECT 127.970 183.470 128.230 183.790 ;
        RECT 128.030 181.750 128.170 183.470 ;
        RECT 133.950 182.450 134.210 182.770 ;
        RECT 127.510 181.430 127.770 181.750 ;
        RECT 127.970 181.430 128.230 181.750 ;
        RECT 126.590 180.750 126.850 181.070 ;
        RECT 122.450 180.410 122.710 180.730 ;
        RECT 123.830 180.410 124.090 180.730 ;
        RECT 122.510 179.030 122.650 180.410 ;
        RECT 123.890 179.960 124.030 180.410 ;
        RECT 123.430 179.820 124.030 179.960 ;
        RECT 123.430 179.030 123.570 179.820 ;
        RECT 126.130 179.730 126.390 180.050 ;
        RECT 126.190 179.030 126.330 179.730 ;
        RECT 122.450 178.710 122.710 179.030 ;
        RECT 123.370 178.710 123.630 179.030 ;
        RECT 126.130 178.710 126.390 179.030 ;
        RECT 121.990 177.690 122.250 178.010 ;
        RECT 121.530 167.150 121.790 167.470 ;
        RECT 121.590 166.790 121.730 167.150 ;
        RECT 121.530 166.470 121.790 166.790 ;
        RECT 120.210 159.250 121.270 159.390 ;
        RECT 117.850 156.270 118.110 156.590 ;
        RECT 118.310 156.270 118.570 156.590 ;
        RECT 116.470 155.930 116.730 156.250 ;
        RECT 116.530 153.870 116.670 155.930 ;
        RECT 116.470 153.550 116.730 153.870 ;
        RECT 117.380 153.695 117.660 154.065 ;
        RECT 117.450 153.530 117.590 153.695 ;
        RECT 117.390 153.210 117.650 153.530 ;
        RECT 117.910 151.830 118.050 156.270 ;
        RECT 117.850 151.510 118.110 151.830 ;
        RECT 118.370 151.490 118.510 156.270 ;
        RECT 118.310 151.170 118.570 151.490 ;
        RECT 115.090 150.830 115.350 151.150 ;
        RECT 116.470 149.810 116.730 150.130 ;
        RECT 113.250 147.770 113.510 148.090 ;
        RECT 113.310 146.390 113.450 147.770 ;
        RECT 114.630 147.090 114.890 147.410 ;
        RECT 114.690 146.390 114.830 147.090 ;
        RECT 113.250 146.070 113.510 146.390 ;
        RECT 114.630 146.070 114.890 146.390 ;
        RECT 116.000 145.535 116.280 145.905 ;
        RECT 116.010 145.390 116.270 145.535 ;
        RECT 116.530 145.030 116.670 149.810 ;
        RECT 118.770 148.790 119.030 149.110 ;
        RECT 116.930 147.430 117.190 147.750 ;
        RECT 115.090 144.710 115.350 145.030 ;
        RECT 116.470 144.710 116.730 145.030 ;
        RECT 113.250 143.350 113.510 143.670 ;
        RECT 110.550 138.050 111.150 138.190 ;
        RECT 109.170 137.550 110.690 137.630 ;
        RECT 109.110 137.490 110.690 137.550 ;
        RECT 109.110 137.230 109.370 137.490 ;
        RECT 110.550 137.210 110.690 137.490 ;
        RECT 109.570 136.890 109.830 137.210 ;
        RECT 110.490 136.890 110.750 137.210 ;
        RECT 108.650 136.210 108.910 136.530 ;
        RECT 108.710 134.830 108.850 136.210 ;
        RECT 108.650 134.510 108.910 134.830 ;
        RECT 108.190 129.750 108.450 130.070 ;
        RECT 107.730 128.390 107.990 128.710 ;
        RECT 106.810 126.350 107.070 126.670 ;
        RECT 107.790 122.930 107.930 128.390 ;
        RECT 108.190 123.970 108.450 124.290 ;
        RECT 107.730 122.610 107.990 122.930 ;
        RECT 105.890 120.910 106.150 121.230 ;
        RECT 105.950 118.510 106.090 120.910 ;
        RECT 105.890 118.190 106.150 118.510 ;
        RECT 107.790 115.190 107.930 122.610 ;
        RECT 108.250 118.510 108.390 123.970 ;
        RECT 108.710 123.950 108.850 134.510 ;
        RECT 109.110 131.450 109.370 131.770 ;
        RECT 109.170 128.710 109.310 131.450 ;
        RECT 109.110 128.390 109.370 128.710 ;
        RECT 108.650 123.630 108.910 123.950 ;
        RECT 109.110 118.870 109.370 119.190 ;
        RECT 108.190 118.190 108.450 118.510 ;
        RECT 108.250 115.790 108.390 118.190 ;
        RECT 108.190 115.470 108.450 115.790 ;
        RECT 107.790 115.050 108.390 115.190 ;
        RECT 106.810 112.750 107.070 113.070 ;
        RECT 106.870 107.630 107.010 112.750 ;
        RECT 107.730 112.070 107.990 112.390 ;
        RECT 106.810 107.310 107.070 107.630 ;
        RECT 106.870 106.610 107.010 107.310 ;
        RECT 106.810 106.290 107.070 106.610 ;
        RECT 107.790 101.170 107.930 112.070 ;
        RECT 107.730 100.850 107.990 101.170 ;
        RECT 108.250 100.230 108.390 115.050 ;
        RECT 109.170 107.290 109.310 118.870 ;
        RECT 109.110 106.970 109.370 107.290 ;
        RECT 109.170 104.570 109.310 106.970 ;
        RECT 109.110 104.480 109.370 104.570 ;
        RECT 108.710 104.340 109.370 104.480 ;
        RECT 108.710 102.190 108.850 104.340 ;
        RECT 109.110 104.250 109.370 104.340 ;
        RECT 108.650 101.870 108.910 102.190 ;
        RECT 109.110 101.870 109.370 102.190 ;
        RECT 105.490 100.090 107.470 100.230 ;
        RECT 104.970 98.810 105.230 99.130 ;
        RECT 105.430 98.470 105.690 98.790 ;
        RECT 104.970 98.130 105.230 98.450 ;
        RECT 105.030 96.410 105.170 98.130 ;
        RECT 104.970 96.090 105.230 96.410 ;
        RECT 105.030 94.030 105.170 96.090 ;
        RECT 104.510 93.710 104.770 94.030 ;
        RECT 104.970 93.710 105.230 94.030 ;
        RECT 101.750 93.030 102.010 93.350 ;
        RECT 104.510 93.030 104.770 93.350 ;
        RECT 99.450 91.330 99.710 91.650 ;
        RECT 101.290 91.330 101.550 91.650 ;
        RECT 97.150 90.990 97.410 91.310 ;
        RECT 97.210 89.890 97.350 90.990 ;
        RECT 96.290 89.750 96.890 89.890 ;
        RECT 97.210 89.750 97.810 89.890 ;
        RECT 96.750 88.250 96.890 89.750 ;
        RECT 97.670 88.590 97.810 89.750 ;
        RECT 97.610 88.270 97.870 88.590 ;
        RECT 99.510 88.250 99.650 91.330 ;
        RECT 101.810 91.310 101.950 93.030 ;
        RECT 101.750 90.990 102.010 91.310 ;
        RECT 104.570 90.290 104.710 93.030 ;
        RECT 104.970 92.865 105.230 93.010 ;
        RECT 104.960 92.495 105.240 92.865 ;
        RECT 105.490 91.310 105.630 98.470 ;
        RECT 105.890 97.110 106.150 97.430 ;
        RECT 105.950 91.990 106.090 97.110 ;
        RECT 106.810 96.770 107.070 97.090 ;
        RECT 106.350 95.750 106.610 96.070 ;
        RECT 106.410 94.225 106.550 95.750 ;
        RECT 106.340 93.855 106.620 94.225 ;
        RECT 106.870 94.030 107.010 96.770 ;
        RECT 106.810 93.710 107.070 94.030 ;
        RECT 106.350 93.430 106.610 93.690 ;
        RECT 106.350 93.370 107.010 93.430 ;
        RECT 106.410 93.290 107.010 93.370 ;
        RECT 105.890 91.670 106.150 91.990 ;
        RECT 106.340 91.815 106.620 92.185 ;
        RECT 106.870 91.990 107.010 93.290 ;
        RECT 107.330 91.990 107.470 100.090 ;
        RECT 107.790 100.090 108.390 100.230 ;
        RECT 106.410 91.310 106.550 91.815 ;
        RECT 106.810 91.670 107.070 91.990 ;
        RECT 107.270 91.670 107.530 91.990 ;
        RECT 107.790 91.390 107.930 100.090 ;
        RECT 108.710 97.430 108.850 101.870 ;
        RECT 109.170 99.130 109.310 101.870 ;
        RECT 109.110 98.810 109.370 99.130 ;
        RECT 108.650 97.340 108.910 97.430 ;
        RECT 108.650 97.200 109.310 97.340 ;
        RECT 108.650 97.110 108.910 97.200 ;
        RECT 108.190 96.430 108.450 96.750 ;
        RECT 108.640 96.575 108.920 96.945 ;
        RECT 105.430 90.990 105.690 91.310 ;
        RECT 106.350 90.990 106.610 91.310 ;
        RECT 107.330 91.250 107.930 91.390 ;
        RECT 100.830 89.970 101.090 90.290 ;
        RECT 104.510 89.970 104.770 90.290 ;
        RECT 100.890 89.270 101.030 89.970 ;
        RECT 105.490 89.890 105.630 90.990 ;
        RECT 105.030 89.750 105.630 89.890 ;
        RECT 100.830 88.950 101.090 89.270 ;
        RECT 100.890 88.250 101.030 88.950 ;
        RECT 101.290 88.610 101.550 88.930 ;
        RECT 59.430 87.930 59.690 88.250 ;
        RECT 67.710 87.930 67.970 88.250 ;
        RECT 69.090 87.930 69.350 88.250 ;
        RECT 76.910 87.930 77.170 88.250 ;
        RECT 77.370 87.930 77.630 88.250 ;
        RECT 77.830 87.930 78.090 88.250 ;
        RECT 83.810 87.930 84.070 88.250 ;
        RECT 88.410 87.930 88.670 88.250 ;
        RECT 92.090 87.930 92.350 88.250 ;
        RECT 93.930 87.930 94.190 88.250 ;
        RECT 96.690 87.930 96.950 88.250 ;
        RECT 99.450 87.930 99.710 88.250 ;
        RECT 100.830 87.930 101.090 88.250 ;
        RECT 32.180 86.715 33.720 87.085 ;
        RECT 59.490 80.020 59.630 87.930 ;
        RECT 65.870 87.250 66.130 87.570 ;
        RECT 65.930 80.020 66.070 87.250 ;
        RECT 69.150 80.020 69.290 87.930 ;
        RECT 72.310 87.250 72.570 87.570 ;
        RECT 75.530 87.250 75.790 87.570 ;
        RECT 78.750 87.250 79.010 87.570 ;
        RECT 81.970 87.250 82.230 87.570 ;
        RECT 85.190 87.250 85.450 87.570 ;
        RECT 88.410 87.250 88.670 87.570 ;
        RECT 91.630 87.250 91.890 87.570 ;
        RECT 94.850 87.250 95.110 87.570 ;
        RECT 98.070 87.250 98.330 87.570 ;
        RECT 72.370 80.020 72.510 87.250 ;
        RECT 75.590 80.020 75.730 87.250 ;
        RECT 78.810 80.020 78.950 87.250 ;
        RECT 82.030 80.020 82.170 87.250 ;
        RECT 85.250 80.020 85.390 87.250 ;
        RECT 88.470 80.020 88.610 87.250 ;
        RECT 91.690 80.020 91.830 87.250 ;
        RECT 94.910 80.020 95.050 87.250 ;
        RECT 98.130 80.020 98.270 87.250 ;
        RECT 101.350 80.020 101.490 88.610 ;
        RECT 105.030 88.590 105.170 89.750 ;
        RECT 104.970 88.270 105.230 88.590 ;
        RECT 106.410 88.250 106.550 90.990 ;
        RECT 107.330 90.290 107.470 91.250 ;
        RECT 107.270 89.970 107.530 90.290 ;
        RECT 106.350 87.930 106.610 88.250 ;
        RECT 108.250 87.910 108.390 96.430 ;
        RECT 108.710 93.690 108.850 96.575 ;
        RECT 108.650 93.370 108.910 93.690 ;
        RECT 109.170 93.010 109.310 97.200 ;
        RECT 109.630 93.010 109.770 136.890 ;
        RECT 110.030 136.210 110.290 136.530 ;
        RECT 110.090 131.770 110.230 136.210 ;
        RECT 110.550 133.810 110.690 136.890 ;
        RECT 110.490 133.490 110.750 133.810 ;
        RECT 110.550 132.110 110.690 133.490 ;
        RECT 110.490 131.790 110.750 132.110 ;
        RECT 110.030 131.450 110.290 131.770 ;
        RECT 110.030 122.610 110.290 122.930 ;
        RECT 110.090 120.890 110.230 122.610 ;
        RECT 110.550 121.230 110.690 131.790 ;
        RECT 111.010 131.090 111.150 138.050 ;
        RECT 111.470 137.890 111.610 138.930 ;
        RECT 111.930 138.850 112.990 138.990 ;
        RECT 111.410 137.570 111.670 137.890 ;
        RECT 111.410 133.830 111.670 134.150 ;
        RECT 110.950 130.770 111.210 131.090 ;
        RECT 110.950 126.010 111.210 126.330 ;
        RECT 111.010 123.610 111.150 126.010 ;
        RECT 110.950 123.290 111.210 123.610 ;
        RECT 111.470 121.310 111.610 133.830 ;
        RECT 111.930 122.930 112.070 138.850 ;
        RECT 113.310 138.190 113.450 143.350 ;
        RECT 113.710 141.990 113.970 142.310 ;
        RECT 113.770 140.950 113.910 141.990 ;
        RECT 114.170 141.650 114.430 141.970 ;
        RECT 114.230 140.950 114.370 141.650 ;
        RECT 113.710 140.630 113.970 140.950 ;
        RECT 114.170 140.630 114.430 140.950 ;
        RECT 115.150 140.270 115.290 144.710 ;
        RECT 115.550 144.370 115.810 144.690 ;
        RECT 115.610 143.670 115.750 144.370 ;
        RECT 115.550 143.350 115.810 143.670 ;
        RECT 115.610 142.650 115.750 143.350 ;
        RECT 115.550 142.330 115.810 142.650 ;
        RECT 116.990 142.310 117.130 147.430 ;
        RECT 117.390 145.390 117.650 145.710 ;
        RECT 117.450 143.670 117.590 145.390 ;
        RECT 117.390 143.350 117.650 143.670 ;
        RECT 116.930 141.990 117.190 142.310 ;
        RECT 116.990 140.350 117.130 141.990 ;
        RECT 118.310 141.650 118.570 141.970 ;
        RECT 116.070 140.270 117.130 140.350 ;
        RECT 113.710 139.950 113.970 140.270 ;
        RECT 115.090 139.950 115.350 140.270 ;
        RECT 116.010 140.210 117.130 140.270 ;
        RECT 116.010 139.950 116.270 140.210 ;
        RECT 112.850 138.050 113.450 138.190 ;
        RECT 113.770 138.190 113.910 139.950 ;
        RECT 113.770 138.050 114.370 138.190 ;
        RECT 112.330 134.850 112.590 135.170 ;
        RECT 112.390 126.670 112.530 134.850 ;
        RECT 112.850 131.090 112.990 138.050 ;
        RECT 113.250 136.890 113.510 137.210 ;
        RECT 112.790 130.770 113.050 131.090 ;
        RECT 112.790 128.050 113.050 128.370 ;
        RECT 112.330 126.350 112.590 126.670 ;
        RECT 111.870 122.610 112.130 122.930 ;
        RECT 110.490 120.910 110.750 121.230 ;
        RECT 111.010 121.170 111.610 121.310 ;
        RECT 112.390 121.230 112.530 126.350 ;
        RECT 112.850 126.330 112.990 128.050 ;
        RECT 112.790 126.010 113.050 126.330 ;
        RECT 110.030 120.570 110.290 120.890 ;
        RECT 110.090 113.410 110.230 120.570 ;
        RECT 111.010 116.130 111.150 121.170 ;
        RECT 112.330 120.910 112.590 121.230 ;
        RECT 111.410 120.570 111.670 120.890 ;
        RECT 111.470 119.190 111.610 120.570 ;
        RECT 111.410 118.870 111.670 119.190 ;
        RECT 112.390 118.850 112.530 120.910 ;
        RECT 112.790 118.870 113.050 119.190 ;
        RECT 112.330 118.760 112.590 118.850 ;
        RECT 111.930 118.620 112.590 118.760 ;
        RECT 111.410 117.170 111.670 117.490 ;
        RECT 110.950 115.810 111.210 116.130 ;
        RECT 110.030 113.090 110.290 113.410 ;
        RECT 110.490 112.750 110.750 113.070 ;
        RECT 110.550 106.950 110.690 112.750 ;
        RECT 110.950 111.790 111.210 112.050 ;
        RECT 111.470 111.790 111.610 117.170 ;
        RECT 111.930 115.450 112.070 118.620 ;
        RECT 112.330 118.530 112.590 118.620 ;
        RECT 112.850 117.830 112.990 118.870 ;
        RECT 112.790 117.510 113.050 117.830 ;
        RECT 112.330 116.150 112.590 116.470 ;
        RECT 111.870 115.130 112.130 115.450 ;
        RECT 111.870 112.750 112.130 113.070 ;
        RECT 110.950 111.730 111.610 111.790 ;
        RECT 111.010 111.650 111.610 111.730 ;
        RECT 111.410 109.010 111.670 109.330 ;
        RECT 110.490 106.630 110.750 106.950 ;
        RECT 110.550 105.250 110.690 106.630 ;
        RECT 110.490 104.930 110.750 105.250 ;
        RECT 110.030 101.870 110.290 102.190 ;
        RECT 110.090 96.750 110.230 101.870 ;
        RECT 110.490 101.190 110.750 101.510 ;
        RECT 110.550 97.090 110.690 101.190 ;
        RECT 110.490 96.945 110.750 97.090 ;
        RECT 110.480 96.830 110.760 96.945 ;
        RECT 110.030 96.430 110.290 96.750 ;
        RECT 110.480 96.690 111.150 96.830 ;
        RECT 110.480 96.575 110.760 96.690 ;
        RECT 110.490 96.090 110.750 96.410 ;
        RECT 110.030 95.750 110.290 96.070 ;
        RECT 109.110 92.690 109.370 93.010 ;
        RECT 109.570 92.690 109.830 93.010 ;
        RECT 108.640 91.815 108.920 92.185 ;
        RECT 108.710 90.970 108.850 91.815 ;
        RECT 109.170 91.310 109.310 92.690 ;
        RECT 109.570 91.670 109.830 91.990 ;
        RECT 109.110 90.990 109.370 91.310 ;
        RECT 108.650 90.650 108.910 90.970 ;
        RECT 109.630 88.930 109.770 91.670 ;
        RECT 109.570 88.610 109.830 88.930 ;
        RECT 110.090 88.250 110.230 95.750 ;
        RECT 110.550 94.225 110.690 96.090 ;
        RECT 110.480 93.855 110.760 94.225 ;
        RECT 110.490 93.370 110.750 93.690 ;
        RECT 110.550 90.290 110.690 93.370 ;
        RECT 111.010 91.650 111.150 96.690 ;
        RECT 110.950 91.330 111.210 91.650 ;
        RECT 111.010 90.825 111.150 91.330 ;
        RECT 110.940 90.455 111.220 90.825 ;
        RECT 110.490 89.970 110.750 90.290 ;
        RECT 111.470 88.250 111.610 109.010 ;
        RECT 111.930 107.030 112.070 112.750 ;
        RECT 112.390 112.640 112.530 116.150 ;
        RECT 112.790 114.790 113.050 115.110 ;
        RECT 112.850 113.750 112.990 114.790 ;
        RECT 112.790 113.430 113.050 113.750 ;
        RECT 112.790 112.640 113.050 112.730 ;
        RECT 112.390 112.500 113.050 112.640 ;
        RECT 112.790 112.410 113.050 112.500 ;
        RECT 112.330 111.730 112.590 112.050 ;
        RECT 112.390 110.010 112.530 111.730 ;
        RECT 112.850 110.010 112.990 112.410 ;
        RECT 112.330 109.690 112.590 110.010 ;
        RECT 112.790 109.690 113.050 110.010 ;
        RECT 111.930 106.890 112.990 107.030 ;
        RECT 112.330 106.290 112.590 106.610 ;
        RECT 111.870 103.910 112.130 104.230 ;
        RECT 111.930 102.530 112.070 103.910 ;
        RECT 111.870 102.210 112.130 102.530 ;
        RECT 112.390 101.590 112.530 106.290 ;
        RECT 112.850 102.870 112.990 106.890 ;
        RECT 112.790 102.550 113.050 102.870 ;
        RECT 111.930 101.450 112.530 101.590 ;
        RECT 111.930 89.890 112.070 101.450 ;
        RECT 112.850 100.150 112.990 102.550 ;
        RECT 112.790 99.830 113.050 100.150 ;
        RECT 112.320 92.495 112.600 92.865 ;
        RECT 112.390 91.310 112.530 92.495 ;
        RECT 113.310 91.990 113.450 136.890 ;
        RECT 113.710 131.450 113.970 131.770 ;
        RECT 113.770 95.730 113.910 131.450 ;
        RECT 114.230 125.650 114.370 138.050 ;
        RECT 115.150 137.890 115.290 139.950 ;
        RECT 114.620 137.375 114.900 137.745 ;
        RECT 115.090 137.570 115.350 137.890 ;
        RECT 114.690 137.210 114.830 137.375 ;
        RECT 116.990 137.210 117.130 140.210 ;
        RECT 117.850 139.610 118.110 139.930 ;
        RECT 114.630 136.890 114.890 137.210 ;
        RECT 114.690 135.510 114.830 136.890 ;
        RECT 116.000 136.695 116.280 137.065 ;
        RECT 116.930 136.890 117.190 137.210 ;
        RECT 114.630 135.190 114.890 135.510 ;
        RECT 114.690 132.110 114.830 135.190 ;
        RECT 114.630 131.790 114.890 132.110 ;
        RECT 115.090 131.450 115.350 131.770 ;
        RECT 115.550 131.450 115.810 131.770 ;
        RECT 115.150 127.260 115.290 131.450 ;
        RECT 115.610 130.070 115.750 131.450 ;
        RECT 115.550 129.750 115.810 130.070 ;
        RECT 115.550 127.260 115.810 127.350 ;
        RECT 115.150 127.120 115.810 127.260 ;
        RECT 115.550 127.030 115.810 127.120 ;
        RECT 114.170 125.330 114.430 125.650 ;
        RECT 115.550 119.890 115.810 120.210 ;
        RECT 115.610 118.510 115.750 119.890 ;
        RECT 114.630 118.420 114.890 118.510 ;
        RECT 114.230 118.280 114.890 118.420 ;
        RECT 114.230 114.770 114.370 118.280 ;
        RECT 114.630 118.190 114.890 118.280 ;
        RECT 115.550 118.190 115.810 118.510 ;
        RECT 114.170 114.450 114.430 114.770 ;
        RECT 114.230 110.010 114.370 114.450 ;
        RECT 115.090 112.750 115.350 113.070 ;
        RECT 115.150 110.350 115.290 112.750 ;
        RECT 115.610 111.030 115.750 118.190 ;
        RECT 115.550 110.710 115.810 111.030 ;
        RECT 116.070 110.590 116.210 136.695 ;
        RECT 116.990 134.150 117.130 136.890 ;
        RECT 117.390 134.510 117.650 134.830 ;
        RECT 116.930 133.830 117.190 134.150 ;
        RECT 117.450 132.790 117.590 134.510 ;
        RECT 117.390 132.470 117.650 132.790 ;
        RECT 116.930 131.110 117.190 131.430 ;
        RECT 116.990 128.280 117.130 131.110 ;
        RECT 117.390 128.960 117.650 129.050 ;
        RECT 117.910 128.960 118.050 139.610 ;
        RECT 118.370 136.530 118.510 141.650 ;
        RECT 118.310 136.210 118.570 136.530 ;
        RECT 118.310 133.490 118.570 133.810 ;
        RECT 118.370 131.770 118.510 133.490 ;
        RECT 118.830 132.450 118.970 148.790 ;
        RECT 118.770 132.130 119.030 132.450 ;
        RECT 118.310 131.450 118.570 131.770 ;
        RECT 119.690 131.450 119.950 131.770 ;
        RECT 119.230 129.750 119.490 130.070 ;
        RECT 117.390 128.820 118.050 128.960 ;
        RECT 117.390 128.730 117.650 128.820 ;
        RECT 116.990 128.140 117.590 128.280 ;
        RECT 117.450 123.950 117.590 128.140 ;
        RECT 117.390 123.630 117.650 123.950 ;
        RECT 116.930 114.790 117.190 115.110 ;
        RECT 116.990 113.410 117.130 114.790 ;
        RECT 116.930 113.265 117.190 113.410 ;
        RECT 116.920 112.895 117.200 113.265 ;
        RECT 117.450 112.640 117.590 123.630 ;
        RECT 117.910 123.610 118.050 128.820 ;
        RECT 119.290 127.010 119.430 129.750 ;
        RECT 119.750 129.390 119.890 131.450 ;
        RECT 119.690 129.070 119.950 129.390 ;
        RECT 119.230 126.690 119.490 127.010 ;
        RECT 117.850 123.290 118.110 123.610 ;
        RECT 117.910 113.750 118.050 123.290 ;
        RECT 118.310 121.250 118.570 121.570 ;
        RECT 118.370 118.510 118.510 121.250 ;
        RECT 118.770 118.870 119.030 119.190 ;
        RECT 118.310 118.190 118.570 118.510 ;
        RECT 118.310 114.450 118.570 114.770 ;
        RECT 117.850 113.430 118.110 113.750 ;
        RECT 116.990 112.500 117.590 112.640 ;
        RECT 116.070 110.450 116.670 110.590 ;
        RECT 115.090 110.030 115.350 110.350 ;
        RECT 114.170 109.690 114.430 110.010 ;
        RECT 115.150 109.750 115.290 110.030 ;
        RECT 114.230 107.630 114.370 109.690 ;
        RECT 115.150 109.610 116.210 109.750 ;
        RECT 116.530 109.670 116.670 110.450 ;
        RECT 114.630 109.010 114.890 109.330 ;
        RECT 114.170 107.310 114.430 107.630 ;
        RECT 114.230 103.890 114.370 107.310 ;
        RECT 114.690 104.230 114.830 109.010 ;
        RECT 115.090 107.310 115.350 107.630 ;
        RECT 114.630 103.910 114.890 104.230 ;
        RECT 114.170 103.570 114.430 103.890 ;
        RECT 115.150 103.745 115.290 107.310 ;
        RECT 115.550 106.290 115.810 106.610 ;
        RECT 115.610 104.230 115.750 106.290 ;
        RECT 115.550 103.910 115.810 104.230 ;
        RECT 115.080 103.375 115.360 103.745 ;
        RECT 114.170 102.550 114.430 102.870 ;
        RECT 114.230 102.190 114.370 102.550 ;
        RECT 114.170 101.870 114.430 102.190 ;
        RECT 115.090 101.870 115.350 102.190 ;
        RECT 115.150 100.150 115.290 101.870 ;
        RECT 115.090 99.830 115.350 100.150 ;
        RECT 115.610 98.790 115.750 103.910 ;
        RECT 116.070 99.130 116.210 109.610 ;
        RECT 116.470 109.350 116.730 109.670 ;
        RECT 116.530 107.630 116.670 109.350 ;
        RECT 116.470 107.310 116.730 107.630 ;
        RECT 116.470 106.630 116.730 106.950 ;
        RECT 116.530 105.590 116.670 106.630 ;
        RECT 116.470 105.270 116.730 105.590 ;
        RECT 116.470 101.870 116.730 102.190 ;
        RECT 116.530 100.150 116.670 101.870 ;
        RECT 116.470 99.830 116.730 100.150 ;
        RECT 116.010 98.810 116.270 99.130 ;
        RECT 115.550 98.470 115.810 98.790 ;
        RECT 115.610 97.430 115.750 98.470 ;
        RECT 116.530 98.450 116.670 99.830 ;
        RECT 116.990 99.810 117.130 112.500 ;
        RECT 118.370 109.670 118.510 114.450 ;
        RECT 118.830 112.390 118.970 118.870 ;
        RECT 118.770 112.070 119.030 112.390 ;
        RECT 118.310 109.350 118.570 109.670 ;
        RECT 118.310 105.270 118.570 105.590 ;
        RECT 118.370 103.890 118.510 105.270 ;
        RECT 118.770 104.250 119.030 104.570 ;
        RECT 118.310 103.570 118.570 103.890 ;
        RECT 118.310 102.550 118.570 102.870 ;
        RECT 116.930 99.490 117.190 99.810 ;
        RECT 116.470 98.130 116.730 98.450 ;
        RECT 115.550 97.110 115.810 97.430 ;
        RECT 115.090 96.770 115.350 97.090 ;
        RECT 114.630 96.430 114.890 96.750 ;
        RECT 113.710 95.410 113.970 95.730 ;
        RECT 113.710 92.690 113.970 93.010 ;
        RECT 113.250 91.670 113.510 91.990 ;
        RECT 112.790 91.330 113.050 91.650 ;
        RECT 112.330 90.990 112.590 91.310 ;
        RECT 112.850 90.290 112.990 91.330 ;
        RECT 113.770 91.310 113.910 92.690 ;
        RECT 114.690 91.310 114.830 96.430 ;
        RECT 115.150 92.185 115.290 96.770 ;
        RECT 115.610 93.690 115.750 97.110 ;
        RECT 116.530 96.750 116.670 98.130 ;
        RECT 118.370 97.430 118.510 102.550 ;
        RECT 118.830 102.530 118.970 104.250 ;
        RECT 118.770 102.210 119.030 102.530 ;
        RECT 118.310 97.110 118.570 97.430 ;
        RECT 118.370 96.750 118.510 97.110 ;
        RECT 116.470 96.430 116.730 96.750 ;
        RECT 118.310 96.430 118.570 96.750 ;
        RECT 118.830 94.030 118.970 102.210 ;
        RECT 119.290 96.410 119.430 126.690 ;
        RECT 119.750 124.630 119.890 129.070 ;
        RECT 120.210 125.990 120.350 159.250 ;
        RECT 120.610 156.270 120.870 156.590 ;
        RECT 121.070 156.270 121.330 156.590 ;
        RECT 120.670 137.065 120.810 156.270 ;
        RECT 121.130 155.910 121.270 156.270 ;
        RECT 121.070 155.590 121.330 155.910 ;
        RECT 121.130 154.210 121.270 155.590 ;
        RECT 121.070 153.890 121.330 154.210 ;
        RECT 121.530 153.550 121.790 153.870 ;
        RECT 121.070 153.210 121.330 153.530 ;
        RECT 121.130 150.470 121.270 153.210 ;
        RECT 121.070 150.150 121.330 150.470 ;
        RECT 121.590 145.905 121.730 153.550 ;
        RECT 122.050 149.110 122.190 177.690 ;
        RECT 122.510 169.510 122.650 178.710 ;
        RECT 123.430 178.350 123.570 178.710 ;
        RECT 123.370 178.030 123.630 178.350 ;
        RECT 124.290 178.030 124.550 178.350 ;
        RECT 125.670 178.030 125.930 178.350 ;
        RECT 123.430 177.330 123.570 178.030 ;
        RECT 123.370 177.010 123.630 177.330 ;
        RECT 122.450 169.190 122.710 169.510 ;
        RECT 122.510 156.840 122.650 169.190 ;
        RECT 122.910 161.370 123.170 161.690 ;
        RECT 122.970 158.970 123.110 161.370 ;
        RECT 122.910 158.650 123.170 158.970 ;
        RECT 122.910 156.840 123.170 156.930 ;
        RECT 122.510 156.700 123.170 156.840 ;
        RECT 122.910 156.610 123.170 156.700 ;
        RECT 123.430 155.910 123.570 177.010 ;
        RECT 124.350 175.970 124.490 178.030 ;
        RECT 124.290 175.650 124.550 175.970 ;
        RECT 125.730 174.610 125.870 178.030 ;
        RECT 125.670 174.290 125.930 174.610 ;
        RECT 126.650 172.910 126.790 180.750 ;
        RECT 134.010 180.730 134.150 182.450 ;
        RECT 134.930 181.945 135.070 185.170 ;
        RECT 134.860 181.575 135.140 181.945 ;
        RECT 133.950 180.410 134.210 180.730 ;
        RECT 131.190 180.070 131.450 180.390 ;
        RECT 131.250 179.030 131.390 180.070 ;
        RECT 135.850 179.030 135.990 185.850 ;
        RECT 136.770 185.345 136.910 187.890 ;
        RECT 136.700 184.975 136.980 185.345 ;
        RECT 137.630 185.170 137.890 185.490 ;
        RECT 136.710 179.730 136.970 180.050 ;
        RECT 131.190 178.710 131.450 179.030 ;
        RECT 135.790 178.710 136.050 179.030 ;
        RECT 136.770 178.350 136.910 179.730 ;
        RECT 137.690 178.545 137.830 185.170 ;
        RECT 136.710 178.030 136.970 178.350 ;
        RECT 137.620 178.175 137.900 178.545 ;
        RECT 127.510 174.970 127.770 175.290 ;
        RECT 127.050 174.290 127.310 174.610 ;
        RECT 126.590 172.590 126.850 172.910 ;
        RECT 125.670 169.870 125.930 170.190 ;
        RECT 123.830 169.530 124.090 169.850 ;
        RECT 123.890 168.150 124.030 169.530 ;
        RECT 123.830 167.830 124.090 168.150 ;
        RECT 125.730 165.430 125.870 169.870 ;
        RECT 126.130 169.530 126.390 169.850 ;
        RECT 125.670 165.110 125.930 165.430 ;
        RECT 124.290 161.710 124.550 162.030 ;
        RECT 124.350 161.010 124.490 161.710 ;
        RECT 124.290 160.690 124.550 161.010 ;
        RECT 125.670 160.690 125.930 161.010 ;
        RECT 125.730 156.590 125.870 160.690 ;
        RECT 123.830 156.270 124.090 156.590 ;
        RECT 125.670 156.270 125.930 156.590 ;
        RECT 123.370 155.590 123.630 155.910 ;
        RECT 121.990 148.790 122.250 149.110 ;
        RECT 123.890 147.410 124.030 156.270 ;
        RECT 126.190 153.530 126.330 169.530 ;
        RECT 126.650 167.470 126.790 172.590 ;
        RECT 126.590 167.150 126.850 167.470 ;
        RECT 126.650 164.410 126.790 167.150 ;
        RECT 126.590 164.090 126.850 164.410 ;
        RECT 126.650 162.030 126.790 164.090 ;
        RECT 126.590 161.710 126.850 162.030 ;
        RECT 127.110 158.710 127.250 174.290 ;
        RECT 127.570 173.590 127.710 174.970 ;
        RECT 128.420 174.775 128.700 175.145 ;
        RECT 134.410 174.970 134.670 175.290 ;
        RECT 128.490 174.610 128.630 174.775 ;
        RECT 128.430 174.290 128.690 174.610 ;
        RECT 129.810 174.290 130.070 174.610 ;
        RECT 130.270 174.290 130.530 174.610 ;
        RECT 127.510 173.270 127.770 173.590 ;
        RECT 129.870 173.250 130.010 174.290 ;
        RECT 129.810 172.930 130.070 173.250 ;
        RECT 130.330 170.870 130.470 174.290 ;
        RECT 134.470 173.590 134.610 174.970 ;
        RECT 134.410 173.270 134.670 173.590 ;
        RECT 136.710 173.270 136.970 173.590 ;
        RECT 132.110 172.930 132.370 173.250 ;
        RECT 130.270 170.550 130.530 170.870 ;
        RECT 128.890 169.190 129.150 169.510 ;
        RECT 127.970 163.410 128.230 163.730 ;
        RECT 128.030 162.030 128.170 163.410 ;
        RECT 127.970 161.710 128.230 162.030 ;
        RECT 127.110 158.570 127.710 158.710 ;
        RECT 126.590 157.970 126.850 158.290 ;
        RECT 127.050 157.970 127.310 158.290 ;
        RECT 126.650 157.270 126.790 157.970 ;
        RECT 127.110 157.270 127.250 157.970 ;
        RECT 126.590 156.950 126.850 157.270 ;
        RECT 127.050 156.950 127.310 157.270 ;
        RECT 127.050 156.270 127.310 156.590 ;
        RECT 126.590 154.230 126.850 154.550 ;
        RECT 126.130 153.210 126.390 153.530 ;
        RECT 124.290 152.870 124.550 153.190 ;
        RECT 124.750 152.870 125.010 153.190 ;
        RECT 124.350 151.830 124.490 152.870 ;
        RECT 124.290 151.510 124.550 151.830 ;
        RECT 124.810 148.090 124.950 152.870 ;
        RECT 126.650 151.490 126.790 154.230 ;
        RECT 126.590 151.170 126.850 151.490 ;
        RECT 124.750 147.770 125.010 148.090 ;
        RECT 123.830 147.090 124.090 147.410 ;
        RECT 124.810 146.390 124.950 147.770 ;
        RECT 124.750 146.070 125.010 146.390 ;
        RECT 121.520 145.535 121.800 145.905 ;
        RECT 126.590 145.730 126.850 146.050 ;
        RECT 122.450 144.370 122.710 144.690 ;
        RECT 122.510 142.310 122.650 144.370 ;
        RECT 123.830 143.010 124.090 143.330 ;
        RECT 123.890 142.310 124.030 143.010 ;
        RECT 124.750 142.330 125.010 142.650 ;
        RECT 122.450 141.990 122.710 142.310 ;
        RECT 123.830 141.990 124.090 142.310 ;
        RECT 121.530 141.650 121.790 141.970 ;
        RECT 121.590 140.610 121.730 141.650 ;
        RECT 121.530 140.290 121.790 140.610 ;
        RECT 123.890 138.190 124.030 141.990 ;
        RECT 123.890 138.050 124.490 138.190 ;
        RECT 120.600 136.695 120.880 137.065 ;
        RECT 121.070 136.890 121.330 137.210 ;
        RECT 121.130 130.070 121.270 136.890 ;
        RECT 122.450 136.550 122.710 136.870 ;
        RECT 122.510 132.790 122.650 136.550 ;
        RECT 123.830 136.210 124.090 136.530 ;
        RECT 123.890 133.810 124.030 136.210 ;
        RECT 123.830 133.490 124.090 133.810 ;
        RECT 122.450 132.470 122.710 132.790 ;
        RECT 122.510 131.430 122.650 132.470 ;
        RECT 123.890 132.110 124.030 133.490 ;
        RECT 123.830 131.790 124.090 132.110 ;
        RECT 122.450 131.110 122.710 131.430 ;
        RECT 121.070 129.750 121.330 130.070 ;
        RECT 120.150 125.670 120.410 125.990 ;
        RECT 119.690 124.310 119.950 124.630 ;
        RECT 119.750 120.890 119.890 124.310 ;
        RECT 121.990 121.250 122.250 121.570 ;
        RECT 119.690 120.570 119.950 120.890 ;
        RECT 119.690 118.190 119.950 118.510 ;
        RECT 119.750 114.770 119.890 118.190 ;
        RECT 122.050 118.170 122.190 121.250 ;
        RECT 122.510 120.550 122.650 131.110 ;
        RECT 124.350 129.730 124.490 138.050 ;
        RECT 124.810 137.210 124.950 142.330 ;
        RECT 126.130 142.220 126.390 142.310 ;
        RECT 126.650 142.220 126.790 145.730 ;
        RECT 126.130 142.080 126.790 142.220 ;
        RECT 126.130 141.990 126.390 142.080 ;
        RECT 125.210 140.290 125.470 140.610 ;
        RECT 125.270 137.890 125.410 140.290 ;
        RECT 125.670 139.950 125.930 140.270 ;
        RECT 126.130 139.950 126.390 140.270 ;
        RECT 125.730 138.230 125.870 139.950 ;
        RECT 125.670 137.910 125.930 138.230 ;
        RECT 125.210 137.570 125.470 137.890 ;
        RECT 124.750 136.890 125.010 137.210 ;
        RECT 124.810 132.110 124.950 136.890 ;
        RECT 126.190 135.170 126.330 139.950 ;
        RECT 126.650 139.930 126.790 142.080 ;
        RECT 126.590 139.610 126.850 139.930 ;
        RECT 127.110 137.550 127.250 156.270 ;
        RECT 127.570 142.650 127.710 158.570 ;
        RECT 127.970 147.090 128.230 147.410 ;
        RECT 128.030 145.710 128.170 147.090 ;
        RECT 127.970 145.390 128.230 145.710 ;
        RECT 128.430 145.390 128.690 145.710 ;
        RECT 128.490 143.330 128.630 145.390 ;
        RECT 128.430 143.010 128.690 143.330 ;
        RECT 127.510 142.330 127.770 142.650 ;
        RECT 127.970 142.330 128.230 142.650 ;
        RECT 127.510 141.650 127.770 141.970 ;
        RECT 127.570 140.270 127.710 141.650 ;
        RECT 128.030 140.270 128.170 142.330 ;
        RECT 128.430 141.990 128.690 142.310 ;
        RECT 128.490 140.950 128.630 141.990 ;
        RECT 128.430 140.630 128.690 140.950 ;
        RECT 127.510 139.950 127.770 140.270 ;
        RECT 127.970 139.950 128.230 140.270 ;
        RECT 128.490 138.190 128.630 140.630 ;
        RECT 127.570 138.050 128.630 138.190 ;
        RECT 127.050 137.230 127.310 137.550 ;
        RECT 126.130 134.850 126.390 135.170 ;
        RECT 127.050 134.170 127.310 134.490 ;
        RECT 126.130 133.830 126.390 134.150 ;
        RECT 125.670 132.130 125.930 132.450 ;
        RECT 124.750 131.790 125.010 132.110 ;
        RECT 124.290 129.410 124.550 129.730 ;
        RECT 124.350 124.710 124.490 129.410 ;
        RECT 124.810 129.390 124.950 131.790 ;
        RECT 125.730 129.390 125.870 132.130 ;
        RECT 126.190 132.110 126.330 133.830 ;
        RECT 126.130 131.790 126.390 132.110 ;
        RECT 126.190 130.070 126.330 131.790 ;
        RECT 126.130 129.750 126.390 130.070 ;
        RECT 124.750 129.070 125.010 129.390 ;
        RECT 125.670 129.070 125.930 129.390 ;
        RECT 125.210 125.330 125.470 125.650 ;
        RECT 124.350 124.570 124.950 124.710 ;
        RECT 124.290 123.630 124.550 123.950 ;
        RECT 124.350 121.910 124.490 123.630 ;
        RECT 124.290 121.590 124.550 121.910 ;
        RECT 124.810 121.230 124.950 124.570 ;
        RECT 124.750 120.910 125.010 121.230 ;
        RECT 122.450 120.230 122.710 120.550 ;
        RECT 121.990 117.850 122.250 118.170 ;
        RECT 119.690 114.450 119.950 114.770 ;
        RECT 120.150 112.410 120.410 112.730 ;
        RECT 121.070 112.410 121.330 112.730 ;
        RECT 120.210 110.350 120.350 112.410 ;
        RECT 120.150 110.030 120.410 110.350 ;
        RECT 121.130 107.290 121.270 112.410 ;
        RECT 122.510 110.010 122.650 120.230 ;
        RECT 124.810 119.190 124.950 120.910 ;
        RECT 125.270 120.890 125.410 125.330 ;
        RECT 126.190 124.710 126.330 129.750 ;
        RECT 126.590 129.070 126.850 129.390 ;
        RECT 126.650 128.710 126.790 129.070 ;
        RECT 127.110 128.710 127.250 134.170 ;
        RECT 127.570 131.770 127.710 138.050 ;
        RECT 128.430 134.510 128.690 134.830 ;
        RECT 128.490 131.770 128.630 134.510 ;
        RECT 127.510 131.450 127.770 131.770 ;
        RECT 128.430 131.450 128.690 131.770 ;
        RECT 128.950 129.390 129.090 169.190 ;
        RECT 129.350 168.850 129.610 169.170 ;
        RECT 129.810 168.850 130.070 169.170 ;
        RECT 130.730 168.850 130.990 169.170 ;
        RECT 129.410 164.750 129.550 168.850 ;
        RECT 129.870 167.810 130.010 168.850 ;
        RECT 129.810 167.490 130.070 167.810 ;
        RECT 129.350 164.430 129.610 164.750 ;
        RECT 130.270 163.410 130.530 163.730 ;
        RECT 130.330 155.910 130.470 163.410 ;
        RECT 130.270 155.590 130.530 155.910 ;
        RECT 130.790 155.570 130.930 168.850 ;
        RECT 131.650 161.370 131.910 161.690 ;
        RECT 131.710 155.910 131.850 161.370 ;
        RECT 131.650 155.590 131.910 155.910 ;
        RECT 130.730 155.250 130.990 155.570 ;
        RECT 129.350 152.530 129.610 152.850 ;
        RECT 129.410 151.830 129.550 152.530 ;
        RECT 129.350 151.510 129.610 151.830 ;
        RECT 132.170 150.130 132.310 172.930 ;
        RECT 135.330 172.590 135.590 172.910 ;
        RECT 134.410 171.570 134.670 171.890 ;
        RECT 133.490 169.530 133.750 169.850 ;
        RECT 133.550 168.150 133.690 169.530 ;
        RECT 133.490 167.830 133.750 168.150 ;
        RECT 134.470 167.470 134.610 171.570 ;
        RECT 134.860 171.375 135.140 171.745 ;
        RECT 134.930 168.150 135.070 171.375 ;
        RECT 135.390 169.850 135.530 172.590 ;
        RECT 135.330 169.530 135.590 169.850 ;
        RECT 136.770 168.345 136.910 173.270 ;
        RECT 134.870 167.830 135.130 168.150 ;
        RECT 136.700 167.975 136.980 168.345 ;
        RECT 134.410 167.150 134.670 167.470 ;
        RECT 135.790 167.150 136.050 167.470 ;
        RECT 133.490 164.090 133.750 164.410 ;
        RECT 133.550 162.710 133.690 164.090 ;
        RECT 135.850 162.710 135.990 167.150 ;
        RECT 136.710 166.130 136.970 166.450 ;
        RECT 136.770 164.945 136.910 166.130 ;
        RECT 136.700 164.575 136.980 164.945 ;
        RECT 133.490 162.390 133.750 162.710 ;
        RECT 135.790 162.390 136.050 162.710 ;
        RECT 136.700 161.175 136.980 161.545 ;
        RECT 136.710 161.030 136.970 161.175 ;
        RECT 135.330 157.970 135.590 158.290 ;
        RECT 135.390 156.590 135.530 157.970 ;
        RECT 138.080 157.775 138.360 158.145 ;
        RECT 135.330 156.270 135.590 156.590 ;
        RECT 136.250 156.270 136.510 156.590 ;
        RECT 132.570 153.550 132.830 153.870 ;
        RECT 132.630 151.150 132.770 153.550 ;
        RECT 133.950 153.210 134.210 153.530 ;
        RECT 134.010 151.830 134.150 153.210 ;
        RECT 134.870 152.530 135.130 152.850 ;
        RECT 133.950 151.510 134.210 151.830 ;
        RECT 134.930 151.345 135.070 152.530 ;
        RECT 132.570 150.830 132.830 151.150 ;
        RECT 134.860 150.975 135.140 151.345 ;
        RECT 132.110 149.810 132.370 150.130 ;
        RECT 129.810 147.770 130.070 148.090 ;
        RECT 129.350 147.430 129.610 147.750 ;
        RECT 129.410 146.390 129.550 147.430 ;
        RECT 129.350 146.070 129.610 146.390 ;
        RECT 129.870 145.905 130.010 147.770 ;
        RECT 136.310 147.410 136.450 156.270 ;
        RECT 136.710 155.250 136.970 155.570 ;
        RECT 136.770 154.745 136.910 155.250 ;
        RECT 136.700 154.375 136.980 154.745 ;
        RECT 138.150 154.550 138.290 157.775 ;
        RECT 138.090 154.230 138.350 154.550 ;
        RECT 136.700 147.575 136.980 147.945 ;
        RECT 136.250 147.090 136.510 147.410 ;
        RECT 134.870 146.070 135.130 146.390 ;
        RECT 129.800 145.535 130.080 145.905 ;
        RECT 130.270 145.730 130.530 146.050 ;
        RECT 129.870 142.650 130.010 145.535 ;
        RECT 129.810 142.330 130.070 142.650 ;
        RECT 129.810 137.570 130.070 137.890 ;
        RECT 129.350 137.230 129.610 137.550 ;
        RECT 128.890 129.070 129.150 129.390 ;
        RECT 126.590 128.390 126.850 128.710 ;
        RECT 127.050 128.390 127.310 128.710 ;
        RECT 125.730 124.570 126.330 124.710 ;
        RECT 125.210 120.570 125.470 120.890 ;
        RECT 122.910 118.870 123.170 119.190 ;
        RECT 124.750 118.870 125.010 119.190 ;
        RECT 122.450 109.690 122.710 110.010 ;
        RECT 122.970 109.670 123.110 118.870 ;
        RECT 123.370 118.190 123.630 118.510 ;
        RECT 124.750 118.420 125.010 118.510 ;
        RECT 125.730 118.420 125.870 124.570 ;
        RECT 126.130 123.860 126.390 123.950 ;
        RECT 126.650 123.860 126.790 128.390 ;
        RECT 127.110 123.950 127.250 128.390 ;
        RECT 127.970 126.010 128.230 126.330 ;
        RECT 127.510 125.670 127.770 125.990 ;
        RECT 126.130 123.720 126.790 123.860 ;
        RECT 126.130 123.630 126.390 123.720 ;
        RECT 127.050 123.630 127.310 123.950 ;
        RECT 127.110 118.510 127.250 123.630 ;
        RECT 124.750 118.280 125.870 118.420 ;
        RECT 124.750 118.190 125.010 118.280 ;
        RECT 123.430 115.450 123.570 118.190 ;
        RECT 125.270 117.830 125.410 118.280 ;
        RECT 126.590 118.190 126.850 118.510 ;
        RECT 127.050 118.190 127.310 118.510 ;
        RECT 126.650 117.910 126.790 118.190 ;
        RECT 127.570 117.910 127.710 125.670 ;
        RECT 128.030 124.390 128.170 126.010 ;
        RECT 128.030 124.250 129.090 124.390 ;
        RECT 125.210 117.510 125.470 117.830 ;
        RECT 126.650 117.770 128.630 117.910 ;
        RECT 125.270 115.450 125.410 117.510 ;
        RECT 127.510 115.470 127.770 115.790 ;
        RECT 123.370 115.130 123.630 115.450 ;
        RECT 125.210 115.130 125.470 115.450 ;
        RECT 126.590 115.130 126.850 115.450 ;
        RECT 122.910 109.350 123.170 109.670 ;
        RECT 123.430 108.390 123.570 115.130 ;
        RECT 124.290 113.090 124.550 113.410 ;
        RECT 124.350 112.585 124.490 113.090 ;
        RECT 125.270 113.070 125.410 115.130 ;
        RECT 125.210 112.750 125.470 113.070 ;
        RECT 126.650 112.640 126.790 115.130 ;
        RECT 127.050 114.450 127.310 114.770 ;
        RECT 127.110 113.410 127.250 114.450 ;
        RECT 127.050 113.090 127.310 113.410 ;
        RECT 127.570 113.070 127.710 115.470 ;
        RECT 127.970 114.790 128.230 115.110 ;
        RECT 128.030 113.070 128.170 114.790 ;
        RECT 127.510 112.750 127.770 113.070 ;
        RECT 127.970 112.750 128.230 113.070 ;
        RECT 124.280 112.215 124.560 112.585 ;
        RECT 126.650 112.500 127.250 112.640 ;
        RECT 122.970 108.250 123.570 108.390 ;
        RECT 122.970 107.630 123.110 108.250 ;
        RECT 124.350 107.630 124.490 112.215 ;
        RECT 125.210 112.070 125.470 112.390 ;
        RECT 125.270 110.350 125.410 112.070 ;
        RECT 125.210 110.030 125.470 110.350 ;
        RECT 122.910 107.310 123.170 107.630 ;
        RECT 123.370 107.310 123.630 107.630 ;
        RECT 123.830 107.310 124.090 107.630 ;
        RECT 124.290 107.310 124.550 107.630 ;
        RECT 126.590 107.540 126.850 107.630 ;
        RECT 127.110 107.540 127.250 112.500 ;
        RECT 126.590 107.400 127.250 107.540 ;
        RECT 126.590 107.310 126.850 107.400 ;
        RECT 120.610 106.970 120.870 107.290 ;
        RECT 121.070 106.970 121.330 107.290 ;
        RECT 120.670 105.785 120.810 106.970 ;
        RECT 120.600 105.415 120.880 105.785 ;
        RECT 121.130 104.570 121.270 106.970 ;
        RECT 121.070 104.250 121.330 104.570 ;
        RECT 122.970 102.190 123.110 107.310 ;
        RECT 123.430 105.590 123.570 107.310 ;
        RECT 123.370 105.270 123.630 105.590 ;
        RECT 122.910 101.870 123.170 102.190 ;
        RECT 122.970 99.130 123.110 101.870 ;
        RECT 123.890 101.850 124.030 107.310 ;
        RECT 126.590 104.930 126.850 105.250 ;
        RECT 124.290 103.630 124.550 103.890 ;
        RECT 124.290 103.570 124.950 103.630 ;
        RECT 125.210 103.570 125.470 103.890 ;
        RECT 126.130 103.570 126.390 103.890 ;
        RECT 124.350 103.490 124.950 103.570 ;
        RECT 124.290 102.210 124.550 102.530 ;
        RECT 123.830 101.530 124.090 101.850 ;
        RECT 123.830 100.850 124.090 101.170 ;
        RECT 123.890 99.470 124.030 100.850 ;
        RECT 124.350 99.470 124.490 102.210 ;
        RECT 123.830 99.150 124.090 99.470 ;
        RECT 124.290 99.150 124.550 99.470 ;
        RECT 122.910 98.810 123.170 99.130 ;
        RECT 123.370 98.360 123.630 98.450 ;
        RECT 122.970 98.220 123.630 98.360 ;
        RECT 122.970 97.430 123.110 98.220 ;
        RECT 123.370 98.130 123.630 98.220 ;
        RECT 120.610 97.110 120.870 97.430 ;
        RECT 122.910 97.110 123.170 97.430 ;
        RECT 123.370 97.110 123.630 97.430 ;
        RECT 119.230 96.090 119.490 96.410 ;
        RECT 120.150 95.410 120.410 95.730 ;
        RECT 118.770 93.710 119.030 94.030 ;
        RECT 115.550 93.370 115.810 93.690 ;
        RECT 115.080 91.815 115.360 92.185 ;
        RECT 113.250 90.990 113.510 91.310 ;
        RECT 113.710 90.990 113.970 91.310 ;
        RECT 114.630 90.990 114.890 91.310 ;
        RECT 113.310 90.825 113.450 90.990 ;
        RECT 113.240 90.455 113.520 90.825 ;
        RECT 112.790 89.970 113.050 90.290 ;
        RECT 113.250 89.970 113.510 90.290 ;
        RECT 111.930 89.750 112.530 89.890 ;
        RECT 112.390 88.590 112.530 89.750 ;
        RECT 112.330 88.270 112.590 88.590 ;
        RECT 113.310 88.250 113.450 89.970 ;
        RECT 110.030 87.930 110.290 88.250 ;
        RECT 111.410 87.930 111.670 88.250 ;
        RECT 113.250 87.930 113.510 88.250 ;
        RECT 108.190 87.590 108.450 87.910 ;
        RECT 113.770 87.570 113.910 90.990 ;
        RECT 115.610 90.290 115.750 93.370 ;
        RECT 116.930 93.030 117.190 93.350 ;
        RECT 116.990 91.990 117.130 93.030 ;
        RECT 118.830 91.990 118.970 93.710 ;
        RECT 120.210 93.690 120.350 95.410 ;
        RECT 120.150 93.370 120.410 93.690 ;
        RECT 116.930 91.670 117.190 91.990 ;
        RECT 118.770 91.670 119.030 91.990 ;
        RECT 120.150 91.670 120.410 91.990 ;
        RECT 118.300 91.135 118.580 91.505 ;
        RECT 120.210 91.310 120.350 91.670 ;
        RECT 118.310 90.990 118.570 91.135 ;
        RECT 119.230 90.990 119.490 91.310 ;
        RECT 120.150 90.990 120.410 91.310 ;
        RECT 115.550 89.970 115.810 90.290 ;
        RECT 114.170 88.950 114.430 89.270 ;
        RECT 104.970 87.250 105.230 87.570 ;
        RECT 107.730 87.250 107.990 87.570 ;
        RECT 110.950 87.250 111.210 87.570 ;
        RECT 113.710 87.250 113.970 87.570 ;
        RECT 105.030 81.870 105.170 87.250 ;
        RECT 104.570 81.730 105.170 81.870 ;
        RECT 104.570 80.020 104.710 81.730 ;
        RECT 107.790 80.020 107.930 87.250 ;
        RECT 111.010 80.020 111.150 87.250 ;
        RECT 114.230 80.020 114.370 88.950 ;
        RECT 119.290 88.930 119.430 90.990 ;
        RECT 120.670 90.970 120.810 97.110 ;
        RECT 122.970 96.750 123.110 97.110 ;
        RECT 121.990 96.430 122.250 96.750 ;
        RECT 122.910 96.430 123.170 96.750 ;
        RECT 122.050 93.010 122.190 96.430 ;
        RECT 123.430 96.150 123.570 97.110 ;
        RECT 122.970 96.010 123.570 96.150 ;
        RECT 122.450 95.410 122.710 95.730 ;
        RECT 121.990 92.690 122.250 93.010 ;
        RECT 122.510 91.650 122.650 95.410 ;
        RECT 122.970 93.010 123.110 96.010 ;
        RECT 123.370 95.410 123.630 95.730 ;
        RECT 123.430 94.710 123.570 95.410 ;
        RECT 123.370 94.390 123.630 94.710 ;
        RECT 122.910 92.690 123.170 93.010 ;
        RECT 122.450 91.330 122.710 91.650 ;
        RECT 120.610 90.650 120.870 90.970 ;
        RECT 119.230 88.610 119.490 88.930 ;
        RECT 122.970 88.250 123.110 92.690 ;
        RECT 123.430 91.650 123.570 94.390 ;
        RECT 123.370 91.330 123.630 91.650 ;
        RECT 123.890 88.250 124.030 99.150 ;
        RECT 124.290 98.470 124.550 98.790 ;
        RECT 124.350 96.750 124.490 98.470 ;
        RECT 124.290 96.430 124.550 96.750 ;
        RECT 124.350 93.260 124.490 96.430 ;
        RECT 124.810 94.370 124.950 103.490 ;
        RECT 125.270 102.190 125.410 103.570 ;
        RECT 125.210 101.870 125.470 102.190 ;
        RECT 126.190 101.510 126.330 103.570 ;
        RECT 126.130 101.190 126.390 101.510 ;
        RECT 126.650 99.130 126.790 104.930 ;
        RECT 127.110 102.190 127.250 107.400 ;
        RECT 127.970 106.290 128.230 106.610 ;
        RECT 127.510 105.270 127.770 105.590 ;
        RECT 127.570 104.230 127.710 105.270 ;
        RECT 128.030 104.230 128.170 106.290 ;
        RECT 127.510 103.910 127.770 104.230 ;
        RECT 127.970 103.910 128.230 104.230 ;
        RECT 127.050 101.870 127.310 102.190 ;
        RECT 127.050 101.190 127.310 101.510 ;
        RECT 127.110 99.130 127.250 101.190 ;
        RECT 128.490 99.130 128.630 117.770 ;
        RECT 128.950 111.030 129.090 124.250 ;
        RECT 129.410 113.750 129.550 137.230 ;
        RECT 129.870 125.990 130.010 137.570 ;
        RECT 130.330 137.550 130.470 145.730 ;
        RECT 133.950 145.390 134.210 145.710 ;
        RECT 133.030 139.950 133.290 140.270 ;
        RECT 133.090 138.230 133.230 139.950 ;
        RECT 133.490 138.930 133.750 139.250 ;
        RECT 133.550 138.230 133.690 138.930 ;
        RECT 131.650 137.910 131.910 138.230 ;
        RECT 133.030 137.910 133.290 138.230 ;
        RECT 133.490 137.910 133.750 138.230 ;
        RECT 130.270 137.230 130.530 137.550 ;
        RECT 131.190 136.890 131.450 137.210 ;
        RECT 131.710 137.120 131.850 137.910 ;
        RECT 134.010 137.745 134.150 145.390 ;
        RECT 134.930 144.545 135.070 146.070 ;
        RECT 136.310 146.050 136.450 147.090 ;
        RECT 136.770 146.390 136.910 147.575 ;
        RECT 136.710 146.070 136.970 146.390 ;
        RECT 136.250 145.730 136.510 146.050 ;
        RECT 134.860 144.175 135.140 144.545 ;
        RECT 135.790 141.650 136.050 141.970 ;
        RECT 135.850 140.270 135.990 141.650 ;
        RECT 135.790 139.950 136.050 140.270 ;
        RECT 134.870 138.930 135.130 139.250 ;
        RECT 133.940 137.375 134.220 137.745 ;
        RECT 132.110 137.120 132.370 137.210 ;
        RECT 131.710 136.980 132.370 137.120 ;
        RECT 130.730 134.850 130.990 135.170 ;
        RECT 130.790 131.430 130.930 134.850 ;
        RECT 130.730 131.110 130.990 131.430 ;
        RECT 131.250 130.070 131.390 136.890 ;
        RECT 131.190 129.750 131.450 130.070 ;
        RECT 131.710 126.670 131.850 136.980 ;
        RECT 132.110 136.890 132.370 136.980 ;
        RECT 134.930 136.870 135.070 138.930 ;
        RECT 136.310 137.210 136.450 145.730 ;
        RECT 136.700 140.775 136.980 141.145 ;
        RECT 136.710 140.630 136.970 140.775 ;
        RECT 136.700 137.375 136.980 137.745 ;
        RECT 136.250 136.890 136.510 137.210 ;
        RECT 134.870 136.550 135.130 136.870 ;
        RECT 135.790 136.210 136.050 136.530 ;
        RECT 135.850 134.830 135.990 136.210 ;
        RECT 136.770 135.510 136.910 137.375 ;
        RECT 136.710 135.190 136.970 135.510 ;
        RECT 135.790 134.510 136.050 134.830 ;
        RECT 135.790 133.830 136.050 134.150 ;
        RECT 136.700 133.975 136.980 134.345 ;
        RECT 134.410 133.490 134.670 133.810 ;
        RECT 134.470 131.770 134.610 133.490 ;
        RECT 134.410 131.450 134.670 131.770 ;
        RECT 132.110 131.110 132.370 131.430 ;
        RECT 132.170 128.370 132.310 131.110 ;
        RECT 132.110 128.050 132.370 128.370 ;
        RECT 131.650 126.350 131.910 126.670 ;
        RECT 132.170 126.330 132.310 128.050 ;
        RECT 135.850 126.330 135.990 133.830 ;
        RECT 136.770 132.790 136.910 133.975 ;
        RECT 136.710 132.470 136.970 132.790 ;
        RECT 136.700 130.575 136.980 130.945 ;
        RECT 136.770 130.070 136.910 130.575 ;
        RECT 136.710 129.750 136.970 130.070 ;
        RECT 136.700 127.175 136.980 127.545 ;
        RECT 136.710 127.030 136.970 127.175 ;
        RECT 132.110 126.010 132.370 126.330 ;
        RECT 133.490 126.070 133.750 126.330 ;
        RECT 133.490 126.010 134.150 126.070 ;
        RECT 135.790 126.010 136.050 126.330 ;
        RECT 129.810 125.670 130.070 125.990 ;
        RECT 133.550 125.930 134.150 126.010 ;
        RECT 129.870 121.570 130.010 125.670 ;
        RECT 134.010 122.930 134.150 125.930 ;
        RECT 134.870 125.330 135.130 125.650 ;
        RECT 134.930 124.145 135.070 125.330 ;
        RECT 134.860 123.775 135.140 124.145 ;
        RECT 133.950 122.610 134.210 122.930 ;
        RECT 129.810 121.250 130.070 121.570 ;
        RECT 134.010 121.230 134.150 122.610 ;
        RECT 133.950 120.910 134.210 121.230 ;
        RECT 133.030 120.230 133.290 120.550 ;
        RECT 130.270 119.890 130.530 120.210 ;
        RECT 130.330 115.450 130.470 119.890 ;
        RECT 132.110 117.510 132.370 117.830 ;
        RECT 130.270 115.130 130.530 115.450 ;
        RECT 129.350 113.430 129.610 113.750 ;
        RECT 131.190 112.750 131.450 113.070 ;
        RECT 128.890 110.710 129.150 111.030 ;
        RECT 130.730 110.710 130.990 111.030 ;
        RECT 130.790 110.010 130.930 110.710 ;
        RECT 131.250 110.690 131.390 112.750 ;
        RECT 131.190 110.370 131.450 110.690 ;
        RECT 131.250 110.010 131.390 110.370 ;
        RECT 130.730 109.690 130.990 110.010 ;
        RECT 131.190 109.690 131.450 110.010 ;
        RECT 129.810 109.010 130.070 109.330 ;
        RECT 129.870 108.310 130.010 109.010 ;
        RECT 129.810 107.990 130.070 108.310 ;
        RECT 130.790 107.540 130.930 109.690 ;
        RECT 131.650 109.350 131.910 109.670 ;
        RECT 131.190 107.540 131.450 107.630 ;
        RECT 130.790 107.400 131.450 107.540 ;
        RECT 130.790 104.570 130.930 107.400 ;
        RECT 131.190 107.310 131.450 107.400 ;
        RECT 131.710 107.290 131.850 109.350 ;
        RECT 131.650 106.970 131.910 107.290 ;
        RECT 131.710 105.785 131.850 106.970 ;
        RECT 131.640 105.415 131.920 105.785 ;
        RECT 130.730 104.250 130.990 104.570 ;
        RECT 131.710 104.230 131.850 105.415 ;
        RECT 132.170 104.570 132.310 117.510 ;
        RECT 133.090 113.750 133.230 120.230 ;
        RECT 133.030 113.430 133.290 113.750 ;
        RECT 132.570 109.690 132.830 110.010 ;
        RECT 132.630 106.950 132.770 109.690 ;
        RECT 132.570 106.630 132.830 106.950 ;
        RECT 133.490 106.290 133.750 106.610 ;
        RECT 133.550 105.105 133.690 106.290 ;
        RECT 133.480 104.735 133.760 105.105 ;
        RECT 132.110 104.250 132.370 104.570 ;
        RECT 131.650 103.910 131.910 104.230 ;
        RECT 126.590 98.810 126.850 99.130 ;
        RECT 127.050 98.810 127.310 99.130 ;
        RECT 128.430 98.810 128.690 99.130 ;
        RECT 132.110 98.470 132.370 98.790 ;
        RECT 131.650 98.360 131.910 98.450 ;
        RECT 131.250 98.220 131.910 98.360 ;
        RECT 125.670 96.770 125.930 97.090 ;
        RECT 125.200 95.895 125.480 96.265 ;
        RECT 124.750 94.050 125.010 94.370 ;
        RECT 125.270 94.030 125.410 95.895 ;
        RECT 125.730 94.710 125.870 96.770 ;
        RECT 125.670 94.390 125.930 94.710 ;
        RECT 125.210 93.710 125.470 94.030 ;
        RECT 127.040 93.855 127.320 94.225 ;
        RECT 127.110 93.350 127.250 93.855 ;
        RECT 131.250 93.690 131.390 98.220 ;
        RECT 131.650 98.130 131.910 98.220 ;
        RECT 132.170 96.750 132.310 98.470 ;
        RECT 131.650 96.430 131.910 96.750 ;
        RECT 132.110 96.430 132.370 96.750 ;
        RECT 131.710 94.710 131.850 96.430 ;
        RECT 131.650 94.390 131.910 94.710 ;
        RECT 128.430 93.370 128.690 93.690 ;
        RECT 130.270 93.370 130.530 93.690 ;
        RECT 131.190 93.370 131.450 93.690 ;
        RECT 125.210 93.260 125.470 93.350 ;
        RECT 124.350 93.120 125.470 93.260 ;
        RECT 124.350 91.990 124.490 93.120 ;
        RECT 125.210 93.030 125.470 93.120 ;
        RECT 127.050 93.030 127.310 93.350 ;
        RECT 127.110 91.990 127.250 93.030 ;
        RECT 124.290 91.670 124.550 91.990 ;
        RECT 127.050 91.670 127.310 91.990 ;
        RECT 127.110 88.250 127.250 91.670 ;
        RECT 128.490 91.650 128.630 93.370 ;
        RECT 130.330 91.990 130.470 93.370 ;
        RECT 130.270 91.670 130.530 91.990 ;
        RECT 128.430 91.330 128.690 91.650 ;
        RECT 134.010 91.310 134.150 120.910 ;
        RECT 135.790 120.570 136.050 120.890 ;
        RECT 134.410 120.230 134.670 120.550 ;
        RECT 134.470 118.510 134.610 120.230 ;
        RECT 135.850 118.510 135.990 120.570 ;
        RECT 136.700 120.375 136.980 120.745 ;
        RECT 136.770 120.210 136.910 120.375 ;
        RECT 136.710 119.890 136.970 120.210 ;
        RECT 134.410 118.190 134.670 118.510 ;
        RECT 135.790 118.190 136.050 118.510 ;
        RECT 138.540 116.975 138.820 117.345 ;
        RECT 136.250 114.450 136.510 114.770 ;
        RECT 135.790 113.430 136.050 113.750 ;
        RECT 134.860 110.175 135.140 110.545 ;
        RECT 134.930 109.330 135.070 110.175 ;
        RECT 135.850 110.010 135.990 113.430 ;
        RECT 136.310 113.070 136.450 114.450 ;
        RECT 136.700 113.575 136.980 113.945 ;
        RECT 138.610 113.750 138.750 116.975 ;
        RECT 136.250 112.750 136.510 113.070 ;
        RECT 135.790 109.690 136.050 110.010 ;
        RECT 134.870 109.010 135.130 109.330 ;
        RECT 135.850 107.970 135.990 109.690 ;
        RECT 136.770 109.330 136.910 113.575 ;
        RECT 138.550 113.430 138.810 113.750 ;
        RECT 136.710 109.010 136.970 109.330 ;
        RECT 135.790 107.650 136.050 107.970 ;
        RECT 134.410 106.630 134.670 106.950 ;
        RECT 136.700 106.775 136.980 107.145 ;
        RECT 134.470 105.590 134.610 106.630 ;
        RECT 135.790 106.290 136.050 106.610 ;
        RECT 134.410 105.270 134.670 105.590 ;
        RECT 134.470 102.870 134.610 105.270 ;
        RECT 135.850 104.570 135.990 106.290 ;
        RECT 136.770 105.590 136.910 106.775 ;
        RECT 136.710 105.270 136.970 105.590 ;
        RECT 135.790 104.250 136.050 104.570 ;
        RECT 135.330 103.910 135.590 104.230 ;
        RECT 134.410 102.550 134.670 102.870 ;
        RECT 135.390 100.150 135.530 103.910 ;
        RECT 136.700 103.375 136.980 103.745 ;
        RECT 136.770 102.870 136.910 103.375 ;
        RECT 136.710 102.550 136.970 102.870 ;
        RECT 135.330 99.830 135.590 100.150 ;
        RECT 136.700 99.975 136.980 100.345 ;
        RECT 134.860 96.575 135.140 96.945 ;
        RECT 135.390 96.750 135.530 99.830 ;
        RECT 134.930 96.070 135.070 96.575 ;
        RECT 135.330 96.430 135.590 96.750 ;
        RECT 136.770 96.070 136.910 99.975 ;
        RECT 134.870 95.750 135.130 96.070 ;
        RECT 136.710 95.750 136.970 96.070 ;
        RECT 136.700 93.175 136.980 93.545 ;
        RECT 136.770 93.010 136.910 93.175 ;
        RECT 136.710 92.690 136.970 93.010 ;
        RECT 132.110 90.990 132.370 91.310 ;
        RECT 133.950 90.990 134.210 91.310 ;
        RECT 132.170 88.250 132.310 90.990 ;
        RECT 136.710 90.145 136.970 90.290 ;
        RECT 136.700 89.775 136.980 90.145 ;
        RECT 117.390 87.930 117.650 88.250 ;
        RECT 122.910 87.930 123.170 88.250 ;
        RECT 123.830 87.930 124.090 88.250 ;
        RECT 127.050 87.930 127.310 88.250 ;
        RECT 132.110 87.930 132.370 88.250 ;
        RECT 117.450 80.020 117.590 87.930 ;
        RECT 120.610 87.250 120.870 87.570 ;
        RECT 123.830 87.250 124.090 87.570 ;
        RECT 127.050 87.250 127.310 87.570 ;
        RECT 130.270 87.250 130.530 87.570 ;
        RECT 120.670 80.020 120.810 87.250 ;
        RECT 123.890 80.020 124.030 87.250 ;
        RECT 127.110 80.020 127.250 87.250 ;
        RECT 130.330 80.020 130.470 87.250 ;
        RECT 59.420 76.020 59.700 80.020 ;
        RECT 65.860 76.020 66.140 80.020 ;
        RECT 69.080 76.020 69.360 80.020 ;
        RECT 72.300 76.020 72.580 80.020 ;
        RECT 75.520 76.020 75.800 80.020 ;
        RECT 78.740 76.020 79.020 80.020 ;
        RECT 81.960 76.020 82.240 80.020 ;
        RECT 85.180 76.020 85.460 80.020 ;
        RECT 88.400 76.020 88.680 80.020 ;
        RECT 91.620 76.020 91.900 80.020 ;
        RECT 94.840 76.020 95.120 80.020 ;
        RECT 98.060 76.020 98.340 80.020 ;
        RECT 101.280 76.020 101.560 80.020 ;
        RECT 104.500 76.020 104.780 80.020 ;
        RECT 107.720 76.020 108.000 80.020 ;
        RECT 110.940 76.020 111.220 80.020 ;
        RECT 114.160 76.020 114.440 80.020 ;
        RECT 117.380 76.020 117.660 80.020 ;
        RECT 120.600 76.020 120.880 80.020 ;
        RECT 123.820 76.020 124.100 80.020 ;
        RECT 127.040 76.020 127.320 80.020 ;
        RECT 130.260 76.020 130.540 80.020 ;
        RECT 26.810 59.165 27.090 63.165 ;
        RECT 30.030 59.165 30.310 63.165 ;
        RECT 33.250 59.165 33.530 63.165 ;
        RECT 36.470 59.165 36.750 63.165 ;
        RECT 39.690 59.165 39.970 63.165 ;
        RECT 26.880 51.290 27.020 59.165 ;
        RECT 30.100 52.730 30.240 59.165 ;
        RECT 30.100 52.590 31.160 52.730 ;
        RECT 28.470 51.455 30.010 51.825 ;
        RECT 26.820 50.970 27.080 51.290 ;
        RECT 18.540 49.950 18.800 50.270 ;
        RECT 23.140 49.950 23.400 50.270 ;
        RECT 23.600 49.950 23.860 50.270 ;
        RECT 18.600 48.570 18.740 49.950 ;
        RECT 23.200 48.570 23.340 49.950 ;
        RECT 18.540 48.250 18.800 48.570 ;
        RECT 23.140 48.250 23.400 48.570 ;
        RECT 23.660 48.085 23.800 49.950 ;
        RECT 25.440 49.270 25.700 49.590 ;
        RECT 30.500 49.270 30.760 49.590 ;
        RECT 25.500 48.230 25.640 49.270 ;
        RECT 23.590 47.715 23.870 48.085 ;
        RECT 25.440 47.910 25.700 48.230 ;
        RECT 26.360 47.570 26.620 47.890 ;
        RECT 27.730 47.715 28.010 48.085 ;
        RECT 24.060 46.550 24.320 46.870 ;
        RECT 24.120 44.830 24.260 46.550 ;
        RECT 24.970 46.355 25.250 46.725 ;
        RECT 24.060 44.510 24.320 44.830 ;
        RECT 16.240 44.170 16.500 44.490 ;
        RECT 13.930 42.955 14.210 43.325 ;
        RECT 16.300 43.130 16.440 44.170 ;
        RECT 21.300 43.830 21.560 44.150 ;
        RECT 21.760 43.830 22.020 44.150 ;
        RECT 13.940 42.810 14.200 42.955 ;
        RECT 16.240 42.810 16.500 43.130 ;
        RECT 21.360 42.450 21.500 43.830 ;
        RECT 21.820 43.130 21.960 43.830 ;
        RECT 24.120 43.130 24.260 44.510 ;
        RECT 21.760 42.810 22.020 43.130 ;
        RECT 24.060 42.810 24.320 43.130 ;
        RECT 21.300 42.130 21.560 42.450 ;
        RECT 19.920 41.790 20.180 42.110 ;
        RECT 16.700 41.450 16.960 41.770 ;
        RECT 16.760 39.730 16.900 41.450 ;
        RECT 16.700 39.410 16.960 39.730 ;
        RECT 19.980 39.050 20.120 41.790 ;
        RECT 24.120 39.390 24.260 42.810 ;
        RECT 21.300 39.070 21.560 39.390 ;
        RECT 24.060 39.070 24.320 39.390 ;
        RECT 19.920 38.730 20.180 39.050 ;
        RECT 14.400 38.390 14.660 38.710 ;
        RECT 19.000 38.390 19.260 38.710 ;
        RECT 14.460 37.350 14.600 38.390 ;
        RECT 14.400 37.030 14.660 37.350 ;
        RECT 13.930 36.155 14.210 36.525 ;
        RECT 14.000 32.250 14.140 36.155 ;
        RECT 14.400 35.670 14.660 35.990 ;
        RECT 14.460 34.290 14.600 35.670 ;
        RECT 19.060 34.970 19.200 38.390 ;
        RECT 19.000 34.650 19.260 34.970 ;
        RECT 14.400 33.970 14.660 34.290 ;
        RECT 13.940 31.930 14.200 32.250 ;
        RECT 14.460 31.570 14.600 33.970 ;
        RECT 19.460 32.950 19.720 33.270 ;
        RECT 19.520 32.250 19.660 32.950 ;
        RECT 19.460 31.930 19.720 32.250 ;
        RECT 14.400 31.250 14.660 31.570 ;
        RECT 19.980 31.230 20.120 38.730 ;
        RECT 21.360 37.010 21.500 39.070 ;
        RECT 25.040 37.350 25.180 46.355 ;
        RECT 26.420 45.850 26.560 47.570 ;
        RECT 26.360 45.530 26.620 45.850 ;
        RECT 26.360 42.810 26.620 43.130 ;
        RECT 27.280 42.810 27.540 43.130 ;
        RECT 26.420 39.730 26.560 42.810 ;
        RECT 27.340 40.410 27.480 42.810 ;
        RECT 27.280 40.090 27.540 40.410 ;
        RECT 26.360 39.410 26.620 39.730 ;
        RECT 24.980 37.030 25.240 37.350 ;
        RECT 21.300 36.690 21.560 37.010 ;
        RECT 27.340 34.970 27.480 40.090 ;
        RECT 27.800 34.970 27.940 47.715 ;
        RECT 28.470 46.015 30.010 46.385 ;
        RECT 30.560 44.830 30.700 49.270 ;
        RECT 31.020 47.210 31.160 52.590 ;
        RECT 33.320 51.290 33.460 59.165 ;
        RECT 33.260 50.970 33.520 51.290 ;
        RECT 31.420 50.630 31.680 50.950 ;
        RECT 30.960 46.890 31.220 47.210 ;
        RECT 31.480 45.850 31.620 50.630 ;
        RECT 36.540 50.270 36.680 59.165 ;
        RECT 39.760 51.290 39.900 59.165 ;
        RECT 47.050 56.555 47.330 56.925 ;
        RECT 44.290 53.155 44.570 53.525 ;
        RECT 39.700 50.970 39.960 51.290 ;
        RECT 38.320 50.630 38.580 50.950 ;
        RECT 33.720 49.950 33.980 50.270 ;
        RECT 36.480 49.950 36.740 50.270 ;
        RECT 31.770 48.735 33.310 49.105 ;
        RECT 33.780 48.570 33.920 49.950 ;
        RECT 34.180 49.270 34.440 49.590 ;
        RECT 33.720 48.250 33.980 48.570 ;
        RECT 34.240 48.230 34.380 49.270 ;
        RECT 34.180 47.910 34.440 48.230 ;
        RECT 38.380 47.890 38.520 50.630 ;
        RECT 44.360 50.270 44.500 53.155 ;
        RECT 47.120 50.270 47.260 56.555 ;
        RECT 41.540 49.950 41.800 50.270 ;
        RECT 44.300 49.950 44.560 50.270 ;
        RECT 45.680 50.125 45.940 50.270 ;
        RECT 40.160 49.270 40.420 49.590 ;
        RECT 35.100 47.570 35.360 47.890 ;
        RECT 36.480 47.570 36.740 47.890 ;
        RECT 38.320 47.570 38.580 47.890 ;
        RECT 31.880 47.230 32.140 47.550 ;
        RECT 31.420 45.530 31.680 45.850 ;
        RECT 31.940 44.830 32.080 47.230 ;
        RECT 34.640 46.550 34.900 46.870 ;
        RECT 34.700 45.170 34.840 46.550 ;
        RECT 34.640 44.850 34.900 45.170 ;
        RECT 35.160 44.830 35.300 47.570 ;
        RECT 36.020 47.230 36.280 47.550 ;
        RECT 30.500 44.510 30.760 44.830 ;
        RECT 30.960 44.510 31.220 44.830 ;
        RECT 31.880 44.510 32.140 44.830 ;
        RECT 33.720 44.510 33.980 44.830 ;
        RECT 34.180 44.510 34.440 44.830 ;
        RECT 35.100 44.510 35.360 44.830 ;
        RECT 30.500 43.830 30.760 44.150 ;
        RECT 28.470 40.575 30.010 40.945 ;
        RECT 28.470 35.135 30.010 35.505 ;
        RECT 27.280 34.650 27.540 34.970 ;
        RECT 27.740 34.650 28.000 34.970 ;
        RECT 22.220 33.630 22.480 33.950 ;
        RECT 19.460 30.910 19.720 31.230 ;
        RECT 19.920 30.910 20.180 31.230 ;
        RECT 14.400 30.570 14.660 30.890 ;
        RECT 13.930 29.355 14.210 29.725 ;
        RECT 14.000 25.450 14.140 29.355 ;
        RECT 14.460 28.850 14.600 30.570 ;
        RECT 16.700 30.230 16.960 30.550 ;
        RECT 14.400 28.530 14.660 28.850 ;
        RECT 16.760 28.170 16.900 30.230 ;
        RECT 16.700 27.850 16.960 28.170 ;
        RECT 14.400 25.470 14.660 25.790 ;
        RECT 13.940 25.130 14.200 25.450 ;
        RECT 14.460 24.090 14.600 25.470 ;
        RECT 19.520 25.450 19.660 30.910 ;
        RECT 22.280 29.530 22.420 33.630 ;
        RECT 27.340 31.910 27.480 34.650 ;
        RECT 30.560 33.950 30.700 43.830 ;
        RECT 31.020 43.130 31.160 44.510 ;
        RECT 31.770 43.295 33.310 43.665 ;
        RECT 30.960 42.810 31.220 43.130 ;
        RECT 30.960 42.130 31.220 42.450 ;
        RECT 31.020 35.990 31.160 42.130 ;
        RECT 31.420 41.110 31.680 41.430 ;
        RECT 31.480 37.090 31.620 41.110 ;
        RECT 33.780 40.410 33.920 44.510 ;
        RECT 33.720 40.090 33.980 40.410 ;
        RECT 34.240 39.810 34.380 44.510 ;
        RECT 36.080 42.790 36.220 47.230 ;
        RECT 36.540 45.850 36.680 47.570 ;
        RECT 37.400 46.550 37.660 46.870 ;
        RECT 36.480 45.530 36.740 45.850 ;
        RECT 36.540 45.250 36.680 45.530 ;
        RECT 36.540 45.110 37.140 45.250 ;
        RECT 36.480 44.170 36.740 44.490 ;
        RECT 36.020 42.470 36.280 42.790 ;
        RECT 34.640 41.790 34.900 42.110 ;
        RECT 33.780 39.670 34.380 39.810 ;
        RECT 33.780 38.710 33.920 39.670 ;
        RECT 34.700 39.390 34.840 41.790 ;
        RECT 35.100 39.750 35.360 40.070 ;
        RECT 34.640 39.070 34.900 39.390 ;
        RECT 34.180 38.730 34.440 39.050 ;
        RECT 33.720 38.390 33.980 38.710 ;
        RECT 31.770 37.855 33.310 38.225 ;
        RECT 31.480 36.950 32.080 37.090 ;
        RECT 31.420 36.350 31.680 36.670 ;
        RECT 30.960 35.670 31.220 35.990 ;
        RECT 27.740 33.630 28.000 33.950 ;
        RECT 30.500 33.630 30.760 33.950 ;
        RECT 27.800 32.250 27.940 33.630 ;
        RECT 27.740 31.930 28.000 32.250 ;
        RECT 25.900 31.590 26.160 31.910 ;
        RECT 27.280 31.590 27.540 31.910 ;
        RECT 22.220 29.210 22.480 29.530 ;
        RECT 21.300 28.190 21.560 28.510 ;
        RECT 19.460 25.130 19.720 25.450 ;
        RECT 19.000 24.790 19.260 25.110 ;
        RECT 14.400 23.770 14.660 24.090 ;
        RECT 14.460 20.690 14.600 23.770 ;
        RECT 17.160 22.410 17.420 22.730 ;
        RECT 17.220 21.370 17.360 22.410 ;
        RECT 19.060 21.370 19.200 24.790 ;
        RECT 19.520 21.370 19.660 25.130 ;
        RECT 21.360 23.410 21.500 28.190 ;
        RECT 22.280 26.130 22.420 29.210 ;
        RECT 22.220 25.810 22.480 26.130 ;
        RECT 25.960 25.790 26.100 31.590 ;
        RECT 27.280 30.570 27.540 30.890 ;
        RECT 27.340 28.170 27.480 30.570 ;
        RECT 28.470 29.695 30.010 30.065 ;
        RECT 27.280 27.850 27.540 28.170 ;
        RECT 21.760 25.470 22.020 25.790 ;
        RECT 25.900 25.470 26.160 25.790 ;
        RECT 21.300 23.090 21.560 23.410 ;
        RECT 21.820 21.370 21.960 25.470 ;
        RECT 17.160 21.050 17.420 21.370 ;
        RECT 19.000 21.050 19.260 21.370 ;
        RECT 19.460 21.050 19.720 21.370 ;
        RECT 21.760 21.050 22.020 21.370 ;
        RECT 24.060 21.050 24.320 21.370 ;
        RECT 14.400 20.370 14.660 20.690 ;
        RECT 11.630 19.835 11.910 20.205 ;
        RECT 11.640 19.690 11.900 19.835 ;
        RECT 24.120 17.630 24.260 21.050 ;
        RECT 25.960 20.350 26.100 25.470 ;
        RECT 30.500 24.790 30.760 25.110 ;
        RECT 28.470 24.255 30.010 24.625 ;
        RECT 30.560 21.370 30.700 24.790 ;
        RECT 31.020 23.070 31.160 35.670 ;
        RECT 31.480 33.950 31.620 36.350 ;
        RECT 31.940 34.630 32.080 36.950 ;
        RECT 31.880 34.310 32.140 34.630 ;
        RECT 31.420 33.630 31.680 33.950 ;
        RECT 31.770 32.415 33.310 32.785 ;
        RECT 33.780 31.230 33.920 38.390 ;
        RECT 34.240 37.690 34.380 38.730 ;
        RECT 34.180 37.370 34.440 37.690 ;
        RECT 35.160 34.290 35.300 39.750 ;
        RECT 35.560 38.730 35.820 39.050 ;
        RECT 35.100 33.970 35.360 34.290 ;
        RECT 34.640 32.160 34.900 32.250 ;
        RECT 35.160 32.160 35.300 33.970 ;
        RECT 34.640 32.020 35.300 32.160 ;
        RECT 34.640 31.930 34.900 32.020 ;
        RECT 33.720 30.910 33.980 31.230 ;
        RECT 34.180 30.910 34.440 31.230 ;
        RECT 34.240 27.830 34.380 30.910 ;
        RECT 35.160 28.930 35.300 32.020 ;
        RECT 35.620 29.190 35.760 38.730 ;
        RECT 36.080 35.990 36.220 42.470 ;
        RECT 36.540 41.770 36.680 44.170 ;
        RECT 36.480 41.450 36.740 41.770 ;
        RECT 36.540 37.690 36.680 41.450 ;
        RECT 36.480 37.370 36.740 37.690 ;
        RECT 36.020 35.670 36.280 35.990 ;
        RECT 36.080 34.630 36.220 35.670 ;
        RECT 36.020 34.310 36.280 34.630 ;
        RECT 36.020 30.570 36.280 30.890 ;
        RECT 34.700 28.850 35.300 28.930 ;
        RECT 35.560 28.870 35.820 29.190 ;
        RECT 34.640 28.790 35.300 28.850 ;
        RECT 34.640 28.530 34.900 28.790 ;
        RECT 31.420 27.510 31.680 27.830 ;
        RECT 34.180 27.510 34.440 27.830 ;
        RECT 31.480 26.130 31.620 27.510 ;
        RECT 31.770 26.975 33.310 27.345 ;
        RECT 31.420 25.810 31.680 26.130 ;
        RECT 31.480 24.090 31.620 25.810 ;
        RECT 31.420 23.770 31.680 24.090 ;
        RECT 30.960 22.750 31.220 23.070 ;
        RECT 30.500 21.050 30.760 21.370 ;
        RECT 31.480 21.030 31.620 23.770 ;
        RECT 31.770 21.535 33.310 21.905 ;
        RECT 31.420 20.770 31.680 21.030 ;
        RECT 30.560 20.710 31.680 20.770 ;
        RECT 30.560 20.630 31.620 20.710 ;
        RECT 25.900 20.030 26.160 20.350 ;
        RECT 28.470 18.815 30.010 19.185 ;
        RECT 24.060 17.310 24.320 17.630 ;
        RECT 29.120 17.540 29.380 17.630 ;
        RECT 30.560 17.540 30.700 20.630 ;
        RECT 31.420 19.350 31.680 19.670 ;
        RECT 29.120 17.400 30.700 17.540 ;
        RECT 29.120 17.310 29.380 17.400 ;
        RECT 31.480 17.290 31.620 19.350 ;
        RECT 34.240 18.650 34.380 27.510 ;
        RECT 36.080 26.470 36.220 30.570 ;
        RECT 37.000 29.530 37.140 45.110 ;
        RECT 37.460 44.830 37.600 46.550 ;
        RECT 37.400 44.510 37.660 44.830 ;
        RECT 40.220 42.450 40.360 49.270 ;
        RECT 41.070 47.800 41.350 48.085 ;
        RECT 40.680 47.715 41.350 47.800 ;
        RECT 40.680 47.660 41.340 47.715 ;
        RECT 40.680 42.790 40.820 47.660 ;
        RECT 41.080 47.570 41.340 47.660 ;
        RECT 41.600 47.210 41.740 49.950 ;
        RECT 45.670 49.755 45.950 50.125 ;
        RECT 47.060 49.950 47.320 50.270 ;
        RECT 43.840 49.270 44.100 49.590 ;
        RECT 46.600 49.270 46.860 49.590 ;
        RECT 41.540 46.890 41.800 47.210 ;
        RECT 41.600 45.850 41.740 46.890 ;
        RECT 43.380 46.550 43.640 46.870 ;
        RECT 41.540 45.530 41.800 45.850 ;
        RECT 43.440 44.830 43.580 46.550 ;
        RECT 43.380 44.510 43.640 44.830 ;
        RECT 43.900 43.130 44.040 49.270 ;
        RECT 44.300 47.570 44.560 47.890 ;
        RECT 44.360 45.850 44.500 47.570 ;
        RECT 44.760 46.890 45.020 47.210 ;
        RECT 44.300 45.530 44.560 45.850 ;
        RECT 44.820 45.250 44.960 46.890 ;
        RECT 44.360 45.110 44.960 45.250 ;
        RECT 43.840 42.810 44.100 43.130 ;
        RECT 40.620 42.470 40.880 42.790 ;
        RECT 41.080 42.470 41.340 42.790 ;
        RECT 40.160 42.130 40.420 42.450 ;
        RECT 38.320 41.110 38.580 41.430 ;
        RECT 38.380 34.970 38.520 41.110 ;
        RECT 39.240 38.390 39.500 38.710 ;
        RECT 39.300 37.010 39.440 38.390 ;
        RECT 40.220 37.010 40.360 42.130 ;
        RECT 41.140 41.770 41.280 42.470 ;
        RECT 43.900 42.450 44.040 42.810 ;
        RECT 43.840 42.130 44.100 42.450 ;
        RECT 41.080 41.450 41.340 41.770 ;
        RECT 41.140 39.390 41.280 41.450 ;
        RECT 42.000 39.750 42.260 40.070 ;
        RECT 41.080 39.070 41.340 39.390 ;
        RECT 39.240 36.690 39.500 37.010 ;
        RECT 40.160 36.690 40.420 37.010 ;
        RECT 38.320 34.650 38.580 34.970 ;
        RECT 37.860 32.950 38.120 33.270 ;
        RECT 36.940 29.210 37.200 29.530 ;
        RECT 36.020 26.150 36.280 26.470 ;
        RECT 36.080 21.370 36.220 26.150 ;
        RECT 37.000 26.130 37.140 29.210 ;
        RECT 36.940 25.810 37.200 26.130 ;
        RECT 36.020 21.050 36.280 21.370 ;
        RECT 37.000 20.350 37.140 25.810 ;
        RECT 37.920 25.790 38.060 32.950 ;
        RECT 38.380 31.570 38.520 34.650 ;
        RECT 42.060 34.370 42.200 39.750 ;
        RECT 42.920 39.410 43.180 39.730 ;
        RECT 42.460 35.670 42.720 35.990 ;
        RECT 41.140 34.230 42.200 34.370 ;
        RECT 41.140 33.950 41.280 34.230 ;
        RECT 41.080 33.630 41.340 33.950 ;
        RECT 42.000 33.630 42.260 33.950 ;
        RECT 40.620 32.950 40.880 33.270 ;
        RECT 42.060 33.125 42.200 33.630 ;
        RECT 42.520 33.610 42.660 35.670 ;
        RECT 42.460 33.290 42.720 33.610 ;
        RECT 40.680 31.570 40.820 32.950 ;
        RECT 41.990 32.755 42.270 33.125 ;
        RECT 42.520 31.910 42.660 33.290 ;
        RECT 42.460 31.590 42.720 31.910 ;
        RECT 38.320 31.250 38.580 31.570 ;
        RECT 40.620 31.250 40.880 31.570 ;
        RECT 39.690 29.355 39.970 29.725 ;
        RECT 37.860 25.470 38.120 25.790 ;
        RECT 37.920 25.110 38.060 25.470 ;
        RECT 37.860 24.790 38.120 25.110 ;
        RECT 39.760 23.070 39.900 29.355 ;
        RECT 42.520 28.850 42.660 31.590 ;
        RECT 42.980 29.530 43.120 39.410 ;
        RECT 43.900 39.390 44.040 42.130 ;
        RECT 44.360 39.390 44.500 45.110 ;
        RECT 44.760 44.510 45.020 44.830 ;
        RECT 44.820 39.925 44.960 44.510 ;
        RECT 45.680 43.830 45.940 44.150 ;
        RECT 46.140 43.830 46.400 44.150 ;
        RECT 45.220 42.130 45.480 42.450 ;
        RECT 45.280 40.410 45.420 42.130 ;
        RECT 45.220 40.090 45.480 40.410 ;
        RECT 44.750 39.555 45.030 39.925 ;
        RECT 45.740 39.810 45.880 43.830 ;
        RECT 46.200 43.130 46.340 43.830 ;
        RECT 46.140 42.810 46.400 43.130 ;
        RECT 46.660 42.450 46.800 49.270 ;
        RECT 47.060 47.570 47.320 47.890 ;
        RECT 47.120 46.725 47.260 47.570 ;
        RECT 47.050 46.355 47.330 46.725 ;
        RECT 47.060 44.510 47.320 44.830 ;
        RECT 47.120 43.325 47.260 44.510 ;
        RECT 47.050 42.955 47.330 43.325 ;
        RECT 46.600 42.130 46.860 42.450 ;
        RECT 46.660 40.070 46.800 42.130 ;
        RECT 45.740 39.670 46.340 39.810 ;
        RECT 46.600 39.750 46.860 40.070 ;
        RECT 46.200 39.390 46.340 39.670 ;
        RECT 43.840 39.070 44.100 39.390 ;
        RECT 44.300 39.070 44.560 39.390 ;
        RECT 45.680 39.070 45.940 39.390 ;
        RECT 46.140 39.070 46.400 39.390 ;
        RECT 44.360 34.630 44.500 39.070 ;
        RECT 44.760 36.690 45.020 37.010 ;
        RECT 44.300 34.310 44.560 34.630 ;
        RECT 44.820 33.950 44.960 36.690 ;
        RECT 45.740 34.970 45.880 39.070 ;
        RECT 46.200 37.010 46.340 39.070 ;
        RECT 46.140 36.690 46.400 37.010 ;
        RECT 47.060 36.690 47.320 37.010 ;
        RECT 47.120 36.525 47.260 36.690 ;
        RECT 47.050 36.155 47.330 36.525 ;
        RECT 45.680 34.650 45.940 34.970 ;
        RECT 44.300 33.630 44.560 33.950 ;
        RECT 44.760 33.630 45.020 33.950 ;
        RECT 44.360 32.250 44.500 33.630 ;
        RECT 45.220 33.290 45.480 33.610 ;
        RECT 44.300 31.930 44.560 32.250 ;
        RECT 43.840 31.250 44.100 31.570 ;
        RECT 44.300 31.250 44.560 31.570 ;
        RECT 42.920 29.210 43.180 29.530 ;
        RECT 42.460 28.530 42.720 28.850 ;
        RECT 40.160 28.190 40.420 28.510 ;
        RECT 42.920 28.190 43.180 28.510 ;
        RECT 40.220 25.110 40.360 28.190 ;
        RECT 41.080 27.510 41.340 27.830 ;
        RECT 41.140 26.810 41.280 27.510 ;
        RECT 41.080 26.490 41.340 26.810 ;
        RECT 42.980 25.790 43.120 28.190 ;
        RECT 43.370 25.955 43.650 26.325 ;
        RECT 43.380 25.810 43.640 25.955 ;
        RECT 42.920 25.470 43.180 25.790 ;
        RECT 40.160 24.790 40.420 25.110 ;
        RECT 38.320 22.750 38.580 23.070 ;
        RECT 39.700 22.750 39.960 23.070 ;
        RECT 36.940 20.030 37.200 20.350 ;
        RECT 37.400 20.030 37.660 20.350 ;
        RECT 34.180 18.330 34.440 18.650 ;
        RECT 37.460 18.310 37.600 20.030 ;
        RECT 38.380 19.525 38.520 22.750 ;
        RECT 38.310 19.155 38.590 19.525 ;
        RECT 37.400 17.990 37.660 18.310 ;
        RECT 37.460 17.630 37.600 17.990 ;
        RECT 40.220 17.630 40.360 24.790 ;
        RECT 42.980 24.090 43.120 25.470 ;
        RECT 43.900 25.110 44.040 31.250 ;
        RECT 43.840 24.790 44.100 25.110 ;
        RECT 42.920 23.770 43.180 24.090 ;
        RECT 43.380 23.430 43.640 23.750 ;
        RECT 41.080 22.925 41.340 23.070 ;
        RECT 41.070 22.555 41.350 22.925 ;
        RECT 42.460 22.070 42.720 22.390 ;
        RECT 42.920 22.070 43.180 22.390 ;
        RECT 42.520 20.350 42.660 22.070 ;
        RECT 42.980 20.690 43.120 22.070 ;
        RECT 42.920 20.370 43.180 20.690 ;
        RECT 42.460 20.030 42.720 20.350 ;
        RECT 42.520 17.970 42.660 20.030 ;
        RECT 43.440 18.310 43.580 23.430 ;
        RECT 43.900 23.070 44.040 24.790 ;
        RECT 44.360 24.090 44.500 31.250 ;
        RECT 44.760 30.910 45.020 31.230 ;
        RECT 44.820 26.810 44.960 30.910 ;
        RECT 45.280 28.510 45.420 33.290 ;
        RECT 46.140 31.250 46.400 31.570 ;
        RECT 45.220 28.190 45.480 28.510 ;
        RECT 45.680 28.190 45.940 28.510 ;
        RECT 44.760 26.490 45.020 26.810 ;
        RECT 45.280 26.470 45.420 28.190 ;
        RECT 45.220 26.150 45.480 26.470 ;
        RECT 44.760 25.810 45.020 26.130 ;
        RECT 44.300 23.770 44.560 24.090 ;
        RECT 44.820 23.070 44.960 25.810 ;
        RECT 43.840 22.750 44.100 23.070 ;
        RECT 44.760 22.750 45.020 23.070 ;
        RECT 43.900 18.650 44.040 22.750 ;
        RECT 45.740 21.370 45.880 28.190 ;
        RECT 46.200 25.790 46.340 31.250 ;
        RECT 46.140 25.470 46.400 25.790 ;
        RECT 47.060 25.130 47.320 25.450 ;
        RECT 46.600 23.090 46.860 23.410 ;
        RECT 46.140 22.750 46.400 23.070 ;
        RECT 45.680 21.050 45.940 21.370 ;
        RECT 46.200 18.650 46.340 22.750 ;
        RECT 43.840 18.330 44.100 18.650 ;
        RECT 46.140 18.330 46.400 18.650 ;
        RECT 43.380 17.990 43.640 18.310 ;
        RECT 42.460 17.650 42.720 17.970 ;
        RECT 37.400 17.310 37.660 17.630 ;
        RECT 40.160 17.310 40.420 17.630 ;
        RECT 42.920 17.310 43.180 17.630 ;
        RECT 31.420 16.970 31.680 17.290 ;
        RECT 26.820 16.630 27.080 16.950 ;
        RECT 29.580 16.630 29.840 16.950 ;
        RECT 33.720 16.630 33.980 16.950 ;
        RECT 39.700 16.630 39.960 16.950 ;
        RECT 26.880 9.400 27.020 16.630 ;
        RECT 29.640 11.250 29.780 16.630 ;
        RECT 31.770 16.095 33.310 16.465 ;
        RECT 33.780 11.250 33.920 16.630 ;
        RECT 29.640 11.110 30.240 11.250 ;
        RECT 30.100 9.400 30.240 11.110 ;
        RECT 33.320 11.110 33.920 11.250 ;
        RECT 33.320 9.400 33.460 11.110 ;
        RECT 39.760 9.400 39.900 16.630 ;
        RECT 42.980 16.125 43.120 17.310 ;
        RECT 42.910 15.755 43.190 16.125 ;
        RECT 46.660 12.725 46.800 23.090 ;
        RECT 47.120 23.070 47.260 25.130 ;
        RECT 47.060 22.750 47.320 23.070 ;
        RECT 47.120 20.350 47.260 22.750 ;
        RECT 47.060 20.030 47.320 20.350 ;
        RECT 46.590 12.355 46.870 12.725 ;
        RECT 26.810 5.400 27.090 9.400 ;
        RECT 30.030 5.400 30.310 9.400 ;
        RECT 33.250 5.400 33.530 9.400 ;
        RECT 39.690 5.400 39.970 9.400 ;
      LAYER met3 ;
        RECT 143.900 225.090 144.220 225.470 ;
        RECT 143.910 224.380 144.210 225.090 ;
        RECT 32.160 211.855 33.740 212.185 ;
        RECT 28.860 209.135 30.440 209.465 ;
        RECT 32.160 206.415 33.740 206.745 ;
        RECT 7.810 205.710 11.810 205.860 ;
        RECT 7.810 205.410 13.020 205.710 ;
        RECT 7.810 205.260 11.810 205.410 ;
        RECT 8.335 204.350 8.665 204.365 ;
        RECT 12.720 204.350 13.020 205.410 ;
        RECT 8.335 204.050 13.020 204.350 ;
        RECT 8.335 204.035 8.665 204.050 ;
        RECT 28.860 203.695 30.440 204.025 ;
        RECT 32.160 200.975 33.740 201.305 ;
        RECT 28.860 198.255 30.440 198.585 ;
        RECT 32.160 195.535 33.740 195.865 ;
        RECT 75.495 193.480 75.825 193.485 ;
        RECT 75.240 193.470 75.825 193.480 ;
        RECT 75.040 193.170 75.825 193.470 ;
        RECT 75.240 193.160 75.825 193.170 ;
        RECT 75.495 193.155 75.825 193.160 ;
        RECT 28.860 192.815 30.440 193.145 ;
        RECT 63.535 191.430 63.865 191.445 ;
        RECT 71.355 191.430 71.685 191.445 ;
        RECT 79.175 191.430 79.505 191.445 ;
        RECT 63.535 191.130 79.505 191.430 ;
        RECT 63.535 191.115 63.865 191.130 ;
        RECT 71.355 191.115 71.685 191.130 ;
        RECT 79.175 191.115 79.505 191.130 ;
        RECT 113.675 191.440 114.005 191.445 ;
        RECT 113.675 191.430 114.260 191.440 ;
        RECT 113.675 191.130 114.460 191.430 ;
        RECT 113.675 191.120 114.260 191.130 ;
        RECT 113.675 191.115 114.005 191.120 ;
        RECT 110.915 190.750 111.245 190.765 ;
        RECT 116.435 190.750 116.765 190.765 ;
        RECT 110.915 190.450 116.765 190.750 ;
        RECT 110.915 190.435 111.245 190.450 ;
        RECT 116.435 190.435 116.765 190.450 ;
        RECT 32.160 190.095 33.740 190.425 ;
        RECT 137.135 188.710 137.465 188.725 ;
        RECT 140.470 188.710 144.470 188.860 ;
        RECT 137.135 188.410 144.470 188.710 ;
        RECT 137.135 188.395 137.465 188.410 ;
        RECT 140.470 188.260 144.470 188.410 ;
        RECT 28.860 187.375 30.440 187.705 ;
        RECT 30.415 186.670 30.745 186.685 ;
        RECT 33.175 186.670 33.505 186.685 ;
        RECT 30.415 186.370 33.505 186.670 ;
        RECT 30.415 186.355 30.745 186.370 ;
        RECT 33.175 186.355 33.505 186.370 ;
        RECT 136.675 185.310 137.005 185.325 ;
        RECT 140.470 185.310 144.470 185.460 ;
        RECT 136.675 185.010 144.470 185.310 ;
        RECT 136.675 184.995 137.005 185.010 ;
        RECT 32.160 184.655 33.740 184.985 ;
        RECT 140.470 184.860 144.470 185.010 ;
        RECT 106.775 184.630 107.105 184.645 ;
        RECT 112.755 184.630 113.085 184.645 ;
        RECT 106.775 184.330 113.085 184.630 ;
        RECT 106.775 184.315 107.105 184.330 ;
        RECT 112.755 184.315 113.085 184.330 ;
        RECT 110.915 183.270 111.245 183.285 ;
        RECT 119.655 183.270 119.985 183.285 ;
        RECT 110.915 182.970 119.985 183.270 ;
        RECT 110.915 182.955 111.245 182.970 ;
        RECT 119.655 182.955 119.985 182.970 ;
        RECT 12.015 182.590 12.345 182.605 ;
        RECT 11.800 182.275 12.345 182.590 ;
        RECT 11.800 182.060 12.100 182.275 ;
        RECT 7.810 181.610 12.100 182.060 ;
        RECT 28.860 181.935 30.440 182.265 ;
        RECT 134.835 181.910 135.165 181.925 ;
        RECT 140.470 181.910 144.470 182.060 ;
        RECT 134.835 181.610 144.470 181.910 ;
        RECT 7.810 181.460 11.810 181.610 ;
        RECT 134.835 181.595 135.165 181.610 ;
        RECT 140.470 181.460 144.470 181.610 ;
        RECT 71.355 181.230 71.685 181.245 ;
        RECT 73.195 181.230 73.525 181.245 ;
        RECT 76.415 181.230 76.745 181.245 ;
        RECT 71.355 180.930 76.745 181.230 ;
        RECT 71.355 180.915 71.685 180.930 ;
        RECT 73.195 180.915 73.525 180.930 ;
        RECT 76.415 180.915 76.745 180.930 ;
        RECT 109.535 180.550 109.865 180.565 ;
        RECT 116.435 180.550 116.765 180.565 ;
        RECT 109.535 180.250 116.765 180.550 ;
        RECT 109.535 180.235 109.865 180.250 ;
        RECT 116.435 180.235 116.765 180.250 ;
        RECT 114.595 179.870 114.925 179.885 ;
        RECT 117.815 179.880 118.145 179.885 ;
        RECT 117.560 179.870 118.145 179.880 ;
        RECT 114.595 179.570 116.980 179.870 ;
        RECT 117.360 179.570 118.145 179.870 ;
        RECT 114.595 179.555 114.925 179.570 ;
        RECT 32.160 179.215 33.740 179.545 ;
        RECT 116.680 179.205 116.980 179.570 ;
        RECT 117.560 179.560 118.145 179.570 ;
        RECT 117.815 179.555 118.145 179.560 ;
        RECT 71.815 179.190 72.145 179.205 ;
        RECT 77.795 179.190 78.125 179.205 ;
        RECT 71.815 178.890 78.125 179.190 ;
        RECT 71.815 178.875 72.145 178.890 ;
        RECT 77.795 178.875 78.125 178.890 ;
        RECT 107.235 179.190 107.565 179.205 ;
        RECT 113.880 179.190 114.260 179.200 ;
        RECT 114.595 179.190 114.925 179.205 ;
        RECT 116.680 179.190 117.225 179.205 ;
        RECT 117.815 179.190 118.145 179.205 ;
        RECT 107.235 178.890 114.925 179.190 ;
        RECT 116.440 178.890 118.145 179.190 ;
        RECT 107.235 178.875 107.565 178.890 ;
        RECT 113.880 178.880 114.260 178.890 ;
        RECT 114.595 178.875 114.925 178.890 ;
        RECT 116.895 178.875 117.225 178.890 ;
        RECT 117.815 178.875 118.145 178.890 ;
        RECT 65.375 178.510 65.705 178.525 ;
        RECT 75.035 178.510 75.365 178.525 ;
        RECT 65.375 178.210 75.365 178.510 ;
        RECT 65.375 178.195 65.705 178.210 ;
        RECT 75.035 178.195 75.365 178.210 ;
        RECT 137.595 178.510 137.925 178.525 ;
        RECT 140.470 178.510 144.470 178.660 ;
        RECT 137.595 178.210 144.470 178.510 ;
        RECT 137.595 178.195 137.925 178.210 ;
        RECT 140.470 178.060 144.470 178.210 ;
        RECT 28.860 176.495 30.440 176.825 ;
        RECT 128.395 175.110 128.725 175.125 ;
        RECT 140.470 175.110 144.470 175.260 ;
        RECT 128.395 174.810 144.470 175.110 ;
        RECT 128.395 174.795 128.725 174.810 ;
        RECT 140.470 174.660 144.470 174.810 ;
        RECT 32.160 173.775 33.740 174.105 ;
        RECT 31.080 172.390 31.460 172.400 ;
        RECT 31.795 172.390 32.125 172.405 ;
        RECT 31.080 172.090 32.125 172.390 ;
        RECT 31.080 172.080 31.460 172.090 ;
        RECT 31.795 172.075 32.125 172.090 ;
        RECT 134.835 171.710 135.165 171.725 ;
        RECT 140.470 171.710 144.470 171.860 ;
        RECT 134.835 171.410 144.470 171.710 ;
        RECT 134.835 171.395 135.165 171.410 ;
        RECT 28.860 171.055 30.440 171.385 ;
        RECT 140.470 171.260 144.470 171.410 ;
        RECT 112.755 170.350 113.085 170.365 ;
        RECT 119.195 170.350 119.525 170.365 ;
        RECT 112.755 170.050 119.525 170.350 ;
        RECT 112.755 170.035 113.085 170.050 ;
        RECT 119.195 170.035 119.525 170.050 ;
        RECT 115.055 169.670 115.385 169.685 ;
        RECT 116.435 169.670 116.765 169.685 ;
        RECT 117.815 169.670 118.145 169.685 ;
        RECT 115.055 169.370 118.145 169.670 ;
        RECT 115.055 169.355 115.385 169.370 ;
        RECT 116.435 169.355 116.765 169.370 ;
        RECT 117.815 169.355 118.145 169.370 ;
        RECT 12.015 168.990 12.345 169.005 ;
        RECT 11.800 168.675 12.345 168.990 ;
        RECT 113.675 168.990 114.005 169.005 ;
        RECT 117.355 168.990 117.685 169.005 ;
        RECT 113.675 168.690 117.685 168.990 ;
        RECT 113.675 168.675 114.005 168.690 ;
        RECT 117.355 168.675 117.685 168.690 ;
        RECT 11.800 168.460 12.100 168.675 ;
        RECT 7.810 168.010 12.100 168.460 ;
        RECT 32.160 168.335 33.740 168.665 ;
        RECT 48.815 168.310 49.145 168.325 ;
        RECT 52.035 168.310 52.365 168.325 ;
        RECT 75.495 168.320 75.825 168.325 ;
        RECT 48.815 168.010 52.365 168.310 ;
        RECT 7.810 167.860 11.810 168.010 ;
        RECT 48.815 167.995 49.145 168.010 ;
        RECT 52.035 167.995 52.365 168.010 ;
        RECT 75.240 168.310 75.825 168.320 ;
        RECT 136.675 168.310 137.005 168.325 ;
        RECT 140.470 168.310 144.470 168.460 ;
        RECT 75.240 168.010 76.050 168.310 ;
        RECT 136.675 168.010 144.470 168.310 ;
        RECT 75.240 168.000 75.825 168.010 ;
        RECT 75.495 167.995 75.825 168.000 ;
        RECT 136.675 167.995 137.005 168.010 ;
        RECT 140.470 167.860 144.470 168.010 ;
        RECT 107.235 167.630 107.565 167.645 ;
        RECT 111.375 167.630 111.705 167.645 ;
        RECT 107.235 167.330 111.705 167.630 ;
        RECT 107.235 167.315 107.565 167.330 ;
        RECT 111.375 167.315 111.705 167.330 ;
        RECT 28.860 165.615 30.440 165.945 ;
        RECT 136.675 164.910 137.005 164.925 ;
        RECT 140.470 164.910 144.470 165.060 ;
        RECT 136.675 164.610 144.470 164.910 ;
        RECT 136.675 164.595 137.005 164.610 ;
        RECT 140.470 164.460 144.470 164.610 ;
        RECT 32.160 162.895 33.740 163.225 ;
        RECT 136.675 161.510 137.005 161.525 ;
        RECT 140.470 161.510 144.470 161.660 ;
        RECT 136.675 161.210 144.470 161.510 ;
        RECT 136.675 161.195 137.005 161.210 ;
        RECT 140.470 161.060 144.470 161.210 ;
        RECT 28.860 160.175 30.440 160.505 ;
        RECT 138.055 158.110 138.385 158.125 ;
        RECT 140.470 158.110 144.470 158.260 ;
        RECT 138.055 157.810 144.470 158.110 ;
        RECT 138.055 157.795 138.385 157.810 ;
        RECT 32.160 157.455 33.740 157.785 ;
        RECT 140.470 157.660 144.470 157.810 ;
        RECT 12.015 155.390 12.345 155.405 ;
        RECT 11.800 155.075 12.345 155.390 ;
        RECT 11.800 154.860 12.100 155.075 ;
        RECT 7.810 154.410 12.100 154.860 ;
        RECT 28.860 154.735 30.440 155.065 ;
        RECT 136.675 154.710 137.005 154.725 ;
        RECT 140.470 154.710 144.470 154.860 ;
        RECT 136.675 154.410 144.470 154.710 ;
        RECT 7.810 154.260 11.810 154.410 ;
        RECT 136.675 154.395 137.005 154.410 ;
        RECT 140.470 154.260 144.470 154.410 ;
        RECT 117.355 154.040 117.685 154.045 ;
        RECT 117.355 154.030 117.940 154.040 ;
        RECT 117.130 153.730 117.940 154.030 ;
        RECT 117.355 153.720 117.940 153.730 ;
        RECT 117.355 153.715 117.685 153.720 ;
        RECT 32.160 152.015 33.740 152.345 ;
        RECT 7.810 151.310 11.810 151.460 ;
        RECT 15.235 151.310 15.565 151.325 ;
        RECT 7.810 151.010 15.565 151.310 ;
        RECT 7.810 150.860 11.810 151.010 ;
        RECT 15.235 150.995 15.565 151.010 ;
        RECT 134.835 151.310 135.165 151.325 ;
        RECT 140.470 151.310 144.470 151.460 ;
        RECT 134.835 151.010 144.470 151.310 ;
        RECT 134.835 150.995 135.165 151.010 ;
        RECT 140.470 150.860 144.470 151.010 ;
        RECT 28.860 149.295 30.440 149.625 ;
        RECT 28.115 147.910 28.445 147.925 ;
        RECT 37.315 147.910 37.645 147.925 ;
        RECT 28.115 147.610 37.645 147.910 ;
        RECT 28.115 147.595 28.445 147.610 ;
        RECT 37.315 147.595 37.645 147.610 ;
        RECT 136.675 147.910 137.005 147.925 ;
        RECT 140.470 147.910 144.470 148.060 ;
        RECT 136.675 147.610 144.470 147.910 ;
        RECT 136.675 147.595 137.005 147.610 ;
        RECT 140.470 147.460 144.470 147.610 ;
        RECT 32.160 146.575 33.740 146.905 ;
        RECT 83.315 145.870 83.645 145.885 ;
        RECT 86.075 145.870 86.405 145.885 ;
        RECT 83.315 145.570 86.405 145.870 ;
        RECT 83.315 145.555 83.645 145.570 ;
        RECT 86.075 145.555 86.405 145.570 ;
        RECT 115.975 145.870 116.305 145.885 ;
        RECT 121.495 145.870 121.825 145.885 ;
        RECT 129.775 145.870 130.105 145.885 ;
        RECT 115.975 145.570 130.105 145.870 ;
        RECT 115.975 145.555 116.305 145.570 ;
        RECT 121.495 145.555 121.825 145.570 ;
        RECT 129.775 145.555 130.105 145.570 ;
        RECT 134.835 144.510 135.165 144.525 ;
        RECT 140.470 144.510 144.470 144.660 ;
        RECT 134.835 144.210 144.470 144.510 ;
        RECT 134.835 144.195 135.165 144.210 ;
        RECT 28.860 143.855 30.440 144.185 ;
        RECT 140.470 144.060 144.470 144.210 ;
        RECT 32.160 141.135 33.740 141.465 ;
        RECT 136.675 141.110 137.005 141.125 ;
        RECT 140.470 141.110 144.470 141.260 ;
        RECT 136.675 140.810 144.470 141.110 ;
        RECT 136.675 140.795 137.005 140.810 ;
        RECT 140.470 140.660 144.470 140.810 ;
        RECT 28.860 138.415 30.440 138.745 ;
        RECT 114.595 137.710 114.925 137.725 ;
        RECT 133.915 137.710 134.245 137.725 ;
        RECT 114.595 137.410 134.245 137.710 ;
        RECT 114.595 137.395 114.925 137.410 ;
        RECT 133.915 137.395 134.245 137.410 ;
        RECT 136.675 137.710 137.005 137.725 ;
        RECT 140.470 137.710 144.470 137.860 ;
        RECT 136.675 137.410 144.470 137.710 ;
        RECT 136.675 137.395 137.005 137.410 ;
        RECT 140.470 137.260 144.470 137.410 ;
        RECT 115.975 137.030 116.305 137.045 ;
        RECT 120.575 137.030 120.905 137.045 ;
        RECT 115.975 136.730 120.905 137.030 ;
        RECT 115.975 136.715 116.305 136.730 ;
        RECT 120.575 136.715 120.905 136.730 ;
        RECT 32.160 135.695 33.740 136.025 ;
        RECT 31.080 134.990 31.460 135.000 ;
        RECT 31.795 134.990 32.125 135.005 ;
        RECT 33.635 134.990 33.965 135.005 ;
        RECT 31.080 134.690 33.965 134.990 ;
        RECT 31.080 134.680 31.460 134.690 ;
        RECT 31.795 134.675 32.125 134.690 ;
        RECT 33.635 134.675 33.965 134.690 ;
        RECT 136.675 134.310 137.005 134.325 ;
        RECT 140.470 134.310 144.470 134.460 ;
        RECT 136.675 134.010 144.470 134.310 ;
        RECT 136.675 133.995 137.005 134.010 ;
        RECT 140.470 133.860 144.470 134.010 ;
        RECT 28.860 132.975 30.440 133.305 ;
        RECT 44.675 131.590 45.005 131.605 ;
        RECT 48.815 131.590 49.145 131.605 ;
        RECT 44.675 131.290 49.145 131.590 ;
        RECT 44.675 131.275 45.005 131.290 ;
        RECT 48.815 131.275 49.145 131.290 ;
        RECT 136.675 130.910 137.005 130.925 ;
        RECT 140.470 130.910 144.470 131.060 ;
        RECT 136.675 130.610 144.470 130.910 ;
        RECT 136.675 130.595 137.005 130.610 ;
        RECT 32.160 130.255 33.740 130.585 ;
        RECT 140.470 130.460 144.470 130.610 ;
        RECT 28.860 127.535 30.440 127.865 ;
        RECT 136.675 127.510 137.005 127.525 ;
        RECT 140.470 127.510 144.470 127.660 ;
        RECT 136.675 127.210 144.470 127.510 ;
        RECT 136.675 127.195 137.005 127.210 ;
        RECT 140.470 127.060 144.470 127.210 ;
        RECT 32.160 124.815 33.740 125.145 ;
        RECT 134.835 124.110 135.165 124.125 ;
        RECT 140.470 124.110 144.470 124.260 ;
        RECT 134.835 123.810 144.470 124.110 ;
        RECT 134.835 123.795 135.165 123.810 ;
        RECT 140.470 123.660 144.470 123.810 ;
        RECT 28.860 122.095 30.440 122.425 ;
        RECT 30.415 120.710 30.745 120.725 ;
        RECT 35.935 120.710 36.265 120.725 ;
        RECT 38.695 120.710 39.025 120.725 ;
        RECT 30.415 120.410 39.025 120.710 ;
        RECT 30.415 120.395 30.745 120.410 ;
        RECT 35.935 120.395 36.265 120.410 ;
        RECT 38.695 120.395 39.025 120.410 ;
        RECT 136.675 120.710 137.005 120.725 ;
        RECT 140.470 120.710 144.470 120.860 ;
        RECT 136.675 120.410 144.470 120.710 ;
        RECT 136.675 120.395 137.005 120.410 ;
        RECT 140.470 120.260 144.470 120.410 ;
        RECT 32.160 119.375 33.740 119.705 ;
        RECT 62.615 117.310 62.945 117.325 ;
        RECT 68.595 117.310 68.925 117.325 ;
        RECT 62.615 117.010 68.925 117.310 ;
        RECT 62.615 116.995 62.945 117.010 ;
        RECT 68.595 116.995 68.925 117.010 ;
        RECT 138.515 117.310 138.845 117.325 ;
        RECT 140.470 117.310 144.470 117.460 ;
        RECT 138.515 117.010 144.470 117.310 ;
        RECT 138.515 116.995 138.845 117.010 ;
        RECT 28.860 116.655 30.440 116.985 ;
        RECT 140.470 116.860 144.470 117.010 ;
        RECT 32.160 113.935 33.740 114.265 ;
        RECT 136.675 113.910 137.005 113.925 ;
        RECT 140.470 113.910 144.470 114.060 ;
        RECT 136.675 113.610 144.470 113.910 ;
        RECT 136.675 113.595 137.005 113.610 ;
        RECT 140.470 113.460 144.470 113.610 ;
        RECT 91.135 113.230 91.465 113.245 ;
        RECT 116.895 113.230 117.225 113.245 ;
        RECT 91.135 112.930 117.225 113.230 ;
        RECT 91.135 112.915 91.465 112.930 ;
        RECT 116.895 112.915 117.225 112.930 ;
        RECT 65.835 112.550 66.165 112.565 ;
        RECT 69.975 112.550 70.305 112.565 ;
        RECT 65.835 112.250 70.305 112.550 ;
        RECT 65.835 112.235 66.165 112.250 ;
        RECT 69.975 112.235 70.305 112.250 ;
        RECT 103.555 112.550 103.885 112.565 ;
        RECT 124.255 112.550 124.585 112.565 ;
        RECT 103.555 112.250 124.585 112.550 ;
        RECT 103.555 112.235 103.885 112.250 ;
        RECT 124.255 112.235 124.585 112.250 ;
        RECT 28.860 111.215 30.440 111.545 ;
        RECT 134.835 110.510 135.165 110.525 ;
        RECT 140.470 110.510 144.470 110.660 ;
        RECT 134.835 110.210 144.470 110.510 ;
        RECT 134.835 110.195 135.165 110.210 ;
        RECT 140.470 110.060 144.470 110.210 ;
        RECT 32.160 108.495 33.740 108.825 ;
        RECT 136.675 107.110 137.005 107.125 ;
        RECT 140.470 107.110 144.470 107.260 ;
        RECT 136.675 106.810 144.470 107.110 ;
        RECT 136.675 106.795 137.005 106.810 ;
        RECT 140.470 106.660 144.470 106.810 ;
        RECT 28.860 105.775 30.440 106.105 ;
        RECT 120.575 105.750 120.905 105.765 ;
        RECT 131.615 105.750 131.945 105.765 ;
        RECT 120.575 105.450 131.945 105.750 ;
        RECT 120.575 105.435 120.905 105.450 ;
        RECT 131.615 105.435 131.945 105.450 ;
        RECT 84.695 105.070 85.025 105.085 ;
        RECT 133.455 105.070 133.785 105.085 ;
        RECT 84.695 104.770 133.785 105.070 ;
        RECT 84.695 104.755 85.025 104.770 ;
        RECT 133.455 104.755 133.785 104.770 ;
        RECT 84.695 103.710 85.025 103.725 ;
        RECT 115.055 103.710 115.385 103.725 ;
        RECT 84.695 103.410 115.385 103.710 ;
        RECT 84.695 103.395 85.025 103.410 ;
        RECT 115.055 103.395 115.385 103.410 ;
        RECT 136.675 103.710 137.005 103.725 ;
        RECT 140.470 103.710 144.470 103.860 ;
        RECT 136.675 103.410 144.470 103.710 ;
        RECT 136.675 103.395 137.005 103.410 ;
        RECT 32.160 103.055 33.740 103.385 ;
        RECT 140.470 103.260 144.470 103.410 ;
        RECT 28.860 100.335 30.440 100.665 ;
        RECT 136.675 100.310 137.005 100.325 ;
        RECT 140.470 100.310 144.470 100.460 ;
        RECT 136.675 100.010 144.470 100.310 ;
        RECT 136.675 99.995 137.005 100.010 ;
        RECT 140.470 99.860 144.470 100.010 ;
        RECT 32.160 97.615 33.740 97.945 ;
        RECT 108.615 96.910 108.945 96.925 ;
        RECT 110.455 96.910 110.785 96.925 ;
        RECT 108.615 96.610 110.785 96.910 ;
        RECT 108.615 96.595 108.945 96.610 ;
        RECT 110.455 96.595 110.785 96.610 ;
        RECT 134.835 96.910 135.165 96.925 ;
        RECT 140.470 96.910 144.470 97.060 ;
        RECT 134.835 96.610 144.470 96.910 ;
        RECT 134.835 96.595 135.165 96.610 ;
        RECT 140.470 96.460 144.470 96.610 ;
        RECT 95.275 96.230 95.605 96.245 ;
        RECT 125.175 96.230 125.505 96.245 ;
        RECT 95.275 95.930 125.505 96.230 ;
        RECT 95.275 95.915 95.605 95.930 ;
        RECT 125.175 95.915 125.505 95.930 ;
        RECT 28.860 94.895 30.440 95.225 ;
        RECT 106.315 94.200 106.645 94.205 ;
        RECT 106.315 94.190 106.900 94.200 ;
        RECT 110.455 94.190 110.785 94.205 ;
        RECT 127.015 94.190 127.345 94.205 ;
        RECT 106.315 93.890 107.100 94.190 ;
        RECT 110.455 93.890 127.345 94.190 ;
        RECT 106.315 93.880 106.900 93.890 ;
        RECT 106.315 93.875 106.645 93.880 ;
        RECT 110.455 93.875 110.785 93.890 ;
        RECT 127.015 93.875 127.345 93.890 ;
        RECT 136.675 93.510 137.005 93.525 ;
        RECT 140.470 93.510 144.470 93.660 ;
        RECT 136.675 93.210 144.470 93.510 ;
        RECT 136.675 93.195 137.005 93.210 ;
        RECT 140.470 93.060 144.470 93.210 ;
        RECT 104.935 92.830 105.265 92.845 ;
        RECT 112.295 92.830 112.625 92.845 ;
        RECT 104.935 92.530 112.625 92.830 ;
        RECT 104.935 92.515 105.265 92.530 ;
        RECT 112.295 92.515 112.625 92.530 ;
        RECT 32.160 92.175 33.740 92.505 ;
        RECT 106.315 92.160 106.645 92.165 ;
        RECT 106.315 92.150 106.900 92.160 ;
        RECT 106.090 91.850 106.900 92.150 ;
        RECT 106.315 91.840 106.900 91.850 ;
        RECT 108.615 92.150 108.945 92.165 ;
        RECT 115.055 92.150 115.385 92.165 ;
        RECT 108.615 91.850 115.385 92.150 ;
        RECT 106.315 91.835 106.645 91.840 ;
        RECT 108.615 91.835 108.945 91.850 ;
        RECT 115.055 91.835 115.385 91.850 ;
        RECT 92.515 91.470 92.845 91.485 ;
        RECT 93.435 91.470 93.765 91.485 ;
        RECT 118.275 91.470 118.605 91.485 ;
        RECT 92.515 91.170 118.605 91.470 ;
        RECT 92.515 91.155 92.845 91.170 ;
        RECT 93.435 91.155 93.765 91.170 ;
        RECT 118.275 91.155 118.605 91.170 ;
        RECT 110.915 90.790 111.245 90.805 ;
        RECT 113.215 90.790 113.545 90.805 ;
        RECT 110.915 90.490 113.545 90.790 ;
        RECT 110.915 90.475 111.245 90.490 ;
        RECT 113.215 90.475 113.545 90.490 ;
        RECT 136.675 90.110 137.005 90.125 ;
        RECT 140.470 90.110 144.470 90.260 ;
        RECT 136.675 89.810 144.470 90.110 ;
        RECT 136.675 89.795 137.005 89.810 ;
        RECT 28.860 89.455 30.440 89.785 ;
        RECT 140.470 89.660 144.470 89.810 ;
        RECT 32.160 86.735 33.740 87.065 ;
        RECT 47.025 56.890 47.355 56.905 ;
        RECT 50.445 56.890 54.445 57.040 ;
        RECT 47.025 56.590 54.445 56.890 ;
        RECT 47.025 56.575 47.355 56.590 ;
        RECT 50.445 56.440 54.445 56.590 ;
        RECT 44.265 53.490 44.595 53.505 ;
        RECT 50.445 53.490 54.445 53.640 ;
        RECT 44.265 53.190 54.445 53.490 ;
        RECT 44.265 53.175 44.595 53.190 ;
        RECT 50.445 53.040 54.445 53.190 ;
        RECT 28.450 51.475 30.030 51.805 ;
        RECT 45.645 50.090 45.975 50.105 ;
        RECT 50.445 50.090 54.445 50.240 ;
        RECT 45.645 49.790 54.445 50.090 ;
        RECT 45.645 49.775 45.975 49.790 ;
        RECT 50.445 49.640 54.445 49.790 ;
        RECT 31.750 48.755 33.330 49.085 ;
        RECT 23.565 48.050 23.895 48.065 ;
        RECT 27.705 48.050 28.035 48.065 ;
        RECT 41.045 48.050 41.375 48.065 ;
        RECT 23.565 47.750 41.375 48.050 ;
        RECT 23.565 47.735 23.895 47.750 ;
        RECT 27.705 47.735 28.035 47.750 ;
        RECT 41.045 47.735 41.375 47.750 ;
        RECT 7.400 46.690 11.400 46.840 ;
        RECT 24.945 46.690 25.275 46.705 ;
        RECT 7.400 46.390 25.275 46.690 ;
        RECT 7.400 46.240 11.400 46.390 ;
        RECT 24.945 46.375 25.275 46.390 ;
        RECT 47.025 46.690 47.355 46.705 ;
        RECT 50.445 46.690 54.445 46.840 ;
        RECT 47.025 46.390 54.445 46.690 ;
        RECT 47.025 46.375 47.355 46.390 ;
        RECT 28.450 46.035 30.030 46.365 ;
        RECT 50.445 46.240 54.445 46.390 ;
        RECT 7.400 43.290 11.400 43.440 ;
        RECT 31.750 43.315 33.330 43.645 ;
        RECT 13.905 43.290 14.235 43.305 ;
        RECT 7.400 42.990 14.235 43.290 ;
        RECT 7.400 42.840 11.400 42.990 ;
        RECT 13.905 42.975 14.235 42.990 ;
        RECT 47.025 43.290 47.355 43.305 ;
        RECT 50.445 43.290 54.445 43.440 ;
        RECT 47.025 42.990 54.445 43.290 ;
        RECT 47.025 42.975 47.355 42.990 ;
        RECT 50.445 42.840 54.445 42.990 ;
        RECT 28.450 40.595 30.030 40.925 ;
        RECT 44.725 39.890 45.055 39.905 ;
        RECT 50.445 39.890 54.445 40.040 ;
        RECT 44.725 39.590 54.445 39.890 ;
        RECT 44.725 39.575 45.055 39.590 ;
        RECT 50.445 39.440 54.445 39.590 ;
        RECT 31.750 37.875 33.330 38.205 ;
        RECT 7.400 36.490 11.400 36.640 ;
        RECT 13.905 36.490 14.235 36.505 ;
        RECT 7.400 36.190 14.235 36.490 ;
        RECT 7.400 36.040 11.400 36.190 ;
        RECT 13.905 36.175 14.235 36.190 ;
        RECT 47.025 36.490 47.355 36.505 ;
        RECT 50.445 36.490 54.445 36.640 ;
        RECT 47.025 36.190 54.445 36.490 ;
        RECT 47.025 36.175 47.355 36.190 ;
        RECT 50.445 36.040 54.445 36.190 ;
        RECT 28.450 35.155 30.030 35.485 ;
        RECT 41.965 33.090 42.295 33.105 ;
        RECT 50.445 33.090 54.445 33.240 ;
        RECT 41.965 32.790 54.445 33.090 ;
        RECT 41.965 32.775 42.295 32.790 ;
        RECT 31.750 32.435 33.330 32.765 ;
        RECT 50.445 32.640 54.445 32.790 ;
        RECT 7.400 29.690 11.400 29.840 ;
        RECT 28.450 29.715 30.030 30.045 ;
        RECT 13.905 29.690 14.235 29.705 ;
        RECT 7.400 29.390 14.235 29.690 ;
        RECT 7.400 29.240 11.400 29.390 ;
        RECT 13.905 29.375 14.235 29.390 ;
        RECT 39.665 29.690 39.995 29.705 ;
        RECT 50.445 29.690 54.445 29.840 ;
        RECT 39.665 29.390 54.445 29.690 ;
        RECT 39.665 29.375 39.995 29.390 ;
        RECT 50.445 29.240 54.445 29.390 ;
        RECT 31.750 26.995 33.330 27.325 ;
        RECT 43.345 26.290 43.675 26.305 ;
        RECT 50.445 26.290 54.445 26.440 ;
        RECT 43.345 25.990 54.445 26.290 ;
        RECT 43.345 25.975 43.675 25.990 ;
        RECT 50.445 25.840 54.445 25.990 ;
        RECT 28.450 24.275 30.030 24.605 ;
        RECT 41.045 22.890 41.375 22.905 ;
        RECT 50.445 22.890 54.445 23.040 ;
        RECT 41.045 22.590 54.445 22.890 ;
        RECT 41.045 22.575 41.375 22.590 ;
        RECT 50.445 22.440 54.445 22.590 ;
        RECT 31.750 21.555 33.330 21.885 ;
        RECT 11.605 20.170 11.935 20.185 ;
        RECT 11.390 19.855 11.935 20.170 ;
        RECT 11.390 19.640 11.690 19.855 ;
        RECT 7.400 19.190 11.690 19.640 ;
        RECT 38.285 19.490 38.615 19.505 ;
        RECT 50.445 19.490 54.445 19.640 ;
        RECT 38.285 19.190 54.445 19.490 ;
        RECT 7.400 19.040 11.400 19.190 ;
        RECT 38.285 19.175 38.615 19.190 ;
        RECT 28.450 18.835 30.030 19.165 ;
        RECT 50.445 19.040 54.445 19.190 ;
        RECT 31.750 16.115 33.330 16.445 ;
        RECT 42.885 16.090 43.215 16.105 ;
        RECT 50.445 16.090 54.445 16.240 ;
        RECT 42.885 15.790 54.445 16.090 ;
        RECT 42.885 15.775 43.215 15.790 ;
        RECT 50.445 15.640 54.445 15.790 ;
        RECT 46.565 12.690 46.895 12.705 ;
        RECT 50.445 12.690 54.445 12.840 ;
        RECT 46.565 12.390 54.445 12.690 ;
        RECT 46.565 12.375 46.895 12.390 ;
        RECT 50.445 12.240 54.445 12.390 ;
      LAYER met4 ;
        RECT 64.090 225.055 64.145 225.385 ;
        RECT 66.455 224.965 66.550 225.295 ;
        RECT 69.305 225.135 69.310 225.465 ;
        RECT 69.610 225.135 69.635 225.465 ;
        RECT 71.995 224.895 72.070 225.225 ;
        RECT 74.785 224.945 74.830 225.275 ;
        RECT 77.515 224.760 77.590 225.085 ;
        RECT 80.295 224.925 80.350 225.255 ;
        RECT 83.025 224.760 83.110 225.085 ;
        RECT 85.795 224.915 85.870 225.245 ;
        RECT 88.535 224.915 88.630 225.245 ;
        RECT 91.350 224.835 91.390 225.165 ;
        RECT 94.125 224.815 94.150 225.145 ;
        RECT 94.450 224.815 94.455 225.145 ;
        RECT 144.130 225.115 144.225 225.445 ;
        RECT 77.515 224.755 77.845 224.760 ;
        RECT 83.025 224.755 83.355 224.760 ;
        RECT 6.000 197.560 6.140 199.160 ;
        RECT 28.850 86.660 30.450 212.260 ;
        RECT 31.105 172.075 31.435 172.405 ;
        RECT 31.120 135.005 31.420 172.075 ;
        RECT 31.105 134.675 31.435 135.005 ;
        RECT 32.150 86.660 33.750 212.260 ;
        RECT 75.265 193.155 75.595 193.485 ;
        RECT 75.280 168.325 75.580 193.155 ;
        RECT 113.905 191.115 114.235 191.445 ;
        RECT 113.920 179.205 114.220 191.115 ;
        RECT 117.585 179.555 117.915 179.885 ;
        RECT 113.905 178.875 114.235 179.205 ;
        RECT 75.265 167.995 75.595 168.325 ;
        RECT 117.600 154.045 117.900 179.555 ;
        RECT 117.585 153.715 117.915 154.045 ;
        RECT 106.545 93.875 106.875 94.205 ;
        RECT 106.560 92.165 106.860 93.875 ;
        RECT 106.545 91.835 106.875 92.165 ;
        RECT 28.440 16.040 30.040 51.880 ;
        RECT 31.740 16.040 33.340 51.880 ;
        RECT 151.950 1.000 152.575 9.470 ;
  END
END tt_um_tim2305_adc_dac
END LIBRARY

