VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_tim2305_adc_dac
  CLASS BLOCK ;
  FOREIGN tt_um_tim2305_adc_dac ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 256.000000 ;
    ANTENNADIFFAREA 4.850000 ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 112.465 219.150 113.275 219.290 ;
        RECT 112.275 218.980 113.275 219.150 ;
        RECT 112.465 217.920 113.275 218.980 ;
        RECT 112.465 217.770 113.275 217.910 ;
        RECT 112.275 217.600 113.275 217.770 ;
        RECT 112.465 212.400 113.275 217.600 ;
        RECT 112.465 212.250 113.275 212.390 ;
        RECT 112.275 212.080 113.275 212.250 ;
        RECT 112.465 208.720 113.275 212.080 ;
        RECT 112.305 208.455 112.415 208.575 ;
        RECT 112.465 208.110 113.145 208.250 ;
        RECT 112.275 207.940 113.145 208.110 ;
        RECT 112.465 207.765 113.145 207.940 ;
        RECT 112.465 206.420 113.375 207.765 ;
        RECT 112.550 205.970 113.335 206.400 ;
        RECT 112.305 205.695 112.415 205.815 ;
        RECT 112.465 204.145 113.375 205.490 ;
        RECT 112.465 203.970 113.145 204.145 ;
        RECT 112.275 203.800 113.145 203.970 ;
        RECT 112.465 203.660 113.145 203.800 ;
        RECT 112.465 203.510 113.145 203.650 ;
        RECT 112.275 203.340 113.145 203.510 ;
      LAYER nwell ;
        RECT 13.190 199.945 92.230 201.550 ;
      LAYER pwell ;
        RECT 112.465 200.135 113.145 203.340 ;
        RECT 13.385 198.745 14.755 199.555 ;
        RECT 14.765 198.745 20.275 199.555 ;
        RECT 20.285 198.745 25.795 199.555 ;
        RECT 26.275 198.830 26.705 199.615 ;
        RECT 26.725 198.745 32.235 199.555 ;
        RECT 32.245 198.745 37.755 199.555 ;
        RECT 37.765 198.745 39.135 199.555 ;
        RECT 39.155 198.830 39.585 199.615 ;
        RECT 39.605 198.745 45.115 199.555 ;
        RECT 45.125 198.745 50.635 199.555 ;
        RECT 50.645 198.745 52.015 199.555 ;
        RECT 52.035 198.830 52.465 199.615 ;
        RECT 52.485 198.745 57.995 199.555 ;
        RECT 58.005 199.425 58.925 199.655 ;
        RECT 58.005 198.745 60.295 199.425 ;
        RECT 60.305 198.745 63.055 199.555 ;
        RECT 63.065 198.745 64.435 199.525 ;
        RECT 64.915 198.830 65.345 199.615 ;
        RECT 65.365 198.745 70.875 199.555 ;
        RECT 70.885 198.745 72.715 199.555 ;
        RECT 72.725 198.745 74.095 199.525 ;
        RECT 74.105 198.745 77.775 199.555 ;
        RECT 77.795 198.830 78.225 199.615 ;
        RECT 78.245 198.745 83.755 199.555 ;
        RECT 83.765 198.745 89.275 199.555 ;
        RECT 89.285 198.745 90.655 199.555 ;
        RECT 90.665 198.745 92.035 199.555 ;
        RECT 112.465 199.225 113.365 200.135 ;
        RECT 13.525 198.535 13.695 198.745 ;
        RECT 14.905 198.535 15.075 198.745 ;
        RECT 20.425 198.535 20.595 198.745 ;
        RECT 25.945 198.695 26.115 198.725 ;
        RECT 25.940 198.585 26.115 198.695 ;
        RECT 25.945 198.535 26.115 198.585 ;
        RECT 26.865 198.555 27.035 198.745 ;
        RECT 31.465 198.535 31.635 198.725 ;
        RECT 32.385 198.555 32.555 198.745 ;
        RECT 36.985 198.535 37.155 198.725 ;
        RECT 37.905 198.555 38.075 198.745 ;
        RECT 38.820 198.585 38.940 198.695 ;
        RECT 39.745 198.535 39.915 198.745 ;
        RECT 43.420 198.535 43.590 198.725 ;
        RECT 43.885 198.535 44.055 198.725 ;
        RECT 45.265 198.555 45.435 198.745 ;
        RECT 46.185 198.535 46.355 198.725 ;
        RECT 50.785 198.555 50.955 198.745 ;
        RECT 52.625 198.555 52.795 198.745 ;
        RECT 53.545 198.535 53.715 198.725 ;
        RECT 57.225 198.535 57.395 198.725 ;
        RECT 59.985 198.555 60.155 198.745 ;
        RECT 60.445 198.555 60.615 198.745 ;
        RECT 63.205 198.555 63.375 198.745 ;
        RECT 64.580 198.585 64.700 198.695 ;
        RECT 65.505 198.535 65.675 198.745 ;
        RECT 67.340 198.585 67.460 198.695 ;
        RECT 71.025 198.555 71.195 198.745 ;
        RECT 73.785 198.555 73.955 198.745 ;
        RECT 74.245 198.555 74.415 198.745 ;
        RECT 74.705 198.535 74.875 198.725 ;
        RECT 75.165 198.535 75.335 198.725 ;
        RECT 78.385 198.555 78.555 198.745 ;
        RECT 80.685 198.535 80.855 198.725 ;
        RECT 83.905 198.555 84.075 198.745 ;
        RECT 86.205 198.535 86.375 198.725 ;
        RECT 89.425 198.555 89.595 198.745 ;
        RECT 89.895 198.580 90.055 198.690 ;
        RECT 91.725 198.535 91.895 198.745 ;
        RECT 13.385 197.725 14.755 198.535 ;
        RECT 14.765 197.725 20.275 198.535 ;
        RECT 20.285 197.725 25.795 198.535 ;
        RECT 25.805 197.725 31.315 198.535 ;
        RECT 31.325 197.725 36.835 198.535 ;
        RECT 36.845 197.725 38.675 198.535 ;
        RECT 39.155 197.665 39.585 198.450 ;
        RECT 39.605 197.725 42.355 198.535 ;
        RECT 42.385 197.625 43.735 198.535 ;
        RECT 43.745 197.855 46.035 198.535 ;
        RECT 46.045 197.855 53.355 198.535 ;
        RECT 45.115 197.625 46.035 197.855 ;
        RECT 49.560 197.635 50.470 197.855 ;
        RECT 52.005 197.625 53.355 197.855 ;
        RECT 53.405 197.725 57.075 198.535 ;
        RECT 57.085 197.855 64.395 198.535 ;
        RECT 60.600 197.635 61.510 197.855 ;
        RECT 63.045 197.625 64.395 197.855 ;
        RECT 64.915 197.665 65.345 198.450 ;
        RECT 65.365 197.725 67.195 198.535 ;
        RECT 67.705 197.855 75.015 198.535 ;
        RECT 67.705 197.625 69.055 197.855 ;
        RECT 70.590 197.635 71.500 197.855 ;
        RECT 75.025 197.725 80.535 198.535 ;
        RECT 80.545 197.725 86.055 198.535 ;
        RECT 86.065 197.725 89.735 198.535 ;
        RECT 90.665 197.725 92.035 198.535 ;
        RECT 112.465 197.690 113.145 199.225 ;
      LAYER nwell ;
        RECT 13.190 194.505 92.230 197.335 ;
      LAYER pwell ;
        RECT 112.465 196.340 113.375 197.690 ;
        RECT 112.465 194.945 113.375 196.290 ;
        RECT 112.465 194.770 113.145 194.945 ;
        RECT 112.275 194.600 113.145 194.770 ;
        RECT 112.465 194.460 113.145 194.600 ;
        RECT 13.385 193.305 14.755 194.115 ;
        RECT 14.765 193.305 20.275 194.115 ;
        RECT 20.285 193.305 25.795 194.115 ;
        RECT 26.275 193.390 26.705 194.175 ;
        RECT 26.725 193.305 32.235 194.115 ;
        RECT 32.245 193.305 37.755 194.115 ;
        RECT 41.740 193.985 42.650 194.205 ;
        RECT 44.185 193.985 45.535 194.215 ;
        RECT 38.225 193.305 45.535 193.985 ;
        RECT 46.045 193.985 46.965 194.215 ;
        RECT 46.045 193.305 48.335 193.985 ;
        RECT 48.345 193.305 49.695 194.215 ;
        RECT 51.095 193.985 52.015 194.215 ;
        RECT 49.725 193.305 52.015 193.985 ;
        RECT 52.035 193.390 52.465 194.175 ;
        RECT 56.000 193.985 56.910 194.205 ;
        RECT 58.445 193.985 59.795 194.215 ;
        RECT 52.485 193.305 59.795 193.985 ;
        RECT 60.785 193.305 62.135 194.215 ;
        RECT 63.085 193.305 64.435 194.215 ;
        RECT 64.445 193.305 65.815 194.115 ;
        RECT 65.845 193.305 67.195 194.215 ;
        RECT 68.575 193.985 69.495 194.215 ;
        RECT 67.205 193.305 69.495 193.985 ;
        RECT 70.465 193.985 71.815 194.215 ;
        RECT 73.350 193.985 74.260 194.205 ;
        RECT 70.465 193.305 77.775 193.985 ;
        RECT 77.795 193.390 78.225 194.175 ;
        RECT 112.310 194.140 112.420 194.300 ;
        RECT 78.245 193.305 83.755 194.115 ;
        RECT 83.765 193.305 89.275 194.115 ;
        RECT 89.285 193.305 90.655 194.115 ;
        RECT 90.665 193.305 92.035 194.115 ;
        RECT 13.525 193.095 13.695 193.305 ;
        RECT 14.905 193.095 15.075 193.305 ;
        RECT 20.425 193.095 20.595 193.305 ;
        RECT 25.945 193.255 26.115 193.285 ;
        RECT 25.940 193.145 26.115 193.255 ;
        RECT 25.945 193.095 26.115 193.145 ;
        RECT 26.865 193.115 27.035 193.305 ;
        RECT 31.465 193.095 31.635 193.285 ;
        RECT 32.385 193.115 32.555 193.305 ;
        RECT 36.985 193.095 37.155 193.285 ;
        RECT 37.900 193.145 38.020 193.255 ;
        RECT 38.365 193.115 38.535 193.305 ;
        RECT 38.820 193.145 38.940 193.255 ;
        RECT 39.745 193.095 39.915 193.285 ;
        RECT 42.965 193.095 43.135 193.285 ;
        RECT 43.430 193.095 43.600 193.285 ;
        RECT 44.805 193.095 44.975 193.285 ;
        RECT 45.720 193.145 45.840 193.255 ;
        RECT 48.025 193.095 48.195 193.305 ;
        RECT 48.490 193.115 48.660 193.305 ;
        RECT 49.865 193.115 50.035 193.305 ;
        RECT 52.625 193.095 52.795 193.305 ;
        RECT 53.085 193.095 53.255 193.285 ;
        RECT 58.605 193.095 58.775 193.285 ;
        RECT 59.995 193.150 60.155 193.260 ;
        RECT 61.820 193.115 61.990 193.305 ;
        RECT 62.295 193.150 62.455 193.260 ;
        RECT 64.120 193.115 64.290 193.305 ;
        RECT 64.585 193.095 64.755 193.305 ;
        RECT 65.505 193.095 65.675 193.285 ;
        RECT 66.880 193.115 67.050 193.305 ;
        RECT 67.345 193.115 67.515 193.305 ;
        RECT 68.725 193.095 68.895 193.285 ;
        RECT 69.655 193.150 69.815 193.260 ;
        RECT 70.565 193.095 70.735 193.285 ;
        RECT 73.785 193.115 73.955 193.285 ;
        RECT 73.790 193.095 73.955 193.115 ;
        RECT 76.085 193.095 76.255 193.285 ;
        RECT 77.465 193.115 77.635 193.305 ;
        RECT 78.385 193.115 78.555 193.305 ;
        RECT 81.605 193.095 81.775 193.285 ;
        RECT 83.905 193.115 84.075 193.305 ;
        RECT 87.125 193.095 87.295 193.285 ;
        RECT 89.425 193.115 89.595 193.305 ;
        RECT 91.725 193.095 91.895 193.305 ;
        RECT 13.385 192.285 14.755 193.095 ;
        RECT 14.765 192.285 20.275 193.095 ;
        RECT 20.285 192.285 25.795 193.095 ;
        RECT 25.805 192.285 31.315 193.095 ;
        RECT 31.325 192.285 36.835 193.095 ;
        RECT 36.845 192.285 38.675 193.095 ;
        RECT 39.155 192.225 39.585 193.010 ;
        RECT 39.605 192.285 40.975 193.095 ;
        RECT 40.985 192.415 43.275 193.095 ;
        RECT 40.985 192.185 41.905 192.415 ;
        RECT 43.285 192.185 44.635 193.095 ;
        RECT 44.665 192.415 47.875 193.095 ;
        RECT 46.740 192.185 47.875 192.415 ;
        RECT 47.900 192.185 49.715 193.095 ;
        RECT 49.725 192.185 52.895 193.095 ;
        RECT 52.945 192.285 58.455 193.095 ;
        RECT 58.465 192.285 62.135 193.095 ;
        RECT 62.155 192.415 64.895 193.095 ;
        RECT 64.915 192.225 65.345 193.010 ;
        RECT 65.365 192.415 68.575 193.095 ;
        RECT 67.440 192.185 68.575 192.415 ;
        RECT 68.600 192.185 70.415 193.095 ;
        RECT 70.425 192.415 73.635 193.095 ;
        RECT 73.790 192.415 75.625 193.095 ;
        RECT 72.500 192.185 73.635 192.415 ;
        RECT 74.695 192.185 75.625 192.415 ;
        RECT 75.945 192.285 81.455 193.095 ;
        RECT 81.465 192.285 86.975 193.095 ;
        RECT 86.985 192.285 90.655 193.095 ;
        RECT 90.665 192.285 92.035 193.095 ;
        RECT 112.550 193.090 113.335 193.520 ;
        RECT 112.310 192.760 112.420 192.920 ;
        RECT 112.465 192.010 113.145 192.150 ;
      LAYER nwell ;
        RECT 13.190 189.065 92.230 191.895 ;
      LAYER pwell ;
        RECT 112.275 191.840 113.145 192.010 ;
        RECT 112.465 191.665 113.145 191.840 ;
        RECT 112.465 190.320 113.375 191.665 ;
        RECT 112.465 189.260 113.245 190.310 ;
        RECT 112.275 189.090 113.245 189.260 ;
        RECT 112.465 188.940 113.245 189.090 ;
        RECT 13.385 187.865 14.755 188.675 ;
        RECT 14.765 187.865 20.275 188.675 ;
        RECT 20.285 187.865 25.795 188.675 ;
        RECT 26.275 187.950 26.705 188.735 ;
        RECT 26.725 187.865 32.235 188.675 ;
        RECT 32.245 187.865 37.755 188.675 ;
        RECT 37.765 187.865 41.435 188.675 ;
        RECT 41.445 188.545 42.365 188.775 ;
        RECT 41.445 187.865 43.735 188.545 ;
        RECT 43.745 187.865 49.255 188.675 ;
        RECT 49.265 187.865 52.015 188.675 ;
        RECT 52.035 187.950 52.465 188.735 ;
        RECT 52.485 187.865 56.155 188.675 ;
        RECT 57.085 187.865 58.900 188.775 ;
        RECT 58.925 187.865 62.135 188.775 ;
        RECT 62.145 187.865 64.895 188.775 ;
        RECT 65.365 188.545 66.285 188.775 ;
        RECT 65.365 187.865 67.655 188.545 ;
        RECT 67.665 187.865 70.415 188.675 ;
        RECT 70.905 187.865 72.255 188.775 ;
        RECT 72.265 187.865 77.775 188.675 ;
        RECT 77.795 187.950 78.225 188.735 ;
        RECT 78.245 187.865 83.755 188.675 ;
        RECT 83.765 187.865 89.275 188.675 ;
        RECT 89.285 187.865 90.655 188.675 ;
        RECT 90.665 187.865 92.035 188.675 ;
        RECT 112.310 188.620 112.420 188.780 ;
        RECT 112.465 187.870 113.145 188.010 ;
        RECT 13.525 187.655 13.695 187.865 ;
        RECT 14.905 187.655 15.075 187.865 ;
        RECT 20.425 187.655 20.595 187.865 ;
        RECT 23.645 187.655 23.815 187.845 ;
        RECT 24.105 187.655 24.275 187.845 ;
        RECT 25.940 187.705 26.060 187.815 ;
        RECT 26.865 187.675 27.035 187.865 ;
        RECT 27.785 187.655 27.955 187.845 ;
        RECT 32.385 187.675 32.555 187.865 ;
        RECT 35.145 187.655 35.315 187.845 ;
        RECT 37.905 187.675 38.075 187.865 ;
        RECT 38.820 187.705 38.940 187.815 ;
        RECT 39.745 187.655 39.915 187.845 ;
        RECT 43.425 187.675 43.595 187.865 ;
        RECT 43.885 187.675 44.055 187.865 ;
        RECT 47.105 187.655 47.275 187.845 ;
        RECT 49.405 187.675 49.575 187.865 ;
        RECT 52.625 187.655 52.795 187.865 ;
        RECT 56.315 187.815 56.475 187.820 ;
        RECT 56.300 187.710 56.475 187.815 ;
        RECT 56.300 187.705 56.420 187.710 ;
        RECT 58.145 187.655 58.315 187.845 ;
        RECT 58.605 187.655 58.775 187.865 ;
        RECT 59.065 187.675 59.235 187.865 ;
        RECT 60.440 187.705 60.560 187.815 ;
        RECT 60.910 187.655 61.080 187.845 ;
        RECT 62.285 187.675 62.455 187.865 ;
        RECT 62.745 187.655 62.915 187.845 ;
        RECT 64.580 187.705 64.700 187.815 ;
        RECT 65.040 187.705 65.160 187.815 ;
        RECT 65.505 187.655 65.675 187.845 ;
        RECT 67.345 187.675 67.515 187.865 ;
        RECT 67.805 187.675 67.975 187.865 ;
        RECT 71.020 187.845 71.190 187.865 ;
        RECT 70.560 187.705 70.680 187.815 ;
        RECT 71.020 187.675 71.195 187.845 ;
        RECT 72.405 187.675 72.575 187.865 ;
        RECT 71.025 187.655 71.195 187.675 ;
        RECT 76.545 187.655 76.715 187.845 ;
        RECT 78.385 187.675 78.555 187.865 ;
        RECT 82.065 187.655 82.235 187.845 ;
        RECT 83.905 187.675 84.075 187.865 ;
        RECT 87.585 187.655 87.755 187.845 ;
        RECT 89.425 187.675 89.595 187.865 ;
        RECT 90.340 187.705 90.460 187.815 ;
        RECT 91.725 187.655 91.895 187.865 ;
        RECT 112.275 187.700 113.145 187.870 ;
        RECT 13.385 186.845 14.755 187.655 ;
        RECT 14.765 186.845 20.275 187.655 ;
        RECT 20.285 186.845 21.655 187.655 ;
        RECT 21.665 186.975 23.955 187.655 ;
        RECT 21.665 186.745 22.585 186.975 ;
        RECT 23.965 186.845 27.635 187.655 ;
        RECT 27.645 186.975 34.955 187.655 ;
        RECT 31.160 186.755 32.070 186.975 ;
        RECT 33.605 186.745 34.955 186.975 ;
        RECT 35.005 186.845 38.675 187.655 ;
        RECT 39.155 186.785 39.585 187.570 ;
        RECT 39.605 186.975 46.915 187.655 ;
        RECT 43.120 186.755 44.030 186.975 ;
        RECT 45.565 186.745 46.915 186.975 ;
        RECT 46.965 186.845 52.475 187.655 ;
        RECT 52.485 186.845 56.155 187.655 ;
        RECT 56.625 186.745 58.440 187.655 ;
        RECT 58.465 186.845 60.295 187.655 ;
        RECT 60.765 186.745 62.595 187.655 ;
        RECT 62.605 186.845 64.435 187.655 ;
        RECT 64.915 186.785 65.345 187.570 ;
        RECT 65.365 186.845 70.875 187.655 ;
        RECT 70.885 186.845 76.395 187.655 ;
        RECT 76.405 186.845 81.915 187.655 ;
        RECT 81.925 186.845 87.435 187.655 ;
        RECT 87.445 186.845 90.195 187.655 ;
        RECT 90.665 186.845 92.035 187.655 ;
      LAYER nwell ;
        RECT 13.190 183.625 92.230 186.455 ;
      LAYER pwell ;
        RECT 112.465 186.190 113.145 187.700 ;
        RECT 112.465 185.260 113.375 186.190 ;
        RECT 112.305 184.995 112.415 185.115 ;
        RECT 112.465 183.730 113.275 184.790 ;
        RECT 112.275 183.560 113.275 183.730 ;
        RECT 112.465 183.420 113.275 183.560 ;
        RECT 13.385 182.425 14.755 183.235 ;
        RECT 14.765 182.425 17.515 183.235 ;
        RECT 17.545 182.425 18.895 183.335 ;
        RECT 18.945 183.105 20.295 183.335 ;
        RECT 21.830 183.105 22.740 183.325 ;
        RECT 18.945 182.425 26.255 183.105 ;
        RECT 26.275 182.510 26.705 183.295 ;
        RECT 27.645 183.105 28.565 183.335 ;
        RECT 27.645 182.425 29.935 183.105 ;
        RECT 29.945 182.425 32.865 183.335 ;
        RECT 33.175 182.425 35.905 183.335 ;
        RECT 36.125 183.245 37.075 183.335 ;
        RECT 36.125 182.425 38.055 183.245 ;
        RECT 38.225 182.425 40.055 183.335 ;
        RECT 40.105 182.425 43.275 183.335 ;
        RECT 43.285 182.425 46.955 183.235 ;
        RECT 46.965 182.425 48.795 183.105 ;
        RECT 48.805 182.425 51.555 183.235 ;
        RECT 52.035 182.510 52.465 183.295 ;
        RECT 52.495 182.425 55.225 183.335 ;
        RECT 55.245 182.425 58.915 183.235 ;
        RECT 59.385 182.425 63.045 183.335 ;
        RECT 63.265 183.245 64.215 183.335 ;
        RECT 63.265 182.425 65.195 183.245 ;
        RECT 65.375 182.425 66.725 183.335 ;
        RECT 67.205 183.135 68.135 183.335 ;
        RECT 69.465 183.135 70.415 183.335 ;
        RECT 67.205 182.655 70.415 183.135 ;
        RECT 67.350 182.455 70.415 182.655 ;
        RECT 13.525 182.215 13.695 182.425 ;
        RECT 14.905 182.215 15.075 182.425 ;
        RECT 17.660 182.235 17.830 182.425 ;
        RECT 20.425 182.215 20.595 182.405 ;
        RECT 24.105 182.235 24.275 182.405 ;
        RECT 24.105 182.215 24.270 182.235 ;
        RECT 24.565 182.215 24.735 182.405 ;
        RECT 25.945 182.235 26.115 182.425 ;
        RECT 26.875 182.270 27.035 182.380 ;
        RECT 29.625 182.235 29.795 182.425 ;
        RECT 30.090 182.375 30.260 182.425 ;
        RECT 30.080 182.265 30.260 182.375 ;
        RECT 30.090 182.235 30.260 182.265 ;
        RECT 33.305 182.215 33.475 182.425 ;
        RECT 37.905 182.405 38.055 182.425 ;
        RECT 33.760 182.265 33.880 182.375 ;
        RECT 34.225 182.215 34.395 182.405 ;
        RECT 37.445 182.215 37.615 182.405 ;
        RECT 37.905 182.235 38.075 182.405 ;
        RECT 39.740 182.370 39.910 182.425 ;
        RECT 39.740 182.260 39.915 182.370 ;
        RECT 39.740 182.235 39.910 182.260 ;
        RECT 40.205 182.235 40.375 182.425 ;
        RECT 40.665 182.215 40.835 182.405 ;
        RECT 43.425 182.235 43.595 182.425 ;
        RECT 44.810 182.215 44.980 182.405 ;
        RECT 45.265 182.235 45.435 182.405 ;
        RECT 45.270 182.215 45.435 182.235 ;
        RECT 47.565 182.215 47.735 182.405 ;
        RECT 48.485 182.235 48.655 182.425 ;
        RECT 48.945 182.235 49.115 182.425 ;
        RECT 51.250 182.215 51.420 182.405 ;
        RECT 51.700 182.265 51.820 182.375 ;
        RECT 52.625 182.235 52.795 182.425 ;
        RECT 55.385 182.235 55.555 182.425 ;
        RECT 57.220 182.215 57.390 182.405 ;
        RECT 57.685 182.215 57.855 182.405 ;
        RECT 59.060 182.265 59.180 182.375 ;
        RECT 61.360 182.265 61.480 182.375 ;
        RECT 13.385 181.405 14.755 182.215 ;
        RECT 14.765 181.405 20.275 182.215 ;
        RECT 20.285 181.405 22.115 182.215 ;
        RECT 22.435 181.535 24.270 182.215 ;
        RECT 22.435 181.305 23.365 181.535 ;
        RECT 24.425 181.405 29.935 182.215 ;
        RECT 30.405 181.535 33.615 182.215 ;
        RECT 30.405 181.305 31.540 181.535 ;
        RECT 34.165 181.305 37.165 182.215 ;
        RECT 37.305 181.405 39.135 182.215 ;
        RECT 39.155 181.345 39.585 182.130 ;
        RECT 40.625 181.305 43.735 182.215 ;
        RECT 43.745 181.305 45.095 182.215 ;
        RECT 45.270 181.535 47.105 182.215 ;
        RECT 47.425 181.535 51.095 182.215 ;
        RECT 46.175 181.305 47.105 181.535 ;
        RECT 50.165 181.305 51.095 181.535 ;
        RECT 51.105 181.305 52.935 182.215 ;
        RECT 53.145 181.305 57.535 182.215 ;
        RECT 57.545 181.305 61.215 182.215 ;
        RECT 61.825 182.185 61.995 182.405 ;
        RECT 62.750 182.235 62.920 182.425 ;
        RECT 65.045 182.405 65.195 182.425 ;
        RECT 65.045 182.235 65.215 182.405 ;
        RECT 65.505 182.235 65.675 182.425 ;
        RECT 66.880 182.265 67.000 182.375 ;
        RECT 67.350 182.235 67.520 182.455 ;
        RECT 69.480 182.425 70.415 182.455 ;
        RECT 70.465 183.105 71.815 183.335 ;
        RECT 73.350 183.105 74.260 183.325 ;
        RECT 70.465 182.425 77.775 183.105 ;
        RECT 77.795 182.510 78.225 183.295 ;
        RECT 78.245 182.425 83.755 183.235 ;
        RECT 83.765 182.425 89.275 183.235 ;
        RECT 89.285 182.425 90.655 183.235 ;
        RECT 90.665 182.425 92.035 183.235 ;
      LAYER nwell ;
        RECT 113.665 183.225 116.495 219.485 ;
      LAYER pwell ;
        RECT 116.885 219.150 117.695 219.290 ;
        RECT 117.905 219.150 118.715 219.290 ;
        RECT 116.885 218.980 118.715 219.150 ;
        RECT 116.885 217.920 117.695 218.980 ;
        RECT 117.905 217.920 118.715 218.980 ;
        RECT 116.785 216.565 117.695 217.910 ;
        RECT 117.015 216.390 117.695 216.565 ;
        RECT 117.905 216.520 118.815 217.870 ;
        RECT 117.015 216.220 117.885 216.390 ;
        RECT 117.015 216.080 117.695 216.220 ;
        RECT 117.740 215.760 117.850 215.920 ;
        RECT 116.785 214.735 117.695 215.150 ;
        RECT 117.905 214.985 118.585 216.520 ;
        RECT 116.785 214.565 117.885 214.735 ;
        RECT 116.785 214.220 117.695 214.565 ;
        RECT 117.015 211.250 117.695 214.220 ;
        RECT 117.905 214.075 118.805 214.985 ;
        RECT 116.885 210.870 117.695 211.010 ;
        RECT 117.905 210.870 118.585 214.075 ;
        RECT 116.885 210.700 118.585 210.870 ;
        RECT 116.885 207.340 117.695 210.700 ;
        RECT 117.905 210.560 118.585 210.700 ;
        RECT 117.905 210.410 118.715 210.550 ;
        RECT 117.715 210.240 118.715 210.410 ;
        RECT 116.885 207.190 117.695 207.330 ;
        RECT 116.885 207.020 117.885 207.190 ;
        RECT 116.885 205.960 117.695 207.020 ;
        RECT 117.905 206.880 118.715 210.240 ;
        RECT 117.745 206.615 117.855 206.735 ;
        RECT 117.990 205.970 118.775 206.400 ;
        RECT 116.785 204.560 117.695 205.910 ;
        RECT 117.905 205.810 118.585 205.950 ;
        RECT 117.715 205.640 118.585 205.810 ;
        RECT 117.015 203.025 117.695 204.560 ;
        RECT 116.795 202.115 117.695 203.025 ;
        RECT 117.015 198.910 117.695 202.115 ;
        RECT 117.015 198.740 117.885 198.910 ;
        RECT 117.015 198.600 117.695 198.740 ;
        RECT 116.785 198.175 117.695 198.590 ;
        RECT 116.785 198.005 117.885 198.175 ;
        RECT 116.785 197.660 117.695 198.005 ;
        RECT 117.015 194.690 117.695 197.660 ;
        RECT 117.905 196.845 118.585 205.640 ;
        RECT 117.905 196.610 118.715 196.750 ;
        RECT 117.715 196.440 118.715 196.610 ;
        RECT 117.905 195.380 118.715 196.440 ;
        RECT 117.905 195.230 118.685 195.370 ;
        RECT 117.715 195.060 118.685 195.230 ;
        RECT 117.740 194.140 117.850 194.300 ;
        RECT 117.905 194.000 118.685 195.060 ;
        RECT 117.905 193.850 118.685 193.990 ;
        RECT 117.715 193.680 118.685 193.850 ;
        RECT 116.825 193.090 117.610 193.520 ;
        RECT 116.785 192.055 117.695 192.975 ;
        RECT 117.905 192.620 118.685 193.680 ;
        RECT 117.905 192.470 118.685 192.610 ;
        RECT 117.715 192.300 118.685 192.470 ;
        RECT 117.015 189.710 117.695 192.055 ;
        RECT 117.905 191.240 118.685 192.300 ;
        RECT 117.905 191.090 118.685 191.230 ;
        RECT 117.715 190.920 118.685 191.090 ;
        RECT 117.905 189.860 118.685 190.920 ;
        RECT 117.015 189.540 117.885 189.710 ;
        RECT 117.015 189.510 117.695 189.540 ;
        RECT 117.740 189.080 117.850 189.240 ;
        RECT 117.905 188.795 118.815 189.830 ;
        RECT 117.715 188.625 118.815 188.795 ;
        RECT 117.905 188.480 118.815 188.625 ;
        RECT 116.785 186.030 117.695 188.470 ;
        RECT 117.905 188.330 118.815 188.390 ;
        RECT 117.715 188.160 118.815 188.330 ;
        RECT 116.785 185.860 117.885 186.030 ;
        RECT 116.785 185.720 117.695 185.860 ;
        RECT 117.740 185.400 117.850 185.560 ;
        RECT 117.905 184.940 118.815 188.160 ;
        RECT 116.885 183.730 117.695 184.790 ;
        RECT 117.905 183.730 118.715 184.790 ;
        RECT 116.885 183.560 118.715 183.730 ;
        RECT 116.885 183.420 117.695 183.560 ;
        RECT 117.905 183.420 118.715 183.560 ;
      LAYER nwell ;
        RECT 119.105 183.225 121.935 219.485 ;
      LAYER pwell ;
        RECT 122.325 219.150 123.135 219.290 ;
        RECT 123.345 219.150 124.155 219.290 ;
        RECT 122.325 218.980 124.155 219.150 ;
        RECT 122.325 217.920 123.135 218.980 ;
        RECT 123.345 217.920 124.155 218.980 ;
        RECT 122.225 216.565 123.135 217.910 ;
        RECT 123.345 217.770 124.025 217.910 ;
        RECT 123.155 217.600 124.025 217.770 ;
        RECT 122.455 216.390 123.135 216.565 ;
        RECT 122.455 216.220 123.325 216.390 ;
        RECT 122.455 216.080 123.135 216.220 ;
        RECT 123.180 215.760 123.290 215.920 ;
        RECT 122.455 215.010 123.135 215.040 ;
        RECT 122.455 214.840 123.325 215.010 ;
        RECT 122.455 212.495 123.135 214.840 ;
        RECT 122.225 211.575 123.135 212.495 ;
        RECT 123.345 214.395 124.025 217.600 ;
        RECT 123.345 213.485 124.245 214.395 ;
        RECT 123.345 211.950 124.025 213.485 ;
        RECT 123.180 211.160 123.290 211.320 ;
        RECT 123.345 210.600 124.255 211.950 ;
        RECT 122.455 210.410 123.135 210.440 ;
        RECT 123.345 210.410 124.155 210.550 ;
        RECT 122.455 210.240 124.155 210.410 ;
        RECT 122.455 207.895 123.135 210.240 ;
        RECT 122.225 206.975 123.135 207.895 ;
        RECT 123.345 206.880 124.155 210.240 ;
        RECT 122.455 203.670 123.135 206.640 ;
        RECT 123.185 206.615 123.295 206.735 ;
        RECT 123.430 205.970 124.215 206.400 ;
        RECT 123.345 205.810 124.025 205.950 ;
        RECT 123.155 205.640 124.025 205.810 ;
        RECT 122.225 203.325 123.135 203.670 ;
        RECT 122.225 203.155 123.325 203.325 ;
        RECT 122.225 202.740 123.135 203.155 ;
        RECT 122.325 202.590 123.135 202.730 ;
        RECT 122.325 202.420 123.325 202.590 ;
        RECT 123.345 202.435 124.025 205.640 ;
        RECT 122.325 200.900 123.135 202.420 ;
        RECT 123.345 201.525 124.245 202.435 ;
        RECT 122.455 200.750 123.135 200.890 ;
        RECT 122.455 200.580 123.325 200.750 ;
        RECT 122.455 197.375 123.135 200.580 ;
        RECT 123.345 199.990 124.025 201.525 ;
        RECT 123.345 198.640 124.255 199.990 ;
        RECT 123.345 198.445 124.025 198.590 ;
        RECT 123.155 198.275 124.025 198.445 ;
        RECT 122.235 196.465 123.135 197.375 ;
        RECT 122.455 194.930 123.135 196.465 ;
        RECT 123.345 196.745 124.025 198.275 ;
        RECT 123.345 195.380 124.255 196.745 ;
        RECT 123.345 195.230 124.155 195.370 ;
        RECT 123.155 195.060 124.155 195.230 ;
        RECT 122.225 193.580 123.135 194.930 ;
        RECT 122.265 193.090 123.050 193.520 ;
        RECT 122.225 192.655 123.135 193.070 ;
        RECT 122.225 192.485 123.325 192.655 ;
        RECT 123.345 192.620 124.155 195.060 ;
        RECT 122.225 192.140 123.135 192.485 ;
        RECT 123.185 192.355 123.295 192.475 ;
        RECT 122.455 189.170 123.135 192.140 ;
        RECT 123.345 192.010 124.025 192.040 ;
        RECT 123.155 191.840 124.025 192.010 ;
        RECT 123.345 189.495 124.025 191.840 ;
        RECT 122.355 188.790 123.135 188.930 ;
        RECT 122.355 188.620 123.325 188.790 ;
        RECT 122.355 187.560 123.135 188.620 ;
        RECT 123.345 188.575 124.255 189.495 ;
        RECT 123.345 188.330 124.255 188.390 ;
        RECT 123.155 188.160 124.255 188.330 ;
        RECT 122.225 186.605 123.135 187.550 ;
        RECT 122.425 185.115 123.105 186.605 ;
        RECT 123.345 185.390 124.255 188.160 ;
        RECT 122.425 184.945 123.325 185.115 ;
        RECT 122.425 184.800 123.105 184.945 ;
        RECT 122.325 183.730 123.135 184.790 ;
        RECT 123.345 183.730 124.155 184.790 ;
        RECT 122.325 183.560 124.155 183.730 ;
        RECT 122.325 183.420 123.135 183.560 ;
        RECT 123.345 183.420 124.155 183.560 ;
      LAYER nwell ;
        RECT 124.545 183.225 127.375 219.485 ;
      LAYER pwell ;
        RECT 127.765 219.150 128.575 219.290 ;
        RECT 128.785 219.150 129.595 219.290 ;
        RECT 127.765 218.980 129.595 219.150 ;
        RECT 127.765 217.920 128.575 218.980 ;
        RECT 128.785 217.920 129.595 218.980 ;
        RECT 127.665 216.565 128.575 217.910 ;
        RECT 128.785 217.770 129.595 217.910 ;
        RECT 128.595 217.600 129.595 217.770 ;
        RECT 127.895 216.390 128.575 216.565 ;
        RECT 128.785 216.540 129.595 217.600 ;
        RECT 128.785 216.390 129.465 216.420 ;
        RECT 127.895 216.220 129.465 216.390 ;
        RECT 127.895 216.080 128.575 216.220 ;
        RECT 128.625 215.815 128.735 215.935 ;
        RECT 127.665 215.195 128.575 215.610 ;
        RECT 127.665 215.025 128.765 215.195 ;
        RECT 127.665 214.680 128.575 215.025 ;
        RECT 127.895 211.710 128.575 214.680 ;
        RECT 128.785 213.875 129.465 216.220 ;
        RECT 128.785 212.955 129.695 213.875 ;
        RECT 128.785 211.835 129.695 212.755 ;
        RECT 127.895 211.330 128.575 211.470 ;
        RECT 127.895 211.160 128.765 211.330 ;
        RECT 127.895 207.955 128.575 211.160 ;
        RECT 128.785 209.490 129.465 211.835 ;
        RECT 128.595 209.320 129.465 209.490 ;
        RECT 128.785 209.290 129.465 209.320 ;
        RECT 128.785 209.030 129.595 209.170 ;
        RECT 128.595 208.860 129.595 209.030 ;
        RECT 127.675 207.045 128.575 207.955 ;
        RECT 127.895 205.510 128.575 207.045 ;
        RECT 128.785 206.420 129.595 208.860 ;
        RECT 128.870 205.970 129.655 206.400 ;
        RECT 127.665 204.160 128.575 205.510 ;
        RECT 128.785 204.895 129.695 205.930 ;
        RECT 128.595 204.725 129.695 204.895 ;
        RECT 128.785 204.580 129.695 204.725 ;
        RECT 127.665 203.695 128.575 204.110 ;
        RECT 127.665 203.525 128.765 203.695 ;
        RECT 127.665 203.180 128.575 203.525 ;
        RECT 127.895 200.210 128.575 203.180 ;
        RECT 128.785 200.750 129.695 204.500 ;
        RECT 128.595 200.580 129.695 200.750 ;
        RECT 128.785 200.440 129.695 200.580 ;
        RECT 127.665 198.955 128.575 199.875 ;
        RECT 127.895 196.610 128.575 198.955 ;
        RECT 128.785 199.415 129.695 200.335 ;
        RECT 128.785 197.070 129.465 199.415 ;
        RECT 128.595 196.900 129.465 197.070 ;
        RECT 128.785 196.870 129.465 196.900 ;
        RECT 128.785 196.610 129.595 196.750 ;
        RECT 127.895 196.440 129.595 196.610 ;
        RECT 127.895 196.410 128.575 196.440 ;
        RECT 127.765 196.150 128.575 196.290 ;
        RECT 127.765 195.980 128.765 196.150 ;
        RECT 127.765 193.540 128.575 195.980 ;
        RECT 128.785 195.380 129.595 196.440 ;
        RECT 128.785 194.420 129.695 195.370 ;
        RECT 127.705 193.090 128.490 193.520 ;
        RECT 127.665 190.175 128.575 192.780 ;
        RECT 128.815 192.015 129.495 194.420 ;
        RECT 128.595 191.845 129.495 192.015 ;
        RECT 128.815 191.700 129.495 191.845 ;
        RECT 128.785 191.545 129.695 191.690 ;
        RECT 128.595 191.375 129.695 191.545 ;
        RECT 128.785 190.340 129.695 191.375 ;
        RECT 127.665 190.160 128.765 190.175 ;
        RECT 128.785 190.160 129.565 190.310 ;
        RECT 127.665 190.005 129.565 190.160 ;
        RECT 127.665 189.860 128.575 190.005 ;
        RECT 128.595 189.990 129.565 190.005 ;
        RECT 128.620 189.540 128.730 189.700 ;
        RECT 128.785 188.940 129.565 189.990 ;
        RECT 127.665 185.570 128.575 188.790 ;
        RECT 128.785 185.570 129.695 188.790 ;
        RECT 127.665 185.400 129.695 185.570 ;
        RECT 127.665 185.340 128.575 185.400 ;
        RECT 128.785 185.340 129.695 185.400 ;
        RECT 128.625 184.995 128.735 185.115 ;
        RECT 127.765 183.730 128.575 184.790 ;
        RECT 128.785 183.730 129.595 184.790 ;
        RECT 127.765 183.560 129.595 183.730 ;
        RECT 127.765 183.420 128.575 183.560 ;
        RECT 128.785 183.420 129.595 183.560 ;
      LAYER nwell ;
        RECT 129.985 183.225 132.815 219.485 ;
      LAYER pwell ;
        RECT 133.205 219.150 134.015 219.290 ;
        RECT 134.225 219.150 135.035 219.290 ;
        RECT 133.205 218.980 135.035 219.150 ;
        RECT 133.205 217.920 134.015 218.980 ;
        RECT 134.225 217.920 135.035 218.980 ;
        RECT 133.105 216.520 134.015 217.870 ;
        RECT 134.225 217.495 135.135 217.910 ;
        RECT 134.035 217.325 135.135 217.495 ;
        RECT 133.335 214.985 134.015 216.520 ;
        RECT 133.115 214.075 134.015 214.985 ;
        RECT 133.335 210.870 134.015 214.075 ;
        RECT 134.225 216.980 135.135 217.325 ;
        RECT 134.225 214.010 134.905 216.980 ;
        RECT 134.225 213.630 134.905 213.770 ;
        RECT 134.035 213.460 134.905 213.630 ;
        RECT 133.335 210.700 134.205 210.870 ;
        RECT 133.335 210.560 134.015 210.700 ;
        RECT 133.205 210.410 134.015 210.550 ;
        RECT 133.205 210.240 134.205 210.410 ;
        RECT 134.225 210.255 134.905 213.460 ;
        RECT 133.205 207.800 134.015 210.240 ;
        RECT 134.225 209.345 135.125 210.255 ;
        RECT 134.225 207.810 134.905 209.345 ;
        RECT 134.065 207.535 134.175 207.655 ;
        RECT 133.335 207.190 134.015 207.330 ;
        RECT 133.335 207.020 134.205 207.190 ;
        RECT 133.335 198.225 134.015 207.020 ;
        RECT 134.225 206.460 135.135 207.810 ;
        RECT 134.310 205.970 135.095 206.400 ;
        RECT 134.225 205.810 134.905 205.950 ;
        RECT 134.035 205.640 134.905 205.810 ;
        RECT 134.225 202.435 134.905 205.640 ;
        RECT 134.225 201.525 135.125 202.435 ;
        RECT 134.225 199.990 134.905 201.525 ;
        RECT 134.225 198.640 135.135 199.990 ;
        RECT 134.065 198.335 134.175 198.455 ;
        RECT 133.105 197.115 134.015 198.035 ;
        RECT 133.335 194.770 134.015 197.115 ;
        RECT 134.225 196.765 135.135 198.130 ;
        RECT 134.225 195.235 134.905 196.765 ;
        RECT 134.035 195.065 134.905 195.235 ;
        RECT 134.225 194.920 134.905 195.065 ;
        RECT 133.335 194.600 134.205 194.770 ;
        RECT 133.335 194.570 134.015 194.600 ;
        RECT 134.060 194.140 134.170 194.300 ;
        RECT 134.225 193.850 135.135 193.910 ;
        RECT 134.035 193.680 135.135 193.850 ;
        RECT 133.145 193.090 133.930 193.520 ;
        RECT 133.305 192.935 133.985 193.060 ;
        RECT 133.305 192.765 134.205 192.935 ;
        RECT 133.305 191.735 133.985 192.765 ;
        RECT 133.105 190.780 134.015 191.735 ;
        RECT 134.225 190.910 135.135 193.680 ;
        RECT 133.205 190.630 134.015 190.770 ;
        RECT 133.205 190.625 134.205 190.630 ;
        RECT 134.225 190.625 135.135 190.770 ;
        RECT 133.205 190.460 135.135 190.625 ;
        RECT 133.205 188.020 134.015 190.460 ;
        RECT 134.035 190.455 135.135 190.460 ;
        RECT 134.225 189.420 135.135 190.455 ;
        RECT 134.065 189.135 134.175 189.255 ;
        RECT 134.225 188.790 135.135 188.850 ;
        RECT 134.035 188.620 135.135 188.790 ;
        RECT 134.065 187.755 134.175 187.875 ;
        RECT 133.105 186.495 134.015 187.530 ;
        RECT 133.105 186.325 134.205 186.495 ;
        RECT 133.105 186.180 134.015 186.325 ;
        RECT 133.235 185.110 134.015 186.170 ;
        RECT 134.225 185.400 135.135 188.620 ;
        RECT 134.065 185.110 134.175 185.115 ;
        RECT 133.235 184.940 134.205 185.110 ;
        RECT 133.235 184.800 134.015 184.940 ;
        RECT 133.205 183.730 134.015 184.790 ;
        RECT 134.225 183.730 135.035 184.790 ;
        RECT 133.205 183.560 135.035 183.730 ;
        RECT 133.205 183.420 134.015 183.560 ;
        RECT 134.225 183.420 135.035 183.560 ;
      LAYER nwell ;
        RECT 135.425 183.225 138.255 219.485 ;
      LAYER pwell ;
        RECT 138.645 219.150 139.455 219.290 ;
        RECT 139.665 219.150 140.475 219.290 ;
        RECT 138.645 218.980 140.475 219.150 ;
        RECT 138.645 217.920 139.455 218.980 ;
        RECT 139.665 217.920 140.475 218.980 ;
        RECT 138.545 216.565 139.455 217.910 ;
        RECT 139.665 217.770 140.345 217.910 ;
        RECT 139.475 217.600 140.345 217.770 ;
        RECT 138.775 216.390 139.455 216.565 ;
        RECT 138.775 216.220 139.645 216.390 ;
        RECT 138.775 216.080 139.455 216.220 ;
        RECT 138.545 215.655 139.455 216.070 ;
        RECT 138.545 215.485 139.645 215.655 ;
        RECT 138.545 215.140 139.455 215.485 ;
        RECT 138.775 212.170 139.455 215.140 ;
        RECT 139.665 214.395 140.345 217.600 ;
        RECT 139.665 213.485 140.565 214.395 ;
        RECT 139.665 211.950 140.345 213.485 ;
        RECT 138.645 211.790 139.455 211.930 ;
        RECT 138.645 211.620 139.645 211.790 ;
        RECT 138.645 210.560 139.455 211.620 ;
        RECT 139.665 210.600 140.575 211.950 ;
        RECT 138.775 201.670 139.455 210.465 ;
        RECT 139.665 209.535 140.575 210.455 ;
        RECT 139.665 207.190 140.345 209.535 ;
        RECT 139.475 207.020 140.345 207.190 ;
        RECT 139.665 206.990 140.345 207.020 ;
        RECT 139.505 206.615 139.615 206.735 ;
        RECT 139.750 205.970 140.535 206.400 ;
        RECT 139.665 205.535 140.575 205.950 ;
        RECT 139.475 205.365 140.575 205.535 ;
        RECT 139.665 205.020 140.575 205.365 ;
        RECT 139.665 202.050 140.345 205.020 ;
        RECT 139.505 201.670 139.615 201.675 ;
        RECT 138.775 201.500 139.645 201.670 ;
        RECT 138.775 201.360 139.455 201.500 ;
        RECT 138.545 200.335 139.455 201.255 ;
        RECT 139.475 201.205 139.645 201.210 ;
        RECT 139.475 201.040 140.345 201.205 ;
        RECT 138.775 197.990 139.455 200.335 ;
        RECT 139.665 200.300 140.345 201.040 ;
        RECT 139.665 199.370 140.575 200.300 ;
        RECT 139.665 197.990 140.575 199.040 ;
        RECT 138.775 197.820 140.575 197.990 ;
        RECT 138.775 197.790 139.455 197.820 ;
        RECT 139.665 197.690 140.575 197.820 ;
        RECT 138.645 197.530 139.455 197.670 ;
        RECT 139.665 197.530 140.345 197.670 ;
        RECT 138.645 197.360 140.345 197.530 ;
        RECT 138.645 196.300 139.455 197.360 ;
        RECT 138.745 196.145 139.425 196.290 ;
        RECT 138.745 195.975 139.645 196.145 ;
        RECT 138.745 194.485 139.425 195.975 ;
        RECT 138.545 193.540 139.455 194.485 ;
        RECT 139.665 194.155 140.345 197.360 ;
        RECT 138.585 193.090 139.370 193.520 ;
        RECT 139.665 193.245 140.565 194.155 ;
        RECT 138.545 192.930 139.455 192.990 ;
        RECT 138.545 192.760 139.645 192.930 ;
        RECT 138.545 189.540 139.455 192.760 ;
        RECT 139.665 191.710 140.345 193.245 ;
        RECT 139.665 190.360 140.575 191.710 ;
        RECT 139.505 190.055 139.615 190.175 ;
        RECT 139.475 189.705 139.645 189.710 ;
        RECT 139.475 189.540 140.345 189.705 ;
        RECT 138.545 189.250 139.455 189.310 ;
        RECT 138.545 189.080 139.645 189.250 ;
        RECT 138.545 185.860 139.455 189.080 ;
        RECT 139.665 188.800 140.345 189.540 ;
        RECT 139.665 187.870 140.575 188.800 ;
        RECT 139.665 187.410 140.445 187.550 ;
        RECT 139.475 187.240 140.445 187.410 ;
        RECT 139.665 186.180 140.445 187.240 ;
        RECT 139.500 185.400 139.610 185.560 ;
        RECT 139.665 185.120 140.445 186.170 ;
        RECT 139.475 184.950 140.445 185.120 ;
        RECT 139.665 184.800 140.445 184.950 ;
        RECT 138.645 183.730 139.455 184.790 ;
        RECT 139.665 183.730 140.475 184.790 ;
        RECT 138.645 183.560 140.475 183.730 ;
        RECT 138.645 183.420 139.455 183.560 ;
        RECT 139.665 183.420 140.475 183.560 ;
      LAYER nwell ;
        RECT 140.865 183.225 143.695 219.485 ;
      LAYER pwell ;
        RECT 144.085 219.150 144.895 219.290 ;
        RECT 145.105 219.150 145.915 219.290 ;
        RECT 144.085 218.980 145.915 219.150 ;
        RECT 144.085 217.920 144.895 218.980 ;
        RECT 145.105 217.920 145.915 218.980 ;
        RECT 144.085 217.770 144.895 217.910 ;
        RECT 145.105 217.770 145.915 217.910 ;
        RECT 144.085 217.600 145.915 217.770 ;
        RECT 144.085 214.240 144.895 217.600 ;
        RECT 144.945 213.975 145.055 214.095 ;
        RECT 143.985 212.380 144.895 213.730 ;
        RECT 145.105 212.400 145.915 217.600 ;
        RECT 144.215 210.845 144.895 212.380 ;
        RECT 144.950 212.080 145.060 212.240 ;
        RECT 145.105 211.330 145.785 211.470 ;
        RECT 144.915 211.160 145.785 211.330 ;
        RECT 143.995 209.935 144.895 210.845 ;
        RECT 144.215 206.730 144.895 209.935 ;
        RECT 145.105 210.985 145.785 211.160 ;
        RECT 145.105 209.640 146.015 210.985 ;
        RECT 145.105 206.730 146.015 209.500 ;
        RECT 144.215 206.560 146.015 206.730 ;
        RECT 144.215 206.420 144.895 206.560 ;
        RECT 145.105 206.500 146.015 206.560 ;
        RECT 144.215 206.270 144.895 206.410 ;
        RECT 144.215 206.100 145.085 206.270 ;
        RECT 144.215 202.895 144.895 206.100 ;
        RECT 145.190 205.970 145.975 206.400 ;
        RECT 144.950 205.640 145.060 205.800 ;
        RECT 145.105 204.890 145.785 204.920 ;
        RECT 144.915 204.720 145.785 204.890 ;
        RECT 143.995 201.985 144.895 202.895 ;
        RECT 144.215 200.450 144.895 201.985 ;
        RECT 145.105 202.375 145.785 204.720 ;
        RECT 145.105 201.455 146.015 202.375 ;
        RECT 144.950 201.040 145.060 201.200 ;
        RECT 143.985 199.100 144.895 200.450 ;
        RECT 145.105 199.085 146.015 200.430 ;
        RECT 145.105 198.910 145.785 199.085 ;
        RECT 144.915 198.740 145.785 198.910 ;
        RECT 143.985 197.810 144.895 198.740 ;
        RECT 145.105 198.600 145.785 198.740 ;
        RECT 145.105 198.450 145.785 198.480 ;
        RECT 144.915 198.280 145.785 198.450 ;
        RECT 144.215 197.070 144.895 197.810 ;
        RECT 144.215 196.905 145.085 197.070 ;
        RECT 144.915 196.900 145.085 196.905 ;
        RECT 144.215 196.610 144.895 196.750 ;
        RECT 144.215 196.440 145.085 196.610 ;
        RECT 144.215 196.265 144.895 196.440 ;
        RECT 143.985 194.920 144.895 196.265 ;
        RECT 145.105 195.935 145.785 198.280 ;
        RECT 145.105 195.015 146.015 195.935 ;
        RECT 143.985 194.770 144.895 194.900 ;
        RECT 143.985 194.760 145.085 194.770 ;
        RECT 145.105 194.760 145.885 194.910 ;
        RECT 143.985 194.600 145.885 194.760 ;
        RECT 143.985 193.550 144.895 194.600 ;
        RECT 144.915 194.590 145.885 194.600 ;
        RECT 145.105 193.540 145.885 194.590 ;
        RECT 144.025 193.090 144.810 193.520 ;
        RECT 145.190 193.090 145.975 193.520 ;
        RECT 143.985 192.930 144.895 192.990 ;
        RECT 143.985 192.760 145.085 192.930 ;
        RECT 143.985 189.990 144.895 192.760 ;
        RECT 145.105 190.805 146.015 192.150 ;
        RECT 145.105 190.630 145.785 190.805 ;
        RECT 144.915 190.460 145.785 190.630 ;
        RECT 145.105 190.320 145.785 190.460 ;
        RECT 145.105 190.170 145.915 190.310 ;
        RECT 144.915 190.000 145.915 190.170 ;
        RECT 144.215 189.710 144.895 189.740 ;
        RECT 144.215 189.540 145.085 189.710 ;
        RECT 144.215 187.195 144.895 189.540 ;
        RECT 145.105 188.940 145.915 190.000 ;
        RECT 145.105 187.870 145.885 188.930 ;
        RECT 144.915 187.700 145.885 187.870 ;
        RECT 145.105 187.560 145.885 187.700 ;
        RECT 143.985 186.275 144.895 187.195 ;
        RECT 145.105 186.490 145.885 187.550 ;
        RECT 144.915 186.320 145.885 186.490 ;
        RECT 145.105 186.180 145.885 186.320 ;
        RECT 144.115 185.120 144.895 186.170 ;
        RECT 145.105 185.120 145.885 186.170 ;
        RECT 144.115 184.950 145.885 185.120 ;
        RECT 144.115 184.800 144.895 184.950 ;
        RECT 145.105 184.800 145.885 184.950 ;
        RECT 144.085 183.730 144.895 184.790 ;
        RECT 145.105 183.730 145.915 184.790 ;
        RECT 144.085 183.560 145.915 183.730 ;
        RECT 144.085 183.420 144.895 183.560 ;
        RECT 145.105 183.420 145.915 183.560 ;
      LAYER nwell ;
        RECT 146.305 183.225 147.910 219.485 ;
      LAYER pwell ;
        RECT 63.950 182.185 64.895 182.215 ;
        RECT 61.825 181.985 64.895 182.185 ;
        RECT 65.365 182.185 66.300 182.215 ;
        RECT 68.260 182.185 68.430 182.405 ;
        RECT 68.725 182.215 68.895 182.405 ;
        RECT 71.025 182.215 71.195 182.405 ;
        RECT 77.465 182.235 77.635 182.425 ;
        RECT 78.385 182.215 78.555 182.425 ;
        RECT 83.905 182.215 84.075 182.425 ;
        RECT 89.425 182.215 89.595 182.425 ;
        RECT 91.725 182.215 91.895 182.425 ;
        RECT 61.685 181.505 64.895 181.985 ;
        RECT 61.685 181.305 62.615 181.505 ;
        RECT 63.950 181.305 64.895 181.505 ;
        RECT 64.915 181.345 65.345 182.130 ;
        RECT 65.365 181.985 68.430 182.185 ;
        RECT 65.365 181.505 68.575 181.985 ;
        RECT 68.585 181.535 70.875 182.215 ;
        RECT 70.885 181.535 78.195 182.215 ;
        RECT 65.365 181.305 66.315 181.505 ;
        RECT 67.645 181.305 68.575 181.505 ;
        RECT 69.955 181.305 70.875 181.535 ;
        RECT 74.400 181.315 75.310 181.535 ;
        RECT 76.845 181.305 78.195 181.535 ;
        RECT 78.245 181.405 83.755 182.215 ;
        RECT 83.765 181.405 89.275 182.215 ;
        RECT 89.285 181.405 90.655 182.215 ;
        RECT 90.665 181.405 92.035 182.215 ;
      LAYER nwell ;
        RECT 13.190 178.185 92.230 181.015 ;
      LAYER pwell ;
        RECT 13.385 176.985 14.755 177.795 ;
        RECT 14.765 176.985 18.435 177.795 ;
        RECT 18.945 177.665 20.295 177.895 ;
        RECT 21.830 177.665 22.740 177.885 ;
        RECT 18.945 176.985 26.255 177.665 ;
        RECT 26.275 177.070 26.705 177.855 ;
        RECT 26.725 177.695 27.655 177.895 ;
        RECT 28.985 177.695 29.935 177.895 ;
        RECT 26.725 177.215 29.935 177.695 ;
        RECT 33.460 177.665 34.370 177.885 ;
        RECT 35.905 177.665 37.255 177.895 ;
        RECT 26.870 177.015 29.935 177.215 ;
        RECT 13.525 176.775 13.695 176.985 ;
        RECT 14.905 176.775 15.075 176.985 ;
        RECT 18.580 176.825 18.700 176.935 ;
        RECT 20.420 176.825 20.540 176.935 ;
        RECT 20.885 176.775 21.055 176.965 ;
        RECT 23.645 176.775 23.815 176.965 ;
        RECT 25.945 176.795 26.115 176.985 ;
        RECT 26.870 176.795 27.040 177.015 ;
        RECT 29.000 176.985 29.935 177.015 ;
        RECT 29.945 176.985 37.255 177.665 ;
        RECT 37.765 177.665 38.695 177.895 ;
        RECT 37.765 176.985 40.515 177.665 ;
        RECT 40.525 176.985 46.035 177.795 ;
        RECT 47.095 177.665 48.025 177.895 ;
        RECT 50.610 177.695 51.555 177.895 ;
        RECT 46.190 176.985 48.025 177.665 ;
        RECT 48.805 177.015 51.555 177.695 ;
        RECT 52.035 177.070 52.465 177.855 ;
        RECT 29.165 176.775 29.335 176.965 ;
        RECT 30.085 176.795 30.255 176.985 ;
        RECT 34.685 176.775 34.855 176.965 ;
        RECT 37.440 176.825 37.560 176.935 ;
        RECT 38.375 176.820 38.535 176.930 ;
        RECT 39.745 176.775 39.915 176.965 ;
        RECT 40.205 176.795 40.375 176.985 ;
        RECT 40.665 176.795 40.835 176.985 ;
        RECT 46.190 176.965 46.355 176.985 ;
        RECT 43.425 176.775 43.595 176.965 ;
        RECT 44.810 176.775 44.980 176.965 ;
        RECT 46.185 176.775 46.355 176.965 ;
        RECT 48.480 176.825 48.600 176.935 ;
        RECT 48.950 176.795 49.120 177.015 ;
        RECT 50.610 176.985 51.555 177.015 ;
        RECT 52.485 176.985 55.695 177.895 ;
        RECT 56.165 176.985 57.515 177.895 ;
        RECT 57.545 177.665 58.465 177.895 ;
        RECT 57.545 176.985 59.835 177.665 ;
        RECT 59.905 176.985 61.675 177.895 ;
        RECT 62.605 176.985 66.080 177.895 ;
        RECT 66.285 176.985 69.955 177.795 ;
        RECT 69.985 176.985 71.335 177.895 ;
        RECT 71.345 176.985 72.695 177.895 ;
        RECT 72.725 176.985 76.395 177.795 ;
        RECT 76.405 176.985 77.775 177.795 ;
        RECT 77.795 177.070 78.225 177.855 ;
        RECT 78.245 176.985 83.755 177.795 ;
        RECT 83.765 176.985 89.275 177.795 ;
        RECT 89.285 176.985 90.655 177.795 ;
        RECT 90.665 176.985 92.035 177.795 ;
        RECT 51.705 176.935 51.875 176.965 ;
        RECT 51.700 176.825 51.875 176.935 ;
        RECT 51.705 176.775 51.875 176.825 ;
        RECT 52.625 176.795 52.795 176.985 ;
        RECT 57.230 176.965 57.400 176.985 ;
        RECT 55.840 176.825 55.960 176.935 ;
        RECT 57.225 176.795 57.400 176.965 ;
        RECT 59.525 176.795 59.695 176.985 ;
        RECT 61.360 176.795 61.530 176.985 ;
        RECT 62.750 176.965 62.920 176.985 ;
        RECT 61.835 176.830 61.995 176.940 ;
        RECT 62.745 176.795 62.920 176.965 ;
        RECT 64.580 176.825 64.700 176.935 ;
        RECT 57.225 176.775 57.395 176.795 ;
        RECT 62.745 176.775 62.915 176.795 ;
        RECT 65.505 176.775 65.675 176.965 ;
        RECT 66.425 176.795 66.595 176.985 ;
        RECT 69.185 176.775 69.355 176.965 ;
        RECT 69.655 176.820 69.815 176.930 ;
        RECT 70.570 176.775 70.740 176.965 ;
        RECT 71.020 176.795 71.190 176.985 ;
        RECT 71.490 176.795 71.660 176.985 ;
        RECT 72.865 176.965 73.035 176.985 ;
        RECT 72.860 176.795 73.035 176.965 ;
        RECT 72.860 176.775 73.030 176.795 ;
        RECT 74.250 176.775 74.420 176.965 ;
        RECT 74.705 176.775 74.875 176.965 ;
        RECT 76.545 176.795 76.715 176.985 ;
        RECT 78.385 176.795 78.555 176.985 ;
        RECT 80.225 176.775 80.395 176.965 ;
        RECT 83.905 176.795 84.075 176.985 ;
        RECT 85.745 176.775 85.915 176.965 ;
        RECT 89.425 176.775 89.595 176.985 ;
        RECT 91.725 176.775 91.895 176.985 ;
        RECT 13.385 175.965 14.755 176.775 ;
        RECT 14.765 175.965 20.275 176.775 ;
        RECT 20.745 176.095 23.495 176.775 ;
        RECT 22.565 175.865 23.495 176.095 ;
        RECT 23.505 175.965 29.015 176.775 ;
        RECT 29.025 175.965 34.535 176.775 ;
        RECT 34.545 175.965 38.215 176.775 ;
        RECT 39.155 175.905 39.585 176.690 ;
        RECT 39.605 175.965 43.275 176.775 ;
        RECT 43.285 175.965 44.655 176.775 ;
        RECT 44.665 175.865 46.015 176.775 ;
        RECT 46.045 175.965 51.555 176.775 ;
        RECT 51.565 175.965 57.075 176.775 ;
        RECT 57.085 175.965 62.595 176.775 ;
        RECT 62.605 175.965 64.435 176.775 ;
        RECT 64.915 175.905 65.345 176.690 ;
        RECT 65.365 175.965 68.115 176.775 ;
        RECT 68.135 175.865 69.485 176.775 ;
        RECT 70.425 175.865 71.775 176.775 ;
        RECT 71.825 175.865 73.175 176.775 ;
        RECT 73.185 175.865 74.535 176.775 ;
        RECT 74.565 175.965 80.075 176.775 ;
        RECT 80.085 175.965 85.595 176.775 ;
        RECT 85.605 175.965 89.275 176.775 ;
        RECT 89.285 175.965 90.655 176.775 ;
        RECT 90.665 175.965 92.035 176.775 ;
      LAYER nwell ;
        RECT 13.190 172.745 92.230 175.575 ;
      LAYER pwell ;
        RECT 13.385 171.545 14.755 172.355 ;
        RECT 14.765 171.545 20.275 172.355 ;
        RECT 20.285 171.545 25.795 172.355 ;
        RECT 26.275 171.630 26.705 172.415 ;
        RECT 26.725 171.545 29.475 172.355 ;
        RECT 31.315 172.225 32.235 172.455 ;
        RECT 29.945 171.545 32.235 172.225 ;
        RECT 32.245 172.225 33.165 172.455 ;
        RECT 32.245 171.545 34.535 172.225 ;
        RECT 34.545 171.545 37.295 172.355 ;
        RECT 42.825 172.225 43.745 172.455 ;
        RECT 45.125 172.225 46.045 172.455 ;
        RECT 38.000 171.545 42.815 172.225 ;
        RECT 42.825 171.545 45.115 172.225 ;
        RECT 45.125 171.545 47.415 172.225 ;
        RECT 47.425 171.545 49.240 172.455 ;
        RECT 49.265 171.545 52.015 172.355 ;
        RECT 52.035 171.630 52.465 172.415 ;
        RECT 52.485 171.545 54.315 172.225 ;
        RECT 54.325 171.545 56.155 172.225 ;
        RECT 56.165 171.545 57.535 172.355 ;
        RECT 57.565 171.545 58.915 172.455 ;
        RECT 58.925 171.545 62.135 172.455 ;
        RECT 62.600 171.775 64.435 172.455 ;
        RECT 62.600 171.545 64.290 171.775 ;
        RECT 64.445 171.545 66.275 172.355 ;
        RECT 66.745 172.225 67.880 172.455 ;
        RECT 70.165 172.365 71.115 172.455 ;
        RECT 66.745 171.545 69.955 172.225 ;
        RECT 70.165 171.545 72.095 172.365 ;
        RECT 74.340 172.225 75.475 172.455 ;
        RECT 72.265 171.545 75.475 172.225 ;
        RECT 75.795 172.225 76.725 172.455 ;
        RECT 75.795 171.545 77.630 172.225 ;
        RECT 77.795 171.630 78.225 172.415 ;
        RECT 81.760 172.225 82.670 172.445 ;
        RECT 84.205 172.225 85.555 172.455 ;
        RECT 78.245 171.545 85.555 172.225 ;
        RECT 85.605 171.545 89.275 172.355 ;
        RECT 89.285 171.545 90.655 172.355 ;
        RECT 90.665 171.545 92.035 172.355 ;
        RECT 13.525 171.335 13.695 171.545 ;
        RECT 14.905 171.335 15.075 171.545 ;
        RECT 20.425 171.335 20.595 171.545 ;
        RECT 22.265 171.335 22.435 171.525 ;
        RECT 25.940 171.385 26.060 171.495 ;
        RECT 26.865 171.355 27.035 171.545 ;
        RECT 29.620 171.335 29.790 171.525 ;
        RECT 30.085 171.355 30.255 171.545 ;
        RECT 31.005 171.335 31.175 171.525 ;
        RECT 34.225 171.355 34.395 171.545 ;
        RECT 34.685 171.355 34.855 171.545 ;
        RECT 37.440 171.385 37.560 171.495 ;
        RECT 38.375 171.380 38.535 171.490 ;
        RECT 39.745 171.335 39.915 171.525 ;
        RECT 42.505 171.355 42.675 171.545 ;
        RECT 44.805 171.355 44.975 171.545 ;
        RECT 47.105 171.355 47.275 171.545 ;
        RECT 48.945 171.355 49.115 171.545 ;
        RECT 49.405 171.355 49.575 171.545 ;
        RECT 49.865 171.335 50.035 171.525 ;
        RECT 52.625 171.355 52.795 171.545 ;
        RECT 55.845 171.355 56.015 171.545 ;
        RECT 56.305 171.355 56.475 171.545 ;
        RECT 58.600 171.355 58.770 171.545 ;
        RECT 59.065 171.335 59.235 171.525 ;
        RECT 59.535 171.380 59.695 171.490 ;
        RECT 61.825 171.335 61.995 171.545 ;
        RECT 62.285 171.335 62.455 171.525 ;
        RECT 64.120 171.355 64.290 171.545 ;
        RECT 64.585 171.355 64.755 171.545 ;
        RECT 65.510 171.335 65.680 171.525 ;
        RECT 66.420 171.385 66.540 171.495 ;
        RECT 69.185 171.335 69.355 171.525 ;
        RECT 69.645 171.355 69.815 171.545 ;
        RECT 71.945 171.525 72.095 171.545 ;
        RECT 71.945 171.355 72.115 171.525 ;
        RECT 72.405 171.355 72.575 171.545 ;
        RECT 77.465 171.525 77.630 171.545 ;
        RECT 77.465 171.355 77.635 171.525 ;
        RECT 77.925 171.335 78.095 171.525 ;
        RECT 78.385 171.335 78.555 171.545 ;
        RECT 83.905 171.335 84.075 171.525 ;
        RECT 85.745 171.355 85.915 171.545 ;
        RECT 89.425 171.335 89.595 171.545 ;
        RECT 91.725 171.335 91.895 171.545 ;
        RECT 13.385 170.525 14.755 171.335 ;
        RECT 14.765 170.525 20.275 171.335 ;
        RECT 20.285 170.525 22.115 171.335 ;
        RECT 22.125 170.655 29.435 171.335 ;
        RECT 25.640 170.435 26.550 170.655 ;
        RECT 28.085 170.425 29.435 170.655 ;
        RECT 29.505 170.425 30.855 171.335 ;
        RECT 30.865 170.655 38.175 171.335 ;
        RECT 34.380 170.435 35.290 170.655 ;
        RECT 36.825 170.425 38.175 170.655 ;
        RECT 39.155 170.465 39.585 171.250 ;
        RECT 39.660 170.425 49.680 171.335 ;
        RECT 49.725 170.655 57.035 171.335 ;
        RECT 53.240 170.435 54.150 170.655 ;
        RECT 55.685 170.425 57.035 170.655 ;
        RECT 57.085 170.425 59.375 171.335 ;
        RECT 60.305 170.655 62.135 171.335 ;
        RECT 60.305 170.425 61.650 170.655 ;
        RECT 62.145 170.525 64.895 171.335 ;
        RECT 64.915 170.465 65.345 171.250 ;
        RECT 65.365 170.655 69.035 171.335 ;
        RECT 65.365 170.425 66.290 170.655 ;
        RECT 69.045 170.525 70.875 171.335 ;
        RECT 70.925 170.655 78.235 171.335 ;
        RECT 70.925 170.425 72.275 170.655 ;
        RECT 73.810 170.435 74.720 170.655 ;
        RECT 78.245 170.525 83.755 171.335 ;
        RECT 83.765 170.525 89.275 171.335 ;
        RECT 89.285 170.525 90.655 171.335 ;
        RECT 90.665 170.525 92.035 171.335 ;
      LAYER nwell ;
        RECT 13.190 167.305 92.230 170.135 ;
      LAYER pwell ;
        RECT 100.450 167.190 106.550 176.980 ;
        RECT 100.450 167.160 106.560 167.190 ;
        RECT 13.385 166.105 14.755 166.915 ;
        RECT 14.765 166.105 20.275 166.915 ;
        RECT 20.285 166.105 22.115 166.915 ;
        RECT 22.585 166.815 23.535 167.015 ;
        RECT 24.865 166.815 25.795 167.015 ;
        RECT 22.585 166.335 25.795 166.815 ;
        RECT 22.585 166.135 25.650 166.335 ;
        RECT 26.275 166.190 26.705 166.975 ;
        RECT 22.585 166.105 23.520 166.135 ;
        RECT 13.525 165.895 13.695 166.105 ;
        RECT 14.905 165.895 15.075 166.105 ;
        RECT 20.425 165.895 20.595 166.105 ;
        RECT 22.260 165.945 22.380 166.055 ;
        RECT 24.105 165.915 24.275 166.085 ;
        RECT 25.480 165.915 25.650 166.135 ;
        RECT 26.735 166.105 29.465 167.015 ;
        RECT 29.650 166.105 33.520 167.015 ;
        RECT 33.625 166.105 35.455 166.915 ;
        RECT 36.515 166.785 37.445 167.015 ;
        RECT 35.610 166.105 37.445 166.785 ;
        RECT 37.815 166.105 40.975 167.015 ;
        RECT 44.500 166.785 45.410 167.005 ;
        RECT 46.945 166.785 48.295 167.015 ;
        RECT 40.985 166.105 48.295 166.785 ;
        RECT 48.540 166.105 52.015 167.015 ;
        RECT 52.035 166.190 52.465 166.975 ;
        RECT 52.505 166.105 53.855 167.015 ;
        RECT 53.875 166.105 55.225 167.015 ;
        RECT 57.065 166.785 57.995 167.015 ;
        RECT 55.245 166.105 57.995 166.785 ;
        RECT 58.005 166.105 62.820 166.785 ;
        RECT 63.105 166.105 66.275 167.015 ;
        RECT 66.285 166.105 68.115 166.915 ;
        RECT 68.635 166.105 71.795 167.015 ;
        RECT 71.805 166.785 72.725 167.015 ;
        RECT 71.805 166.105 74.095 166.785 ;
        RECT 74.105 166.105 77.775 166.915 ;
        RECT 77.795 166.190 78.225 166.975 ;
        RECT 78.245 166.105 83.755 166.915 ;
        RECT 83.765 166.105 89.275 166.915 ;
        RECT 89.285 166.105 90.655 166.915 ;
        RECT 90.665 166.105 92.035 166.915 ;
        RECT 100.650 166.760 101.810 167.160 ;
        RECT 25.940 165.945 26.060 166.055 ;
        RECT 26.865 165.915 27.035 166.105 ;
        RECT 29.650 166.085 29.795 166.105 ;
        RECT 24.110 165.895 24.275 165.915 ;
        RECT 29.165 165.895 29.335 166.085 ;
        RECT 29.625 165.915 29.795 166.085 ;
        RECT 33.765 165.915 33.935 166.105 ;
        RECT 35.610 166.085 35.775 166.105 ;
        RECT 34.225 165.895 34.395 166.085 ;
        RECT 34.685 165.895 34.855 166.085 ;
        RECT 35.605 165.915 35.775 166.085 ;
        RECT 37.445 165.895 37.615 166.085 ;
        RECT 37.905 165.915 38.075 166.105 ;
        RECT 39.745 165.895 39.915 166.085 ;
        RECT 41.125 165.915 41.295 166.105 ;
        RECT 45.265 165.895 45.435 166.085 ;
        RECT 50.785 165.895 50.955 166.085 ;
        RECT 51.700 165.915 51.870 166.105 ;
        RECT 52.620 165.915 52.790 166.105 ;
        RECT 54.005 165.915 54.175 166.105 ;
        RECT 55.385 165.915 55.555 166.105 ;
        RECT 56.305 165.895 56.475 166.085 ;
        RECT 58.145 165.915 58.315 166.105 ;
        RECT 62.280 165.945 62.400 166.055 ;
        RECT 58.170 165.895 58.315 165.915 ;
        RECT 62.750 165.895 62.920 166.085 ;
        RECT 63.205 165.915 63.375 166.105 ;
        RECT 65.505 165.895 65.675 166.085 ;
        RECT 66.425 165.915 66.595 166.105 ;
        RECT 68.260 165.945 68.380 166.055 ;
        RECT 68.725 165.895 68.895 166.105 ;
        RECT 73.785 165.895 73.955 166.105 ;
        RECT 74.245 165.915 74.415 166.105 ;
        RECT 78.385 165.915 78.555 166.105 ;
        RECT 79.305 165.895 79.475 166.085 ;
        RECT 83.905 165.915 84.075 166.105 ;
        RECT 84.825 165.895 84.995 166.085 ;
        RECT 89.425 165.915 89.595 166.105 ;
        RECT 90.340 165.945 90.460 166.055 ;
        RECT 91.725 165.895 91.895 166.105 ;
        RECT 13.385 165.085 14.755 165.895 ;
        RECT 14.765 165.085 20.275 165.895 ;
        RECT 20.285 165.085 23.955 165.895 ;
        RECT 24.110 165.215 25.945 165.895 ;
        RECT 25.015 164.985 25.945 165.215 ;
        RECT 26.265 165.215 29.475 165.895 ;
        RECT 29.720 165.215 34.535 165.895 ;
        RECT 26.265 164.985 27.400 165.215 ;
        RECT 34.555 164.985 37.285 165.895 ;
        RECT 37.305 165.085 39.135 165.895 ;
        RECT 39.155 165.025 39.585 165.810 ;
        RECT 39.605 165.085 45.115 165.895 ;
        RECT 45.125 165.085 50.635 165.895 ;
        RECT 50.645 165.085 56.155 165.895 ;
        RECT 56.165 165.085 57.995 165.895 ;
        RECT 58.170 164.985 62.040 165.895 ;
        RECT 62.750 165.665 64.440 165.895 ;
        RECT 62.605 164.985 64.440 165.665 ;
        RECT 64.915 165.025 65.345 165.810 ;
        RECT 65.365 165.215 68.105 165.895 ;
        RECT 68.585 165.215 73.400 165.895 ;
        RECT 73.645 165.085 79.155 165.895 ;
        RECT 79.165 165.085 84.675 165.895 ;
        RECT 84.685 165.085 90.195 165.895 ;
        RECT 90.665 165.085 92.035 165.895 ;
        RECT 103.770 165.080 106.560 167.160 ;
      LAYER nwell ;
        RECT 13.190 161.865 92.230 164.695 ;
        RECT 101.660 162.970 106.500 165.080 ;
        RECT 107.780 164.740 117.970 176.990 ;
      LAYER pwell ;
        RECT 120.330 167.140 126.430 176.930 ;
        RECT 120.330 167.110 126.440 167.140 ;
        RECT 120.530 166.710 121.690 167.110 ;
        RECT 123.650 165.030 126.440 167.110 ;
      LAYER nwell ;
        RECT 121.540 162.920 126.380 165.030 ;
        RECT 127.660 164.690 137.850 176.940 ;
      LAYER pwell ;
        RECT 140.360 167.190 146.460 176.980 ;
        RECT 140.360 167.160 146.470 167.190 ;
        RECT 140.560 166.760 141.720 167.160 ;
        RECT 143.680 165.080 146.470 167.160 ;
      LAYER nwell ;
        RECT 141.570 162.970 146.410 165.080 ;
        RECT 147.690 164.740 157.880 176.990 ;
      LAYER pwell ;
        RECT 13.385 160.665 14.755 161.475 ;
        RECT 14.765 160.665 20.275 161.475 ;
        RECT 20.285 160.665 25.795 161.475 ;
        RECT 26.275 160.750 26.705 161.535 ;
        RECT 26.725 161.375 27.655 161.575 ;
        RECT 28.985 161.375 29.935 161.575 ;
        RECT 26.725 160.895 29.935 161.375 ;
        RECT 30.995 161.345 31.925 161.575 ;
        RECT 26.870 160.695 29.935 160.895 ;
        RECT 13.525 160.455 13.695 160.665 ;
        RECT 14.905 160.455 15.075 160.665 ;
        RECT 20.425 160.455 20.595 160.665 ;
        RECT 24.100 160.505 24.220 160.615 ;
        RECT 25.940 160.505 26.060 160.615 ;
        RECT 26.870 160.475 27.040 160.695 ;
        RECT 29.000 160.665 29.935 160.695 ;
        RECT 30.090 160.665 31.925 161.345 ;
        RECT 32.855 160.665 36.510 161.575 ;
        RECT 36.845 160.665 39.595 161.575 ;
        RECT 40.525 160.665 43.635 161.575 ;
        RECT 43.745 160.665 46.495 161.475 ;
        RECT 46.965 160.665 48.795 161.345 ;
        RECT 48.805 160.665 51.725 161.575 ;
        RECT 52.035 160.750 52.465 161.535 ;
        RECT 52.485 160.665 53.855 161.475 ;
        RECT 54.175 161.345 55.105 161.575 ;
        RECT 56.650 161.345 57.995 161.575 ;
        RECT 54.175 160.665 56.010 161.345 ;
        RECT 56.165 160.665 57.995 161.345 ;
        RECT 58.945 160.665 60.295 161.575 ;
        RECT 60.305 160.665 63.515 161.575 ;
        RECT 63.980 160.895 65.815 161.575 ;
        RECT 63.980 160.665 65.670 160.895 ;
        RECT 65.825 160.665 67.655 161.475 ;
        RECT 67.705 160.665 70.875 161.575 ;
        RECT 73.625 161.345 74.555 161.575 ;
        RECT 70.885 160.665 74.555 161.345 ;
        RECT 74.565 160.665 77.315 161.475 ;
        RECT 77.795 160.750 78.225 161.535 ;
        RECT 78.245 160.665 83.755 161.475 ;
        RECT 83.765 160.665 89.275 161.475 ;
        RECT 89.285 160.665 90.655 161.475 ;
        RECT 90.665 160.665 92.035 161.475 ;
        RECT 30.090 160.645 30.255 160.665 ;
        RECT 32.855 160.645 33.015 160.665 ;
        RECT 30.085 160.475 30.255 160.645 ;
        RECT 31.465 160.455 31.635 160.645 ;
        RECT 31.935 160.500 32.095 160.610 ;
        RECT 32.380 160.505 32.500 160.615 ;
        RECT 32.845 160.455 33.015 160.645 ;
        RECT 35.605 160.455 35.775 160.645 ;
        RECT 36.985 160.475 37.155 160.665 ;
        RECT 37.440 160.505 37.560 160.615 ;
        RECT 37.900 160.455 38.070 160.645 ;
        RECT 39.755 160.615 39.915 160.620 ;
        RECT 39.740 160.510 39.915 160.615 ;
        RECT 39.740 160.505 39.860 160.510 ;
        RECT 40.205 160.455 40.375 160.645 ;
        RECT 43.425 160.475 43.595 160.665 ;
        RECT 43.885 160.475 44.055 160.665 ;
        RECT 46.640 160.505 46.760 160.615 ;
        RECT 47.565 160.455 47.735 160.645 ;
        RECT 48.485 160.475 48.655 160.665 ;
        RECT 48.950 160.475 49.120 160.665 ;
        RECT 52.625 160.475 52.795 160.665 ;
        RECT 55.845 160.645 56.010 160.665 ;
        RECT 54.925 160.455 55.095 160.645 ;
        RECT 55.845 160.475 56.015 160.645 ;
        RECT 56.305 160.455 56.475 160.665 ;
        RECT 58.155 160.510 58.315 160.620 ;
        RECT 59.065 160.455 59.235 160.645 ;
        RECT 59.980 160.475 60.150 160.665 ;
        RECT 60.445 160.475 60.615 160.665 ;
        RECT 65.500 160.645 65.670 160.665 ;
        RECT 64.580 160.505 64.700 160.615 ;
        RECT 65.500 160.475 65.675 160.645 ;
        RECT 65.965 160.475 66.135 160.665 ;
        RECT 67.805 160.475 67.975 160.665 ;
        RECT 65.505 160.455 65.675 160.475 ;
        RECT 71.025 160.455 71.195 160.665 ;
        RECT 72.860 160.505 72.980 160.615 ;
        RECT 73.325 160.455 73.495 160.645 ;
        RECT 74.705 160.475 74.875 160.665 ;
        RECT 77.460 160.505 77.580 160.615 ;
        RECT 78.385 160.475 78.555 160.665 ;
        RECT 80.685 160.455 80.855 160.645 ;
        RECT 83.905 160.475 84.075 160.665 ;
        RECT 86.205 160.455 86.375 160.645 ;
        RECT 89.425 160.475 89.595 160.665 ;
        RECT 89.895 160.500 90.055 160.610 ;
        RECT 91.725 160.455 91.895 160.665 ;
        RECT 13.385 159.645 14.755 160.455 ;
        RECT 14.765 159.645 20.275 160.455 ;
        RECT 20.285 159.645 23.955 160.455 ;
        RECT 24.465 159.775 31.775 160.455 ;
        RECT 24.465 159.545 25.815 159.775 ;
        RECT 27.350 159.555 28.260 159.775 ;
        RECT 32.705 159.545 35.455 160.455 ;
        RECT 35.465 159.645 37.295 160.455 ;
        RECT 37.785 159.545 39.135 160.455 ;
        RECT 39.155 159.585 39.585 160.370 ;
        RECT 40.065 159.775 47.375 160.455 ;
        RECT 47.425 159.775 54.735 160.455 ;
        RECT 43.580 159.555 44.490 159.775 ;
        RECT 46.025 159.545 47.375 159.775 ;
        RECT 50.940 159.555 51.850 159.775 ;
        RECT 53.385 159.545 54.735 159.775 ;
        RECT 54.785 159.645 56.155 160.455 ;
        RECT 56.165 159.545 58.915 160.455 ;
        RECT 58.925 159.645 64.435 160.455 ;
        RECT 64.915 159.585 65.345 160.370 ;
        RECT 65.365 159.645 70.875 160.455 ;
        RECT 70.885 159.645 72.715 160.455 ;
        RECT 73.185 159.775 80.495 160.455 ;
        RECT 76.700 159.555 77.610 159.775 ;
        RECT 79.145 159.545 80.495 159.775 ;
        RECT 80.545 159.645 86.055 160.455 ;
        RECT 86.065 159.645 89.735 160.455 ;
        RECT 90.665 159.645 92.035 160.455 ;
      LAYER nwell ;
        RECT 13.190 156.425 92.230 159.255 ;
      LAYER pwell ;
        RECT 13.385 155.225 14.755 156.035 ;
        RECT 14.765 155.225 20.275 156.035 ;
        RECT 20.285 155.225 25.795 156.035 ;
        RECT 26.275 155.310 26.705 156.095 ;
        RECT 26.725 155.225 28.075 156.135 ;
        RECT 33.365 156.045 34.315 156.135 ;
        RECT 28.105 155.225 31.775 156.035 ;
        RECT 31.785 155.225 33.155 156.035 ;
        RECT 33.365 155.225 35.295 156.045 ;
        RECT 35.465 155.225 39.135 156.035 ;
        RECT 39.145 155.225 40.515 156.035 ;
        RECT 40.525 155.905 41.455 156.135 ;
        RECT 40.525 155.225 44.195 155.905 ;
        RECT 44.205 155.225 45.575 156.035 ;
        RECT 48.325 155.905 49.255 156.135 ;
        RECT 45.585 155.225 49.255 155.905 ;
        RECT 49.265 155.225 52.015 156.035 ;
        RECT 52.035 155.310 52.465 156.095 ;
        RECT 52.485 155.225 54.315 156.035 ;
        RECT 54.325 155.905 55.250 156.135 ;
        RECT 58.005 155.935 58.955 156.135 ;
        RECT 54.325 155.225 57.995 155.905 ;
        RECT 58.005 155.255 61.675 155.935 ;
        RECT 58.005 155.225 58.955 155.255 ;
        RECT 13.525 155.015 13.695 155.225 ;
        RECT 14.905 155.015 15.075 155.225 ;
        RECT 20.425 155.015 20.595 155.225 ;
        RECT 22.260 155.065 22.380 155.175 ;
        RECT 22.725 155.015 22.895 155.205 ;
        RECT 25.940 155.065 26.060 155.175 ;
        RECT 26.865 155.035 27.035 155.205 ;
        RECT 26.865 155.015 27.030 155.035 ;
        RECT 27.325 155.015 27.495 155.205 ;
        RECT 27.790 155.035 27.960 155.225 ;
        RECT 28.245 155.035 28.415 155.225 ;
        RECT 31.925 155.035 32.095 155.225 ;
        RECT 35.145 155.205 35.295 155.225 ;
        RECT 34.685 155.015 34.855 155.205 ;
        RECT 35.145 155.035 35.315 155.205 ;
        RECT 35.605 155.035 35.775 155.225 ;
        RECT 38.375 155.060 38.535 155.170 ;
        RECT 39.285 155.035 39.455 155.225 ;
        RECT 39.745 155.015 39.915 155.205 ;
        RECT 43.885 155.035 44.055 155.225 ;
        RECT 44.345 155.035 44.515 155.225 ;
        RECT 45.265 155.015 45.435 155.205 ;
        RECT 45.725 155.035 45.895 155.225 ;
        RECT 48.945 155.015 49.115 155.205 ;
        RECT 49.405 155.035 49.575 155.225 ;
        RECT 50.330 155.015 50.500 155.205 ;
        RECT 51.705 155.015 51.875 155.205 ;
        RECT 52.625 155.035 52.795 155.225 ;
        RECT 54.470 155.035 54.640 155.225 ;
        RECT 13.385 154.205 14.755 155.015 ;
        RECT 14.765 154.205 20.275 155.015 ;
        RECT 20.285 154.205 22.115 155.015 ;
        RECT 22.585 154.335 24.875 155.015 ;
        RECT 23.955 154.105 24.875 154.335 ;
        RECT 25.195 154.335 27.030 155.015 ;
        RECT 27.185 154.335 34.495 155.015 ;
        RECT 25.195 154.105 26.125 154.335 ;
        RECT 30.700 154.115 31.610 154.335 ;
        RECT 33.145 154.105 34.495 154.335 ;
        RECT 34.545 154.205 38.215 155.015 ;
        RECT 39.155 154.145 39.585 154.930 ;
        RECT 39.605 154.205 45.115 155.015 ;
        RECT 45.125 154.205 48.795 155.015 ;
        RECT 48.805 154.205 50.175 155.015 ;
        RECT 50.185 154.105 51.535 155.015 ;
        RECT 51.645 154.105 54.645 155.015 ;
        RECT 54.930 154.985 55.100 155.205 ;
        RECT 57.685 155.015 57.855 155.205 ;
        RECT 61.360 155.170 61.530 155.255 ;
        RECT 61.685 155.225 64.895 156.135 ;
        RECT 64.905 155.225 68.015 156.135 ;
        RECT 68.125 155.225 71.235 156.135 ;
        RECT 71.825 155.225 73.175 156.135 ;
        RECT 75.925 155.905 76.855 156.135 ;
        RECT 73.185 155.225 76.855 155.905 ;
        RECT 77.795 155.310 78.225 156.095 ;
        RECT 81.760 155.905 82.670 156.125 ;
        RECT 84.205 155.905 85.555 156.135 ;
        RECT 78.245 155.225 85.555 155.905 ;
        RECT 85.605 155.225 89.275 156.035 ;
        RECT 89.285 155.225 90.655 156.035 ;
        RECT 90.665 155.225 92.035 156.035 ;
        RECT 61.360 155.060 61.535 155.170 ;
        RECT 61.360 155.035 61.530 155.060 ;
        RECT 61.815 155.035 61.985 155.225 ;
        RECT 56.590 154.985 57.535 155.015 ;
        RECT 54.785 154.305 57.535 154.985 ;
        RECT 56.590 154.105 57.535 154.305 ;
        RECT 57.545 154.205 61.215 155.015 ;
        RECT 62.145 154.985 63.100 155.015 ;
        RECT 64.130 154.985 64.300 155.205 ;
        RECT 64.580 155.065 64.700 155.175 ;
        RECT 65.515 155.060 65.675 155.170 ;
        RECT 67.805 155.035 67.975 155.225 ;
        RECT 66.285 154.985 67.240 155.015 ;
        RECT 68.270 154.985 68.440 155.205 ;
        RECT 68.735 155.060 68.895 155.170 ;
        RECT 71.025 155.035 71.195 155.225 ;
        RECT 72.860 155.205 73.030 155.225 ;
        RECT 71.480 155.065 71.600 155.175 ;
        RECT 72.405 155.015 72.575 155.205 ;
        RECT 72.860 155.035 73.035 155.205 ;
        RECT 73.325 155.035 73.495 155.225 ;
        RECT 72.865 155.015 73.035 155.035 ;
        RECT 76.545 155.015 76.715 155.205 ;
        RECT 77.015 155.070 77.175 155.180 ;
        RECT 78.385 155.015 78.555 155.225 ;
        RECT 78.845 155.015 79.015 155.205 ;
        RECT 84.365 155.015 84.535 155.205 ;
        RECT 85.745 155.035 85.915 155.225 ;
        RECT 89.425 155.035 89.595 155.225 ;
        RECT 89.895 155.060 90.055 155.170 ;
        RECT 91.725 155.015 91.895 155.225 ;
        RECT 62.145 154.305 64.425 154.985 ;
        RECT 62.145 154.105 63.100 154.305 ;
        RECT 64.915 154.145 65.345 154.930 ;
        RECT 66.285 154.305 68.565 154.985 ;
        RECT 69.505 154.335 72.715 155.015 ;
        RECT 66.285 154.105 67.240 154.305 ;
        RECT 69.505 154.105 70.640 154.335 ;
        RECT 72.725 154.205 74.555 155.015 ;
        RECT 74.565 154.335 76.855 155.015 ;
        RECT 74.565 154.105 75.485 154.335 ;
        RECT 76.865 154.105 78.680 155.015 ;
        RECT 78.705 154.205 84.215 155.015 ;
        RECT 84.225 154.205 89.735 155.015 ;
        RECT 90.665 154.205 92.035 155.015 ;
      LAYER nwell ;
        RECT 13.190 150.985 92.230 153.815 ;
      LAYER pwell ;
        RECT 100.450 152.190 106.550 161.980 ;
        RECT 100.450 152.160 106.560 152.190 ;
        RECT 100.650 151.760 101.810 152.160 ;
        RECT 13.385 149.785 14.755 150.595 ;
        RECT 14.765 149.785 18.435 150.595 ;
        RECT 22.420 150.465 23.330 150.685 ;
        RECT 24.865 150.465 26.215 150.695 ;
        RECT 18.905 149.785 26.215 150.465 ;
        RECT 26.275 149.870 26.705 150.655 ;
        RECT 26.735 149.785 29.465 150.695 ;
        RECT 29.485 149.785 32.235 150.595 ;
        RECT 32.245 149.785 35.900 150.695 ;
        RECT 35.925 149.785 37.295 150.595 ;
        RECT 37.760 150.015 39.595 150.695 ;
        RECT 37.760 149.785 39.450 150.015 ;
        RECT 40.105 149.785 43.275 150.695 ;
        RECT 43.285 149.785 44.655 150.595 ;
        RECT 44.765 149.785 47.875 150.695 ;
        RECT 47.885 149.785 49.255 150.595 ;
        RECT 51.070 150.495 52.015 150.695 ;
        RECT 49.265 149.815 52.015 150.495 ;
        RECT 52.035 149.870 52.465 150.655 ;
        RECT 13.525 149.575 13.695 149.785 ;
        RECT 14.905 149.575 15.075 149.785 ;
        RECT 18.580 149.625 18.700 149.735 ;
        RECT 19.045 149.595 19.215 149.785 ;
        RECT 13.385 148.765 14.755 149.575 ;
        RECT 14.765 148.765 20.275 149.575 ;
        RECT 20.285 149.545 21.220 149.575 ;
        RECT 23.180 149.545 23.350 149.765 ;
        RECT 23.640 149.625 23.760 149.735 ;
        RECT 25.945 149.575 26.115 149.765 ;
        RECT 26.405 149.575 26.575 149.765 ;
        RECT 26.865 149.595 27.035 149.785 ;
        RECT 29.625 149.595 29.795 149.785 ;
        RECT 31.930 149.575 32.100 149.765 ;
        RECT 32.390 149.595 32.560 149.785 ;
        RECT 35.145 149.575 35.315 149.765 ;
        RECT 36.065 149.595 36.235 149.785 ;
        RECT 38.820 149.625 38.940 149.735 ;
        RECT 39.280 149.595 39.450 149.785 ;
        RECT 39.740 149.625 39.860 149.735 ;
        RECT 40.205 149.595 40.375 149.785 ;
        RECT 43.425 149.595 43.595 149.785 ;
        RECT 44.805 149.595 44.975 149.785 ;
        RECT 46.645 149.575 46.815 149.765 ;
        RECT 47.105 149.575 47.275 149.765 ;
        RECT 48.025 149.595 48.195 149.785 ;
        RECT 48.940 149.625 49.060 149.735 ;
        RECT 49.410 149.595 49.580 149.815 ;
        RECT 51.070 149.785 52.015 149.815 ;
        RECT 52.485 149.785 60.045 150.695 ;
        RECT 60.305 149.785 63.960 150.695 ;
        RECT 63.985 149.785 65.335 150.695 ;
        RECT 65.365 149.785 70.875 150.595 ;
        RECT 70.885 149.785 73.635 150.595 ;
        RECT 73.665 149.785 75.015 150.695 ;
        RECT 75.025 149.785 76.375 150.695 ;
        RECT 76.405 149.785 77.775 150.595 ;
        RECT 77.795 149.870 78.225 150.655 ;
        RECT 78.245 149.785 83.755 150.595 ;
        RECT 83.765 149.785 89.275 150.595 ;
        RECT 89.285 149.785 90.655 150.595 ;
        RECT 90.665 149.785 92.035 150.595 ;
        RECT 103.770 150.080 106.560 152.160 ;
        RECT 51.705 149.575 51.875 149.765 ;
        RECT 52.165 149.575 52.335 149.765 ;
        RECT 52.630 149.595 52.800 149.785 ;
        RECT 57.685 149.575 57.855 149.765 ;
        RECT 59.065 149.595 59.235 149.765 ;
        RECT 60.450 149.595 60.620 149.785 ;
        RECT 59.070 149.575 59.235 149.595 ;
        RECT 61.370 149.575 61.540 149.765 ;
        RECT 65.050 149.595 65.220 149.785 ;
        RECT 65.505 149.765 65.675 149.785 ;
        RECT 71.025 149.765 71.195 149.785 ;
        RECT 65.505 149.595 65.680 149.765 ;
        RECT 65.510 149.575 65.680 149.595 ;
        RECT 71.020 149.595 71.195 149.765 ;
        RECT 71.020 149.575 71.190 149.595 ;
        RECT 71.485 149.575 71.655 149.765 ;
        RECT 74.700 149.595 74.870 149.785 ;
        RECT 75.170 149.765 75.340 149.785 ;
        RECT 75.165 149.595 75.340 149.765 ;
        RECT 76.545 149.595 76.715 149.785 ;
        RECT 78.385 149.595 78.555 149.785 ;
        RECT 75.165 149.575 75.335 149.595 ;
        RECT 82.525 149.575 82.695 149.765 ;
        RECT 83.905 149.595 84.075 149.785 ;
        RECT 88.045 149.575 88.215 149.765 ;
        RECT 89.425 149.595 89.595 149.785 ;
        RECT 91.725 149.575 91.895 149.785 ;
        RECT 20.285 149.345 23.350 149.545 ;
        RECT 20.285 148.865 23.495 149.345 ;
        RECT 20.285 148.665 21.235 148.865 ;
        RECT 22.565 148.665 23.495 148.865 ;
        RECT 23.965 148.895 26.255 149.575 ;
        RECT 23.965 148.665 24.885 148.895 ;
        RECT 26.265 148.765 31.775 149.575 ;
        RECT 31.785 148.665 34.850 149.575 ;
        RECT 35.005 148.765 38.675 149.575 ;
        RECT 39.155 148.705 39.585 149.490 ;
        RECT 39.645 148.895 46.955 149.575 ;
        RECT 39.645 148.665 40.995 148.895 ;
        RECT 42.530 148.675 43.440 148.895 ;
        RECT 46.965 148.765 48.795 149.575 ;
        RECT 49.275 148.665 52.005 149.575 ;
        RECT 52.025 148.765 57.535 149.575 ;
        RECT 57.545 148.765 58.915 149.575 ;
        RECT 59.070 148.895 60.905 149.575 ;
        RECT 59.975 148.665 60.905 148.895 ;
        RECT 61.225 148.665 64.700 149.575 ;
        RECT 64.915 148.705 65.345 149.490 ;
        RECT 65.365 148.665 68.840 149.575 ;
        RECT 69.500 149.345 71.190 149.575 ;
        RECT 69.500 148.665 71.335 149.345 ;
        RECT 71.345 148.895 75.015 149.575 ;
        RECT 75.025 148.895 82.335 149.575 ;
        RECT 74.085 148.665 75.015 148.895 ;
        RECT 78.540 148.675 79.450 148.895 ;
        RECT 80.985 148.665 82.335 148.895 ;
        RECT 82.385 148.765 87.895 149.575 ;
        RECT 87.905 148.765 90.655 149.575 ;
        RECT 90.665 148.765 92.035 149.575 ;
      LAYER nwell ;
        RECT 13.190 145.545 92.230 148.375 ;
        RECT 101.660 147.970 106.500 150.080 ;
        RECT 107.780 149.740 117.970 161.990 ;
      LAYER pwell ;
        RECT 120.330 152.190 126.430 161.980 ;
        RECT 120.330 152.160 126.440 152.190 ;
        RECT 120.530 151.760 121.690 152.160 ;
        RECT 123.650 150.080 126.440 152.160 ;
      LAYER nwell ;
        RECT 121.540 147.970 126.380 150.080 ;
        RECT 127.660 149.740 137.850 161.990 ;
      LAYER pwell ;
        RECT 140.410 152.140 146.510 161.930 ;
        RECT 140.410 152.110 146.520 152.140 ;
        RECT 140.610 151.710 141.770 152.110 ;
        RECT 143.730 150.030 146.520 152.110 ;
      LAYER nwell ;
        RECT 141.620 147.920 146.460 150.030 ;
        RECT 147.740 149.690 157.930 161.940 ;
      LAYER pwell ;
        RECT 13.385 144.345 14.755 145.155 ;
        RECT 14.765 144.345 20.275 145.155 ;
        RECT 20.285 144.345 25.795 145.155 ;
        RECT 26.275 144.430 26.705 145.215 ;
        RECT 26.725 144.345 28.095 145.155 ;
        RECT 28.125 144.345 29.475 145.255 ;
        RECT 30.415 144.345 33.145 145.255 ;
        RECT 35.820 145.025 36.740 145.255 ;
        RECT 37.895 145.025 38.825 145.255 ;
        RECT 33.275 144.345 36.740 145.025 ;
        RECT 36.990 144.345 38.825 145.025 ;
        RECT 39.155 144.345 40.505 145.255 ;
        RECT 43.265 145.025 44.195 145.255 ;
        RECT 40.525 144.345 44.195 145.025 ;
        RECT 44.205 144.345 49.715 145.155 ;
        RECT 49.725 144.345 51.555 145.155 ;
        RECT 52.035 144.430 52.465 145.215 ;
        RECT 59.605 145.165 60.555 145.255 ;
        RECT 52.485 144.345 57.995 145.155 ;
        RECT 58.625 144.345 60.555 145.165 ;
        RECT 60.765 145.055 61.695 145.255 ;
        RECT 63.030 145.055 63.975 145.255 ;
        RECT 60.765 144.575 63.975 145.055 ;
        RECT 60.905 144.375 63.975 144.575 ;
        RECT 13.525 144.135 13.695 144.345 ;
        RECT 14.905 144.135 15.075 144.345 ;
        RECT 20.425 144.135 20.595 144.345 ;
        RECT 25.025 144.155 25.195 144.325 ;
        RECT 25.485 144.155 25.655 144.325 ;
        RECT 25.940 144.185 26.060 144.295 ;
        RECT 26.865 144.155 27.035 144.345 ;
        RECT 25.025 144.135 25.175 144.155 ;
        RECT 13.385 143.325 14.755 144.135 ;
        RECT 14.765 143.325 20.275 144.135 ;
        RECT 20.285 143.325 23.035 144.135 ;
        RECT 23.245 143.315 25.175 144.135 ;
        RECT 25.490 144.135 25.655 144.155 ;
        RECT 25.490 143.455 27.325 144.135 ;
        RECT 27.790 144.105 27.960 144.325 ;
        RECT 28.240 144.155 28.410 144.345 ;
        RECT 29.635 144.190 29.795 144.300 ;
        RECT 30.545 144.155 30.715 144.345 ;
        RECT 31.465 144.135 31.635 144.325 ;
        RECT 33.305 144.155 33.475 144.345 ;
        RECT 36.990 144.325 37.155 144.345 ;
        RECT 36.525 144.155 36.695 144.325 ;
        RECT 36.985 144.155 37.155 144.325 ;
        RECT 39.285 144.155 39.455 144.345 ;
        RECT 36.675 144.135 36.695 144.155 ;
        RECT 39.745 144.135 39.915 144.325 ;
        RECT 40.665 144.155 40.835 144.345 ;
        RECT 43.425 144.135 43.595 144.325 ;
        RECT 43.895 144.180 44.055 144.290 ;
        RECT 44.345 144.155 44.515 144.345 ;
        RECT 45.720 144.135 45.890 144.325 ;
        RECT 46.185 144.135 46.355 144.325 ;
        RECT 48.020 144.185 48.140 144.295 ;
        RECT 49.400 144.135 49.570 144.325 ;
        RECT 49.865 144.155 50.035 144.345 ;
        RECT 51.245 144.135 51.415 144.325 ;
        RECT 51.700 144.185 51.820 144.295 ;
        RECT 52.625 144.155 52.795 144.345 ;
        RECT 58.625 144.325 58.775 144.345 ;
        RECT 58.140 144.185 58.260 144.295 ;
        RECT 58.605 144.135 58.775 144.325 ;
        RECT 59.075 144.180 59.235 144.290 ;
        RECT 59.985 144.135 60.155 144.325 ;
        RECT 60.905 144.155 61.075 144.375 ;
        RECT 63.030 144.345 63.975 144.375 ;
        RECT 63.985 144.345 67.145 145.255 ;
        RECT 72.275 145.025 75.275 145.255 ;
        RECT 67.205 144.345 72.020 145.025 ;
        RECT 72.275 144.935 76.855 145.025 ;
        RECT 72.265 144.575 76.855 144.935 ;
        RECT 72.265 144.385 73.195 144.575 ;
        RECT 72.275 144.345 73.195 144.385 ;
        RECT 75.285 144.345 76.855 144.575 ;
        RECT 77.795 144.430 78.225 145.215 ;
        RECT 78.245 144.345 79.615 145.125 ;
        RECT 79.625 144.345 85.135 145.155 ;
        RECT 85.145 144.345 90.655 145.155 ;
        RECT 90.665 144.345 92.035 145.155 ;
        RECT 63.205 144.135 63.375 144.325 ;
        RECT 65.505 144.135 65.675 144.325 ;
        RECT 66.885 144.155 67.055 144.345 ;
        RECT 67.345 144.155 67.515 144.345 ;
        RECT 68.265 144.135 68.435 144.325 ;
        RECT 70.105 144.135 70.275 144.325 ;
        RECT 76.545 144.155 76.715 144.345 ;
        RECT 77.015 144.190 77.175 144.300 ;
        RECT 77.465 144.135 77.635 144.325 ;
        RECT 79.305 144.155 79.475 144.345 ;
        RECT 79.765 144.155 79.935 144.345 ;
        RECT 82.985 144.135 83.155 144.325 ;
        RECT 85.285 144.155 85.455 144.345 ;
        RECT 88.505 144.135 88.675 144.325 ;
        RECT 90.340 144.185 90.460 144.295 ;
        RECT 91.725 144.135 91.895 144.345 ;
        RECT 30.365 144.105 31.315 144.135 ;
        RECT 23.245 143.225 24.195 143.315 ;
        RECT 26.395 143.225 27.325 143.455 ;
        RECT 27.645 143.425 31.315 144.105 ;
        RECT 31.325 143.455 36.140 144.135 ;
        RECT 36.675 143.455 39.125 144.135 ;
        RECT 30.365 143.225 31.315 143.425 ;
        RECT 37.165 143.225 39.125 143.455 ;
        RECT 39.155 143.265 39.585 144.050 ;
        RECT 39.605 143.325 41.695 144.135 ;
        RECT 42.365 143.355 43.735 144.135 ;
        RECT 44.685 143.225 46.035 144.135 ;
        RECT 46.045 143.325 47.875 144.135 ;
        RECT 48.365 143.225 49.715 144.135 ;
        RECT 49.725 143.455 51.555 144.135 ;
        RECT 51.605 143.455 58.915 144.135 ;
        RECT 51.605 143.225 52.955 143.455 ;
        RECT 54.490 143.235 55.400 143.455 ;
        RECT 59.845 143.225 63.055 144.135 ;
        RECT 63.065 143.325 64.895 144.135 ;
        RECT 64.915 143.265 65.345 144.050 ;
        RECT 65.365 143.225 68.115 144.135 ;
        RECT 68.125 143.325 69.955 144.135 ;
        RECT 69.965 143.455 77.275 144.135 ;
        RECT 73.480 143.235 74.390 143.455 ;
        RECT 75.925 143.225 77.275 143.455 ;
        RECT 77.325 143.325 82.835 144.135 ;
        RECT 82.845 143.325 88.355 144.135 ;
        RECT 88.365 143.325 90.195 144.135 ;
        RECT 90.665 143.325 92.035 144.135 ;
      LAYER nwell ;
        RECT 13.190 140.105 92.230 142.935 ;
      LAYER pwell ;
        RECT 13.385 138.905 14.755 139.715 ;
        RECT 14.765 138.905 18.435 139.715 ;
        RECT 22.420 139.585 23.330 139.805 ;
        RECT 24.865 139.585 26.215 139.815 ;
        RECT 18.905 138.905 26.215 139.585 ;
        RECT 26.275 138.990 26.705 139.775 ;
        RECT 29.065 139.585 30.415 139.815 ;
        RECT 31.950 139.585 32.860 139.805 ;
        RECT 36.480 139.585 37.400 139.815 ;
        RECT 27.185 138.905 29.015 139.585 ;
        RECT 29.065 138.905 36.375 139.585 ;
        RECT 36.480 138.905 39.945 139.585 ;
        RECT 40.065 138.905 41.895 139.715 ;
        RECT 45.420 139.585 46.330 139.805 ;
        RECT 47.865 139.585 49.215 139.815 ;
        RECT 51.095 139.585 52.015 139.815 ;
        RECT 41.905 138.905 49.215 139.585 ;
        RECT 49.725 138.905 52.015 139.585 ;
        RECT 52.035 138.990 52.465 139.775 ;
        RECT 55.225 139.585 56.155 139.815 ;
        RECT 52.485 138.905 56.155 139.585 ;
        RECT 56.180 138.905 57.995 139.815 ;
        RECT 58.240 138.905 63.055 139.585 ;
        RECT 63.065 138.905 64.435 139.715 ;
        RECT 64.445 139.585 65.580 139.815 ;
        RECT 64.445 138.905 67.655 139.585 ;
        RECT 67.665 138.905 73.175 139.715 ;
        RECT 73.185 138.905 76.855 139.715 ;
        RECT 77.795 138.990 78.225 139.775 ;
        RECT 78.245 138.905 83.755 139.715 ;
        RECT 83.765 138.905 89.275 139.715 ;
        RECT 89.285 138.905 90.655 139.715 ;
        RECT 90.665 138.905 92.035 139.715 ;
        RECT 13.525 138.695 13.695 138.905 ;
        RECT 14.905 138.715 15.075 138.905 ;
        RECT 16.285 138.695 16.455 138.885 ;
        RECT 16.745 138.695 16.915 138.885 ;
        RECT 18.580 138.745 18.700 138.855 ;
        RECT 19.045 138.715 19.215 138.905 ;
        RECT 20.435 138.740 20.595 138.850 ;
        RECT 13.385 137.885 14.755 138.695 ;
        RECT 14.765 138.015 16.595 138.695 ;
        RECT 14.765 137.785 16.110 138.015 ;
        RECT 16.605 137.885 20.275 138.695 ;
        RECT 21.205 138.665 22.140 138.695 ;
        RECT 24.100 138.665 24.270 138.885 ;
        RECT 24.565 138.695 24.735 138.885 ;
        RECT 25.945 138.715 26.115 138.885 ;
        RECT 26.860 138.745 26.980 138.855 ;
        RECT 27.325 138.715 27.495 138.905 ;
        RECT 25.950 138.695 26.115 138.715 ;
        RECT 28.245 138.695 28.415 138.885 ;
        RECT 30.545 138.695 30.715 138.885 ;
        RECT 36.065 138.715 36.235 138.905 ;
        RECT 37.905 138.695 38.075 138.885 ;
        RECT 39.745 138.715 39.915 138.905 ;
        RECT 40.205 138.715 40.375 138.905 ;
        RECT 40.665 138.695 40.835 138.885 ;
        RECT 42.045 138.715 42.215 138.905 ;
        RECT 48.945 138.695 49.115 138.885 ;
        RECT 49.400 138.745 49.520 138.855 ;
        RECT 49.865 138.715 50.035 138.905 ;
        RECT 52.165 138.695 52.335 138.885 ;
        RECT 52.625 138.715 52.795 138.905 ;
        RECT 53.540 138.695 53.710 138.885 ;
        RECT 54.005 138.695 54.175 138.885 ;
        RECT 56.305 138.715 56.475 138.905 ;
        RECT 57.680 138.745 57.800 138.855 ;
        RECT 58.145 138.695 58.315 138.885 ;
        RECT 61.365 138.695 61.535 138.885 ;
        RECT 62.745 138.715 62.915 138.905 ;
        RECT 63.205 138.715 63.375 138.905 ;
        RECT 65.505 138.695 65.675 138.885 ;
        RECT 67.345 138.715 67.515 138.905 ;
        RECT 67.805 138.715 67.975 138.905 ;
        RECT 68.260 138.695 68.430 138.885 ;
        RECT 68.725 138.695 68.895 138.885 ;
        RECT 70.105 138.695 70.275 138.885 ;
        RECT 73.325 138.715 73.495 138.905 ;
        RECT 77.015 138.750 77.175 138.860 ;
        RECT 78.385 138.715 78.555 138.905 ;
        RECT 80.685 138.695 80.855 138.885 ;
        RECT 81.145 138.695 81.315 138.885 ;
        RECT 83.905 138.715 84.075 138.905 ;
        RECT 86.665 138.695 86.835 138.885 ;
        RECT 89.425 138.715 89.595 138.905 ;
        RECT 90.340 138.745 90.460 138.855 ;
        RECT 91.725 138.695 91.895 138.905 ;
        RECT 21.205 138.465 24.270 138.665 ;
        RECT 21.205 137.985 24.415 138.465 ;
        RECT 21.205 137.785 22.155 137.985 ;
        RECT 23.485 137.785 24.415 137.985 ;
        RECT 24.425 137.885 25.795 138.695 ;
        RECT 25.950 138.015 27.785 138.695 ;
        RECT 28.105 138.015 30.395 138.695 ;
        RECT 30.405 138.015 37.715 138.695 ;
        RECT 26.855 137.785 27.785 138.015 ;
        RECT 29.475 137.785 30.395 138.015 ;
        RECT 33.920 137.795 34.830 138.015 ;
        RECT 36.365 137.785 37.715 138.015 ;
        RECT 37.765 137.885 39.135 138.695 ;
        RECT 39.155 137.825 39.585 138.610 ;
        RECT 40.525 138.015 45.340 138.695 ;
        RECT 45.585 138.015 49.255 138.695 ;
        RECT 49.265 138.015 52.475 138.695 ;
        RECT 45.585 137.785 46.515 138.015 ;
        RECT 49.265 137.785 50.400 138.015 ;
        RECT 52.505 137.785 53.855 138.695 ;
        RECT 53.865 137.885 57.535 138.695 ;
        RECT 58.055 137.785 61.215 138.695 ;
        RECT 61.225 137.885 64.895 138.695 ;
        RECT 64.915 137.825 65.345 138.610 ;
        RECT 65.365 137.885 67.195 138.695 ;
        RECT 67.225 137.785 68.575 138.695 ;
        RECT 68.585 137.885 69.955 138.695 ;
        RECT 69.965 138.015 73.635 138.695 ;
        RECT 72.705 137.785 73.635 138.015 ;
        RECT 73.685 138.015 80.995 138.695 ;
        RECT 73.685 137.785 75.035 138.015 ;
        RECT 76.570 137.795 77.480 138.015 ;
        RECT 81.005 137.885 86.515 138.695 ;
        RECT 86.525 137.885 90.195 138.695 ;
        RECT 90.665 137.885 92.035 138.695 ;
      LAYER nwell ;
        RECT 13.190 134.665 92.230 137.495 ;
      LAYER pwell ;
        RECT 100.450 137.140 106.550 146.930 ;
        RECT 100.450 137.110 106.560 137.140 ;
        RECT 100.650 136.710 101.810 137.110 ;
        RECT 103.770 135.030 106.560 137.110 ;
        RECT 13.385 133.465 14.755 134.275 ;
        RECT 14.765 133.465 20.275 134.275 ;
        RECT 20.285 133.465 25.795 134.275 ;
        RECT 26.275 133.550 26.705 134.335 ;
        RECT 26.725 133.465 30.395 134.275 ;
        RECT 31.325 133.465 33.415 134.275 ;
        RECT 34.100 133.465 35.915 134.375 ;
        RECT 35.925 133.465 37.755 134.275 ;
        RECT 41.740 134.145 42.650 134.365 ;
        RECT 44.185 134.145 45.535 134.375 ;
        RECT 38.225 133.465 45.535 134.145 ;
        RECT 45.585 133.465 51.095 134.275 ;
        RECT 52.035 133.550 52.465 134.335 ;
        RECT 52.485 133.465 54.315 134.145 ;
        RECT 54.325 133.465 57.995 134.275 ;
        RECT 60.745 134.145 61.675 134.375 ;
        RECT 58.005 133.465 61.675 134.145 ;
        RECT 61.705 133.465 63.055 134.375 ;
        RECT 63.545 133.465 64.895 134.375 ;
        RECT 65.825 134.145 66.745 134.375 ;
        RECT 65.825 133.465 68.115 134.145 ;
        RECT 68.140 133.465 69.955 134.375 ;
        RECT 70.925 133.465 74.095 134.375 ;
        RECT 74.105 133.465 77.775 134.275 ;
        RECT 77.795 133.550 78.225 134.335 ;
        RECT 78.245 133.465 83.755 134.275 ;
        RECT 83.765 133.465 89.275 134.275 ;
        RECT 89.285 133.465 90.655 134.275 ;
        RECT 90.665 133.465 92.035 134.275 ;
        RECT 13.525 133.255 13.695 133.465 ;
        RECT 14.905 133.255 15.075 133.465 ;
        RECT 20.425 133.255 20.595 133.465 ;
        RECT 25.945 133.415 26.115 133.445 ;
        RECT 25.940 133.305 26.115 133.415 ;
        RECT 25.945 133.255 26.115 133.305 ;
        RECT 26.865 133.275 27.035 133.465 ;
        RECT 13.385 132.445 14.755 133.255 ;
        RECT 14.765 132.445 20.275 133.255 ;
        RECT 20.285 132.445 25.795 133.255 ;
        RECT 25.805 132.445 27.175 133.255 ;
        RECT 27.185 133.225 28.120 133.255 ;
        RECT 30.080 133.225 30.250 133.445 ;
        RECT 30.555 133.415 30.715 133.420 ;
        RECT 30.540 133.310 30.715 133.415 ;
        RECT 30.540 133.305 30.660 133.310 ;
        RECT 31.005 133.255 31.175 133.445 ;
        RECT 31.465 133.275 31.635 133.465 ;
        RECT 34.225 133.275 34.395 133.465 ;
        RECT 34.695 133.300 34.855 133.410 ;
        RECT 35.605 133.255 35.775 133.445 ;
        RECT 36.065 133.275 36.235 133.465 ;
        RECT 37.900 133.305 38.020 133.415 ;
        RECT 38.365 133.275 38.535 133.465 ;
        RECT 39.745 133.255 39.915 133.445 ;
        RECT 41.585 133.255 41.755 133.445 ;
        RECT 45.725 133.275 45.895 133.465 ;
        RECT 46.185 133.255 46.355 133.445 ;
        RECT 47.570 133.255 47.740 133.445 ;
        RECT 48.035 133.300 48.195 133.410 ;
        RECT 48.945 133.255 49.115 133.445 ;
        RECT 51.255 133.310 51.415 133.420 ;
        RECT 52.165 133.255 52.335 133.445 ;
        RECT 54.005 133.275 54.175 133.465 ;
        RECT 54.465 133.275 54.635 133.465 ;
        RECT 55.845 133.255 56.015 133.445 ;
        RECT 57.685 133.255 57.855 133.445 ;
        RECT 58.145 133.275 58.315 133.465 ;
        RECT 62.740 133.275 62.910 133.465 ;
        RECT 63.200 133.305 63.320 133.415 ;
        RECT 64.580 133.275 64.750 133.465 ;
        RECT 65.055 133.310 65.215 133.420 ;
        RECT 65.515 133.300 65.675 133.410 ;
        RECT 66.425 133.255 66.595 133.445 ;
        RECT 67.805 133.275 67.975 133.465 ;
        RECT 68.265 133.275 68.435 133.465 ;
        RECT 70.115 133.310 70.275 133.420 ;
        RECT 71.025 133.275 71.195 133.465 ;
        RECT 73.785 133.255 73.955 133.445 ;
        RECT 74.245 133.275 74.415 133.465 ;
        RECT 78.385 133.275 78.555 133.465 ;
        RECT 79.305 133.255 79.475 133.445 ;
        RECT 83.905 133.275 84.075 133.465 ;
        RECT 84.825 133.255 84.995 133.445 ;
        RECT 89.425 133.275 89.595 133.465 ;
        RECT 90.340 133.305 90.460 133.415 ;
        RECT 91.725 133.255 91.895 133.465 ;
        RECT 27.185 133.025 30.250 133.225 ;
        RECT 27.185 132.545 30.395 133.025 ;
        RECT 30.975 132.575 34.440 133.255 ;
        RECT 35.575 132.575 39.040 133.255 ;
        RECT 27.185 132.345 28.135 132.545 ;
        RECT 29.465 132.345 30.395 132.545 ;
        RECT 33.520 132.345 34.440 132.575 ;
        RECT 38.120 132.345 39.040 132.575 ;
        RECT 39.155 132.385 39.585 133.170 ;
        RECT 39.620 132.345 41.435 133.255 ;
        RECT 41.445 132.445 42.815 133.255 ;
        RECT 42.920 132.575 46.385 133.255 ;
        RECT 42.920 132.345 43.840 132.575 ;
        RECT 46.505 132.345 47.855 133.255 ;
        RECT 48.845 132.345 52.015 133.255 ;
        RECT 52.025 132.575 55.695 133.255 ;
        RECT 54.765 132.345 55.695 132.575 ;
        RECT 55.705 132.445 57.535 133.255 ;
        RECT 57.545 132.575 64.855 133.255 ;
        RECT 61.060 132.355 61.970 132.575 ;
        RECT 63.505 132.345 64.855 132.575 ;
        RECT 64.915 132.385 65.345 133.170 ;
        RECT 66.285 132.575 73.595 133.255 ;
        RECT 69.800 132.355 70.710 132.575 ;
        RECT 72.245 132.345 73.595 132.575 ;
        RECT 73.645 132.445 79.155 133.255 ;
        RECT 79.165 132.445 84.675 133.255 ;
        RECT 84.685 132.445 90.195 133.255 ;
        RECT 90.665 132.445 92.035 133.255 ;
      LAYER nwell ;
        RECT 101.660 132.920 106.500 135.030 ;
        RECT 107.780 134.690 117.970 146.940 ;
      LAYER pwell ;
        RECT 120.330 137.140 126.430 146.930 ;
        RECT 120.330 137.110 126.440 137.140 ;
        RECT 120.530 136.710 121.690 137.110 ;
        RECT 123.650 135.030 126.440 137.110 ;
      LAYER nwell ;
        RECT 121.540 132.920 126.380 135.030 ;
        RECT 127.660 134.690 137.850 146.940 ;
      LAYER pwell ;
        RECT 140.360 137.140 146.460 146.930 ;
        RECT 140.360 137.110 146.470 137.140 ;
        RECT 140.560 136.710 141.720 137.110 ;
        RECT 143.680 135.030 146.470 137.110 ;
      LAYER nwell ;
        RECT 141.570 132.920 146.410 135.030 ;
        RECT 147.690 134.690 157.880 146.940 ;
        RECT 13.190 129.225 92.230 132.055 ;
      LAYER pwell ;
        RECT 13.385 128.025 14.755 128.835 ;
        RECT 14.765 128.025 20.275 128.835 ;
        RECT 20.285 128.025 25.795 128.835 ;
        RECT 26.275 128.110 26.705 128.895 ;
        RECT 26.765 128.705 28.115 128.935 ;
        RECT 29.650 128.705 30.560 128.925 ;
        RECT 34.395 128.705 35.325 128.935 ;
        RECT 39.900 128.705 40.810 128.925 ;
        RECT 42.345 128.705 43.695 128.935 ;
        RECT 46.495 128.705 47.415 128.935 ;
        RECT 26.765 128.025 34.075 128.705 ;
        RECT 34.395 128.025 36.230 128.705 ;
        RECT 36.385 128.025 43.695 128.705 ;
        RECT 43.830 128.025 47.415 128.705 ;
        RECT 47.520 128.705 48.440 128.935 ;
        RECT 47.520 128.025 50.985 128.705 ;
        RECT 52.035 128.110 52.465 128.895 ;
        RECT 52.485 128.025 53.835 128.935 ;
        RECT 57.380 128.705 58.290 128.925 ;
        RECT 59.825 128.705 61.175 128.935 ;
        RECT 53.865 128.025 61.175 128.705 ;
        RECT 61.225 128.025 64.895 128.835 ;
        RECT 68.105 128.705 69.035 128.935 ;
        RECT 65.365 128.025 69.035 128.705 ;
        RECT 69.045 128.025 74.555 128.835 ;
        RECT 74.565 128.025 77.315 128.835 ;
        RECT 77.795 128.110 78.225 128.895 ;
        RECT 78.245 128.025 83.755 128.835 ;
        RECT 83.765 128.025 89.275 128.835 ;
        RECT 89.285 128.025 90.655 128.835 ;
        RECT 90.665 128.025 92.035 128.835 ;
        RECT 13.525 127.815 13.695 128.025 ;
        RECT 14.905 127.815 15.075 128.025 ;
        RECT 20.425 127.815 20.595 128.025 ;
        RECT 25.945 127.975 26.115 128.005 ;
        RECT 25.940 127.865 26.115 127.975 ;
        RECT 25.945 127.815 26.115 127.865 ;
        RECT 33.765 127.835 33.935 128.025 ;
        RECT 36.065 128.005 36.230 128.025 ;
        RECT 35.605 127.815 35.775 128.005 ;
        RECT 36.065 127.835 36.235 128.005 ;
        RECT 36.525 127.835 36.695 128.025 ;
        RECT 38.825 127.815 38.995 128.005 ;
        RECT 39.755 127.860 39.915 127.970 ;
        RECT 40.665 127.815 40.835 128.005 ;
        RECT 47.100 127.835 47.270 128.025 ;
        RECT 47.560 127.815 47.730 128.005 ;
        RECT 48.025 127.815 48.195 128.005 ;
        RECT 50.785 127.835 50.955 128.025 ;
        RECT 51.255 127.870 51.415 127.980 ;
        RECT 53.550 127.835 53.720 128.025 ;
        RECT 54.005 127.835 54.175 128.025 ;
        RECT 55.385 127.815 55.555 128.005 ;
        RECT 60.905 127.815 61.075 128.005 ;
        RECT 61.365 127.835 61.535 128.025 ;
        RECT 64.580 127.865 64.700 127.975 ;
        RECT 65.040 127.865 65.160 127.975 ;
        RECT 65.505 127.815 65.675 128.025 ;
        RECT 69.185 127.835 69.355 128.025 ;
        RECT 71.025 127.815 71.195 128.005 ;
        RECT 74.705 127.835 74.875 128.025 ;
        RECT 76.545 127.815 76.715 128.005 ;
        RECT 77.460 127.865 77.580 127.975 ;
        RECT 78.385 127.835 78.555 128.025 ;
        RECT 82.065 127.815 82.235 128.005 ;
        RECT 83.905 127.835 84.075 128.025 ;
        RECT 87.585 127.815 87.755 128.005 ;
        RECT 89.425 127.835 89.595 128.025 ;
        RECT 90.340 127.865 90.460 127.975 ;
        RECT 91.725 127.815 91.895 128.025 ;
        RECT 13.385 127.005 14.755 127.815 ;
        RECT 14.765 127.005 20.275 127.815 ;
        RECT 20.285 127.005 25.795 127.815 ;
        RECT 25.805 127.005 28.555 127.815 ;
        RECT 28.605 127.135 35.915 127.815 ;
        RECT 28.605 126.905 29.955 127.135 ;
        RECT 31.490 126.915 32.400 127.135 ;
        RECT 35.925 126.905 39.035 127.815 ;
        RECT 39.155 126.945 39.585 127.730 ;
        RECT 40.635 127.135 44.100 127.815 ;
        RECT 44.290 127.135 47.875 127.815 ;
        RECT 47.885 127.135 55.195 127.815 ;
        RECT 43.180 126.905 44.100 127.135 ;
        RECT 46.955 126.905 47.875 127.135 ;
        RECT 51.400 126.915 52.310 127.135 ;
        RECT 53.845 126.905 55.195 127.135 ;
        RECT 55.245 127.005 60.755 127.815 ;
        RECT 60.765 127.005 64.435 127.815 ;
        RECT 64.915 126.945 65.345 127.730 ;
        RECT 65.365 127.005 70.875 127.815 ;
        RECT 70.885 127.005 76.395 127.815 ;
        RECT 76.405 127.005 81.915 127.815 ;
        RECT 81.925 127.005 87.435 127.815 ;
        RECT 87.445 127.005 90.195 127.815 ;
        RECT 90.665 127.005 92.035 127.815 ;
      LAYER nwell ;
        RECT 13.190 123.785 92.230 126.615 ;
      LAYER pwell ;
        RECT 13.385 122.585 14.755 123.395 ;
        RECT 14.765 122.585 20.275 123.395 ;
        RECT 20.285 122.585 25.795 123.395 ;
        RECT 26.275 122.670 26.705 123.455 ;
        RECT 26.725 122.585 28.095 123.395 ;
        RECT 30.760 123.265 31.680 123.495 ;
        RECT 28.215 122.585 31.680 123.265 ;
        RECT 31.785 122.585 34.535 123.395 ;
        RECT 35.015 122.585 38.675 123.495 ;
        RECT 38.715 122.585 41.435 123.495 ;
        RECT 44.960 123.265 45.870 123.485 ;
        RECT 47.405 123.265 48.755 123.495 ;
        RECT 50.140 123.295 51.095 123.495 ;
        RECT 41.445 122.585 48.755 123.265 ;
        RECT 48.815 122.615 51.095 123.295 ;
        RECT 52.035 122.670 52.465 123.455 ;
        RECT 13.525 122.375 13.695 122.585 ;
        RECT 14.905 122.375 15.075 122.585 ;
        RECT 20.425 122.375 20.595 122.585 ;
        RECT 23.185 122.375 23.355 122.565 ;
        RECT 25.940 122.425 26.060 122.535 ;
        RECT 26.865 122.395 27.035 122.585 ;
        RECT 28.245 122.395 28.415 122.585 ;
        RECT 30.545 122.375 30.715 122.565 ;
        RECT 31.925 122.395 32.095 122.585 ;
        RECT 34.680 122.425 34.800 122.535 ;
        RECT 35.140 122.395 35.310 122.585 ;
        RECT 36.065 122.375 36.235 122.565 ;
        RECT 38.820 122.425 38.940 122.535 ;
        RECT 39.745 122.375 39.915 122.565 ;
        RECT 41.125 122.395 41.295 122.585 ;
        RECT 41.585 122.395 41.755 122.585 ;
        RECT 47.105 122.395 47.275 122.565 ;
        RECT 47.105 122.375 47.270 122.395 ;
        RECT 48.485 122.375 48.655 122.565 ;
        RECT 48.940 122.395 49.110 122.615 ;
        RECT 50.140 122.585 51.095 122.615 ;
        RECT 52.485 122.585 55.225 123.265 ;
        RECT 55.245 122.585 57.075 123.395 ;
        RECT 57.180 123.265 58.100 123.495 ;
        RECT 57.180 122.585 60.645 123.265 ;
        RECT 60.765 122.585 62.595 123.395 ;
        RECT 62.700 123.265 63.620 123.495 ;
        RECT 62.700 122.585 66.165 123.265 ;
        RECT 66.285 122.585 69.760 123.495 ;
        RECT 69.965 122.585 75.475 123.395 ;
        RECT 75.485 122.585 77.315 123.395 ;
        RECT 77.795 122.670 78.225 123.455 ;
        RECT 78.245 122.585 83.755 123.395 ;
        RECT 83.765 122.585 89.275 123.395 ;
        RECT 89.285 122.585 90.655 123.395 ;
        RECT 90.665 122.585 92.035 123.395 ;
        RECT 49.860 122.375 50.030 122.565 ;
        RECT 50.325 122.375 50.495 122.565 ;
        RECT 51.255 122.430 51.415 122.540 ;
        RECT 52.625 122.395 52.795 122.585 ;
        RECT 54.005 122.375 54.175 122.565 ;
        RECT 55.385 122.375 55.555 122.585 ;
        RECT 60.445 122.395 60.615 122.585 ;
        RECT 60.905 122.395 61.075 122.585 ;
        RECT 62.750 122.375 62.920 122.565 ;
        RECT 64.135 122.420 64.295 122.530 ;
        RECT 65.505 122.375 65.675 122.565 ;
        RECT 65.965 122.395 66.135 122.585 ;
        RECT 66.430 122.395 66.600 122.585 ;
        RECT 70.105 122.395 70.275 122.585 ;
        RECT 74.245 122.375 74.415 122.565 ;
        RECT 74.705 122.375 74.875 122.565 ;
        RECT 75.625 122.395 75.795 122.585 ;
        RECT 77.460 122.425 77.580 122.535 ;
        RECT 78.385 122.395 78.555 122.585 ;
        RECT 80.225 122.375 80.395 122.565 ;
        RECT 83.905 122.395 84.075 122.585 ;
        RECT 85.745 122.375 85.915 122.565 ;
        RECT 89.425 122.375 89.595 122.585 ;
        RECT 91.725 122.375 91.895 122.585 ;
        RECT 13.385 121.565 14.755 122.375 ;
        RECT 14.765 121.565 20.275 122.375 ;
        RECT 20.285 121.565 23.035 122.375 ;
        RECT 23.045 121.695 30.355 122.375 ;
        RECT 26.560 121.475 27.470 121.695 ;
        RECT 29.005 121.465 30.355 121.695 ;
        RECT 30.405 121.565 35.915 122.375 ;
        RECT 35.925 121.565 38.675 122.375 ;
        RECT 39.155 121.505 39.585 122.290 ;
        RECT 39.605 121.565 45.115 122.375 ;
        RECT 45.435 121.695 47.270 122.375 ;
        RECT 45.435 121.465 46.365 121.695 ;
        RECT 47.435 121.465 48.785 122.375 ;
        RECT 48.825 121.465 50.175 122.375 ;
        RECT 50.185 121.565 53.855 122.375 ;
        RECT 53.865 121.565 55.235 122.375 ;
        RECT 55.245 121.695 62.555 122.375 ;
        RECT 58.760 121.475 59.670 121.695 ;
        RECT 61.205 121.465 62.555 121.695 ;
        RECT 62.605 121.465 63.955 122.375 ;
        RECT 64.915 121.505 65.345 122.290 ;
        RECT 65.365 121.565 67.195 122.375 ;
        RECT 67.245 121.695 74.555 122.375 ;
        RECT 67.245 121.465 68.595 121.695 ;
        RECT 70.130 121.475 71.040 121.695 ;
        RECT 74.565 121.565 80.075 122.375 ;
        RECT 80.085 121.565 85.595 122.375 ;
        RECT 85.605 121.565 89.275 122.375 ;
        RECT 89.285 121.565 90.655 122.375 ;
        RECT 90.665 121.565 92.035 122.375 ;
        RECT 100.450 122.140 106.550 131.930 ;
        RECT 100.450 122.110 106.560 122.140 ;
        RECT 100.650 121.710 101.810 122.110 ;
      LAYER nwell ;
        RECT 13.190 118.345 92.230 121.175 ;
      LAYER pwell ;
        RECT 103.770 120.030 106.560 122.110 ;
        RECT 13.385 117.145 14.755 117.955 ;
        RECT 14.765 117.145 16.135 117.955 ;
        RECT 16.185 117.825 17.535 118.055 ;
        RECT 19.070 117.825 19.980 118.045 ;
        RECT 16.185 117.145 23.495 117.825 ;
        RECT 23.505 117.145 26.255 118.055 ;
        RECT 26.275 117.230 26.705 118.015 ;
        RECT 30.240 117.825 31.150 118.045 ;
        RECT 32.685 117.825 34.035 118.055 ;
        RECT 26.725 117.145 34.035 117.825 ;
        RECT 34.180 117.825 35.100 118.055 ;
        RECT 38.320 117.825 39.240 118.055 ;
        RECT 34.180 117.145 37.645 117.825 ;
        RECT 38.320 117.145 41.785 117.825 ;
        RECT 41.905 117.145 47.415 117.955 ;
        RECT 47.425 117.145 51.095 117.955 ;
        RECT 52.035 117.230 52.465 118.015 ;
        RECT 56.000 117.825 56.910 118.045 ;
        RECT 58.445 117.825 59.795 118.055 ;
        RECT 63.820 117.825 64.730 118.045 ;
        RECT 66.265 117.825 67.615 118.055 ;
        RECT 52.485 117.145 59.795 117.825 ;
        RECT 60.305 117.145 67.615 117.825 ;
        RECT 67.760 117.825 68.680 118.055 ;
        RECT 67.760 117.145 71.225 117.825 ;
        RECT 71.345 117.145 74.555 118.055 ;
        RECT 74.565 117.145 77.315 117.955 ;
        RECT 77.795 117.230 78.225 118.015 ;
        RECT 78.245 117.145 83.755 117.955 ;
        RECT 83.765 117.145 89.275 117.955 ;
        RECT 89.285 117.145 90.655 117.955 ;
        RECT 90.665 117.145 92.035 117.955 ;
      LAYER nwell ;
        RECT 101.660 117.920 106.500 120.030 ;
        RECT 107.780 119.690 117.970 131.940 ;
      LAYER pwell ;
        RECT 120.330 122.200 126.430 131.990 ;
        RECT 120.330 122.170 126.440 122.200 ;
        RECT 120.530 121.770 121.690 122.170 ;
        RECT 123.650 120.090 126.440 122.170 ;
      LAYER nwell ;
        RECT 121.540 117.980 126.380 120.090 ;
        RECT 127.660 119.750 137.850 132.000 ;
      LAYER pwell ;
        RECT 140.360 122.200 146.460 131.990 ;
        RECT 140.360 122.170 146.470 122.200 ;
        RECT 140.560 121.770 141.720 122.170 ;
        RECT 143.680 120.090 146.470 122.170 ;
      LAYER nwell ;
        RECT 141.570 117.980 146.410 120.090 ;
        RECT 147.690 119.750 157.880 132.000 ;
      LAYER pwell ;
        RECT 13.525 116.935 13.695 117.145 ;
        RECT 14.905 116.935 15.075 117.145 ;
        RECT 16.745 116.935 16.915 117.125 ;
        RECT 22.265 116.935 22.435 117.125 ;
        RECT 23.185 116.955 23.355 117.145 ;
        RECT 23.645 116.955 23.815 117.145 ;
        RECT 24.105 116.935 24.275 117.125 ;
        RECT 26.865 116.955 27.035 117.145 ;
        RECT 27.785 116.935 27.955 117.125 ;
        RECT 31.465 116.935 31.635 117.125 ;
        RECT 31.930 116.935 32.100 117.125 ;
        RECT 33.305 116.935 33.475 117.125 ;
        RECT 36.070 116.935 36.240 117.125 ;
        RECT 37.445 116.955 37.615 117.145 ;
        RECT 37.900 116.985 38.020 117.095 ;
        RECT 39.740 116.985 39.860 117.095 ;
        RECT 41.130 116.935 41.300 117.125 ;
        RECT 41.585 116.935 41.755 117.145 ;
        RECT 42.045 116.955 42.215 117.145 ;
        RECT 45.260 116.935 45.430 117.125 ;
        RECT 47.565 116.955 47.735 117.145 ;
        RECT 49.865 116.935 50.035 117.125 ;
        RECT 50.325 116.935 50.495 117.125 ;
        RECT 51.255 116.990 51.415 117.100 ;
        RECT 52.625 116.955 52.795 117.145 ;
        RECT 57.685 116.935 57.855 117.125 ;
        RECT 59.980 116.985 60.100 117.095 ;
        RECT 60.445 116.955 60.615 117.145 ;
        RECT 63.205 116.935 63.375 117.125 ;
        RECT 65.500 116.985 65.620 117.095 ;
        RECT 66.890 116.935 67.060 117.125 ;
        RECT 67.345 116.935 67.515 117.125 ;
        RECT 68.730 116.935 68.900 117.125 ;
        RECT 70.105 116.935 70.275 117.125 ;
        RECT 71.025 116.955 71.195 117.145 ;
        RECT 71.485 116.955 71.655 117.145 ;
        RECT 71.940 116.985 72.060 117.095 ;
        RECT 72.405 116.935 72.575 117.125 ;
        RECT 74.705 116.955 74.875 117.145 ;
        RECT 75.165 116.935 75.335 117.125 ;
        RECT 77.460 116.985 77.580 117.095 ;
        RECT 78.385 116.955 78.555 117.145 ;
        RECT 80.685 116.935 80.855 117.125 ;
        RECT 83.905 116.955 84.075 117.145 ;
        RECT 86.205 116.935 86.375 117.125 ;
        RECT 88.965 116.935 89.135 117.125 ;
        RECT 89.425 116.955 89.595 117.145 ;
        RECT 91.725 116.935 91.895 117.145 ;
        RECT 13.385 116.125 14.755 116.935 ;
        RECT 14.765 116.255 16.595 116.935 ;
        RECT 16.605 116.125 22.115 116.935 ;
        RECT 22.125 116.125 23.955 116.935 ;
        RECT 23.980 116.025 25.795 116.935 ;
        RECT 25.805 116.255 28.095 116.935 ;
        RECT 28.200 116.255 31.665 116.935 ;
        RECT 25.805 116.025 26.725 116.255 ;
        RECT 28.200 116.025 29.120 116.255 ;
        RECT 31.785 116.025 33.135 116.935 ;
        RECT 33.165 116.125 35.915 116.935 ;
        RECT 35.925 116.025 38.845 116.935 ;
        RECT 39.155 116.065 39.585 116.850 ;
        RECT 40.065 116.025 41.415 116.935 ;
        RECT 41.555 116.255 45.020 116.935 ;
        RECT 44.100 116.025 45.020 116.255 ;
        RECT 45.145 116.025 46.495 116.935 ;
        RECT 46.600 116.255 50.065 116.935 ;
        RECT 50.185 116.255 57.495 116.935 ;
        RECT 46.600 116.025 47.520 116.255 ;
        RECT 53.700 116.035 54.610 116.255 ;
        RECT 56.145 116.025 57.495 116.255 ;
        RECT 57.545 116.125 63.055 116.935 ;
        RECT 63.065 116.125 64.895 116.935 ;
        RECT 64.915 116.065 65.345 116.850 ;
        RECT 65.825 116.025 67.175 116.935 ;
        RECT 67.205 116.125 68.575 116.935 ;
        RECT 68.585 116.025 69.935 116.935 ;
        RECT 69.965 116.125 71.795 116.935 ;
        RECT 72.265 116.255 75.015 116.935 ;
        RECT 74.085 116.025 75.015 116.255 ;
        RECT 75.025 116.125 80.535 116.935 ;
        RECT 80.545 116.125 86.055 116.935 ;
        RECT 86.065 116.125 88.815 116.935 ;
        RECT 88.825 116.255 90.655 116.935 ;
        RECT 89.310 116.025 90.655 116.255 ;
        RECT 90.665 116.125 92.035 116.935 ;
      LAYER nwell ;
        RECT 13.190 112.905 92.230 115.735 ;
      LAYER pwell ;
        RECT 13.385 111.705 14.755 112.515 ;
        RECT 15.425 112.385 19.355 112.615 ;
        RECT 14.940 111.705 19.355 112.385 ;
        RECT 19.460 112.385 20.380 112.615 ;
        RECT 19.460 111.705 22.925 112.385 ;
        RECT 23.045 111.705 25.795 112.515 ;
        RECT 26.275 111.790 26.705 112.575 ;
        RECT 26.725 111.705 32.235 112.515 ;
        RECT 32.245 111.705 34.075 112.515 ;
        RECT 38.060 112.385 38.970 112.605 ;
        RECT 40.505 112.385 41.855 112.615 ;
        RECT 34.545 111.705 41.855 112.385 ;
        RECT 41.915 111.705 44.645 112.615 ;
        RECT 48.180 112.385 49.090 112.605 ;
        RECT 50.625 112.385 51.975 112.615 ;
        RECT 44.665 111.705 51.975 112.385 ;
        RECT 52.035 111.790 52.465 112.575 ;
        RECT 52.485 111.705 55.235 112.515 ;
        RECT 55.245 112.415 56.175 112.615 ;
        RECT 57.505 112.415 58.455 112.615 ;
        RECT 55.245 111.935 58.455 112.415 ;
        RECT 61.980 112.385 62.890 112.605 ;
        RECT 64.425 112.385 65.775 112.615 ;
        RECT 55.390 111.735 58.455 111.935 ;
        RECT 13.525 111.495 13.695 111.705 ;
        RECT 14.940 111.685 15.050 111.705 ;
        RECT 14.880 111.515 15.075 111.685 ;
        RECT 14.905 111.495 15.075 111.515 ;
        RECT 16.290 111.495 16.460 111.685 ;
        RECT 18.125 111.495 18.295 111.685 ;
        RECT 21.805 111.495 21.975 111.685 ;
        RECT 22.725 111.515 22.895 111.705 ;
        RECT 23.185 111.515 23.355 111.705 ;
        RECT 25.940 111.545 26.060 111.655 ;
        RECT 26.865 111.515 27.035 111.705 ;
        RECT 29.170 111.495 29.340 111.685 ;
        RECT 30.555 111.540 30.715 111.650 ;
        RECT 31.465 111.495 31.635 111.685 ;
        RECT 32.385 111.515 32.555 111.705 ;
        RECT 34.220 111.545 34.340 111.655 ;
        RECT 34.685 111.515 34.855 111.705 ;
        RECT 38.820 111.545 38.940 111.655 ;
        RECT 13.385 110.685 14.755 111.495 ;
        RECT 14.765 110.685 16.135 111.495 ;
        RECT 16.145 110.585 17.975 111.495 ;
        RECT 18.095 110.815 21.560 111.495 ;
        RECT 21.665 110.815 28.975 111.495 ;
        RECT 20.640 110.585 21.560 110.815 ;
        RECT 25.180 110.595 26.090 110.815 ;
        RECT 27.625 110.585 28.975 110.815 ;
        RECT 29.025 110.585 30.375 111.495 ;
        RECT 31.325 110.815 38.635 111.495 ;
        RECT 39.740 111.465 39.910 111.685 ;
        RECT 42.045 111.655 42.215 111.705 ;
        RECT 44.805 111.685 44.975 111.705 ;
        RECT 42.040 111.545 42.215 111.655 ;
        RECT 42.045 111.515 42.215 111.545 ;
        RECT 42.505 111.515 42.675 111.685 ;
        RECT 44.805 111.515 44.980 111.685 ;
        RECT 42.510 111.495 42.675 111.515 ;
        RECT 44.810 111.495 44.980 111.515 ;
        RECT 46.645 111.495 46.815 111.685 ;
        RECT 48.025 111.495 48.195 111.685 ;
        RECT 52.625 111.515 52.795 111.705 ;
        RECT 53.545 111.495 53.715 111.685 ;
        RECT 55.390 111.655 55.560 111.735 ;
        RECT 57.520 111.705 58.455 111.735 ;
        RECT 58.465 111.705 65.775 112.385 ;
        RECT 65.825 111.705 67.175 112.615 ;
        RECT 67.205 111.705 68.575 112.515 ;
        RECT 68.595 111.705 69.945 112.615 ;
        RECT 70.005 112.385 71.355 112.615 ;
        RECT 72.890 112.385 73.800 112.605 ;
        RECT 70.005 111.705 77.315 112.385 ;
        RECT 77.795 111.790 78.225 112.575 ;
        RECT 78.245 111.705 83.755 112.515 ;
        RECT 83.765 111.705 87.435 112.515 ;
        RECT 87.445 111.705 88.815 112.485 ;
        RECT 89.310 112.385 90.655 112.615 ;
        RECT 88.825 111.705 90.655 112.385 ;
        RECT 90.665 111.705 92.035 112.515 ;
        RECT 55.380 111.545 55.560 111.655 ;
        RECT 55.390 111.515 55.560 111.545 ;
        RECT 55.850 111.495 56.020 111.685 ;
        RECT 58.605 111.515 58.775 111.705 ;
        RECT 59.985 111.495 60.155 111.685 ;
        RECT 61.820 111.545 61.940 111.655 ;
        RECT 64.585 111.495 64.755 111.685 ;
        RECT 65.505 111.495 65.675 111.685 ;
        RECT 65.970 111.515 66.140 111.705 ;
        RECT 67.345 111.515 67.515 111.705 ;
        RECT 69.195 111.540 69.355 111.650 ;
        RECT 69.645 111.515 69.815 111.705 ;
        RECT 73.325 111.495 73.495 111.685 ;
        RECT 73.785 111.495 73.955 111.685 ;
        RECT 76.085 111.495 76.255 111.685 ;
        RECT 77.005 111.515 77.175 111.705 ;
        RECT 77.460 111.545 77.580 111.655 ;
        RECT 78.385 111.515 78.555 111.705 ;
        RECT 79.765 111.495 79.935 111.685 ;
        RECT 83.905 111.515 84.075 111.705 ;
        RECT 87.585 111.515 87.755 111.705 ;
        RECT 88.965 111.515 89.135 111.705 ;
        RECT 90.345 111.495 90.515 111.685 ;
        RECT 91.725 111.495 91.895 111.705 ;
        RECT 40.940 111.465 41.895 111.495 ;
        RECT 34.840 110.595 35.750 110.815 ;
        RECT 37.285 110.585 38.635 110.815 ;
        RECT 39.155 110.625 39.585 111.410 ;
        RECT 39.615 110.785 41.895 111.465 ;
        RECT 42.510 110.815 44.345 111.495 ;
        RECT 40.940 110.585 41.895 110.785 ;
        RECT 43.415 110.585 44.345 110.815 ;
        RECT 44.665 110.585 46.495 111.495 ;
        RECT 46.515 110.585 47.865 111.495 ;
        RECT 47.885 110.685 53.395 111.495 ;
        RECT 53.405 110.685 55.235 111.495 ;
        RECT 55.705 110.815 59.800 111.495 ;
        RECT 56.190 110.585 59.800 110.815 ;
        RECT 59.845 110.685 61.675 111.495 ;
        RECT 62.145 110.585 64.895 111.495 ;
        RECT 64.915 110.625 65.345 111.410 ;
        RECT 65.365 110.815 69.035 111.495 ;
        RECT 68.105 110.585 69.035 110.815 ;
        RECT 70.060 110.815 73.525 111.495 ;
        RECT 70.060 110.585 70.980 110.815 ;
        RECT 73.645 110.585 75.935 111.495 ;
        RECT 75.945 110.685 79.615 111.495 ;
        RECT 79.625 110.815 86.935 111.495 ;
        RECT 83.140 110.595 84.050 110.815 ;
        RECT 85.585 110.585 86.935 110.815 ;
        RECT 87.080 110.815 90.545 111.495 ;
        RECT 87.080 110.585 88.000 110.815 ;
        RECT 90.665 110.685 92.035 111.495 ;
      LAYER nwell ;
        RECT 13.190 107.465 92.230 110.295 ;
      LAYER pwell ;
        RECT 100.400 107.200 106.500 116.990 ;
        RECT 13.385 106.265 14.755 107.075 ;
        RECT 18.280 106.945 19.190 107.165 ;
        RECT 20.725 106.945 22.075 107.175 ;
        RECT 14.765 106.265 22.075 106.945 ;
        RECT 22.125 106.265 23.955 107.175 ;
        RECT 24.275 106.945 25.205 107.175 ;
        RECT 24.275 106.265 26.110 106.945 ;
        RECT 26.275 106.350 26.705 107.135 ;
        RECT 29.015 106.975 30.370 107.175 ;
        RECT 27.690 106.945 30.370 106.975 ;
        RECT 30.865 106.975 31.820 107.175 ;
        RECT 27.690 106.295 30.855 106.945 ;
        RECT 29.015 106.265 30.855 106.295 ;
        RECT 30.865 106.295 33.145 106.975 ;
        RECT 30.865 106.265 31.820 106.295 ;
        RECT 13.525 106.055 13.695 106.265 ;
        RECT 14.905 106.215 15.075 106.265 ;
        RECT 14.900 106.105 15.075 106.215 ;
        RECT 14.905 106.075 15.075 106.105 ;
        RECT 15.370 106.055 15.540 106.245 ;
        RECT 20.425 106.055 20.595 106.245 ;
        RECT 20.895 106.100 21.055 106.210 ;
        RECT 21.800 106.055 21.970 106.245 ;
        RECT 22.270 106.075 22.440 106.265 ;
        RECT 25.945 106.245 26.110 106.265 ;
        RECT 23.195 106.055 23.365 106.245 ;
        RECT 24.560 106.105 24.680 106.215 ;
        RECT 25.945 106.075 26.115 106.245 ;
        RECT 26.400 106.055 26.570 106.245 ;
        RECT 26.865 106.055 27.035 106.245 ;
        RECT 30.545 106.075 30.715 106.265 ;
        RECT 31.465 106.055 31.635 106.245 ;
        RECT 31.925 106.055 32.095 106.245 ;
        RECT 32.850 106.075 33.020 106.295 ;
        RECT 33.165 106.265 34.995 107.075 ;
        RECT 35.485 106.265 36.835 107.175 ;
        RECT 36.845 106.975 37.790 107.175 ;
        RECT 39.125 106.975 40.055 107.175 ;
        RECT 36.845 106.495 40.055 106.975 ;
        RECT 40.160 106.945 41.080 107.175 ;
        RECT 44.885 107.085 45.835 107.175 ;
        RECT 36.845 106.295 39.915 106.495 ;
        RECT 36.845 106.265 37.790 106.295 ;
        RECT 33.305 106.075 33.475 106.265 ;
        RECT 35.140 106.105 35.260 106.215 ;
        RECT 35.600 106.075 35.770 106.265 ;
        RECT 39.745 106.075 39.915 106.295 ;
        RECT 40.160 106.265 43.625 106.945 ;
        RECT 43.905 106.265 45.835 107.085 ;
        RECT 46.045 106.265 49.715 107.075 ;
        RECT 51.095 106.945 52.015 107.175 ;
        RECT 49.725 106.265 52.015 106.945 ;
        RECT 52.035 106.350 52.465 107.135 ;
        RECT 52.485 106.265 61.590 106.945 ;
        RECT 61.685 106.265 65.355 107.075 ;
        RECT 66.295 106.265 67.645 107.175 ;
        RECT 67.665 106.265 69.035 107.075 ;
        RECT 69.045 106.975 69.995 107.175 ;
        RECT 71.325 106.975 72.255 107.175 ;
        RECT 73.600 106.975 74.555 107.175 ;
        RECT 69.045 106.495 72.255 106.975 ;
        RECT 69.045 106.295 72.110 106.495 ;
        RECT 72.275 106.295 74.555 106.975 ;
        RECT 69.045 106.265 69.980 106.295 ;
        RECT 43.425 106.245 43.595 106.265 ;
        RECT 43.905 106.245 44.055 106.265 ;
        RECT 42.045 106.055 42.215 106.245 ;
        RECT 43.420 106.075 43.595 106.245 ;
        RECT 43.420 106.055 43.590 106.075 ;
        RECT 43.885 106.055 44.055 106.245 ;
        RECT 46.185 106.075 46.355 106.265 ;
        RECT 49.865 106.075 50.035 106.265 ;
        RECT 51.255 106.100 51.415 106.210 ;
        RECT 52.625 106.075 52.795 106.265 ;
        RECT 55.385 106.055 55.555 106.245 ;
        RECT 55.840 106.105 55.960 106.215 ;
        RECT 56.305 106.055 56.475 106.245 ;
        RECT 58.605 106.055 58.775 106.245 ;
        RECT 61.825 106.075 61.995 106.265 ;
        RECT 62.285 106.055 62.455 106.245 ;
        RECT 65.510 106.055 65.680 106.245 ;
        RECT 66.425 106.075 66.595 106.265 ;
        RECT 67.345 106.055 67.515 106.245 ;
        RECT 67.805 106.075 67.975 106.265 ;
        RECT 71.940 106.075 72.110 106.295 ;
        RECT 72.400 106.075 72.570 106.295 ;
        RECT 73.600 106.265 74.555 106.295 ;
        RECT 74.565 106.265 76.755 107.175 ;
        RECT 77.795 106.350 78.225 107.135 ;
        RECT 78.245 106.495 80.080 107.175 ;
        RECT 78.390 106.265 80.080 106.495 ;
        RECT 80.545 106.265 81.915 107.075 ;
        RECT 81.925 106.945 82.855 107.175 ;
        RECT 100.400 107.170 106.510 107.200 ;
        RECT 81.925 106.265 85.825 106.945 ;
        RECT 86.065 106.265 87.435 107.075 ;
        RECT 87.445 106.265 88.815 107.045 ;
        RECT 88.825 106.265 90.655 107.075 ;
        RECT 90.665 106.265 92.035 107.075 ;
        RECT 100.600 106.770 101.760 107.170 ;
        RECT 72.860 106.105 72.980 106.215 ;
        RECT 73.330 106.055 73.500 106.245 ;
        RECT 74.710 106.075 74.880 106.265 ;
        RECT 77.015 106.110 77.175 106.220 ;
        RECT 78.390 106.075 78.560 106.265 ;
        RECT 78.840 106.055 79.010 106.245 ;
        RECT 80.685 106.055 80.855 106.265 ;
        RECT 81.145 106.055 81.315 106.245 ;
        RECT 82.340 106.075 82.510 106.265 ;
        RECT 84.825 106.055 84.995 106.245 ;
        RECT 86.205 106.075 86.375 106.265 ;
        RECT 87.585 106.075 87.755 106.265 ;
        RECT 88.965 106.075 89.135 106.265 ;
        RECT 89.425 106.055 89.595 106.245 ;
        RECT 89.895 106.100 90.055 106.210 ;
        RECT 91.725 106.055 91.895 106.265 ;
        RECT 13.385 105.245 14.755 106.055 ;
        RECT 15.225 105.145 18.895 106.055 ;
        RECT 18.905 105.375 20.735 106.055 ;
        RECT 18.905 105.145 20.250 105.375 ;
        RECT 21.685 105.145 23.035 106.055 ;
        RECT 23.045 105.275 24.415 106.055 ;
        RECT 24.885 105.145 26.715 106.055 ;
        RECT 26.725 105.245 28.095 106.055 ;
        RECT 28.200 105.375 31.665 106.055 ;
        RECT 31.785 105.375 39.095 106.055 ;
        RECT 28.200 105.145 29.120 105.375 ;
        RECT 35.300 105.155 36.210 105.375 ;
        RECT 37.745 105.145 39.095 105.375 ;
        RECT 39.155 105.185 39.585 105.970 ;
        RECT 39.615 105.145 42.345 106.055 ;
        RECT 42.385 105.145 43.735 106.055 ;
        RECT 43.745 105.375 51.055 106.055 ;
        RECT 47.260 105.155 48.170 105.375 ;
        RECT 49.705 105.145 51.055 105.375 ;
        RECT 52.120 105.375 55.585 106.055 ;
        RECT 56.165 105.375 58.455 106.055 ;
        RECT 58.575 105.375 62.040 106.055 ;
        RECT 52.120 105.145 53.040 105.375 ;
        RECT 57.535 105.145 58.455 105.375 ;
        RECT 61.120 105.145 62.040 105.375 ;
        RECT 62.145 105.245 64.895 106.055 ;
        RECT 64.915 105.185 65.345 105.970 ;
        RECT 65.365 105.145 67.195 106.055 ;
        RECT 67.205 105.245 72.715 106.055 ;
        RECT 73.185 105.375 75.460 106.055 ;
        RECT 74.090 105.145 75.460 105.375 ;
        RECT 75.680 105.145 79.155 106.055 ;
        RECT 79.165 105.375 80.995 106.055 ;
        RECT 79.165 105.145 80.510 105.375 ;
        RECT 81.005 105.245 84.675 106.055 ;
        RECT 84.685 105.245 86.055 106.055 ;
        RECT 86.160 105.375 89.625 106.055 ;
        RECT 86.160 105.145 87.080 105.375 ;
        RECT 90.665 105.245 92.035 106.055 ;
        RECT 103.720 105.090 106.510 107.170 ;
      LAYER nwell ;
        RECT 13.190 102.025 92.230 104.855 ;
        RECT 101.610 102.980 106.450 105.090 ;
        RECT 107.730 104.750 117.920 117.000 ;
      LAYER pwell ;
        RECT 120.330 107.200 126.430 116.990 ;
        RECT 120.330 107.170 126.440 107.200 ;
        RECT 120.530 106.770 121.690 107.170 ;
        RECT 123.650 105.090 126.440 107.170 ;
      LAYER nwell ;
        RECT 121.540 102.980 126.380 105.090 ;
        RECT 127.660 104.750 137.850 117.000 ;
      LAYER pwell ;
        RECT 140.360 107.200 146.460 116.990 ;
        RECT 140.360 107.170 146.470 107.200 ;
        RECT 140.560 106.770 141.720 107.170 ;
        RECT 143.680 105.090 146.470 107.170 ;
      LAYER nwell ;
        RECT 141.570 102.980 146.410 105.090 ;
        RECT 147.690 104.750 157.880 117.000 ;
      LAYER pwell ;
        RECT 13.385 100.825 14.755 101.635 ;
        RECT 14.765 100.825 16.595 101.505 ;
        RECT 17.545 100.825 18.895 101.735 ;
        RECT 21.560 101.505 22.480 101.735 ;
        RECT 19.015 100.825 22.480 101.505 ;
        RECT 23.145 100.825 26.255 101.735 ;
        RECT 26.275 100.910 26.705 101.695 ;
        RECT 30.240 101.505 31.150 101.725 ;
        RECT 32.685 101.505 34.035 101.735 ;
        RECT 26.725 100.825 34.035 101.505 ;
        RECT 34.085 100.825 37.755 101.635 ;
        RECT 38.225 100.825 39.575 101.735 ;
        RECT 40.065 100.825 43.275 101.735 ;
        RECT 43.285 100.825 46.785 101.735 ;
        RECT 46.965 100.825 50.635 101.635 ;
        RECT 50.655 100.825 52.005 101.735 ;
        RECT 52.035 100.910 52.465 101.695 ;
        RECT 53.445 101.505 54.795 101.735 ;
        RECT 56.330 101.505 57.240 101.725 ;
        RECT 60.765 101.505 61.695 101.735 ;
        RECT 65.390 101.505 66.735 101.735 ;
        RECT 53.445 100.825 60.755 101.505 ;
        RECT 60.765 100.825 64.665 101.505 ;
        RECT 64.905 100.825 66.735 101.505 ;
        RECT 66.745 100.825 68.095 101.735 ;
        RECT 68.125 100.825 71.795 101.635 ;
        RECT 72.725 100.825 74.075 101.735 ;
        RECT 74.105 100.825 77.315 101.735 ;
        RECT 77.795 100.910 78.225 101.695 ;
        RECT 78.245 100.825 80.075 101.635 ;
        RECT 84.060 101.505 84.970 101.725 ;
        RECT 86.505 101.505 87.855 101.735 ;
        RECT 80.545 100.825 87.855 101.505 ;
        RECT 87.905 100.825 90.655 101.635 ;
        RECT 90.665 100.825 92.035 101.635 ;
        RECT 13.525 100.615 13.695 100.825 ;
        RECT 14.905 100.615 15.075 100.825 ;
        RECT 16.755 100.670 16.915 100.780 ;
        RECT 17.660 100.635 17.830 100.825 ;
        RECT 19.045 100.635 19.215 100.825 ;
        RECT 22.720 100.665 22.840 100.775 ;
        RECT 23.185 100.635 23.355 100.825 ;
        RECT 25.485 100.615 25.655 100.805 ;
        RECT 25.940 100.615 26.110 100.805 ;
        RECT 26.865 100.635 27.035 100.825 ;
        RECT 27.325 100.615 27.495 100.805 ;
        RECT 32.845 100.615 33.015 100.805 ;
        RECT 34.225 100.635 34.395 100.825 ;
        RECT 37.900 100.665 38.020 100.775 ;
        RECT 38.375 100.660 38.535 100.770 ;
        RECT 39.290 100.635 39.460 100.825 ;
        RECT 39.745 100.775 39.915 100.805 ;
        RECT 39.740 100.665 39.915 100.775 ;
        RECT 39.745 100.615 39.915 100.665 ;
        RECT 40.195 100.635 40.365 100.825 ;
        RECT 46.650 100.805 46.785 100.825 ;
        RECT 42.500 100.665 42.620 100.775 ;
        RECT 43.240 100.615 43.410 100.805 ;
        RECT 46.650 100.635 46.820 100.805 ;
        RECT 47.105 100.615 47.275 100.825 ;
        RECT 51.705 100.635 51.875 100.825 ;
        RECT 52.635 100.670 52.795 100.780 ;
        RECT 57.220 100.615 57.390 100.805 ;
        RECT 57.685 100.615 57.855 100.805 ;
        RECT 60.445 100.635 60.615 100.825 ;
        RECT 61.180 100.635 61.350 100.825 ;
        RECT 65.045 100.635 65.215 100.825 ;
        RECT 65.780 100.615 65.950 100.805 ;
        RECT 66.890 100.635 67.060 100.825 ;
        RECT 68.265 100.635 68.435 100.825 ;
        RECT 69.645 100.615 69.815 100.805 ;
        RECT 71.480 100.665 71.600 100.775 ;
        RECT 71.955 100.670 72.115 100.780 ;
        RECT 73.790 100.635 73.960 100.825 ;
        RECT 77.005 100.805 77.175 100.825 ;
        RECT 74.705 100.615 74.875 100.805 ;
        RECT 77.000 100.635 77.175 100.805 ;
        RECT 77.460 100.665 77.580 100.775 ;
        RECT 78.385 100.635 78.555 100.825 ;
        RECT 77.000 100.615 77.170 100.635 ;
        RECT 13.385 99.805 14.755 100.615 ;
        RECT 14.765 99.935 22.075 100.615 ;
        RECT 18.280 99.715 19.190 99.935 ;
        RECT 20.725 99.705 22.075 99.935 ;
        RECT 22.125 99.935 25.795 100.615 ;
        RECT 22.125 99.705 23.055 99.935 ;
        RECT 25.825 99.705 27.175 100.615 ;
        RECT 27.185 99.805 32.695 100.615 ;
        RECT 32.705 99.805 38.215 100.615 ;
        RECT 39.155 99.745 39.585 100.530 ;
        RECT 39.605 99.805 42.355 100.615 ;
        RECT 42.825 99.935 46.725 100.615 ;
        RECT 46.965 99.935 54.275 100.615 ;
        RECT 42.825 99.705 43.755 99.935 ;
        RECT 50.480 99.715 51.390 99.935 ;
        RECT 52.925 99.705 54.275 99.935 ;
        RECT 54.420 99.705 57.535 100.615 ;
        RECT 57.545 99.935 64.855 100.615 ;
        RECT 61.060 99.715 61.970 99.935 ;
        RECT 63.505 99.705 64.855 99.935 ;
        RECT 64.915 99.745 65.345 100.530 ;
        RECT 65.365 99.935 69.265 100.615 ;
        RECT 65.365 99.705 66.295 99.935 ;
        RECT 69.505 99.805 71.335 100.615 ;
        RECT 71.935 99.705 74.935 100.615 ;
        RECT 75.105 99.705 77.315 100.615 ;
        RECT 77.325 100.585 78.280 100.615 ;
        RECT 79.310 100.585 79.480 100.805 ;
        RECT 79.770 100.615 79.940 100.805 ;
        RECT 80.220 100.665 80.340 100.775 ;
        RECT 80.685 100.635 80.855 100.825 ;
        RECT 82.060 100.665 82.180 100.775 ;
        RECT 82.800 100.615 82.970 100.805 ;
        RECT 86.665 100.615 86.835 100.805 ;
        RECT 88.045 100.635 88.215 100.825 ;
        RECT 90.340 100.665 90.460 100.775 ;
        RECT 91.725 100.615 91.895 100.825 ;
        RECT 77.325 99.905 79.605 100.585 ;
        RECT 79.625 99.935 81.900 100.615 ;
        RECT 77.325 99.705 78.280 99.905 ;
        RECT 80.530 99.705 81.900 99.935 ;
        RECT 82.385 99.935 86.285 100.615 ;
        RECT 82.385 99.705 83.315 99.935 ;
        RECT 86.525 99.805 90.195 100.615 ;
        RECT 90.665 99.805 92.035 100.615 ;
      LAYER nwell ;
        RECT 13.190 96.585 92.230 99.415 ;
      LAYER pwell ;
        RECT 13.385 95.385 14.755 96.195 ;
        RECT 14.765 95.385 18.435 96.195 ;
        RECT 18.445 95.385 20.275 96.295 ;
        RECT 20.380 96.065 21.300 96.295 ;
        RECT 20.380 95.385 23.845 96.065 ;
        RECT 23.965 95.385 25.795 96.195 ;
        RECT 26.275 95.470 26.705 96.255 ;
        RECT 26.725 95.385 32.235 96.195 ;
        RECT 32.245 95.385 34.075 96.195 ;
        RECT 37.600 96.065 38.510 96.285 ;
        RECT 40.045 96.065 41.395 96.295 ;
        RECT 34.085 95.385 41.395 96.065 ;
        RECT 41.540 96.065 42.460 96.295 ;
        RECT 41.540 95.385 45.005 96.065 ;
        RECT 45.125 95.385 47.875 96.195 ;
        RECT 47.885 96.065 48.815 96.295 ;
        RECT 47.885 95.385 51.785 96.065 ;
        RECT 52.035 95.470 52.465 96.255 ;
        RECT 52.485 96.065 53.415 96.295 ;
        RECT 52.485 95.385 56.385 96.065 ;
        RECT 56.625 95.385 60.295 96.195 ;
        RECT 60.305 95.385 61.675 96.195 ;
        RECT 64.340 96.065 65.260 96.295 ;
        RECT 61.795 95.385 65.260 96.065 ;
        RECT 65.365 95.385 67.195 96.195 ;
        RECT 67.205 96.065 68.125 96.295 ;
        RECT 67.205 95.385 69.495 96.065 ;
        RECT 69.505 95.385 70.855 96.295 ;
        RECT 70.885 95.385 73.635 96.195 ;
        RECT 75.440 96.095 76.395 96.295 ;
        RECT 74.115 95.415 76.395 96.095 ;
        RECT 13.525 95.175 13.695 95.385 ;
        RECT 14.905 95.175 15.075 95.385 ;
        RECT 16.560 95.175 16.730 95.365 ;
        RECT 18.590 95.195 18.760 95.385 ;
        RECT 20.420 95.225 20.540 95.335 ;
        RECT 13.385 94.365 14.755 95.175 ;
        RECT 14.765 94.365 16.135 95.175 ;
        RECT 16.145 94.495 20.045 95.175 ;
        RECT 20.885 95.145 21.055 95.365 ;
        RECT 23.645 95.175 23.815 95.385 ;
        RECT 24.105 95.195 24.275 95.385 ;
        RECT 25.940 95.225 26.060 95.335 ;
        RECT 26.405 95.175 26.575 95.365 ;
        RECT 26.865 95.195 27.035 95.385 ;
        RECT 32.385 95.195 32.555 95.385 ;
        RECT 34.225 95.195 34.395 95.385 ;
        RECT 35.420 95.175 35.590 95.365 ;
        RECT 39.740 95.225 39.860 95.335 ;
        RECT 40.480 95.175 40.650 95.365 ;
        RECT 44.345 95.175 44.515 95.365 ;
        RECT 44.805 95.195 44.975 95.385 ;
        RECT 45.265 95.195 45.435 95.385 ;
        RECT 46.645 95.175 46.815 95.365 ;
        RECT 48.300 95.195 48.470 95.385 ;
        RECT 52.165 95.175 52.335 95.365 ;
        RECT 52.900 95.195 53.070 95.385 ;
        RECT 54.920 95.225 55.040 95.335 ;
        RECT 56.765 95.195 56.935 95.385 ;
        RECT 60.445 95.195 60.615 95.385 ;
        RECT 61.825 95.195 61.995 95.385 ;
        RECT 62.285 95.175 62.455 95.365 ;
        RECT 62.745 95.175 62.915 95.365 ;
        RECT 64.580 95.225 64.700 95.335 ;
        RECT 65.505 95.195 65.675 95.385 ;
        RECT 69.185 95.365 69.355 95.385 ;
        RECT 68.265 95.175 68.435 95.365 ;
        RECT 68.720 95.225 68.840 95.335 ;
        RECT 69.175 95.195 69.355 95.365 ;
        RECT 69.650 95.195 69.820 95.385 ;
        RECT 71.025 95.195 71.195 95.385 ;
        RECT 69.175 95.175 69.345 95.195 ;
        RECT 72.405 95.175 72.575 95.365 ;
        RECT 73.780 95.225 73.900 95.335 ;
        RECT 22.085 95.145 23.465 95.175 ;
        RECT 16.145 94.265 17.075 94.495 ;
        RECT 20.760 94.465 23.465 95.145 ;
        RECT 22.085 94.265 23.465 94.465 ;
        RECT 23.505 94.365 26.255 95.175 ;
        RECT 26.265 94.495 33.995 95.175 ;
        RECT 29.780 94.275 30.690 94.495 ;
        RECT 32.225 94.265 33.995 94.495 ;
        RECT 35.005 94.495 38.905 95.175 ;
        RECT 35.005 94.265 35.935 94.495 ;
        RECT 39.155 94.305 39.585 95.090 ;
        RECT 40.065 94.495 43.965 95.175 ;
        RECT 44.205 94.495 46.495 95.175 ;
        RECT 40.065 94.265 40.995 94.495 ;
        RECT 45.575 94.265 46.495 94.495 ;
        RECT 46.505 94.365 52.015 95.175 ;
        RECT 52.025 94.365 54.775 95.175 ;
        RECT 55.285 94.495 62.595 95.175 ;
        RECT 55.285 94.265 56.635 94.495 ;
        RECT 58.170 94.275 59.080 94.495 ;
        RECT 62.605 94.365 64.435 95.175 ;
        RECT 64.915 94.305 65.345 95.090 ;
        RECT 65.365 94.265 68.575 95.175 ;
        RECT 69.045 94.265 72.255 95.175 ;
        RECT 72.265 94.365 74.095 95.175 ;
        RECT 74.240 95.145 74.410 95.415 ;
        RECT 75.440 95.385 76.395 95.415 ;
        RECT 76.405 95.385 77.775 96.195 ;
        RECT 77.795 95.470 78.225 96.255 ;
        RECT 82.365 96.065 83.295 96.295 ;
        RECT 79.395 95.385 83.295 96.065 ;
        RECT 83.305 95.385 88.815 96.195 ;
        RECT 88.825 95.385 90.655 96.195 ;
        RECT 90.665 95.385 92.035 96.195 ;
        RECT 76.545 95.195 76.715 95.385 ;
        RECT 78.395 95.230 78.555 95.340 ;
        RECT 78.855 95.220 79.015 95.330 ;
        RECT 76.550 95.175 76.715 95.195 ;
        RECT 79.765 95.175 79.935 95.365 ;
        RECT 82.710 95.195 82.880 95.385 ;
        RECT 82.985 95.175 83.155 95.365 ;
        RECT 83.445 95.195 83.615 95.385 ;
        RECT 88.505 95.175 88.675 95.365 ;
        RECT 88.965 95.195 89.135 95.385 ;
        RECT 90.340 95.225 90.460 95.335 ;
        RECT 91.725 95.175 91.895 95.385 ;
        RECT 75.440 95.145 76.395 95.175 ;
        RECT 74.115 94.465 76.395 95.145 ;
        RECT 76.550 94.495 78.385 95.175 ;
        RECT 75.440 94.265 76.395 94.465 ;
        RECT 77.455 94.265 78.385 94.495 ;
        RECT 79.625 94.265 82.835 95.175 ;
        RECT 82.845 94.365 88.355 95.175 ;
        RECT 88.365 94.365 90.195 95.175 ;
        RECT 90.665 94.365 92.035 95.175 ;
      LAYER nwell ;
        RECT 13.190 91.145 92.230 93.975 ;
        RECT 99.800 92.735 112.970 100.575 ;
      LAYER pwell ;
        RECT 134.270 96.400 158.480 102.920 ;
        RECT 13.385 89.945 14.755 90.755 ;
        RECT 18.280 90.625 19.190 90.845 ;
        RECT 20.725 90.625 22.495 90.855 ;
        RECT 24.875 90.625 25.795 90.855 ;
        RECT 14.765 89.945 22.495 90.625 ;
        RECT 23.505 89.945 25.795 90.625 ;
        RECT 26.275 90.030 26.705 90.815 ;
        RECT 27.185 90.625 28.115 90.855 ;
        RECT 27.185 89.945 31.085 90.625 ;
        RECT 31.325 89.945 36.835 90.755 ;
        RECT 36.845 89.945 40.515 90.755 ;
        RECT 43.180 90.625 44.100 90.855 ;
        RECT 40.635 89.945 44.100 90.625 ;
        RECT 44.205 89.945 46.035 90.755 ;
        RECT 49.225 90.655 50.175 90.855 ;
        RECT 46.505 89.975 50.175 90.655 ;
        RECT 13.525 89.735 13.695 89.945 ;
        RECT 14.905 89.735 15.075 89.945 ;
        RECT 16.740 89.785 16.860 89.895 ;
        RECT 13.385 88.925 14.755 89.735 ;
        RECT 14.765 88.925 16.595 89.735 ;
        RECT 17.065 89.705 18.020 89.735 ;
        RECT 19.050 89.705 19.220 89.925 ;
        RECT 19.505 89.735 19.675 89.925 ;
        RECT 22.735 89.790 22.895 89.900 ;
        RECT 23.645 89.755 23.815 89.945 ;
        RECT 26.865 89.895 27.035 89.925 ;
        RECT 25.940 89.785 26.060 89.895 ;
        RECT 26.860 89.785 27.035 89.895 ;
        RECT 26.865 89.735 27.035 89.785 ;
        RECT 27.600 89.755 27.770 89.945 ;
        RECT 29.165 89.735 29.335 89.925 ;
        RECT 31.465 89.755 31.635 89.945 ;
        RECT 31.925 89.735 32.095 89.925 ;
        RECT 36.985 89.755 37.155 89.945 ;
        RECT 40.020 89.735 40.190 89.925 ;
        RECT 40.665 89.755 40.835 89.945 ;
        RECT 43.885 89.735 44.055 89.925 ;
        RECT 44.345 89.755 44.515 89.945 ;
        RECT 45.730 89.735 45.900 89.925 ;
        RECT 46.180 89.785 46.300 89.895 ;
        RECT 46.650 89.755 46.820 89.975 ;
        RECT 49.225 89.945 50.175 89.975 ;
        RECT 50.185 89.945 52.015 90.755 ;
        RECT 52.035 90.030 52.465 90.815 ;
        RECT 52.485 89.945 57.995 90.755 ;
        RECT 58.005 89.945 63.515 90.755 ;
        RECT 63.525 89.945 67.195 90.755 ;
        RECT 67.305 89.945 69.495 90.855 ;
        RECT 69.505 89.945 71.335 90.755 ;
        RECT 72.715 90.625 73.635 90.855 ;
        RECT 71.345 89.945 73.635 90.625 ;
        RECT 73.645 89.945 77.315 90.755 ;
        RECT 77.795 90.030 78.225 90.815 ;
        RECT 78.245 89.945 80.455 90.855 ;
        RECT 80.555 89.945 81.905 90.855 ;
        RECT 81.925 89.945 85.595 90.755 ;
        RECT 85.605 89.945 86.975 90.755 ;
        RECT 87.080 90.625 88.000 90.855 ;
        RECT 87.080 89.945 90.545 90.625 ;
        RECT 90.665 89.945 92.035 90.755 ;
        RECT 50.325 89.755 50.495 89.945 ;
        RECT 17.065 89.025 19.345 89.705 ;
        RECT 19.365 89.055 26.675 89.735 ;
        RECT 26.725 89.055 29.015 89.735 ;
        RECT 17.065 88.825 18.020 89.025 ;
        RECT 22.880 88.835 23.790 89.055 ;
        RECT 25.325 88.825 26.675 89.055 ;
        RECT 28.095 88.825 29.015 89.055 ;
        RECT 29.025 88.925 31.775 89.735 ;
        RECT 31.785 89.055 39.095 89.735 ;
        RECT 35.300 88.835 36.210 89.055 ;
        RECT 37.745 88.825 39.095 89.055 ;
        RECT 39.155 88.865 39.585 89.650 ;
        RECT 39.605 89.055 43.505 89.735 ;
        RECT 39.605 88.825 40.535 89.055 ;
        RECT 43.745 88.925 45.575 89.735 ;
        RECT 45.585 88.825 49.060 89.735 ;
        RECT 49.265 89.705 50.200 89.735 ;
        RECT 52.160 89.705 52.330 89.925 ;
        RECT 52.625 89.755 52.795 89.945 ;
        RECT 54.925 89.735 55.095 89.925 ;
        RECT 55.385 89.735 55.555 89.925 ;
        RECT 57.225 89.735 57.395 89.925 ;
        RECT 58.145 89.755 58.315 89.945 ;
        RECT 63.665 89.755 63.835 89.945 ;
        RECT 64.580 89.785 64.700 89.895 ;
        RECT 65.510 89.735 65.680 89.925 ;
        RECT 69.180 89.890 69.350 89.945 ;
        RECT 69.180 89.780 69.355 89.890 ;
        RECT 69.180 89.755 69.350 89.780 ;
        RECT 69.645 89.755 69.815 89.945 ;
        RECT 70.105 89.735 70.275 89.925 ;
        RECT 71.485 89.755 71.655 89.945 ;
        RECT 72.870 89.735 73.040 89.925 ;
        RECT 73.785 89.755 73.955 89.945 ;
        RECT 74.705 89.735 74.875 89.925 ;
        RECT 77.460 89.785 77.580 89.895 ;
        RECT 77.925 89.735 78.095 89.925 ;
        RECT 78.390 89.755 78.560 89.945 ;
        RECT 81.140 89.785 81.260 89.895 ;
        RECT 81.605 89.735 81.775 89.945 ;
        RECT 82.065 89.755 82.235 89.945 ;
        RECT 85.745 89.755 85.915 89.945 ;
        RECT 88.965 89.735 89.135 89.925 ;
        RECT 90.345 89.755 90.515 89.945 ;
        RECT 91.725 89.735 91.895 89.945 ;
        RECT 49.265 89.505 52.330 89.705 ;
        RECT 49.265 89.025 52.475 89.505 ;
        RECT 49.265 88.825 50.215 89.025 ;
        RECT 51.545 88.825 52.475 89.025 ;
        RECT 52.485 89.055 55.235 89.735 ;
        RECT 52.485 88.825 53.415 89.055 ;
        RECT 55.245 88.925 57.075 89.735 ;
        RECT 57.085 89.055 64.395 89.735 ;
        RECT 60.600 88.835 61.510 89.055 ;
        RECT 63.045 88.825 64.395 89.055 ;
        RECT 64.915 88.865 65.345 89.650 ;
        RECT 65.365 88.825 69.035 89.735 ;
        RECT 69.965 89.055 72.715 89.735 ;
        RECT 71.785 88.825 72.715 89.055 ;
        RECT 72.725 88.825 74.555 89.735 ;
        RECT 74.565 88.925 77.315 89.735 ;
        RECT 77.785 88.825 80.995 89.735 ;
        RECT 81.465 89.055 88.775 89.735 ;
        RECT 88.825 89.055 90.655 89.735 ;
        RECT 84.980 88.835 85.890 89.055 ;
        RECT 87.425 88.825 88.775 89.055 ;
        RECT 89.310 88.825 90.655 89.055 ;
        RECT 90.665 88.925 92.035 89.735 ;
      LAYER nwell ;
        RECT 13.190 85.705 92.230 88.535 ;
      LAYER pwell ;
        RECT 99.810 88.235 112.980 92.025 ;
        RECT 13.385 84.505 14.755 85.315 ;
        RECT 14.765 84.505 18.435 85.315 ;
        RECT 18.445 84.505 19.815 85.315 ;
        RECT 20.875 85.185 21.805 85.415 ;
        RECT 19.970 84.505 21.805 85.185 ;
        RECT 22.325 85.325 23.275 85.415 ;
        RECT 22.325 84.505 24.255 85.325 ;
        RECT 24.895 84.505 26.245 85.415 ;
        RECT 26.275 84.590 26.705 85.375 ;
        RECT 31.160 85.185 32.070 85.405 ;
        RECT 33.605 85.185 35.375 85.415 ;
        RECT 27.645 84.505 35.375 85.185 ;
        RECT 35.465 84.505 39.135 85.315 ;
        RECT 40.160 85.185 41.080 85.415 ;
        RECT 43.745 85.215 44.675 85.415 ;
        RECT 46.005 85.215 46.955 85.415 ;
        RECT 40.160 84.505 43.625 85.185 ;
        RECT 43.745 84.735 46.955 85.215 ;
        RECT 43.890 84.535 46.955 84.735 ;
        RECT 13.525 84.295 13.695 84.505 ;
        RECT 14.905 84.295 15.075 84.505 ;
        RECT 18.585 84.315 18.755 84.505 ;
        RECT 19.970 84.485 20.135 84.505 ;
        RECT 24.105 84.485 24.255 84.505 ;
        RECT 19.965 84.315 20.135 84.485 ;
        RECT 20.425 84.295 20.595 84.485 ;
        RECT 24.105 84.315 24.275 84.485 ;
        RECT 24.560 84.345 24.680 84.455 ;
        RECT 25.025 84.315 25.195 84.505 ;
        RECT 25.945 84.295 26.115 84.485 ;
        RECT 26.875 84.350 27.035 84.460 ;
        RECT 27.785 84.455 27.955 84.505 ;
        RECT 27.780 84.345 27.955 84.455 ;
        RECT 27.785 84.315 27.955 84.345 ;
        RECT 28.520 84.295 28.690 84.485 ;
        RECT 32.385 84.295 32.555 84.485 ;
        RECT 35.605 84.315 35.775 84.505 ;
        RECT 37.905 84.295 38.075 84.485 ;
        RECT 39.295 84.350 39.455 84.460 ;
        RECT 39.745 84.295 39.915 84.485 ;
        RECT 43.425 84.315 43.595 84.505 ;
        RECT 43.890 84.315 44.060 84.535 ;
        RECT 46.020 84.505 46.955 84.535 ;
        RECT 47.885 85.185 48.815 85.415 ;
        RECT 47.885 84.505 50.635 85.185 ;
        RECT 50.645 84.505 52.015 85.315 ;
        RECT 52.035 84.590 52.465 85.375 ;
        RECT 52.485 85.185 53.415 85.415 ;
        RECT 60.600 85.185 61.510 85.405 ;
        RECT 63.045 85.185 64.395 85.415 ;
        RECT 52.485 84.505 56.385 85.185 ;
        RECT 57.085 84.505 64.395 85.185 ;
        RECT 64.445 84.505 67.655 85.415 ;
        RECT 67.975 85.185 68.905 85.415 ;
        RECT 67.975 84.505 69.810 85.185 ;
        RECT 69.965 84.505 71.315 85.415 ;
        RECT 71.345 84.505 72.715 85.315 ;
        RECT 72.725 84.505 74.555 85.415 ;
        RECT 76.535 85.185 77.465 85.415 ;
        RECT 75.630 84.505 77.465 85.185 ;
        RECT 77.795 84.590 78.225 85.375 ;
        RECT 78.395 84.505 82.050 85.415 ;
        RECT 83.305 85.185 84.235 85.415 ;
        RECT 83.305 84.505 87.205 85.185 ;
        RECT 87.445 84.505 88.815 85.285 ;
        RECT 88.825 84.505 90.655 85.315 ;
        RECT 90.665 84.505 92.035 85.315 ;
        RECT 47.115 84.350 47.275 84.460 ;
        RECT 13.385 83.485 14.755 84.295 ;
        RECT 14.765 83.485 20.275 84.295 ;
        RECT 20.285 83.485 25.795 84.295 ;
        RECT 25.805 83.485 27.635 84.295 ;
        RECT 28.105 83.615 32.005 84.295 ;
        RECT 28.105 83.385 29.035 83.615 ;
        RECT 32.245 83.485 37.755 84.295 ;
        RECT 37.765 83.485 39.135 84.295 ;
        RECT 39.155 83.425 39.585 84.210 ;
        RECT 39.605 83.615 46.915 84.295 ;
        RECT 43.120 83.395 44.030 83.615 ;
        RECT 45.565 83.385 46.915 83.615 ;
        RECT 46.965 84.265 47.910 84.295 ;
        RECT 49.400 84.265 49.570 84.485 ;
        RECT 49.860 84.345 49.980 84.455 ;
        RECT 50.325 84.295 50.495 84.505 ;
        RECT 50.785 84.315 50.955 84.505 ;
        RECT 52.900 84.315 53.070 84.505 ;
        RECT 56.760 84.345 56.880 84.455 ;
        RECT 57.225 84.315 57.395 84.505 ;
        RECT 60.905 84.295 61.075 84.485 ;
        RECT 61.365 84.295 61.535 84.485 ;
        RECT 64.575 84.315 64.745 84.505 ;
        RECT 69.645 84.485 69.810 84.505 ;
        RECT 65.515 84.340 65.675 84.450 ;
        RECT 46.965 83.585 49.715 84.265 ;
        RECT 50.185 83.615 57.495 84.295 ;
        RECT 46.965 83.385 47.910 83.585 ;
        RECT 53.700 83.395 54.610 83.615 ;
        RECT 56.145 83.385 57.495 83.615 ;
        RECT 57.640 83.615 61.105 84.295 ;
        RECT 57.640 83.385 58.560 83.615 ;
        RECT 61.225 83.485 64.895 84.295 ;
        RECT 66.430 84.265 66.600 84.485 ;
        RECT 69.645 84.315 69.815 84.485 ;
        RECT 71.030 84.315 71.200 84.505 ;
        RECT 71.485 84.315 71.655 84.505 ;
        RECT 71.945 84.295 72.115 84.485 ;
        RECT 72.405 84.295 72.575 84.485 ;
        RECT 72.870 84.315 73.040 84.505 ;
        RECT 75.630 84.485 75.795 84.505 ;
        RECT 78.395 84.485 78.555 84.505 ;
        RECT 74.715 84.350 74.875 84.460 ;
        RECT 75.625 84.315 75.795 84.485 ;
        RECT 77.005 84.295 77.175 84.485 ;
        RECT 77.465 84.295 77.635 84.485 ;
        RECT 78.385 84.315 78.555 84.485 ;
        RECT 82.535 84.350 82.695 84.460 ;
        RECT 82.985 84.295 83.155 84.485 ;
        RECT 83.720 84.315 83.890 84.505 ;
        RECT 85.745 84.295 85.915 84.485 ;
        RECT 87.585 84.315 87.755 84.505 ;
        RECT 88.965 84.315 89.135 84.505 ;
        RECT 90.345 84.295 90.515 84.485 ;
        RECT 91.725 84.295 91.895 84.505 ;
        RECT 68.560 84.265 69.495 84.295 ;
        RECT 64.915 83.425 65.345 84.210 ;
        RECT 66.430 84.065 69.495 84.265 ;
        RECT 66.285 83.585 69.495 84.065 ;
        RECT 66.285 83.385 67.215 83.585 ;
        RECT 68.545 83.385 69.495 83.585 ;
        RECT 69.505 83.615 72.255 84.295 ;
        RECT 69.505 83.385 70.435 83.615 ;
        RECT 72.265 83.485 75.015 84.295 ;
        RECT 75.025 83.615 77.315 84.295 ;
        RECT 75.025 83.385 75.945 83.615 ;
        RECT 77.325 83.485 82.835 84.295 ;
        RECT 82.845 83.485 85.595 84.295 ;
        RECT 85.605 83.515 86.975 84.295 ;
        RECT 87.080 83.615 90.545 84.295 ;
        RECT 87.080 83.385 88.000 83.615 ;
        RECT 90.665 83.485 92.035 84.295 ;
      LAYER nwell ;
        RECT 13.190 80.265 92.230 83.095 ;
      LAYER pwell ;
        RECT 99.810 80.745 113.660 87.965 ;
      LAYER nwell ;
        RECT 117.410 82.420 129.660 92.610 ;
      LAYER pwell ;
        RECT 127.210 81.190 129.320 81.200 ;
        RECT 17.265 79.885 18.215 79.975 ;
        RECT 13.385 79.065 14.755 79.875 ;
        RECT 14.765 79.065 16.595 79.875 ;
        RECT 17.265 79.065 19.195 79.885 ;
        RECT 19.365 79.065 20.715 79.975 ;
        RECT 20.745 79.065 22.095 79.975 ;
        RECT 23.045 79.775 23.975 79.975 ;
        RECT 25.310 79.775 26.255 79.975 ;
        RECT 23.045 79.295 26.255 79.775 ;
        RECT 23.185 79.095 26.255 79.295 ;
        RECT 26.275 79.150 26.705 79.935 ;
        RECT 13.525 78.855 13.695 79.065 ;
        RECT 14.905 78.875 15.075 79.065 ;
        RECT 19.045 79.045 19.195 79.065 ;
        RECT 15.825 78.855 15.995 79.045 ;
        RECT 16.740 78.905 16.860 79.015 ;
        RECT 19.045 78.875 19.215 79.045 ;
        RECT 20.430 78.875 20.600 79.065 ;
        RECT 20.890 78.875 21.060 79.065 ;
        RECT 22.275 78.910 22.435 79.020 ;
        RECT 23.185 78.855 23.355 79.095 ;
        RECT 25.310 79.065 26.255 79.095 ;
        RECT 26.725 79.065 28.095 79.875 ;
        RECT 28.105 79.745 29.035 79.975 ;
        RECT 28.105 79.065 32.005 79.745 ;
        RECT 32.245 79.065 37.755 79.875 ;
        RECT 41.885 79.745 42.815 79.975 ;
        RECT 38.915 79.065 42.815 79.745 ;
        RECT 42.825 79.065 44.655 79.875 ;
        RECT 44.760 79.745 45.680 79.975 ;
        RECT 51.000 79.745 51.920 79.975 ;
        RECT 44.760 79.065 48.225 79.745 ;
        RECT 48.455 79.065 51.920 79.745 ;
        RECT 52.035 79.150 52.465 79.935 ;
        RECT 52.485 79.745 53.405 79.975 ;
        RECT 54.785 79.745 55.715 79.975 ;
        RECT 52.485 79.065 54.775 79.745 ;
        RECT 54.785 79.065 58.685 79.745 ;
        RECT 58.925 79.065 64.435 79.875 ;
        RECT 67.100 79.745 68.020 79.975 ;
        RECT 69.495 79.745 70.415 79.975 ;
        RECT 64.555 79.065 68.020 79.745 ;
        RECT 68.125 79.065 70.415 79.745 ;
        RECT 70.425 79.065 73.175 79.875 ;
        RECT 73.795 79.065 77.450 79.975 ;
        RECT 77.795 79.150 78.225 79.935 ;
        RECT 78.245 79.065 81.455 79.975 ;
        RECT 84.980 79.745 85.890 79.965 ;
        RECT 87.425 79.745 88.775 79.975 ;
        RECT 89.310 79.745 90.655 79.975 ;
        RECT 81.465 79.065 88.775 79.745 ;
        RECT 88.825 79.065 90.655 79.745 ;
        RECT 90.665 79.065 92.035 79.875 ;
        RECT 13.385 78.045 14.755 78.855 ;
        RECT 15.685 78.175 22.995 78.855 ;
        RECT 19.200 77.955 20.110 78.175 ;
        RECT 21.645 77.945 22.995 78.175 ;
        RECT 23.045 78.045 24.875 78.855 ;
        RECT 25.025 78.825 25.195 79.045 ;
        RECT 26.865 78.875 27.035 79.065 ;
        RECT 28.240 78.905 28.360 79.015 ;
        RECT 28.520 78.875 28.690 79.065 ;
        RECT 28.705 78.855 28.875 79.045 ;
        RECT 32.385 78.875 32.555 79.065 ;
        RECT 36.525 78.855 36.695 79.045 ;
        RECT 37.915 78.910 38.075 79.020 ;
        RECT 39.745 78.855 39.915 79.045 ;
        RECT 42.230 78.875 42.400 79.065 ;
        RECT 42.965 78.875 43.135 79.065 ;
        RECT 47.100 78.905 47.220 79.015 ;
        RECT 48.025 78.875 48.195 79.065 ;
        RECT 48.485 78.875 48.655 79.065 ;
        RECT 54.465 78.855 54.635 79.065 ;
        RECT 54.925 78.855 55.095 79.045 ;
        RECT 55.200 78.875 55.370 79.065 ;
        RECT 59.065 78.875 59.235 79.065 ;
        RECT 64.585 78.855 64.755 79.065 ;
        RECT 65.505 78.855 65.675 79.045 ;
        RECT 68.265 78.875 68.435 79.065 ;
        RECT 68.730 78.855 68.900 79.045 ;
        RECT 70.565 78.875 70.735 79.065 ;
        RECT 73.795 79.045 73.955 79.065 ;
        RECT 71.955 78.900 72.115 79.010 ;
        RECT 73.320 78.905 73.440 79.015 ;
        RECT 73.785 78.875 73.955 79.045 ;
        RECT 75.165 78.855 75.335 79.045 ;
        RECT 77.925 78.855 78.095 79.045 ;
        RECT 78.385 78.855 78.555 79.065 ;
        RECT 81.605 78.875 81.775 79.065 ;
        RECT 82.065 78.855 82.235 79.045 ;
        RECT 83.720 78.855 83.890 79.045 ;
        RECT 87.585 78.855 87.755 79.045 ;
        RECT 88.965 78.855 89.135 79.065 ;
        RECT 91.725 78.855 91.895 79.065 ;
        RECT 27.150 78.825 28.095 78.855 ;
        RECT 25.025 78.625 28.095 78.825 ;
        RECT 24.885 78.145 28.095 78.625 ;
        RECT 28.565 78.175 36.295 78.855 ;
        RECT 24.885 77.945 25.815 78.145 ;
        RECT 27.150 77.945 28.095 78.145 ;
        RECT 32.080 77.955 32.990 78.175 ;
        RECT 34.525 77.945 36.295 78.175 ;
        RECT 36.385 78.045 39.135 78.855 ;
        RECT 39.155 77.985 39.585 78.770 ;
        RECT 39.605 78.175 46.915 78.855 ;
        RECT 43.120 77.955 44.030 78.175 ;
        RECT 45.565 77.945 46.915 78.175 ;
        RECT 47.465 78.175 54.775 78.855 ;
        RECT 47.465 77.945 48.815 78.175 ;
        RECT 50.350 77.955 51.260 78.175 ;
        RECT 54.785 78.045 57.535 78.855 ;
        RECT 57.585 78.175 64.895 78.855 ;
        RECT 57.585 77.945 58.935 78.175 ;
        RECT 60.470 77.955 61.380 78.175 ;
        RECT 64.915 77.985 65.345 78.770 ;
        RECT 65.445 77.945 68.445 78.855 ;
        RECT 68.585 77.945 71.505 78.855 ;
        RECT 72.735 77.945 75.465 78.855 ;
        RECT 75.495 77.945 78.225 78.855 ;
        RECT 78.245 78.045 81.915 78.855 ;
        RECT 81.925 78.045 83.295 78.855 ;
        RECT 83.305 78.175 87.205 78.855 ;
        RECT 83.305 77.945 84.235 78.175 ;
        RECT 87.445 78.075 88.815 78.855 ;
        RECT 88.825 78.045 90.655 78.855 ;
        RECT 90.665 78.045 92.035 78.855 ;
      LAYER nwell ;
        RECT 13.190 74.825 92.230 77.655 ;
      LAYER pwell ;
        RECT 99.810 74.755 110.700 80.745 ;
        RECT 117.420 78.410 129.320 81.190 ;
        RECT 117.420 76.450 127.240 78.410 ;
        RECT 117.420 75.290 127.640 76.450 ;
      LAYER nwell ;
        RECT 129.320 76.300 131.430 81.140 ;
        RECT 134.240 78.800 139.890 84.990 ;
      LAYER pwell ;
        RECT 134.230 75.340 139.880 78.440 ;
        RECT 117.420 75.090 127.240 75.290 ;
        RECT 13.385 73.625 14.755 74.435 ;
        RECT 14.765 73.625 16.595 74.435 ;
        RECT 16.915 74.305 17.845 74.535 ;
        RECT 19.365 74.335 20.295 74.535 ;
        RECT 21.625 74.335 22.575 74.535 ;
        RECT 16.915 73.625 18.750 74.305 ;
        RECT 19.365 73.855 22.575 74.335 ;
        RECT 23.045 74.335 23.975 74.535 ;
        RECT 25.310 74.335 26.255 74.535 ;
        RECT 23.045 73.855 26.255 74.335 ;
        RECT 13.525 73.415 13.695 73.625 ;
        RECT 14.905 73.575 15.075 73.625 ;
        RECT 18.585 73.605 18.750 73.625 ;
        RECT 19.510 73.655 22.575 73.855 ;
        RECT 14.900 73.465 15.075 73.575 ;
        RECT 14.905 73.435 15.075 73.465 ;
        RECT 15.640 73.415 15.810 73.605 ;
        RECT 18.585 73.435 18.755 73.605 ;
        RECT 19.040 73.465 19.160 73.575 ;
        RECT 19.510 73.435 19.680 73.655 ;
        RECT 21.640 73.625 22.575 73.655 ;
        RECT 23.185 73.655 26.255 73.855 ;
        RECT 26.275 73.710 26.705 74.495 ;
        RECT 19.780 73.415 19.950 73.605 ;
        RECT 22.720 73.465 22.840 73.575 ;
        RECT 23.185 73.435 23.355 73.655 ;
        RECT 25.310 73.625 26.255 73.655 ;
        RECT 26.725 73.625 28.555 74.435 ;
        RECT 32.540 74.305 33.450 74.525 ;
        RECT 34.985 74.305 36.755 74.535 ;
        RECT 29.025 73.625 36.755 74.305 ;
        RECT 36.845 73.625 40.515 74.435 ;
        RECT 42.365 74.305 43.295 74.535 ;
        RECT 46.505 74.305 47.435 74.535 ;
        RECT 40.990 73.625 42.355 74.305 ;
        RECT 42.365 73.625 46.265 74.305 ;
        RECT 46.505 73.625 50.405 74.305 ;
        RECT 50.645 73.625 52.015 74.435 ;
        RECT 52.035 73.710 52.465 74.495 ;
        RECT 52.485 74.305 53.415 74.535 ;
        RECT 57.125 74.305 58.475 74.535 ;
        RECT 60.010 74.305 60.920 74.525 ;
        RECT 67.100 74.305 68.020 74.535 ;
        RECT 52.485 73.625 56.385 74.305 ;
        RECT 57.125 73.625 64.435 74.305 ;
        RECT 64.555 73.625 68.020 74.305 ;
        RECT 68.125 73.625 71.335 74.535 ;
        RECT 72.485 74.445 73.435 74.535 ;
        RECT 71.505 73.625 73.435 74.445 ;
        RECT 73.645 73.625 74.995 74.535 ;
        RECT 75.970 74.305 77.315 74.535 ;
        RECT 75.485 73.625 77.315 74.305 ;
        RECT 77.795 73.710 78.225 74.495 ;
        RECT 78.245 73.625 80.995 74.435 ;
        RECT 84.980 74.305 85.890 74.525 ;
        RECT 87.425 74.305 88.775 74.535 ;
        RECT 89.310 74.305 90.655 74.535 ;
        RECT 81.465 73.625 88.775 74.305 ;
        RECT 88.825 73.625 90.655 74.305 ;
        RECT 90.665 73.625 92.035 74.435 ;
        RECT 23.655 73.460 23.815 73.570 ;
        RECT 26.865 73.435 27.035 73.625 ;
        RECT 27.970 73.415 28.140 73.605 ;
        RECT 28.705 73.575 28.875 73.605 ;
        RECT 28.700 73.465 28.875 73.575 ;
        RECT 28.705 73.415 28.875 73.465 ;
        RECT 29.165 73.435 29.335 73.625 ;
        RECT 33.765 73.415 33.935 73.605 ;
        RECT 36.985 73.435 37.155 73.625 ;
        RECT 39.755 73.460 39.915 73.570 ;
        RECT 40.665 73.415 40.835 73.605 ;
        RECT 42.780 73.435 42.950 73.625 ;
        RECT 45.725 73.415 45.895 73.605 ;
        RECT 46.920 73.435 47.090 73.625 ;
        RECT 48.485 73.415 48.655 73.605 ;
        RECT 50.785 73.435 50.955 73.625 ;
        RECT 52.900 73.435 53.070 73.625 ;
        RECT 56.120 73.415 56.290 73.605 ;
        RECT 56.760 73.465 56.880 73.575 ;
        RECT 63.205 73.415 63.375 73.605 ;
        RECT 63.665 73.415 63.835 73.605 ;
        RECT 64.125 73.435 64.295 73.625 ;
        RECT 64.585 73.435 64.755 73.625 ;
        RECT 65.505 73.435 65.675 73.605 ;
        RECT 68.265 73.435 68.435 73.625 ;
        RECT 71.505 73.605 71.655 73.625 ;
        RECT 69.650 73.415 69.820 73.605 ;
        RECT 71.030 73.415 71.200 73.605 ;
        RECT 71.485 73.435 71.655 73.605 ;
        RECT 72.400 73.415 72.570 73.605 ;
        RECT 72.875 73.460 73.035 73.570 ;
        RECT 73.785 73.415 73.955 73.605 ;
        RECT 74.710 73.435 74.880 73.625 ;
        RECT 75.160 73.465 75.280 73.575 ;
        RECT 75.625 73.435 75.795 73.625 ;
        RECT 77.460 73.465 77.580 73.575 ;
        RECT 78.385 73.435 78.555 73.625 ;
        RECT 80.220 73.415 80.390 73.605 ;
        RECT 80.685 73.415 80.855 73.605 ;
        RECT 81.140 73.465 81.260 73.575 ;
        RECT 81.605 73.435 81.775 73.625 ;
        RECT 82.520 73.465 82.640 73.575 ;
        RECT 83.260 73.415 83.430 73.605 ;
        RECT 88.965 73.435 89.135 73.625 ;
        RECT 90.345 73.415 90.515 73.605 ;
        RECT 91.725 73.415 91.895 73.625 ;
        RECT 13.385 72.605 14.755 73.415 ;
        RECT 15.225 72.735 19.125 73.415 ;
        RECT 19.365 72.735 23.265 73.415 ;
        RECT 24.655 72.735 28.555 73.415 ;
        RECT 28.565 72.735 33.380 73.415 ;
        RECT 15.225 72.505 16.155 72.735 ;
        RECT 19.365 72.505 20.295 72.735 ;
        RECT 27.625 72.505 28.555 72.735 ;
        RECT 33.625 72.605 39.135 73.415 ;
        RECT 39.155 72.545 39.585 73.330 ;
        RECT 40.525 72.735 45.340 73.415 ;
        RECT 45.585 72.605 48.335 73.415 ;
        RECT 48.345 72.735 55.655 73.415 ;
        RECT 51.860 72.515 52.770 72.735 ;
        RECT 54.305 72.505 55.655 72.735 ;
        RECT 55.705 72.735 59.605 73.415 ;
        RECT 59.940 72.735 63.405 73.415 ;
        RECT 55.705 72.505 56.635 72.735 ;
        RECT 59.940 72.505 60.860 72.735 ;
        RECT 63.525 72.605 64.895 73.415 ;
        RECT 64.915 72.545 65.345 73.330 ;
        RECT 65.770 72.735 68.195 73.415 ;
        RECT 68.585 72.505 69.935 73.415 ;
        RECT 69.965 72.505 71.315 73.415 ;
        RECT 71.365 72.505 72.715 73.415 ;
        RECT 73.645 72.505 76.855 73.415 ;
        RECT 77.060 72.505 80.535 73.415 ;
        RECT 80.545 72.605 82.375 73.415 ;
        RECT 82.845 72.735 86.745 73.415 ;
        RECT 87.080 72.735 90.545 73.415 ;
        RECT 82.845 72.505 83.775 72.735 ;
        RECT 87.080 72.505 88.000 72.735 ;
        RECT 90.665 72.605 92.035 73.415 ;
      LAYER nwell ;
        RECT 13.190 69.385 92.230 72.215 ;
      LAYER pwell ;
        RECT 13.385 68.185 14.755 68.995 ;
        RECT 18.280 68.865 19.190 69.085 ;
        RECT 20.725 68.865 22.495 69.095 ;
        RECT 14.765 68.185 22.495 68.865 ;
        RECT 22.585 68.185 26.255 68.995 ;
        RECT 26.275 68.270 26.705 69.055 ;
        RECT 30.240 68.865 31.150 69.085 ;
        RECT 32.685 68.865 34.455 69.095 ;
        RECT 26.725 68.185 34.455 68.865 ;
        RECT 34.545 68.185 36.375 68.995 ;
        RECT 36.385 68.865 37.315 69.095 ;
        RECT 44.040 68.865 44.950 69.085 ;
        RECT 46.485 68.865 47.835 69.095 ;
        RECT 36.385 68.185 40.285 68.865 ;
        RECT 40.525 68.185 47.835 68.865 ;
        RECT 47.885 68.865 48.815 69.095 ;
        RECT 47.885 68.185 51.785 68.865 ;
        RECT 52.035 68.270 52.465 69.055 ;
        RECT 52.580 68.865 53.500 69.095 ;
        RECT 52.580 68.185 56.045 68.865 ;
        RECT 56.165 68.185 59.835 68.995 ;
        RECT 68.480 68.865 69.400 69.095 ;
        RECT 60.765 68.185 65.580 68.865 ;
        RECT 65.935 68.185 69.400 68.865 ;
        RECT 69.705 69.005 70.655 69.095 ;
        RECT 69.705 68.185 71.635 69.005 ;
        RECT 71.815 68.185 73.165 69.095 ;
        RECT 73.205 68.185 74.555 69.095 ;
        RECT 75.900 68.895 76.855 69.095 ;
        RECT 74.575 68.215 76.855 68.895 ;
        RECT 77.795 68.270 78.225 69.055 ;
        RECT 13.525 67.975 13.695 68.185 ;
        RECT 14.905 67.995 15.075 68.185 ;
        RECT 16.285 67.975 16.455 68.165 ;
        RECT 16.755 68.020 16.915 68.130 ;
        RECT 17.665 67.975 17.835 68.165 ;
        RECT 22.725 67.995 22.895 68.185 ;
        RECT 26.865 67.995 27.035 68.185 ;
        RECT 28.890 67.975 29.060 68.165 ;
        RECT 29.625 67.975 29.795 68.165 ;
        RECT 34.685 67.995 34.855 68.185 ;
        RECT 35.145 67.975 35.315 68.165 ;
        RECT 36.800 67.995 36.970 68.185 ;
        RECT 38.820 68.025 38.940 68.135 ;
        RECT 39.740 68.025 39.860 68.135 ;
        RECT 40.665 67.995 40.835 68.185 ;
        RECT 43.425 67.975 43.595 68.165 ;
        RECT 46.655 67.975 46.825 68.165 ;
        RECT 47.105 67.975 47.275 68.165 ;
        RECT 48.300 67.995 48.470 68.185 ;
        RECT 51.705 67.975 51.875 68.165 ;
        RECT 52.175 68.020 52.335 68.130 ;
        RECT 53.360 67.975 53.530 68.165 ;
        RECT 55.845 67.995 56.015 68.185 ;
        RECT 56.305 67.995 56.475 68.185 ;
        RECT 59.995 68.030 60.155 68.140 ;
        RECT 60.905 67.995 61.075 68.185 ;
        RECT 64.125 67.975 64.295 68.165 ;
        RECT 64.580 68.025 64.700 68.135 ;
        RECT 65.780 67.975 65.950 68.165 ;
        RECT 65.965 67.995 66.135 68.185 ;
        RECT 71.485 68.165 71.635 68.185 ;
        RECT 72.865 68.165 73.035 68.185 ;
        RECT 69.645 67.975 69.815 68.165 ;
        RECT 71.485 67.995 71.655 68.165 ;
        RECT 72.400 68.025 72.520 68.135 ;
        RECT 72.860 67.995 73.035 68.165 ;
        RECT 73.320 67.995 73.490 68.185 ;
        RECT 74.700 67.995 74.870 68.215 ;
        RECT 75.900 68.185 76.855 68.215 ;
        RECT 79.165 68.185 82.375 69.095 ;
        RECT 82.385 68.185 85.135 68.995 ;
        RECT 85.145 68.865 86.490 69.095 ;
        RECT 87.080 68.865 88.000 69.095 ;
        RECT 85.145 68.185 86.975 68.865 ;
        RECT 87.080 68.185 90.545 68.865 ;
        RECT 90.665 68.185 92.035 68.995 ;
        RECT 78.380 68.140 78.550 68.165 ;
        RECT 77.015 68.030 77.175 68.140 ;
        RECT 78.380 68.030 78.555 68.140 ;
        RECT 13.385 67.165 14.755 67.975 ;
        RECT 14.765 67.295 16.595 67.975 ;
        RECT 17.525 67.295 25.255 67.975 ;
        RECT 25.575 67.295 29.475 67.975 ;
        RECT 14.765 67.065 16.110 67.295 ;
        RECT 21.040 67.075 21.950 67.295 ;
        RECT 23.485 67.065 25.255 67.295 ;
        RECT 28.545 67.065 29.475 67.295 ;
        RECT 29.485 67.165 34.995 67.975 ;
        RECT 35.005 67.165 38.675 67.975 ;
        RECT 39.155 67.105 39.585 67.890 ;
        RECT 40.160 67.295 43.625 67.975 ;
        RECT 40.160 67.065 41.080 67.295 ;
        RECT 43.745 67.065 46.955 67.975 ;
        RECT 46.965 67.165 48.335 67.975 ;
        RECT 48.440 67.295 51.905 67.975 ;
        RECT 52.945 67.295 56.845 67.975 ;
        RECT 57.125 67.295 64.435 67.975 ;
        RECT 48.440 67.065 49.360 67.295 ;
        RECT 52.945 67.065 53.875 67.295 ;
        RECT 57.125 67.065 58.475 67.295 ;
        RECT 60.010 67.075 60.920 67.295 ;
        RECT 64.915 67.105 65.345 67.890 ;
        RECT 65.365 67.295 69.265 67.975 ;
        RECT 65.365 67.065 66.295 67.295 ;
        RECT 69.505 67.165 72.255 67.975 ;
        RECT 72.860 67.945 73.030 67.995 ;
        RECT 78.380 67.975 78.550 68.030 ;
        RECT 78.845 67.975 79.015 68.165 ;
        RECT 79.305 67.995 79.475 68.185 ;
        RECT 82.065 67.975 82.235 68.165 ;
        RECT 82.525 67.995 82.695 68.185 ;
        RECT 86.665 67.995 86.835 68.185 ;
        RECT 90.345 67.975 90.515 68.185 ;
        RECT 91.725 67.975 91.895 68.185 ;
        RECT 74.060 67.945 75.015 67.975 ;
        RECT 72.735 67.265 75.015 67.945 ;
        RECT 74.060 67.065 75.015 67.265 ;
        RECT 75.220 67.065 78.695 67.975 ;
        RECT 78.705 67.065 81.915 67.975 ;
        RECT 81.925 67.295 89.235 67.975 ;
        RECT 85.440 67.075 86.350 67.295 ;
        RECT 87.885 67.065 89.235 67.295 ;
        RECT 89.285 67.195 90.655 67.975 ;
        RECT 90.665 67.165 92.035 67.975 ;
      LAYER nwell ;
        RECT 13.190 63.945 92.230 66.775 ;
      LAYER pwell ;
        RECT 13.385 62.745 14.755 63.555 ;
        RECT 14.765 63.425 16.110 63.655 ;
        RECT 16.605 63.425 17.950 63.655 ;
        RECT 14.765 62.745 16.595 63.425 ;
        RECT 16.605 62.745 18.435 63.425 ;
        RECT 18.445 62.745 19.815 63.555 ;
        RECT 19.825 63.425 21.170 63.655 ;
        RECT 19.825 62.745 21.655 63.425 ;
        RECT 21.665 62.745 25.335 63.555 ;
        RECT 26.275 62.830 26.705 63.615 ;
        RECT 26.725 62.745 30.200 63.655 ;
        RECT 31.455 63.425 32.385 63.655 ;
        RECT 30.550 62.745 32.385 63.425 ;
        RECT 32.705 62.745 34.535 63.555 ;
        RECT 38.060 63.425 38.970 63.645 ;
        RECT 40.505 63.425 41.855 63.655 ;
        RECT 34.545 62.745 41.855 63.425 ;
        RECT 41.905 62.745 44.655 63.555 ;
        RECT 44.665 63.425 45.595 63.655 ;
        RECT 44.665 62.745 48.565 63.425 ;
        RECT 49.275 62.745 52.015 63.425 ;
        RECT 52.035 62.830 52.465 63.615 ;
        RECT 56.000 63.425 56.910 63.645 ;
        RECT 58.445 63.425 59.795 63.655 ;
        RECT 52.485 62.745 59.795 63.425 ;
        RECT 59.940 63.425 60.860 63.655 ;
        RECT 66.180 63.425 67.100 63.655 ;
        RECT 59.940 62.745 63.405 63.425 ;
        RECT 63.635 62.745 67.100 63.425 ;
        RECT 67.205 62.745 69.035 63.655 ;
        RECT 76.535 63.425 77.465 63.655 ;
        RECT 69.965 62.745 74.780 63.425 ;
        RECT 75.630 62.745 77.465 63.425 ;
        RECT 77.795 62.830 78.225 63.615 ;
        RECT 78.245 62.745 80.075 63.555 ;
        RECT 82.740 63.425 83.660 63.655 ;
        RECT 80.195 62.745 83.660 63.425 ;
        RECT 83.765 63.425 84.695 63.655 ;
        RECT 89.310 63.425 90.655 63.655 ;
        RECT 83.765 62.745 87.665 63.425 ;
        RECT 88.825 62.745 90.655 63.425 ;
        RECT 90.665 62.745 92.035 63.555 ;
        RECT 13.525 62.535 13.695 62.745 ;
        RECT 14.905 62.535 15.075 62.725 ;
        RECT 16.285 62.555 16.455 62.745 ;
        RECT 18.125 62.555 18.295 62.745 ;
        RECT 16.290 62.535 16.455 62.555 ;
        RECT 18.585 62.535 18.755 62.745 ;
        RECT 21.345 62.555 21.515 62.745 ;
        RECT 21.805 62.555 21.975 62.745 ;
        RECT 24.130 62.555 24.300 62.725 ;
        RECT 24.130 62.535 24.240 62.555 ;
        RECT 24.565 62.535 24.735 62.725 ;
        RECT 25.495 62.590 25.655 62.700 ;
        RECT 26.870 62.555 27.040 62.745 ;
        RECT 30.550 62.725 30.715 62.745 ;
        RECT 30.545 62.555 30.715 62.725 ;
        RECT 31.925 62.535 32.095 62.725 ;
        RECT 32.845 62.555 33.015 62.745 ;
        RECT 34.685 62.555 34.855 62.745 ;
        RECT 39.745 62.535 39.915 62.725 ;
        RECT 42.045 62.555 42.215 62.745 ;
        RECT 42.505 62.535 42.675 62.725 ;
        RECT 45.080 62.555 45.250 62.745 ;
        RECT 48.940 62.585 49.060 62.695 ;
        RECT 49.865 62.535 50.035 62.725 ;
        RECT 51.705 62.555 51.875 62.745 ;
        RECT 52.625 62.555 52.795 62.745 ;
        RECT 55.110 62.535 55.280 62.725 ;
        RECT 55.845 62.535 56.015 62.725 ;
        RECT 63.205 62.555 63.375 62.745 ;
        RECT 63.665 62.555 63.835 62.745 ;
        RECT 64.585 62.535 64.755 62.725 ;
        RECT 68.265 62.535 68.435 62.725 ;
        RECT 68.720 62.555 68.890 62.745 ;
        RECT 70.105 62.725 70.275 62.745 ;
        RECT 75.630 62.725 75.795 62.745 ;
        RECT 69.195 62.590 69.355 62.700 ;
        RECT 69.650 62.535 69.820 62.725 ;
        RECT 70.105 62.555 70.280 62.725 ;
        RECT 75.160 62.585 75.280 62.695 ;
        RECT 75.625 62.555 75.795 62.725 ;
        RECT 78.385 62.555 78.555 62.745 ;
        RECT 80.225 62.555 80.395 62.745 ;
        RECT 70.110 62.535 70.280 62.555 ;
        RECT 81.140 62.535 81.310 62.725 ;
        RECT 82.535 62.580 82.695 62.690 ;
        RECT 83.720 62.535 83.890 62.725 ;
        RECT 84.180 62.555 84.350 62.745 ;
        RECT 88.055 62.590 88.215 62.700 ;
        RECT 88.505 62.535 88.675 62.725 ;
        RECT 88.965 62.535 89.135 62.745 ;
        RECT 91.725 62.535 91.895 62.745 ;
        RECT 13.385 61.725 14.755 62.535 ;
        RECT 14.765 61.725 16.135 62.535 ;
        RECT 16.290 61.855 18.125 62.535 ;
        RECT 17.195 61.625 18.125 61.855 ;
        RECT 18.445 61.725 19.815 62.535 ;
        RECT 19.825 61.855 24.240 62.535 ;
        RECT 24.425 61.855 31.735 62.535 ;
        RECT 31.785 61.855 39.095 62.535 ;
        RECT 19.825 61.625 23.755 61.855 ;
        RECT 27.940 61.635 28.850 61.855 ;
        RECT 30.385 61.625 31.735 61.855 ;
        RECT 35.300 61.635 36.210 61.855 ;
        RECT 37.745 61.625 39.095 61.855 ;
        RECT 39.155 61.665 39.585 62.450 ;
        RECT 39.605 61.725 42.355 62.535 ;
        RECT 42.365 61.855 49.675 62.535 ;
        RECT 45.880 61.635 46.790 61.855 ;
        RECT 48.325 61.625 49.675 61.855 ;
        RECT 49.725 61.725 51.555 62.535 ;
        RECT 51.795 61.855 55.695 62.535 ;
        RECT 54.765 61.625 55.695 61.855 ;
        RECT 55.705 61.725 57.535 62.535 ;
        RECT 57.585 61.855 64.895 62.535 ;
        RECT 57.585 61.625 58.935 61.855 ;
        RECT 60.470 61.635 61.380 61.855 ;
        RECT 64.915 61.665 65.345 62.450 ;
        RECT 65.365 61.625 68.575 62.535 ;
        RECT 68.585 61.625 69.935 62.535 ;
        RECT 69.965 61.625 80.975 62.535 ;
        RECT 81.025 61.625 82.375 62.535 ;
        RECT 83.305 61.855 87.205 62.535 ;
        RECT 83.305 61.625 84.235 61.855 ;
        RECT 87.445 61.755 88.815 62.535 ;
        RECT 88.825 61.855 90.655 62.535 ;
        RECT 89.310 61.625 90.655 61.855 ;
        RECT 90.665 61.725 92.035 62.535 ;
      LAYER nwell ;
        RECT 13.190 58.505 92.230 61.335 ;
      LAYER pwell ;
        RECT 13.385 57.305 14.755 58.115 ;
        RECT 14.765 57.985 16.110 58.215 ;
        RECT 20.120 57.985 21.030 58.205 ;
        RECT 22.565 57.985 23.915 58.215 ;
        RECT 14.765 57.305 16.595 57.985 ;
        RECT 16.605 57.305 23.915 57.985 ;
        RECT 23.965 57.305 25.795 58.115 ;
        RECT 26.275 57.390 26.705 58.175 ;
        RECT 27.775 57.985 28.705 58.215 ;
        RECT 26.870 57.305 28.705 57.985 ;
        RECT 29.680 57.305 33.155 58.215 ;
        RECT 33.165 57.305 34.995 58.115 ;
        RECT 38.520 57.985 39.430 58.205 ;
        RECT 40.965 57.985 42.315 58.215 ;
        RECT 35.005 57.305 42.315 57.985 ;
        RECT 42.365 57.985 43.295 58.215 ;
        RECT 50.165 57.985 51.095 58.215 ;
        RECT 42.365 57.305 46.265 57.985 ;
        RECT 47.195 57.305 51.095 57.985 ;
        RECT 52.035 57.390 52.465 58.175 ;
        RECT 52.485 57.305 56.155 58.115 ;
        RECT 56.165 57.985 57.095 58.215 ;
        RECT 56.165 57.305 60.065 57.985 ;
        RECT 60.305 57.305 65.815 58.115 ;
        RECT 65.825 57.305 69.035 58.215 ;
        RECT 69.065 57.305 70.415 58.215 ;
        RECT 70.425 57.305 73.345 58.215 ;
        RECT 73.795 57.305 77.450 58.215 ;
        RECT 77.795 57.390 78.225 58.175 ;
        RECT 78.245 57.305 81.455 58.215 ;
        RECT 85.440 57.985 86.350 58.205 ;
        RECT 87.885 57.985 89.235 58.215 ;
        RECT 81.925 57.305 89.235 57.985 ;
        RECT 89.285 57.305 90.655 58.085 ;
        RECT 90.665 57.305 92.035 58.115 ;
        RECT 13.525 57.095 13.695 57.305 ;
        RECT 16.285 57.285 16.455 57.305 ;
        RECT 14.905 57.095 15.075 57.285 ;
        RECT 16.285 57.115 16.460 57.285 ;
        RECT 16.745 57.115 16.915 57.305 ;
        RECT 16.290 57.095 16.460 57.115 ;
        RECT 19.970 57.095 20.140 57.285 ;
        RECT 24.105 57.115 24.275 57.305 ;
        RECT 26.870 57.285 27.035 57.305 ;
        RECT 25.940 57.145 26.060 57.255 ;
        RECT 26.415 57.095 26.585 57.285 ;
        RECT 26.865 57.115 27.035 57.285 ;
        RECT 29.160 57.145 29.280 57.255 ;
        RECT 30.080 57.095 30.250 57.285 ;
        RECT 30.545 57.095 30.715 57.285 ;
        RECT 32.840 57.115 33.010 57.305 ;
        RECT 33.305 57.115 33.475 57.305 ;
        RECT 35.145 57.115 35.315 57.305 ;
        RECT 37.905 57.095 38.075 57.285 ;
        RECT 40.020 57.095 40.190 57.285 ;
        RECT 42.780 57.115 42.950 57.305 ;
        RECT 46.640 57.145 46.760 57.255 ;
        RECT 47.105 57.095 47.275 57.285 ;
        RECT 47.555 57.095 47.725 57.285 ;
        RECT 50.510 57.115 50.680 57.305 ;
        RECT 50.785 57.095 50.955 57.285 ;
        RECT 51.255 57.150 51.415 57.260 ;
        RECT 52.625 57.115 52.795 57.305 ;
        RECT 52.900 57.095 53.070 57.285 ;
        RECT 56.580 57.115 56.750 57.305 ;
        RECT 59.985 57.095 60.155 57.285 ;
        RECT 60.445 57.255 60.615 57.305 ;
        RECT 60.440 57.145 60.615 57.255 ;
        RECT 60.445 57.115 60.615 57.145 ;
        RECT 64.125 57.095 64.295 57.285 ;
        RECT 64.580 57.145 64.700 57.255 ;
        RECT 65.505 57.095 65.675 57.285 ;
        RECT 68.725 57.115 68.895 57.305 ;
        RECT 69.180 57.115 69.350 57.305 ;
        RECT 70.570 57.285 70.740 57.305 ;
        RECT 73.795 57.285 73.955 57.305 ;
        RECT 70.560 57.115 70.740 57.285 ;
        RECT 70.560 57.095 70.730 57.115 ;
        RECT 72.400 57.095 72.570 57.285 ;
        RECT 72.875 57.140 73.035 57.250 ;
        RECT 73.785 57.115 73.955 57.285 ;
        RECT 77.000 57.095 77.170 57.285 ;
        RECT 78.385 57.115 78.555 57.305 ;
        RECT 79.765 57.115 79.935 57.285 ;
        RECT 80.220 57.145 80.340 57.255 ;
        RECT 79.765 57.095 79.785 57.115 ;
        RECT 80.685 57.095 80.855 57.285 ;
        RECT 81.600 57.145 81.720 57.255 ;
        RECT 82.065 57.115 82.235 57.305 ;
        RECT 88.055 57.140 88.215 57.250 ;
        RECT 88.965 57.095 89.135 57.285 ;
        RECT 90.345 57.115 90.515 57.305 ;
        RECT 91.725 57.095 91.895 57.305 ;
        RECT 13.385 56.285 14.755 57.095 ;
        RECT 14.765 56.285 16.135 57.095 ;
        RECT 16.145 56.185 19.620 57.095 ;
        RECT 19.825 56.185 23.300 57.095 ;
        RECT 23.505 56.185 26.715 57.095 ;
        RECT 26.920 56.185 30.395 57.095 ;
        RECT 30.405 56.415 37.715 57.095 ;
        RECT 33.920 56.195 34.830 56.415 ;
        RECT 36.365 56.185 37.715 56.415 ;
        RECT 37.765 56.285 39.135 57.095 ;
        RECT 39.155 56.225 39.585 57.010 ;
        RECT 39.605 56.415 43.505 57.095 ;
        RECT 43.840 56.415 47.305 57.095 ;
        RECT 39.605 56.185 40.535 56.415 ;
        RECT 43.840 56.185 44.760 56.415 ;
        RECT 47.425 56.185 50.635 57.095 ;
        RECT 50.645 56.285 52.475 57.095 ;
        RECT 52.485 56.415 56.385 57.095 ;
        RECT 56.720 56.415 60.185 57.095 ;
        RECT 60.860 56.415 64.325 57.095 ;
        RECT 52.485 56.185 53.415 56.415 ;
        RECT 56.720 56.185 57.640 56.415 ;
        RECT 60.860 56.185 61.780 56.415 ;
        RECT 64.915 56.225 65.345 57.010 ;
        RECT 65.475 56.415 68.940 57.095 ;
        RECT 68.020 56.185 68.940 56.415 ;
        RECT 69.045 56.185 70.875 57.095 ;
        RECT 70.885 56.185 72.715 57.095 ;
        RECT 73.730 56.415 77.315 57.095 ;
        RECT 76.395 56.185 77.315 56.415 ;
        RECT 77.335 56.415 79.785 57.095 ;
        RECT 80.545 56.415 87.855 57.095 ;
        RECT 88.825 56.415 90.655 57.095 ;
        RECT 77.335 56.185 79.295 56.415 ;
        RECT 84.060 56.195 84.970 56.415 ;
        RECT 86.505 56.185 87.855 56.415 ;
        RECT 89.310 56.185 90.655 56.415 ;
        RECT 90.665 56.285 92.035 57.095 ;
      LAYER nwell ;
        RECT 13.190 53.065 92.230 55.895 ;
      LAYER pwell ;
        RECT 13.385 51.865 14.755 52.675 ;
        RECT 15.815 52.545 16.745 52.775 ;
        RECT 20.580 52.545 21.490 52.765 ;
        RECT 23.025 52.545 24.375 52.775 ;
        RECT 14.910 51.865 16.745 52.545 ;
        RECT 17.065 51.865 24.375 52.545 ;
        RECT 24.425 51.865 26.255 52.675 ;
        RECT 26.275 51.950 26.705 52.735 ;
        RECT 26.725 51.865 31.540 52.545 ;
        RECT 31.785 51.865 34.995 52.775 ;
        RECT 35.005 51.865 40.515 52.675 ;
        RECT 40.525 51.865 46.035 52.675 ;
        RECT 46.045 51.865 48.795 52.675 ;
        RECT 48.805 51.865 52.015 52.775 ;
        RECT 52.035 51.950 52.465 52.735 ;
        RECT 56.920 52.545 57.830 52.765 ;
        RECT 59.365 52.545 60.715 52.775 ;
        RECT 53.405 51.865 60.715 52.545 ;
        RECT 60.805 52.545 62.155 52.775 ;
        RECT 63.690 52.545 64.600 52.765 ;
        RECT 68.165 52.545 69.515 52.775 ;
        RECT 71.050 52.545 71.960 52.765 ;
        RECT 60.805 51.865 68.115 52.545 ;
        RECT 68.165 51.865 75.475 52.545 ;
        RECT 75.505 51.865 76.855 52.775 ;
        RECT 77.795 51.950 78.225 52.735 ;
        RECT 78.340 52.545 79.260 52.775 ;
        RECT 82.385 52.545 83.315 52.775 ;
        RECT 86.620 52.545 87.540 52.775 ;
        RECT 78.340 51.865 81.805 52.545 ;
        RECT 82.385 51.865 86.285 52.545 ;
        RECT 86.620 51.865 90.085 52.545 ;
        RECT 90.665 51.865 92.035 52.675 ;
        RECT 13.525 51.655 13.695 51.865 ;
        RECT 14.910 51.845 15.075 51.865 ;
        RECT 14.905 51.675 15.075 51.845 ;
        RECT 16.285 51.655 16.455 51.845 ;
        RECT 17.205 51.675 17.375 51.865 ;
        RECT 18.125 51.655 18.295 51.845 ;
        RECT 18.585 51.655 18.755 51.845 ;
        RECT 24.100 51.705 24.220 51.815 ;
        RECT 24.565 51.675 24.735 51.865 ;
        RECT 26.865 51.675 27.035 51.865 ;
        RECT 24.570 51.655 24.735 51.675 ;
        RECT 31.465 51.655 31.635 51.845 ;
        RECT 31.925 51.675 32.095 51.845 ;
        RECT 31.930 51.655 32.095 51.675 ;
        RECT 34.225 51.655 34.395 51.845 ;
        RECT 34.695 51.675 34.865 51.865 ;
        RECT 35.145 51.675 35.315 51.865 ;
        RECT 38.825 51.675 38.995 51.845 ;
        RECT 39.740 51.705 39.860 51.815 ;
        RECT 40.195 51.655 40.365 51.845 ;
        RECT 40.665 51.675 40.835 51.865 ;
        RECT 43.420 51.705 43.540 51.815 ;
        RECT 43.885 51.655 44.055 51.845 ;
        RECT 46.185 51.675 46.355 51.865 ;
        RECT 48.935 51.675 49.105 51.865 ;
        RECT 51.245 51.655 51.415 51.845 ;
        RECT 52.635 51.710 52.795 51.820 ;
        RECT 53.545 51.675 53.715 51.865 ;
        RECT 58.880 51.655 59.050 51.845 ;
        RECT 62.745 51.655 62.915 51.845 ;
        RECT 64.580 51.705 64.700 51.815 ;
        RECT 65.505 51.655 65.675 51.845 ;
        RECT 67.805 51.675 67.975 51.865 ;
        RECT 71.025 51.655 71.195 51.845 ;
        RECT 75.165 51.675 75.335 51.865 ;
        RECT 75.620 51.675 75.790 51.865 ;
        RECT 76.545 51.655 76.715 51.845 ;
        RECT 77.015 51.710 77.175 51.820 ;
        RECT 78.385 51.655 78.555 51.845 ;
        RECT 79.765 51.655 79.935 51.845 ;
        RECT 81.605 51.675 81.775 51.865 ;
        RECT 82.060 51.705 82.180 51.815 ;
        RECT 82.800 51.675 82.970 51.865 ;
        RECT 85.285 51.655 85.455 51.845 ;
        RECT 88.960 51.705 89.080 51.815 ;
        RECT 89.885 51.675 90.055 51.865 ;
        RECT 90.345 51.815 90.515 51.845 ;
        RECT 90.340 51.705 90.515 51.815 ;
        RECT 90.345 51.655 90.515 51.705 ;
        RECT 91.725 51.655 91.895 51.865 ;
        RECT 13.385 50.845 14.755 51.655 ;
        RECT 14.765 50.975 16.595 51.655 ;
        RECT 16.605 50.975 18.435 51.655 ;
        RECT 14.765 50.745 16.110 50.975 ;
        RECT 16.605 50.745 17.950 50.975 ;
        RECT 18.445 50.845 23.955 51.655 ;
        RECT 24.570 50.975 26.405 51.655 ;
        RECT 26.960 50.975 31.775 51.655 ;
        RECT 31.930 50.975 33.765 51.655 ;
        RECT 25.475 50.745 26.405 50.975 ;
        RECT 32.835 50.745 33.765 50.975 ;
        RECT 34.085 50.845 35.915 51.655 ;
        RECT 36.305 50.975 38.730 51.655 ;
        RECT 39.155 50.785 39.585 51.570 ;
        RECT 40.065 50.745 43.275 51.655 ;
        RECT 43.745 50.975 51.055 51.655 ;
        RECT 51.105 50.975 58.415 51.655 ;
        RECT 47.260 50.755 48.170 50.975 ;
        RECT 49.705 50.745 51.055 50.975 ;
        RECT 54.620 50.755 55.530 50.975 ;
        RECT 57.065 50.745 58.415 50.975 ;
        RECT 58.465 50.975 62.365 51.655 ;
        RECT 58.465 50.745 59.395 50.975 ;
        RECT 62.605 50.845 64.435 51.655 ;
        RECT 64.915 50.785 65.345 51.570 ;
        RECT 65.365 50.845 70.875 51.655 ;
        RECT 70.885 50.845 76.395 51.655 ;
        RECT 76.405 50.845 78.235 51.655 ;
        RECT 78.255 50.745 79.605 51.655 ;
        RECT 79.625 50.845 85.135 51.655 ;
        RECT 85.145 50.845 88.815 51.655 ;
        RECT 89.285 50.875 90.655 51.655 ;
        RECT 90.665 50.845 92.035 51.655 ;
      LAYER nwell ;
        RECT 13.190 47.625 92.230 50.455 ;
      LAYER pwell ;
        RECT 13.385 46.425 14.755 47.235 ;
        RECT 14.765 47.105 16.110 47.335 ;
        RECT 14.765 46.425 16.595 47.105 ;
        RECT 17.720 46.425 21.195 47.335 ;
        RECT 21.205 47.105 22.550 47.335 ;
        RECT 21.205 46.425 23.035 47.105 ;
        RECT 23.045 46.425 25.795 47.235 ;
        RECT 26.275 46.510 26.705 47.295 ;
        RECT 27.380 46.425 30.855 47.335 ;
        RECT 34.380 47.105 35.290 47.325 ;
        RECT 36.825 47.105 38.175 47.335 ;
        RECT 41.740 47.105 42.650 47.325 ;
        RECT 44.185 47.105 45.535 47.335 ;
        RECT 30.865 46.425 38.175 47.105 ;
        RECT 38.225 46.425 45.535 47.105 ;
        RECT 45.585 47.105 46.515 47.335 ;
        RECT 45.585 46.425 49.485 47.105 ;
        RECT 49.725 46.425 51.555 47.235 ;
        RECT 52.035 46.510 52.465 47.295 ;
        RECT 52.580 47.105 53.500 47.335 ;
        RECT 57.505 47.135 58.915 47.335 ;
        RECT 52.580 46.425 56.045 47.105 ;
        RECT 56.180 46.455 58.915 47.135 ;
        RECT 13.525 46.215 13.695 46.425 ;
        RECT 14.905 46.215 15.075 46.405 ;
        RECT 16.285 46.235 16.455 46.425 ;
        RECT 16.755 46.270 16.915 46.380 ;
        RECT 16.290 46.215 16.455 46.235 ;
        RECT 18.585 46.215 18.755 46.405 ;
        RECT 20.880 46.235 21.050 46.425 ;
        RECT 22.725 46.235 22.895 46.425 ;
        RECT 23.185 46.235 23.355 46.425 ;
        RECT 25.945 46.375 26.115 46.405 ;
        RECT 25.940 46.265 26.115 46.375 ;
        RECT 26.860 46.265 26.980 46.375 ;
        RECT 25.945 46.235 26.115 46.265 ;
        RECT 30.540 46.235 30.710 46.425 ;
        RECT 31.005 46.235 31.175 46.425 ;
        RECT 25.950 46.215 26.115 46.235 ;
        RECT 31.460 46.215 31.630 46.405 ;
        RECT 31.925 46.215 32.095 46.405 ;
        RECT 38.365 46.235 38.535 46.425 ;
        RECT 39.745 46.215 39.915 46.405 ;
        RECT 46.000 46.235 46.170 46.425 ;
        RECT 48.025 46.215 48.195 46.405 ;
        RECT 48.485 46.215 48.655 46.405 ;
        RECT 49.865 46.235 50.035 46.425 ;
        RECT 51.250 46.215 51.420 46.405 ;
        RECT 51.700 46.265 51.820 46.375 ;
        RECT 54.925 46.215 55.095 46.405 ;
        RECT 55.845 46.235 56.015 46.425 ;
        RECT 56.305 46.235 56.475 46.455 ;
        RECT 57.520 46.425 58.915 46.455 ;
        RECT 58.925 46.425 60.755 47.105 ;
        RECT 60.765 46.425 62.135 47.235 ;
        RECT 62.145 46.425 65.355 47.335 ;
        RECT 66.025 47.105 69.955 47.335 ;
        RECT 65.540 46.425 69.955 47.105 ;
        RECT 69.965 46.425 73.175 47.335 ;
        RECT 73.495 47.105 74.425 47.335 ;
        RECT 73.495 46.425 75.330 47.105 ;
        RECT 75.485 46.425 77.315 47.235 ;
        RECT 77.795 46.510 78.225 47.295 ;
        RECT 78.440 46.425 81.915 47.335 ;
        RECT 81.925 46.425 87.435 47.235 ;
        RECT 87.445 46.425 90.195 47.235 ;
        RECT 90.665 46.425 92.035 47.235 ;
        RECT 56.765 46.215 56.935 46.405 ;
        RECT 59.065 46.235 59.235 46.425 ;
        RECT 59.535 46.260 59.695 46.370 ;
        RECT 60.905 46.235 61.075 46.425 ;
        RECT 62.280 46.215 62.450 46.405 ;
        RECT 62.745 46.215 62.915 46.405 ;
        RECT 64.580 46.265 64.700 46.375 ;
        RECT 65.045 46.235 65.215 46.425 ;
        RECT 65.540 46.405 65.650 46.425 ;
        RECT 65.480 46.235 65.675 46.405 ;
        RECT 68.725 46.235 68.895 46.405 ;
        RECT 65.505 46.215 65.675 46.235 ;
        RECT 69.185 46.215 69.355 46.405 ;
        RECT 70.105 46.235 70.275 46.425 ;
        RECT 75.165 46.405 75.330 46.425 ;
        RECT 74.245 46.215 74.415 46.405 ;
        RECT 75.165 46.235 75.335 46.405 ;
        RECT 75.625 46.235 75.795 46.425 ;
        RECT 81.600 46.405 81.770 46.425 ;
        RECT 77.460 46.265 77.580 46.375 ;
        RECT 81.600 46.235 81.775 46.405 ;
        RECT 82.065 46.235 82.235 46.425 ;
        RECT 81.605 46.215 81.775 46.235 ;
        RECT 87.125 46.215 87.295 46.405 ;
        RECT 87.585 46.235 87.755 46.425 ;
        RECT 88.965 46.215 89.135 46.405 ;
        RECT 90.340 46.265 90.460 46.375 ;
        RECT 91.725 46.215 91.895 46.425 ;
        RECT 13.385 45.405 14.755 46.215 ;
        RECT 14.765 45.405 16.135 46.215 ;
        RECT 16.290 45.535 18.125 46.215 ;
        RECT 18.445 45.535 25.755 46.215 ;
        RECT 25.950 45.535 27.785 46.215 ;
        RECT 17.195 45.305 18.125 45.535 ;
        RECT 21.960 45.315 22.870 45.535 ;
        RECT 24.405 45.305 25.755 45.535 ;
        RECT 26.855 45.305 27.785 45.535 ;
        RECT 28.300 45.305 31.775 46.215 ;
        RECT 31.785 45.535 39.095 46.215 ;
        RECT 35.300 45.315 36.210 45.535 ;
        RECT 37.745 45.305 39.095 45.535 ;
        RECT 39.155 45.345 39.585 46.130 ;
        RECT 39.605 45.535 44.420 46.215 ;
        RECT 44.760 45.535 48.225 46.215 ;
        RECT 48.345 45.535 51.085 46.215 ;
        RECT 44.760 45.305 45.680 45.535 ;
        RECT 51.110 45.305 54.695 46.215 ;
        RECT 54.785 45.405 56.615 46.215 ;
        RECT 56.625 45.405 58.715 46.215 ;
        RECT 60.405 45.305 62.595 46.215 ;
        RECT 62.605 45.405 64.435 46.215 ;
        RECT 64.915 45.345 65.345 46.130 ;
        RECT 65.365 45.405 67.195 46.215 ;
        RECT 67.205 45.535 68.570 46.215 ;
        RECT 69.045 45.535 73.860 46.215 ;
        RECT 74.105 45.535 81.415 46.215 ;
        RECT 77.620 45.315 78.530 45.535 ;
        RECT 80.065 45.305 81.415 45.535 ;
        RECT 81.465 45.405 86.975 46.215 ;
        RECT 86.985 45.405 88.815 46.215 ;
        RECT 88.825 45.535 90.655 46.215 ;
        RECT 89.310 45.305 90.655 45.535 ;
        RECT 90.665 45.405 92.035 46.215 ;
      LAYER nwell ;
        RECT 13.190 42.185 92.230 45.015 ;
      LAYER pwell ;
        RECT 13.385 40.985 14.755 41.795 ;
        RECT 18.280 41.665 19.190 41.885 ;
        RECT 20.725 41.665 22.075 41.895 ;
        RECT 14.765 40.985 22.075 41.665 ;
        RECT 22.125 41.665 23.470 41.895 ;
        RECT 22.125 40.985 23.955 41.665 ;
        RECT 23.965 40.985 25.795 41.795 ;
        RECT 26.275 41.070 26.705 41.855 ;
        RECT 26.725 40.985 29.935 41.895 ;
        RECT 29.960 41.665 31.330 41.895 ;
        RECT 29.960 40.985 32.235 41.665 ;
        RECT 32.255 40.985 33.605 41.895 ;
        RECT 33.625 40.985 39.135 41.795 ;
        RECT 39.605 41.665 40.535 41.895 ;
        RECT 48.180 41.665 49.090 41.885 ;
        RECT 50.625 41.665 51.975 41.895 ;
        RECT 39.605 40.985 43.505 41.665 ;
        RECT 44.665 40.985 51.975 41.665 ;
        RECT 52.035 41.070 52.465 41.855 ;
        RECT 52.495 40.985 53.845 41.895 ;
        RECT 57.380 41.665 58.290 41.885 ;
        RECT 59.825 41.665 61.175 41.895 ;
        RECT 65.660 41.665 66.570 41.885 ;
        RECT 68.105 41.665 69.455 41.895 ;
        RECT 53.865 40.985 61.175 41.665 ;
        RECT 62.145 40.985 69.455 41.665 ;
        RECT 70.620 40.985 74.095 41.895 ;
        RECT 75.155 41.665 76.085 41.895 ;
        RECT 74.250 40.985 76.085 41.665 ;
        RECT 76.405 40.985 77.775 41.795 ;
        RECT 77.795 41.070 78.225 41.855 ;
        RECT 81.760 41.665 82.670 41.885 ;
        RECT 84.205 41.665 85.555 41.895 ;
        RECT 78.245 40.985 85.555 41.665 ;
        RECT 85.605 40.985 89.275 41.795 ;
        RECT 89.285 40.985 90.655 41.795 ;
        RECT 90.665 40.985 92.035 41.795 ;
        RECT 13.525 40.775 13.695 40.985 ;
        RECT 14.905 40.795 15.075 40.985 ;
        RECT 15.830 40.775 16.000 40.965 ;
        RECT 21.345 40.795 21.515 40.965 ;
        RECT 21.345 40.775 21.510 40.795 ;
        RECT 21.805 40.775 21.975 40.965 ;
        RECT 23.645 40.795 23.815 40.985 ;
        RECT 24.105 40.795 24.275 40.985 ;
        RECT 25.025 40.775 25.195 40.965 ;
        RECT 25.940 40.825 26.060 40.935 ;
        RECT 28.700 40.825 28.820 40.935 ;
        RECT 29.170 40.775 29.340 40.965 ;
        RECT 29.635 40.795 29.805 40.985 ;
        RECT 30.545 40.775 30.715 40.965 ;
        RECT 31.920 40.795 32.090 40.985 ;
        RECT 32.385 40.795 32.555 40.985 ;
        RECT 33.765 40.795 33.935 40.985 ;
        RECT 33.765 40.775 33.915 40.795 ;
        RECT 34.225 40.775 34.395 40.965 ;
        RECT 37.905 40.775 38.075 40.965 ;
        RECT 39.280 40.825 39.400 40.935 ;
        RECT 39.745 40.775 39.915 40.965 ;
        RECT 40.020 40.795 40.190 40.985 ;
        RECT 41.575 40.775 41.745 40.965 ;
        RECT 43.895 40.830 44.055 40.940 ;
        RECT 44.805 40.775 44.975 40.985 ;
        RECT 47.560 40.825 47.680 40.935 ;
        RECT 48.300 40.775 48.470 40.965 ;
        RECT 52.625 40.795 52.795 40.985 ;
        RECT 54.005 40.795 54.175 40.985 ;
        RECT 13.385 39.965 14.755 40.775 ;
        RECT 15.685 39.865 19.160 40.775 ;
        RECT 19.675 40.095 21.510 40.775 ;
        RECT 19.675 39.865 20.605 40.095 ;
        RECT 21.665 39.865 24.875 40.775 ;
        RECT 24.885 39.965 28.555 40.775 ;
        RECT 29.025 39.865 30.375 40.775 ;
        RECT 30.405 39.965 31.775 40.775 ;
        RECT 31.985 39.955 33.915 40.775 ;
        RECT 34.085 39.965 37.755 40.775 ;
        RECT 37.765 39.965 39.135 40.775 ;
        RECT 31.985 39.865 32.935 39.955 ;
        RECT 39.155 39.905 39.585 40.690 ;
        RECT 39.605 39.965 41.435 40.775 ;
        RECT 41.445 39.865 44.655 40.775 ;
        RECT 44.665 39.965 47.415 40.775 ;
        RECT 47.885 40.095 51.785 40.775 ;
        RECT 52.025 40.745 53.420 40.775 ;
        RECT 54.465 40.745 54.635 40.965 ;
        RECT 54.920 40.825 55.040 40.935 ;
        RECT 56.305 40.775 56.475 40.965 ;
        RECT 61.365 40.775 61.535 40.965 ;
        RECT 61.825 40.795 61.995 40.965 ;
        RECT 62.285 40.795 62.455 40.985 ;
        RECT 64.580 40.825 64.700 40.935 ;
        RECT 61.855 40.775 61.995 40.795 ;
        RECT 65.510 40.775 65.680 40.965 ;
        RECT 69.180 40.825 69.300 40.935 ;
        RECT 69.645 40.795 69.815 40.965 ;
        RECT 69.650 40.775 69.815 40.795 ;
        RECT 71.950 40.775 72.120 40.965 ;
        RECT 73.780 40.795 73.950 40.985 ;
        RECT 74.250 40.965 74.415 40.985 ;
        RECT 74.245 40.795 74.415 40.965 ;
        RECT 74.265 40.775 74.415 40.795 ;
        RECT 76.545 40.775 76.715 40.985 ;
        RECT 78.385 40.795 78.555 40.985 ;
        RECT 83.440 40.775 83.610 40.965 ;
        RECT 84.815 40.775 84.985 40.965 ;
        RECT 85.285 40.775 85.455 40.965 ;
        RECT 85.745 40.795 85.915 40.985 ;
        RECT 89.425 40.795 89.595 40.985 ;
        RECT 91.725 40.775 91.895 40.985 ;
        RECT 47.885 39.865 48.815 40.095 ;
        RECT 52.025 40.065 54.760 40.745 ;
        RECT 52.025 39.865 53.435 40.065 ;
        RECT 55.255 39.865 56.605 40.775 ;
        RECT 56.860 40.095 61.675 40.775 ;
        RECT 61.855 39.955 64.425 40.775 ;
        RECT 62.835 39.865 64.425 39.955 ;
        RECT 64.915 39.905 65.345 40.690 ;
        RECT 65.365 39.865 68.840 40.775 ;
        RECT 69.650 40.095 71.485 40.775 ;
        RECT 70.555 39.865 71.485 40.095 ;
        RECT 71.805 39.865 73.995 40.775 ;
        RECT 74.265 39.955 76.195 40.775 ;
        RECT 76.405 39.965 80.075 40.775 ;
        RECT 75.245 39.865 76.195 39.955 ;
        RECT 80.280 39.865 83.755 40.775 ;
        RECT 83.765 39.995 85.135 40.775 ;
        RECT 85.145 39.965 90.655 40.775 ;
        RECT 90.665 39.965 92.035 40.775 ;
      LAYER nwell ;
        RECT 13.190 36.745 92.230 39.575 ;
      LAYER pwell ;
        RECT 13.385 35.545 14.755 36.355 ;
        RECT 14.765 35.545 17.515 36.355 ;
        RECT 21.500 36.225 22.410 36.445 ;
        RECT 23.945 36.225 25.295 36.455 ;
        RECT 17.985 35.545 25.295 36.225 ;
        RECT 26.275 35.630 26.705 36.415 ;
        RECT 27.035 36.225 27.965 36.455 ;
        RECT 27.035 35.545 28.870 36.225 ;
        RECT 30.140 35.545 33.615 36.455 ;
        RECT 33.725 35.545 35.915 36.455 ;
        RECT 35.925 35.545 37.755 36.355 ;
        RECT 37.805 36.225 39.155 36.455 ;
        RECT 40.690 36.225 41.600 36.445 ;
        RECT 37.805 35.545 45.115 36.225 ;
        RECT 45.125 35.545 48.600 36.455 ;
        RECT 48.805 35.545 51.555 36.355 ;
        RECT 52.035 35.630 52.465 36.415 ;
        RECT 52.485 35.545 55.235 36.355 ;
        RECT 55.245 36.225 56.175 36.455 ;
        RECT 59.480 36.225 60.400 36.455 ;
        RECT 55.245 35.545 59.145 36.225 ;
        RECT 59.480 35.545 62.945 36.225 ;
        RECT 63.065 35.545 64.895 36.225 ;
        RECT 64.905 35.545 70.415 36.355 ;
        RECT 70.425 35.545 74.095 36.355 ;
        RECT 74.105 35.545 75.475 36.355 ;
        RECT 76.535 36.225 77.465 36.455 ;
        RECT 75.630 35.545 77.465 36.225 ;
        RECT 77.795 35.630 78.225 36.415 ;
        RECT 79.360 35.545 82.835 36.455 ;
        RECT 86.360 36.225 87.270 36.445 ;
        RECT 88.805 36.225 90.155 36.455 ;
        RECT 82.845 35.545 90.155 36.225 ;
        RECT 90.665 35.545 92.035 36.355 ;
        RECT 13.525 35.335 13.695 35.545 ;
        RECT 14.905 35.335 15.075 35.545 ;
        RECT 17.660 35.385 17.780 35.495 ;
        RECT 18.125 35.355 18.295 35.545 ;
        RECT 28.705 35.525 28.870 35.545 ;
        RECT 20.435 35.380 20.595 35.490 ;
        RECT 21.350 35.335 21.520 35.525 ;
        RECT 25.025 35.335 25.195 35.525 ;
        RECT 25.495 35.390 25.655 35.500 ;
        RECT 26.865 35.335 27.035 35.525 ;
        RECT 28.705 35.355 28.875 35.525 ;
        RECT 29.175 35.390 29.335 35.500 ;
        RECT 28.710 35.335 28.875 35.355 ;
        RECT 31.005 35.335 31.175 35.525 ;
        RECT 33.300 35.355 33.470 35.545 ;
        RECT 35.600 35.355 35.770 35.545 ;
        RECT 36.065 35.355 36.235 35.545 ;
        RECT 38.375 35.380 38.535 35.490 ;
        RECT 39.745 35.335 39.915 35.525 ;
        RECT 42.965 35.355 43.135 35.525 ;
        RECT 44.805 35.355 44.975 35.545 ;
        RECT 45.270 35.525 45.440 35.545 ;
        RECT 45.265 35.355 45.440 35.525 ;
        RECT 48.945 35.355 49.115 35.545 ;
        RECT 52.625 35.525 52.795 35.545 ;
        RECT 42.970 35.335 43.135 35.355 ;
        RECT 45.265 35.335 45.435 35.355 ;
        RECT 50.785 35.335 50.955 35.525 ;
        RECT 51.700 35.385 51.820 35.495 ;
        RECT 52.625 35.355 52.800 35.525 ;
        RECT 55.660 35.355 55.830 35.545 ;
        RECT 52.630 35.335 52.800 35.355 ;
        RECT 56.305 35.335 56.475 35.525 ;
        RECT 57.685 35.335 57.855 35.525 ;
        RECT 62.745 35.355 62.915 35.545 ;
        RECT 63.205 35.355 63.375 35.545 ;
        RECT 65.045 35.355 65.215 35.545 ;
        RECT 65.505 35.335 65.675 35.525 ;
        RECT 69.180 35.385 69.300 35.495 ;
        RECT 70.565 35.355 70.735 35.545 ;
        RECT 71.945 35.355 72.115 35.525 ;
        RECT 71.945 35.335 72.085 35.355 ;
        RECT 72.410 35.335 72.580 35.525 ;
        RECT 74.245 35.355 74.415 35.545 ;
        RECT 75.630 35.525 75.795 35.545 ;
        RECT 74.705 35.335 74.875 35.525 ;
        RECT 75.625 35.355 75.795 35.525 ;
        RECT 76.540 35.385 76.660 35.495 ;
        RECT 77.005 35.355 77.175 35.525 ;
        RECT 78.395 35.390 78.555 35.500 ;
        RECT 77.010 35.335 77.175 35.355 ;
        RECT 82.065 35.335 82.235 35.525 ;
        RECT 82.520 35.490 82.690 35.545 ;
        RECT 82.520 35.380 82.695 35.490 ;
        RECT 82.520 35.355 82.690 35.380 ;
        RECT 82.985 35.355 83.155 35.545 ;
        RECT 83.445 35.335 83.615 35.525 ;
        RECT 90.340 35.385 90.460 35.495 ;
        RECT 91.725 35.335 91.895 35.545 ;
        RECT 13.385 34.525 14.755 35.335 ;
        RECT 14.765 34.525 20.275 35.335 ;
        RECT 21.205 34.425 24.680 35.335 ;
        RECT 24.885 34.655 26.715 35.335 ;
        RECT 25.370 34.425 26.715 34.655 ;
        RECT 26.725 34.525 28.555 35.335 ;
        RECT 28.710 34.655 30.545 35.335 ;
        RECT 30.865 34.655 38.175 35.335 ;
        RECT 29.615 34.425 30.545 34.655 ;
        RECT 34.380 34.435 35.290 34.655 ;
        RECT 36.825 34.425 38.175 34.655 ;
        RECT 39.155 34.465 39.585 35.250 ;
        RECT 39.605 34.425 42.815 35.335 ;
        RECT 42.970 34.655 44.805 35.335 ;
        RECT 43.875 34.425 44.805 34.655 ;
        RECT 45.125 34.525 50.635 35.335 ;
        RECT 50.645 34.525 52.475 35.335 ;
        RECT 52.490 34.425 56.075 35.335 ;
        RECT 56.165 34.525 57.535 35.335 ;
        RECT 57.545 34.655 64.855 35.335 ;
        RECT 61.060 34.435 61.970 34.655 ;
        RECT 63.505 34.425 64.855 34.655 ;
        RECT 64.915 34.465 65.345 35.250 ;
        RECT 65.365 34.525 69.035 35.335 ;
        RECT 69.515 34.515 72.085 35.335 ;
        RECT 69.515 34.425 71.105 34.515 ;
        RECT 72.265 34.425 74.455 35.335 ;
        RECT 74.565 34.525 76.395 35.335 ;
        RECT 77.010 34.655 78.845 35.335 ;
        RECT 77.915 34.425 78.845 34.655 ;
        RECT 79.165 34.425 82.375 35.335 ;
        RECT 83.305 34.655 90.615 35.335 ;
        RECT 86.820 34.435 87.730 34.655 ;
        RECT 89.265 34.425 90.615 34.655 ;
        RECT 90.665 34.525 92.035 35.335 ;
      LAYER nwell ;
        RECT 13.190 31.305 92.230 34.135 ;
      LAYER pwell ;
        RECT 13.385 30.105 14.755 30.915 ;
        RECT 14.765 30.785 16.110 31.015 ;
        RECT 17.375 30.785 18.305 31.015 ;
        RECT 14.765 30.105 16.595 30.785 ;
        RECT 17.375 30.105 19.210 30.785 ;
        RECT 19.365 30.105 21.195 30.915 ;
        RECT 21.665 30.105 25.140 31.015 ;
        RECT 26.275 30.190 26.705 30.975 ;
        RECT 26.725 30.105 32.235 30.915 ;
        RECT 32.245 30.105 37.755 30.915 ;
        RECT 37.765 30.105 43.275 30.915 ;
        RECT 45.255 30.785 46.185 31.015 ;
        RECT 44.350 30.105 46.185 30.785 ;
        RECT 46.505 30.105 48.335 30.915 ;
        RECT 48.805 30.105 52.015 31.015 ;
        RECT 52.035 30.190 52.465 30.975 ;
        RECT 52.485 30.105 53.855 30.915 ;
        RECT 54.060 30.105 57.535 31.015 ;
        RECT 57.855 30.785 58.785 31.015 ;
        RECT 63.360 30.785 64.270 31.005 ;
        RECT 65.805 30.785 67.155 31.015 ;
        RECT 57.855 30.105 59.690 30.785 ;
        RECT 59.845 30.105 67.155 30.785 ;
        RECT 67.515 30.785 68.445 31.015 ;
        RECT 73.020 30.785 73.930 31.005 ;
        RECT 75.465 30.785 76.815 31.015 ;
        RECT 67.515 30.105 69.350 30.785 ;
        RECT 69.505 30.105 76.815 30.785 ;
        RECT 77.795 30.190 78.225 30.975 ;
        RECT 79.755 30.785 80.685 31.015 ;
        RECT 78.850 30.105 80.685 30.785 ;
        RECT 81.005 30.105 86.515 30.915 ;
        RECT 86.525 30.105 88.355 30.915 ;
        RECT 89.310 30.785 90.655 31.015 ;
        RECT 88.825 30.105 90.655 30.785 ;
        RECT 90.665 30.105 92.035 30.915 ;
        RECT 13.525 29.895 13.695 30.105 ;
        RECT 14.900 29.945 15.020 30.055 ;
        RECT 15.370 29.895 15.540 30.085 ;
        RECT 16.285 29.915 16.455 30.105 ;
        RECT 19.045 30.085 19.210 30.105 ;
        RECT 16.740 29.945 16.860 30.055 ;
        RECT 19.045 29.895 19.215 30.085 ;
        RECT 19.505 29.915 19.675 30.105 ;
        RECT 21.340 29.945 21.460 30.055 ;
        RECT 21.810 29.915 21.980 30.105 ;
        RECT 25.495 29.950 25.655 30.060 ;
        RECT 26.865 29.915 27.035 30.105 ;
        RECT 28.245 29.915 28.415 30.085 ;
        RECT 28.700 29.945 28.820 30.055 ;
        RECT 28.245 29.895 28.410 29.915 ;
        RECT 29.170 29.895 29.340 30.085 ;
        RECT 32.385 29.915 32.555 30.105 ;
        RECT 32.840 29.945 32.960 30.055 ;
        RECT 36.520 29.895 36.690 30.085 ;
        RECT 36.985 29.915 37.155 30.085 ;
        RECT 37.905 29.915 38.075 30.105 ;
        RECT 44.350 30.085 44.515 30.105 ;
        RECT 36.990 29.895 37.155 29.915 ;
        RECT 39.745 29.895 39.915 30.085 ;
        RECT 42.505 29.895 42.675 30.085 ;
        RECT 43.435 29.950 43.595 30.060 ;
        RECT 44.345 29.915 44.515 30.085 ;
        RECT 46.645 29.915 46.815 30.105 ;
        RECT 48.480 29.945 48.600 30.055 ;
        RECT 48.945 29.915 49.115 30.105 ;
        RECT 49.865 29.895 50.035 30.085 ;
        RECT 51.245 29.895 51.415 30.085 ;
        RECT 52.625 29.915 52.795 30.105 ;
        RECT 57.220 29.915 57.390 30.105 ;
        RECT 59.525 30.085 59.690 30.105 ;
        RECT 58.600 29.945 58.720 30.055 ;
        RECT 59.070 29.895 59.240 30.085 ;
        RECT 59.525 29.915 59.695 30.085 ;
        RECT 59.985 29.915 60.155 30.105 ;
        RECT 69.185 30.085 69.350 30.105 ;
        RECT 64.585 29.915 64.755 30.085 ;
        RECT 65.515 29.940 65.675 30.050 ;
        RECT 64.585 29.895 64.750 29.915 ;
        RECT 69.185 29.895 69.355 30.085 ;
        RECT 69.645 29.915 69.815 30.105 ;
        RECT 78.850 30.085 79.015 30.105 ;
        RECT 72.860 29.895 73.030 30.085 ;
        RECT 73.325 29.895 73.495 30.085 ;
        RECT 75.160 29.945 75.280 30.055 ;
        RECT 75.625 29.895 75.795 30.085 ;
        RECT 77.015 29.950 77.175 30.060 ;
        RECT 78.380 29.945 78.500 30.055 ;
        RECT 78.845 29.915 79.015 30.085 ;
        RECT 81.145 29.915 81.315 30.105 ;
        RECT 85.745 29.895 85.915 30.085 ;
        RECT 86.205 29.895 86.375 30.085 ;
        RECT 86.665 29.915 86.835 30.105 ;
        RECT 88.500 29.945 88.620 30.055 ;
        RECT 88.965 29.915 89.135 30.105 ;
        RECT 89.895 29.940 90.055 30.050 ;
        RECT 91.725 29.895 91.895 30.105 ;
        RECT 13.385 29.085 14.755 29.895 ;
        RECT 15.225 28.985 18.700 29.895 ;
        RECT 18.905 29.215 26.215 29.895 ;
        RECT 22.420 28.995 23.330 29.215 ;
        RECT 24.865 28.985 26.215 29.215 ;
        RECT 26.575 29.215 28.410 29.895 ;
        RECT 26.575 28.985 27.505 29.215 ;
        RECT 29.025 28.985 32.500 29.895 ;
        RECT 33.360 28.985 36.835 29.895 ;
        RECT 36.990 29.215 38.825 29.895 ;
        RECT 37.895 28.985 38.825 29.215 ;
        RECT 39.155 29.025 39.585 29.810 ;
        RECT 39.605 29.085 42.355 29.895 ;
        RECT 42.365 29.215 49.675 29.895 ;
        RECT 45.880 28.995 46.790 29.215 ;
        RECT 48.325 28.985 49.675 29.215 ;
        RECT 49.725 29.085 51.095 29.895 ;
        RECT 51.105 29.215 58.415 29.895 ;
        RECT 54.620 28.995 55.530 29.215 ;
        RECT 57.065 28.985 58.415 29.215 ;
        RECT 58.925 28.985 62.400 29.895 ;
        RECT 62.915 29.215 64.750 29.895 ;
        RECT 62.915 28.985 63.845 29.215 ;
        RECT 64.915 29.025 65.345 29.810 ;
        RECT 66.285 28.985 69.495 29.895 ;
        RECT 69.700 28.985 73.175 29.895 ;
        RECT 73.185 29.085 75.015 29.895 ;
        RECT 75.485 29.215 82.795 29.895 ;
        RECT 79.000 28.995 79.910 29.215 ;
        RECT 81.445 28.985 82.795 29.215 ;
        RECT 82.845 28.985 86.055 29.895 ;
        RECT 86.065 29.085 89.735 29.895 ;
        RECT 90.665 29.085 92.035 29.895 ;
      LAYER nwell ;
        RECT 13.190 25.865 92.230 28.695 ;
      LAYER pwell ;
        RECT 13.385 24.665 14.755 25.475 ;
        RECT 18.280 25.345 19.190 25.565 ;
        RECT 20.725 25.345 22.075 25.575 ;
        RECT 14.765 24.665 22.075 25.345 ;
        RECT 22.125 24.665 25.335 25.575 ;
        RECT 26.275 24.750 26.705 25.535 ;
        RECT 26.725 24.665 28.095 25.475 ;
        RECT 31.620 25.345 32.530 25.565 ;
        RECT 34.065 25.345 35.415 25.575 ;
        RECT 38.980 25.345 39.890 25.565 ;
        RECT 41.425 25.345 42.775 25.575 ;
        RECT 28.105 24.665 35.415 25.345 ;
        RECT 35.465 24.665 42.775 25.345 ;
        RECT 43.745 24.665 47.220 25.575 ;
        RECT 47.425 24.665 49.255 25.475 ;
        RECT 50.775 25.345 51.705 25.575 ;
        RECT 49.870 24.665 51.705 25.345 ;
        RECT 52.035 24.750 52.465 25.535 ;
        RECT 52.485 24.665 55.960 25.575 ;
        RECT 56.165 24.665 57.995 25.475 ;
        RECT 58.005 25.345 59.350 25.575 ;
        RECT 58.005 24.665 59.835 25.345 ;
        RECT 59.845 24.665 65.355 25.475 ;
        RECT 65.365 24.665 70.875 25.475 ;
        RECT 70.885 24.665 74.555 25.475 ;
        RECT 76.535 25.345 77.465 25.575 ;
        RECT 75.630 24.665 77.465 25.345 ;
        RECT 77.795 24.750 78.225 25.535 ;
        RECT 78.245 24.665 81.720 25.575 ;
        RECT 81.925 24.665 83.295 25.475 ;
        RECT 86.820 25.345 87.730 25.565 ;
        RECT 89.265 25.345 90.615 25.575 ;
        RECT 83.305 24.665 90.615 25.345 ;
        RECT 90.665 24.665 92.035 25.475 ;
        RECT 13.525 24.455 13.695 24.665 ;
        RECT 14.905 24.475 15.075 24.665 ;
        RECT 16.285 24.455 16.455 24.645 ;
        RECT 16.745 24.455 16.915 24.645 ;
        RECT 19.505 24.455 19.675 24.645 ;
        RECT 21.345 24.455 21.515 24.645 ;
        RECT 21.815 24.500 21.975 24.610 ;
        RECT 22.265 24.475 22.435 24.665 ;
        RECT 22.725 24.455 22.895 24.645 ;
        RECT 25.495 24.510 25.655 24.620 ;
        RECT 25.945 24.455 26.115 24.645 ;
        RECT 26.865 24.475 27.035 24.665 ;
        RECT 27.795 24.500 27.955 24.610 ;
        RECT 28.245 24.475 28.415 24.665 ;
        RECT 28.705 24.475 28.875 24.645 ;
        RECT 28.710 24.455 28.875 24.475 ;
        RECT 31.005 24.455 31.175 24.645 ;
        RECT 35.605 24.475 35.775 24.665 ;
        RECT 36.525 24.455 36.695 24.645 ;
        RECT 39.745 24.455 39.915 24.645 ;
        RECT 41.585 24.455 41.755 24.645 ;
        RECT 42.975 24.510 43.135 24.620 ;
        RECT 43.890 24.475 44.060 24.665 ;
        RECT 44.805 24.455 44.975 24.645 ;
        RECT 46.185 24.455 46.355 24.645 ;
        RECT 47.565 24.475 47.735 24.665 ;
        RECT 49.870 24.645 50.035 24.665 ;
        RECT 49.405 24.615 49.575 24.645 ;
        RECT 49.400 24.505 49.575 24.615 ;
        RECT 49.405 24.455 49.575 24.505 ;
        RECT 49.865 24.475 50.035 24.645 ;
        RECT 52.630 24.475 52.800 24.665 ;
        RECT 54.925 24.455 55.095 24.645 ;
        RECT 56.305 24.475 56.475 24.665 ;
        RECT 58.600 24.505 58.720 24.615 ;
        RECT 59.070 24.455 59.240 24.645 ;
        RECT 59.525 24.475 59.695 24.665 ;
        RECT 59.985 24.475 60.155 24.665 ;
        RECT 64.585 24.475 64.755 24.645 ;
        RECT 65.505 24.475 65.675 24.665 ;
        RECT 64.585 24.455 64.750 24.475 ;
        RECT 68.265 24.455 68.435 24.645 ;
        RECT 68.730 24.455 68.900 24.645 ;
        RECT 71.025 24.475 71.195 24.665 ;
        RECT 75.630 24.645 75.795 24.665 ;
        RECT 74.245 24.475 74.415 24.645 ;
        RECT 74.245 24.455 74.410 24.475 ;
        RECT 74.705 24.455 74.875 24.645 ;
        RECT 75.625 24.475 75.795 24.645 ;
        RECT 76.540 24.505 76.660 24.615 ;
        RECT 78.390 24.475 78.560 24.665 ;
        RECT 79.765 24.455 79.935 24.645 ;
        RECT 82.065 24.475 82.235 24.665 ;
        RECT 83.445 24.645 83.615 24.665 ;
        RECT 83.440 24.475 83.615 24.645 ;
        RECT 83.440 24.455 83.610 24.475 ;
        RECT 83.905 24.455 84.075 24.645 ;
        RECT 85.285 24.455 85.455 24.645 ;
        RECT 87.125 24.455 87.295 24.645 ;
        RECT 90.345 24.455 90.515 24.645 ;
        RECT 91.725 24.455 91.895 24.665 ;
        RECT 13.385 23.645 14.755 24.455 ;
        RECT 14.765 23.775 16.595 24.455 ;
        RECT 14.765 23.545 16.110 23.775 ;
        RECT 16.605 23.645 17.975 24.455 ;
        RECT 17.985 23.775 19.815 24.455 ;
        RECT 19.825 23.775 21.655 24.455 ;
        RECT 17.985 23.545 19.330 23.775 ;
        RECT 19.825 23.545 21.170 23.775 ;
        RECT 22.585 23.545 25.795 24.455 ;
        RECT 25.805 23.775 27.635 24.455 ;
        RECT 28.710 23.775 30.545 24.455 ;
        RECT 26.290 23.545 27.635 23.775 ;
        RECT 29.615 23.545 30.545 23.775 ;
        RECT 30.865 23.645 36.375 24.455 ;
        RECT 36.385 23.645 39.135 24.455 ;
        RECT 39.155 23.585 39.585 24.370 ;
        RECT 39.605 23.645 41.435 24.455 ;
        RECT 41.445 23.545 44.655 24.455 ;
        RECT 44.665 23.645 46.035 24.455 ;
        RECT 46.045 23.545 49.255 24.455 ;
        RECT 49.265 23.645 54.775 24.455 ;
        RECT 54.785 23.645 58.455 24.455 ;
        RECT 58.925 23.545 62.400 24.455 ;
        RECT 62.915 23.775 64.750 24.455 ;
        RECT 62.915 23.545 63.845 23.775 ;
        RECT 64.915 23.585 65.345 24.370 ;
        RECT 65.365 23.545 68.575 24.455 ;
        RECT 68.585 23.545 72.060 24.455 ;
        RECT 72.575 23.775 74.410 24.455 ;
        RECT 72.575 23.545 73.505 23.775 ;
        RECT 74.565 23.645 76.395 24.455 ;
        RECT 76.865 23.545 80.075 24.455 ;
        RECT 80.280 23.545 83.755 24.455 ;
        RECT 83.765 23.645 85.135 24.455 ;
        RECT 85.145 23.775 86.975 24.455 ;
        RECT 86.985 23.775 88.815 24.455 ;
        RECT 85.630 23.545 86.975 23.775 ;
        RECT 87.470 23.545 88.815 23.775 ;
        RECT 88.825 23.775 90.655 24.455 ;
        RECT 88.825 23.545 90.170 23.775 ;
        RECT 90.665 23.645 92.035 24.455 ;
      LAYER nwell ;
        RECT 13.190 20.425 92.230 23.255 ;
      LAYER pwell ;
        RECT 13.385 19.225 14.755 20.035 ;
        RECT 15.225 19.225 18.700 20.135 ;
        RECT 19.825 19.905 21.170 20.135 ;
        RECT 19.825 19.225 21.655 19.905 ;
        RECT 21.665 19.225 25.140 20.135 ;
        RECT 26.275 19.310 26.705 20.095 ;
        RECT 27.380 19.225 30.855 20.135 ;
        RECT 31.060 19.225 34.535 20.135 ;
        RECT 38.060 19.905 38.970 20.125 ;
        RECT 40.505 19.905 41.855 20.135 ;
        RECT 34.545 19.225 41.855 19.905 ;
        RECT 42.825 19.225 46.300 20.135 ;
        RECT 46.505 19.225 48.335 20.035 ;
        RECT 48.345 19.225 51.820 20.135 ;
        RECT 52.035 19.310 52.465 20.095 ;
        RECT 52.485 19.225 54.315 20.035 ;
        RECT 54.785 19.225 58.260 20.135 ;
        RECT 61.980 19.905 62.890 20.125 ;
        RECT 64.425 19.905 65.775 20.135 ;
        RECT 69.340 19.905 70.250 20.125 ;
        RECT 71.785 19.905 73.135 20.135 ;
        RECT 58.465 19.225 65.775 19.905 ;
        RECT 65.825 19.225 73.135 19.905 ;
        RECT 73.185 19.225 76.660 20.135 ;
        RECT 77.795 19.310 78.225 20.095 ;
        RECT 78.900 19.225 82.375 20.135 ;
        RECT 82.580 19.225 86.055 20.135 ;
        RECT 86.550 19.905 87.895 20.135 ;
        RECT 88.390 19.905 89.735 20.135 ;
        RECT 86.065 19.225 87.895 19.905 ;
        RECT 87.905 19.225 89.735 19.905 ;
        RECT 90.665 19.225 92.035 20.035 ;
        RECT 13.525 19.015 13.695 19.225 ;
        RECT 14.900 19.170 15.020 19.175 ;
        RECT 14.900 19.065 15.075 19.170 ;
        RECT 14.915 19.060 15.075 19.065 ;
        RECT 15.370 19.035 15.540 19.225 ;
        RECT 15.825 19.035 15.995 19.205 ;
        RECT 15.830 19.015 15.995 19.035 ;
        RECT 18.125 19.015 18.295 19.205 ;
        RECT 19.055 19.070 19.215 19.180 ;
        RECT 19.505 19.015 19.675 19.205 ;
        RECT 21.345 19.035 21.515 19.225 ;
        RECT 21.810 19.035 21.980 19.225 ;
        RECT 25.495 19.070 25.655 19.180 ;
        RECT 26.865 19.175 27.035 19.205 ;
        RECT 26.860 19.065 27.035 19.175 ;
        RECT 26.865 19.035 27.035 19.065 ;
        RECT 26.870 19.015 27.035 19.035 ;
        RECT 29.165 19.015 29.335 19.205 ;
        RECT 30.540 19.035 30.710 19.225 ;
        RECT 34.220 19.035 34.390 19.225 ;
        RECT 34.685 19.035 34.855 19.225 ;
        RECT 38.365 19.035 38.535 19.205 ;
        RECT 38.820 19.065 38.940 19.175 ;
        RECT 39.740 19.065 39.860 19.175 ;
        RECT 42.055 19.070 42.215 19.180 ;
        RECT 42.970 19.035 43.140 19.225 ;
        RECT 46.645 19.035 46.815 19.225 ;
        RECT 38.365 19.015 38.530 19.035 ;
        RECT 47.105 19.015 47.275 19.205 ;
        RECT 47.560 19.065 47.680 19.175 ;
        RECT 48.025 19.015 48.195 19.205 ;
        RECT 48.490 19.035 48.660 19.225 ;
        RECT 52.625 19.035 52.795 19.225 ;
        RECT 54.460 19.065 54.580 19.175 ;
        RECT 54.930 19.035 55.100 19.225 ;
        RECT 55.385 19.015 55.555 19.205 ;
        RECT 58.605 19.035 58.775 19.225 ;
        RECT 64.585 19.035 64.755 19.205 ;
        RECT 65.965 19.035 66.135 19.225 ;
        RECT 64.585 19.015 64.750 19.035 ;
        RECT 68.265 19.015 68.435 19.205 ;
        RECT 68.725 19.015 68.895 19.205 ;
        RECT 70.105 19.015 70.275 19.205 ;
        RECT 73.330 19.035 73.500 19.225 ;
        RECT 77.015 19.070 77.175 19.180 ;
        RECT 77.465 19.035 77.635 19.205 ;
        RECT 78.380 19.065 78.500 19.175 ;
        RECT 77.470 19.015 77.635 19.035 ;
        RECT 79.765 19.015 79.935 19.205 ;
        RECT 81.145 19.015 81.315 19.205 ;
        RECT 82.060 19.035 82.230 19.225 ;
        RECT 85.740 19.035 85.910 19.225 ;
        RECT 86.205 19.035 86.375 19.225 ;
        RECT 88.045 19.035 88.215 19.225 ;
        RECT 88.505 19.015 88.675 19.205 ;
        RECT 89.895 19.070 90.055 19.180 ;
        RECT 90.340 19.065 90.460 19.175 ;
        RECT 91.725 19.015 91.895 19.225 ;
        RECT 13.385 18.205 14.755 19.015 ;
        RECT 15.830 18.335 17.665 19.015 ;
        RECT 16.735 18.105 17.665 18.335 ;
        RECT 17.985 18.205 19.355 19.015 ;
        RECT 19.365 18.335 26.675 19.015 ;
        RECT 26.870 18.335 28.705 19.015 ;
        RECT 29.025 18.335 36.335 19.015 ;
        RECT 22.880 18.115 23.790 18.335 ;
        RECT 25.325 18.105 26.675 18.335 ;
        RECT 27.775 18.105 28.705 18.335 ;
        RECT 32.540 18.115 33.450 18.335 ;
        RECT 34.985 18.105 36.335 18.335 ;
        RECT 36.695 18.335 38.530 19.015 ;
        RECT 36.695 18.105 37.625 18.335 ;
        RECT 39.155 18.145 39.585 18.930 ;
        RECT 40.105 18.335 47.415 19.015 ;
        RECT 47.885 18.335 55.195 19.015 ;
        RECT 55.245 18.335 62.555 19.015 ;
        RECT 40.105 18.105 41.455 18.335 ;
        RECT 42.990 18.115 43.900 18.335 ;
        RECT 51.400 18.115 52.310 18.335 ;
        RECT 53.845 18.105 55.195 18.335 ;
        RECT 58.760 18.115 59.670 18.335 ;
        RECT 61.205 18.105 62.555 18.335 ;
        RECT 62.915 18.335 64.750 19.015 ;
        RECT 62.915 18.105 63.845 18.335 ;
        RECT 64.915 18.145 65.345 18.930 ;
        RECT 65.365 18.105 68.575 19.015 ;
        RECT 68.585 18.205 69.955 19.015 ;
        RECT 69.965 18.335 77.275 19.015 ;
        RECT 77.470 18.335 79.305 19.015 ;
        RECT 73.480 18.115 74.390 18.335 ;
        RECT 75.925 18.105 77.275 18.335 ;
        RECT 78.375 18.105 79.305 18.335 ;
        RECT 79.625 18.205 80.995 19.015 ;
        RECT 81.005 18.335 88.315 19.015 ;
        RECT 88.365 18.335 90.195 19.015 ;
        RECT 84.520 18.115 85.430 18.335 ;
        RECT 86.965 18.105 88.315 18.335 ;
        RECT 88.850 18.105 90.195 18.335 ;
        RECT 90.665 18.205 92.035 19.015 ;
      LAYER nwell ;
        RECT 13.190 14.985 92.230 17.815 ;
      LAYER pwell ;
        RECT 13.385 13.785 14.755 14.595 ;
        RECT 18.280 14.465 19.190 14.685 ;
        RECT 20.725 14.465 22.075 14.695 ;
        RECT 14.765 13.785 22.075 14.465 ;
        RECT 23.355 14.465 24.285 14.695 ;
        RECT 23.355 13.785 25.190 14.465 ;
        RECT 26.275 13.870 26.705 14.655 ;
        RECT 27.645 14.465 28.990 14.695 ;
        RECT 29.945 14.465 31.290 14.695 ;
        RECT 31.785 14.465 33.130 14.695 ;
        RECT 33.625 14.465 34.970 14.695 ;
        RECT 35.465 14.465 36.810 14.695 ;
        RECT 37.305 14.465 38.650 14.695 ;
        RECT 27.645 13.785 29.475 14.465 ;
        RECT 29.945 13.785 31.775 14.465 ;
        RECT 31.785 13.785 33.615 14.465 ;
        RECT 33.625 13.785 35.455 14.465 ;
        RECT 35.465 13.785 37.295 14.465 ;
        RECT 37.305 13.785 39.135 14.465 ;
        RECT 39.155 13.870 39.585 14.655 ;
        RECT 40.525 13.785 43.735 14.695 ;
        RECT 44.795 14.465 45.725 14.695 ;
        RECT 43.890 13.785 45.725 14.465 ;
        RECT 46.045 14.465 47.390 14.695 ;
        RECT 48.370 14.465 49.715 14.695 ;
        RECT 50.775 14.465 51.705 14.695 ;
        RECT 46.045 13.785 47.875 14.465 ;
        RECT 47.885 13.785 49.715 14.465 ;
        RECT 49.870 13.785 51.705 14.465 ;
        RECT 52.035 13.870 52.465 14.655 ;
        RECT 53.405 14.465 54.750 14.695 ;
        RECT 53.405 13.785 55.235 14.465 ;
        RECT 55.245 13.785 56.615 14.595 ;
        RECT 56.625 14.465 57.970 14.695 ;
        RECT 56.625 13.785 58.455 14.465 ;
        RECT 58.465 13.785 59.835 14.595 ;
        RECT 60.330 14.465 61.675 14.695 ;
        RECT 59.845 13.785 61.675 14.465 ;
        RECT 61.685 13.785 63.055 14.595 ;
        RECT 63.065 14.465 64.410 14.695 ;
        RECT 63.065 13.785 64.895 14.465 ;
        RECT 64.915 13.870 65.345 14.655 ;
        RECT 66.285 14.465 67.630 14.695 ;
        RECT 66.285 13.785 68.115 14.465 ;
        RECT 68.125 13.785 69.495 14.595 ;
        RECT 69.505 14.465 70.850 14.695 ;
        RECT 69.505 13.785 71.335 14.465 ;
        RECT 71.345 13.785 72.715 14.595 ;
        RECT 73.210 14.465 74.555 14.695 ;
        RECT 72.725 13.785 74.555 14.465 ;
        RECT 74.565 13.785 75.935 14.595 ;
        RECT 75.945 14.465 77.290 14.695 ;
        RECT 75.945 13.785 77.775 14.465 ;
        RECT 77.795 13.870 78.225 14.655 ;
        RECT 79.295 14.465 80.225 14.695 ;
        RECT 81.595 14.465 82.525 14.695 ;
        RECT 86.820 14.465 87.730 14.685 ;
        RECT 89.265 14.465 90.615 14.695 ;
        RECT 78.390 13.785 80.225 14.465 ;
        RECT 80.690 13.785 82.525 14.465 ;
        RECT 83.305 13.785 90.615 14.465 ;
        RECT 90.665 13.785 92.035 14.595 ;
        RECT 13.525 13.595 13.695 13.785 ;
        RECT 14.905 13.595 15.075 13.785 ;
        RECT 25.025 13.765 25.190 13.785 ;
        RECT 22.275 13.630 22.435 13.740 ;
        RECT 25.025 13.595 25.195 13.765 ;
        RECT 25.495 13.630 25.655 13.740 ;
        RECT 26.875 13.630 27.035 13.740 ;
        RECT 29.165 13.595 29.335 13.785 ;
        RECT 29.620 13.625 29.740 13.735 ;
        RECT 31.465 13.595 31.635 13.785 ;
        RECT 33.305 13.595 33.475 13.785 ;
        RECT 35.145 13.595 35.315 13.785 ;
        RECT 36.985 13.595 37.155 13.785 ;
        RECT 38.825 13.595 38.995 13.785 ;
        RECT 39.755 13.630 39.915 13.740 ;
        RECT 40.665 13.595 40.835 13.785 ;
        RECT 43.890 13.765 44.055 13.785 ;
        RECT 43.885 13.595 44.055 13.765 ;
        RECT 47.565 13.595 47.735 13.785 ;
        RECT 48.025 13.595 48.195 13.785 ;
        RECT 49.870 13.765 50.035 13.785 ;
        RECT 49.865 13.595 50.035 13.765 ;
        RECT 52.635 13.630 52.795 13.740 ;
        RECT 54.925 13.595 55.095 13.785 ;
        RECT 55.385 13.595 55.555 13.785 ;
        RECT 58.145 13.595 58.315 13.785 ;
        RECT 58.605 13.595 58.775 13.785 ;
        RECT 59.985 13.595 60.155 13.785 ;
        RECT 61.825 13.595 61.995 13.785 ;
        RECT 64.585 13.595 64.755 13.785 ;
        RECT 65.515 13.630 65.675 13.740 ;
        RECT 67.805 13.595 67.975 13.785 ;
        RECT 68.265 13.595 68.435 13.785 ;
        RECT 71.025 13.595 71.195 13.785 ;
        RECT 71.485 13.595 71.655 13.785 ;
        RECT 72.865 13.595 73.035 13.785 ;
        RECT 74.705 13.595 74.875 13.785 ;
        RECT 77.465 13.595 77.635 13.785 ;
        RECT 78.390 13.765 78.555 13.785 ;
        RECT 80.690 13.765 80.855 13.785 ;
        RECT 78.385 13.595 78.555 13.765 ;
        RECT 80.685 13.595 80.855 13.765 ;
        RECT 82.980 13.625 83.100 13.735 ;
        RECT 83.445 13.595 83.615 13.785 ;
        RECT 91.725 13.595 91.895 13.785 ;
      LAYER li1 ;
        RECT 112.275 219.210 112.445 219.295 ;
        RECT 114.995 219.210 115.165 219.295 ;
        RECT 117.715 219.210 117.885 219.295 ;
        RECT 120.435 219.210 120.605 219.295 ;
        RECT 123.155 219.210 123.325 219.295 ;
        RECT 125.875 219.210 126.045 219.295 ;
        RECT 128.595 219.210 128.765 219.295 ;
        RECT 131.315 219.210 131.485 219.295 ;
        RECT 134.035 219.210 134.205 219.295 ;
        RECT 136.755 219.210 136.925 219.295 ;
        RECT 139.475 219.210 139.645 219.295 ;
        RECT 142.195 219.210 142.365 219.295 ;
        RECT 144.915 219.210 145.085 219.295 ;
        RECT 147.635 219.210 147.805 219.295 ;
        RECT 112.275 218.690 113.735 219.210 ;
        RECT 112.275 218.000 113.195 218.690 ;
        RECT 113.905 218.520 116.255 219.210 ;
        RECT 116.425 218.690 119.175 219.210 ;
        RECT 113.365 218.000 116.795 218.520 ;
        RECT 116.965 218.000 118.635 218.690 ;
        RECT 119.345 218.520 121.695 219.210 ;
        RECT 121.865 218.690 124.615 219.210 ;
        RECT 118.805 218.000 122.235 218.520 ;
        RECT 122.405 218.000 124.075 218.690 ;
        RECT 124.785 218.520 127.135 219.210 ;
        RECT 127.305 218.690 130.055 219.210 ;
        RECT 124.245 218.000 127.675 218.520 ;
        RECT 127.845 218.000 129.515 218.690 ;
        RECT 130.225 218.520 132.575 219.210 ;
        RECT 132.745 218.690 135.495 219.210 ;
        RECT 129.685 218.000 133.115 218.520 ;
        RECT 133.285 218.000 134.955 218.690 ;
        RECT 135.665 218.520 138.015 219.210 ;
        RECT 138.185 218.690 140.935 219.210 ;
        RECT 135.125 218.000 138.555 218.520 ;
        RECT 138.725 218.000 140.395 218.690 ;
        RECT 141.105 218.520 143.455 219.210 ;
        RECT 143.625 218.690 146.375 219.210 ;
        RECT 140.565 218.000 143.995 218.520 ;
        RECT 144.165 218.000 145.835 218.690 ;
        RECT 146.545 218.520 147.805 219.210 ;
        RECT 146.005 218.000 147.805 218.520 ;
        RECT 112.275 217.830 112.445 218.000 ;
        RECT 114.995 217.830 115.165 218.000 ;
        RECT 112.275 216.245 112.990 217.830 ;
        RECT 114.560 217.825 115.165 217.830 ;
        RECT 117.715 217.825 117.885 218.000 ;
        RECT 114.560 217.565 116.315 217.825 ;
        RECT 116.875 217.565 117.885 217.825 ;
        RECT 118.540 217.780 119.375 217.830 ;
        RECT 114.560 216.965 115.165 217.565 ;
        RECT 115.335 217.220 117.545 217.390 ;
        RECT 115.335 217.135 116.240 217.220 ;
        RECT 116.970 217.135 117.545 217.220 ;
        RECT 117.715 217.280 117.885 217.565 ;
        RECT 118.105 217.770 119.375 217.780 ;
        RECT 120.435 217.825 120.605 218.000 ;
        RECT 123.155 217.825 123.325 218.000 ;
        RECT 125.875 217.825 126.045 218.000 ;
        RECT 128.595 217.830 128.765 218.000 ;
        RECT 131.315 217.830 131.485 218.000 ;
        RECT 128.595 217.825 130.055 217.830 ;
        RECT 118.105 217.660 120.220 217.770 ;
        RECT 118.105 217.605 118.665 217.660 ;
        RECT 119.245 217.615 120.220 217.660 ;
        RECT 118.105 217.450 118.625 217.605 ;
        RECT 117.715 217.110 118.495 217.280 ;
        RECT 116.475 216.965 116.805 217.050 ;
        RECT 117.715 216.965 117.885 217.110 ;
        RECT 114.560 216.635 115.925 216.965 ;
        RECT 116.095 216.795 117.165 216.965 ;
        RECT 112.275 215.905 113.820 216.245 ;
        RECT 112.275 212.485 112.990 215.905 ;
        RECT 114.560 214.560 115.165 216.635 ;
        RECT 116.095 216.420 116.265 216.795 ;
        RECT 115.335 216.250 116.265 216.420 ;
        RECT 116.445 216.160 116.815 216.515 ;
        RECT 116.995 216.420 117.165 216.795 ;
        RECT 117.335 216.635 117.885 216.965 ;
        RECT 118.795 216.940 119.125 217.490 ;
        RECT 119.295 217.440 120.220 217.615 ;
        RECT 120.435 217.565 121.755 217.825 ;
        RECT 122.315 217.565 123.325 217.825 ;
        RECT 123.585 217.570 124.045 217.740 ;
        RECT 120.435 217.270 120.605 217.565 ;
        RECT 123.155 217.400 123.325 217.565 ;
        RECT 119.425 217.100 120.605 217.270 ;
        RECT 120.775 217.220 122.985 217.390 ;
        RECT 120.775 217.135 121.680 217.220 ;
        RECT 122.410 217.135 122.985 217.220 ;
        RECT 116.995 216.250 117.545 216.420 ;
        RECT 117.715 216.350 117.885 216.635 ;
        RECT 118.100 216.930 119.125 216.940 ;
        RECT 120.435 216.965 120.605 217.100 ;
        RECT 123.155 217.070 123.705 217.400 ;
        RECT 123.875 217.305 124.045 217.570 ;
        RECT 124.215 217.475 124.865 217.825 ;
        RECT 125.035 217.570 125.705 217.740 ;
        RECT 125.035 217.305 125.205 217.570 ;
        RECT 125.875 217.565 127.195 217.825 ;
        RECT 127.755 217.565 130.055 217.825 ;
        RECT 125.875 217.400 126.045 217.565 ;
        RECT 123.875 217.075 125.205 217.305 ;
        RECT 125.375 217.070 126.045 217.400 ;
        RECT 126.215 217.220 128.425 217.390 ;
        RECT 126.215 217.135 127.120 217.220 ;
        RECT 127.850 217.135 128.425 217.220 ;
        RECT 128.595 217.310 130.055 217.565 ;
        RECT 121.915 216.965 122.245 217.050 ;
        RECT 123.155 216.965 123.325 217.070 ;
        RECT 118.100 216.740 120.265 216.930 ;
        RECT 118.100 216.610 118.625 216.740 ;
        RECT 119.330 216.590 120.265 216.740 ;
        RECT 120.435 216.635 121.365 216.965 ;
        RECT 121.535 216.795 122.605 216.965 ;
        RECT 117.715 216.140 118.415 216.350 ;
        RECT 115.335 214.895 117.545 215.065 ;
        RECT 115.335 214.730 116.305 214.895 ;
        RECT 116.975 214.810 117.545 214.895 ;
        RECT 116.475 214.640 116.805 214.725 ;
        RECT 117.715 214.640 117.885 216.140 ;
        RECT 118.795 215.865 119.125 216.570 ;
        RECT 119.330 216.035 119.705 216.590 ;
        RECT 120.435 216.360 120.605 216.635 ;
        RECT 121.535 216.420 121.705 216.795 ;
        RECT 119.935 216.045 120.605 216.360 ;
        RECT 120.775 216.250 121.705 216.420 ;
        RECT 121.885 216.160 122.255 216.515 ;
        RECT 122.435 216.420 122.605 216.795 ;
        RECT 122.775 216.635 123.325 216.965 ;
        RECT 125.875 216.965 126.045 217.070 ;
        RECT 127.355 216.965 127.685 217.050 ;
        RECT 128.595 216.965 129.515 217.310 ;
        RECT 130.225 217.270 131.485 217.830 ;
        RECT 132.545 217.780 133.380 217.830 ;
        RECT 132.545 217.770 133.815 217.780 ;
        RECT 131.700 217.660 133.815 217.770 ;
        RECT 131.700 217.615 132.675 217.660 ;
        RECT 131.700 217.440 132.625 217.615 ;
        RECT 133.255 217.605 133.815 217.660 ;
        RECT 130.225 217.140 132.495 217.270 ;
        RECT 123.585 216.715 125.705 216.900 ;
        RECT 123.155 216.460 123.325 216.635 ;
        RECT 125.875 216.635 126.805 216.965 ;
        RECT 126.975 216.795 128.045 216.965 ;
        RECT 122.435 216.250 122.985 216.420 ;
        RECT 123.155 216.210 123.785 216.460 ;
        RECT 123.955 216.265 124.905 216.545 ;
        RECT 125.875 216.475 126.045 216.635 ;
        RECT 125.415 216.210 126.045 216.475 ;
        RECT 126.975 216.420 127.145 216.795 ;
        RECT 126.215 216.250 127.145 216.420 ;
        RECT 118.165 215.695 120.135 215.865 ;
        RECT 118.165 215.080 118.335 215.695 ;
        RECT 118.505 215.205 119.795 215.525 ;
        RECT 118.505 215.060 118.835 215.205 ;
        RECT 114.560 214.425 116.305 214.560 ;
        RECT 116.475 214.470 117.145 214.640 ;
        RECT 113.310 214.390 116.305 214.425 ;
        RECT 113.310 214.075 115.165 214.390 ;
        RECT 116.475 214.220 116.805 214.245 ;
        RECT 114.560 212.485 115.165 214.075 ;
        RECT 112.275 212.310 112.445 212.485 ;
        RECT 114.995 212.310 115.165 212.485 ;
        RECT 112.275 210.660 113.735 212.310 ;
        RECT 113.905 212.020 115.165 212.310 ;
        RECT 115.335 214.050 116.805 214.220 ;
        RECT 115.335 212.360 115.505 214.050 ;
        RECT 116.975 213.885 117.145 214.470 ;
        RECT 117.315 214.325 117.885 214.640 ;
        RECT 118.165 214.675 118.335 214.910 ;
        RECT 119.045 214.845 119.765 215.035 ;
        RECT 119.965 214.980 120.135 215.695 ;
        RECT 119.935 214.675 120.265 214.755 ;
        RECT 118.165 214.505 120.265 214.675 ;
        RECT 117.315 214.310 118.385 214.325 ;
        RECT 117.715 213.955 118.385 214.310 ;
        RECT 118.565 214.045 118.865 214.505 ;
        RECT 120.435 214.500 120.605 216.045 ;
        RECT 120.775 214.670 121.455 214.955 ;
        RECT 120.435 214.335 121.065 214.500 ;
        RECT 119.045 214.165 119.375 214.335 ;
        RECT 119.635 214.230 121.065 214.335 ;
        RECT 119.635 214.165 120.605 214.230 ;
        RECT 116.975 213.880 117.545 213.885 ;
        RECT 115.675 213.710 117.545 213.880 ;
        RECT 115.675 212.755 115.845 213.710 ;
        RECT 116.015 213.370 116.985 213.540 ;
        RECT 116.015 212.720 116.185 213.370 ;
        RECT 117.180 213.355 117.545 213.710 ;
        RECT 117.205 213.165 117.375 213.170 ;
        RECT 116.385 212.890 117.545 213.165 ;
        RECT 116.015 212.530 117.545 212.720 ;
        RECT 115.335 212.190 116.360 212.360 ;
        RECT 117.715 212.350 117.885 213.955 ;
        RECT 118.565 213.845 118.895 214.045 ;
        RECT 119.115 213.995 119.375 214.165 ;
        RECT 119.115 213.825 120.160 213.995 ;
        RECT 119.115 213.635 119.285 213.825 ;
        RECT 118.165 213.465 119.285 213.635 ;
        RECT 118.165 212.960 118.335 213.465 ;
        RECT 119.455 213.295 119.820 213.655 ;
        RECT 118.535 213.125 119.820 213.295 ;
        RECT 118.535 212.770 118.755 213.125 ;
        RECT 118.165 212.600 118.335 212.765 ;
        RECT 118.925 212.715 119.520 212.955 ;
        RECT 119.990 212.890 120.160 213.825 ;
        RECT 118.165 212.545 118.605 212.600 ;
        RECT 119.710 212.545 120.265 212.680 ;
        RECT 118.165 212.430 120.265 212.545 ;
        RECT 120.435 212.440 120.605 214.165 ;
        RECT 121.235 214.210 121.455 214.670 ;
        RECT 121.625 214.380 122.185 215.070 ;
        RECT 122.355 214.670 122.985 214.955 ;
        RECT 122.355 214.210 122.525 214.670 ;
        RECT 123.155 214.515 123.325 216.210 ;
        RECT 123.915 216.040 125.280 216.095 ;
        RECT 123.605 215.925 125.705 216.040 ;
        RECT 123.605 215.870 124.045 215.925 ;
        RECT 123.605 215.705 123.775 215.870 ;
        RECT 125.150 215.790 125.705 215.925 ;
        RECT 123.605 215.005 123.775 215.510 ;
        RECT 123.975 215.345 124.195 215.700 ;
        RECT 124.365 215.515 124.960 215.755 ;
        RECT 123.975 215.175 125.260 215.345 ;
        RECT 123.605 214.835 124.725 215.005 ;
        RECT 124.555 214.645 124.725 214.835 ;
        RECT 124.895 214.815 125.260 215.175 ;
        RECT 125.430 214.645 125.600 215.580 ;
        RECT 123.155 214.500 123.825 214.515 ;
        RECT 122.695 214.230 123.825 214.500 ;
        RECT 121.235 214.000 122.525 214.210 ;
        RECT 123.155 214.145 123.825 214.230 ;
        RECT 124.005 214.425 124.335 214.625 ;
        RECT 124.555 214.475 125.600 214.645 ;
        RECT 125.875 215.020 126.045 216.210 ;
        RECT 127.325 216.160 127.695 216.515 ;
        RECT 127.875 216.420 128.045 216.795 ;
        RECT 128.215 216.635 129.515 216.965 ;
        RECT 128.595 216.620 129.515 216.635 ;
        RECT 129.685 217.100 132.495 217.140 ;
        RECT 129.685 216.620 131.485 217.100 ;
        RECT 132.795 216.940 133.125 217.490 ;
        RECT 133.295 217.450 133.815 217.605 ;
        RECT 134.035 217.400 134.205 218.000 ;
        RECT 136.755 217.825 136.925 218.000 ;
        RECT 139.475 217.825 139.645 218.000 ;
        RECT 142.195 217.830 142.365 218.000 ;
        RECT 144.915 217.830 145.085 218.000 ;
        RECT 147.635 217.830 147.805 218.000 ;
        RECT 134.375 217.655 136.585 217.825 ;
        RECT 134.375 217.570 134.945 217.655 ;
        RECT 135.615 217.490 136.585 217.655 ;
        RECT 136.755 217.565 138.075 217.825 ;
        RECT 138.635 217.565 139.645 217.825 ;
        RECT 139.905 217.570 140.365 217.740 ;
        RECT 135.115 217.400 135.445 217.485 ;
        RECT 134.035 217.280 134.605 217.400 ;
        RECT 133.425 217.110 134.605 217.280 ;
        RECT 134.035 217.070 134.605 217.110 ;
        RECT 134.775 217.230 135.445 217.400 ;
        RECT 136.755 217.320 136.925 217.565 ;
        RECT 139.475 217.400 139.645 217.565 ;
        RECT 132.795 216.930 133.820 216.940 ;
        RECT 127.875 216.250 128.425 216.420 ;
        RECT 128.595 215.880 128.765 216.620 ;
        RECT 128.935 216.050 129.565 216.335 ;
        RECT 128.595 215.610 129.225 215.880 ;
        RECT 126.215 215.355 128.425 215.525 ;
        RECT 126.215 215.190 127.185 215.355 ;
        RECT 127.855 215.270 128.425 215.355 ;
        RECT 127.355 215.100 127.685 215.185 ;
        RECT 128.595 215.100 128.765 215.610 ;
        RECT 129.395 215.590 129.565 216.050 ;
        RECT 129.735 215.760 130.295 216.450 ;
        RECT 131.315 216.360 131.485 216.620 ;
        RECT 131.655 216.740 133.820 216.930 ;
        RECT 131.655 216.590 132.590 216.740 ;
        RECT 133.295 216.610 133.820 216.740 ;
        RECT 130.465 216.050 131.145 216.335 ;
        RECT 130.465 215.590 130.685 216.050 ;
        RECT 131.315 216.045 131.985 216.360 ;
        RECT 131.315 215.880 131.485 216.045 ;
        RECT 132.215 216.035 132.590 216.590 ;
        RECT 130.855 215.610 131.485 215.880 ;
        RECT 132.795 215.865 133.125 216.570 ;
        RECT 134.035 216.350 134.205 217.070 ;
        RECT 134.775 216.645 134.945 217.230 ;
        RECT 135.615 217.150 136.925 217.320 ;
        RECT 135.115 216.980 135.445 217.005 ;
        RECT 135.115 216.810 136.585 216.980 ;
        RECT 133.505 216.140 134.205 216.350 ;
        RECT 129.395 215.380 130.685 215.590 ;
        RECT 125.875 214.850 127.185 215.020 ;
        RECT 127.355 214.930 128.025 215.100 ;
        RECT 120.775 213.430 122.985 213.830 ;
        RECT 120.775 212.960 121.455 213.240 ;
        RECT 121.235 212.565 121.455 212.960 ;
        RECT 121.625 212.735 122.185 213.430 ;
        RECT 122.355 212.960 122.985 213.240 ;
        RECT 122.355 212.565 122.525 212.960 ;
        RECT 118.475 212.375 119.840 212.430 ;
        RECT 113.905 211.850 115.925 212.020 ;
        RECT 113.905 210.930 115.165 211.850 ;
        RECT 115.515 211.440 115.925 211.615 ;
        RECT 116.170 211.610 116.360 212.190 ;
        RECT 116.735 211.620 116.905 212.330 ;
        RECT 117.180 212.260 117.885 212.350 ;
        RECT 120.435 212.260 121.065 212.440 ;
        RECT 117.180 212.010 118.345 212.260 ;
        RECT 117.180 211.840 117.885 212.010 ;
        RECT 118.515 211.925 119.465 212.205 ;
        RECT 119.975 212.115 121.065 212.260 ;
        RECT 121.235 212.115 122.525 212.565 ;
        RECT 123.155 212.440 123.325 214.145 ;
        RECT 124.005 213.965 124.305 214.425 ;
        RECT 124.555 214.305 124.815 214.475 ;
        RECT 125.875 214.305 126.045 214.850 ;
        RECT 127.355 214.680 127.685 214.705 ;
        RECT 124.485 214.135 124.815 214.305 ;
        RECT 125.075 214.135 126.045 214.305 ;
        RECT 123.605 213.795 125.705 213.965 ;
        RECT 123.605 213.560 123.775 213.795 ;
        RECT 125.375 213.715 125.705 213.795 ;
        RECT 124.485 213.435 125.205 213.625 ;
        RECT 123.605 212.775 123.775 213.390 ;
        RECT 123.945 213.265 124.275 213.410 ;
        RECT 123.945 212.945 125.235 213.265 ;
        RECT 125.405 212.775 125.575 213.490 ;
        RECT 123.605 212.605 125.575 212.775 ;
        RECT 122.695 212.330 123.325 212.440 ;
        RECT 122.695 212.120 123.855 212.330 ;
        RECT 122.695 212.115 123.325 212.120 ;
        RECT 119.975 211.995 120.605 212.115 ;
        RECT 121.915 212.010 122.245 212.115 ;
        RECT 116.735 211.440 117.510 211.620 ;
        RECT 115.515 211.375 117.510 211.440 ;
        RECT 117.715 211.400 117.885 211.840 ;
        RECT 118.145 211.570 120.265 211.755 ;
        RECT 120.435 211.400 120.605 211.995 ;
        RECT 120.775 211.840 121.745 211.945 ;
        RECT 122.415 211.840 122.985 211.945 ;
        RECT 120.775 211.560 122.985 211.840 ;
        RECT 115.515 211.100 116.905 211.375 ;
        RECT 117.715 211.070 118.265 211.400 ;
        RECT 118.435 211.165 119.765 211.395 ;
        RECT 117.715 210.930 117.885 211.070 ;
        RECT 112.275 208.800 113.215 210.660 ;
        RECT 113.905 210.490 116.255 210.930 ;
        RECT 113.385 209.110 116.255 210.490 ;
        RECT 116.425 210.470 117.885 210.930 ;
        RECT 118.435 210.900 118.605 211.165 ;
        RECT 118.145 210.730 118.605 210.900 ;
        RECT 118.775 210.645 119.425 210.995 ;
        RECT 119.595 210.900 119.765 211.165 ;
        RECT 119.935 211.070 120.605 211.400 ;
        RECT 119.595 210.730 120.265 210.900 ;
        RECT 120.435 210.470 120.605 211.070 ;
        RECT 123.155 211.360 123.325 212.115 ;
        RECT 124.235 211.900 124.565 212.605 ;
        RECT 125.875 212.480 126.045 214.135 ;
        RECT 126.215 214.510 127.685 214.680 ;
        RECT 126.215 212.820 126.385 214.510 ;
        RECT 127.855 214.345 128.025 214.930 ;
        RECT 128.195 214.770 128.765 215.100 ;
        RECT 128.935 214.810 131.145 215.210 ;
        RECT 127.855 214.340 128.425 214.345 ;
        RECT 126.555 214.170 128.425 214.340 ;
        RECT 126.555 213.215 126.725 214.170 ;
        RECT 126.895 213.830 127.865 214.000 ;
        RECT 126.895 213.180 127.065 213.830 ;
        RECT 128.060 213.815 128.425 214.170 ;
        RECT 128.595 213.820 128.765 214.770 ;
        RECT 128.935 214.340 129.565 214.620 ;
        RECT 129.395 213.945 129.565 214.340 ;
        RECT 129.735 214.115 130.295 214.810 ;
        RECT 130.465 214.340 131.145 214.620 ;
        RECT 130.465 213.945 130.685 214.340 ;
        RECT 128.085 213.625 128.255 213.630 ;
        RECT 127.265 213.350 128.425 213.625 ;
        RECT 128.595 213.495 129.225 213.820 ;
        RECT 129.395 213.495 130.685 213.945 ;
        RECT 131.315 214.335 131.485 215.610 ;
        RECT 131.785 215.695 133.755 215.865 ;
        RECT 131.785 214.980 131.955 215.695 ;
        RECT 132.125 215.205 133.415 215.525 ;
        RECT 133.085 215.060 133.415 215.205 ;
        RECT 133.585 215.080 133.755 215.695 ;
        RECT 134.035 215.110 134.205 216.140 ;
        RECT 134.375 216.640 134.945 216.645 ;
        RECT 134.375 216.470 136.245 216.640 ;
        RECT 134.375 216.115 134.740 216.470 ;
        RECT 134.935 216.130 135.905 216.300 ;
        RECT 134.545 215.925 134.715 215.930 ;
        RECT 134.375 215.650 135.535 215.925 ;
        RECT 135.735 215.480 135.905 216.130 ;
        RECT 136.075 215.515 136.245 216.470 ;
        RECT 134.375 215.290 135.905 215.480 ;
        RECT 136.415 215.120 136.585 216.810 ;
        RECT 132.155 214.845 132.875 215.035 ;
        RECT 131.655 214.675 131.985 214.755 ;
        RECT 133.585 214.675 133.755 214.910 ;
        RECT 131.655 214.505 133.755 214.675 ;
        RECT 134.035 214.600 134.740 215.110 ;
        RECT 131.315 214.165 132.285 214.335 ;
        RECT 132.545 214.165 132.875 214.335 ;
        RECT 131.315 213.820 131.485 214.165 ;
        RECT 132.545 213.995 132.805 214.165 ;
        RECT 133.055 214.045 133.355 214.505 ;
        RECT 134.035 214.325 134.205 214.600 ;
        RECT 135.015 214.380 135.185 215.090 ;
        RECT 130.855 213.495 131.485 213.820 ;
        RECT 126.895 212.990 128.425 213.180 ;
        RECT 126.215 212.650 127.240 212.820 ;
        RECT 128.595 212.810 128.765 213.495 ;
        RECT 129.675 213.390 130.005 213.495 ;
        RECT 128.935 213.220 129.505 213.325 ;
        RECT 130.175 213.220 131.145 213.325 ;
        RECT 128.935 212.940 131.145 213.220 ;
        RECT 124.770 211.880 125.145 212.435 ;
        RECT 125.875 212.425 126.805 212.480 ;
        RECT 125.375 212.310 126.805 212.425 ;
        RECT 125.375 212.110 126.045 212.310 ;
        RECT 123.540 211.730 124.065 211.860 ;
        RECT 124.770 211.730 125.705 211.880 ;
        RECT 123.540 211.540 125.705 211.730 ;
        RECT 123.540 211.530 124.565 211.540 ;
        RECT 123.155 211.190 123.935 211.360 ;
        RECT 123.155 210.470 123.325 211.190 ;
        RECT 123.545 210.865 124.065 211.020 ;
        RECT 124.235 210.980 124.565 211.530 ;
        RECT 125.875 211.370 126.045 212.110 ;
        RECT 126.395 211.900 126.805 212.075 ;
        RECT 127.050 212.070 127.240 212.650 ;
        RECT 127.615 212.080 127.785 212.790 ;
        RECT 128.060 212.300 128.765 212.810 ;
        RECT 128.935 212.490 131.145 212.770 ;
        RECT 128.935 212.385 129.505 212.490 ;
        RECT 130.175 212.385 131.145 212.490 ;
        RECT 128.595 212.215 128.765 212.300 ;
        RECT 129.675 212.215 130.005 212.320 ;
        RECT 131.315 212.260 131.485 213.495 ;
        RECT 131.760 213.825 132.805 213.995 ;
        RECT 133.025 213.845 133.355 214.045 ;
        RECT 133.535 213.955 134.205 214.325 ;
        RECT 134.410 214.200 135.185 214.380 ;
        RECT 135.560 214.950 136.585 215.120 ;
        RECT 136.755 216.965 136.925 217.150 ;
        RECT 137.095 217.220 139.305 217.390 ;
        RECT 137.095 217.135 138.000 217.220 ;
        RECT 138.730 217.135 139.305 217.220 ;
        RECT 139.475 217.070 140.025 217.400 ;
        RECT 140.195 217.305 140.365 217.570 ;
        RECT 140.535 217.475 141.185 217.825 ;
        RECT 141.355 217.570 142.025 217.740 ;
        RECT 141.355 217.305 141.525 217.570 ;
        RECT 142.195 217.400 143.455 217.830 ;
        RECT 140.195 217.075 141.525 217.305 ;
        RECT 141.695 217.070 143.455 217.400 ;
        RECT 138.235 216.965 138.565 217.050 ;
        RECT 139.475 216.965 139.645 217.070 ;
        RECT 136.755 216.635 137.685 216.965 ;
        RECT 137.855 216.795 138.925 216.965 ;
        RECT 136.755 215.480 136.925 216.635 ;
        RECT 137.855 216.420 138.025 216.795 ;
        RECT 137.095 216.250 138.025 216.420 ;
        RECT 138.205 216.160 138.575 216.515 ;
        RECT 138.755 216.420 138.925 216.795 ;
        RECT 139.095 216.635 139.645 216.965 ;
        RECT 139.905 216.715 142.025 216.900 ;
        RECT 139.475 216.460 139.645 216.635 ;
        RECT 138.755 216.250 139.305 216.420 ;
        RECT 139.475 216.210 140.105 216.460 ;
        RECT 140.275 216.265 141.225 216.545 ;
        RECT 142.195 216.475 143.455 217.070 ;
        RECT 141.735 216.210 143.455 216.475 ;
        RECT 137.095 215.815 139.305 215.985 ;
        RECT 137.095 215.650 138.065 215.815 ;
        RECT 138.735 215.730 139.305 215.815 ;
        RECT 138.235 215.560 138.565 215.645 ;
        RECT 139.475 215.560 139.645 216.210 ;
        RECT 140.235 216.040 141.600 216.095 ;
        RECT 139.925 215.925 142.025 216.040 ;
        RECT 139.925 215.870 140.365 215.925 ;
        RECT 139.925 215.705 140.095 215.870 ;
        RECT 141.470 215.790 142.025 215.925 ;
        RECT 142.195 216.010 143.455 216.210 ;
        RECT 143.625 216.245 145.630 217.830 ;
        RECT 143.625 216.180 146.460 216.245 ;
        RECT 136.755 215.310 138.065 215.480 ;
        RECT 138.235 215.390 138.905 215.560 ;
        RECT 135.560 214.370 135.750 214.950 ;
        RECT 136.755 214.780 136.925 215.310 ;
        RECT 138.235 215.140 138.565 215.165 ;
        RECT 135.995 214.610 136.925 214.780 ;
        RECT 135.995 214.200 136.405 214.375 ;
        RECT 134.410 214.135 136.405 214.200 ;
        RECT 131.760 212.890 131.930 213.825 ;
        RECT 132.100 213.295 132.465 213.655 ;
        RECT 132.635 213.635 132.805 213.825 ;
        RECT 132.635 213.465 133.755 213.635 ;
        RECT 132.100 213.125 133.385 213.295 ;
        RECT 132.400 212.715 132.995 212.955 ;
        RECT 133.165 212.770 133.385 213.125 ;
        RECT 133.585 212.960 133.755 213.465 ;
        RECT 134.035 213.260 134.205 213.955 ;
        RECT 135.015 213.860 136.405 214.135 ;
        RECT 134.465 213.430 134.925 213.600 ;
        RECT 134.035 212.930 134.585 213.260 ;
        RECT 134.755 213.165 134.925 213.430 ;
        RECT 135.095 213.335 135.745 213.685 ;
        RECT 135.915 213.430 136.585 213.600 ;
        RECT 135.915 213.165 136.085 213.430 ;
        RECT 136.755 213.260 136.925 214.610 ;
        RECT 134.755 212.935 136.085 213.165 ;
        RECT 136.255 212.940 136.925 213.260 ;
        RECT 137.095 214.970 138.565 215.140 ;
        RECT 137.095 213.280 137.265 214.970 ;
        RECT 138.735 214.805 138.905 215.390 ;
        RECT 139.075 215.230 139.645 215.560 ;
        RECT 138.735 214.800 139.305 214.805 ;
        RECT 137.435 214.630 139.305 214.800 ;
        RECT 137.435 213.675 137.605 214.630 ;
        RECT 137.775 214.290 138.745 214.460 ;
        RECT 137.775 213.640 137.945 214.290 ;
        RECT 138.940 214.275 139.305 214.630 ;
        RECT 139.475 214.515 139.645 215.230 ;
        RECT 139.925 215.005 140.095 215.510 ;
        RECT 140.295 215.345 140.515 215.700 ;
        RECT 140.685 215.515 141.280 215.755 ;
        RECT 140.295 215.175 141.580 215.345 ;
        RECT 139.925 214.835 141.045 215.005 ;
        RECT 140.875 214.645 141.045 214.835 ;
        RECT 141.215 214.815 141.580 215.175 ;
        RECT 141.750 214.645 141.920 215.580 ;
        RECT 139.475 214.145 140.145 214.515 ;
        RECT 140.325 214.425 140.655 214.625 ;
        RECT 140.875 214.475 141.920 214.645 ;
        RECT 138.965 214.085 139.135 214.090 ;
        RECT 138.145 213.810 139.305 214.085 ;
        RECT 137.775 213.450 139.305 213.640 ;
        RECT 137.095 213.110 138.120 213.280 ;
        RECT 139.475 213.270 139.645 214.145 ;
        RECT 140.325 213.965 140.625 214.425 ;
        RECT 140.875 214.305 141.135 214.475 ;
        RECT 142.195 214.320 143.975 216.010 ;
        RECT 144.145 215.905 146.460 216.180 ;
        RECT 144.145 214.320 145.630 215.905 ;
        RECT 147.200 214.425 147.805 217.830 ;
        RECT 142.195 214.305 142.365 214.320 ;
        RECT 140.805 214.135 141.135 214.305 ;
        RECT 141.395 214.135 142.365 214.305 ;
        RECT 139.925 213.795 142.025 213.965 ;
        RECT 139.925 213.560 140.095 213.795 ;
        RECT 141.695 213.715 142.025 213.795 ;
        RECT 140.805 213.435 141.525 213.625 ;
        RECT 136.255 212.930 137.685 212.940 ;
        RECT 131.655 212.545 132.210 212.680 ;
        RECT 133.585 212.600 133.755 212.765 ;
        RECT 133.315 212.545 133.755 212.600 ;
        RECT 131.655 212.430 133.755 212.545 ;
        RECT 132.080 212.375 133.445 212.430 ;
        RECT 134.035 212.320 134.205 212.930 ;
        RECT 136.755 212.770 137.685 212.930 ;
        RECT 134.465 212.575 136.585 212.760 ;
        RECT 134.035 212.260 134.665 212.320 ;
        RECT 131.315 212.215 131.945 212.260 ;
        RECT 127.615 211.900 128.390 212.080 ;
        RECT 126.395 211.835 128.390 211.900 ;
        RECT 128.595 211.890 129.225 212.215 ;
        RECT 126.395 211.560 127.785 211.835 ;
        RECT 124.865 211.200 126.045 211.370 ;
        RECT 123.545 210.810 124.105 210.865 ;
        RECT 124.735 210.855 125.660 211.030 ;
        RECT 124.685 210.810 125.660 210.855 ;
        RECT 123.545 210.700 125.660 210.810 ;
        RECT 125.875 210.960 126.045 211.200 ;
        RECT 126.215 211.130 126.885 211.300 ;
        RECT 123.545 210.690 124.815 210.700 ;
        RECT 123.980 210.640 124.815 210.690 ;
        RECT 125.875 210.630 126.545 210.960 ;
        RECT 126.715 210.865 126.885 211.130 ;
        RECT 127.055 211.035 127.705 211.385 ;
        RECT 127.875 211.130 128.335 211.300 ;
        RECT 127.875 210.865 128.045 211.130 ;
        RECT 128.595 210.960 128.765 211.890 ;
        RECT 129.395 211.765 130.685 212.215 ;
        RECT 130.855 211.995 131.945 212.215 ;
        RECT 130.855 211.890 131.485 211.995 ;
        RECT 132.455 211.925 133.405 212.205 ;
        RECT 133.575 212.070 134.665 212.260 ;
        RECT 134.835 212.125 135.785 212.405 ;
        RECT 136.755 212.335 136.925 212.770 ;
        RECT 136.295 212.070 136.925 212.335 ;
        RECT 133.575 212.010 134.205 212.070 ;
        RECT 129.395 211.370 129.565 211.765 ;
        RECT 128.935 211.090 129.565 211.370 ;
        RECT 126.715 210.635 128.045 210.865 ;
        RECT 128.215 210.630 128.765 210.960 ;
        RECT 129.735 210.900 130.295 211.595 ;
        RECT 130.465 211.370 130.685 211.765 ;
        RECT 131.315 211.400 131.485 211.890 ;
        RECT 131.655 211.570 133.775 211.755 ;
        RECT 134.035 211.400 134.205 212.010 ;
        RECT 134.795 211.900 136.160 211.955 ;
        RECT 134.485 211.785 136.585 211.900 ;
        RECT 134.485 211.730 134.925 211.785 ;
        RECT 134.485 211.565 134.655 211.730 ;
        RECT 136.030 211.650 136.585 211.785 ;
        RECT 136.755 211.850 136.925 212.070 ;
        RECT 137.275 212.360 137.685 212.535 ;
        RECT 137.930 212.530 138.120 213.110 ;
        RECT 138.495 212.540 138.665 213.250 ;
        RECT 138.940 212.760 139.645 213.270 ;
        RECT 138.495 212.360 139.270 212.540 ;
        RECT 137.275 212.295 139.270 212.360 ;
        RECT 139.475 212.330 139.645 212.760 ;
        RECT 139.925 212.775 140.095 213.390 ;
        RECT 140.265 213.265 140.595 213.410 ;
        RECT 140.265 212.945 141.555 213.265 ;
        RECT 141.725 212.775 141.895 213.490 ;
        RECT 139.925 212.605 141.895 212.775 ;
        RECT 142.195 213.130 142.365 214.135 ;
        RECT 143.425 213.640 144.260 213.690 ;
        RECT 143.425 213.630 144.695 213.640 ;
        RECT 142.580 213.520 144.695 213.630 ;
        RECT 142.580 213.475 143.555 213.520 ;
        RECT 142.580 213.300 143.505 213.475 ;
        RECT 144.135 213.465 144.695 213.520 ;
        RECT 142.195 212.960 143.375 213.130 ;
        RECT 137.275 212.020 138.665 212.295 ;
        RECT 139.475 212.120 140.175 212.330 ;
        RECT 139.475 211.850 139.645 212.120 ;
        RECT 140.555 211.900 140.885 212.605 ;
        RECT 141.090 211.880 141.465 212.435 ;
        RECT 142.195 212.425 142.365 212.960 ;
        RECT 143.675 212.800 144.005 213.350 ;
        RECT 144.175 213.310 144.695 213.465 ;
        RECT 144.915 213.140 145.630 214.320 ;
        RECT 145.950 214.075 147.805 214.425 ;
        RECT 144.305 212.970 145.630 213.140 ;
        RECT 143.675 212.790 144.700 212.800 ;
        RECT 142.535 212.600 144.700 212.790 ;
        RECT 142.535 212.450 143.470 212.600 ;
        RECT 144.175 212.470 144.700 212.600 ;
        RECT 144.915 212.485 145.630 212.970 ;
        RECT 147.200 212.485 147.805 214.075 ;
        RECT 141.695 212.220 142.365 212.425 ;
        RECT 141.695 212.110 142.865 212.220 ;
        RECT 142.195 211.905 142.865 212.110 ;
        RECT 130.465 211.090 131.145 211.370 ;
        RECT 131.315 211.070 131.985 211.400 ;
        RECT 132.155 211.165 133.485 211.395 ;
        RECT 125.875 210.470 126.045 210.630 ;
        RECT 116.425 209.280 119.175 210.470 ;
        RECT 113.385 208.800 116.775 209.110 ;
        RECT 112.275 207.695 112.445 208.800 ;
        RECT 112.615 207.910 113.165 208.080 ;
        RECT 112.275 207.365 112.825 207.695 ;
        RECT 112.995 207.535 113.165 207.910 ;
        RECT 113.345 207.815 113.715 208.170 ;
        RECT 113.895 207.910 114.825 208.080 ;
        RECT 113.895 207.535 114.065 207.910 ;
        RECT 114.995 207.695 116.775 208.800 ;
        RECT 112.995 207.365 114.065 207.535 ;
        RECT 114.235 207.420 116.775 207.695 ;
        RECT 116.945 208.820 119.175 209.280 ;
        RECT 119.345 209.900 120.605 210.470 ;
        RECT 120.775 210.070 121.455 210.355 ;
        RECT 119.345 209.630 121.065 209.900 ;
        RECT 116.945 207.420 118.655 208.820 ;
        RECT 119.345 208.650 120.605 209.630 ;
        RECT 121.235 209.610 121.455 210.070 ;
        RECT 121.625 209.780 122.185 210.470 ;
        RECT 122.355 210.070 122.985 210.355 ;
        RECT 122.355 209.610 122.525 210.070 ;
        RECT 123.155 209.900 124.615 210.470 ;
        RECT 122.695 209.630 124.615 209.900 ;
        RECT 121.235 209.400 122.525 209.610 ;
        RECT 120.775 208.830 122.985 209.230 ;
        RECT 114.235 207.365 115.165 207.420 ;
        RECT 112.275 206.765 112.445 207.365 ;
        RECT 113.355 207.280 113.685 207.365 ;
        RECT 114.995 207.250 115.165 207.365 ;
        RECT 117.715 207.250 118.655 207.420 ;
        RECT 112.615 207.110 113.190 207.195 ;
        RECT 113.920 207.110 114.825 207.195 ;
        RECT 112.615 206.940 114.825 207.110 ;
        RECT 114.995 206.765 116.255 207.250 ;
        RECT 112.275 206.505 113.285 206.765 ;
        RECT 113.845 206.560 116.255 206.765 ;
        RECT 116.425 206.960 118.655 207.250 ;
        RECT 118.825 207.840 120.605 208.650 ;
        RECT 120.775 208.360 121.455 208.640 ;
        RECT 121.235 207.965 121.455 208.360 ;
        RECT 121.625 208.135 122.185 208.830 ;
        RECT 123.155 208.820 124.615 209.630 ;
        RECT 124.785 210.035 126.045 210.470 ;
        RECT 126.215 210.275 128.335 210.460 ;
        RECT 124.785 209.770 126.505 210.035 ;
        RECT 127.015 209.825 127.965 210.105 ;
        RECT 128.595 210.100 128.765 210.630 ;
        RECT 128.935 210.500 131.145 210.900 ;
        RECT 131.315 210.470 131.485 211.070 ;
        RECT 132.155 210.900 132.325 211.165 ;
        RECT 131.655 210.730 132.325 210.900 ;
        RECT 132.495 210.645 133.145 210.995 ;
        RECT 133.315 210.900 133.485 211.165 ;
        RECT 133.655 211.070 134.205 211.400 ;
        RECT 133.315 210.730 133.775 210.900 ;
        RECT 134.035 210.470 134.205 211.070 ;
        RECT 134.485 210.865 134.655 211.370 ;
        RECT 134.855 211.205 135.075 211.560 ;
        RECT 135.245 211.375 135.840 211.615 ;
        RECT 134.855 211.035 136.140 211.205 ;
        RECT 134.485 210.695 135.605 210.865 ;
        RECT 135.435 210.505 135.605 210.695 ;
        RECT 135.775 210.675 136.140 211.035 ;
        RECT 136.310 210.505 136.480 211.440 ;
        RECT 129.395 210.120 130.685 210.330 ;
        RECT 128.595 210.020 129.225 210.100 ;
        RECT 128.135 209.830 129.225 210.020 ;
        RECT 128.135 209.770 128.765 209.830 ;
        RECT 122.355 208.360 122.985 208.640 ;
        RECT 122.355 207.965 122.525 208.360 ;
        RECT 118.825 207.515 121.065 207.840 ;
        RECT 121.235 207.515 122.525 207.965 ;
        RECT 123.155 207.840 124.095 208.820 ;
        RECT 124.785 208.650 126.045 209.770 ;
        RECT 126.640 209.600 128.005 209.655 ;
        RECT 126.215 209.485 128.315 209.600 ;
        RECT 126.215 209.350 126.770 209.485 ;
        RECT 127.875 209.430 128.315 209.485 ;
        RECT 122.695 207.515 124.095 207.840 ;
        RECT 118.825 206.960 120.605 207.515 ;
        RECT 121.915 207.410 122.245 207.515 ;
        RECT 120.775 207.240 121.745 207.345 ;
        RECT 122.415 207.240 122.985 207.345 ;
        RECT 120.775 206.960 122.985 207.240 ;
        RECT 123.155 206.960 124.095 207.515 ;
        RECT 124.265 207.865 126.045 208.650 ;
        RECT 126.320 208.205 126.490 209.140 ;
        RECT 126.960 209.075 127.555 209.315 ;
        RECT 128.145 209.265 128.315 209.430 ;
        RECT 127.725 208.905 127.945 209.260 ;
        RECT 128.595 209.090 128.765 209.770 ;
        RECT 129.395 209.660 129.565 210.120 ;
        RECT 128.935 209.375 129.565 209.660 ;
        RECT 129.735 209.260 130.295 209.950 ;
        RECT 130.465 209.660 130.685 210.120 ;
        RECT 131.315 210.100 132.575 210.470 ;
        RECT 130.855 209.830 132.575 210.100 ;
        RECT 130.465 209.375 131.145 209.660 ;
        RECT 131.315 209.090 132.575 209.830 ;
        RECT 132.745 210.375 134.205 210.470 ;
        RECT 132.745 210.005 134.705 210.375 ;
        RECT 134.885 210.285 135.215 210.485 ;
        RECT 135.435 210.335 136.480 210.505 ;
        RECT 136.755 211.160 138.015 211.850 ;
        RECT 138.185 211.360 139.645 211.850 ;
        RECT 139.860 211.730 140.385 211.860 ;
        RECT 141.090 211.730 142.025 211.880 ;
        RECT 139.860 211.540 142.025 211.730 ;
        RECT 139.860 211.530 140.885 211.540 ;
        RECT 138.185 211.330 140.255 211.360 ;
        RECT 138.725 211.190 140.255 211.330 ;
        RECT 136.755 210.640 138.555 211.160 ;
        RECT 138.725 210.640 139.645 211.190 ;
        RECT 139.865 210.865 140.385 211.020 ;
        RECT 140.555 210.980 140.885 211.530 ;
        RECT 142.195 211.370 142.365 211.905 ;
        RECT 143.095 211.895 143.470 212.450 ;
        RECT 143.675 211.725 144.005 212.430 ;
        RECT 144.915 212.210 145.085 212.485 ;
        RECT 144.385 212.000 145.085 212.210 ;
        RECT 141.185 211.200 142.365 211.370 ;
        RECT 139.865 210.810 140.425 210.865 ;
        RECT 141.055 210.855 141.980 211.030 ;
        RECT 141.005 210.810 141.980 210.855 ;
        RECT 139.865 210.700 141.980 210.810 ;
        RECT 139.865 210.690 141.135 210.700 ;
        RECT 140.300 210.640 141.135 210.690 ;
        RECT 136.755 210.380 136.925 210.640 ;
        RECT 139.475 210.380 139.645 210.640 ;
        RECT 132.745 209.260 134.205 210.005 ;
        RECT 134.885 209.825 135.185 210.285 ;
        RECT 135.435 210.165 135.695 210.335 ;
        RECT 136.755 210.165 137.670 210.380 ;
        RECT 135.365 209.995 135.695 210.165 ;
        RECT 135.955 210.110 137.670 210.165 ;
        RECT 135.955 209.995 136.925 210.110 ;
        RECT 134.485 209.655 136.585 209.825 ;
        RECT 134.485 209.420 134.655 209.655 ;
        RECT 136.255 209.575 136.585 209.655 ;
        RECT 135.365 209.295 136.085 209.485 ;
        RECT 136.755 209.480 136.925 209.995 ;
        RECT 137.840 209.940 138.825 210.380 ;
        RECT 138.995 210.080 139.645 210.380 ;
        RECT 139.815 210.190 142.025 210.470 ;
        RECT 139.815 210.085 140.385 210.190 ;
        RECT 141.055 210.085 142.025 210.190 ;
        RECT 142.195 210.195 142.365 211.200 ;
        RECT 142.665 211.555 144.635 211.725 ;
        RECT 142.665 210.840 142.835 211.555 ;
        RECT 143.005 211.065 144.295 211.385 ;
        RECT 143.965 210.920 144.295 211.065 ;
        RECT 144.465 210.940 144.635 211.555 ;
        RECT 144.915 210.915 145.085 212.000 ;
        RECT 145.255 211.130 145.805 211.300 ;
        RECT 143.035 210.705 143.755 210.895 ;
        RECT 142.535 210.535 142.865 210.615 ;
        RECT 144.465 210.535 144.635 210.770 ;
        RECT 142.535 210.365 144.635 210.535 ;
        RECT 144.915 210.585 145.465 210.915 ;
        RECT 145.635 210.755 145.805 211.130 ;
        RECT 145.985 211.035 146.355 211.390 ;
        RECT 146.535 211.130 147.465 211.300 ;
        RECT 146.535 210.755 146.705 211.130 ;
        RECT 147.635 210.915 147.805 212.485 ;
        RECT 145.635 210.585 146.705 210.755 ;
        RECT 146.875 210.585 147.805 210.915 ;
        RECT 137.100 209.910 138.825 209.940 ;
        RECT 139.475 209.915 139.645 210.080 ;
        RECT 142.195 210.025 143.165 210.195 ;
        RECT 143.425 210.025 143.755 210.195 ;
        RECT 140.555 209.915 140.885 210.020 ;
        RECT 142.195 209.915 142.365 210.025 ;
        RECT 137.100 209.650 139.280 209.910 ;
        RECT 126.660 208.735 127.945 208.905 ;
        RECT 126.660 208.375 127.025 208.735 ;
        RECT 128.145 208.565 128.315 209.070 ;
        RECT 127.195 208.395 128.315 208.565 ;
        RECT 127.195 208.205 127.365 208.395 ;
        RECT 126.320 208.035 127.365 208.205 ;
        RECT 127.105 207.865 127.365 208.035 ;
        RECT 127.585 207.985 127.915 208.185 ;
        RECT 128.595 208.075 130.055 209.090 ;
        RECT 124.265 207.695 126.845 207.865 ;
        RECT 127.105 207.695 127.435 207.865 ;
        RECT 124.265 206.960 126.045 207.695 ;
        RECT 127.615 207.525 127.915 207.985 ;
        RECT 128.095 207.880 130.055 208.075 ;
        RECT 130.225 207.880 133.095 209.090 ;
        RECT 133.265 208.190 134.205 209.260 ;
        RECT 134.485 208.635 134.655 209.250 ;
        RECT 134.825 209.125 135.155 209.270 ;
        RECT 134.825 208.805 136.115 209.125 ;
        RECT 136.285 208.635 136.455 209.350 ;
        RECT 134.485 208.465 136.455 208.635 ;
        RECT 136.755 209.225 137.655 209.480 ;
        RECT 136.755 208.610 136.930 209.225 ;
        RECT 137.840 209.215 138.825 209.650 ;
        RECT 139.475 209.590 140.105 209.915 ;
        RECT 139.475 209.480 139.645 209.590 ;
        RECT 138.995 209.220 139.645 209.480 ;
        RECT 137.840 209.040 138.065 209.215 ;
        RECT 137.100 208.780 138.065 209.040 ;
        RECT 133.265 207.980 134.735 208.190 ;
        RECT 133.265 207.880 134.205 207.980 ;
        RECT 128.095 207.705 129.535 207.880 ;
        RECT 130.225 207.710 131.485 207.880 ;
        RECT 126.215 207.355 128.315 207.525 ;
        RECT 126.215 207.275 126.545 207.355 ;
        RECT 116.425 206.730 117.885 206.960 ;
        RECT 113.845 206.505 116.795 206.560 ;
        RECT 112.275 206.330 112.445 206.505 ;
        RECT 114.995 206.330 116.795 206.505 ;
        RECT 112.275 206.040 113.170 206.330 ;
        RECT 113.830 206.040 116.795 206.330 ;
        RECT 116.965 206.330 117.885 206.730 ;
        RECT 120.435 206.330 120.605 206.960 ;
        RECT 116.965 206.040 118.610 206.330 ;
        RECT 119.270 206.040 120.605 206.330 ;
        RECT 120.955 206.515 122.345 206.790 ;
        RECT 120.955 206.450 122.950 206.515 ;
        RECT 120.955 206.275 121.365 206.450 ;
        RECT 112.275 205.405 112.445 206.040 ;
        RECT 114.995 205.405 115.165 206.040 ;
        RECT 117.715 205.870 117.885 206.040 ;
        RECT 120.435 205.870 121.365 206.040 ;
        RECT 116.225 205.820 117.060 205.870 ;
        RECT 116.225 205.810 117.495 205.820 ;
        RECT 115.380 205.700 117.495 205.810 ;
        RECT 115.380 205.655 116.355 205.700 ;
        RECT 115.380 205.480 116.305 205.655 ;
        RECT 116.935 205.645 117.495 205.700 ;
        RECT 112.275 205.145 113.285 205.405 ;
        RECT 113.845 205.310 115.165 205.405 ;
        RECT 113.845 205.145 116.175 205.310 ;
        RECT 112.275 204.545 112.445 205.145 ;
        RECT 114.995 205.140 116.175 205.145 ;
        RECT 112.615 204.800 114.825 204.970 ;
        RECT 112.615 204.715 113.190 204.800 ;
        RECT 113.920 204.715 114.825 204.800 ;
        RECT 113.355 204.545 113.685 204.630 ;
        RECT 114.995 204.545 115.165 205.140 ;
        RECT 116.475 204.980 116.805 205.530 ;
        RECT 116.975 205.490 117.495 205.645 ;
        RECT 117.715 205.565 118.395 205.870 ;
        RECT 117.715 205.320 117.885 205.565 ;
        RECT 118.565 205.555 119.125 205.870 ;
        RECT 120.435 205.860 120.605 205.870 ;
        RECT 119.625 205.565 120.605 205.860 ;
        RECT 121.610 205.700 121.800 206.280 ;
        RECT 117.105 205.150 117.885 205.320 ;
        RECT 116.475 204.970 117.500 204.980 ;
        RECT 115.335 204.780 117.500 204.970 ;
        RECT 115.335 204.630 116.270 204.780 ;
        RECT 116.975 204.650 117.500 204.780 ;
        RECT 117.715 204.965 117.885 205.150 ;
        RECT 118.065 205.140 120.265 205.385 ;
        RECT 118.065 205.135 119.125 205.140 ;
        RECT 117.715 204.705 118.410 204.965 ;
        RECT 112.275 204.215 112.825 204.545 ;
        RECT 112.995 204.375 114.065 204.545 ;
        RECT 112.275 203.140 112.445 204.215 ;
        RECT 112.995 204.000 113.165 204.375 ;
        RECT 112.615 203.830 113.165 204.000 ;
        RECT 113.345 203.740 113.715 204.095 ;
        RECT 113.895 204.000 114.065 204.375 ;
        RECT 114.235 204.400 115.165 204.545 ;
        RECT 114.235 204.215 115.665 204.400 ;
        RECT 114.995 204.085 115.665 204.215 ;
        RECT 113.895 203.830 114.825 204.000 ;
        RECT 112.705 203.310 113.165 203.480 ;
        RECT 112.275 202.810 112.825 203.140 ;
        RECT 112.995 203.045 113.165 203.310 ;
        RECT 113.335 203.215 113.985 203.565 ;
        RECT 114.155 203.310 114.825 203.480 ;
        RECT 114.155 203.045 114.325 203.310 ;
        RECT 114.995 203.140 115.165 204.085 ;
        RECT 115.895 204.075 116.270 204.630 ;
        RECT 116.475 203.905 116.805 204.610 ;
        RECT 117.715 204.390 117.885 204.705 ;
        RECT 118.875 204.525 119.125 205.135 ;
        RECT 120.435 204.965 120.605 205.565 ;
        RECT 119.625 204.705 120.605 204.965 ;
        RECT 117.185 204.180 117.885 204.390 ;
        RECT 118.065 204.275 120.260 204.525 ;
        RECT 117.715 204.105 117.885 204.180 ;
        RECT 112.995 202.815 114.325 203.045 ;
        RECT 114.495 202.810 115.165 203.140 ;
        RECT 115.465 203.735 117.435 203.905 ;
        RECT 115.465 203.020 115.635 203.735 ;
        RECT 115.805 203.245 117.095 203.565 ;
        RECT 116.765 203.100 117.095 203.245 ;
        RECT 117.265 203.120 117.435 203.735 ;
        RECT 117.715 203.845 118.445 204.105 ;
        RECT 117.715 203.245 117.885 203.845 ;
        RECT 118.080 203.415 118.705 203.675 ;
        RECT 115.835 202.885 116.555 203.075 ;
        RECT 117.715 202.985 118.365 203.245 ;
        RECT 112.275 202.200 112.445 202.810 ;
        RECT 112.705 202.455 114.825 202.640 ;
        RECT 114.995 202.375 115.165 202.810 ;
        RECT 115.335 202.715 115.665 202.795 ;
        RECT 117.265 202.715 117.435 202.950 ;
        RECT 115.335 202.545 117.435 202.715 ;
        RECT 112.275 201.950 112.905 202.200 ;
        RECT 113.075 202.005 114.025 202.285 ;
        RECT 114.995 202.215 115.965 202.375 ;
        RECT 114.535 202.205 115.965 202.215 ;
        RECT 116.225 202.205 116.555 202.375 ;
        RECT 114.535 201.950 115.165 202.205 ;
        RECT 116.225 202.035 116.485 202.205 ;
        RECT 116.735 202.085 117.035 202.545 ;
        RECT 117.715 202.385 117.885 202.985 ;
        RECT 118.535 202.815 118.705 203.415 ;
        RECT 118.080 202.555 118.705 202.815 ;
        RECT 117.715 202.365 118.365 202.385 ;
        RECT 13.380 201.275 92.040 201.445 ;
        RECT 13.465 200.185 14.675 201.275 ;
        RECT 14.845 200.840 20.190 201.275 ;
        RECT 20.365 200.840 25.710 201.275 ;
        RECT 13.465 199.475 13.985 200.015 ;
        RECT 14.155 199.645 14.675 200.185 ;
        RECT 13.465 198.725 14.675 199.475 ;
        RECT 16.430 199.270 16.770 200.100 ;
        RECT 18.250 199.590 18.600 200.840 ;
        RECT 21.950 199.270 22.290 200.100 ;
        RECT 23.770 199.590 24.120 200.840 ;
        RECT 26.345 200.110 26.635 201.275 ;
        RECT 26.805 200.840 32.150 201.275 ;
        RECT 32.325 200.840 37.670 201.275 ;
        RECT 14.845 198.725 20.190 199.270 ;
        RECT 20.365 198.725 25.710 199.270 ;
        RECT 26.345 198.725 26.635 199.450 ;
        RECT 28.390 199.270 28.730 200.100 ;
        RECT 30.210 199.590 30.560 200.840 ;
        RECT 33.910 199.270 34.250 200.100 ;
        RECT 35.730 199.590 36.080 200.840 ;
        RECT 37.845 200.185 39.055 201.275 ;
        RECT 37.845 199.475 38.365 200.015 ;
        RECT 38.535 199.645 39.055 200.185 ;
        RECT 39.225 200.110 39.515 201.275 ;
        RECT 39.685 200.840 45.030 201.275 ;
        RECT 45.205 200.840 50.550 201.275 ;
        RECT 26.805 198.725 32.150 199.270 ;
        RECT 32.325 198.725 37.670 199.270 ;
        RECT 37.845 198.725 39.055 199.475 ;
        RECT 39.225 198.725 39.515 199.450 ;
        RECT 41.270 199.270 41.610 200.100 ;
        RECT 43.090 199.590 43.440 200.840 ;
        RECT 46.790 199.270 47.130 200.100 ;
        RECT 48.610 199.590 48.960 200.840 ;
        RECT 50.725 200.185 51.935 201.275 ;
        RECT 50.725 199.475 51.245 200.015 ;
        RECT 51.415 199.645 51.935 200.185 ;
        RECT 52.105 200.110 52.395 201.275 ;
        RECT 52.565 200.840 57.910 201.275 ;
        RECT 39.685 198.725 45.030 199.270 ;
        RECT 45.205 198.725 50.550 199.270 ;
        RECT 50.725 198.725 51.935 199.475 ;
        RECT 52.105 198.725 52.395 199.450 ;
        RECT 54.150 199.270 54.490 200.100 ;
        RECT 55.970 199.590 56.320 200.840 ;
        RECT 58.085 200.405 58.360 201.105 ;
        RECT 58.530 200.730 58.785 201.275 ;
        RECT 58.955 200.765 59.435 201.105 ;
        RECT 59.610 200.720 60.215 201.275 ;
        RECT 59.600 200.620 60.215 200.720 ;
        RECT 59.600 200.595 59.785 200.620 ;
        RECT 58.085 199.375 58.255 200.405 ;
        RECT 58.530 200.275 59.285 200.525 ;
        RECT 59.455 200.350 59.785 200.595 ;
        RECT 58.530 200.240 59.300 200.275 ;
        RECT 58.530 200.230 59.315 200.240 ;
        RECT 58.425 200.215 59.320 200.230 ;
        RECT 58.425 200.200 59.340 200.215 ;
        RECT 58.425 200.190 59.360 200.200 ;
        RECT 58.425 200.180 59.385 200.190 ;
        RECT 58.425 200.150 59.455 200.180 ;
        RECT 58.425 200.120 59.475 200.150 ;
        RECT 58.425 200.090 59.495 200.120 ;
        RECT 58.425 200.065 59.525 200.090 ;
        RECT 58.425 200.030 59.560 200.065 ;
        RECT 58.425 200.025 59.590 200.030 ;
        RECT 58.425 199.630 58.655 200.025 ;
        RECT 59.200 200.020 59.590 200.025 ;
        RECT 59.225 200.010 59.590 200.020 ;
        RECT 59.240 200.005 59.590 200.010 ;
        RECT 59.255 200.000 59.590 200.005 ;
        RECT 59.955 200.000 60.215 200.450 ;
        RECT 60.385 200.185 62.975 201.275 ;
        RECT 59.255 199.995 60.215 200.000 ;
        RECT 59.265 199.985 60.215 199.995 ;
        RECT 59.275 199.980 60.215 199.985 ;
        RECT 59.285 199.970 60.215 199.980 ;
        RECT 59.290 199.960 60.215 199.970 ;
        RECT 59.295 199.955 60.215 199.960 ;
        RECT 59.305 199.940 60.215 199.955 ;
        RECT 59.310 199.925 60.215 199.940 ;
        RECT 59.320 199.900 60.215 199.925 ;
        RECT 58.825 199.430 59.155 199.855 ;
        RECT 52.565 198.725 57.910 199.270 ;
        RECT 58.085 198.895 58.345 199.375 ;
        RECT 58.515 198.725 58.765 199.265 ;
        RECT 58.935 198.945 59.155 199.430 ;
        RECT 59.325 199.830 60.215 199.900 ;
        RECT 59.325 199.105 59.495 199.830 ;
        RECT 59.665 199.275 60.215 199.660 ;
        RECT 60.385 199.495 61.595 200.015 ;
        RECT 61.765 199.665 62.975 200.185 ;
        RECT 63.235 200.345 63.405 201.105 ;
        RECT 63.585 200.515 63.915 201.275 ;
        RECT 63.235 200.175 63.900 200.345 ;
        RECT 64.085 200.200 64.355 201.105 ;
        RECT 63.730 200.030 63.900 200.175 ;
        RECT 63.165 199.625 63.495 199.995 ;
        RECT 63.730 199.700 64.015 200.030 ;
        RECT 59.325 198.935 60.215 199.105 ;
        RECT 60.385 198.725 62.975 199.495 ;
        RECT 63.730 199.445 63.900 199.700 ;
        RECT 63.235 199.275 63.900 199.445 ;
        RECT 64.185 199.400 64.355 200.200 ;
        RECT 64.985 200.110 65.275 201.275 ;
        RECT 65.445 200.840 70.790 201.275 ;
        RECT 63.235 198.895 63.405 199.275 ;
        RECT 63.585 198.725 63.915 199.105 ;
        RECT 64.095 198.895 64.355 199.400 ;
        RECT 64.985 198.725 65.275 199.450 ;
        RECT 67.030 199.270 67.370 200.100 ;
        RECT 68.850 199.590 69.200 200.840 ;
        RECT 70.965 200.185 72.635 201.275 ;
        RECT 70.965 199.495 71.715 200.015 ;
        RECT 71.885 199.665 72.635 200.185 ;
        RECT 72.805 200.200 73.075 201.105 ;
        RECT 73.245 200.515 73.575 201.275 ;
        RECT 73.755 200.345 73.925 201.105 ;
        RECT 65.445 198.725 70.790 199.270 ;
        RECT 70.965 198.725 72.635 199.495 ;
        RECT 72.805 199.400 72.975 200.200 ;
        RECT 73.260 200.175 73.925 200.345 ;
        RECT 74.185 200.185 77.695 201.275 ;
        RECT 73.260 200.030 73.430 200.175 ;
        RECT 73.145 199.700 73.430 200.030 ;
        RECT 73.260 199.445 73.430 199.700 ;
        RECT 73.665 199.625 73.995 199.995 ;
        RECT 74.185 199.495 75.835 200.015 ;
        RECT 76.005 199.665 77.695 200.185 ;
        RECT 77.865 200.110 78.155 201.275 ;
        RECT 78.325 200.840 83.670 201.275 ;
        RECT 83.845 200.840 89.190 201.275 ;
        RECT 72.805 198.895 73.065 199.400 ;
        RECT 73.260 199.275 73.925 199.445 ;
        RECT 73.245 198.725 73.575 199.105 ;
        RECT 73.755 198.895 73.925 199.275 ;
        RECT 74.185 198.725 77.695 199.495 ;
        RECT 77.865 198.725 78.155 199.450 ;
        RECT 79.910 199.270 80.250 200.100 ;
        RECT 81.730 199.590 82.080 200.840 ;
        RECT 85.430 199.270 85.770 200.100 ;
        RECT 87.250 199.590 87.600 200.840 ;
        RECT 89.365 200.185 90.575 201.275 ;
        RECT 89.365 199.475 89.885 200.015 ;
        RECT 90.055 199.645 90.575 200.185 ;
        RECT 90.745 200.185 91.955 201.275 ;
        RECT 112.275 200.255 112.445 201.950 ;
        RECT 113.035 201.780 114.400 201.835 ;
        RECT 112.725 201.665 114.825 201.780 ;
        RECT 112.725 201.610 113.165 201.665 ;
        RECT 112.725 201.445 112.895 201.610 ;
        RECT 114.270 201.530 114.825 201.665 ;
        RECT 112.725 200.745 112.895 201.250 ;
        RECT 113.095 201.085 113.315 201.440 ;
        RECT 113.485 201.255 114.080 201.495 ;
        RECT 113.095 200.915 114.380 201.085 ;
        RECT 112.725 200.575 113.845 200.745 ;
        RECT 113.675 200.385 113.845 200.575 ;
        RECT 114.015 200.555 114.380 200.915 ;
        RECT 114.550 200.385 114.720 201.320 ;
        RECT 90.745 199.645 91.265 200.185 ;
        RECT 91.435 199.475 91.955 200.015 ;
        RECT 78.325 198.725 83.670 199.270 ;
        RECT 83.845 198.725 89.190 199.270 ;
        RECT 89.365 198.725 90.575 199.475 ;
        RECT 90.745 198.725 91.955 199.475 ;
        RECT 112.275 199.885 112.945 200.255 ;
        RECT 113.125 200.165 113.455 200.365 ;
        RECT 113.675 200.215 114.720 200.385 ;
        RECT 114.995 200.300 115.165 201.950 ;
        RECT 115.440 201.865 116.485 202.035 ;
        RECT 116.705 201.885 117.035 202.085 ;
        RECT 117.215 202.125 118.365 202.365 ;
        RECT 117.215 201.995 117.885 202.125 ;
        RECT 115.440 200.930 115.610 201.865 ;
        RECT 115.780 201.335 116.145 201.695 ;
        RECT 116.315 201.675 116.485 201.865 ;
        RECT 116.315 201.505 117.435 201.675 ;
        RECT 115.780 201.165 117.065 201.335 ;
        RECT 116.080 200.755 116.675 200.995 ;
        RECT 116.845 200.810 117.065 201.165 ;
        RECT 117.265 201.000 117.435 201.505 ;
        RECT 117.715 201.525 117.885 201.995 ;
        RECT 118.535 201.955 118.705 202.555 ;
        RECT 118.080 201.695 118.705 201.955 ;
        RECT 117.715 201.280 118.365 201.525 ;
        RECT 115.335 200.585 115.890 200.720 ;
        RECT 117.265 200.640 117.435 200.805 ;
        RECT 116.995 200.585 117.435 200.640 ;
        RECT 115.335 200.470 117.435 200.585 ;
        RECT 117.715 200.665 117.885 201.280 ;
        RECT 118.535 201.110 118.705 201.695 ;
        RECT 118.080 200.835 118.705 201.110 ;
        RECT 115.760 200.415 117.125 200.470 ;
        RECT 117.715 200.420 118.365 200.665 ;
        RECT 117.715 200.300 117.885 200.420 ;
        RECT 13.380 198.555 92.040 198.725 ;
        RECT 13.465 197.805 14.675 198.555 ;
        RECT 14.845 198.010 20.190 198.555 ;
        RECT 20.365 198.010 25.710 198.555 ;
        RECT 25.885 198.010 31.230 198.555 ;
        RECT 31.405 198.010 36.750 198.555 ;
        RECT 13.465 197.265 13.985 197.805 ;
        RECT 14.155 197.095 14.675 197.635 ;
        RECT 16.430 197.180 16.770 198.010 ;
        RECT 13.465 196.005 14.675 197.095 ;
        RECT 18.250 196.440 18.600 197.690 ;
        RECT 21.950 197.180 22.290 198.010 ;
        RECT 23.770 196.440 24.120 197.690 ;
        RECT 27.470 197.180 27.810 198.010 ;
        RECT 29.290 196.440 29.640 197.690 ;
        RECT 32.990 197.180 33.330 198.010 ;
        RECT 36.925 197.785 38.595 198.555 ;
        RECT 39.225 197.830 39.515 198.555 ;
        RECT 39.685 197.785 42.275 198.555 ;
        RECT 34.810 196.440 35.160 197.690 ;
        RECT 36.925 197.265 37.675 197.785 ;
        RECT 37.845 197.095 38.595 197.615 ;
        RECT 39.685 197.265 40.895 197.785 ;
        RECT 42.455 197.745 42.725 198.555 ;
        RECT 42.895 197.745 43.225 198.385 ;
        RECT 43.395 197.745 43.635 198.555 ;
        RECT 43.825 198.175 44.715 198.345 ;
        RECT 14.845 196.005 20.190 196.440 ;
        RECT 20.365 196.005 25.710 196.440 ;
        RECT 25.885 196.005 31.230 196.440 ;
        RECT 31.405 196.005 36.750 196.440 ;
        RECT 36.925 196.005 38.595 197.095 ;
        RECT 39.225 196.005 39.515 197.170 ;
        RECT 41.065 197.095 42.275 197.615 ;
        RECT 42.445 197.315 42.795 197.565 ;
        RECT 42.965 197.145 43.135 197.745 ;
        RECT 43.825 197.620 44.375 198.005 ;
        RECT 43.305 197.315 43.655 197.565 ;
        RECT 44.545 197.450 44.715 198.175 ;
        RECT 43.825 197.380 44.715 197.450 ;
        RECT 44.885 197.850 45.105 198.335 ;
        RECT 45.275 198.015 45.525 198.555 ;
        RECT 45.695 197.905 45.955 198.385 ;
        RECT 44.885 197.425 45.215 197.850 ;
        RECT 43.825 197.355 44.720 197.380 ;
        RECT 43.825 197.340 44.730 197.355 ;
        RECT 43.825 197.325 44.735 197.340 ;
        RECT 43.825 197.320 44.745 197.325 ;
        RECT 43.825 197.310 44.750 197.320 ;
        RECT 43.825 197.300 44.755 197.310 ;
        RECT 43.825 197.295 44.765 197.300 ;
        RECT 43.825 197.285 44.775 197.295 ;
        RECT 43.825 197.280 44.785 197.285 ;
        RECT 39.685 196.005 42.275 197.095 ;
        RECT 42.455 196.005 42.785 197.145 ;
        RECT 42.965 196.975 43.645 197.145 ;
        RECT 43.315 196.190 43.645 196.975 ;
        RECT 43.825 196.830 44.085 197.280 ;
        RECT 44.450 197.275 44.785 197.280 ;
        RECT 44.450 197.270 44.800 197.275 ;
        RECT 44.450 197.260 44.815 197.270 ;
        RECT 44.450 197.255 44.840 197.260 ;
        RECT 45.385 197.255 45.615 197.650 ;
        RECT 44.450 197.250 45.615 197.255 ;
        RECT 44.480 197.215 45.615 197.250 ;
        RECT 44.515 197.190 45.615 197.215 ;
        RECT 44.545 197.160 45.615 197.190 ;
        RECT 44.565 197.130 45.615 197.160 ;
        RECT 44.585 197.100 45.615 197.130 ;
        RECT 44.655 197.090 45.615 197.100 ;
        RECT 44.680 197.080 45.615 197.090 ;
        RECT 44.700 197.065 45.615 197.080 ;
        RECT 44.720 197.050 45.615 197.065 ;
        RECT 44.725 197.040 45.510 197.050 ;
        RECT 44.740 197.005 45.510 197.040 ;
        RECT 44.255 196.685 44.585 196.930 ;
        RECT 44.755 196.755 45.510 197.005 ;
        RECT 45.785 196.875 45.955 197.905 ;
        RECT 46.215 198.005 46.385 198.295 ;
        RECT 46.555 198.175 46.885 198.555 ;
        RECT 46.215 197.835 46.880 198.005 ;
        RECT 46.130 197.015 46.480 197.665 ;
        RECT 44.255 196.660 44.440 196.685 ;
        RECT 43.825 196.560 44.440 196.660 ;
        RECT 43.825 196.005 44.430 196.560 ;
        RECT 44.605 196.175 45.085 196.515 ;
        RECT 45.255 196.005 45.510 196.550 ;
        RECT 45.680 196.175 45.955 196.875 ;
        RECT 46.650 196.845 46.880 197.835 ;
        RECT 46.215 196.675 46.880 196.845 ;
        RECT 46.215 196.175 46.385 196.675 ;
        RECT 46.555 196.005 46.885 196.505 ;
        RECT 47.055 196.175 47.240 198.295 ;
        RECT 47.495 198.095 47.745 198.555 ;
        RECT 47.915 198.105 48.250 198.275 ;
        RECT 48.445 198.105 49.120 198.275 ;
        RECT 47.915 197.965 48.085 198.105 ;
        RECT 47.410 196.975 47.690 197.925 ;
        RECT 47.860 197.835 48.085 197.965 ;
        RECT 47.860 196.730 48.030 197.835 ;
        RECT 48.255 197.685 48.780 197.905 ;
        RECT 48.200 196.920 48.440 197.515 ;
        RECT 48.610 196.985 48.780 197.685 ;
        RECT 48.950 197.325 49.120 198.105 ;
        RECT 49.440 198.055 49.810 198.555 ;
        RECT 49.990 198.105 50.395 198.275 ;
        RECT 50.565 198.105 51.350 198.275 ;
        RECT 49.990 197.875 50.160 198.105 ;
        RECT 49.330 197.575 50.160 197.875 ;
        RECT 50.545 197.605 51.010 197.935 ;
        RECT 49.330 197.545 49.530 197.575 ;
        RECT 49.650 197.325 49.820 197.395 ;
        RECT 48.950 197.155 49.820 197.325 ;
        RECT 49.310 197.065 49.820 197.155 ;
        RECT 47.860 196.600 48.165 196.730 ;
        RECT 48.610 196.620 49.140 196.985 ;
        RECT 47.480 196.005 47.745 196.465 ;
        RECT 47.915 196.175 48.165 196.600 ;
        RECT 49.310 196.450 49.480 197.065 ;
        RECT 48.375 196.280 49.480 196.450 ;
        RECT 49.650 196.005 49.820 196.805 ;
        RECT 49.990 196.505 50.160 197.575 ;
        RECT 50.330 196.675 50.520 197.395 ;
        RECT 50.690 196.645 51.010 197.605 ;
        RECT 51.180 197.645 51.350 198.105 ;
        RECT 51.625 198.025 51.835 198.555 ;
        RECT 52.095 197.815 52.425 198.340 ;
        RECT 52.595 197.945 52.765 198.555 ;
        RECT 52.935 197.900 53.265 198.335 ;
        RECT 52.935 197.815 53.315 197.900 ;
        RECT 52.225 197.645 52.425 197.815 ;
        RECT 53.090 197.775 53.315 197.815 ;
        RECT 51.180 197.315 52.055 197.645 ;
        RECT 52.225 197.315 52.975 197.645 ;
        RECT 49.990 196.175 50.240 196.505 ;
        RECT 51.180 196.475 51.350 197.315 ;
        RECT 52.225 197.110 52.415 197.315 ;
        RECT 53.145 197.195 53.315 197.775 ;
        RECT 53.485 197.785 56.995 198.555 ;
        RECT 57.255 198.005 57.425 198.295 ;
        RECT 57.595 198.175 57.925 198.555 ;
        RECT 57.255 197.835 57.920 198.005 ;
        RECT 53.485 197.265 55.135 197.785 ;
        RECT 53.100 197.145 53.315 197.195 ;
        RECT 51.520 196.735 52.415 197.110 ;
        RECT 52.925 197.065 53.315 197.145 ;
        RECT 55.305 197.095 56.995 197.615 ;
        RECT 50.465 196.305 51.350 196.475 ;
        RECT 51.530 196.005 51.845 196.505 ;
        RECT 52.075 196.175 52.415 196.735 ;
        RECT 52.585 196.005 52.755 197.015 ;
        RECT 52.925 196.220 53.255 197.065 ;
        RECT 53.485 196.005 56.995 197.095 ;
        RECT 57.170 197.015 57.520 197.665 ;
        RECT 57.690 196.845 57.920 197.835 ;
        RECT 57.255 196.675 57.920 196.845 ;
        RECT 57.255 196.175 57.425 196.675 ;
        RECT 57.595 196.005 57.925 196.505 ;
        RECT 58.095 196.175 58.280 198.295 ;
        RECT 58.535 198.095 58.785 198.555 ;
        RECT 58.955 198.105 59.290 198.275 ;
        RECT 59.485 198.105 60.160 198.275 ;
        RECT 58.955 197.965 59.125 198.105 ;
        RECT 58.450 196.975 58.730 197.925 ;
        RECT 58.900 197.835 59.125 197.965 ;
        RECT 58.900 196.730 59.070 197.835 ;
        RECT 59.295 197.685 59.820 197.905 ;
        RECT 59.240 196.920 59.480 197.515 ;
        RECT 59.650 196.985 59.820 197.685 ;
        RECT 59.990 197.325 60.160 198.105 ;
        RECT 60.480 198.055 60.850 198.555 ;
        RECT 61.030 198.105 61.435 198.275 ;
        RECT 61.605 198.105 62.390 198.275 ;
        RECT 61.030 197.875 61.200 198.105 ;
        RECT 60.370 197.575 61.200 197.875 ;
        RECT 61.585 197.605 62.050 197.935 ;
        RECT 60.370 197.545 60.570 197.575 ;
        RECT 60.690 197.325 60.860 197.395 ;
        RECT 59.990 197.155 60.860 197.325 ;
        RECT 60.350 197.065 60.860 197.155 ;
        RECT 58.900 196.600 59.205 196.730 ;
        RECT 59.650 196.620 60.180 196.985 ;
        RECT 58.520 196.005 58.785 196.465 ;
        RECT 58.955 196.175 59.205 196.600 ;
        RECT 60.350 196.450 60.520 197.065 ;
        RECT 59.415 196.280 60.520 196.450 ;
        RECT 60.690 196.005 60.860 196.805 ;
        RECT 61.030 196.505 61.200 197.575 ;
        RECT 61.370 196.675 61.560 197.395 ;
        RECT 61.730 196.645 62.050 197.605 ;
        RECT 62.220 197.645 62.390 198.105 ;
        RECT 62.665 198.025 62.875 198.555 ;
        RECT 63.135 197.815 63.465 198.340 ;
        RECT 63.635 197.945 63.805 198.555 ;
        RECT 63.975 197.900 64.305 198.335 ;
        RECT 63.975 197.815 64.355 197.900 ;
        RECT 64.985 197.830 65.275 198.555 ;
        RECT 63.265 197.645 63.465 197.815 ;
        RECT 64.130 197.775 64.355 197.815 ;
        RECT 62.220 197.315 63.095 197.645 ;
        RECT 63.265 197.315 64.015 197.645 ;
        RECT 61.030 196.175 61.280 196.505 ;
        RECT 62.220 196.475 62.390 197.315 ;
        RECT 63.265 197.110 63.455 197.315 ;
        RECT 64.185 197.195 64.355 197.775 ;
        RECT 65.445 197.785 67.115 198.555 ;
        RECT 67.795 197.900 68.125 198.335 ;
        RECT 68.295 197.945 68.465 198.555 ;
        RECT 67.745 197.815 68.125 197.900 ;
        RECT 68.635 197.815 68.965 198.340 ;
        RECT 69.225 198.025 69.435 198.555 ;
        RECT 69.710 198.105 70.495 198.275 ;
        RECT 70.665 198.105 71.070 198.275 ;
        RECT 65.445 197.265 66.195 197.785 ;
        RECT 67.745 197.775 67.970 197.815 ;
        RECT 64.140 197.145 64.355 197.195 ;
        RECT 62.560 196.735 63.455 197.110 ;
        RECT 63.965 197.065 64.355 197.145 ;
        RECT 61.505 196.305 62.390 196.475 ;
        RECT 62.570 196.005 62.885 196.505 ;
        RECT 63.115 196.175 63.455 196.735 ;
        RECT 63.625 196.005 63.795 197.015 ;
        RECT 63.965 196.220 64.295 197.065 ;
        RECT 64.985 196.005 65.275 197.170 ;
        RECT 66.365 197.095 67.115 197.615 ;
        RECT 65.445 196.005 67.115 197.095 ;
        RECT 67.745 197.195 67.915 197.775 ;
        RECT 68.635 197.645 68.835 197.815 ;
        RECT 69.710 197.645 69.880 198.105 ;
        RECT 68.085 197.315 68.835 197.645 ;
        RECT 69.005 197.315 69.880 197.645 ;
        RECT 67.745 197.145 67.960 197.195 ;
        RECT 67.745 197.065 68.135 197.145 ;
        RECT 67.805 196.220 68.135 197.065 ;
        RECT 68.645 197.110 68.835 197.315 ;
        RECT 68.305 196.005 68.475 197.015 ;
        RECT 68.645 196.735 69.540 197.110 ;
        RECT 68.645 196.175 68.985 196.735 ;
        RECT 69.215 196.005 69.530 196.505 ;
        RECT 69.710 196.475 69.880 197.315 ;
        RECT 70.050 197.605 70.515 197.935 ;
        RECT 70.900 197.875 71.070 198.105 ;
        RECT 71.250 198.055 71.620 198.555 ;
        RECT 71.940 198.105 72.615 198.275 ;
        RECT 72.810 198.105 73.145 198.275 ;
        RECT 70.050 196.645 70.370 197.605 ;
        RECT 70.900 197.575 71.730 197.875 ;
        RECT 70.540 196.675 70.730 197.395 ;
        RECT 70.900 196.505 71.070 197.575 ;
        RECT 71.530 197.545 71.730 197.575 ;
        RECT 71.240 197.325 71.410 197.395 ;
        RECT 71.940 197.325 72.110 198.105 ;
        RECT 72.975 197.965 73.145 198.105 ;
        RECT 73.315 198.095 73.565 198.555 ;
        RECT 71.240 197.155 72.110 197.325 ;
        RECT 72.280 197.685 72.805 197.905 ;
        RECT 72.975 197.835 73.200 197.965 ;
        RECT 71.240 197.065 71.750 197.155 ;
        RECT 69.710 196.305 70.595 196.475 ;
        RECT 70.820 196.175 71.070 196.505 ;
        RECT 71.240 196.005 71.410 196.805 ;
        RECT 71.580 196.450 71.750 197.065 ;
        RECT 72.280 196.985 72.450 197.685 ;
        RECT 71.920 196.620 72.450 196.985 ;
        RECT 72.620 196.920 72.860 197.515 ;
        RECT 73.030 196.730 73.200 197.835 ;
        RECT 73.370 196.975 73.650 197.925 ;
        RECT 72.895 196.600 73.200 196.730 ;
        RECT 71.580 196.280 72.685 196.450 ;
        RECT 72.895 196.175 73.145 196.600 ;
        RECT 73.315 196.005 73.580 196.465 ;
        RECT 73.820 196.175 74.005 198.295 ;
        RECT 74.175 198.175 74.505 198.555 ;
        RECT 74.675 198.005 74.845 198.295 ;
        RECT 75.105 198.010 80.450 198.555 ;
        RECT 80.625 198.010 85.970 198.555 ;
        RECT 74.180 197.835 74.845 198.005 ;
        RECT 74.180 196.845 74.410 197.835 ;
        RECT 74.580 197.015 74.930 197.665 ;
        RECT 76.690 197.180 77.030 198.010 ;
        RECT 74.180 196.675 74.845 196.845 ;
        RECT 74.175 196.005 74.505 196.505 ;
        RECT 74.675 196.175 74.845 196.675 ;
        RECT 78.510 196.440 78.860 197.690 ;
        RECT 82.210 197.180 82.550 198.010 ;
        RECT 86.145 197.785 89.655 198.555 ;
        RECT 90.745 197.805 91.955 198.555 ;
        RECT 84.030 196.440 84.380 197.690 ;
        RECT 86.145 197.265 87.795 197.785 ;
        RECT 87.965 197.095 89.655 197.615 ;
        RECT 75.105 196.005 80.450 196.440 ;
        RECT 80.625 196.005 85.970 196.440 ;
        RECT 86.145 196.005 89.655 197.095 ;
        RECT 90.745 197.095 91.265 197.635 ;
        RECT 91.435 197.265 91.955 197.805 ;
        RECT 112.275 198.070 112.445 199.885 ;
        RECT 113.125 199.705 113.425 200.165 ;
        RECT 113.675 200.045 113.935 200.215 ;
        RECT 114.995 200.045 115.625 200.300 ;
        RECT 113.605 199.875 113.935 200.045 ;
        RECT 114.195 200.035 115.625 200.045 ;
        RECT 114.195 199.875 115.165 200.035 ;
        RECT 116.135 199.965 117.085 200.245 ;
        RECT 117.255 200.050 117.885 200.300 ;
        RECT 118.535 200.250 118.705 200.835 ;
        RECT 112.725 199.535 114.825 199.705 ;
        RECT 112.725 199.300 112.895 199.535 ;
        RECT 114.495 199.455 114.825 199.535 ;
        RECT 114.995 199.440 115.165 199.875 ;
        RECT 117.715 199.810 117.885 200.050 ;
        RECT 118.080 199.990 118.705 200.250 ;
        RECT 115.335 199.610 117.455 199.795 ;
        RECT 117.715 199.560 118.365 199.810 ;
        RECT 117.715 199.440 117.885 199.560 ;
        RECT 113.605 199.175 114.325 199.365 ;
        RECT 112.725 198.515 112.895 199.130 ;
        RECT 113.065 199.005 113.395 199.150 ;
        RECT 113.065 198.685 114.355 199.005 ;
        RECT 114.525 198.515 114.695 199.230 ;
        RECT 112.725 198.345 114.695 198.515 ;
        RECT 114.995 199.110 115.665 199.440 ;
        RECT 115.835 199.205 117.165 199.435 ;
        RECT 112.275 197.860 112.975 198.070 ;
        RECT 112.275 197.100 112.445 197.860 ;
        RECT 113.355 197.640 113.685 198.345 ;
        RECT 113.890 197.620 114.265 198.175 ;
        RECT 114.995 198.165 115.165 199.110 ;
        RECT 115.835 198.940 116.005 199.205 ;
        RECT 115.335 198.770 116.005 198.940 ;
        RECT 116.175 198.685 116.825 199.035 ;
        RECT 116.995 198.940 117.165 199.205 ;
        RECT 117.335 199.110 117.885 199.440 ;
        RECT 118.535 199.390 118.705 199.990 ;
        RECT 118.080 199.130 118.705 199.390 ;
        RECT 117.715 198.950 117.885 199.110 ;
        RECT 116.995 198.770 117.455 198.940 ;
        RECT 117.715 198.700 118.365 198.950 ;
        RECT 115.335 198.335 117.545 198.505 ;
        RECT 115.335 198.170 116.305 198.335 ;
        RECT 116.975 198.250 117.545 198.335 ;
        RECT 114.495 198.000 115.165 198.165 ;
        RECT 116.475 198.080 116.805 198.165 ;
        RECT 117.715 198.090 117.885 198.700 ;
        RECT 118.535 198.530 118.705 199.130 ;
        RECT 118.080 198.270 118.705 198.530 ;
        RECT 118.535 198.095 118.705 198.270 ;
        RECT 118.875 198.265 119.125 204.275 ;
        RECT 120.435 204.105 120.605 204.705 ;
        RECT 119.635 203.845 120.605 204.105 ;
        RECT 119.295 203.415 120.260 203.675 ;
        RECT 120.430 203.500 120.605 203.845 ;
        RECT 120.775 205.530 121.800 205.700 ;
        RECT 122.175 206.270 122.950 206.450 ;
        RECT 123.155 206.330 123.325 206.960 ;
        RECT 125.875 206.330 126.045 206.960 ;
        RECT 122.175 205.560 122.345 206.270 ;
        RECT 123.155 206.050 124.050 206.330 ;
        RECT 122.620 206.040 124.050 206.050 ;
        RECT 124.710 206.040 126.045 206.330 ;
        RECT 126.345 206.335 126.515 207.050 ;
        RECT 126.715 206.995 127.435 207.185 ;
        RECT 128.145 207.120 128.315 207.355 ;
        RECT 127.645 206.825 127.975 206.970 ;
        RECT 126.685 206.505 127.975 206.825 ;
        RECT 128.145 206.335 128.315 206.950 ;
        RECT 126.345 206.165 128.315 206.335 ;
        RECT 128.595 206.500 129.535 207.705 ;
        RECT 129.705 207.240 131.485 207.710 ;
        RECT 134.035 207.250 134.205 207.880 ;
        RECT 135.115 207.760 135.445 208.465 ;
        RECT 136.755 208.365 137.655 208.610 ;
        RECT 135.650 207.740 136.025 208.295 ;
        RECT 136.755 208.285 136.930 208.365 ;
        RECT 136.255 207.970 136.930 208.285 ;
        RECT 137.825 208.180 138.065 208.780 ;
        RECT 136.755 207.750 136.930 207.970 ;
        RECT 137.100 207.920 138.065 208.180 ;
        RECT 134.420 207.590 134.945 207.720 ;
        RECT 135.650 207.590 136.585 207.740 ;
        RECT 134.420 207.400 136.585 207.590 ;
        RECT 136.755 207.505 137.655 207.750 ;
        RECT 134.420 207.390 135.445 207.400 ;
        RECT 129.705 206.945 132.295 207.240 ;
        RECT 129.705 206.500 131.485 206.945 ;
        RECT 132.795 206.935 133.355 207.250 ;
        RECT 133.525 207.220 134.205 207.250 ;
        RECT 133.525 207.050 134.815 207.220 ;
        RECT 133.525 206.945 134.205 207.050 ;
        RECT 131.655 206.520 133.855 206.765 ;
        RECT 128.595 206.330 128.765 206.500 ;
        RECT 131.315 206.345 131.485 206.500 ;
        RECT 132.795 206.515 133.855 206.520 ;
        RECT 131.315 206.330 132.295 206.345 ;
        RECT 122.620 205.540 123.325 206.040 ;
        RECT 125.875 205.985 126.045 206.040 ;
        RECT 123.585 205.610 124.045 205.780 ;
        RECT 120.775 203.840 120.945 205.530 ;
        RECT 123.155 205.440 123.325 205.540 ;
        RECT 121.455 205.170 122.985 205.360 ;
        RECT 121.115 204.180 121.285 205.135 ;
        RECT 121.455 204.520 121.625 205.170 ;
        RECT 123.155 205.110 123.705 205.440 ;
        RECT 123.875 205.345 124.045 205.610 ;
        RECT 124.215 205.515 124.865 205.865 ;
        RECT 125.035 205.610 125.705 205.780 ;
        RECT 125.875 205.670 126.545 205.985 ;
        RECT 125.035 205.345 125.205 205.610 ;
        RECT 125.875 205.440 126.045 205.670 ;
        RECT 126.775 205.440 127.150 205.995 ;
        RECT 127.355 205.460 127.685 206.165 ;
        RECT 128.595 206.040 129.490 206.330 ;
        RECT 130.150 206.085 132.295 206.330 ;
        RECT 130.150 206.040 131.485 206.085 ;
        RECT 128.595 205.890 128.765 206.040 ;
        RECT 128.065 205.860 128.765 205.890 ;
        RECT 128.065 205.680 129.575 205.860 ;
        RECT 128.595 205.590 129.575 205.680 ;
        RECT 123.875 205.115 125.205 205.345 ;
        RECT 125.375 205.110 126.045 205.440 ;
        RECT 121.825 204.725 122.985 205.000 ;
        RECT 121.965 204.720 122.135 204.725 ;
        RECT 121.455 204.350 122.425 204.520 ;
        RECT 122.620 204.180 122.985 204.535 ;
        RECT 121.115 204.010 122.985 204.180 ;
        RECT 122.415 204.005 122.985 204.010 ;
        RECT 123.155 204.500 123.325 205.110 ;
        RECT 123.585 204.755 125.705 204.940 ;
        RECT 125.875 204.930 126.045 205.110 ;
        RECT 126.215 205.290 127.150 205.440 ;
        RECT 127.855 205.290 128.380 205.420 ;
        RECT 126.215 205.100 128.380 205.290 ;
        RECT 127.355 205.090 128.380 205.100 ;
        RECT 125.875 204.760 127.055 204.930 ;
        RECT 123.155 204.250 123.785 204.500 ;
        RECT 123.955 204.305 124.905 204.585 ;
        RECT 125.875 204.515 126.045 204.760 ;
        RECT 125.415 204.250 126.045 204.515 ;
        RECT 126.260 204.415 127.185 204.590 ;
        RECT 127.355 204.540 127.685 205.090 ;
        RECT 128.595 204.920 128.765 205.590 ;
        RECT 129.755 205.520 130.005 205.870 ;
        RECT 131.315 205.860 131.485 206.040 ;
        RECT 132.795 205.905 133.045 206.515 ;
        RECT 134.035 206.345 134.205 206.945 ;
        RECT 134.425 206.725 134.945 206.880 ;
        RECT 135.115 206.840 135.445 207.390 ;
        RECT 136.755 207.230 136.930 207.505 ;
        RECT 137.825 207.320 138.065 207.920 ;
        RECT 135.745 207.060 136.930 207.230 ;
        RECT 137.100 207.060 138.065 207.320 ;
        RECT 136.755 206.890 136.930 207.060 ;
        RECT 134.425 206.670 134.985 206.725 ;
        RECT 135.615 206.715 136.540 206.890 ;
        RECT 135.565 206.670 136.540 206.715 ;
        RECT 134.425 206.560 136.540 206.670 ;
        RECT 136.755 206.645 137.655 206.890 ;
        RECT 134.425 206.550 135.695 206.560 ;
        RECT 134.860 206.500 135.695 206.550 ;
        RECT 133.510 206.330 134.205 206.345 ;
        RECT 136.755 206.330 136.930 206.645 ;
        RECT 137.825 206.475 138.065 207.060 ;
        RECT 133.510 206.085 134.930 206.330 ;
        RECT 134.035 206.040 134.930 206.085 ;
        RECT 135.590 206.045 136.930 206.330 ;
        RECT 137.100 206.215 138.065 206.475 ;
        RECT 135.590 206.040 137.655 206.045 ;
        RECT 130.175 205.530 131.485 205.860 ;
        RECT 131.660 205.655 133.855 205.905 ;
        RECT 131.315 205.485 131.485 205.530 ;
        RECT 128.935 205.350 129.575 205.420 ;
        RECT 128.935 205.180 130.345 205.350 ;
        RECT 128.935 205.090 129.575 205.180 ;
        RECT 127.985 204.750 129.575 204.920 ;
        RECT 128.595 204.680 129.575 204.750 ;
        RECT 127.855 204.425 128.375 204.580 ;
        RECT 126.260 204.370 127.235 204.415 ;
        RECT 127.815 204.370 128.375 204.425 ;
        RECT 126.260 204.260 128.375 204.370 ;
        RECT 120.775 203.670 122.245 203.840 ;
        RECT 121.915 203.645 122.245 203.670 ;
        RECT 119.295 202.815 119.535 203.415 ;
        RECT 120.430 203.330 121.745 203.500 ;
        RECT 122.415 203.420 122.585 204.005 ;
        RECT 123.155 203.580 123.325 204.250 ;
        RECT 123.915 204.080 125.280 204.135 ;
        RECT 123.605 203.965 125.705 204.080 ;
        RECT 123.605 203.910 124.045 203.965 ;
        RECT 123.605 203.745 123.775 203.910 ;
        RECT 125.150 203.830 125.705 203.965 ;
        RECT 120.430 203.245 120.605 203.330 ;
        RECT 119.705 202.985 120.605 203.245 ;
        RECT 121.915 203.250 122.585 203.420 ;
        RECT 122.755 203.250 123.325 203.580 ;
        RECT 121.915 203.165 122.245 203.250 ;
        RECT 119.295 202.555 120.260 202.815 ;
        RECT 120.430 202.650 120.605 202.985 ;
        RECT 120.775 202.995 121.745 203.160 ;
        RECT 122.415 202.995 122.985 203.080 ;
        RECT 120.775 202.825 122.985 202.995 ;
        RECT 123.155 202.650 123.325 203.250 ;
        RECT 123.605 203.045 123.775 203.550 ;
        RECT 123.975 203.385 124.195 203.740 ;
        RECT 124.365 203.555 124.960 203.795 ;
        RECT 123.975 203.215 125.260 203.385 ;
        RECT 123.605 202.875 124.725 203.045 ;
        RECT 124.555 202.685 124.725 202.875 ;
        RECT 124.895 202.855 125.260 203.215 ;
        RECT 125.430 202.685 125.600 203.620 ;
        RECT 119.295 201.955 119.535 202.555 ;
        RECT 120.430 202.385 121.695 202.650 ;
        RECT 119.705 202.125 121.695 202.385 ;
        RECT 119.295 201.695 120.260 201.955 ;
        RECT 120.430 201.730 121.695 202.125 ;
        RECT 121.865 202.555 123.325 202.650 ;
        RECT 121.865 202.185 123.825 202.555 ;
        RECT 124.005 202.465 124.335 202.665 ;
        RECT 124.555 202.515 125.600 202.685 ;
        RECT 125.875 203.520 126.045 204.250 ;
        RECT 127.105 204.250 128.375 204.260 ;
        RECT 127.105 204.200 127.940 204.250 ;
        RECT 126.215 203.855 128.425 204.025 ;
        RECT 126.215 203.690 127.185 203.855 ;
        RECT 127.855 203.770 128.425 203.855 ;
        RECT 128.595 203.890 128.765 204.680 ;
        RECT 129.755 204.660 130.005 205.010 ;
        RECT 130.175 205.000 130.345 205.180 ;
        RECT 131.315 205.225 132.285 205.485 ;
        RECT 130.175 204.670 131.130 205.000 ;
        RECT 131.315 204.625 131.490 205.225 ;
        RECT 131.660 204.795 132.625 205.055 ;
        RECT 128.935 204.060 129.585 204.390 ;
        RECT 127.355 203.600 127.685 203.685 ;
        RECT 128.595 203.600 129.225 203.890 ;
        RECT 125.875 203.350 127.185 203.520 ;
        RECT 127.355 203.430 128.025 203.600 ;
        RECT 121.865 201.900 123.325 202.185 ;
        RECT 124.005 202.005 124.305 202.465 ;
        RECT 124.555 202.345 124.815 202.515 ;
        RECT 125.875 202.345 126.045 203.350 ;
        RECT 127.355 203.180 127.685 203.205 ;
        RECT 124.485 202.175 124.815 202.345 ;
        RECT 125.075 202.175 126.045 202.345 ;
        RECT 119.295 201.095 119.535 201.695 ;
        RECT 120.430 201.525 122.215 201.730 ;
        RECT 119.705 201.265 122.215 201.525 ;
        RECT 119.295 200.835 120.260 201.095 ;
        RECT 120.430 200.980 122.215 201.265 ;
        RECT 122.385 200.980 123.325 201.900 ;
        RECT 123.605 201.835 125.705 202.005 ;
        RECT 123.605 201.600 123.775 201.835 ;
        RECT 125.375 201.755 125.705 201.835 ;
        RECT 124.485 201.475 125.205 201.665 ;
        RECT 119.295 200.250 119.535 200.835 ;
        RECT 120.430 200.665 120.605 200.980 ;
        RECT 119.705 200.420 120.605 200.665 ;
        RECT 120.775 200.550 121.445 200.720 ;
        RECT 120.430 200.380 120.605 200.420 ;
        RECT 119.295 199.990 120.260 200.250 ;
        RECT 120.430 200.050 121.105 200.380 ;
        RECT 121.275 200.285 121.445 200.550 ;
        RECT 121.615 200.455 122.265 200.805 ;
        RECT 122.435 200.550 122.895 200.720 ;
        RECT 122.435 200.285 122.605 200.550 ;
        RECT 123.155 200.380 123.325 200.980 ;
        RECT 123.605 200.815 123.775 201.430 ;
        RECT 123.945 201.305 124.275 201.450 ;
        RECT 123.945 200.985 125.235 201.305 ;
        RECT 125.405 200.815 125.575 201.530 ;
        RECT 123.605 200.645 125.575 200.815 ;
        RECT 125.875 200.980 126.045 202.175 ;
        RECT 126.215 203.010 127.685 203.180 ;
        RECT 126.215 201.320 126.385 203.010 ;
        RECT 127.855 202.845 128.025 203.430 ;
        RECT 128.195 203.560 129.225 203.600 ;
        RECT 128.195 203.270 128.765 203.560 ;
        RECT 129.415 203.345 129.585 204.060 ;
        RECT 129.755 203.920 130.005 204.430 ;
        RECT 131.315 204.370 132.215 204.625 ;
        RECT 130.195 204.365 132.215 204.370 ;
        RECT 130.195 204.040 131.490 204.365 ;
        RECT 132.385 204.195 132.625 204.795 ;
        RECT 131.315 203.765 131.490 204.040 ;
        RECT 131.660 203.935 132.625 204.195 ;
        RECT 127.855 202.840 128.425 202.845 ;
        RECT 126.555 202.670 128.425 202.840 ;
        RECT 126.555 201.715 126.725 202.670 ;
        RECT 126.895 202.330 127.865 202.500 ;
        RECT 126.895 201.680 127.065 202.330 ;
        RECT 128.060 202.315 128.425 202.670 ;
        RECT 128.595 202.815 128.765 203.270 ;
        RECT 128.935 203.015 129.585 203.345 ;
        RECT 129.755 203.340 131.070 203.710 ;
        RECT 131.315 203.505 132.215 203.765 ;
        RECT 128.595 202.485 129.225 202.815 ;
        RECT 127.405 202.125 127.575 202.130 ;
        RECT 127.265 201.850 128.425 202.125 ;
        RECT 126.895 201.490 128.425 201.680 ;
        RECT 128.595 201.320 128.765 202.485 ;
        RECT 129.415 202.260 129.585 203.015 ;
        RECT 129.755 202.840 131.070 203.170 ;
        RECT 131.315 202.905 131.490 203.505 ;
        RECT 132.385 203.335 132.625 203.935 ;
        RECT 131.660 203.075 132.625 203.335 ;
        RECT 131.315 202.645 132.215 202.905 ;
        RECT 129.755 202.300 131.070 202.630 ;
        RECT 129.095 202.090 129.585 202.260 ;
        RECT 128.950 201.590 129.585 201.920 ;
        RECT 129.755 201.710 129.965 202.130 ;
        RECT 131.315 202.045 131.490 202.645 ;
        RECT 132.385 202.475 132.625 203.075 ;
        RECT 131.660 202.215 132.625 202.475 ;
        RECT 130.135 201.780 131.145 202.030 ;
        RECT 131.315 201.800 132.215 202.045 ;
        RECT 129.395 201.540 129.585 201.590 ;
        RECT 130.135 201.540 130.425 201.780 ;
        RECT 131.315 201.610 131.490 201.800 ;
        RECT 132.385 201.630 132.625 202.215 ;
        RECT 126.215 201.150 127.240 201.320 ;
        RECT 128.595 201.310 129.225 201.320 ;
        RECT 125.875 200.810 126.805 200.980 ;
        RECT 121.275 200.055 122.605 200.285 ;
        RECT 122.775 200.370 123.325 200.380 ;
        RECT 122.775 200.160 123.855 200.370 ;
        RECT 122.775 200.050 123.325 200.160 ;
        RECT 119.295 199.390 119.535 199.990 ;
        RECT 120.430 199.805 120.605 200.050 ;
        RECT 119.705 199.560 120.605 199.805 ;
        RECT 120.775 199.695 122.895 199.880 ;
        RECT 120.430 199.455 120.605 199.560 ;
        RECT 119.295 199.130 120.260 199.390 ;
        RECT 120.430 199.190 121.065 199.455 ;
        RECT 121.575 199.245 122.525 199.525 ;
        RECT 123.155 199.440 123.325 200.050 ;
        RECT 124.235 199.940 124.565 200.645 ;
        RECT 124.770 199.920 125.145 200.475 ;
        RECT 125.875 200.465 126.045 200.810 ;
        RECT 125.375 200.150 126.045 200.465 ;
        RECT 123.540 199.770 124.065 199.900 ;
        RECT 124.770 199.770 125.705 199.920 ;
        RECT 123.540 199.580 125.705 199.770 ;
        RECT 123.540 199.570 124.565 199.580 ;
        RECT 122.695 199.400 123.325 199.440 ;
        RECT 122.695 199.230 123.935 199.400 ;
        RECT 122.695 199.190 123.325 199.230 ;
        RECT 119.295 198.530 119.535 199.130 ;
        RECT 120.430 198.945 120.605 199.190 ;
        RECT 121.200 199.020 122.565 199.075 ;
        RECT 119.705 198.700 120.605 198.945 ;
        RECT 120.775 198.905 122.875 199.020 ;
        RECT 120.775 198.770 121.330 198.905 ;
        RECT 122.435 198.850 122.875 198.905 ;
        RECT 119.295 198.270 120.260 198.530 ;
        RECT 119.295 198.095 119.520 198.270 ;
        RECT 117.715 198.080 118.365 198.090 ;
        RECT 114.495 197.850 116.305 198.000 ;
        RECT 116.475 197.910 117.145 198.080 ;
        RECT 114.995 197.830 116.305 197.850 ;
        RECT 112.660 197.470 113.185 197.600 ;
        RECT 113.890 197.470 114.825 197.620 ;
        RECT 112.660 197.280 114.825 197.470 ;
        RECT 112.660 197.270 113.685 197.280 ;
        RECT 90.745 196.005 91.955 197.095 ;
        RECT 112.275 196.930 113.055 197.100 ;
        RECT 112.275 196.205 112.445 196.930 ;
        RECT 112.665 196.605 113.185 196.760 ;
        RECT 113.355 196.720 113.685 197.270 ;
        RECT 114.995 197.110 115.165 197.830 ;
        RECT 116.475 197.660 116.805 197.685 ;
        RECT 113.985 196.940 115.165 197.110 ;
        RECT 112.665 196.550 113.225 196.605 ;
        RECT 113.855 196.595 114.780 196.770 ;
        RECT 113.805 196.550 114.780 196.595 ;
        RECT 112.665 196.440 114.780 196.550 ;
        RECT 112.665 196.430 113.935 196.440 ;
        RECT 113.100 196.380 113.935 196.430 ;
        RECT 114.995 196.205 115.165 196.940 ;
        RECT 13.380 195.835 92.040 196.005 ;
        RECT 112.275 195.945 113.285 196.205 ;
        RECT 113.845 195.945 115.165 196.205 ;
        RECT 13.465 194.745 14.675 195.835 ;
        RECT 14.845 195.400 20.190 195.835 ;
        RECT 20.365 195.400 25.710 195.835 ;
        RECT 13.465 194.035 13.985 194.575 ;
        RECT 14.155 194.205 14.675 194.745 ;
        RECT 13.465 193.285 14.675 194.035 ;
        RECT 16.430 193.830 16.770 194.660 ;
        RECT 18.250 194.150 18.600 195.400 ;
        RECT 21.950 193.830 22.290 194.660 ;
        RECT 23.770 194.150 24.120 195.400 ;
        RECT 26.345 194.670 26.635 195.835 ;
        RECT 26.805 195.400 32.150 195.835 ;
        RECT 32.325 195.400 37.670 195.835 ;
        RECT 14.845 193.285 20.190 193.830 ;
        RECT 20.365 193.285 25.710 193.830 ;
        RECT 26.345 193.285 26.635 194.010 ;
        RECT 28.390 193.830 28.730 194.660 ;
        RECT 30.210 194.150 30.560 195.400 ;
        RECT 33.910 193.830 34.250 194.660 ;
        RECT 35.730 194.150 36.080 195.400 ;
        RECT 38.395 195.165 38.565 195.665 ;
        RECT 38.735 195.335 39.065 195.835 ;
        RECT 38.395 194.995 39.060 195.165 ;
        RECT 38.310 194.175 38.660 194.825 ;
        RECT 38.830 194.005 39.060 194.995 ;
        RECT 38.395 193.835 39.060 194.005 ;
        RECT 26.805 193.285 32.150 193.830 ;
        RECT 32.325 193.285 37.670 193.830 ;
        RECT 38.395 193.545 38.565 193.835 ;
        RECT 38.735 193.285 39.065 193.665 ;
        RECT 39.235 193.545 39.420 195.665 ;
        RECT 39.660 195.375 39.925 195.835 ;
        RECT 40.095 195.240 40.345 195.665 ;
        RECT 40.555 195.390 41.660 195.560 ;
        RECT 40.040 195.110 40.345 195.240 ;
        RECT 39.590 193.915 39.870 194.865 ;
        RECT 40.040 194.005 40.210 195.110 ;
        RECT 40.380 194.325 40.620 194.920 ;
        RECT 40.790 194.855 41.320 195.220 ;
        RECT 40.790 194.155 40.960 194.855 ;
        RECT 41.490 194.775 41.660 195.390 ;
        RECT 41.830 195.035 42.000 195.835 ;
        RECT 42.170 195.335 42.420 195.665 ;
        RECT 42.645 195.365 43.530 195.535 ;
        RECT 41.490 194.685 42.000 194.775 ;
        RECT 40.040 193.875 40.265 194.005 ;
        RECT 40.435 193.935 40.960 194.155 ;
        RECT 41.130 194.515 42.000 194.685 ;
        RECT 39.675 193.285 39.925 193.745 ;
        RECT 40.095 193.735 40.265 193.875 ;
        RECT 41.130 193.735 41.300 194.515 ;
        RECT 41.830 194.445 42.000 194.515 ;
        RECT 41.510 194.265 41.710 194.295 ;
        RECT 42.170 194.265 42.340 195.335 ;
        RECT 42.510 194.445 42.700 195.165 ;
        RECT 41.510 193.965 42.340 194.265 ;
        RECT 42.870 194.235 43.190 195.195 ;
        RECT 40.095 193.565 40.430 193.735 ;
        RECT 40.625 193.565 41.300 193.735 ;
        RECT 41.620 193.285 41.990 193.785 ;
        RECT 42.170 193.735 42.340 193.965 ;
        RECT 42.725 193.905 43.190 194.235 ;
        RECT 43.360 194.525 43.530 195.365 ;
        RECT 43.710 195.335 44.025 195.835 ;
        RECT 44.255 195.105 44.595 195.665 ;
        RECT 43.700 194.730 44.595 195.105 ;
        RECT 44.765 194.825 44.935 195.835 ;
        RECT 44.405 194.525 44.595 194.730 ;
        RECT 45.105 194.775 45.435 195.620 ;
        RECT 46.125 194.965 46.400 195.665 ;
        RECT 46.570 195.290 46.825 195.835 ;
        RECT 46.995 195.325 47.475 195.665 ;
        RECT 47.650 195.280 48.255 195.835 ;
        RECT 47.640 195.180 48.255 195.280 ;
        RECT 47.640 195.155 47.825 195.180 ;
        RECT 45.105 194.695 45.495 194.775 ;
        RECT 45.280 194.645 45.495 194.695 ;
        RECT 43.360 194.195 44.235 194.525 ;
        RECT 44.405 194.195 45.155 194.525 ;
        RECT 43.360 193.735 43.530 194.195 ;
        RECT 44.405 194.025 44.605 194.195 ;
        RECT 45.325 194.065 45.495 194.645 ;
        RECT 45.270 194.025 45.495 194.065 ;
        RECT 42.170 193.565 42.575 193.735 ;
        RECT 42.745 193.565 43.530 193.735 ;
        RECT 43.805 193.285 44.015 193.815 ;
        RECT 44.275 193.500 44.605 194.025 ;
        RECT 45.115 193.940 45.495 194.025 ;
        RECT 44.775 193.285 44.945 193.895 ;
        RECT 45.115 193.505 45.445 193.940 ;
        RECT 46.125 193.935 46.295 194.965 ;
        RECT 46.570 194.835 47.325 195.085 ;
        RECT 47.495 194.910 47.825 195.155 ;
        RECT 46.570 194.800 47.340 194.835 ;
        RECT 46.570 194.790 47.355 194.800 ;
        RECT 46.465 194.775 47.360 194.790 ;
        RECT 46.465 194.760 47.380 194.775 ;
        RECT 46.465 194.750 47.400 194.760 ;
        RECT 46.465 194.740 47.425 194.750 ;
        RECT 46.465 194.710 47.495 194.740 ;
        RECT 46.465 194.680 47.515 194.710 ;
        RECT 46.465 194.650 47.535 194.680 ;
        RECT 46.465 194.625 47.565 194.650 ;
        RECT 46.465 194.590 47.600 194.625 ;
        RECT 46.465 194.585 47.630 194.590 ;
        RECT 46.465 194.190 46.695 194.585 ;
        RECT 47.240 194.580 47.630 194.585 ;
        RECT 47.265 194.570 47.630 194.580 ;
        RECT 47.280 194.565 47.630 194.570 ;
        RECT 47.295 194.560 47.630 194.565 ;
        RECT 47.995 194.560 48.255 195.010 ;
        RECT 48.435 194.865 48.765 195.650 ;
        RECT 48.435 194.695 49.115 194.865 ;
        RECT 49.295 194.695 49.625 195.835 ;
        RECT 49.805 195.280 50.410 195.835 ;
        RECT 50.585 195.325 51.065 195.665 ;
        RECT 51.235 195.290 51.490 195.835 ;
        RECT 49.805 195.180 50.420 195.280 ;
        RECT 50.235 195.155 50.420 195.180 ;
        RECT 47.295 194.555 48.255 194.560 ;
        RECT 47.305 194.545 48.255 194.555 ;
        RECT 47.315 194.540 48.255 194.545 ;
        RECT 47.325 194.530 48.255 194.540 ;
        RECT 47.330 194.520 48.255 194.530 ;
        RECT 47.335 194.515 48.255 194.520 ;
        RECT 47.345 194.500 48.255 194.515 ;
        RECT 47.350 194.485 48.255 194.500 ;
        RECT 47.360 194.460 48.255 194.485 ;
        RECT 46.865 193.990 47.195 194.415 ;
        RECT 46.125 193.455 46.385 193.935 ;
        RECT 46.555 193.285 46.805 193.825 ;
        RECT 46.975 193.505 47.195 193.990 ;
        RECT 47.365 194.390 48.255 194.460 ;
        RECT 47.365 193.665 47.535 194.390 ;
        RECT 48.425 194.275 48.775 194.525 ;
        RECT 47.705 193.835 48.255 194.220 ;
        RECT 48.945 194.095 49.115 194.695 ;
        RECT 49.805 194.560 50.065 195.010 ;
        RECT 50.235 194.910 50.565 195.155 ;
        RECT 50.735 194.835 51.490 195.085 ;
        RECT 51.660 194.965 51.935 195.665 ;
        RECT 50.720 194.800 51.490 194.835 ;
        RECT 50.705 194.790 51.490 194.800 ;
        RECT 50.700 194.775 51.595 194.790 ;
        RECT 50.680 194.760 51.595 194.775 ;
        RECT 50.660 194.750 51.595 194.760 ;
        RECT 50.635 194.740 51.595 194.750 ;
        RECT 50.565 194.710 51.595 194.740 ;
        RECT 50.545 194.680 51.595 194.710 ;
        RECT 50.525 194.650 51.595 194.680 ;
        RECT 50.495 194.625 51.595 194.650 ;
        RECT 50.460 194.590 51.595 194.625 ;
        RECT 50.430 194.585 51.595 194.590 ;
        RECT 50.430 194.580 50.820 194.585 ;
        RECT 50.430 194.570 50.795 194.580 ;
        RECT 50.430 194.565 50.780 194.570 ;
        RECT 50.430 194.560 50.765 194.565 ;
        RECT 49.805 194.555 50.765 194.560 ;
        RECT 49.805 194.545 50.755 194.555 ;
        RECT 49.805 194.540 50.745 194.545 ;
        RECT 49.805 194.530 50.735 194.540 ;
        RECT 49.285 194.275 49.635 194.525 ;
        RECT 49.805 194.520 50.730 194.530 ;
        RECT 49.805 194.515 50.725 194.520 ;
        RECT 49.805 194.500 50.715 194.515 ;
        RECT 49.805 194.485 50.710 194.500 ;
        RECT 49.805 194.460 50.700 194.485 ;
        RECT 49.805 194.390 50.695 194.460 ;
        RECT 47.365 193.495 48.255 193.665 ;
        RECT 48.445 193.285 48.685 194.095 ;
        RECT 48.855 193.455 49.185 194.095 ;
        RECT 49.355 193.285 49.625 194.095 ;
        RECT 49.805 193.835 50.355 194.220 ;
        RECT 50.525 193.665 50.695 194.390 ;
        RECT 49.805 193.495 50.695 193.665 ;
        RECT 50.865 193.990 51.195 194.415 ;
        RECT 51.365 194.190 51.595 194.585 ;
        RECT 50.865 193.505 51.085 193.990 ;
        RECT 51.765 193.935 51.935 194.965 ;
        RECT 52.105 194.670 52.395 195.835 ;
        RECT 52.655 195.165 52.825 195.665 ;
        RECT 52.995 195.335 53.325 195.835 ;
        RECT 52.655 194.995 53.320 195.165 ;
        RECT 52.570 194.175 52.920 194.825 ;
        RECT 51.255 193.285 51.505 193.825 ;
        RECT 51.675 193.455 51.935 193.935 ;
        RECT 52.105 193.285 52.395 194.010 ;
        RECT 53.090 194.005 53.320 194.995 ;
        RECT 52.655 193.835 53.320 194.005 ;
        RECT 52.655 193.545 52.825 193.835 ;
        RECT 52.995 193.285 53.325 193.665 ;
        RECT 53.495 193.545 53.680 195.665 ;
        RECT 53.920 195.375 54.185 195.835 ;
        RECT 54.355 195.240 54.605 195.665 ;
        RECT 54.815 195.390 55.920 195.560 ;
        RECT 54.300 195.110 54.605 195.240 ;
        RECT 53.850 193.915 54.130 194.865 ;
        RECT 54.300 194.005 54.470 195.110 ;
        RECT 54.640 194.325 54.880 194.920 ;
        RECT 55.050 194.855 55.580 195.220 ;
        RECT 55.050 194.155 55.220 194.855 ;
        RECT 55.750 194.775 55.920 195.390 ;
        RECT 56.090 195.035 56.260 195.835 ;
        RECT 56.430 195.335 56.680 195.665 ;
        RECT 56.905 195.365 57.790 195.535 ;
        RECT 55.750 194.685 56.260 194.775 ;
        RECT 54.300 193.875 54.525 194.005 ;
        RECT 54.695 193.935 55.220 194.155 ;
        RECT 55.390 194.515 56.260 194.685 ;
        RECT 53.935 193.285 54.185 193.745 ;
        RECT 54.355 193.735 54.525 193.875 ;
        RECT 55.390 193.735 55.560 194.515 ;
        RECT 56.090 194.445 56.260 194.515 ;
        RECT 55.770 194.265 55.970 194.295 ;
        RECT 56.430 194.265 56.600 195.335 ;
        RECT 56.770 194.445 56.960 195.165 ;
        RECT 55.770 193.965 56.600 194.265 ;
        RECT 57.130 194.235 57.450 195.195 ;
        RECT 54.355 193.565 54.690 193.735 ;
        RECT 54.885 193.565 55.560 193.735 ;
        RECT 55.880 193.285 56.250 193.785 ;
        RECT 56.430 193.735 56.600 193.965 ;
        RECT 56.985 193.905 57.450 194.235 ;
        RECT 57.620 194.525 57.790 195.365 ;
        RECT 57.970 195.335 58.285 195.835 ;
        RECT 58.515 195.105 58.855 195.665 ;
        RECT 57.960 194.730 58.855 195.105 ;
        RECT 59.025 194.825 59.195 195.835 ;
        RECT 58.665 194.525 58.855 194.730 ;
        RECT 59.365 194.775 59.695 195.620 ;
        RECT 59.365 194.695 59.755 194.775 ;
        RECT 60.855 194.695 61.185 195.835 ;
        RECT 61.715 194.865 62.045 195.650 ;
        RECT 61.365 194.695 62.045 194.865 ;
        RECT 63.155 194.695 63.485 195.835 ;
        RECT 64.015 194.865 64.345 195.650 ;
        RECT 63.665 194.695 64.345 194.865 ;
        RECT 64.525 194.745 65.735 195.835 ;
        RECT 59.540 194.645 59.755 194.695 ;
        RECT 57.620 194.195 58.495 194.525 ;
        RECT 58.665 194.195 59.415 194.525 ;
        RECT 57.620 193.735 57.790 194.195 ;
        RECT 58.665 194.025 58.865 194.195 ;
        RECT 59.585 194.065 59.755 194.645 ;
        RECT 60.845 194.275 61.195 194.525 ;
        RECT 61.365 194.095 61.535 194.695 ;
        RECT 61.705 194.275 62.055 194.525 ;
        RECT 63.145 194.275 63.495 194.525 ;
        RECT 63.665 194.095 63.835 194.695 ;
        RECT 64.005 194.275 64.355 194.525 ;
        RECT 59.530 194.025 59.755 194.065 ;
        RECT 56.430 193.565 56.835 193.735 ;
        RECT 57.005 193.565 57.790 193.735 ;
        RECT 58.065 193.285 58.275 193.815 ;
        RECT 58.535 193.500 58.865 194.025 ;
        RECT 59.375 193.940 59.755 194.025 ;
        RECT 59.035 193.285 59.205 193.895 ;
        RECT 59.375 193.505 59.705 193.940 ;
        RECT 60.855 193.285 61.125 194.095 ;
        RECT 61.295 193.455 61.625 194.095 ;
        RECT 61.795 193.285 62.035 194.095 ;
        RECT 63.155 193.285 63.425 194.095 ;
        RECT 63.595 193.455 63.925 194.095 ;
        RECT 64.095 193.285 64.335 194.095 ;
        RECT 64.525 194.035 65.045 194.575 ;
        RECT 65.215 194.205 65.735 194.745 ;
        RECT 65.915 194.695 66.245 195.835 ;
        RECT 66.775 194.865 67.105 195.650 ;
        RECT 67.285 195.280 67.890 195.835 ;
        RECT 68.065 195.325 68.545 195.665 ;
        RECT 68.715 195.290 68.970 195.835 ;
        RECT 67.285 195.180 67.900 195.280 ;
        RECT 67.715 195.155 67.900 195.180 ;
        RECT 66.425 194.695 67.105 194.865 ;
        RECT 65.905 194.275 66.255 194.525 ;
        RECT 66.425 194.095 66.595 194.695 ;
        RECT 67.285 194.560 67.545 195.010 ;
        RECT 67.715 194.910 68.045 195.155 ;
        RECT 68.215 194.835 68.970 195.085 ;
        RECT 69.140 194.965 69.415 195.665 ;
        RECT 68.200 194.800 68.970 194.835 ;
        RECT 68.185 194.790 68.970 194.800 ;
        RECT 68.180 194.775 69.075 194.790 ;
        RECT 68.160 194.760 69.075 194.775 ;
        RECT 68.140 194.750 69.075 194.760 ;
        RECT 68.115 194.740 69.075 194.750 ;
        RECT 68.045 194.710 69.075 194.740 ;
        RECT 68.025 194.680 69.075 194.710 ;
        RECT 68.005 194.650 69.075 194.680 ;
        RECT 67.975 194.625 69.075 194.650 ;
        RECT 67.940 194.590 69.075 194.625 ;
        RECT 67.910 194.585 69.075 194.590 ;
        RECT 67.910 194.580 68.300 194.585 ;
        RECT 67.910 194.570 68.275 194.580 ;
        RECT 67.910 194.565 68.260 194.570 ;
        RECT 67.910 194.560 68.245 194.565 ;
        RECT 67.285 194.555 68.245 194.560 ;
        RECT 67.285 194.545 68.235 194.555 ;
        RECT 67.285 194.540 68.225 194.545 ;
        RECT 67.285 194.530 68.215 194.540 ;
        RECT 66.765 194.275 67.115 194.525 ;
        RECT 67.285 194.520 68.210 194.530 ;
        RECT 67.285 194.515 68.205 194.520 ;
        RECT 67.285 194.500 68.195 194.515 ;
        RECT 67.285 194.485 68.190 194.500 ;
        RECT 67.285 194.460 68.180 194.485 ;
        RECT 67.285 194.390 68.175 194.460 ;
        RECT 64.525 193.285 65.735 194.035 ;
        RECT 65.915 193.285 66.185 194.095 ;
        RECT 66.355 193.455 66.685 194.095 ;
        RECT 66.855 193.285 67.095 194.095 ;
        RECT 67.285 193.835 67.835 194.220 ;
        RECT 68.005 193.665 68.175 194.390 ;
        RECT 67.285 193.495 68.175 193.665 ;
        RECT 68.345 193.990 68.675 194.415 ;
        RECT 68.845 194.190 69.075 194.585 ;
        RECT 68.345 193.505 68.565 193.990 ;
        RECT 69.245 193.935 69.415 194.965 ;
        RECT 70.565 194.775 70.895 195.620 ;
        RECT 71.065 194.825 71.235 195.835 ;
        RECT 71.405 195.105 71.745 195.665 ;
        RECT 71.975 195.335 72.290 195.835 ;
        RECT 72.470 195.365 73.355 195.535 ;
        RECT 70.505 194.695 70.895 194.775 ;
        RECT 71.405 194.730 72.300 195.105 ;
        RECT 70.505 194.645 70.720 194.695 ;
        RECT 70.505 194.065 70.675 194.645 ;
        RECT 71.405 194.525 71.595 194.730 ;
        RECT 72.470 194.525 72.640 195.365 ;
        RECT 73.580 195.335 73.830 195.665 ;
        RECT 70.845 194.195 71.595 194.525 ;
        RECT 71.765 194.195 72.640 194.525 ;
        RECT 70.505 194.025 70.730 194.065 ;
        RECT 71.395 194.025 71.595 194.195 ;
        RECT 70.505 193.940 70.885 194.025 ;
        RECT 68.735 193.285 68.985 193.825 ;
        RECT 69.155 193.455 69.415 193.935 ;
        RECT 70.555 193.505 70.885 193.940 ;
        RECT 71.055 193.285 71.225 193.895 ;
        RECT 71.395 193.500 71.725 194.025 ;
        RECT 71.985 193.285 72.195 193.815 ;
        RECT 72.470 193.735 72.640 194.195 ;
        RECT 72.810 194.235 73.130 195.195 ;
        RECT 73.300 194.445 73.490 195.165 ;
        RECT 73.660 194.265 73.830 195.335 ;
        RECT 74.000 195.035 74.170 195.835 ;
        RECT 74.340 195.390 75.445 195.560 ;
        RECT 74.340 194.775 74.510 195.390 ;
        RECT 75.655 195.240 75.905 195.665 ;
        RECT 76.075 195.375 76.340 195.835 ;
        RECT 74.680 194.855 75.210 195.220 ;
        RECT 75.655 195.110 75.960 195.240 ;
        RECT 74.000 194.685 74.510 194.775 ;
        RECT 74.000 194.515 74.870 194.685 ;
        RECT 74.000 194.445 74.170 194.515 ;
        RECT 74.290 194.265 74.490 194.295 ;
        RECT 72.810 193.905 73.275 194.235 ;
        RECT 73.660 193.965 74.490 194.265 ;
        RECT 73.660 193.735 73.830 193.965 ;
        RECT 72.470 193.565 73.255 193.735 ;
        RECT 73.425 193.565 73.830 193.735 ;
        RECT 74.010 193.285 74.380 193.785 ;
        RECT 74.700 193.735 74.870 194.515 ;
        RECT 75.040 194.155 75.210 194.855 ;
        RECT 75.380 194.325 75.620 194.920 ;
        RECT 75.040 193.935 75.565 194.155 ;
        RECT 75.790 194.005 75.960 195.110 ;
        RECT 75.735 193.875 75.960 194.005 ;
        RECT 76.130 193.915 76.410 194.865 ;
        RECT 75.735 193.735 75.905 193.875 ;
        RECT 74.700 193.565 75.375 193.735 ;
        RECT 75.570 193.565 75.905 193.735 ;
        RECT 76.075 193.285 76.325 193.745 ;
        RECT 76.580 193.545 76.765 195.665 ;
        RECT 76.935 195.335 77.265 195.835 ;
        RECT 77.435 195.165 77.605 195.665 ;
        RECT 76.940 194.995 77.605 195.165 ;
        RECT 76.940 194.005 77.170 194.995 ;
        RECT 77.340 194.175 77.690 194.825 ;
        RECT 77.865 194.670 78.155 195.835 ;
        RECT 78.325 195.400 83.670 195.835 ;
        RECT 83.845 195.400 89.190 195.835 ;
        RECT 76.940 193.835 77.605 194.005 ;
        RECT 76.935 193.285 77.265 193.665 ;
        RECT 77.435 193.545 77.605 193.835 ;
        RECT 77.865 193.285 78.155 194.010 ;
        RECT 79.910 193.830 80.250 194.660 ;
        RECT 81.730 194.150 82.080 195.400 ;
        RECT 85.430 193.830 85.770 194.660 ;
        RECT 87.250 194.150 87.600 195.400 ;
        RECT 89.365 194.745 90.575 195.835 ;
        RECT 89.365 194.035 89.885 194.575 ;
        RECT 90.055 194.205 90.575 194.745 ;
        RECT 90.745 194.745 91.955 195.835 ;
        RECT 112.275 195.345 112.445 195.945 ;
        RECT 112.615 195.600 114.825 195.770 ;
        RECT 112.615 195.515 113.190 195.600 ;
        RECT 113.920 195.515 114.825 195.600 ;
        RECT 114.995 195.460 115.165 195.945 ;
        RECT 115.335 197.490 116.805 197.660 ;
        RECT 115.335 195.800 115.505 197.490 ;
        RECT 116.975 197.325 117.145 197.910 ;
        RECT 117.315 197.830 118.365 198.080 ;
        RECT 117.315 197.750 117.885 197.830 ;
        RECT 116.975 197.320 117.545 197.325 ;
        RECT 115.675 197.150 117.545 197.320 ;
        RECT 115.675 196.195 115.845 197.150 ;
        RECT 116.015 196.810 116.985 196.980 ;
        RECT 116.015 196.160 116.185 196.810 ;
        RECT 117.180 196.795 117.545 197.150 ;
        RECT 117.715 197.230 117.885 197.750 ;
        RECT 118.535 197.660 119.520 198.095 ;
        RECT 120.430 198.085 120.605 198.700 ;
        RECT 119.705 197.830 120.605 198.085 ;
        RECT 118.080 197.400 120.260 197.660 ;
        RECT 118.535 197.370 120.260 197.400 ;
        RECT 117.715 196.930 118.365 197.230 ;
        RECT 118.535 196.930 119.520 197.370 ;
        RECT 120.435 197.285 120.605 197.830 ;
        RECT 120.880 197.625 121.050 198.560 ;
        RECT 121.520 198.495 122.115 198.735 ;
        RECT 122.705 198.685 122.875 198.850 ;
        RECT 122.285 198.325 122.505 198.680 ;
        RECT 123.155 198.500 123.325 199.190 ;
        RECT 123.545 198.905 124.065 199.060 ;
        RECT 124.235 199.020 124.565 199.570 ;
        RECT 125.875 199.410 126.045 200.150 ;
        RECT 126.395 200.400 126.805 200.575 ;
        RECT 127.050 200.570 127.240 201.150 ;
        RECT 127.615 200.580 127.785 201.290 ;
        RECT 128.060 201.150 129.225 201.310 ;
        RECT 129.395 201.280 130.425 201.540 ;
        RECT 130.595 201.280 131.490 201.610 ;
        RECT 131.660 201.370 132.625 201.630 ;
        RECT 129.395 201.170 129.965 201.280 ;
        RECT 128.060 200.800 128.765 201.150 ;
        RECT 129.755 200.960 129.965 201.170 ;
        RECT 131.315 201.185 131.490 201.280 ;
        RECT 127.615 200.400 128.390 200.580 ;
        RECT 126.395 200.335 128.390 200.400 ;
        RECT 126.395 200.060 127.785 200.335 ;
        RECT 126.215 199.610 128.425 199.890 ;
        RECT 126.215 199.505 127.185 199.610 ;
        RECT 127.855 199.505 128.425 199.610 ;
        RECT 128.595 199.795 128.765 200.800 ;
        RECT 128.935 200.790 129.565 200.860 ;
        RECT 130.135 200.790 131.145 201.045 ;
        RECT 128.935 200.520 131.145 200.790 ;
        RECT 131.315 200.940 132.215 201.185 ;
        RECT 128.935 200.070 131.145 200.350 ;
        RECT 128.935 199.965 129.505 200.070 ;
        RECT 130.175 199.965 131.145 200.070 ;
        RECT 131.315 200.325 131.490 200.940 ;
        RECT 132.385 200.770 132.625 201.370 ;
        RECT 131.660 200.510 132.625 200.770 ;
        RECT 131.315 200.080 132.215 200.325 ;
        RECT 129.675 199.795 130.005 199.900 ;
        RECT 131.315 199.795 131.490 200.080 ;
        RECT 132.385 199.910 132.625 200.510 ;
        RECT 128.595 199.470 129.225 199.795 ;
        RECT 124.865 199.335 126.045 199.410 ;
        RECT 127.355 199.335 127.685 199.440 ;
        RECT 128.595 199.335 128.765 199.470 ;
        RECT 124.865 199.240 126.505 199.335 ;
        RECT 123.545 198.850 124.105 198.905 ;
        RECT 124.735 198.895 125.660 199.070 ;
        RECT 124.685 198.850 125.660 198.895 ;
        RECT 123.545 198.740 125.660 198.850 ;
        RECT 125.875 199.010 126.505 199.240 ;
        RECT 123.545 198.730 124.815 198.740 ;
        RECT 123.980 198.680 124.815 198.730 ;
        RECT 121.220 198.155 122.505 198.325 ;
        RECT 121.220 197.795 121.585 198.155 ;
        RECT 122.705 197.985 122.875 198.490 ;
        RECT 121.755 197.815 122.875 197.985 ;
        RECT 123.155 198.170 123.830 198.500 ;
        RECT 124.685 198.445 124.855 198.450 ;
        RECT 121.755 197.625 121.925 197.815 ;
        RECT 120.880 197.455 121.925 197.625 ;
        RECT 121.665 197.285 121.925 197.455 ;
        RECT 122.145 197.405 122.475 197.605 ;
        RECT 123.155 197.495 123.325 198.170 ;
        RECT 124.005 198.145 124.855 198.445 ;
        RECT 125.025 198.250 125.685 198.420 ;
        RECT 123.520 197.975 123.895 198.000 ;
        RECT 125.025 197.975 125.255 198.250 ;
        RECT 125.875 198.080 126.045 199.010 ;
        RECT 126.675 198.885 127.965 199.335 ;
        RECT 128.135 199.010 128.765 199.335 ;
        RECT 126.675 198.490 126.895 198.885 ;
        RECT 126.215 198.210 126.895 198.490 ;
        RECT 123.520 197.760 125.255 197.975 ;
        RECT 120.435 197.200 121.405 197.285 ;
        RECT 119.690 197.115 121.405 197.200 ;
        RECT 121.665 197.115 121.995 197.285 ;
        RECT 119.690 196.930 120.605 197.115 ;
        RECT 122.175 196.945 122.475 197.405 ;
        RECT 122.655 197.125 123.325 197.495 ;
        RECT 124.045 197.740 125.255 197.760 ;
        RECT 125.425 197.750 126.045 198.080 ;
        RECT 127.065 198.020 127.625 198.715 ;
        RECT 127.795 198.490 127.965 198.885 ;
        RECT 127.795 198.210 128.425 198.490 ;
        RECT 123.510 197.310 123.850 197.480 ;
        RECT 124.045 197.420 124.375 197.740 ;
        RECT 117.715 196.670 117.885 196.930 ;
        RECT 120.435 196.670 120.605 196.930 ;
        RECT 120.775 196.775 122.875 196.945 ;
        RECT 120.775 196.695 121.105 196.775 ;
        RECT 116.525 196.605 116.695 196.610 ;
        RECT 116.385 196.330 117.545 196.605 ;
        RECT 116.015 195.970 117.545 196.160 ;
        RECT 117.715 196.150 119.175 196.670 ;
        RECT 115.335 195.630 116.360 195.800 ;
        RECT 117.715 195.790 118.635 196.150 ;
        RECT 119.345 195.980 120.605 196.670 ;
        RECT 113.355 195.345 113.685 195.430 ;
        RECT 114.995 195.345 115.925 195.460 ;
        RECT 112.275 195.015 112.825 195.345 ;
        RECT 112.995 195.175 114.065 195.345 ;
        RECT 90.745 194.205 91.265 194.745 ;
        RECT 91.435 194.035 91.955 194.575 ;
        RECT 78.325 193.285 83.670 193.830 ;
        RECT 83.845 193.285 89.190 193.830 ;
        RECT 89.365 193.285 90.575 194.035 ;
        RECT 90.745 193.285 91.955 194.035 ;
        RECT 112.275 193.450 112.445 195.015 ;
        RECT 112.995 194.800 113.165 195.175 ;
        RECT 112.615 194.630 113.165 194.800 ;
        RECT 113.345 194.540 113.715 194.895 ;
        RECT 113.895 194.800 114.065 195.175 ;
        RECT 114.235 195.290 115.925 195.345 ;
        RECT 114.235 195.015 115.165 195.290 ;
        RECT 113.895 194.630 114.825 194.800 ;
        RECT 114.995 193.450 115.165 195.015 ;
        RECT 115.515 194.880 115.925 195.055 ;
        RECT 116.170 195.050 116.360 195.630 ;
        RECT 116.735 195.060 116.905 195.770 ;
        RECT 117.180 195.460 118.635 195.790 ;
        RECT 118.805 195.460 120.605 195.980 ;
        RECT 120.905 195.755 121.075 196.470 ;
        RECT 121.275 196.415 121.995 196.605 ;
        RECT 122.705 196.540 122.875 196.775 ;
        RECT 123.155 196.720 123.325 197.125 ;
        RECT 123.655 197.250 123.850 197.310 ;
        RECT 124.545 197.265 125.660 197.550 ;
        RECT 124.545 197.250 124.715 197.265 ;
        RECT 123.655 197.080 124.715 197.250 ;
        RECT 125.875 197.220 126.045 197.750 ;
        RECT 126.215 197.620 128.425 198.020 ;
        RECT 128.595 197.680 128.765 199.010 ;
        RECT 129.395 199.345 130.685 199.795 ;
        RECT 130.855 199.470 131.490 199.795 ;
        RECT 131.660 199.650 132.625 199.910 ;
        RECT 129.395 198.950 129.565 199.345 ;
        RECT 128.935 198.670 129.565 198.950 ;
        RECT 129.735 198.480 130.295 199.175 ;
        RECT 130.465 198.950 130.685 199.345 ;
        RECT 131.315 199.465 131.490 199.470 ;
        RECT 132.400 199.475 132.625 199.650 ;
        RECT 132.795 199.645 133.045 205.655 ;
        RECT 134.035 205.485 134.205 206.040 ;
        RECT 134.465 205.610 134.925 205.780 ;
        RECT 133.475 205.440 134.205 205.485 ;
        RECT 133.475 205.225 134.585 205.440 ;
        RECT 134.035 205.110 134.585 205.225 ;
        RECT 134.755 205.345 134.925 205.610 ;
        RECT 135.095 205.515 135.745 205.865 ;
        RECT 136.755 205.785 137.655 206.040 ;
        RECT 135.915 205.610 136.585 205.780 ;
        RECT 135.915 205.345 136.085 205.610 ;
        RECT 136.755 205.440 136.930 205.785 ;
        RECT 137.825 205.615 138.065 206.215 ;
        RECT 134.755 205.115 136.085 205.345 ;
        RECT 136.255 205.185 136.930 205.440 ;
        RECT 137.100 205.355 138.065 205.615 ;
        RECT 136.255 205.110 137.655 205.185 ;
        RECT 133.215 204.795 133.840 205.055 ;
        RECT 133.215 204.195 133.385 204.795 ;
        RECT 134.035 204.625 134.205 205.110 ;
        RECT 134.465 204.755 136.585 204.940 ;
        RECT 136.755 204.925 137.655 205.110 ;
        RECT 133.555 204.500 134.205 204.625 ;
        RECT 133.555 204.365 134.665 204.500 ;
        RECT 134.035 204.250 134.665 204.365 ;
        RECT 134.835 204.305 135.785 204.585 ;
        RECT 136.755 204.515 136.930 204.925 ;
        RECT 137.825 204.755 138.065 205.355 ;
        RECT 136.295 204.325 136.930 204.515 ;
        RECT 137.100 204.495 138.065 204.755 ;
        RECT 136.295 204.250 137.655 204.325 ;
        RECT 133.215 203.935 133.840 204.195 ;
        RECT 133.215 203.335 133.385 203.935 ;
        RECT 134.035 203.765 134.205 204.250 ;
        RECT 134.795 204.080 136.160 204.135 ;
        RECT 133.555 203.505 134.205 203.765 ;
        RECT 134.485 203.965 136.585 204.080 ;
        RECT 134.485 203.910 134.925 203.965 ;
        RECT 134.485 203.745 134.655 203.910 ;
        RECT 136.030 203.830 136.585 203.965 ;
        RECT 136.755 204.065 137.655 204.250 ;
        RECT 133.215 203.075 133.840 203.335 ;
        RECT 133.215 202.490 133.385 203.075 ;
        RECT 134.035 202.905 134.205 203.505 ;
        RECT 133.555 202.660 134.205 202.905 ;
        RECT 134.485 203.045 134.655 203.550 ;
        RECT 134.855 203.385 135.075 203.740 ;
        RECT 135.245 203.555 135.840 203.795 ;
        RECT 134.855 203.215 136.140 203.385 ;
        RECT 134.485 202.875 135.605 203.045 ;
        RECT 135.435 202.685 135.605 202.875 ;
        RECT 135.775 202.855 136.140 203.215 ;
        RECT 136.310 202.685 136.480 203.620 ;
        RECT 134.035 202.555 134.205 202.660 ;
        RECT 133.215 202.215 133.840 202.490 ;
        RECT 133.215 201.630 133.385 202.215 ;
        RECT 134.035 202.185 134.705 202.555 ;
        RECT 134.885 202.465 135.215 202.665 ;
        RECT 135.435 202.515 136.480 202.685 ;
        RECT 136.755 203.465 136.930 204.065 ;
        RECT 137.825 203.895 138.065 204.495 ;
        RECT 137.100 203.635 138.065 203.895 ;
        RECT 136.755 203.205 137.725 203.465 ;
        RECT 136.755 202.605 136.925 203.205 ;
        RECT 138.235 203.035 138.485 209.045 ;
        RECT 138.655 209.040 138.825 209.215 ;
        RECT 138.655 208.780 139.280 209.040 ;
        RECT 138.655 208.180 138.825 208.780 ;
        RECT 139.475 208.610 139.645 209.220 ;
        RECT 140.275 209.465 141.565 209.915 ;
        RECT 141.735 209.590 142.365 209.915 ;
        RECT 143.425 209.855 143.685 210.025 ;
        RECT 143.935 209.905 144.235 210.365 ;
        RECT 144.915 210.185 145.085 210.585 ;
        RECT 145.995 210.500 146.325 210.585 ;
        RECT 140.275 209.070 140.445 209.465 ;
        RECT 139.815 208.790 140.445 209.070 ;
        RECT 138.995 208.360 139.645 208.610 ;
        RECT 140.615 208.600 141.175 209.295 ;
        RECT 141.345 209.070 141.565 209.465 ;
        RECT 141.345 208.790 142.025 209.070 ;
        RECT 138.655 207.920 139.280 208.180 ;
        RECT 138.655 207.320 138.825 207.920 ;
        RECT 139.475 207.800 139.645 208.360 ;
        RECT 139.815 208.200 142.025 208.600 ;
        RECT 142.195 208.120 142.365 209.590 ;
        RECT 142.640 209.685 143.685 209.855 ;
        RECT 143.905 209.705 144.235 209.905 ;
        RECT 144.415 209.985 145.085 210.185 ;
        RECT 145.255 210.330 145.830 210.415 ;
        RECT 146.560 210.330 147.465 210.415 ;
        RECT 145.255 210.160 147.465 210.330 ;
        RECT 147.635 209.985 147.805 210.585 ;
        RECT 144.415 209.815 145.925 209.985 ;
        RECT 144.915 209.725 145.925 209.815 ;
        RECT 146.485 209.725 147.805 209.985 ;
        RECT 142.640 208.750 142.810 209.685 ;
        RECT 142.980 209.155 143.345 209.515 ;
        RECT 143.515 209.495 143.685 209.685 ;
        RECT 143.515 209.325 144.635 209.495 ;
        RECT 142.980 208.985 144.265 209.155 ;
        RECT 143.280 208.575 143.875 208.815 ;
        RECT 144.045 208.630 144.265 208.985 ;
        RECT 144.465 208.820 144.635 209.325 ;
        RECT 142.535 208.405 143.090 208.540 ;
        RECT 144.465 208.460 144.635 208.625 ;
        RECT 144.195 208.405 144.635 208.460 ;
        RECT 142.535 208.290 144.635 208.405 ;
        RECT 144.915 208.490 145.085 209.725 ;
        RECT 145.255 209.380 146.665 209.550 ;
        RECT 147.635 209.540 147.805 209.725 ;
        RECT 145.255 209.060 145.825 209.380 ;
        RECT 145.255 208.660 145.825 208.890 ;
        RECT 145.995 208.805 146.325 209.210 ;
        RECT 146.495 209.030 146.665 209.380 ;
        RECT 146.835 209.210 147.805 209.540 ;
        RECT 146.495 208.780 147.465 209.030 ;
        RECT 142.960 208.235 144.325 208.290 ;
        RECT 144.915 208.120 145.485 208.490 ;
        RECT 140.275 207.820 141.565 208.030 ;
        RECT 139.475 207.750 140.105 207.800 ;
        RECT 138.995 207.530 140.105 207.750 ;
        RECT 138.995 207.500 139.645 207.530 ;
        RECT 138.655 207.060 139.280 207.320 ;
        RECT 138.655 206.475 138.825 207.060 ;
        RECT 139.475 206.890 139.645 207.500 ;
        RECT 140.275 207.360 140.445 207.820 ;
        RECT 139.815 207.075 140.445 207.360 ;
        RECT 140.615 206.960 141.175 207.650 ;
        RECT 141.345 207.360 141.565 207.820 ;
        RECT 142.195 207.855 142.825 208.120 ;
        RECT 144.455 208.070 145.485 208.120 ;
        RECT 142.195 207.800 142.365 207.855 ;
        RECT 141.735 207.530 142.365 207.800 ;
        RECT 143.335 207.785 144.285 208.065 ;
        RECT 144.455 207.870 145.085 208.070 ;
        RECT 145.655 207.900 145.825 208.660 ;
        RECT 145.995 208.340 147.125 208.590 ;
        RECT 141.345 207.075 142.025 207.360 ;
        RECT 142.195 207.260 142.365 207.530 ;
        RECT 142.535 207.430 144.655 207.615 ;
        RECT 144.915 207.560 145.085 207.870 ;
        RECT 145.255 207.730 145.825 207.900 ;
        RECT 145.995 207.940 147.125 208.140 ;
        RECT 145.995 207.895 146.325 207.940 ;
        RECT 147.295 207.770 147.465 208.780 ;
        RECT 144.915 207.260 145.825 207.560 ;
        RECT 145.995 207.320 146.275 207.710 ;
        RECT 146.445 207.600 147.465 207.770 ;
        RECT 138.995 206.645 139.645 206.890 ;
        RECT 138.655 206.200 139.280 206.475 ;
        RECT 139.475 206.330 139.645 206.645 ;
        RECT 142.195 206.930 142.865 207.260 ;
        RECT 143.035 207.025 144.365 207.255 ;
        RECT 142.195 206.330 142.365 206.930 ;
        RECT 143.035 206.760 143.205 207.025 ;
        RECT 142.535 206.590 143.205 206.760 ;
        RECT 143.375 206.505 144.025 206.855 ;
        RECT 144.195 206.760 144.365 207.025 ;
        RECT 144.535 207.110 145.825 207.260 ;
        RECT 146.445 207.150 146.615 207.600 ;
        RECT 147.635 207.430 147.805 209.210 ;
        RECT 144.535 206.930 145.085 207.110 ;
        RECT 145.995 206.980 146.615 207.150 ;
        RECT 146.785 207.115 147.805 207.430 ;
        RECT 144.195 206.590 144.655 206.760 ;
        RECT 138.655 205.615 138.825 206.200 ;
        RECT 139.475 206.040 140.370 206.330 ;
        RECT 141.030 206.040 142.365 206.330 ;
        RECT 144.915 206.330 145.085 206.930 ;
        RECT 145.265 206.810 145.825 206.940 ;
        RECT 146.835 206.810 147.465 206.940 ;
        RECT 145.265 206.500 147.465 206.810 ;
        RECT 147.635 206.330 147.805 207.115 ;
        RECT 142.535 206.070 143.205 206.240 ;
        RECT 139.475 206.030 139.645 206.040 ;
        RECT 138.995 205.785 139.645 206.030 ;
        RECT 142.195 205.900 142.365 206.040 ;
        RECT 138.655 205.355 139.280 205.615 ;
        RECT 139.475 205.440 139.645 205.785 ;
        RECT 139.815 205.695 142.025 205.865 ;
        RECT 139.815 205.610 140.385 205.695 ;
        RECT 141.055 205.530 142.025 205.695 ;
        RECT 142.195 205.570 142.865 205.900 ;
        RECT 143.035 205.805 143.205 206.070 ;
        RECT 143.375 205.975 144.025 206.325 ;
        RECT 144.195 206.070 144.655 206.240 ;
        RECT 144.195 205.805 144.365 206.070 ;
        RECT 144.915 206.040 145.810 206.330 ;
        RECT 146.470 206.040 147.805 206.330 ;
        RECT 144.915 205.900 145.085 206.040 ;
        RECT 143.035 205.575 144.365 205.805 ;
        RECT 144.535 205.570 145.085 205.900 ;
        RECT 140.555 205.440 140.885 205.525 ;
        RECT 138.655 204.755 138.825 205.355 ;
        RECT 139.475 205.185 140.045 205.440 ;
        RECT 138.995 205.110 140.045 205.185 ;
        RECT 140.215 205.270 140.885 205.440 ;
        RECT 142.195 205.360 142.365 205.570 ;
        RECT 138.995 204.925 139.645 205.110 ;
        RECT 138.655 204.495 139.280 204.755 ;
        RECT 138.655 203.895 138.825 204.495 ;
        RECT 139.475 204.325 139.645 204.925 ;
        RECT 140.215 204.685 140.385 205.270 ;
        RECT 141.055 205.190 142.365 205.360 ;
        RECT 142.535 205.215 144.655 205.400 ;
        RECT 140.555 205.020 140.885 205.045 ;
        RECT 140.555 204.850 142.025 205.020 ;
        RECT 138.995 204.065 139.645 204.325 ;
        RECT 139.815 204.680 140.385 204.685 ;
        RECT 139.815 204.510 141.685 204.680 ;
        RECT 139.815 204.155 140.180 204.510 ;
        RECT 140.375 204.170 141.345 204.340 ;
        RECT 138.655 203.635 139.280 203.895 ;
        RECT 139.475 203.465 139.645 204.065 ;
        RECT 140.665 203.965 140.835 203.970 ;
        RECT 139.815 203.690 140.975 203.965 ;
        RECT 141.175 203.520 141.345 204.170 ;
        RECT 141.515 203.555 141.685 204.510 ;
        RECT 138.915 203.205 139.645 203.465 ;
        RECT 139.815 203.330 141.345 203.520 ;
        RECT 139.475 203.150 139.645 203.205 ;
        RECT 141.855 203.160 142.025 204.850 ;
        RECT 137.100 202.785 139.295 203.035 ;
        RECT 134.035 202.045 134.205 202.185 ;
        RECT 133.555 201.800 134.205 202.045 ;
        RECT 134.885 202.005 135.185 202.465 ;
        RECT 135.435 202.345 135.695 202.515 ;
        RECT 136.755 202.345 137.735 202.605 ;
        RECT 135.365 202.175 135.695 202.345 ;
        RECT 135.955 202.175 136.925 202.345 ;
        RECT 133.215 201.370 133.840 201.630 ;
        RECT 133.215 200.770 133.385 201.370 ;
        RECT 134.035 201.190 134.205 201.800 ;
        RECT 134.485 201.835 136.585 202.005 ;
        RECT 134.485 201.600 134.655 201.835 ;
        RECT 136.255 201.755 136.585 201.835 ;
        RECT 136.755 201.745 136.925 202.175 ;
        RECT 138.235 202.175 138.485 202.785 ;
        RECT 139.475 202.640 140.180 203.150 ;
        RECT 139.475 202.605 139.645 202.640 ;
        RECT 138.950 202.345 139.645 202.605 ;
        RECT 140.455 202.420 140.625 203.130 ;
        RECT 138.235 202.170 139.295 202.175 ;
        RECT 137.095 201.925 139.295 202.170 ;
        RECT 135.365 201.475 136.085 201.665 ;
        RECT 133.555 200.940 134.205 201.190 ;
        RECT 133.215 200.510 133.840 200.770 ;
        RECT 133.215 199.910 133.385 200.510 ;
        RECT 134.035 200.370 134.205 200.940 ;
        RECT 134.485 200.815 134.655 201.430 ;
        RECT 134.825 201.305 135.155 201.450 ;
        RECT 134.825 200.985 136.115 201.305 ;
        RECT 136.285 200.815 136.455 201.530 ;
        RECT 134.485 200.645 136.455 200.815 ;
        RECT 136.755 201.450 137.735 201.745 ;
        RECT 136.755 200.715 136.925 201.450 ;
        RECT 138.235 201.440 138.795 201.755 ;
        RECT 139.475 201.745 139.645 202.345 ;
        RECT 139.850 202.240 140.625 202.420 ;
        RECT 141.000 202.990 142.025 203.160 ;
        RECT 142.195 204.975 142.365 205.190 ;
        RECT 142.195 204.710 142.825 204.975 ;
        RECT 143.335 204.765 144.285 205.045 ;
        RECT 144.915 204.960 145.085 205.570 ;
        RECT 144.455 204.710 145.085 204.960 ;
        RECT 141.000 202.410 141.190 202.990 ;
        RECT 142.195 202.820 142.365 204.710 ;
        RECT 142.960 204.540 144.325 204.595 ;
        RECT 142.535 204.425 144.635 204.540 ;
        RECT 142.535 204.290 143.090 204.425 ;
        RECT 144.195 204.370 144.635 204.425 ;
        RECT 142.640 203.145 142.810 204.080 ;
        RECT 143.280 204.015 143.875 204.255 ;
        RECT 144.465 204.205 144.635 204.370 ;
        RECT 144.915 204.380 145.085 204.710 ;
        RECT 145.255 204.550 145.885 204.835 ;
        RECT 144.045 203.845 144.265 204.200 ;
        RECT 144.915 204.110 145.545 204.380 ;
        RECT 142.980 203.675 144.265 203.845 ;
        RECT 142.980 203.315 143.345 203.675 ;
        RECT 144.465 203.505 144.635 204.010 ;
        RECT 143.515 203.335 144.635 203.505 ;
        RECT 143.515 203.145 143.685 203.335 ;
        RECT 142.640 202.975 143.685 203.145 ;
        RECT 141.435 202.805 142.365 202.820 ;
        RECT 143.425 202.805 143.685 202.975 ;
        RECT 143.905 202.925 144.235 203.125 ;
        RECT 144.915 203.015 145.085 204.110 ;
        RECT 145.715 204.090 145.885 204.550 ;
        RECT 146.055 204.260 146.615 204.950 ;
        RECT 146.785 204.550 147.465 204.835 ;
        RECT 146.785 204.090 147.005 204.550 ;
        RECT 147.635 204.380 147.805 206.040 ;
        RECT 147.175 204.110 147.805 204.380 ;
        RECT 145.715 203.880 147.005 204.090 ;
        RECT 145.255 203.310 147.465 203.710 ;
        RECT 141.435 202.650 143.165 202.805 ;
        RECT 142.195 202.635 143.165 202.650 ;
        RECT 143.425 202.635 143.755 202.805 ;
        RECT 141.435 202.240 141.845 202.415 ;
        RECT 139.850 202.175 141.845 202.240 ;
        RECT 140.455 201.900 141.845 202.175 ;
        RECT 138.965 201.440 139.645 201.745 ;
        RECT 137.095 200.990 139.305 201.270 ;
        RECT 137.095 200.885 138.065 200.990 ;
        RECT 138.735 200.885 139.305 200.990 ;
        RECT 139.475 201.105 139.645 201.440 ;
        RECT 139.475 200.865 140.155 201.105 ;
        RECT 138.235 200.715 138.565 200.820 ;
        RECT 139.475 200.715 139.645 200.865 ;
        RECT 140.325 200.855 140.885 201.210 ;
        RECT 134.035 200.330 134.735 200.370 ;
        RECT 133.555 200.160 134.735 200.330 ;
        RECT 133.555 200.080 134.205 200.160 ;
        RECT 133.215 199.650 133.840 199.910 ;
        RECT 133.215 199.475 133.385 199.650 ;
        RECT 131.315 199.210 132.215 199.465 ;
        RECT 130.465 198.670 131.145 198.950 ;
        RECT 131.315 198.580 131.485 199.210 ;
        RECT 132.400 199.040 133.385 199.475 ;
        RECT 134.035 199.470 134.205 200.080 ;
        RECT 135.115 199.940 135.445 200.645 ;
        RECT 135.650 199.920 136.025 200.475 ;
        RECT 136.755 200.465 137.385 200.715 ;
        RECT 136.255 200.390 137.385 200.465 ;
        RECT 136.255 200.150 136.925 200.390 ;
        RECT 134.420 199.770 134.945 199.900 ;
        RECT 135.650 199.770 136.585 199.920 ;
        RECT 134.420 199.580 136.585 199.770 ;
        RECT 134.420 199.570 135.445 199.580 ;
        RECT 133.555 199.400 134.205 199.470 ;
        RECT 133.555 199.230 134.815 199.400 ;
        RECT 133.555 199.210 134.205 199.230 ;
        RECT 131.660 198.780 133.840 199.040 ;
        RECT 131.660 198.750 133.385 198.780 ;
        RECT 128.935 198.080 131.145 198.480 ;
        RECT 131.315 198.310 132.230 198.580 ;
        RECT 132.400 198.310 133.385 198.750 ;
        RECT 134.035 198.610 134.205 199.210 ;
        RECT 134.425 198.905 134.945 199.060 ;
        RECT 135.115 199.020 135.445 199.570 ;
        RECT 136.755 199.410 136.925 200.150 ;
        RECT 137.555 200.265 138.845 200.715 ;
        RECT 139.015 200.390 139.645 200.715 ;
        RECT 141.055 200.695 141.400 201.085 ;
        RECT 142.195 200.925 142.365 202.635 ;
        RECT 143.935 202.465 144.235 202.925 ;
        RECT 144.415 202.645 145.085 203.015 ;
        RECT 145.255 202.840 145.885 203.120 ;
        RECT 142.535 202.295 144.635 202.465 ;
        RECT 142.535 202.215 142.865 202.295 ;
        RECT 142.665 201.275 142.835 201.990 ;
        RECT 143.035 201.935 143.755 202.125 ;
        RECT 144.465 202.060 144.635 202.295 ;
        RECT 144.915 202.320 145.085 202.645 ;
        RECT 145.715 202.445 145.885 202.840 ;
        RECT 146.055 202.615 146.615 203.310 ;
        RECT 146.785 202.840 147.465 203.120 ;
        RECT 146.785 202.445 147.005 202.840 ;
        RECT 144.915 201.995 145.545 202.320 ;
        RECT 145.715 201.995 147.005 202.445 ;
        RECT 147.635 202.320 147.805 204.110 ;
        RECT 147.175 201.995 147.805 202.320 ;
        RECT 143.965 201.765 144.295 201.910 ;
        RECT 143.005 201.445 144.295 201.765 ;
        RECT 144.465 201.275 144.635 201.890 ;
        RECT 142.665 201.105 144.635 201.275 ;
        RECT 141.055 200.685 141.225 200.695 ;
        RECT 139.825 200.515 141.225 200.685 ;
        RECT 139.825 200.405 140.155 200.515 ;
        RECT 137.555 199.870 137.775 200.265 ;
        RECT 137.095 199.590 137.775 199.870 ;
        RECT 135.745 199.240 136.925 199.410 ;
        RECT 137.945 199.400 138.505 200.095 ;
        RECT 138.675 199.870 138.845 200.265 ;
        RECT 139.475 200.175 139.645 200.390 ;
        RECT 139.475 199.960 140.155 200.175 ;
        RECT 140.325 200.080 140.885 200.345 ;
        RECT 138.675 199.590 139.305 199.870 ;
        RECT 134.425 198.850 134.985 198.905 ;
        RECT 135.615 198.895 136.540 199.070 ;
        RECT 135.565 198.850 136.540 198.895 ;
        RECT 134.425 198.740 136.540 198.850 ;
        RECT 134.425 198.730 135.695 198.740 ;
        RECT 134.860 198.680 135.695 198.730 ;
        RECT 133.555 198.310 134.205 198.610 ;
        RECT 129.395 197.700 130.685 197.910 ;
        RECT 126.675 197.240 127.965 197.450 ;
        RECT 122.205 196.245 122.535 196.390 ;
        RECT 121.245 195.925 122.535 196.245 ;
        RECT 122.705 195.755 122.875 196.370 ;
        RECT 120.905 195.585 122.875 195.755 ;
        RECT 123.155 196.320 123.820 196.720 ;
        RECT 124.185 196.690 124.715 197.080 ;
        RECT 123.155 195.730 123.325 196.320 ;
        RECT 124.185 196.260 124.565 196.690 ;
        RECT 124.885 196.395 125.195 197.090 ;
        RECT 125.875 197.085 126.505 197.220 ;
        RECT 125.405 196.950 126.505 197.085 ;
        RECT 125.405 196.400 126.045 196.950 ;
        RECT 126.675 196.780 126.895 197.240 ;
        RECT 126.215 196.495 126.895 196.780 ;
        RECT 123.495 196.090 124.015 196.150 ;
        RECT 124.820 196.090 125.605 196.220 ;
        RECT 123.495 195.915 125.605 196.090 ;
        RECT 125.875 196.210 126.045 196.400 ;
        RECT 127.065 196.380 127.625 197.070 ;
        RECT 127.795 196.780 127.965 197.240 ;
        RECT 128.595 197.410 129.225 197.680 ;
        RECT 128.595 197.220 128.765 197.410 ;
        RECT 129.395 197.240 129.565 197.700 ;
        RECT 128.135 196.950 128.765 197.220 ;
        RECT 128.935 196.955 129.565 197.240 ;
        RECT 127.795 196.495 128.425 196.780 ;
        RECT 128.595 196.670 128.765 196.950 ;
        RECT 129.735 196.840 130.295 197.530 ;
        RECT 130.465 197.240 130.685 197.700 ;
        RECT 131.315 197.680 131.485 198.310 ;
        RECT 134.035 198.050 134.205 198.310 ;
        RECT 136.755 198.600 136.925 199.240 ;
        RECT 137.095 199.000 139.305 199.400 ;
        RECT 139.475 198.910 139.645 199.960 ;
        RECT 141.055 199.830 141.225 200.515 ;
        RECT 142.195 200.610 142.865 200.925 ;
        RECT 142.195 200.210 142.365 200.610 ;
        RECT 143.095 200.380 143.470 200.935 ;
        RECT 143.675 200.400 144.005 201.105 ;
        RECT 144.915 200.830 145.085 201.995 ;
        RECT 145.995 201.890 146.325 201.995 ;
        RECT 145.255 201.720 145.825 201.825 ;
        RECT 146.495 201.720 147.465 201.825 ;
        RECT 145.255 201.440 147.465 201.720 ;
        RECT 144.385 200.620 145.085 200.830 ;
        RECT 141.395 199.880 142.365 200.210 ;
        RECT 142.535 200.230 143.470 200.380 ;
        RECT 144.175 200.230 144.700 200.360 ;
        RECT 142.535 200.040 144.700 200.230 ;
        RECT 139.815 199.490 140.385 199.790 ;
        RECT 140.555 199.660 141.225 199.830 ;
        RECT 142.195 199.870 142.365 199.880 ;
        RECT 143.675 200.030 144.700 200.040 ;
        RECT 144.915 200.345 145.085 200.620 ;
        RECT 147.635 200.345 147.805 201.995 ;
        RECT 144.915 200.085 145.925 200.345 ;
        RECT 146.485 200.085 147.805 200.345 ;
        RECT 141.405 199.490 142.025 199.710 ;
        RECT 139.815 199.175 142.025 199.490 ;
        RECT 142.195 199.700 143.375 199.870 ;
        RECT 142.195 198.910 142.365 199.700 ;
        RECT 142.580 199.355 143.505 199.530 ;
        RECT 143.675 199.480 144.005 200.030 ;
        RECT 144.915 199.860 145.085 200.085 ;
        RECT 144.305 199.690 145.085 199.860 ;
        RECT 144.175 199.365 144.695 199.520 ;
        RECT 142.580 199.310 143.555 199.355 ;
        RECT 144.135 199.310 144.695 199.365 ;
        RECT 142.580 199.200 144.695 199.310 ;
        RECT 143.425 199.190 144.695 199.200 ;
        RECT 144.915 199.485 145.085 199.690 ;
        RECT 145.255 199.740 147.465 199.910 ;
        RECT 145.255 199.655 145.830 199.740 ;
        RECT 146.560 199.655 147.465 199.740 ;
        RECT 145.995 199.485 146.325 199.570 ;
        RECT 147.635 199.485 147.805 200.085 ;
        RECT 143.425 199.140 144.260 199.190 ;
        RECT 144.915 199.155 145.465 199.485 ;
        RECT 145.635 199.315 146.705 199.485 ;
        RECT 137.555 198.620 138.845 198.830 ;
        RECT 136.755 198.330 137.385 198.600 ;
        RECT 136.755 198.050 136.925 198.330 ;
        RECT 137.555 198.160 137.775 198.620 ;
        RECT 130.855 197.495 131.485 197.680 ;
        RECT 131.655 197.770 133.865 198.050 ;
        RECT 131.655 197.665 132.625 197.770 ;
        RECT 133.295 197.665 133.865 197.770 ;
        RECT 134.035 197.780 134.840 198.050 ;
        RECT 135.800 197.780 136.925 198.050 ;
        RECT 137.095 197.875 137.775 198.160 ;
        RECT 132.795 197.495 133.125 197.600 ;
        RECT 134.035 197.495 134.205 197.780 ;
        RECT 130.855 197.410 131.945 197.495 ;
        RECT 130.465 196.955 131.145 197.240 ;
        RECT 131.315 197.170 131.945 197.410 ;
        RECT 131.315 196.670 131.485 197.170 ;
        RECT 128.595 196.210 130.055 196.670 ;
        RECT 125.875 195.730 127.135 196.210 ;
        RECT 117.180 195.280 117.885 195.460 ;
        RECT 116.735 194.880 117.510 195.060 ;
        RECT 115.515 194.815 117.510 194.880 ;
        RECT 117.715 194.850 117.885 195.280 ;
        RECT 120.435 195.405 120.605 195.460 ;
        RECT 118.055 195.030 118.605 195.200 ;
        RECT 115.515 194.540 116.905 194.815 ;
        RECT 117.715 194.520 118.265 194.850 ;
        RECT 118.435 194.705 118.605 195.030 ;
        RECT 118.785 194.940 119.155 195.270 ;
        RECT 119.335 195.030 120.265 195.200 ;
        RECT 120.435 195.090 121.105 195.405 ;
        RECT 119.335 194.705 119.505 195.030 ;
        RECT 120.435 194.850 120.605 195.090 ;
        RECT 121.335 194.860 121.710 195.415 ;
        RECT 121.915 194.880 122.245 195.585 ;
        RECT 123.155 195.460 123.960 195.730 ;
        RECT 124.920 195.460 127.135 195.730 ;
        RECT 123.155 195.310 123.325 195.460 ;
        RECT 122.625 195.290 123.325 195.310 ;
        RECT 125.875 195.290 127.135 195.460 ;
        RECT 122.625 195.100 124.615 195.290 ;
        RECT 118.435 194.535 119.505 194.705 ;
        RECT 117.715 193.470 117.885 194.520 ;
        RECT 118.860 194.420 119.190 194.535 ;
        RECT 119.675 194.520 120.605 194.850 ;
        RECT 120.775 194.710 121.710 194.860 ;
        RECT 122.415 194.710 122.940 194.840 ;
        RECT 120.775 194.520 122.940 194.710 ;
        RECT 120.435 194.350 120.605 194.520 ;
        RECT 121.915 194.510 122.940 194.520 ;
        RECT 118.055 194.250 118.560 194.340 ;
        RECT 119.360 194.250 120.265 194.350 ;
        RECT 118.055 194.080 120.265 194.250 ;
        RECT 120.435 194.180 121.615 194.350 ;
        RECT 118.055 193.650 118.605 193.820 ;
        RECT 117.715 193.450 118.265 193.470 ;
        RECT 13.380 193.115 92.040 193.285 ;
        RECT 112.275 193.160 113.170 193.450 ;
        RECT 113.830 193.160 116.330 193.450 ;
        RECT 116.990 193.160 118.265 193.450 ;
        RECT 13.465 192.365 14.675 193.115 ;
        RECT 14.845 192.570 20.190 193.115 ;
        RECT 20.365 192.570 25.710 193.115 ;
        RECT 25.885 192.570 31.230 193.115 ;
        RECT 31.405 192.570 36.750 193.115 ;
        RECT 13.465 191.825 13.985 192.365 ;
        RECT 14.155 191.655 14.675 192.195 ;
        RECT 16.430 191.740 16.770 192.570 ;
        RECT 13.465 190.565 14.675 191.655 ;
        RECT 18.250 191.000 18.600 192.250 ;
        RECT 21.950 191.740 22.290 192.570 ;
        RECT 23.770 191.000 24.120 192.250 ;
        RECT 27.470 191.740 27.810 192.570 ;
        RECT 29.290 191.000 29.640 192.250 ;
        RECT 32.990 191.740 33.330 192.570 ;
        RECT 36.925 192.345 38.595 193.115 ;
        RECT 39.225 192.390 39.515 193.115 ;
        RECT 39.685 192.365 40.895 193.115 ;
        RECT 41.065 192.465 41.325 192.945 ;
        RECT 41.495 192.575 41.745 193.115 ;
        RECT 34.810 191.000 35.160 192.250 ;
        RECT 36.925 191.825 37.675 192.345 ;
        RECT 37.845 191.655 38.595 192.175 ;
        RECT 39.685 191.825 40.205 192.365 ;
        RECT 14.845 190.565 20.190 191.000 ;
        RECT 20.365 190.565 25.710 191.000 ;
        RECT 25.885 190.565 31.230 191.000 ;
        RECT 31.405 190.565 36.750 191.000 ;
        RECT 36.925 190.565 38.595 191.655 ;
        RECT 39.225 190.565 39.515 191.730 ;
        RECT 40.375 191.655 40.895 192.195 ;
        RECT 39.685 190.565 40.895 191.655 ;
        RECT 41.065 191.435 41.235 192.465 ;
        RECT 41.915 192.410 42.135 192.895 ;
        RECT 41.405 191.815 41.635 192.210 ;
        RECT 41.805 191.985 42.135 192.410 ;
        RECT 42.305 192.735 43.195 192.905 ;
        RECT 42.305 192.010 42.475 192.735 ;
        RECT 42.645 192.180 43.195 192.565 ;
        RECT 43.385 192.305 43.625 193.115 ;
        RECT 43.795 192.305 44.125 192.945 ;
        RECT 44.295 192.305 44.565 193.115 ;
        RECT 44.830 192.615 45.325 192.945 ;
        RECT 42.305 191.940 43.195 192.010 ;
        RECT 42.300 191.915 43.195 191.940 ;
        RECT 42.290 191.900 43.195 191.915 ;
        RECT 42.285 191.885 43.195 191.900 ;
        RECT 42.275 191.880 43.195 191.885 ;
        RECT 42.270 191.870 43.195 191.880 ;
        RECT 43.365 191.875 43.715 192.125 ;
        RECT 42.265 191.860 43.195 191.870 ;
        RECT 42.255 191.855 43.195 191.860 ;
        RECT 42.245 191.845 43.195 191.855 ;
        RECT 42.235 191.840 43.195 191.845 ;
        RECT 42.235 191.835 42.570 191.840 ;
        RECT 42.220 191.830 42.570 191.835 ;
        RECT 42.205 191.820 42.570 191.830 ;
        RECT 42.180 191.815 42.570 191.820 ;
        RECT 41.405 191.810 42.570 191.815 ;
        RECT 41.405 191.775 42.540 191.810 ;
        RECT 41.405 191.750 42.505 191.775 ;
        RECT 41.405 191.720 42.475 191.750 ;
        RECT 41.405 191.690 42.455 191.720 ;
        RECT 41.405 191.660 42.435 191.690 ;
        RECT 41.405 191.650 42.365 191.660 ;
        RECT 41.405 191.640 42.340 191.650 ;
        RECT 41.405 191.625 42.320 191.640 ;
        RECT 41.405 191.610 42.300 191.625 ;
        RECT 41.510 191.600 42.295 191.610 ;
        RECT 41.510 191.565 42.280 191.600 ;
        RECT 41.065 190.735 41.340 191.435 ;
        RECT 41.510 191.315 42.265 191.565 ;
        RECT 42.435 191.245 42.765 191.490 ;
        RECT 42.935 191.390 43.195 191.840 ;
        RECT 43.885 191.705 44.055 192.305 ;
        RECT 44.225 191.875 44.575 192.125 ;
        RECT 43.375 191.535 44.055 191.705 ;
        RECT 42.580 191.220 42.765 191.245 ;
        RECT 42.580 191.120 43.195 191.220 ;
        RECT 41.510 190.565 41.765 191.110 ;
        RECT 41.935 190.735 42.415 191.075 ;
        RECT 42.590 190.565 43.195 191.120 ;
        RECT 43.375 190.750 43.705 191.535 ;
        RECT 44.235 190.565 44.565 191.705 ;
        RECT 44.745 191.125 44.985 192.435 ;
        RECT 45.155 191.705 45.325 192.615 ;
        RECT 45.545 191.875 45.895 192.840 ;
        RECT 46.075 191.875 46.375 192.845 ;
        RECT 46.555 191.875 46.835 192.845 ;
        RECT 47.015 192.315 47.285 193.115 ;
        RECT 47.455 192.395 47.795 192.905 ;
        RECT 47.990 192.725 48.320 193.115 ;
        RECT 48.490 192.555 48.715 192.935 ;
        RECT 47.030 191.875 47.360 192.125 ;
        RECT 47.030 191.705 47.345 191.875 ;
        RECT 45.155 191.535 47.345 191.705 ;
        RECT 44.750 190.565 45.085 190.945 ;
        RECT 45.255 190.735 45.505 191.535 ;
        RECT 45.725 190.565 46.055 191.285 ;
        RECT 46.240 190.735 46.490 191.535 ;
        RECT 46.955 190.565 47.285 191.365 ;
        RECT 47.535 190.995 47.795 192.395 ;
        RECT 47.975 191.875 48.215 192.525 ;
        RECT 48.385 192.375 48.715 192.555 ;
        RECT 48.385 191.705 48.560 192.375 ;
        RECT 48.915 192.205 49.145 192.825 ;
        RECT 49.325 192.385 49.625 193.115 ;
        RECT 49.805 192.280 50.095 193.115 ;
        RECT 50.265 192.715 51.220 192.885 ;
        RECT 51.635 192.725 51.965 193.115 ;
        RECT 48.730 191.875 49.145 192.205 ;
        RECT 49.325 191.875 49.620 192.205 ;
        RECT 50.265 191.835 50.435 192.715 ;
        RECT 52.135 192.545 52.305 192.865 ;
        RECT 52.475 192.725 52.805 193.115 ;
        RECT 53.025 192.570 58.370 193.115 ;
        RECT 50.605 192.375 52.855 192.545 ;
        RECT 50.605 191.875 50.835 192.375 ;
        RECT 51.005 191.955 51.380 192.125 ;
        RECT 47.455 190.735 47.795 190.995 ;
        RECT 47.975 191.515 48.560 191.705 ;
        RECT 47.975 190.745 48.250 191.515 ;
        RECT 48.730 191.345 49.625 191.675 ;
        RECT 48.420 191.175 49.625 191.345 ;
        RECT 48.420 190.745 48.750 191.175 ;
        RECT 48.920 190.565 49.115 191.005 ;
        RECT 49.295 190.745 49.625 191.175 ;
        RECT 49.805 191.665 50.435 191.835 ;
        RECT 51.210 191.755 51.380 191.955 ;
        RECT 51.550 191.925 52.100 192.125 ;
        RECT 52.270 191.755 52.515 192.205 ;
        RECT 49.805 190.735 50.125 191.665 ;
        RECT 51.210 191.585 52.515 191.755 ;
        RECT 52.685 191.415 52.855 192.375 ;
        RECT 54.610 191.740 54.950 192.570 ;
        RECT 58.545 192.345 62.055 193.115 ;
        RECT 62.285 192.635 62.565 193.115 ;
        RECT 62.735 192.465 62.995 192.855 ;
        RECT 63.170 192.635 63.425 193.115 ;
        RECT 63.595 192.465 63.890 192.855 ;
        RECT 64.070 192.635 64.345 193.115 ;
        RECT 64.515 192.615 64.815 192.945 ;
        RECT 50.305 191.245 51.545 191.415 ;
        RECT 50.305 190.735 50.705 191.245 ;
        RECT 50.875 190.565 51.045 191.075 ;
        RECT 51.215 190.735 51.545 191.245 ;
        RECT 51.715 190.565 51.885 191.415 ;
        RECT 52.475 190.735 52.855 191.415 ;
        RECT 56.430 191.000 56.780 192.250 ;
        RECT 58.545 191.825 60.195 192.345 ;
        RECT 62.240 192.295 63.890 192.465 ;
        RECT 60.365 191.655 62.055 192.175 ;
        RECT 53.025 190.565 58.370 191.000 ;
        RECT 58.545 190.565 62.055 191.655 ;
        RECT 62.240 191.785 62.645 192.295 ;
        RECT 62.815 191.955 63.955 192.125 ;
        RECT 62.240 191.615 62.995 191.785 ;
        RECT 62.280 190.565 62.565 191.435 ;
        RECT 62.735 191.365 62.995 191.615 ;
        RECT 63.785 191.705 63.955 191.955 ;
        RECT 64.125 191.875 64.475 192.445 ;
        RECT 64.645 191.705 64.815 192.615 ;
        RECT 64.985 192.390 65.275 193.115 ;
        RECT 65.530 192.615 66.025 192.945 ;
        RECT 63.785 191.535 64.815 191.705 ;
        RECT 62.735 191.195 63.855 191.365 ;
        RECT 62.735 190.735 62.995 191.195 ;
        RECT 63.170 190.565 63.425 191.025 ;
        RECT 63.595 190.735 63.855 191.195 ;
        RECT 64.025 190.565 64.335 191.365 ;
        RECT 64.505 190.735 64.815 191.535 ;
        RECT 64.985 190.565 65.275 191.730 ;
        RECT 65.445 191.125 65.685 192.435 ;
        RECT 65.855 191.705 66.025 192.615 ;
        RECT 66.245 191.875 66.595 192.840 ;
        RECT 66.775 191.875 67.075 192.845 ;
        RECT 67.255 191.875 67.535 192.845 ;
        RECT 67.715 192.315 67.985 193.115 ;
        RECT 68.155 192.395 68.495 192.905 ;
        RECT 68.690 192.725 69.020 193.115 ;
        RECT 69.190 192.555 69.415 192.935 ;
        RECT 67.730 191.875 68.060 192.125 ;
        RECT 67.730 191.705 68.045 191.875 ;
        RECT 65.855 191.535 68.045 191.705 ;
        RECT 65.450 190.565 65.785 190.945 ;
        RECT 65.955 190.735 66.205 191.535 ;
        RECT 66.425 190.565 66.755 191.285 ;
        RECT 66.940 190.735 67.190 191.535 ;
        RECT 67.655 190.565 67.985 191.365 ;
        RECT 68.235 190.995 68.495 192.395 ;
        RECT 68.675 191.875 68.915 192.525 ;
        RECT 69.085 192.375 69.415 192.555 ;
        RECT 69.085 191.705 69.260 192.375 ;
        RECT 69.615 192.205 69.845 192.825 ;
        RECT 70.025 192.385 70.325 193.115 ;
        RECT 70.590 192.615 71.085 192.945 ;
        RECT 69.430 191.875 69.845 192.205 ;
        RECT 70.025 191.875 70.320 192.205 ;
        RECT 68.155 190.735 68.495 190.995 ;
        RECT 68.675 191.515 69.260 191.705 ;
        RECT 68.675 190.745 68.950 191.515 ;
        RECT 69.430 191.345 70.325 191.675 ;
        RECT 69.120 191.175 70.325 191.345 ;
        RECT 69.120 190.745 69.450 191.175 ;
        RECT 69.620 190.565 69.815 191.005 ;
        RECT 69.995 190.745 70.325 191.175 ;
        RECT 70.505 191.125 70.745 192.435 ;
        RECT 70.915 191.705 71.085 192.615 ;
        RECT 71.305 191.875 71.655 192.840 ;
        RECT 71.835 191.875 72.135 192.845 ;
        RECT 72.315 191.875 72.595 192.845 ;
        RECT 72.775 192.315 73.045 193.115 ;
        RECT 73.215 192.395 73.555 192.905 ;
        RECT 73.890 192.605 74.130 193.115 ;
        RECT 74.310 192.605 74.590 192.935 ;
        RECT 74.820 192.605 75.035 193.115 ;
        RECT 72.790 191.875 73.120 192.125 ;
        RECT 72.790 191.705 73.105 191.875 ;
        RECT 70.915 191.535 73.105 191.705 ;
        RECT 70.510 190.565 70.845 190.945 ;
        RECT 71.015 190.735 71.265 191.535 ;
        RECT 71.485 190.565 71.815 191.285 ;
        RECT 72.000 190.735 72.250 191.535 ;
        RECT 72.715 190.565 73.045 191.365 ;
        RECT 73.295 190.995 73.555 192.395 ;
        RECT 73.785 191.875 74.140 192.435 ;
        RECT 74.310 191.705 74.480 192.605 ;
        RECT 74.650 191.875 74.915 192.435 ;
        RECT 75.205 192.375 75.820 192.945 ;
        RECT 76.025 192.570 81.370 193.115 ;
        RECT 81.545 192.570 86.890 193.115 ;
        RECT 75.165 191.705 75.335 192.205 ;
        RECT 73.910 191.535 75.335 191.705 ;
        RECT 73.910 191.360 74.300 191.535 ;
        RECT 73.215 190.735 73.555 190.995 ;
        RECT 74.785 190.565 75.115 191.365 ;
        RECT 75.505 191.355 75.820 192.375 ;
        RECT 77.610 191.740 77.950 192.570 ;
        RECT 75.285 190.735 75.820 191.355 ;
        RECT 79.430 191.000 79.780 192.250 ;
        RECT 83.130 191.740 83.470 192.570 ;
        RECT 87.065 192.345 90.575 193.115 ;
        RECT 90.745 192.365 91.955 193.115 ;
        RECT 84.950 191.000 85.300 192.250 ;
        RECT 87.065 191.825 88.715 192.345 ;
        RECT 88.885 191.655 90.575 192.175 ;
        RECT 76.025 190.565 81.370 191.000 ;
        RECT 81.545 190.565 86.890 191.000 ;
        RECT 87.065 190.565 90.575 191.655 ;
        RECT 90.745 191.655 91.265 192.195 ;
        RECT 91.435 191.825 91.955 192.365 ;
        RECT 90.745 190.565 91.955 191.655 ;
        RECT 112.275 191.595 112.445 193.160 ;
        RECT 114.995 192.435 115.165 193.160 ;
        RECT 117.715 193.140 118.265 193.160 ;
        RECT 118.435 193.325 118.605 193.650 ;
        RECT 118.785 193.560 119.155 193.890 ;
        RECT 119.335 193.650 120.265 193.820 ;
        RECT 119.335 193.325 119.505 193.650 ;
        RECT 120.435 193.470 120.605 194.180 ;
        RECT 120.820 193.835 121.745 194.010 ;
        RECT 121.915 193.960 122.245 194.510 ;
        RECT 123.155 194.340 124.615 195.100 ;
        RECT 122.545 194.170 124.615 194.340 ;
        RECT 123.155 194.080 124.615 194.170 ;
        RECT 124.785 194.830 127.135 195.290 ;
        RECT 127.305 196.150 130.055 196.210 ;
        RECT 127.305 195.460 129.515 196.150 ;
        RECT 130.225 195.980 131.485 196.670 ;
        RECT 132.115 197.045 133.405 197.495 ;
        RECT 133.575 197.190 134.205 197.495 ;
        RECT 134.375 197.420 136.485 197.595 ;
        RECT 134.375 197.360 134.895 197.420 ;
        RECT 135.700 197.290 136.485 197.420 ;
        RECT 136.755 197.590 136.925 197.780 ;
        RECT 137.945 197.760 138.505 198.450 ;
        RECT 138.675 198.160 138.845 198.620 ;
        RECT 139.475 198.700 140.465 198.910 ;
        RECT 141.055 198.700 142.365 198.910 ;
        RECT 139.475 198.600 139.645 198.700 ;
        RECT 139.015 198.330 139.645 198.600 ;
        RECT 138.675 197.875 139.305 198.160 ;
        RECT 139.475 198.030 139.645 198.330 ;
        RECT 139.815 198.280 142.025 198.530 ;
        RECT 139.815 198.200 140.445 198.280 ;
        RECT 141.045 198.200 142.025 198.280 ;
        RECT 142.195 198.230 142.365 198.700 ;
        RECT 142.535 198.620 144.745 198.935 ;
        RECT 142.535 198.400 143.155 198.620 ;
        RECT 143.335 198.280 144.005 198.450 ;
        RECT 144.175 198.320 144.745 198.620 ;
        RECT 139.475 197.800 140.465 198.030 ;
        RECT 139.475 197.590 139.645 197.800 ;
        RECT 140.635 197.780 140.885 198.110 ;
        RECT 142.195 198.030 143.165 198.230 ;
        RECT 141.055 197.900 143.165 198.030 ;
        RECT 141.055 197.800 142.365 197.900 ;
        RECT 133.575 197.170 134.700 197.190 ;
        RECT 132.115 196.650 132.335 197.045 ;
        RECT 131.655 196.370 132.335 196.650 ;
        RECT 132.505 196.180 133.065 196.875 ;
        RECT 133.235 196.650 133.405 197.045 ;
        RECT 134.035 196.790 134.700 197.170 ;
        RECT 135.065 196.820 135.445 197.250 ;
        RECT 133.235 196.370 133.865 196.650 ;
        RECT 129.685 195.460 131.485 195.980 ;
        RECT 131.655 195.780 133.865 196.180 ;
        RECT 127.305 195.000 128.765 195.460 ;
        RECT 131.315 195.380 131.485 195.460 ;
        RECT 132.115 195.400 133.405 195.610 ;
        RECT 129.095 195.120 131.145 195.290 ;
        RECT 129.095 195.015 129.440 195.120 ;
        RECT 130.175 195.015 131.145 195.120 ;
        RECT 131.315 195.110 131.945 195.380 ;
        RECT 122.415 193.845 122.935 194.000 ;
        RECT 120.820 193.790 121.795 193.835 ;
        RECT 122.375 193.790 122.935 193.845 ;
        RECT 120.820 193.680 122.935 193.790 ;
        RECT 121.665 193.670 122.935 193.680 ;
        RECT 121.665 193.620 122.500 193.670 ;
        RECT 118.435 193.155 119.505 193.325 ;
        RECT 119.675 193.450 120.605 193.470 ;
        RECT 123.155 193.450 124.095 194.080 ;
        RECT 124.785 193.910 127.655 194.830 ;
        RECT 119.675 193.160 121.770 193.450 ;
        RECT 122.430 193.160 124.095 193.450 ;
        RECT 115.335 192.710 117.545 192.990 ;
        RECT 115.335 192.605 116.305 192.710 ;
        RECT 116.975 192.605 117.545 192.710 ;
        RECT 116.475 192.435 116.805 192.540 ;
        RECT 117.715 192.435 117.885 193.140 ;
        RECT 118.860 193.040 119.190 193.155 ;
        RECT 119.675 193.140 120.605 193.160 ;
        RECT 118.055 192.870 118.560 192.960 ;
        RECT 119.360 192.870 120.265 192.970 ;
        RECT 118.055 192.700 120.265 192.870 ;
        RECT 114.995 192.110 115.625 192.435 ;
        RECT 112.615 191.810 113.165 191.980 ;
        RECT 112.275 191.265 112.825 191.595 ;
        RECT 112.995 191.435 113.165 191.810 ;
        RECT 113.345 191.715 113.715 192.070 ;
        RECT 113.895 191.810 114.825 191.980 ;
        RECT 113.895 191.435 114.065 191.810 ;
        RECT 114.995 191.595 115.165 192.110 ;
        RECT 112.995 191.265 114.065 191.435 ;
        RECT 114.235 191.265 115.165 191.595 ;
        RECT 115.795 191.985 117.085 192.435 ;
        RECT 117.255 192.110 117.885 192.435 ;
        RECT 118.055 192.270 118.605 192.440 ;
        RECT 115.795 191.590 116.015 191.985 ;
        RECT 115.335 191.310 116.015 191.590 ;
        RECT 112.275 190.665 112.445 191.265 ;
        RECT 113.355 191.180 113.685 191.265 ;
        RECT 112.615 191.010 113.190 191.095 ;
        RECT 113.920 191.010 114.825 191.095 ;
        RECT 112.615 190.840 114.825 191.010 ;
        RECT 114.995 190.665 115.165 191.265 ;
        RECT 116.185 191.120 116.745 191.815 ;
        RECT 116.915 191.590 117.085 191.985 ;
        RECT 117.715 192.090 117.885 192.110 ;
        RECT 117.715 191.760 118.265 192.090 ;
        RECT 118.435 191.945 118.605 192.270 ;
        RECT 118.785 192.180 119.155 192.510 ;
        RECT 120.435 192.480 120.605 193.140 ;
        RECT 120.775 192.815 122.985 192.985 ;
        RECT 120.775 192.650 121.745 192.815 ;
        RECT 122.415 192.730 122.985 192.815 ;
        RECT 123.155 192.700 124.095 193.160 ;
        RECT 124.265 193.620 127.655 193.910 ;
        RECT 127.825 194.825 128.765 195.000 ;
        RECT 129.675 194.845 130.005 194.950 ;
        RECT 127.825 194.445 129.165 194.825 ;
        RECT 129.335 194.675 130.345 194.845 ;
        RECT 131.315 194.805 131.485 195.110 ;
        RECT 132.115 194.940 132.335 195.400 ;
        RECT 127.825 193.935 128.765 194.445 ;
        RECT 129.335 194.275 129.505 194.675 ;
        RECT 128.985 194.105 129.505 194.275 ;
        RECT 129.675 194.125 130.005 194.505 ;
        RECT 130.175 194.355 130.345 194.675 ;
        RECT 130.515 194.525 131.485 194.805 ;
        RECT 131.655 194.655 132.335 194.940 ;
        RECT 132.505 194.540 133.065 195.230 ;
        RECT 133.235 194.940 133.405 195.400 ;
        RECT 134.035 195.380 134.205 196.790 ;
        RECT 135.065 196.430 135.595 196.820 ;
        RECT 134.535 196.260 135.595 196.430 ;
        RECT 135.765 196.420 136.075 197.115 ;
        RECT 136.755 197.110 138.015 197.590 ;
        RECT 136.285 196.900 138.015 197.110 ;
        RECT 138.185 197.160 139.645 197.590 ;
        RECT 139.905 197.330 140.365 197.500 ;
        RECT 138.185 197.070 140.025 197.160 ;
        RECT 136.285 196.425 138.555 196.900 ;
        RECT 134.535 196.200 134.730 196.260 ;
        RECT 134.390 196.030 134.730 196.200 ;
        RECT 135.425 196.245 135.595 196.260 ;
        RECT 136.755 196.380 138.555 196.425 ;
        RECT 138.725 196.830 140.025 197.070 ;
        RECT 140.195 197.065 140.365 197.330 ;
        RECT 140.535 197.235 141.185 197.585 ;
        RECT 141.355 197.330 142.025 197.500 ;
        RECT 141.355 197.065 141.525 197.330 ;
        RECT 142.195 197.160 142.365 197.800 ;
        RECT 143.335 197.595 143.505 198.280 ;
        RECT 144.915 198.150 145.085 199.155 ;
        RECT 145.635 198.940 145.805 199.315 ;
        RECT 145.255 198.770 145.805 198.940 ;
        RECT 145.985 198.680 146.355 199.035 ;
        RECT 146.535 198.940 146.705 199.315 ;
        RECT 146.875 199.155 147.805 199.485 ;
        RECT 146.535 198.770 147.465 198.940 ;
        RECT 143.675 197.765 144.235 198.030 ;
        RECT 144.405 197.940 145.085 198.150 ;
        RECT 145.255 198.110 145.885 198.395 ;
        RECT 144.405 197.935 145.545 197.940 ;
        RECT 144.405 197.595 144.735 197.705 ;
        RECT 143.335 197.425 144.735 197.595 ;
        RECT 144.915 197.670 145.545 197.935 ;
        RECT 143.335 197.415 143.505 197.425 ;
        RECT 140.195 196.835 141.525 197.065 ;
        RECT 141.695 196.830 142.365 197.160 ;
        RECT 143.160 197.025 143.505 197.415 ;
        RECT 143.675 196.900 144.235 197.255 ;
        RECT 144.915 197.245 145.085 197.670 ;
        RECT 145.715 197.650 145.885 198.110 ;
        RECT 146.055 197.820 146.615 198.510 ;
        RECT 146.785 198.110 147.465 198.395 ;
        RECT 146.785 197.650 147.005 198.110 ;
        RECT 147.635 197.940 147.805 199.155 ;
        RECT 147.175 197.670 147.805 197.940 ;
        RECT 145.715 197.440 147.005 197.650 ;
        RECT 144.405 197.005 145.085 197.245 ;
        RECT 138.725 196.380 139.645 196.830 ;
        RECT 139.905 196.475 142.025 196.660 ;
        RECT 134.925 195.770 135.255 196.090 ;
        RECT 135.425 195.960 136.540 196.245 ;
        RECT 134.925 195.750 136.135 195.770 ;
        RECT 136.755 195.760 136.925 196.380 ;
        RECT 139.475 196.220 139.645 196.380 ;
        RECT 134.400 195.535 136.135 195.750 ;
        RECT 134.400 195.510 134.775 195.535 ;
        RECT 133.575 195.340 134.205 195.380 ;
        RECT 133.575 195.110 134.710 195.340 ;
        RECT 134.035 195.010 134.710 195.110 ;
        RECT 134.885 195.065 135.735 195.365 ;
        RECT 135.905 195.260 136.135 195.535 ;
        RECT 136.305 195.430 136.925 195.760 ;
        RECT 135.905 195.090 136.565 195.260 ;
        RECT 134.885 195.060 135.055 195.065 ;
        RECT 133.235 194.655 133.865 194.940 ;
        RECT 130.175 194.185 130.635 194.355 ;
        RECT 127.825 193.620 129.165 193.935 ;
        RECT 124.265 193.450 126.045 193.620 ;
        RECT 128.595 193.605 129.165 193.620 ;
        RECT 128.595 193.450 128.765 193.605 ;
        RECT 124.265 193.160 127.210 193.450 ;
        RECT 127.870 193.160 128.765 193.450 ;
        RECT 129.335 193.430 129.505 194.105 ;
        RECT 128.985 193.260 129.505 193.430 ;
        RECT 129.675 193.215 130.295 193.955 ;
        RECT 124.265 192.700 126.045 193.160 ;
        RECT 128.595 193.060 128.765 193.160 ;
        RECT 121.915 192.560 122.245 192.645 ;
        RECT 123.155 192.560 123.325 192.700 ;
        RECT 119.335 192.270 120.265 192.440 ;
        RECT 120.435 192.310 121.745 192.480 ;
        RECT 121.915 192.390 122.585 192.560 ;
        RECT 119.335 191.945 119.505 192.270 ;
        RECT 120.435 192.090 120.605 192.310 ;
        RECT 121.915 192.140 122.245 192.165 ;
        RECT 118.435 191.775 119.505 191.945 ;
        RECT 116.915 191.310 117.545 191.590 ;
        RECT 115.335 190.720 117.545 191.120 ;
        RECT 13.380 190.395 92.040 190.565 ;
        RECT 112.275 190.405 113.285 190.665 ;
        RECT 113.845 190.405 115.165 190.665 ;
        RECT 117.715 190.710 117.885 191.760 ;
        RECT 118.860 191.660 119.190 191.775 ;
        RECT 119.675 191.760 120.605 192.090 ;
        RECT 118.055 191.490 118.560 191.580 ;
        RECT 119.360 191.490 120.265 191.590 ;
        RECT 118.055 191.320 120.265 191.490 ;
        RECT 118.055 190.890 118.605 191.060 ;
        RECT 13.465 189.305 14.675 190.395 ;
        RECT 14.845 189.960 20.190 190.395 ;
        RECT 20.365 189.960 25.710 190.395 ;
        RECT 13.465 188.595 13.985 189.135 ;
        RECT 14.155 188.765 14.675 189.305 ;
        RECT 13.465 187.845 14.675 188.595 ;
        RECT 16.430 188.390 16.770 189.220 ;
        RECT 18.250 188.710 18.600 189.960 ;
        RECT 21.950 188.390 22.290 189.220 ;
        RECT 23.770 188.710 24.120 189.960 ;
        RECT 26.345 189.230 26.635 190.395 ;
        RECT 26.805 189.960 32.150 190.395 ;
        RECT 32.325 189.960 37.670 190.395 ;
        RECT 14.845 187.845 20.190 188.390 ;
        RECT 20.365 187.845 25.710 188.390 ;
        RECT 26.345 187.845 26.635 188.570 ;
        RECT 28.390 188.390 28.730 189.220 ;
        RECT 30.210 188.710 30.560 189.960 ;
        RECT 33.910 188.390 34.250 189.220 ;
        RECT 35.730 188.710 36.080 189.960 ;
        RECT 37.845 189.305 41.355 190.395 ;
        RECT 37.845 188.615 39.495 189.135 ;
        RECT 39.665 188.785 41.355 189.305 ;
        RECT 41.525 189.525 41.800 190.225 ;
        RECT 41.970 189.850 42.225 190.395 ;
        RECT 42.395 189.885 42.875 190.225 ;
        RECT 43.050 189.840 43.655 190.395 ;
        RECT 43.825 189.960 49.170 190.395 ;
        RECT 43.040 189.740 43.655 189.840 ;
        RECT 43.040 189.715 43.225 189.740 ;
        RECT 26.805 187.845 32.150 188.390 ;
        RECT 32.325 187.845 37.670 188.390 ;
        RECT 37.845 187.845 41.355 188.615 ;
        RECT 41.525 188.495 41.695 189.525 ;
        RECT 41.970 189.395 42.725 189.645 ;
        RECT 42.895 189.470 43.225 189.715 ;
        RECT 41.970 189.360 42.740 189.395 ;
        RECT 41.970 189.350 42.755 189.360 ;
        RECT 41.865 189.335 42.760 189.350 ;
        RECT 41.865 189.320 42.780 189.335 ;
        RECT 41.865 189.310 42.800 189.320 ;
        RECT 41.865 189.300 42.825 189.310 ;
        RECT 41.865 189.270 42.895 189.300 ;
        RECT 41.865 189.240 42.915 189.270 ;
        RECT 41.865 189.210 42.935 189.240 ;
        RECT 41.865 189.185 42.965 189.210 ;
        RECT 41.865 189.150 43.000 189.185 ;
        RECT 41.865 189.145 43.030 189.150 ;
        RECT 41.865 188.750 42.095 189.145 ;
        RECT 42.640 189.140 43.030 189.145 ;
        RECT 42.665 189.130 43.030 189.140 ;
        RECT 42.680 189.125 43.030 189.130 ;
        RECT 42.695 189.120 43.030 189.125 ;
        RECT 43.395 189.120 43.655 189.570 ;
        RECT 42.695 189.115 43.655 189.120 ;
        RECT 42.705 189.105 43.655 189.115 ;
        RECT 42.715 189.100 43.655 189.105 ;
        RECT 42.725 189.090 43.655 189.100 ;
        RECT 42.730 189.080 43.655 189.090 ;
        RECT 42.735 189.075 43.655 189.080 ;
        RECT 42.745 189.060 43.655 189.075 ;
        RECT 42.750 189.045 43.655 189.060 ;
        RECT 42.760 189.020 43.655 189.045 ;
        RECT 42.265 188.550 42.595 188.975 ;
        RECT 41.525 188.015 41.785 188.495 ;
        RECT 41.955 187.845 42.205 188.385 ;
        RECT 42.375 188.065 42.595 188.550 ;
        RECT 42.765 188.950 43.655 189.020 ;
        RECT 42.765 188.225 42.935 188.950 ;
        RECT 43.105 188.395 43.655 188.780 ;
        RECT 45.410 188.390 45.750 189.220 ;
        RECT 47.230 188.710 47.580 189.960 ;
        RECT 49.345 189.305 51.935 190.395 ;
        RECT 49.345 188.615 50.555 189.135 ;
        RECT 50.725 188.785 51.935 189.305 ;
        RECT 52.105 189.230 52.395 190.395 ;
        RECT 52.565 189.305 56.075 190.395 ;
        RECT 52.565 188.615 54.215 189.135 ;
        RECT 54.385 188.785 56.075 189.305 ;
        RECT 57.175 189.785 57.505 190.215 ;
        RECT 57.685 189.955 57.880 190.395 ;
        RECT 58.050 189.785 58.380 190.215 ;
        RECT 57.175 189.615 58.380 189.785 ;
        RECT 57.175 189.285 58.070 189.615 ;
        RECT 58.550 189.445 58.825 190.215 ;
        RECT 58.240 189.255 58.825 189.445 ;
        RECT 57.180 188.755 57.475 189.085 ;
        RECT 57.655 188.755 58.070 189.085 ;
        RECT 42.765 188.055 43.655 188.225 ;
        RECT 43.825 187.845 49.170 188.390 ;
        RECT 49.345 187.845 51.935 188.615 ;
        RECT 52.105 187.845 52.395 188.570 ;
        RECT 52.565 187.845 56.075 188.615 ;
        RECT 57.175 187.845 57.475 188.575 ;
        RECT 57.655 188.135 57.885 188.755 ;
        RECT 58.240 188.585 58.415 189.255 ;
        RECT 58.085 188.405 58.415 188.585 ;
        RECT 58.585 188.435 58.825 189.085 ;
        RECT 58.085 188.025 58.310 188.405 ;
        RECT 58.480 187.845 58.810 188.235 ;
        RECT 59.005 188.125 59.285 190.225 ;
        RECT 59.475 189.635 60.260 190.395 ;
        RECT 60.655 189.565 61.040 190.225 ;
        RECT 60.655 189.465 61.065 189.565 ;
        RECT 59.455 189.255 61.065 189.465 ;
        RECT 61.365 189.375 61.565 190.165 ;
        RECT 59.455 188.655 59.730 189.255 ;
        RECT 61.235 189.205 61.565 189.375 ;
        RECT 61.735 189.215 62.055 190.395 ;
        RECT 61.235 189.085 61.415 189.205 ;
        RECT 59.900 188.835 60.255 189.085 ;
        RECT 60.450 189.035 60.915 189.085 ;
        RECT 60.445 188.865 60.915 189.035 ;
        RECT 60.450 188.835 60.915 188.865 ;
        RECT 61.085 188.835 61.415 189.085 ;
        RECT 61.590 188.835 62.055 189.035 ;
        RECT 62.225 188.790 62.505 190.225 ;
        RECT 62.675 189.620 63.385 190.395 ;
        RECT 63.555 189.450 63.885 190.225 ;
        RECT 62.735 189.235 63.885 189.450 ;
        RECT 59.455 188.475 60.705 188.655 ;
        RECT 60.340 188.405 60.705 188.475 ;
        RECT 60.875 188.455 62.055 188.625 ;
        RECT 59.515 187.845 59.685 188.305 ;
        RECT 60.875 188.235 61.205 188.455 ;
        RECT 59.955 188.055 61.205 188.235 ;
        RECT 61.375 187.845 61.545 188.285 ;
        RECT 61.715 188.040 62.055 188.455 ;
        RECT 62.225 188.015 62.565 188.790 ;
        RECT 62.735 188.665 63.020 189.235 ;
        RECT 63.205 188.835 63.675 189.065 ;
        RECT 64.080 189.035 64.295 190.150 ;
        RECT 64.475 189.675 64.805 190.395 ;
        RECT 65.445 189.525 65.720 190.225 ;
        RECT 65.890 189.850 66.145 190.395 ;
        RECT 66.315 189.885 66.795 190.225 ;
        RECT 66.970 189.840 67.575 190.395 ;
        RECT 66.960 189.740 67.575 189.840 ;
        RECT 66.960 189.715 67.145 189.740 ;
        RECT 64.585 189.035 64.815 189.375 ;
        RECT 63.845 188.855 64.295 189.035 ;
        RECT 63.845 188.835 64.175 188.855 ;
        RECT 64.485 188.835 64.815 189.035 ;
        RECT 62.735 188.475 63.445 188.665 ;
        RECT 63.145 188.335 63.445 188.475 ;
        RECT 63.635 188.475 64.815 188.665 ;
        RECT 63.635 188.395 63.965 188.475 ;
        RECT 63.145 188.325 63.460 188.335 ;
        RECT 63.145 188.315 63.470 188.325 ;
        RECT 63.145 188.310 63.480 188.315 ;
        RECT 62.735 187.845 62.905 188.305 ;
        RECT 63.145 188.300 63.485 188.310 ;
        RECT 63.145 188.295 63.490 188.300 ;
        RECT 63.145 188.285 63.495 188.295 ;
        RECT 63.145 188.280 63.500 188.285 ;
        RECT 63.145 188.015 63.505 188.280 ;
        RECT 64.135 187.845 64.305 188.305 ;
        RECT 64.475 188.015 64.815 188.475 ;
        RECT 65.445 188.495 65.615 189.525 ;
        RECT 65.890 189.395 66.645 189.645 ;
        RECT 66.815 189.470 67.145 189.715 ;
        RECT 65.890 189.360 66.660 189.395 ;
        RECT 65.890 189.350 66.675 189.360 ;
        RECT 65.785 189.335 66.680 189.350 ;
        RECT 65.785 189.320 66.700 189.335 ;
        RECT 65.785 189.310 66.720 189.320 ;
        RECT 65.785 189.300 66.745 189.310 ;
        RECT 65.785 189.270 66.815 189.300 ;
        RECT 65.785 189.240 66.835 189.270 ;
        RECT 65.785 189.210 66.855 189.240 ;
        RECT 65.785 189.185 66.885 189.210 ;
        RECT 65.785 189.150 66.920 189.185 ;
        RECT 65.785 189.145 66.950 189.150 ;
        RECT 65.785 188.750 66.015 189.145 ;
        RECT 66.560 189.140 66.950 189.145 ;
        RECT 66.585 189.130 66.950 189.140 ;
        RECT 66.600 189.125 66.950 189.130 ;
        RECT 66.615 189.120 66.950 189.125 ;
        RECT 67.315 189.120 67.575 189.570 ;
        RECT 67.745 189.305 70.335 190.395 ;
        RECT 66.615 189.115 67.575 189.120 ;
        RECT 66.625 189.105 67.575 189.115 ;
        RECT 66.635 189.100 67.575 189.105 ;
        RECT 66.645 189.090 67.575 189.100 ;
        RECT 66.650 189.080 67.575 189.090 ;
        RECT 66.655 189.075 67.575 189.080 ;
        RECT 66.665 189.060 67.575 189.075 ;
        RECT 66.670 189.045 67.575 189.060 ;
        RECT 66.680 189.020 67.575 189.045 ;
        RECT 66.185 188.550 66.515 188.975 ;
        RECT 65.445 188.015 65.705 188.495 ;
        RECT 65.875 187.845 66.125 188.385 ;
        RECT 66.295 188.065 66.515 188.550 ;
        RECT 66.685 188.950 67.575 189.020 ;
        RECT 66.685 188.225 66.855 188.950 ;
        RECT 67.025 188.395 67.575 188.780 ;
        RECT 67.745 188.615 68.955 189.135 ;
        RECT 69.125 188.785 70.335 189.305 ;
        RECT 70.965 189.255 71.245 190.395 ;
        RECT 71.415 189.245 71.745 190.225 ;
        RECT 71.915 189.255 72.175 190.395 ;
        RECT 72.345 189.960 77.690 190.395 ;
        RECT 70.975 188.815 71.310 189.085 ;
        RECT 71.480 188.645 71.650 189.245 ;
        RECT 71.820 188.835 72.155 189.085 ;
        RECT 66.685 188.055 67.575 188.225 ;
        RECT 67.745 187.845 70.335 188.615 ;
        RECT 70.965 187.845 71.275 188.645 ;
        RECT 71.480 188.015 72.175 188.645 ;
        RECT 73.930 188.390 74.270 189.220 ;
        RECT 75.750 188.710 76.100 189.960 ;
        RECT 77.865 189.230 78.155 190.395 ;
        RECT 78.325 189.960 83.670 190.395 ;
        RECT 83.845 189.960 89.190 190.395 ;
        RECT 72.345 187.845 77.690 188.390 ;
        RECT 77.865 187.845 78.155 188.570 ;
        RECT 79.910 188.390 80.250 189.220 ;
        RECT 81.730 188.710 82.080 189.960 ;
        RECT 85.430 188.390 85.770 189.220 ;
        RECT 87.250 188.710 87.600 189.960 ;
        RECT 89.365 189.305 90.575 190.395 ;
        RECT 89.365 188.595 89.885 189.135 ;
        RECT 90.055 188.765 90.575 189.305 ;
        RECT 90.745 189.305 91.955 190.395 ;
        RECT 112.275 189.790 112.445 190.405 ;
        RECT 114.995 190.320 115.165 190.405 ;
        RECT 115.795 190.340 117.085 190.550 ;
        RECT 112.615 190.050 114.825 190.230 ;
        RECT 112.615 189.970 113.120 190.050 ;
        RECT 113.920 189.960 114.825 190.050 ;
        RECT 114.995 190.050 115.625 190.320 ;
        RECT 112.275 189.460 112.825 189.790 ;
        RECT 113.420 189.775 113.750 189.880 ;
        RECT 114.995 189.790 115.165 190.050 ;
        RECT 115.795 189.880 116.015 190.340 ;
        RECT 112.995 189.605 114.065 189.775 ;
        RECT 90.745 188.765 91.265 189.305 ;
        RECT 91.435 188.595 91.955 189.135 ;
        RECT 78.325 187.845 83.670 188.390 ;
        RECT 83.845 187.845 89.190 188.390 ;
        RECT 89.365 187.845 90.575 188.595 ;
        RECT 90.745 187.845 91.955 188.595 ;
        RECT 112.275 187.925 112.445 189.460 ;
        RECT 112.995 189.280 113.165 189.605 ;
        RECT 112.615 189.110 113.165 189.280 ;
        RECT 113.345 189.040 113.715 189.380 ;
        RECT 113.895 189.280 114.065 189.605 ;
        RECT 114.235 189.460 115.165 189.790 ;
        RECT 115.335 189.595 116.015 189.880 ;
        RECT 116.185 189.480 116.745 190.170 ;
        RECT 116.915 189.880 117.085 190.340 ;
        RECT 117.715 190.380 118.265 190.710 ;
        RECT 118.435 190.565 118.605 190.890 ;
        RECT 118.785 190.800 119.155 191.130 ;
        RECT 119.335 190.890 120.265 191.060 ;
        RECT 119.335 190.565 119.505 190.890 ;
        RECT 120.435 190.710 120.605 191.760 ;
        RECT 118.435 190.395 119.505 190.565 ;
        RECT 117.715 190.320 117.885 190.380 ;
        RECT 117.255 190.050 117.885 190.320 ;
        RECT 118.860 190.280 119.190 190.395 ;
        RECT 119.675 190.380 120.605 190.710 ;
        RECT 116.915 189.595 117.545 189.880 ;
        RECT 117.715 189.760 117.885 190.050 ;
        RECT 118.055 190.110 118.560 190.200 ;
        RECT 119.360 190.110 120.265 190.210 ;
        RECT 118.055 189.940 120.265 190.110 ;
        RECT 120.435 189.940 120.605 190.380 ;
        RECT 120.775 191.970 122.245 192.140 ;
        RECT 120.775 190.280 120.945 191.970 ;
        RECT 122.415 191.805 122.585 192.390 ;
        RECT 122.755 192.230 123.325 192.560 ;
        RECT 122.415 191.800 122.985 191.805 ;
        RECT 121.115 191.630 122.985 191.800 ;
        RECT 121.115 190.675 121.285 191.630 ;
        RECT 121.455 191.290 122.425 191.460 ;
        RECT 121.455 190.640 121.625 191.290 ;
        RECT 122.620 191.275 122.985 191.630 ;
        RECT 123.155 191.500 123.325 192.230 ;
        RECT 123.495 191.670 124.125 191.955 ;
        RECT 123.155 191.230 123.785 191.500 ;
        RECT 122.645 191.085 122.815 191.090 ;
        RECT 121.825 190.810 122.985 191.085 ;
        RECT 121.455 190.450 122.985 190.640 ;
        RECT 120.775 190.110 121.800 190.280 ;
        RECT 123.155 190.270 123.325 191.230 ;
        RECT 123.955 191.210 124.125 191.670 ;
        RECT 124.295 191.380 124.855 192.070 ;
        RECT 125.025 191.670 125.705 191.955 ;
        RECT 125.875 191.700 126.045 192.700 ;
        RECT 126.685 192.690 128.025 192.815 ;
        RECT 126.255 192.645 128.025 192.690 ;
        RECT 128.595 192.730 129.265 193.060 ;
        RECT 130.465 193.045 130.635 194.185 ;
        RECT 128.595 192.660 128.765 192.730 ;
        RECT 126.255 192.360 126.855 192.645 ;
        RECT 127.025 192.230 127.685 192.475 ;
        RECT 126.265 191.930 126.855 192.180 ;
        RECT 127.855 192.160 128.025 192.645 ;
        RECT 128.195 192.330 128.765 192.660 ;
        RECT 129.675 192.535 130.005 192.945 ;
        RECT 130.175 192.725 130.635 193.045 ;
        RECT 125.025 191.210 125.245 191.670 ;
        RECT 125.875 191.500 126.515 191.700 ;
        RECT 125.415 191.370 126.515 191.500 ;
        RECT 125.415 191.230 126.045 191.370 ;
        RECT 123.955 191.000 125.245 191.210 ;
        RECT 123.495 190.430 125.705 190.830 ;
        RECT 125.875 190.700 126.045 191.230 ;
        RECT 126.685 191.140 126.855 191.930 ;
        RECT 127.025 191.750 127.685 192.015 ;
        RECT 127.855 191.830 128.365 192.160 ;
        RECT 128.595 192.120 128.765 192.330 ;
        RECT 128.985 192.530 130.005 192.535 ;
        RECT 128.985 192.290 130.600 192.530 ;
        RECT 130.805 192.305 131.095 194.355 ;
        RECT 131.315 193.450 131.485 194.525 ;
        RECT 134.035 193.450 134.205 195.010 ;
        RECT 136.755 194.380 136.925 195.430 ;
        RECT 137.145 194.550 137.435 196.205 ;
        RECT 137.605 195.885 138.065 196.205 ;
        RECT 137.605 194.785 137.775 195.885 ;
        RECT 138.235 195.855 138.805 196.205 ;
        RECT 139.475 196.200 140.105 196.220 ;
        RECT 138.975 195.970 140.105 196.200 ;
        RECT 140.275 196.025 141.225 196.305 ;
        RECT 142.195 196.235 142.365 196.830 ;
        RECT 142.535 196.410 143.465 196.580 ;
        RECT 141.735 196.195 142.365 196.235 ;
        RECT 141.735 195.970 143.125 196.195 ;
        RECT 138.975 195.870 139.645 195.970 ;
        RECT 137.945 194.975 138.565 195.685 ;
        RECT 138.735 195.500 139.255 195.670 ;
        RECT 137.605 194.615 138.065 194.785 ;
        RECT 136.755 194.100 137.725 194.380 ;
        RECT 137.895 194.230 138.065 194.615 ;
        RECT 138.235 194.400 138.565 194.805 ;
        RECT 138.735 194.800 138.905 195.500 ;
        RECT 139.475 195.300 139.645 195.870 ;
        RECT 142.195 195.865 143.125 195.970 ;
        RECT 143.295 196.035 143.465 196.410 ;
        RECT 143.645 196.315 144.015 196.670 ;
        RECT 144.195 196.410 144.745 196.580 ;
        RECT 144.195 196.035 144.365 196.410 ;
        RECT 144.915 196.195 145.085 197.005 ;
        RECT 145.255 196.870 147.465 197.270 ;
        RECT 145.255 196.400 145.885 196.680 ;
        RECT 143.295 195.865 144.365 196.035 ;
        RECT 144.535 195.880 145.085 196.195 ;
        RECT 145.715 196.005 145.885 196.400 ;
        RECT 146.055 196.175 146.615 196.870 ;
        RECT 146.785 196.400 147.465 196.680 ;
        RECT 146.785 196.005 147.005 196.400 ;
        RECT 144.535 195.865 145.545 195.880 ;
        RECT 140.235 195.800 141.600 195.855 ;
        RECT 139.925 195.685 142.025 195.800 ;
        RECT 139.925 195.630 140.365 195.685 ;
        RECT 139.925 195.465 140.095 195.630 ;
        RECT 141.470 195.550 142.025 195.685 ;
        RECT 139.075 194.970 139.645 195.300 ;
        RECT 138.735 194.630 139.255 194.800 ;
        RECT 138.735 194.230 138.905 194.630 ;
        RECT 139.475 194.460 139.645 194.970 ;
        RECT 139.925 194.765 140.095 195.270 ;
        RECT 140.295 195.105 140.515 195.460 ;
        RECT 140.685 195.275 141.280 195.515 ;
        RECT 140.295 194.935 141.580 195.105 ;
        RECT 139.925 194.595 141.045 194.765 ;
        RECT 134.385 193.600 136.585 193.910 ;
        RECT 134.385 193.470 134.945 193.600 ;
        RECT 135.955 193.470 136.585 193.600 ;
        RECT 131.315 193.160 132.650 193.450 ;
        RECT 133.310 193.300 134.205 193.450 ;
        RECT 136.755 193.450 136.925 194.100 ;
        RECT 137.895 194.060 138.905 194.230 ;
        RECT 139.075 194.275 139.645 194.460 ;
        RECT 140.875 194.405 141.045 194.595 ;
        RECT 141.215 194.575 141.580 194.935 ;
        RECT 141.750 194.405 141.920 195.340 ;
        RECT 139.075 194.080 140.145 194.275 ;
        RECT 138.235 193.960 138.565 194.060 ;
        RECT 139.475 193.905 140.145 194.080 ;
        RECT 140.325 194.185 140.655 194.385 ;
        RECT 140.875 194.235 141.920 194.405 ;
        RECT 142.195 195.265 142.365 195.865 ;
        RECT 143.675 195.780 144.005 195.865 ;
        RECT 142.535 195.610 143.440 195.695 ;
        RECT 144.170 195.610 144.745 195.695 ;
        RECT 142.535 195.440 144.745 195.610 ;
        RECT 144.915 195.555 145.545 195.865 ;
        RECT 145.715 195.555 147.005 196.005 ;
        RECT 147.635 195.880 147.805 197.670 ;
        RECT 147.175 195.555 147.805 195.880 ;
        RECT 144.915 195.265 145.085 195.555 ;
        RECT 145.995 195.450 146.325 195.555 ;
        RECT 142.195 195.005 143.515 195.265 ;
        RECT 144.075 195.005 145.085 195.265 ;
        RECT 142.195 194.790 142.365 195.005 ;
        RECT 142.195 194.560 143.505 194.790 ;
        RECT 137.095 193.790 138.065 193.890 ;
        RECT 138.800 193.790 139.145 193.890 ;
        RECT 137.095 193.620 139.145 193.790 ;
        RECT 139.475 193.450 139.645 193.905 ;
        RECT 140.325 193.725 140.625 194.185 ;
        RECT 140.875 194.065 141.135 194.235 ;
        RECT 142.195 194.065 142.365 194.560 ;
        RECT 143.675 194.480 143.925 194.810 ;
        RECT 144.915 194.790 145.085 195.005 ;
        RECT 145.255 195.280 145.825 195.385 ;
        RECT 146.495 195.280 147.465 195.385 ;
        RECT 145.255 195.000 147.465 195.280 ;
        RECT 144.095 194.560 145.085 194.790 ;
        RECT 145.255 194.570 145.805 194.740 ;
        RECT 144.915 194.390 145.085 194.560 ;
        RECT 140.805 193.895 141.135 194.065 ;
        RECT 141.395 193.895 142.365 194.065 ;
        RECT 142.535 194.310 143.515 194.390 ;
        RECT 144.115 194.310 144.745 194.390 ;
        RECT 142.535 194.060 144.745 194.310 ;
        RECT 144.915 194.060 145.465 194.390 ;
        RECT 145.635 194.245 145.805 194.570 ;
        RECT 145.985 194.470 146.355 194.810 ;
        RECT 146.535 194.570 147.465 194.750 ;
        RECT 146.535 194.245 146.705 194.570 ;
        RECT 147.635 194.390 147.805 195.555 ;
        RECT 145.635 194.075 146.705 194.245 ;
        RECT 142.195 193.890 142.365 193.895 ;
        RECT 144.915 193.890 145.085 194.060 ;
        RECT 146.060 193.970 146.390 194.075 ;
        RECT 146.875 194.060 147.805 194.390 ;
        RECT 133.310 193.160 134.945 193.300 ;
        RECT 135.115 193.260 135.735 193.430 ;
        RECT 136.755 193.295 138.090 193.450 ;
        RECT 131.315 192.120 131.485 193.160 ;
        RECT 127.025 191.270 127.685 191.555 ;
        RECT 126.265 190.890 126.855 191.140 ;
        RECT 127.025 190.880 127.685 191.095 ;
        RECT 127.355 190.790 127.685 190.880 ;
        RECT 125.875 190.450 127.185 190.700 ;
        RECT 127.855 190.620 128.025 191.830 ;
        RECT 128.595 191.780 129.265 192.120 ;
        RECT 129.435 191.780 130.005 192.120 ;
        RECT 130.240 191.780 131.485 192.120 ;
        RECT 131.705 191.800 131.995 192.990 ;
        RECT 132.165 192.645 132.625 192.970 ;
        RECT 132.795 192.645 133.125 192.990 ;
        RECT 133.295 192.720 133.815 192.975 ;
        RECT 134.035 192.850 134.945 193.160 ;
        RECT 132.165 191.970 132.335 192.645 ;
        RECT 132.505 192.280 133.125 192.475 ;
        RECT 132.165 191.800 132.625 191.970 ;
        RECT 128.595 191.590 128.765 191.780 ;
        RECT 131.315 191.630 131.485 191.780 ;
        RECT 128.595 191.350 129.575 191.590 ;
        RECT 128.595 190.780 128.765 191.350 ;
        RECT 129.755 191.260 130.005 191.610 ;
        RECT 130.175 191.270 131.130 191.600 ;
        RECT 131.315 191.350 132.285 191.630 ;
        RECT 132.455 191.480 132.625 191.800 ;
        RECT 132.795 191.650 133.125 192.280 ;
        RECT 133.295 192.050 133.465 192.720 ;
        RECT 134.035 192.550 134.205 192.850 ;
        RECT 135.115 192.700 135.395 193.090 ;
        RECT 135.565 192.810 135.735 193.260 ;
        RECT 135.905 193.160 138.090 193.295 ;
        RECT 138.750 193.160 139.645 193.450 ;
        RECT 139.925 193.555 142.025 193.725 ;
        RECT 139.925 193.320 140.095 193.555 ;
        RECT 141.695 193.475 142.025 193.555 ;
        RECT 142.195 193.680 143.505 193.890 ;
        RECT 144.095 193.680 145.085 193.890 ;
        RECT 142.195 193.450 142.365 193.680 ;
        RECT 144.915 193.450 145.085 193.680 ;
        RECT 145.255 193.800 145.760 193.880 ;
        RECT 146.560 193.800 147.465 193.890 ;
        RECT 145.255 193.620 147.465 193.800 ;
        RECT 147.635 193.450 147.805 194.060 ;
        RECT 140.805 193.195 141.525 193.385 ;
        RECT 135.905 192.980 136.925 193.160 ;
        RECT 133.635 192.340 134.205 192.550 ;
        RECT 134.375 192.510 134.945 192.680 ;
        RECT 135.565 192.640 136.585 192.810 ;
        RECT 133.635 192.220 134.605 192.340 ;
        RECT 133.295 191.880 133.815 192.050 ;
        RECT 134.035 191.920 134.605 192.220 ;
        RECT 133.295 191.480 133.465 191.880 ;
        RECT 134.035 191.710 134.205 191.920 ;
        RECT 134.775 191.750 134.945 192.510 ;
        RECT 135.115 192.470 135.445 192.515 ;
        RECT 135.115 192.270 136.245 192.470 ;
        RECT 135.115 191.820 136.245 192.070 ;
        RECT 128.935 191.090 129.575 191.180 ;
        RECT 130.175 191.090 130.345 191.270 ;
        RECT 128.935 190.920 130.345 191.090 ;
        RECT 128.935 190.850 129.575 190.920 ;
        RECT 127.355 190.450 128.025 190.620 ;
        RECT 128.195 190.680 128.765 190.780 ;
        RECT 128.195 190.450 129.575 190.680 ;
        RECT 120.435 189.770 121.365 189.940 ;
        RECT 117.715 189.490 118.695 189.760 ;
        RECT 113.895 189.100 114.825 189.280 ;
        RECT 114.995 188.380 115.165 189.460 ;
        RECT 117.715 188.820 117.885 189.490 ;
        RECT 118.875 189.420 119.125 189.770 ;
        RECT 120.435 189.760 120.605 189.770 ;
        RECT 119.295 189.430 120.605 189.760 ;
        RECT 118.055 189.250 118.695 189.320 ;
        RECT 118.055 189.080 119.465 189.250 ;
        RECT 118.055 188.990 118.695 189.080 ;
        RECT 117.715 188.580 118.695 188.820 ;
        RECT 114.995 188.050 115.885 188.380 ;
        RECT 116.185 188.160 116.725 188.390 ;
        RECT 116.525 188.060 116.725 188.160 ;
        RECT 116.895 188.050 117.545 188.390 ;
        RECT 13.380 187.675 92.040 187.845 ;
        RECT 13.465 186.925 14.675 187.675 ;
        RECT 14.845 187.130 20.190 187.675 ;
        RECT 13.465 186.385 13.985 186.925 ;
        RECT 14.155 186.215 14.675 186.755 ;
        RECT 16.430 186.300 16.770 187.130 ;
        RECT 20.365 186.925 21.575 187.675 ;
        RECT 21.745 187.025 22.005 187.505 ;
        RECT 22.175 187.135 22.425 187.675 ;
        RECT 13.465 185.125 14.675 186.215 ;
        RECT 18.250 185.560 18.600 186.810 ;
        RECT 20.365 186.385 20.885 186.925 ;
        RECT 21.055 186.215 21.575 186.755 ;
        RECT 14.845 185.125 20.190 185.560 ;
        RECT 20.365 185.125 21.575 186.215 ;
        RECT 21.745 185.995 21.915 187.025 ;
        RECT 22.595 186.970 22.815 187.455 ;
        RECT 22.085 186.375 22.315 186.770 ;
        RECT 22.485 186.545 22.815 186.970 ;
        RECT 22.985 187.295 23.875 187.465 ;
        RECT 22.985 186.570 23.155 187.295 ;
        RECT 23.325 186.740 23.875 187.125 ;
        RECT 24.045 186.905 27.555 187.675 ;
        RECT 27.815 187.125 27.985 187.415 ;
        RECT 28.155 187.295 28.485 187.675 ;
        RECT 27.815 186.955 28.480 187.125 ;
        RECT 22.985 186.500 23.875 186.570 ;
        RECT 22.980 186.475 23.875 186.500 ;
        RECT 22.970 186.460 23.875 186.475 ;
        RECT 22.965 186.445 23.875 186.460 ;
        RECT 22.955 186.440 23.875 186.445 ;
        RECT 22.950 186.430 23.875 186.440 ;
        RECT 22.945 186.420 23.875 186.430 ;
        RECT 22.935 186.415 23.875 186.420 ;
        RECT 22.925 186.405 23.875 186.415 ;
        RECT 22.915 186.400 23.875 186.405 ;
        RECT 22.915 186.395 23.250 186.400 ;
        RECT 22.900 186.390 23.250 186.395 ;
        RECT 22.885 186.380 23.250 186.390 ;
        RECT 22.860 186.375 23.250 186.380 ;
        RECT 22.085 186.370 23.250 186.375 ;
        RECT 22.085 186.335 23.220 186.370 ;
        RECT 22.085 186.310 23.185 186.335 ;
        RECT 22.085 186.280 23.155 186.310 ;
        RECT 22.085 186.250 23.135 186.280 ;
        RECT 22.085 186.220 23.115 186.250 ;
        RECT 22.085 186.210 23.045 186.220 ;
        RECT 22.085 186.200 23.020 186.210 ;
        RECT 22.085 186.185 23.000 186.200 ;
        RECT 22.085 186.170 22.980 186.185 ;
        RECT 22.190 186.160 22.975 186.170 ;
        RECT 22.190 186.125 22.960 186.160 ;
        RECT 21.745 185.295 22.020 185.995 ;
        RECT 22.190 185.875 22.945 186.125 ;
        RECT 23.115 185.805 23.445 186.050 ;
        RECT 23.615 185.950 23.875 186.400 ;
        RECT 24.045 186.385 25.695 186.905 ;
        RECT 25.865 186.215 27.555 186.735 ;
        RECT 23.260 185.780 23.445 185.805 ;
        RECT 23.260 185.680 23.875 185.780 ;
        RECT 22.190 185.125 22.445 185.670 ;
        RECT 22.615 185.295 23.095 185.635 ;
        RECT 23.270 185.125 23.875 185.680 ;
        RECT 24.045 185.125 27.555 186.215 ;
        RECT 27.730 186.135 28.080 186.785 ;
        RECT 28.250 185.965 28.480 186.955 ;
        RECT 27.815 185.795 28.480 185.965 ;
        RECT 27.815 185.295 27.985 185.795 ;
        RECT 28.155 185.125 28.485 185.625 ;
        RECT 28.655 185.295 28.840 187.415 ;
        RECT 29.095 187.215 29.345 187.675 ;
        RECT 29.515 187.225 29.850 187.395 ;
        RECT 30.045 187.225 30.720 187.395 ;
        RECT 29.515 187.085 29.685 187.225 ;
        RECT 29.010 186.095 29.290 187.045 ;
        RECT 29.460 186.955 29.685 187.085 ;
        RECT 29.460 185.850 29.630 186.955 ;
        RECT 29.855 186.805 30.380 187.025 ;
        RECT 29.800 186.040 30.040 186.635 ;
        RECT 30.210 186.105 30.380 186.805 ;
        RECT 30.550 186.445 30.720 187.225 ;
        RECT 31.040 187.175 31.410 187.675 ;
        RECT 31.590 187.225 31.995 187.395 ;
        RECT 32.165 187.225 32.950 187.395 ;
        RECT 31.590 186.995 31.760 187.225 ;
        RECT 30.930 186.695 31.760 186.995 ;
        RECT 32.145 186.725 32.610 187.055 ;
        RECT 30.930 186.665 31.130 186.695 ;
        RECT 31.250 186.445 31.420 186.515 ;
        RECT 30.550 186.275 31.420 186.445 ;
        RECT 30.910 186.185 31.420 186.275 ;
        RECT 29.460 185.720 29.765 185.850 ;
        RECT 30.210 185.740 30.740 186.105 ;
        RECT 29.080 185.125 29.345 185.585 ;
        RECT 29.515 185.295 29.765 185.720 ;
        RECT 30.910 185.570 31.080 186.185 ;
        RECT 29.975 185.400 31.080 185.570 ;
        RECT 31.250 185.125 31.420 185.925 ;
        RECT 31.590 185.625 31.760 186.695 ;
        RECT 31.930 185.795 32.120 186.515 ;
        RECT 32.290 185.765 32.610 186.725 ;
        RECT 32.780 186.765 32.950 187.225 ;
        RECT 33.225 187.145 33.435 187.675 ;
        RECT 33.695 186.935 34.025 187.460 ;
        RECT 34.195 187.065 34.365 187.675 ;
        RECT 34.535 187.020 34.865 187.455 ;
        RECT 34.535 186.935 34.915 187.020 ;
        RECT 33.825 186.765 34.025 186.935 ;
        RECT 34.690 186.895 34.915 186.935 ;
        RECT 32.780 186.435 33.655 186.765 ;
        RECT 33.825 186.435 34.575 186.765 ;
        RECT 31.590 185.295 31.840 185.625 ;
        RECT 32.780 185.595 32.950 186.435 ;
        RECT 33.825 186.230 34.015 186.435 ;
        RECT 34.745 186.315 34.915 186.895 ;
        RECT 35.085 186.905 38.595 187.675 ;
        RECT 39.225 186.950 39.515 187.675 ;
        RECT 39.775 187.125 39.945 187.415 ;
        RECT 40.115 187.295 40.445 187.675 ;
        RECT 39.775 186.955 40.440 187.125 ;
        RECT 35.085 186.385 36.735 186.905 ;
        RECT 34.700 186.265 34.915 186.315 ;
        RECT 33.120 185.855 34.015 186.230 ;
        RECT 34.525 186.185 34.915 186.265 ;
        RECT 36.905 186.215 38.595 186.735 ;
        RECT 32.065 185.425 32.950 185.595 ;
        RECT 33.130 185.125 33.445 185.625 ;
        RECT 33.675 185.295 34.015 185.855 ;
        RECT 34.185 185.125 34.355 186.135 ;
        RECT 34.525 185.340 34.855 186.185 ;
        RECT 35.085 185.125 38.595 186.215 ;
        RECT 39.225 185.125 39.515 186.290 ;
        RECT 39.690 186.135 40.040 186.785 ;
        RECT 40.210 185.965 40.440 186.955 ;
        RECT 39.775 185.795 40.440 185.965 ;
        RECT 39.775 185.295 39.945 185.795 ;
        RECT 40.115 185.125 40.445 185.625 ;
        RECT 40.615 185.295 40.800 187.415 ;
        RECT 41.055 187.215 41.305 187.675 ;
        RECT 41.475 187.225 41.810 187.395 ;
        RECT 42.005 187.225 42.680 187.395 ;
        RECT 41.475 187.085 41.645 187.225 ;
        RECT 40.970 186.095 41.250 187.045 ;
        RECT 41.420 186.955 41.645 187.085 ;
        RECT 41.420 185.850 41.590 186.955 ;
        RECT 41.815 186.805 42.340 187.025 ;
        RECT 41.760 186.040 42.000 186.635 ;
        RECT 42.170 186.105 42.340 186.805 ;
        RECT 42.510 186.445 42.680 187.225 ;
        RECT 43.000 187.175 43.370 187.675 ;
        RECT 43.550 187.225 43.955 187.395 ;
        RECT 44.125 187.225 44.910 187.395 ;
        RECT 43.550 186.995 43.720 187.225 ;
        RECT 42.890 186.695 43.720 186.995 ;
        RECT 44.105 186.725 44.570 187.055 ;
        RECT 42.890 186.665 43.090 186.695 ;
        RECT 43.210 186.445 43.380 186.515 ;
        RECT 42.510 186.275 43.380 186.445 ;
        RECT 42.870 186.185 43.380 186.275 ;
        RECT 41.420 185.720 41.725 185.850 ;
        RECT 42.170 185.740 42.700 186.105 ;
        RECT 41.040 185.125 41.305 185.585 ;
        RECT 41.475 185.295 41.725 185.720 ;
        RECT 42.870 185.570 43.040 186.185 ;
        RECT 41.935 185.400 43.040 185.570 ;
        RECT 43.210 185.125 43.380 185.925 ;
        RECT 43.550 185.625 43.720 186.695 ;
        RECT 43.890 185.795 44.080 186.515 ;
        RECT 44.250 185.765 44.570 186.725 ;
        RECT 44.740 186.765 44.910 187.225 ;
        RECT 45.185 187.145 45.395 187.675 ;
        RECT 45.655 186.935 45.985 187.460 ;
        RECT 46.155 187.065 46.325 187.675 ;
        RECT 46.495 187.020 46.825 187.455 ;
        RECT 47.045 187.130 52.390 187.675 ;
        RECT 46.495 186.935 46.875 187.020 ;
        RECT 45.785 186.765 45.985 186.935 ;
        RECT 46.650 186.895 46.875 186.935 ;
        RECT 44.740 186.435 45.615 186.765 ;
        RECT 45.785 186.435 46.535 186.765 ;
        RECT 43.550 185.295 43.800 185.625 ;
        RECT 44.740 185.595 44.910 186.435 ;
        RECT 45.785 186.230 45.975 186.435 ;
        RECT 46.705 186.315 46.875 186.895 ;
        RECT 46.660 186.265 46.875 186.315 ;
        RECT 48.630 186.300 48.970 187.130 ;
        RECT 52.565 186.905 56.075 187.675 ;
        RECT 56.715 186.945 57.015 187.675 ;
        RECT 45.080 185.855 45.975 186.230 ;
        RECT 46.485 186.185 46.875 186.265 ;
        RECT 44.025 185.425 44.910 185.595 ;
        RECT 45.090 185.125 45.405 185.625 ;
        RECT 45.635 185.295 45.975 185.855 ;
        RECT 46.145 185.125 46.315 186.135 ;
        RECT 46.485 185.340 46.815 186.185 ;
        RECT 50.450 185.560 50.800 186.810 ;
        RECT 52.565 186.385 54.215 186.905 ;
        RECT 57.195 186.765 57.425 187.385 ;
        RECT 57.625 187.115 57.850 187.495 ;
        RECT 58.020 187.285 58.350 187.675 ;
        RECT 57.625 186.935 57.955 187.115 ;
        RECT 54.385 186.215 56.075 186.735 ;
        RECT 56.720 186.435 57.015 186.765 ;
        RECT 57.195 186.435 57.610 186.765 ;
        RECT 57.780 186.265 57.955 186.935 ;
        RECT 58.125 186.435 58.365 187.085 ;
        RECT 58.545 186.905 60.215 187.675 ;
        RECT 60.850 187.145 61.140 187.495 ;
        RECT 61.335 187.315 61.665 187.675 ;
        RECT 61.835 187.145 62.065 187.450 ;
        RECT 60.850 186.975 62.065 187.145 ;
        RECT 58.545 186.385 59.295 186.905 ;
        RECT 62.255 186.805 62.425 187.370 ;
        RECT 47.045 185.125 52.390 185.560 ;
        RECT 52.565 185.125 56.075 186.215 ;
        RECT 56.715 185.905 57.610 186.235 ;
        RECT 57.780 186.075 58.365 186.265 ;
        RECT 59.465 186.215 60.215 186.735 ;
        RECT 60.910 186.655 61.170 186.765 ;
        RECT 60.905 186.485 61.170 186.655 ;
        RECT 60.910 186.435 61.170 186.485 ;
        RECT 61.350 186.435 61.735 186.765 ;
        RECT 61.905 186.635 62.425 186.805 ;
        RECT 62.685 186.905 64.355 187.675 ;
        RECT 64.985 186.950 65.275 187.675 ;
        RECT 65.445 187.130 70.790 187.675 ;
        RECT 70.965 187.130 76.310 187.675 ;
        RECT 76.485 187.130 81.830 187.675 ;
        RECT 82.005 187.130 87.350 187.675 ;
        RECT 56.715 185.735 57.920 185.905 ;
        RECT 56.715 185.305 57.045 185.735 ;
        RECT 57.225 185.125 57.420 185.565 ;
        RECT 57.590 185.305 57.920 185.735 ;
        RECT 58.090 185.305 58.365 186.075 ;
        RECT 58.545 185.125 60.215 186.215 ;
        RECT 60.850 185.125 61.170 186.265 ;
        RECT 61.350 185.385 61.545 186.435 ;
        RECT 61.905 186.255 62.075 186.635 ;
        RECT 61.725 185.975 62.075 186.255 ;
        RECT 62.265 186.105 62.510 186.465 ;
        RECT 62.685 186.385 63.435 186.905 ;
        RECT 63.605 186.215 64.355 186.735 ;
        RECT 67.030 186.300 67.370 187.130 ;
        RECT 61.725 185.295 62.055 185.975 ;
        RECT 62.255 185.125 62.510 185.925 ;
        RECT 62.685 185.125 64.355 186.215 ;
        RECT 64.985 185.125 65.275 186.290 ;
        RECT 68.850 185.560 69.200 186.810 ;
        RECT 72.550 186.300 72.890 187.130 ;
        RECT 74.370 185.560 74.720 186.810 ;
        RECT 78.070 186.300 78.410 187.130 ;
        RECT 79.890 185.560 80.240 186.810 ;
        RECT 83.590 186.300 83.930 187.130 ;
        RECT 87.525 186.905 90.115 187.675 ;
        RECT 90.745 186.925 91.955 187.675 ;
        RECT 85.410 185.560 85.760 186.810 ;
        RECT 87.525 186.385 88.735 186.905 ;
        RECT 88.905 186.215 90.115 186.735 ;
        RECT 65.445 185.125 70.790 185.560 ;
        RECT 70.965 185.125 76.310 185.560 ;
        RECT 76.485 185.125 81.830 185.560 ;
        RECT 82.005 185.125 87.350 185.560 ;
        RECT 87.525 185.125 90.115 186.215 ;
        RECT 90.745 186.215 91.265 186.755 ;
        RECT 91.435 186.385 91.955 186.925 ;
        RECT 112.275 187.590 112.950 187.925 ;
        RECT 90.745 185.125 91.955 186.215 ;
        RECT 112.275 186.165 112.445 187.590 ;
        RECT 113.125 187.570 113.975 187.870 ;
        RECT 114.145 187.670 114.805 187.840 ;
        RECT 112.640 187.400 113.015 187.420 ;
        RECT 114.145 187.400 114.375 187.670 ;
        RECT 114.995 187.500 115.165 188.050 ;
        RECT 115.410 187.750 116.705 187.870 ;
        RECT 115.410 187.655 116.725 187.750 ;
        RECT 112.640 187.180 114.375 187.400 ;
        RECT 113.165 187.165 114.375 187.180 ;
        RECT 114.545 187.170 115.165 187.500 ;
        RECT 112.630 186.730 112.970 186.900 ;
        RECT 113.165 186.865 113.495 187.165 ;
        RECT 112.775 186.695 112.970 186.730 ;
        RECT 113.665 186.710 114.780 186.995 ;
        RECT 114.995 186.960 115.165 187.170 ;
        RECT 115.335 187.130 116.325 187.460 ;
        RECT 116.525 187.420 116.725 187.655 ;
        RECT 116.895 187.540 117.085 188.050 ;
        RECT 117.715 187.880 117.885 188.580 ;
        RECT 118.875 188.560 119.125 188.910 ;
        RECT 119.295 188.900 119.465 189.080 ;
        RECT 119.295 188.570 120.250 188.900 ;
        RECT 120.435 188.410 120.605 189.430 ;
        RECT 120.955 189.360 121.365 189.535 ;
        RECT 121.610 189.530 121.800 190.110 ;
        RECT 122.175 189.540 122.345 190.250 ;
        RECT 122.620 189.760 123.325 190.270 ;
        RECT 123.495 189.960 124.125 190.240 ;
        RECT 122.175 189.360 122.950 189.540 ;
        RECT 120.955 189.295 122.950 189.360 ;
        RECT 123.155 189.440 123.325 189.760 ;
        RECT 123.955 189.565 124.125 189.960 ;
        RECT 124.295 189.735 124.855 190.430 ;
        RECT 125.025 189.960 125.705 190.240 ;
        RECT 125.025 189.565 125.245 189.960 ;
        RECT 120.955 189.020 122.345 189.295 ;
        RECT 123.155 189.115 123.785 189.440 ;
        RECT 123.955 189.115 125.245 189.565 ;
        RECT 125.875 189.440 126.045 190.450 ;
        RECT 127.355 190.310 127.685 190.450 ;
        RECT 128.595 190.410 129.575 190.450 ;
        RECT 126.255 190.140 127.105 190.280 ;
        RECT 127.870 190.140 128.380 190.280 ;
        RECT 126.255 189.950 128.380 190.140 ;
        RECT 125.415 189.115 126.045 189.440 ;
        RECT 120.775 188.590 121.705 188.760 ;
        RECT 118.250 188.135 120.265 188.390 ;
        RECT 118.250 188.030 118.625 188.135 ;
        RECT 119.280 188.050 120.265 188.135 ;
        RECT 120.435 188.080 121.365 188.410 ;
        RECT 121.535 188.265 121.705 188.590 ;
        RECT 121.885 188.500 122.255 188.830 ;
        RECT 122.435 188.590 122.985 188.760 ;
        RECT 122.435 188.265 122.605 188.590 ;
        RECT 123.155 188.410 123.325 189.115 ;
        RECT 124.235 189.010 124.565 189.115 ;
        RECT 123.495 188.840 124.065 188.945 ;
        RECT 124.735 188.840 125.705 188.945 ;
        RECT 123.495 188.560 125.705 188.840 ;
        RECT 125.875 188.635 126.045 189.115 ;
        RECT 128.595 189.790 128.765 190.410 ;
        RECT 129.755 190.400 130.005 190.750 ;
        RECT 131.315 190.740 131.485 191.350 ;
        RECT 132.455 191.310 133.465 191.480 ;
        RECT 133.635 191.330 134.205 191.710 ;
        RECT 134.375 191.520 134.945 191.750 ;
        RECT 136.415 191.630 136.585 192.640 ;
        RECT 132.795 191.205 133.125 191.310 ;
        RECT 131.655 191.035 132.625 191.140 ;
        RECT 133.360 191.035 133.705 191.140 ;
        RECT 131.655 190.865 133.705 191.035 ;
        RECT 130.175 190.690 131.485 190.740 ;
        RECT 134.035 190.690 134.205 191.330 ;
        RECT 134.375 191.030 134.945 191.350 ;
        RECT 135.115 191.200 135.445 191.605 ;
        RECT 135.615 191.380 136.585 191.630 ;
        RECT 136.755 192.480 136.925 192.980 ;
        RECT 137.095 192.735 139.110 192.990 ;
        RECT 137.095 192.650 138.080 192.735 ;
        RECT 138.735 192.630 139.110 192.735 ;
        RECT 138.235 192.480 138.565 192.565 ;
        RECT 136.755 192.070 137.355 192.480 ;
        RECT 137.525 192.215 138.565 192.480 ;
        RECT 139.475 192.365 139.645 193.160 ;
        RECT 139.925 192.535 140.095 193.150 ;
        RECT 140.265 193.025 140.595 193.170 ;
        RECT 140.265 192.705 141.555 193.025 ;
        RECT 141.725 192.535 141.895 193.250 ;
        RECT 139.925 192.365 141.895 192.535 ;
        RECT 142.195 193.160 143.530 193.450 ;
        RECT 144.190 193.160 145.810 193.450 ;
        RECT 146.470 193.160 147.805 193.450 ;
        RECT 142.195 192.375 142.365 193.160 ;
        RECT 142.535 192.680 144.735 192.990 ;
        RECT 142.535 192.550 143.165 192.680 ;
        RECT 144.175 192.550 144.735 192.680 ;
        RECT 135.615 191.030 135.785 191.380 ;
        RECT 136.755 191.325 136.925 192.070 ;
        RECT 136.755 191.200 137.345 191.325 ;
        RECT 134.375 190.860 135.785 191.030 ;
        RECT 135.955 190.995 137.345 191.200 ;
        RECT 137.525 191.205 137.695 192.215 ;
        RECT 138.735 192.195 139.645 192.365 ;
        RECT 139.475 192.090 139.645 192.195 ;
        RECT 137.865 191.545 138.035 192.000 ;
        RECT 138.235 191.715 138.565 192.045 ;
        RECT 138.735 191.745 139.110 191.915 ;
        RECT 139.475 191.880 140.175 192.090 ;
        RECT 138.735 191.545 138.905 191.745 ;
        RECT 137.865 191.375 138.905 191.545 ;
        RECT 137.525 191.035 139.305 191.205 ;
        RECT 139.475 191.120 139.645 191.880 ;
        RECT 140.555 191.660 140.885 192.365 ;
        RECT 141.090 191.640 141.465 192.195 ;
        RECT 142.195 192.185 143.215 192.375 ;
        RECT 141.695 192.060 143.215 192.185 ;
        RECT 143.385 192.340 144.005 192.510 ;
        RECT 144.915 192.380 145.085 193.160 ;
        RECT 141.695 191.870 142.365 192.060 ;
        RECT 143.385 191.890 143.555 192.340 ;
        RECT 139.860 191.490 140.385 191.620 ;
        RECT 141.090 191.490 142.025 191.640 ;
        RECT 139.860 191.300 142.025 191.490 ;
        RECT 139.860 191.290 140.885 191.300 ;
        RECT 135.955 190.870 136.925 190.995 ;
        RECT 130.175 190.410 132.575 190.690 ;
        RECT 128.935 189.970 129.485 190.140 ;
        RECT 128.595 189.460 129.145 189.790 ;
        RECT 129.315 189.645 129.485 189.970 ;
        RECT 129.665 189.870 130.035 190.210 ;
        RECT 130.215 189.970 131.145 190.150 ;
        RECT 130.215 189.645 130.385 189.970 ;
        RECT 131.315 189.790 132.575 190.410 ;
        RECT 129.315 189.475 130.385 189.645 ;
        RECT 121.535 188.095 122.605 188.265 ;
        RECT 117.255 187.765 117.885 187.880 ;
        RECT 118.795 187.880 119.125 187.965 ;
        RECT 120.435 187.880 120.605 188.080 ;
        RECT 121.850 187.980 122.180 188.095 ;
        RECT 122.775 188.080 123.325 188.410 ;
        RECT 117.255 187.710 118.625 187.765 ;
        RECT 117.715 187.595 118.625 187.710 ;
        RECT 118.795 187.615 119.835 187.880 ;
        RECT 113.665 186.695 113.835 186.710 ;
        RECT 112.775 186.525 113.835 186.695 ;
        RECT 112.275 185.770 112.940 186.165 ;
        RECT 113.305 186.135 113.835 186.525 ;
        RECT 13.380 184.955 92.040 185.125 ;
        RECT 13.465 183.865 14.675 184.955 ;
        RECT 14.845 183.865 17.435 184.955 ;
        RECT 13.465 183.155 13.985 183.695 ;
        RECT 14.155 183.325 14.675 183.865 ;
        RECT 14.845 183.175 16.055 183.695 ;
        RECT 16.225 183.345 17.435 183.865 ;
        RECT 17.605 183.815 17.885 184.955 ;
        RECT 18.055 183.805 18.385 184.785 ;
        RECT 18.555 183.815 18.815 184.955 ;
        RECT 19.045 183.895 19.375 184.740 ;
        RECT 19.545 183.945 19.715 184.955 ;
        RECT 19.885 184.225 20.225 184.785 ;
        RECT 20.455 184.455 20.770 184.955 ;
        RECT 20.950 184.485 21.835 184.655 ;
        RECT 18.985 183.815 19.375 183.895 ;
        RECT 19.885 183.850 20.780 184.225 ;
        RECT 17.615 183.375 17.950 183.645 ;
        RECT 18.120 183.205 18.290 183.805 ;
        RECT 18.985 183.765 19.200 183.815 ;
        RECT 18.460 183.395 18.795 183.645 ;
        RECT 13.465 182.405 14.675 183.155 ;
        RECT 14.845 182.405 17.435 183.175 ;
        RECT 17.605 182.405 17.915 183.205 ;
        RECT 18.120 182.575 18.815 183.205 ;
        RECT 18.985 183.185 19.155 183.765 ;
        RECT 19.885 183.645 20.075 183.850 ;
        RECT 20.950 183.645 21.120 184.485 ;
        RECT 22.060 184.455 22.310 184.785 ;
        RECT 19.325 183.315 20.075 183.645 ;
        RECT 20.245 183.315 21.120 183.645 ;
        RECT 18.985 183.145 19.210 183.185 ;
        RECT 19.875 183.145 20.075 183.315 ;
        RECT 18.985 183.060 19.365 183.145 ;
        RECT 19.035 182.625 19.365 183.060 ;
        RECT 19.535 182.405 19.705 183.015 ;
        RECT 19.875 182.620 20.205 183.145 ;
        RECT 20.465 182.405 20.675 182.935 ;
        RECT 20.950 182.855 21.120 183.315 ;
        RECT 21.290 183.355 21.610 184.315 ;
        RECT 21.780 183.565 21.970 184.285 ;
        RECT 22.140 183.385 22.310 184.455 ;
        RECT 22.480 184.155 22.650 184.955 ;
        RECT 22.820 184.510 23.925 184.680 ;
        RECT 22.820 183.895 22.990 184.510 ;
        RECT 24.135 184.360 24.385 184.785 ;
        RECT 24.555 184.495 24.820 184.955 ;
        RECT 23.160 183.975 23.690 184.340 ;
        RECT 24.135 184.230 24.440 184.360 ;
        RECT 22.480 183.805 22.990 183.895 ;
        RECT 22.480 183.635 23.350 183.805 ;
        RECT 22.480 183.565 22.650 183.635 ;
        RECT 22.770 183.385 22.970 183.415 ;
        RECT 21.290 183.025 21.755 183.355 ;
        RECT 22.140 183.085 22.970 183.385 ;
        RECT 22.140 182.855 22.310 183.085 ;
        RECT 20.950 182.685 21.735 182.855 ;
        RECT 21.905 182.685 22.310 182.855 ;
        RECT 22.490 182.405 22.860 182.905 ;
        RECT 23.180 182.855 23.350 183.635 ;
        RECT 23.520 183.275 23.690 183.975 ;
        RECT 23.860 183.445 24.100 184.040 ;
        RECT 23.520 183.055 24.045 183.275 ;
        RECT 24.270 183.125 24.440 184.230 ;
        RECT 24.215 182.995 24.440 183.125 ;
        RECT 24.610 183.035 24.890 183.985 ;
        RECT 24.215 182.855 24.385 182.995 ;
        RECT 23.180 182.685 23.855 182.855 ;
        RECT 24.050 182.685 24.385 182.855 ;
        RECT 24.555 182.405 24.805 182.865 ;
        RECT 25.060 182.665 25.245 184.785 ;
        RECT 25.415 184.455 25.745 184.955 ;
        RECT 25.915 184.285 26.085 184.785 ;
        RECT 25.420 184.115 26.085 184.285 ;
        RECT 25.420 183.125 25.650 184.115 ;
        RECT 25.820 183.295 26.170 183.945 ;
        RECT 26.345 183.790 26.635 184.955 ;
        RECT 27.725 184.085 28.000 184.785 ;
        RECT 28.170 184.410 28.425 184.955 ;
        RECT 28.595 184.445 29.075 184.785 ;
        RECT 29.250 184.400 29.855 184.955 ;
        RECT 29.240 184.300 29.855 184.400 ;
        RECT 29.240 184.275 29.425 184.300 ;
        RECT 25.420 182.955 26.085 183.125 ;
        RECT 25.415 182.405 25.745 182.785 ;
        RECT 25.915 182.665 26.085 182.955 ;
        RECT 26.345 182.405 26.635 183.130 ;
        RECT 27.725 183.055 27.895 184.085 ;
        RECT 28.170 183.955 28.925 184.205 ;
        RECT 29.095 184.030 29.425 184.275 ;
        RECT 28.170 183.920 28.940 183.955 ;
        RECT 28.170 183.910 28.955 183.920 ;
        RECT 28.065 183.895 28.960 183.910 ;
        RECT 28.065 183.880 28.980 183.895 ;
        RECT 28.065 183.870 29.000 183.880 ;
        RECT 28.065 183.860 29.025 183.870 ;
        RECT 28.065 183.830 29.095 183.860 ;
        RECT 28.065 183.800 29.115 183.830 ;
        RECT 28.065 183.770 29.135 183.800 ;
        RECT 28.065 183.745 29.165 183.770 ;
        RECT 28.065 183.710 29.200 183.745 ;
        RECT 28.065 183.705 29.230 183.710 ;
        RECT 28.065 183.310 28.295 183.705 ;
        RECT 28.840 183.700 29.230 183.705 ;
        RECT 28.865 183.690 29.230 183.700 ;
        RECT 28.880 183.685 29.230 183.690 ;
        RECT 28.895 183.680 29.230 183.685 ;
        RECT 29.595 183.680 29.855 184.130 ;
        RECT 28.895 183.675 29.855 183.680 ;
        RECT 28.905 183.665 29.855 183.675 ;
        RECT 28.915 183.660 29.855 183.665 ;
        RECT 28.925 183.650 29.855 183.660 ;
        RECT 28.930 183.640 29.855 183.650 ;
        RECT 28.935 183.635 29.855 183.640 ;
        RECT 28.945 183.620 29.855 183.635 ;
        RECT 28.950 183.605 29.855 183.620 ;
        RECT 28.960 183.580 29.855 183.605 ;
        RECT 28.465 183.110 28.795 183.535 ;
        RECT 27.725 182.575 27.985 183.055 ;
        RECT 28.155 182.405 28.405 182.945 ;
        RECT 28.575 182.625 28.795 183.110 ;
        RECT 28.965 183.510 29.855 183.580 ;
        RECT 30.035 183.895 30.365 184.745 ;
        RECT 28.965 182.785 29.135 183.510 ;
        RECT 29.305 182.955 29.855 183.340 ;
        RECT 30.035 183.130 30.225 183.895 ;
        RECT 30.535 183.815 30.785 184.955 ;
        RECT 30.975 184.315 31.225 184.735 ;
        RECT 31.455 184.485 31.785 184.955 ;
        RECT 32.015 184.315 32.265 184.735 ;
        RECT 30.975 184.145 32.265 184.315 ;
        RECT 32.445 184.315 32.775 184.745 ;
        RECT 32.445 184.145 32.900 184.315 ;
        RECT 30.965 183.645 31.180 183.975 ;
        RECT 30.395 183.315 30.705 183.645 ;
        RECT 30.875 183.315 31.180 183.645 ;
        RECT 31.355 183.315 31.640 183.975 ;
        RECT 31.835 183.315 32.100 183.975 ;
        RECT 32.315 183.315 32.560 183.975 ;
        RECT 30.535 183.145 30.705 183.315 ;
        RECT 32.730 183.145 32.900 184.145 ;
        RECT 28.965 182.615 29.855 182.785 ;
        RECT 30.035 182.620 30.365 183.130 ;
        RECT 30.535 182.975 32.900 183.145 ;
        RECT 30.535 182.405 30.865 182.805 ;
        RECT 31.915 182.635 32.245 182.975 ;
        RECT 32.415 182.405 32.745 182.805 ;
        RECT 33.255 182.585 33.515 184.775 ;
        RECT 33.685 184.225 34.025 184.955 ;
        RECT 34.205 184.045 34.475 184.775 ;
        RECT 33.705 183.825 34.475 184.045 ;
        RECT 34.655 184.065 34.885 184.775 ;
        RECT 35.055 184.245 35.385 184.955 ;
        RECT 35.555 184.065 35.815 184.775 ;
        RECT 34.655 183.825 35.815 184.065 ;
        RECT 36.005 184.235 36.465 184.785 ;
        RECT 36.655 184.235 36.985 184.955 ;
        RECT 33.705 183.155 33.995 183.825 ;
        RECT 34.175 183.335 34.640 183.645 ;
        RECT 34.820 183.335 35.345 183.645 ;
        RECT 33.705 182.955 34.935 183.155 ;
        RECT 33.775 182.405 34.445 182.775 ;
        RECT 34.625 182.585 34.935 182.955 ;
        RECT 35.115 182.695 35.345 183.335 ;
        RECT 35.525 183.315 35.825 183.645 ;
        RECT 35.525 182.405 35.815 183.135 ;
        RECT 36.005 182.865 36.255 184.235 ;
        RECT 37.185 184.065 37.485 184.615 ;
        RECT 37.655 184.285 37.935 184.955 ;
        RECT 36.545 183.895 37.485 184.065 ;
        RECT 36.545 183.645 36.715 183.895 ;
        RECT 37.855 183.645 38.120 184.005 ;
        RECT 38.315 183.985 38.645 184.785 ;
        RECT 38.815 184.155 39.045 184.955 ;
        RECT 39.215 183.985 39.545 184.785 ;
        RECT 38.315 183.815 39.545 183.985 ;
        RECT 39.715 183.815 39.970 184.955 ;
        RECT 40.145 184.105 40.525 184.785 ;
        RECT 41.115 184.105 41.285 184.955 ;
        RECT 41.455 184.275 41.785 184.785 ;
        RECT 41.955 184.445 42.125 184.955 ;
        RECT 42.295 184.275 42.695 184.785 ;
        RECT 41.455 184.105 42.695 184.275 ;
        RECT 36.425 183.315 36.715 183.645 ;
        RECT 36.885 183.395 37.225 183.645 ;
        RECT 37.445 183.395 38.120 183.645 ;
        RECT 38.305 183.315 38.615 183.645 ;
        RECT 36.545 183.225 36.715 183.315 ;
        RECT 36.545 183.035 37.935 183.225 ;
        RECT 36.005 182.575 36.565 182.865 ;
        RECT 36.735 182.405 36.985 182.865 ;
        RECT 37.605 182.675 37.935 183.035 ;
        RECT 38.315 182.915 38.645 183.145 ;
        RECT 38.820 183.085 39.195 183.645 ;
        RECT 39.365 182.915 39.545 183.815 ;
        RECT 39.730 183.065 39.950 183.645 ;
        RECT 40.145 183.145 40.315 184.105 ;
        RECT 40.485 183.765 41.790 183.935 ;
        RECT 42.875 183.855 43.195 184.785 ;
        RECT 43.365 183.865 46.875 184.955 ;
        RECT 47.050 184.530 47.385 184.955 ;
        RECT 47.555 184.350 47.740 184.755 ;
        RECT 40.485 183.315 40.730 183.765 ;
        RECT 40.900 183.395 41.450 183.595 ;
        RECT 41.620 183.565 41.790 183.765 ;
        RECT 42.565 183.685 43.195 183.855 ;
        RECT 41.620 183.395 41.995 183.565 ;
        RECT 42.165 183.145 42.395 183.645 ;
        RECT 40.145 182.975 42.395 183.145 ;
        RECT 38.315 182.575 39.545 182.915 ;
        RECT 39.715 182.405 39.970 182.895 ;
        RECT 40.195 182.405 40.525 182.795 ;
        RECT 40.695 182.655 40.865 182.975 ;
        RECT 42.565 182.805 42.735 183.685 ;
        RECT 41.035 182.405 41.365 182.795 ;
        RECT 41.780 182.635 42.735 182.805 ;
        RECT 42.905 182.405 43.195 183.240 ;
        RECT 43.365 183.175 45.015 183.695 ;
        RECT 45.185 183.345 46.875 183.865 ;
        RECT 47.075 184.175 47.740 184.350 ;
        RECT 47.945 184.175 48.275 184.955 ;
        RECT 43.365 182.405 46.875 183.175 ;
        RECT 47.075 183.145 47.415 184.175 ;
        RECT 48.445 183.985 48.715 184.755 ;
        RECT 47.585 183.815 48.715 183.985 ;
        RECT 48.885 183.865 51.475 184.955 ;
        RECT 47.585 183.315 47.835 183.815 ;
        RECT 47.075 182.975 47.760 183.145 ;
        RECT 48.015 183.065 48.375 183.645 ;
        RECT 47.050 182.405 47.385 182.805 ;
        RECT 47.555 182.575 47.760 182.975 ;
        RECT 48.545 182.905 48.715 183.815 ;
        RECT 47.970 182.405 48.245 182.885 ;
        RECT 48.455 182.575 48.715 182.905 ;
        RECT 48.885 183.175 50.095 183.695 ;
        RECT 50.265 183.345 51.475 183.865 ;
        RECT 52.105 183.790 52.395 184.955 ;
        RECT 48.885 182.405 51.475 183.175 ;
        RECT 52.105 182.405 52.395 183.130 ;
        RECT 52.575 182.585 52.835 184.775 ;
        RECT 53.005 184.225 53.345 184.955 ;
        RECT 53.525 184.045 53.795 184.775 ;
        RECT 53.025 183.825 53.795 184.045 ;
        RECT 53.975 184.065 54.205 184.775 ;
        RECT 54.375 184.245 54.705 184.955 ;
        RECT 54.875 184.065 55.135 184.775 ;
        RECT 53.975 183.825 55.135 184.065 ;
        RECT 55.325 183.865 58.835 184.955 ;
        RECT 53.025 183.155 53.315 183.825 ;
        RECT 53.495 183.335 53.960 183.645 ;
        RECT 54.140 183.335 54.665 183.645 ;
        RECT 53.025 182.955 54.255 183.155 ;
        RECT 53.095 182.405 53.765 182.775 ;
        RECT 53.945 182.585 54.255 182.955 ;
        RECT 54.435 182.695 54.665 183.335 ;
        RECT 54.845 183.315 55.145 183.645 ;
        RECT 55.325 183.175 56.975 183.695 ;
        RECT 57.145 183.345 58.835 183.865 ;
        RECT 59.465 183.985 59.755 184.785 ;
        RECT 59.925 184.155 60.160 184.955 ;
        RECT 60.345 184.615 61.880 184.785 ;
        RECT 60.345 183.985 60.675 184.615 ;
        RECT 59.465 183.815 60.675 183.985 ;
        RECT 59.465 183.315 59.710 183.645 ;
        RECT 54.845 182.405 55.135 183.135 ;
        RECT 55.325 182.405 58.835 183.175 ;
        RECT 59.880 183.145 60.050 183.815 ;
        RECT 60.845 183.645 61.080 184.390 ;
        RECT 60.220 183.315 60.620 183.645 ;
        RECT 60.790 183.315 61.080 183.645 ;
        RECT 61.270 183.645 61.540 184.390 ;
        RECT 61.710 183.985 61.880 184.615 ;
        RECT 62.050 184.155 62.455 184.955 ;
        RECT 61.710 183.815 62.455 183.985 ;
        RECT 61.270 183.315 61.610 183.645 ;
        RECT 61.780 183.315 62.115 183.645 ;
        RECT 62.285 183.315 62.455 183.815 ;
        RECT 62.625 183.390 62.975 184.785 ;
        RECT 59.465 182.575 60.050 183.145 ;
        RECT 60.300 182.975 61.695 183.145 ;
        RECT 60.300 182.630 60.630 182.975 ;
        RECT 60.845 182.405 61.220 182.805 ;
        RECT 61.400 182.630 61.695 182.975 ;
        RECT 61.865 182.405 62.535 183.145 ;
        RECT 62.705 182.575 62.975 183.390 ;
        RECT 63.145 184.235 63.605 184.785 ;
        RECT 63.795 184.235 64.125 184.955 ;
        RECT 63.145 182.865 63.395 184.235 ;
        RECT 64.325 184.065 64.625 184.615 ;
        RECT 64.795 184.285 65.075 184.955 ;
        RECT 63.685 183.895 64.625 184.065 ;
        RECT 63.685 183.645 63.855 183.895 ;
        RECT 64.995 183.645 65.260 184.005 ;
        RECT 65.485 183.815 65.715 184.955 ;
        RECT 65.885 183.805 66.215 184.785 ;
        RECT 66.385 183.815 66.595 184.955 ;
        RECT 67.285 184.445 67.545 184.955 ;
        RECT 63.565 183.315 63.855 183.645 ;
        RECT 64.025 183.395 64.365 183.645 ;
        RECT 64.585 183.395 65.260 183.645 ;
        RECT 65.465 183.395 65.795 183.645 ;
        RECT 63.685 183.225 63.855 183.315 ;
        RECT 63.685 183.035 65.075 183.225 ;
        RECT 63.145 182.575 63.705 182.865 ;
        RECT 63.875 182.405 64.125 182.865 ;
        RECT 64.745 182.675 65.075 183.035 ;
        RECT 65.485 182.405 65.715 183.225 ;
        RECT 65.965 183.205 66.215 183.805 ;
        RECT 67.285 183.395 67.625 184.275 ;
        RECT 67.795 183.565 67.965 184.785 ;
        RECT 68.205 184.450 68.820 184.955 ;
        RECT 68.205 183.915 68.455 184.280 ;
        RECT 68.625 184.275 68.820 184.450 ;
        RECT 68.990 184.445 69.465 184.785 ;
        RECT 69.635 184.410 69.850 184.955 ;
        RECT 68.625 184.085 68.955 184.275 ;
        RECT 69.175 183.915 69.890 184.210 ;
        RECT 70.060 184.085 70.335 184.785 ;
        RECT 68.205 183.745 69.995 183.915 ;
        RECT 67.795 183.315 68.590 183.565 ;
        RECT 67.795 183.225 68.045 183.315 ;
        RECT 65.885 182.575 66.215 183.205 ;
        RECT 66.385 182.405 66.595 183.225 ;
        RECT 67.285 182.405 67.545 183.225 ;
        RECT 67.715 182.805 68.045 183.225 ;
        RECT 68.760 182.890 69.015 183.745 ;
        RECT 68.225 182.625 69.015 182.890 ;
        RECT 69.185 183.045 69.595 183.565 ;
        RECT 69.765 183.315 69.995 183.745 ;
        RECT 70.165 183.055 70.335 184.085 ;
        RECT 70.565 183.895 70.895 184.740 ;
        RECT 71.065 183.945 71.235 184.955 ;
        RECT 71.405 184.225 71.745 184.785 ;
        RECT 71.975 184.455 72.290 184.955 ;
        RECT 72.470 184.485 73.355 184.655 ;
        RECT 70.505 183.815 70.895 183.895 ;
        RECT 71.405 183.850 72.300 184.225 ;
        RECT 70.505 183.765 70.720 183.815 ;
        RECT 70.505 183.185 70.675 183.765 ;
        RECT 71.405 183.645 71.595 183.850 ;
        RECT 72.470 183.645 72.640 184.485 ;
        RECT 73.580 184.455 73.830 184.785 ;
        RECT 70.845 183.315 71.595 183.645 ;
        RECT 71.765 183.315 72.640 183.645 ;
        RECT 70.505 183.145 70.730 183.185 ;
        RECT 71.395 183.145 71.595 183.315 ;
        RECT 70.505 183.060 70.885 183.145 ;
        RECT 69.185 182.625 69.385 183.045 ;
        RECT 69.575 182.405 69.905 182.865 ;
        RECT 70.075 182.575 70.335 183.055 ;
        RECT 70.555 182.625 70.885 183.060 ;
        RECT 71.055 182.405 71.225 183.015 ;
        RECT 71.395 182.620 71.725 183.145 ;
        RECT 71.985 182.405 72.195 182.935 ;
        RECT 72.470 182.855 72.640 183.315 ;
        RECT 72.810 183.355 73.130 184.315 ;
        RECT 73.300 183.565 73.490 184.285 ;
        RECT 73.660 183.385 73.830 184.455 ;
        RECT 74.000 184.155 74.170 184.955 ;
        RECT 74.340 184.510 75.445 184.680 ;
        RECT 74.340 183.895 74.510 184.510 ;
        RECT 75.655 184.360 75.905 184.785 ;
        RECT 76.075 184.495 76.340 184.955 ;
        RECT 74.680 183.975 75.210 184.340 ;
        RECT 75.655 184.230 75.960 184.360 ;
        RECT 74.000 183.805 74.510 183.895 ;
        RECT 74.000 183.635 74.870 183.805 ;
        RECT 74.000 183.565 74.170 183.635 ;
        RECT 74.290 183.385 74.490 183.415 ;
        RECT 72.810 183.025 73.275 183.355 ;
        RECT 73.660 183.085 74.490 183.385 ;
        RECT 73.660 182.855 73.830 183.085 ;
        RECT 72.470 182.685 73.255 182.855 ;
        RECT 73.425 182.685 73.830 182.855 ;
        RECT 74.010 182.405 74.380 182.905 ;
        RECT 74.700 182.855 74.870 183.635 ;
        RECT 75.040 183.275 75.210 183.975 ;
        RECT 75.380 183.445 75.620 184.040 ;
        RECT 75.040 183.055 75.565 183.275 ;
        RECT 75.790 183.125 75.960 184.230 ;
        RECT 75.735 182.995 75.960 183.125 ;
        RECT 76.130 183.035 76.410 183.985 ;
        RECT 75.735 182.855 75.905 182.995 ;
        RECT 74.700 182.685 75.375 182.855 ;
        RECT 75.570 182.685 75.905 182.855 ;
        RECT 76.075 182.405 76.325 182.865 ;
        RECT 76.580 182.665 76.765 184.785 ;
        RECT 76.935 184.455 77.265 184.955 ;
        RECT 77.435 184.285 77.605 184.785 ;
        RECT 76.940 184.115 77.605 184.285 ;
        RECT 76.940 183.125 77.170 184.115 ;
        RECT 77.340 183.295 77.690 183.945 ;
        RECT 77.865 183.790 78.155 184.955 ;
        RECT 78.325 184.520 83.670 184.955 ;
        RECT 83.845 184.520 89.190 184.955 ;
        RECT 76.940 182.955 77.605 183.125 ;
        RECT 76.935 182.405 77.265 182.785 ;
        RECT 77.435 182.665 77.605 182.955 ;
        RECT 77.865 182.405 78.155 183.130 ;
        RECT 79.910 182.950 80.250 183.780 ;
        RECT 81.730 183.270 82.080 184.520 ;
        RECT 85.430 182.950 85.770 183.780 ;
        RECT 87.250 183.270 87.600 184.520 ;
        RECT 89.365 183.865 90.575 184.955 ;
        RECT 89.365 183.155 89.885 183.695 ;
        RECT 90.055 183.325 90.575 183.865 ;
        RECT 90.745 183.865 91.955 184.955 ;
        RECT 112.275 184.710 112.445 185.770 ;
        RECT 113.305 185.710 113.685 186.135 ;
        RECT 114.005 185.840 114.315 186.535 ;
        RECT 114.995 186.530 115.940 186.960 ;
        RECT 114.525 186.250 115.940 186.530 ;
        RECT 116.110 186.595 116.325 187.130 ;
        RECT 116.495 186.780 116.725 187.250 ;
        RECT 116.895 187.210 117.165 187.540 ;
        RECT 117.280 187.075 117.545 187.080 ;
        RECT 117.275 187.070 117.545 187.075 ;
        RECT 117.265 187.065 117.545 187.070 ;
        RECT 117.260 187.060 117.545 187.065 ;
        RECT 117.250 187.055 117.545 187.060 ;
        RECT 117.245 187.045 117.545 187.055 ;
        RECT 117.235 187.035 117.545 187.045 ;
        RECT 117.225 187.020 117.545 187.035 ;
        RECT 116.895 186.720 117.545 187.020 ;
        RECT 116.895 186.595 117.085 186.720 ;
        RECT 116.110 186.310 117.085 186.595 ;
        RECT 117.715 186.480 117.885 187.595 ;
        RECT 118.250 187.145 118.625 187.315 ;
        RECT 118.455 186.945 118.625 187.145 ;
        RECT 118.795 187.115 119.125 187.445 ;
        RECT 119.325 186.945 119.495 187.400 ;
        RECT 118.455 186.775 119.495 186.945 ;
        RECT 119.665 186.605 119.835 187.615 ;
        RECT 120.005 187.470 120.605 187.880 ;
        RECT 120.775 187.810 121.680 187.910 ;
        RECT 122.480 187.810 122.985 187.900 ;
        RECT 120.775 187.640 122.985 187.810 ;
        RECT 123.155 187.780 123.325 188.080 ;
        RECT 123.505 188.080 125.705 188.390 ;
        RECT 123.505 187.950 124.065 188.080 ;
        RECT 125.075 187.950 125.705 188.080 ;
        RECT 125.875 188.305 127.145 188.635 ;
        RECT 120.435 186.990 120.605 187.470 ;
        RECT 120.775 187.300 122.825 187.470 ;
        RECT 120.775 187.200 121.745 187.300 ;
        RECT 122.480 187.200 122.825 187.300 ;
        RECT 123.155 187.330 124.065 187.780 ;
        RECT 124.235 187.740 124.855 187.910 ;
        RECT 125.875 187.775 126.045 188.305 ;
        RECT 127.395 188.205 127.605 188.850 ;
        RECT 127.775 188.365 128.410 188.695 ;
        RECT 121.915 187.030 122.245 187.130 ;
        RECT 120.435 186.725 121.405 186.990 ;
        RECT 117.255 186.310 117.885 186.480 ;
        RECT 118.055 186.435 119.835 186.605 ;
        RECT 114.525 185.845 115.165 186.250 ;
        RECT 116.770 186.080 117.545 186.140 ;
        RECT 112.615 185.535 113.135 185.600 ;
        RECT 113.940 185.535 114.725 185.665 ;
        RECT 112.615 185.360 114.725 185.535 ;
        RECT 114.995 184.710 115.165 185.845 ;
        RECT 115.335 185.800 117.545 186.080 ;
        RECT 117.715 185.705 117.885 186.310 ;
        RECT 118.055 185.875 118.705 186.205 ;
        RECT 117.715 185.535 118.355 185.705 ;
        RECT 117.715 184.710 117.885 185.535 ;
        RECT 118.535 185.365 118.705 185.875 ;
        RECT 118.875 185.695 119.085 186.265 ;
        RECT 119.255 186.225 119.835 186.435 ;
        RECT 120.015 186.710 121.405 186.725 ;
        RECT 121.575 186.860 122.585 187.030 ;
        RECT 123.155 187.010 123.325 187.330 ;
        RECT 124.235 187.180 124.515 187.570 ;
        RECT 124.685 187.290 124.855 187.740 ;
        RECT 125.025 187.460 126.045 187.775 ;
        RECT 126.215 187.505 127.225 187.830 ;
        RECT 125.875 187.335 126.045 187.460 ;
        RECT 120.015 186.395 120.605 186.710 ;
        RECT 119.255 185.900 120.265 186.225 ;
        RECT 118.070 185.035 118.705 185.365 ;
        RECT 118.875 184.880 119.085 185.525 ;
        RECT 120.435 185.425 120.605 186.395 ;
        RECT 119.335 185.095 120.605 185.425 ;
        RECT 120.435 184.710 120.605 185.095 ;
        RECT 120.825 184.885 121.115 186.540 ;
        RECT 121.575 186.475 121.745 186.860 ;
        RECT 121.285 186.305 121.745 186.475 ;
        RECT 121.285 185.205 121.455 186.305 ;
        RECT 121.915 186.285 122.245 186.690 ;
        RECT 122.415 186.460 122.585 186.860 ;
        RECT 122.755 186.820 123.325 187.010 ;
        RECT 123.495 186.990 124.065 187.160 ;
        RECT 124.685 187.120 125.705 187.290 ;
        RECT 122.755 186.630 123.725 186.820 ;
        RECT 122.415 186.290 122.935 186.460 ;
        RECT 123.155 186.400 123.725 186.630 ;
        RECT 121.625 185.405 122.245 186.115 ;
        RECT 122.415 185.590 122.585 186.290 ;
        RECT 123.155 186.120 123.325 186.400 ;
        RECT 123.895 186.230 124.065 186.990 ;
        RECT 124.235 186.950 124.565 186.995 ;
        RECT 124.235 186.750 125.365 186.950 ;
        RECT 124.235 186.300 125.365 186.550 ;
        RECT 122.755 185.790 123.325 186.120 ;
        RECT 123.495 186.000 124.065 186.230 ;
        RECT 125.535 186.110 125.705 187.120 ;
        RECT 122.415 185.420 122.935 185.590 ;
        RECT 121.285 184.885 121.745 185.205 ;
        RECT 121.915 184.885 122.485 185.235 ;
        RECT 123.155 185.220 123.325 185.790 ;
        RECT 123.495 185.510 124.065 185.830 ;
        RECT 124.235 185.680 124.565 186.085 ;
        RECT 124.735 185.860 125.705 186.110 ;
        RECT 125.875 187.005 126.465 187.335 ;
        RECT 126.645 187.295 127.225 187.505 ;
        RECT 127.395 187.465 127.605 188.035 ;
        RECT 127.775 187.855 127.945 188.365 ;
        RECT 128.595 188.195 128.765 189.460 ;
        RECT 129.740 189.370 130.070 189.475 ;
        RECT 130.555 189.460 132.575 189.790 ;
        RECT 132.745 190.670 134.205 190.690 ;
        RECT 132.745 190.430 135.015 190.670 ;
        RECT 132.745 189.760 134.205 190.430 ;
        RECT 135.195 190.340 135.445 190.690 ;
        RECT 135.615 190.350 136.570 190.680 ;
        RECT 134.375 190.170 135.015 190.260 ;
        RECT 135.615 190.170 135.785 190.350 ;
        RECT 134.375 190.000 135.785 190.170 ;
        RECT 136.755 190.025 136.925 190.870 ;
        RECT 137.525 190.825 138.105 191.035 ;
        RECT 139.475 190.950 140.255 191.120 ;
        RECT 137.095 190.500 138.105 190.825 ;
        RECT 138.275 190.295 138.485 190.865 ;
        RECT 138.655 190.475 139.305 190.805 ;
        RECT 134.375 189.930 135.015 190.000 ;
        RECT 132.745 189.490 135.015 189.760 ;
        RECT 132.745 189.480 134.205 189.490 ;
        RECT 135.195 189.480 135.445 189.830 ;
        RECT 136.755 189.820 138.025 190.025 ;
        RECT 135.615 189.695 138.025 189.820 ;
        RECT 135.615 189.490 136.925 189.695 ;
        RECT 131.315 189.310 132.575 189.460 ;
        RECT 128.935 189.200 129.440 189.280 ;
        RECT 130.240 189.200 131.145 189.290 ;
        RECT 128.935 189.020 131.145 189.200 ;
        RECT 128.950 188.365 129.585 188.695 ;
        RECT 128.125 188.025 129.235 188.195 ;
        RECT 127.775 187.525 128.425 187.855 ;
        RECT 126.645 187.125 128.425 187.295 ;
        RECT 125.875 186.260 126.045 187.005 ;
        RECT 124.735 185.510 124.905 185.860 ;
        RECT 125.875 185.850 126.475 186.260 ;
        RECT 126.645 186.115 126.815 187.125 ;
        RECT 126.985 186.785 128.025 186.955 ;
        RECT 126.985 186.330 127.155 186.785 ;
        RECT 127.355 186.285 127.685 186.615 ;
        RECT 127.855 186.585 128.025 186.785 ;
        RECT 127.855 186.415 128.230 186.585 ;
        RECT 128.595 186.135 128.765 188.025 ;
        RECT 129.415 187.855 129.585 188.365 ;
        RECT 129.755 188.205 129.965 188.850 ;
        RECT 131.315 188.635 133.095 189.310 ;
        RECT 130.215 188.305 133.095 188.635 ;
        RECT 131.315 188.100 133.095 188.305 ;
        RECT 133.265 188.225 134.205 189.480 ;
        RECT 134.570 188.595 136.585 188.850 ;
        RECT 134.570 188.490 134.945 188.595 ;
        RECT 135.600 188.510 136.585 188.595 ;
        RECT 136.755 188.800 136.925 189.490 ;
        RECT 138.275 189.480 138.485 190.125 ;
        RECT 138.655 189.965 138.825 190.475 ;
        RECT 139.475 190.305 139.645 190.950 ;
        RECT 139.865 190.625 140.385 190.780 ;
        RECT 140.555 190.740 140.885 191.290 ;
        RECT 142.195 191.130 142.365 191.870 ;
        RECT 141.185 190.960 142.365 191.130 ;
        RECT 139.865 190.570 140.425 190.625 ;
        RECT 141.055 190.615 141.980 190.790 ;
        RECT 141.005 190.570 141.980 190.615 ;
        RECT 139.865 190.460 141.980 190.570 ;
        RECT 139.865 190.450 141.135 190.460 ;
        RECT 140.300 190.400 141.135 190.450 ;
        RECT 139.005 190.135 139.645 190.305 ;
        RECT 138.655 189.635 139.290 189.965 ;
        RECT 139.475 189.605 139.645 190.135 ;
        RECT 142.195 190.280 142.365 190.960 ;
        RECT 142.535 191.720 143.555 191.890 ;
        RECT 143.725 191.780 144.005 192.170 ;
        RECT 144.175 192.065 145.085 192.380 ;
        RECT 147.635 192.065 147.805 193.160 ;
        RECT 144.175 191.930 145.925 192.065 ;
        RECT 144.915 191.805 145.925 191.930 ;
        RECT 146.485 191.805 147.805 192.065 ;
        RECT 142.535 190.710 142.705 191.720 ;
        RECT 143.675 191.550 144.005 191.595 ;
        RECT 142.875 191.350 144.005 191.550 ;
        RECT 144.175 191.590 144.745 191.760 ;
        RECT 142.875 190.900 144.005 191.150 ;
        RECT 144.175 190.830 144.345 191.590 ;
        RECT 144.915 191.420 145.085 191.805 ;
        RECT 144.515 191.205 145.085 191.420 ;
        RECT 145.255 191.460 147.465 191.630 ;
        RECT 145.255 191.375 145.830 191.460 ;
        RECT 146.560 191.375 147.465 191.460 ;
        RECT 145.995 191.205 146.325 191.290 ;
        RECT 147.635 191.205 147.805 191.805 ;
        RECT 144.515 191.000 145.465 191.205 ;
        RECT 144.915 190.875 145.465 191.000 ;
        RECT 145.635 191.035 146.705 191.205 ;
        RECT 142.535 190.460 143.505 190.710 ;
        RECT 142.195 189.950 143.165 190.280 ;
        RECT 143.335 190.110 143.505 190.460 ;
        RECT 143.675 190.280 144.005 190.685 ;
        RECT 144.175 190.600 144.745 190.830 ;
        RECT 144.175 190.110 144.745 190.430 ;
        RECT 139.475 189.365 140.155 189.605 ;
        RECT 137.095 189.055 139.110 189.310 ;
        RECT 137.095 188.970 138.080 189.055 ;
        RECT 138.735 188.950 139.110 189.055 ;
        RECT 138.235 188.800 138.565 188.885 ;
        RECT 135.115 188.340 135.445 188.425 ;
        RECT 136.755 188.390 137.355 188.800 ;
        RECT 137.525 188.535 138.565 188.800 ;
        RECT 139.475 188.685 139.645 189.365 ;
        RECT 140.325 189.355 140.885 189.710 ;
        RECT 141.055 189.195 141.400 189.585 ;
        RECT 142.195 189.200 142.365 189.950 ;
        RECT 143.335 189.940 144.745 190.110 ;
        RECT 144.915 190.230 145.085 190.875 ;
        RECT 145.635 190.660 145.805 191.035 ;
        RECT 145.255 190.490 145.805 190.660 ;
        RECT 145.985 190.400 146.355 190.755 ;
        RECT 146.535 190.660 146.705 191.035 ;
        RECT 146.875 190.875 147.805 191.205 ;
        RECT 146.535 190.490 147.465 190.660 ;
        RECT 147.635 190.230 147.805 190.875 ;
        RECT 142.535 189.370 143.215 189.655 ;
        RECT 141.055 189.185 141.225 189.195 ;
        RECT 139.825 189.015 141.225 189.185 ;
        RECT 139.825 188.905 140.155 189.015 ;
        RECT 138.735 188.675 139.645 188.685 ;
        RECT 136.755 188.340 136.925 188.390 ;
        RECT 133.265 188.100 134.945 188.225 ;
        RECT 128.935 187.525 129.585 187.855 ;
        RECT 129.755 187.465 129.965 188.035 ;
        RECT 130.135 187.505 131.145 187.830 ;
        RECT 130.135 187.295 130.715 187.505 ;
        RECT 131.315 187.460 131.485 188.100 ;
        RECT 134.035 188.055 134.945 188.100 ;
        RECT 135.115 188.075 136.155 188.340 ;
        RECT 131.315 187.335 132.625 187.460 ;
        RECT 128.935 187.125 130.715 187.295 ;
        RECT 129.335 186.785 130.375 186.955 ;
        RECT 129.335 186.585 129.505 186.785 ;
        RECT 129.130 186.415 129.505 186.585 ;
        RECT 129.675 186.285 130.005 186.615 ;
        RECT 130.205 186.330 130.375 186.785 ;
        RECT 126.645 185.850 127.685 186.115 ;
        RECT 127.855 185.965 129.505 186.135 ;
        RECT 130.545 186.115 130.715 187.125 ;
        RECT 130.895 187.130 132.625 187.335 ;
        RECT 130.895 187.005 131.485 187.130 ;
        RECT 132.795 187.120 133.045 187.470 ;
        RECT 134.035 187.460 134.205 188.055 ;
        RECT 134.570 187.605 134.945 187.775 ;
        RECT 133.225 187.190 134.205 187.460 ;
        RECT 134.775 187.405 134.945 187.605 ;
        RECT 135.115 187.575 135.445 187.905 ;
        RECT 135.645 187.405 135.815 187.860 ;
        RECT 134.775 187.235 135.815 187.405 ;
        RECT 131.315 186.260 131.485 187.005 ;
        RECT 133.225 186.950 133.865 187.020 ;
        RECT 132.455 186.780 133.865 186.950 ;
        RECT 132.455 186.600 132.625 186.780 ;
        RECT 133.225 186.690 133.865 186.780 ;
        RECT 131.670 186.270 132.625 186.600 ;
        RECT 132.795 186.260 133.045 186.610 ;
        RECT 134.035 186.520 134.205 187.190 ;
        RECT 135.985 187.065 136.155 188.075 ;
        RECT 136.325 187.930 136.925 188.340 ;
        RECT 136.755 187.645 136.925 187.930 ;
        RECT 136.755 187.315 137.345 187.645 ;
        RECT 137.525 187.525 137.695 188.535 ;
        RECT 138.735 188.515 140.155 188.675 ;
        RECT 140.325 188.580 140.885 188.845 ;
        RECT 139.475 188.460 140.155 188.515 ;
        RECT 137.865 187.865 138.035 188.320 ;
        RECT 138.235 188.035 138.565 188.365 ;
        RECT 138.735 188.065 139.110 188.235 ;
        RECT 138.735 187.865 138.905 188.065 ;
        RECT 137.865 187.695 138.905 187.865 ;
        RECT 137.525 187.355 139.305 187.525 ;
        RECT 136.755 187.185 136.925 187.315 ;
        RECT 134.375 186.895 136.155 187.065 ;
        RECT 133.225 186.280 134.205 186.520 ;
        RECT 134.375 186.335 135.025 186.665 ;
        RECT 125.875 185.680 126.045 185.850 ;
        RECT 127.355 185.765 127.685 185.850 ;
        RECT 123.495 185.340 124.905 185.510 ;
        RECT 125.075 185.350 126.045 185.680 ;
        RECT 122.655 184.890 123.325 185.220 ;
        RECT 123.155 184.710 123.325 184.890 ;
        RECT 125.875 184.710 126.045 185.350 ;
        RECT 126.215 185.595 127.200 185.680 ;
        RECT 127.855 185.595 128.230 185.700 ;
        RECT 126.215 185.570 128.230 185.595 ;
        RECT 126.215 185.400 128.255 185.570 ;
        RECT 126.215 185.340 128.230 185.400 ;
        RECT 128.595 184.710 128.765 185.965 ;
        RECT 129.675 185.850 130.715 186.115 ;
        RECT 130.885 185.850 131.485 186.260 ;
        RECT 134.035 186.165 134.205 186.280 ;
        RECT 129.675 185.765 130.005 185.850 ;
        RECT 129.130 185.595 129.505 185.700 ;
        RECT 130.160 185.595 131.145 185.680 ;
        RECT 129.130 185.340 131.145 185.595 ;
        RECT 131.315 185.650 131.485 185.850 ;
        RECT 131.655 185.920 133.865 186.090 ;
        RECT 131.655 185.820 132.560 185.920 ;
        RECT 133.360 185.830 133.865 185.920 ;
        RECT 134.035 185.995 134.675 186.165 ;
        RECT 131.315 185.320 132.245 185.650 ;
        RECT 132.730 185.635 133.060 185.750 ;
        RECT 134.035 185.650 134.205 185.995 ;
        RECT 134.855 185.825 135.025 186.335 ;
        RECT 135.195 186.155 135.405 186.725 ;
        RECT 135.575 186.685 136.155 186.895 ;
        RECT 136.335 186.855 136.925 187.185 ;
        RECT 137.525 187.145 138.105 187.355 ;
        RECT 135.575 186.360 136.585 186.685 ;
        RECT 136.755 186.345 136.925 186.855 ;
        RECT 137.095 186.820 138.105 187.145 ;
        RECT 138.275 186.615 138.485 187.185 ;
        RECT 138.655 186.795 139.305 187.125 ;
        RECT 139.475 187.030 139.645 188.460 ;
        RECT 141.055 188.330 141.225 189.015 ;
        RECT 142.195 188.930 142.825 189.200 ;
        RECT 142.195 188.710 142.365 188.930 ;
        RECT 141.395 188.380 142.365 188.710 ;
        RECT 142.995 188.910 143.215 189.370 ;
        RECT 143.385 189.080 143.945 189.770 ;
        RECT 144.915 189.710 146.375 190.230 ;
        RECT 144.115 189.370 144.745 189.655 ;
        RECT 144.115 188.910 144.285 189.370 ;
        RECT 144.915 189.200 145.835 189.710 ;
        RECT 146.545 189.540 147.805 190.230 ;
        RECT 144.455 189.020 145.835 189.200 ;
        RECT 146.005 189.020 147.805 189.540 ;
        RECT 144.455 188.930 145.085 189.020 ;
        RECT 142.995 188.700 144.285 188.910 ;
        RECT 139.815 187.990 140.385 188.290 ;
        RECT 140.555 188.160 141.225 188.330 ;
        RECT 141.405 187.990 142.025 188.210 ;
        RECT 139.815 187.675 142.025 187.990 ;
        RECT 139.815 187.210 140.365 187.380 ;
        RECT 136.755 186.015 138.025 186.345 ;
        RECT 132.415 185.465 133.485 185.635 ;
        RECT 131.315 184.710 131.485 185.320 ;
        RECT 132.415 185.140 132.585 185.465 ;
        RECT 131.655 184.970 132.585 185.140 ;
        RECT 132.765 184.900 133.135 185.230 ;
        RECT 133.315 185.140 133.485 185.465 ;
        RECT 133.655 185.320 134.205 185.650 ;
        RECT 134.390 185.495 135.025 185.825 ;
        RECT 135.195 185.340 135.405 185.985 ;
        RECT 136.755 185.885 136.925 186.015 ;
        RECT 135.655 185.555 136.925 185.885 ;
        RECT 138.275 185.800 138.485 186.445 ;
        RECT 138.655 186.285 138.825 186.795 ;
        RECT 139.475 186.700 140.025 187.030 ;
        RECT 140.195 186.885 140.365 187.210 ;
        RECT 140.545 187.120 140.915 187.450 ;
        RECT 141.095 187.210 142.025 187.380 ;
        RECT 141.095 186.885 141.265 187.210 ;
        RECT 142.195 187.140 142.365 188.380 ;
        RECT 142.535 188.130 144.745 188.530 ;
        RECT 144.915 188.410 145.085 188.930 ;
        RECT 145.255 188.680 147.465 188.850 ;
        RECT 145.255 188.590 145.760 188.680 ;
        RECT 146.560 188.580 147.465 188.680 ;
        RECT 142.535 187.660 143.215 187.940 ;
        RECT 142.995 187.265 143.215 187.660 ;
        RECT 143.385 187.435 143.945 188.130 ;
        RECT 144.915 188.080 145.465 188.410 ;
        RECT 146.060 188.395 146.390 188.510 ;
        RECT 147.635 188.410 147.805 189.020 ;
        RECT 145.635 188.225 146.705 188.395 ;
        RECT 144.115 187.660 144.745 187.940 ;
        RECT 144.115 187.265 144.285 187.660 ;
        RECT 142.195 187.030 142.825 187.140 ;
        RECT 140.195 186.715 141.265 186.885 ;
        RECT 141.435 186.815 142.825 187.030 ;
        RECT 142.995 186.815 144.285 187.265 ;
        RECT 144.915 187.140 145.085 188.080 ;
        RECT 145.635 187.900 145.805 188.225 ;
        RECT 145.255 187.730 145.805 187.900 ;
        RECT 145.985 187.660 146.355 187.990 ;
        RECT 146.535 187.900 146.705 188.225 ;
        RECT 146.875 188.080 147.805 188.410 ;
        RECT 146.535 187.730 147.465 187.900 ;
        RECT 145.255 187.300 147.465 187.470 ;
        RECT 145.255 187.210 145.760 187.300 ;
        RECT 146.560 187.200 147.465 187.300 ;
        RECT 144.455 187.030 145.085 187.140 ;
        RECT 144.455 186.815 145.465 187.030 ;
        RECT 146.060 187.015 146.390 187.130 ;
        RECT 147.635 187.030 147.805 188.080 ;
        RECT 139.475 186.625 139.645 186.700 ;
        RECT 139.005 186.455 139.645 186.625 ;
        RECT 140.620 186.600 140.950 186.715 ;
        RECT 141.435 186.700 142.365 186.815 ;
        RECT 143.675 186.710 144.005 186.815 ;
        RECT 138.655 185.955 139.290 186.285 ;
        RECT 133.315 184.970 133.865 185.140 ;
        RECT 134.035 184.710 134.205 185.320 ;
        RECT 136.755 184.710 136.925 185.555 ;
        RECT 139.475 185.650 139.645 186.455 ;
        RECT 139.815 186.430 140.320 186.520 ;
        RECT 141.120 186.430 142.025 186.530 ;
        RECT 139.815 186.260 142.025 186.430 ;
        RECT 139.815 185.910 142.025 186.090 ;
        RECT 139.815 185.830 140.320 185.910 ;
        RECT 141.120 185.820 142.025 185.910 ;
        RECT 139.475 185.320 140.025 185.650 ;
        RECT 140.620 185.635 140.950 185.740 ;
        RECT 142.195 185.650 142.365 186.700 ;
        RECT 144.915 186.700 145.465 186.815 ;
        RECT 145.635 186.845 146.705 187.015 ;
        RECT 142.535 186.540 143.505 186.645 ;
        RECT 144.175 186.540 144.745 186.645 ;
        RECT 142.535 186.260 144.745 186.540 ;
        RECT 142.535 185.910 144.745 186.090 ;
        RECT 142.535 185.820 143.440 185.910 ;
        RECT 144.240 185.830 144.745 185.910 ;
        RECT 140.195 185.465 141.265 185.635 ;
        RECT 139.475 184.710 139.645 185.320 ;
        RECT 140.195 185.140 140.365 185.465 ;
        RECT 139.815 184.970 140.365 185.140 ;
        RECT 140.545 184.900 140.915 185.240 ;
        RECT 141.095 185.140 141.265 185.465 ;
        RECT 141.435 185.320 143.125 185.650 ;
        RECT 143.610 185.635 143.940 185.740 ;
        RECT 144.915 185.650 145.085 186.700 ;
        RECT 145.635 186.520 145.805 186.845 ;
        RECT 145.255 186.350 145.805 186.520 ;
        RECT 145.985 186.280 146.355 186.610 ;
        RECT 146.535 186.520 146.705 186.845 ;
        RECT 146.875 186.700 147.805 187.030 ;
        RECT 146.535 186.350 147.465 186.520 ;
        RECT 145.255 185.910 147.465 186.090 ;
        RECT 145.255 185.830 145.760 185.910 ;
        RECT 146.560 185.820 147.465 185.910 ;
        RECT 143.295 185.465 144.365 185.635 ;
        RECT 141.095 184.960 142.025 185.140 ;
        RECT 142.195 184.710 142.365 185.320 ;
        RECT 143.295 185.140 143.465 185.465 ;
        RECT 142.535 184.960 143.465 185.140 ;
        RECT 143.645 184.900 144.015 185.240 ;
        RECT 144.195 185.140 144.365 185.465 ;
        RECT 144.535 185.320 145.465 185.650 ;
        RECT 146.060 185.635 146.390 185.740 ;
        RECT 147.635 185.650 147.805 186.700 ;
        RECT 145.635 185.465 146.705 185.635 ;
        RECT 144.195 184.970 144.745 185.140 ;
        RECT 144.915 184.710 145.085 185.320 ;
        RECT 145.635 185.140 145.805 185.465 ;
        RECT 145.255 184.970 145.805 185.140 ;
        RECT 145.985 184.900 146.355 185.240 ;
        RECT 146.535 185.140 146.705 185.465 ;
        RECT 146.875 185.320 147.805 185.650 ;
        RECT 146.535 184.960 147.465 185.140 ;
        RECT 147.635 184.710 147.805 185.320 ;
        RECT 112.275 184.020 113.195 184.710 ;
        RECT 113.365 184.190 116.795 184.710 ;
        RECT 90.745 183.325 91.265 183.865 ;
        RECT 91.435 183.155 91.955 183.695 ;
        RECT 112.275 183.500 113.735 184.020 ;
        RECT 113.905 183.500 116.255 184.190 ;
        RECT 116.965 184.020 118.635 184.710 ;
        RECT 118.805 184.190 122.235 184.710 ;
        RECT 116.425 183.500 119.175 184.020 ;
        RECT 119.345 183.500 121.695 184.190 ;
        RECT 122.405 184.020 124.075 184.710 ;
        RECT 124.245 184.190 127.675 184.710 ;
        RECT 121.865 183.500 124.615 184.020 ;
        RECT 124.785 183.500 127.135 184.190 ;
        RECT 127.845 184.020 129.515 184.710 ;
        RECT 129.685 184.190 133.115 184.710 ;
        RECT 127.305 183.500 130.055 184.020 ;
        RECT 130.225 183.500 132.575 184.190 ;
        RECT 133.285 184.020 134.955 184.710 ;
        RECT 135.125 184.190 138.555 184.710 ;
        RECT 132.745 183.500 135.495 184.020 ;
        RECT 135.665 183.500 138.015 184.190 ;
        RECT 138.725 184.020 140.395 184.710 ;
        RECT 140.565 184.190 143.995 184.710 ;
        RECT 138.185 183.500 140.935 184.020 ;
        RECT 141.105 183.500 143.455 184.190 ;
        RECT 144.165 184.020 145.835 184.710 ;
        RECT 146.005 184.190 147.805 184.710 ;
        RECT 143.625 183.500 146.375 184.020 ;
        RECT 146.545 183.500 147.805 184.190 ;
        RECT 112.275 183.415 112.445 183.500 ;
        RECT 114.995 183.415 115.165 183.500 ;
        RECT 117.715 183.415 117.885 183.500 ;
        RECT 120.435 183.415 120.605 183.500 ;
        RECT 123.155 183.415 123.325 183.500 ;
        RECT 125.875 183.415 126.045 183.500 ;
        RECT 128.595 183.415 128.765 183.500 ;
        RECT 131.315 183.415 131.485 183.500 ;
        RECT 134.035 183.415 134.205 183.500 ;
        RECT 136.755 183.415 136.925 183.500 ;
        RECT 139.475 183.415 139.645 183.500 ;
        RECT 142.195 183.415 142.365 183.500 ;
        RECT 144.915 183.415 145.085 183.500 ;
        RECT 147.635 183.415 147.805 183.500 ;
        RECT 78.325 182.405 83.670 182.950 ;
        RECT 83.845 182.405 89.190 182.950 ;
        RECT 89.365 182.405 90.575 183.155 ;
        RECT 90.745 182.405 91.955 183.155 ;
        RECT 13.380 182.235 92.040 182.405 ;
        RECT 13.465 181.485 14.675 182.235 ;
        RECT 14.845 181.690 20.190 182.235 ;
        RECT 13.465 180.945 13.985 181.485 ;
        RECT 14.155 180.775 14.675 181.315 ;
        RECT 16.430 180.860 16.770 181.690 ;
        RECT 20.365 181.465 22.035 182.235 ;
        RECT 22.240 181.495 22.855 182.065 ;
        RECT 23.025 181.725 23.240 182.235 ;
        RECT 23.470 181.725 23.750 182.055 ;
        RECT 23.930 181.725 24.170 182.235 ;
        RECT 13.465 179.685 14.675 180.775 ;
        RECT 18.250 180.120 18.600 181.370 ;
        RECT 20.365 180.945 21.115 181.465 ;
        RECT 21.285 180.775 22.035 181.295 ;
        RECT 14.845 179.685 20.190 180.120 ;
        RECT 20.365 179.685 22.035 180.775 ;
        RECT 22.240 180.475 22.555 181.495 ;
        RECT 22.725 180.825 22.895 181.325 ;
        RECT 23.145 180.995 23.410 181.555 ;
        RECT 23.580 180.825 23.750 181.725 ;
        RECT 24.505 181.690 29.850 182.235 ;
        RECT 23.920 180.995 24.275 181.555 ;
        RECT 26.090 180.860 26.430 181.690 ;
        RECT 30.485 181.515 30.825 182.025 ;
        RECT 22.725 180.655 24.150 180.825 ;
        RECT 22.240 179.855 22.775 180.475 ;
        RECT 22.945 179.685 23.275 180.485 ;
        RECT 23.760 180.480 24.150 180.655 ;
        RECT 27.910 180.120 28.260 181.370 ;
        RECT 24.505 179.685 29.850 180.120 ;
        RECT 30.485 180.115 30.745 181.515 ;
        RECT 30.995 181.435 31.265 182.235 ;
        RECT 30.920 180.995 31.250 181.245 ;
        RECT 31.445 180.995 31.725 181.965 ;
        RECT 31.905 180.995 32.205 181.965 ;
        RECT 32.385 180.995 32.735 181.960 ;
        RECT 32.955 181.735 33.450 182.065 ;
        RECT 30.935 180.825 31.250 180.995 ;
        RECT 32.955 180.825 33.125 181.735 ;
        RECT 30.935 180.655 33.125 180.825 ;
        RECT 30.485 179.855 30.825 180.115 ;
        RECT 30.995 179.685 31.325 180.485 ;
        RECT 31.790 179.855 32.040 180.655 ;
        RECT 32.225 179.685 32.555 180.405 ;
        RECT 32.775 179.855 33.025 180.655 ;
        RECT 33.295 180.245 33.535 181.555 ;
        RECT 34.165 181.495 34.605 182.055 ;
        RECT 34.775 181.495 35.225 182.235 ;
        RECT 35.395 181.665 35.565 182.065 ;
        RECT 35.735 181.835 36.155 182.235 ;
        RECT 36.325 181.665 36.555 182.065 ;
        RECT 35.395 181.495 36.555 181.665 ;
        RECT 36.725 181.495 37.215 182.065 ;
        RECT 34.165 180.485 34.475 181.495 ;
        RECT 34.645 180.875 34.815 181.325 ;
        RECT 34.985 181.045 35.375 181.325 ;
        RECT 35.560 180.995 35.805 181.325 ;
        RECT 34.645 180.705 35.435 180.875 ;
        RECT 33.195 179.685 33.530 180.065 ;
        RECT 34.165 179.855 34.605 180.485 ;
        RECT 34.780 179.685 35.095 180.535 ;
        RECT 35.265 180.025 35.435 180.705 ;
        RECT 35.605 180.195 35.805 180.995 ;
        RECT 36.005 180.195 36.255 181.325 ;
        RECT 36.470 180.995 36.875 181.325 ;
        RECT 37.045 180.825 37.215 181.495 ;
        RECT 37.385 181.465 39.055 182.235 ;
        RECT 39.225 181.510 39.515 182.235 ;
        RECT 40.605 181.495 41.070 182.040 ;
        RECT 37.385 180.945 38.135 181.465 ;
        RECT 36.445 180.655 37.215 180.825 ;
        RECT 38.305 180.775 39.055 181.295 ;
        RECT 36.445 180.025 36.695 180.655 ;
        RECT 35.265 179.855 36.695 180.025 ;
        RECT 36.875 179.685 37.205 180.485 ;
        RECT 37.385 179.685 39.055 180.775 ;
        RECT 39.225 179.685 39.515 180.850 ;
        RECT 40.605 180.535 40.775 181.495 ;
        RECT 41.575 181.415 41.745 182.235 ;
        RECT 41.915 181.585 42.245 182.065 ;
        RECT 42.415 181.845 42.765 182.235 ;
        RECT 42.935 181.665 43.165 182.065 ;
        RECT 42.655 181.585 43.165 181.665 ;
        RECT 41.915 181.495 43.165 181.585 ;
        RECT 43.335 181.495 43.655 181.975 ;
        RECT 41.915 181.415 42.825 181.495 ;
        RECT 40.945 180.875 41.190 181.325 ;
        RECT 41.450 181.045 42.145 181.245 ;
        RECT 42.315 181.075 42.915 181.245 ;
        RECT 42.315 180.875 42.485 181.075 ;
        RECT 43.145 180.905 43.315 181.325 ;
        RECT 40.945 180.705 42.485 180.875 ;
        RECT 42.655 180.735 43.315 180.905 ;
        RECT 42.655 180.535 42.825 180.735 ;
        RECT 43.485 180.565 43.655 181.495 ;
        RECT 43.825 181.435 44.520 182.065 ;
        RECT 44.725 181.435 45.035 182.235 ;
        RECT 45.370 181.725 45.610 182.235 ;
        RECT 45.790 181.725 46.070 182.055 ;
        RECT 46.300 181.725 46.515 182.235 ;
        RECT 44.345 181.385 44.520 181.435 ;
        RECT 43.845 180.995 44.180 181.245 ;
        RECT 44.350 180.835 44.520 181.385 ;
        RECT 44.690 180.995 45.025 181.265 ;
        RECT 45.265 180.995 45.620 181.555 ;
        RECT 40.605 180.365 42.825 180.535 ;
        RECT 42.995 180.365 43.655 180.565 ;
        RECT 40.605 179.685 40.905 180.195 ;
        RECT 41.075 179.855 41.405 180.365 ;
        RECT 42.995 180.195 43.165 180.365 ;
        RECT 41.575 179.685 42.205 180.195 ;
        RECT 42.785 180.025 43.165 180.195 ;
        RECT 43.335 179.685 43.635 180.195 ;
        RECT 43.825 179.685 44.085 180.825 ;
        RECT 44.255 179.855 44.585 180.835 ;
        RECT 45.790 180.825 45.960 181.725 ;
        RECT 46.130 180.995 46.395 181.555 ;
        RECT 46.685 181.495 47.300 182.065 ;
        RECT 47.590 181.665 47.765 182.065 ;
        RECT 47.935 181.855 48.265 182.235 ;
        RECT 48.510 181.735 48.740 182.065 ;
        RECT 47.590 181.495 48.220 181.665 ;
        RECT 46.645 180.825 46.815 181.325 ;
        RECT 44.755 179.685 45.035 180.825 ;
        RECT 45.390 180.655 46.815 180.825 ;
        RECT 45.390 180.480 45.780 180.655 ;
        RECT 46.265 179.685 46.595 180.485 ;
        RECT 46.985 180.475 47.300 181.495 ;
        RECT 48.050 181.325 48.220 181.495 ;
        RECT 47.505 180.645 47.870 181.325 ;
        RECT 48.050 180.995 48.400 181.325 ;
        RECT 48.050 180.475 48.220 180.995 ;
        RECT 46.765 179.855 47.300 180.475 ;
        RECT 47.590 180.305 48.220 180.475 ;
        RECT 48.570 180.445 48.740 181.735 ;
        RECT 48.940 180.625 49.220 181.900 ;
        RECT 49.445 181.895 49.715 181.900 ;
        RECT 49.405 181.725 49.715 181.895 ;
        RECT 50.175 181.855 50.505 182.235 ;
        RECT 50.675 181.980 51.010 182.025 ;
        RECT 49.445 180.625 49.715 181.725 ;
        RECT 49.905 180.625 50.245 181.655 ;
        RECT 50.675 181.515 51.015 181.980 ;
        RECT 51.190 181.705 51.480 182.055 ;
        RECT 51.675 181.875 52.005 182.235 ;
        RECT 52.175 181.705 52.405 182.010 ;
        RECT 51.190 181.535 52.405 181.705 ;
        RECT 52.595 181.895 52.765 181.930 ;
        RECT 52.595 181.725 52.795 181.895 ;
        RECT 50.415 180.995 50.675 181.325 ;
        RECT 50.415 180.445 50.585 180.995 ;
        RECT 50.845 180.825 51.015 181.515 ;
        RECT 52.595 181.365 52.765 181.725 ;
        RECT 53.165 181.640 53.485 182.065 ;
        RECT 53.655 181.810 53.985 182.235 ;
        RECT 54.155 181.815 55.245 182.065 ;
        RECT 55.435 181.815 56.525 182.065 ;
        RECT 54.155 181.640 54.325 181.815 ;
        RECT 53.165 181.470 54.325 181.640 ;
        RECT 54.495 181.475 56.185 181.645 ;
        RECT 56.355 181.640 56.525 181.815 ;
        RECT 56.695 181.810 57.025 182.235 ;
        RECT 57.195 181.640 57.445 182.065 ;
        RECT 51.250 181.215 51.510 181.325 ;
        RECT 51.245 181.045 51.510 181.215 ;
        RECT 51.250 180.995 51.510 181.045 ;
        RECT 51.690 180.995 52.075 181.325 ;
        RECT 52.245 181.195 52.765 181.365 ;
        RECT 53.040 181.215 54.150 181.245 ;
        RECT 47.590 179.855 47.765 180.305 ;
        RECT 48.570 180.275 50.585 180.445 ;
        RECT 47.935 179.685 48.265 180.125 ;
        RECT 48.570 179.855 48.740 180.275 ;
        RECT 48.975 179.685 49.645 180.095 ;
        RECT 49.860 179.855 50.030 180.275 ;
        RECT 50.230 179.685 50.560 180.095 ;
        RECT 50.755 179.855 51.015 180.825 ;
        RECT 51.190 179.685 51.510 180.825 ;
        RECT 51.690 179.945 51.885 180.995 ;
        RECT 52.245 180.815 52.415 181.195 ;
        RECT 53.040 181.045 54.175 181.215 ;
        RECT 54.440 181.045 55.095 181.245 ;
        RECT 52.065 180.535 52.415 180.815 ;
        RECT 52.605 180.665 52.850 181.025 ;
        RECT 55.380 180.835 55.670 181.475 ;
        RECT 56.355 181.470 57.445 181.640 ;
        RECT 57.625 181.650 57.935 182.065 ;
        RECT 58.130 181.855 58.460 182.235 ;
        RECT 58.630 181.895 60.035 182.065 ;
        RECT 58.630 181.665 58.800 181.895 ;
        RECT 55.840 181.045 56.470 181.245 ;
        RECT 56.760 181.215 57.390 181.245 ;
        RECT 56.760 181.045 57.395 181.215 ;
        RECT 53.235 180.665 55.165 180.835 ;
        RECT 52.065 179.855 52.395 180.535 ;
        RECT 52.595 179.685 52.850 180.485 ;
        RECT 53.235 179.855 53.565 180.665 ;
        RECT 53.735 179.685 53.905 180.495 ;
        RECT 54.075 179.855 54.405 180.665 ;
        RECT 54.575 179.685 54.745 180.495 ;
        RECT 54.915 180.025 55.165 180.665 ;
        RECT 55.380 180.665 57.445 180.835 ;
        RECT 55.380 180.195 55.765 180.665 ;
        RECT 55.935 180.025 56.105 180.495 ;
        RECT 56.275 180.195 56.605 180.665 ;
        RECT 56.775 180.025 57.025 180.495 ;
        RECT 54.915 179.855 57.025 180.025 ;
        RECT 57.195 179.855 57.445 180.665 ;
        RECT 57.625 180.535 57.795 181.650 ;
        RECT 58.105 181.495 58.800 181.665 ;
        RECT 59.865 181.665 60.035 181.895 ;
        RECT 60.305 181.835 60.635 182.235 ;
        RECT 60.875 181.665 61.045 182.065 ;
        RECT 58.105 181.325 58.275 181.495 ;
        RECT 57.965 180.995 58.275 181.325 ;
        RECT 58.445 180.995 58.780 181.325 ;
        RECT 59.050 180.995 59.245 181.570 ;
        RECT 59.505 181.325 59.695 181.555 ;
        RECT 59.865 181.495 61.045 181.665 ;
        RECT 61.765 181.415 62.025 182.235 ;
        RECT 62.195 181.415 62.525 181.835 ;
        RECT 62.705 181.665 62.965 182.065 ;
        RECT 63.135 181.835 63.465 182.235 ;
        RECT 63.635 181.665 63.805 182.015 ;
        RECT 63.975 181.835 64.350 182.235 ;
        RECT 62.705 181.495 64.370 181.665 ;
        RECT 64.540 181.560 64.815 181.905 ;
        RECT 62.275 181.325 62.525 181.415 ;
        RECT 64.200 181.325 64.370 181.495 ;
        RECT 59.505 180.995 59.850 181.325 ;
        RECT 60.160 180.995 60.635 181.325 ;
        RECT 60.890 180.995 61.075 181.325 ;
        RECT 61.770 180.995 62.105 181.245 ;
        RECT 62.275 180.995 62.990 181.325 ;
        RECT 63.205 180.995 64.030 181.325 ;
        RECT 64.200 180.995 64.475 181.325 ;
        RECT 58.105 180.825 58.275 180.995 ;
        RECT 58.105 180.655 61.045 180.825 ;
        RECT 57.625 179.895 57.965 180.535 ;
        RECT 58.555 180.315 60.115 180.485 ;
        RECT 58.135 179.685 58.380 180.145 ;
        RECT 58.555 179.855 58.805 180.315 ;
        RECT 58.995 179.685 59.665 180.065 ;
        RECT 59.865 179.855 60.115 180.315 ;
        RECT 60.875 179.855 61.045 180.655 ;
        RECT 61.765 179.685 62.025 180.825 ;
        RECT 62.275 180.435 62.445 180.995 ;
        RECT 62.705 180.535 63.035 180.825 ;
        RECT 63.205 180.705 63.450 180.995 ;
        RECT 64.200 180.825 64.370 180.995 ;
        RECT 64.645 180.825 64.815 181.560 ;
        RECT 64.985 181.510 65.275 182.235 ;
        RECT 65.445 181.585 65.705 182.065 ;
        RECT 65.875 181.775 66.205 182.235 ;
        RECT 66.395 181.595 66.595 182.015 ;
        RECT 63.710 180.655 64.370 180.825 ;
        RECT 63.710 180.535 63.880 180.655 ;
        RECT 62.705 180.365 63.880 180.535 ;
        RECT 62.265 179.865 63.880 180.195 ;
        RECT 64.050 179.685 64.330 180.485 ;
        RECT 64.540 179.855 64.815 180.825 ;
        RECT 64.985 179.685 65.275 180.850 ;
        RECT 65.445 180.555 65.615 181.585 ;
        RECT 65.785 180.895 66.015 181.325 ;
        RECT 66.185 181.075 66.595 181.595 ;
        RECT 66.765 181.750 67.555 182.015 ;
        RECT 66.765 180.895 67.020 181.750 ;
        RECT 67.735 181.415 68.065 181.835 ;
        RECT 68.235 181.415 68.495 182.235 ;
        RECT 68.665 181.855 69.555 182.025 ;
        RECT 67.735 181.325 67.985 181.415 ;
        RECT 67.190 181.075 67.985 181.325 ;
        RECT 68.665 181.300 69.215 181.685 ;
        RECT 65.785 180.725 67.575 180.895 ;
        RECT 65.445 179.855 65.720 180.555 ;
        RECT 65.890 180.430 66.605 180.725 ;
        RECT 66.825 180.365 67.155 180.555 ;
        RECT 65.930 179.685 66.145 180.230 ;
        RECT 66.315 179.855 66.790 180.195 ;
        RECT 66.960 180.190 67.155 180.365 ;
        RECT 67.325 180.360 67.575 180.725 ;
        RECT 66.960 179.685 67.575 180.190 ;
        RECT 67.815 179.855 67.985 181.075 ;
        RECT 68.155 180.365 68.495 181.245 ;
        RECT 69.385 181.130 69.555 181.855 ;
        RECT 68.665 181.060 69.555 181.130 ;
        RECT 69.725 181.530 69.945 182.015 ;
        RECT 70.115 181.695 70.365 182.235 ;
        RECT 70.535 181.585 70.795 182.065 ;
        RECT 69.725 181.105 70.055 181.530 ;
        RECT 68.665 181.035 69.560 181.060 ;
        RECT 68.665 181.020 69.570 181.035 ;
        RECT 68.665 181.005 69.575 181.020 ;
        RECT 68.665 181.000 69.585 181.005 ;
        RECT 68.665 180.990 69.590 181.000 ;
        RECT 68.665 180.980 69.595 180.990 ;
        RECT 68.665 180.975 69.605 180.980 ;
        RECT 68.665 180.965 69.615 180.975 ;
        RECT 68.665 180.960 69.625 180.965 ;
        RECT 68.665 180.510 68.925 180.960 ;
        RECT 69.290 180.955 69.625 180.960 ;
        RECT 69.290 180.950 69.640 180.955 ;
        RECT 69.290 180.940 69.655 180.950 ;
        RECT 69.290 180.935 69.680 180.940 ;
        RECT 70.225 180.935 70.455 181.330 ;
        RECT 69.290 180.930 70.455 180.935 ;
        RECT 69.320 180.895 70.455 180.930 ;
        RECT 69.355 180.870 70.455 180.895 ;
        RECT 69.385 180.840 70.455 180.870 ;
        RECT 69.405 180.810 70.455 180.840 ;
        RECT 69.425 180.780 70.455 180.810 ;
        RECT 69.495 180.770 70.455 180.780 ;
        RECT 69.520 180.760 70.455 180.770 ;
        RECT 69.540 180.745 70.455 180.760 ;
        RECT 69.560 180.730 70.455 180.745 ;
        RECT 69.565 180.720 70.350 180.730 ;
        RECT 69.580 180.685 70.350 180.720 ;
        RECT 69.095 180.365 69.425 180.610 ;
        RECT 69.595 180.435 70.350 180.685 ;
        RECT 70.625 180.555 70.795 181.585 ;
        RECT 71.055 181.685 71.225 181.975 ;
        RECT 71.395 181.855 71.725 182.235 ;
        RECT 71.055 181.515 71.720 181.685 ;
        RECT 70.970 180.695 71.320 181.345 ;
        RECT 69.095 180.340 69.280 180.365 ;
        RECT 68.665 180.240 69.280 180.340 ;
        RECT 68.235 179.685 68.495 180.195 ;
        RECT 68.665 179.685 69.270 180.240 ;
        RECT 69.445 179.855 69.925 180.195 ;
        RECT 70.095 179.685 70.350 180.230 ;
        RECT 70.520 179.855 70.795 180.555 ;
        RECT 71.490 180.525 71.720 181.515 ;
        RECT 71.055 180.355 71.720 180.525 ;
        RECT 71.055 179.855 71.225 180.355 ;
        RECT 71.395 179.685 71.725 180.185 ;
        RECT 71.895 179.855 72.080 181.975 ;
        RECT 72.335 181.775 72.585 182.235 ;
        RECT 72.755 181.785 73.090 181.955 ;
        RECT 73.285 181.785 73.960 181.955 ;
        RECT 72.755 181.645 72.925 181.785 ;
        RECT 72.250 180.655 72.530 181.605 ;
        RECT 72.700 181.515 72.925 181.645 ;
        RECT 72.700 180.410 72.870 181.515 ;
        RECT 73.095 181.365 73.620 181.585 ;
        RECT 73.040 180.600 73.280 181.195 ;
        RECT 73.450 180.665 73.620 181.365 ;
        RECT 73.790 181.005 73.960 181.785 ;
        RECT 74.280 181.735 74.650 182.235 ;
        RECT 74.830 181.785 75.235 181.955 ;
        RECT 75.405 181.785 76.190 181.955 ;
        RECT 74.830 181.555 75.000 181.785 ;
        RECT 74.170 181.255 75.000 181.555 ;
        RECT 75.385 181.285 75.850 181.615 ;
        RECT 74.170 181.225 74.370 181.255 ;
        RECT 74.490 181.005 74.660 181.075 ;
        RECT 73.790 180.835 74.660 181.005 ;
        RECT 74.150 180.745 74.660 180.835 ;
        RECT 72.700 180.280 73.005 180.410 ;
        RECT 73.450 180.300 73.980 180.665 ;
        RECT 72.320 179.685 72.585 180.145 ;
        RECT 72.755 179.855 73.005 180.280 ;
        RECT 74.150 180.130 74.320 180.745 ;
        RECT 73.215 179.960 74.320 180.130 ;
        RECT 74.490 179.685 74.660 180.485 ;
        RECT 74.830 180.185 75.000 181.255 ;
        RECT 75.170 180.355 75.360 181.075 ;
        RECT 75.530 180.325 75.850 181.285 ;
        RECT 76.020 181.325 76.190 181.785 ;
        RECT 76.465 181.705 76.675 182.235 ;
        RECT 76.935 181.495 77.265 182.020 ;
        RECT 77.435 181.625 77.605 182.235 ;
        RECT 77.775 181.580 78.105 182.015 ;
        RECT 78.325 181.690 83.670 182.235 ;
        RECT 83.845 181.690 89.190 182.235 ;
        RECT 77.775 181.495 78.155 181.580 ;
        RECT 77.065 181.325 77.265 181.495 ;
        RECT 77.930 181.455 78.155 181.495 ;
        RECT 76.020 180.995 76.895 181.325 ;
        RECT 77.065 180.995 77.815 181.325 ;
        RECT 74.830 179.855 75.080 180.185 ;
        RECT 76.020 180.155 76.190 180.995 ;
        RECT 77.065 180.790 77.255 180.995 ;
        RECT 77.985 180.875 78.155 181.455 ;
        RECT 77.940 180.825 78.155 180.875 ;
        RECT 79.910 180.860 80.250 181.690 ;
        RECT 76.360 180.415 77.255 180.790 ;
        RECT 77.765 180.745 78.155 180.825 ;
        RECT 75.305 179.985 76.190 180.155 ;
        RECT 76.370 179.685 76.685 180.185 ;
        RECT 76.915 179.855 77.255 180.415 ;
        RECT 77.425 179.685 77.595 180.695 ;
        RECT 77.765 179.900 78.095 180.745 ;
        RECT 81.730 180.120 82.080 181.370 ;
        RECT 85.430 180.860 85.770 181.690 ;
        RECT 89.365 181.485 90.575 182.235 ;
        RECT 90.745 181.485 91.955 182.235 ;
        RECT 87.250 180.120 87.600 181.370 ;
        RECT 89.365 180.945 89.885 181.485 ;
        RECT 90.055 180.775 90.575 181.315 ;
        RECT 78.325 179.685 83.670 180.120 ;
        RECT 83.845 179.685 89.190 180.120 ;
        RECT 89.365 179.685 90.575 180.775 ;
        RECT 90.745 180.775 91.265 181.315 ;
        RECT 91.435 180.945 91.955 181.485 ;
        RECT 90.745 179.685 91.955 180.775 ;
        RECT 13.380 179.515 92.040 179.685 ;
        RECT 13.465 178.425 14.675 179.515 ;
        RECT 14.845 178.425 18.355 179.515 ;
        RECT 19.045 178.455 19.375 179.300 ;
        RECT 19.545 178.505 19.715 179.515 ;
        RECT 19.885 178.785 20.225 179.345 ;
        RECT 20.455 179.015 20.770 179.515 ;
        RECT 20.950 179.045 21.835 179.215 ;
        RECT 13.465 177.715 13.985 178.255 ;
        RECT 14.155 177.885 14.675 178.425 ;
        RECT 14.845 177.735 16.495 178.255 ;
        RECT 16.665 177.905 18.355 178.425 ;
        RECT 18.985 178.375 19.375 178.455 ;
        RECT 19.885 178.410 20.780 178.785 ;
        RECT 18.985 178.325 19.200 178.375 ;
        RECT 18.985 177.745 19.155 178.325 ;
        RECT 19.885 178.205 20.075 178.410 ;
        RECT 20.950 178.205 21.120 179.045 ;
        RECT 22.060 179.015 22.310 179.345 ;
        RECT 19.325 177.875 20.075 178.205 ;
        RECT 20.245 177.875 21.120 178.205 ;
        RECT 13.465 176.965 14.675 177.715 ;
        RECT 14.845 176.965 18.355 177.735 ;
        RECT 18.985 177.705 19.210 177.745 ;
        RECT 19.875 177.705 20.075 177.875 ;
        RECT 18.985 177.620 19.365 177.705 ;
        RECT 19.035 177.185 19.365 177.620 ;
        RECT 19.535 176.965 19.705 177.575 ;
        RECT 19.875 177.180 20.205 177.705 ;
        RECT 20.465 176.965 20.675 177.495 ;
        RECT 20.950 177.415 21.120 177.875 ;
        RECT 21.290 177.915 21.610 178.875 ;
        RECT 21.780 178.125 21.970 178.845 ;
        RECT 22.140 177.945 22.310 179.015 ;
        RECT 22.480 178.715 22.650 179.515 ;
        RECT 22.820 179.070 23.925 179.240 ;
        RECT 22.820 178.455 22.990 179.070 ;
        RECT 24.135 178.920 24.385 179.345 ;
        RECT 24.555 179.055 24.820 179.515 ;
        RECT 23.160 178.535 23.690 178.900 ;
        RECT 24.135 178.790 24.440 178.920 ;
        RECT 22.480 178.365 22.990 178.455 ;
        RECT 22.480 178.195 23.350 178.365 ;
        RECT 22.480 178.125 22.650 178.195 ;
        RECT 22.770 177.945 22.970 177.975 ;
        RECT 21.290 177.585 21.755 177.915 ;
        RECT 22.140 177.645 22.970 177.945 ;
        RECT 22.140 177.415 22.310 177.645 ;
        RECT 20.950 177.245 21.735 177.415 ;
        RECT 21.905 177.245 22.310 177.415 ;
        RECT 22.490 176.965 22.860 177.465 ;
        RECT 23.180 177.415 23.350 178.195 ;
        RECT 23.520 177.835 23.690 178.535 ;
        RECT 23.860 178.005 24.100 178.600 ;
        RECT 23.520 177.615 24.045 177.835 ;
        RECT 24.270 177.685 24.440 178.790 ;
        RECT 24.215 177.555 24.440 177.685 ;
        RECT 24.610 177.595 24.890 178.545 ;
        RECT 24.215 177.415 24.385 177.555 ;
        RECT 23.180 177.245 23.855 177.415 ;
        RECT 24.050 177.245 24.385 177.415 ;
        RECT 24.555 176.965 24.805 177.425 ;
        RECT 25.060 177.225 25.245 179.345 ;
        RECT 25.415 179.015 25.745 179.515 ;
        RECT 25.915 178.845 26.085 179.345 ;
        RECT 25.420 178.675 26.085 178.845 ;
        RECT 25.420 177.685 25.650 178.675 ;
        RECT 25.820 177.855 26.170 178.505 ;
        RECT 26.345 178.350 26.635 179.515 ;
        RECT 26.805 179.005 27.065 179.515 ;
        RECT 26.805 177.955 27.145 178.835 ;
        RECT 27.315 178.125 27.485 179.345 ;
        RECT 27.725 179.010 28.340 179.515 ;
        RECT 27.725 178.475 27.975 178.840 ;
        RECT 28.145 178.835 28.340 179.010 ;
        RECT 28.510 179.005 28.985 179.345 ;
        RECT 29.155 178.970 29.370 179.515 ;
        RECT 28.145 178.645 28.475 178.835 ;
        RECT 28.695 178.475 29.410 178.770 ;
        RECT 29.580 178.645 29.855 179.345 ;
        RECT 30.115 178.845 30.285 179.345 ;
        RECT 30.455 179.015 30.785 179.515 ;
        RECT 30.115 178.675 30.780 178.845 ;
        RECT 27.725 178.305 29.515 178.475 ;
        RECT 27.315 177.875 28.110 178.125 ;
        RECT 27.315 177.785 27.565 177.875 ;
        RECT 25.420 177.515 26.085 177.685 ;
        RECT 25.415 176.965 25.745 177.345 ;
        RECT 25.915 177.225 26.085 177.515 ;
        RECT 26.345 176.965 26.635 177.690 ;
        RECT 26.805 176.965 27.065 177.785 ;
        RECT 27.235 177.365 27.565 177.785 ;
        RECT 28.280 177.450 28.535 178.305 ;
        RECT 27.745 177.185 28.535 177.450 ;
        RECT 28.705 177.605 29.115 178.125 ;
        RECT 29.285 177.875 29.515 178.305 ;
        RECT 29.685 177.615 29.855 178.645 ;
        RECT 30.030 177.855 30.380 178.505 ;
        RECT 30.550 177.685 30.780 178.675 ;
        RECT 28.705 177.185 28.905 177.605 ;
        RECT 29.095 176.965 29.425 177.425 ;
        RECT 29.595 177.135 29.855 177.615 ;
        RECT 30.115 177.515 30.780 177.685 ;
        RECT 30.115 177.225 30.285 177.515 ;
        RECT 30.455 176.965 30.785 177.345 ;
        RECT 30.955 177.225 31.140 179.345 ;
        RECT 31.380 179.055 31.645 179.515 ;
        RECT 31.815 178.920 32.065 179.345 ;
        RECT 32.275 179.070 33.380 179.240 ;
        RECT 31.760 178.790 32.065 178.920 ;
        RECT 31.310 177.595 31.590 178.545 ;
        RECT 31.760 177.685 31.930 178.790 ;
        RECT 32.100 178.005 32.340 178.600 ;
        RECT 32.510 178.535 33.040 178.900 ;
        RECT 32.510 177.835 32.680 178.535 ;
        RECT 33.210 178.455 33.380 179.070 ;
        RECT 33.550 178.715 33.720 179.515 ;
        RECT 33.890 179.015 34.140 179.345 ;
        RECT 34.365 179.045 35.250 179.215 ;
        RECT 33.210 178.365 33.720 178.455 ;
        RECT 31.760 177.555 31.985 177.685 ;
        RECT 32.155 177.615 32.680 177.835 ;
        RECT 32.850 178.195 33.720 178.365 ;
        RECT 31.395 176.965 31.645 177.425 ;
        RECT 31.815 177.415 31.985 177.555 ;
        RECT 32.850 177.415 33.020 178.195 ;
        RECT 33.550 178.125 33.720 178.195 ;
        RECT 33.230 177.945 33.430 177.975 ;
        RECT 33.890 177.945 34.060 179.015 ;
        RECT 34.230 178.125 34.420 178.845 ;
        RECT 33.230 177.645 34.060 177.945 ;
        RECT 34.590 177.915 34.910 178.875 ;
        RECT 31.815 177.245 32.150 177.415 ;
        RECT 32.345 177.245 33.020 177.415 ;
        RECT 33.340 176.965 33.710 177.465 ;
        RECT 33.890 177.415 34.060 177.645 ;
        RECT 34.445 177.585 34.910 177.915 ;
        RECT 35.080 178.205 35.250 179.045 ;
        RECT 35.430 179.015 35.745 179.515 ;
        RECT 35.975 178.785 36.315 179.345 ;
        RECT 35.420 178.410 36.315 178.785 ;
        RECT 36.485 178.505 36.655 179.515 ;
        RECT 36.125 178.205 36.315 178.410 ;
        RECT 36.825 178.455 37.155 179.300 ;
        RECT 37.865 178.460 38.170 179.245 ;
        RECT 38.350 179.045 39.035 179.515 ;
        RECT 38.345 178.525 39.040 178.835 ;
        RECT 36.825 178.375 37.215 178.455 ;
        RECT 37.000 178.325 37.215 178.375 ;
        RECT 35.080 177.875 35.955 178.205 ;
        RECT 36.125 177.875 36.875 178.205 ;
        RECT 35.080 177.415 35.250 177.875 ;
        RECT 36.125 177.705 36.325 177.875 ;
        RECT 37.045 177.745 37.215 178.325 ;
        RECT 36.990 177.705 37.215 177.745 ;
        RECT 33.890 177.245 34.295 177.415 ;
        RECT 34.465 177.245 35.250 177.415 ;
        RECT 35.525 176.965 35.735 177.495 ;
        RECT 35.995 177.180 36.325 177.705 ;
        RECT 36.835 177.620 37.215 177.705 ;
        RECT 37.865 177.655 38.040 178.460 ;
        RECT 39.215 178.355 39.500 179.300 ;
        RECT 39.675 179.065 40.005 179.515 ;
        RECT 40.175 178.895 40.345 179.325 ;
        RECT 40.605 179.080 45.950 179.515 ;
        RECT 38.640 178.205 39.500 178.355 ;
        RECT 38.215 178.185 39.500 178.205 ;
        RECT 39.670 178.665 40.345 178.895 ;
        RECT 38.215 177.825 39.200 178.185 ;
        RECT 39.670 178.015 39.905 178.665 ;
        RECT 36.495 176.965 36.665 177.575 ;
        RECT 36.835 177.185 37.165 177.620 ;
        RECT 37.865 177.135 38.105 177.655 ;
        RECT 39.030 177.490 39.200 177.825 ;
        RECT 39.370 177.685 39.905 178.015 ;
        RECT 39.685 177.535 39.905 177.685 ;
        RECT 40.075 177.645 40.375 178.495 ;
        RECT 38.275 176.965 38.670 177.460 ;
        RECT 39.030 177.295 39.405 177.490 ;
        RECT 39.235 177.150 39.405 177.295 ;
        RECT 39.685 177.160 39.925 177.535 ;
        RECT 42.190 177.510 42.530 178.340 ;
        RECT 44.010 177.830 44.360 179.080 ;
        RECT 46.310 178.545 46.700 178.720 ;
        RECT 47.185 178.715 47.515 179.515 ;
        RECT 47.685 178.725 48.220 179.345 ;
        RECT 48.890 179.005 50.545 179.295 ;
        RECT 46.310 178.375 47.735 178.545 ;
        RECT 46.185 177.645 46.540 178.205 ;
        RECT 40.095 176.965 40.430 177.470 ;
        RECT 40.605 176.965 45.950 177.510 ;
        RECT 46.710 177.475 46.880 178.375 ;
        RECT 47.050 177.645 47.315 178.205 ;
        RECT 47.565 177.875 47.735 178.375 ;
        RECT 47.905 177.705 48.220 178.725 ;
        RECT 48.890 178.665 50.480 178.835 ;
        RECT 50.715 178.715 50.995 179.515 ;
        RECT 48.890 178.375 49.210 178.665 ;
        RECT 50.310 178.545 50.480 178.665 ;
        RECT 49.405 178.325 50.120 178.495 ;
        RECT 50.310 178.375 51.035 178.545 ;
        RECT 51.205 178.375 51.475 179.345 ;
        RECT 46.290 176.965 46.530 177.475 ;
        RECT 46.710 177.145 46.990 177.475 ;
        RECT 47.220 176.965 47.435 177.475 ;
        RECT 47.605 177.135 48.220 177.705 ;
        RECT 48.890 177.635 49.240 178.205 ;
        RECT 49.410 177.875 50.120 178.325 ;
        RECT 50.865 178.205 51.035 178.375 ;
        RECT 50.290 177.875 50.695 178.205 ;
        RECT 50.865 177.875 51.135 178.205 ;
        RECT 50.865 177.705 51.035 177.875 ;
        RECT 49.425 177.535 51.035 177.705 ;
        RECT 51.305 177.640 51.475 178.375 ;
        RECT 52.105 178.350 52.395 179.515 ;
        RECT 48.895 176.965 49.225 177.465 ;
        RECT 49.425 177.185 49.595 177.535 ;
        RECT 49.795 176.965 50.125 177.365 ;
        RECT 50.295 177.185 50.465 177.535 ;
        RECT 50.635 176.965 51.015 177.365 ;
        RECT 51.205 177.295 51.475 177.640 ;
        RECT 52.105 176.965 52.395 177.690 ;
        RECT 52.565 177.245 52.845 179.345 ;
        RECT 53.035 178.755 53.820 179.515 ;
        RECT 54.215 178.685 54.600 179.345 ;
        RECT 54.215 178.585 54.625 178.685 ;
        RECT 53.015 178.375 54.625 178.585 ;
        RECT 54.925 178.495 55.125 179.285 ;
        RECT 53.015 177.775 53.290 178.375 ;
        RECT 54.795 178.325 55.125 178.495 ;
        RECT 55.295 178.335 55.615 179.515 ;
        RECT 56.245 178.375 56.505 179.515 ;
        RECT 56.675 178.365 57.005 179.345 ;
        RECT 57.175 178.375 57.455 179.515 ;
        RECT 57.625 178.645 57.900 179.345 ;
        RECT 58.070 178.970 58.325 179.515 ;
        RECT 58.495 179.005 58.975 179.345 ;
        RECT 59.150 178.960 59.755 179.515 ;
        RECT 59.140 178.860 59.755 178.960 ;
        RECT 59.140 178.835 59.325 178.860 ;
        RECT 54.795 178.205 54.975 178.325 ;
        RECT 53.460 177.955 53.815 178.205 ;
        RECT 54.010 178.155 54.475 178.205 ;
        RECT 54.005 177.985 54.475 178.155 ;
        RECT 54.010 177.955 54.475 177.985 ;
        RECT 54.645 177.955 54.975 178.205 ;
        RECT 55.150 177.955 55.615 178.155 ;
        RECT 56.265 177.955 56.600 178.205 ;
        RECT 53.015 177.595 54.265 177.775 ;
        RECT 56.770 177.765 56.940 178.365 ;
        RECT 57.110 177.935 57.445 178.205 ;
        RECT 53.900 177.525 54.265 177.595 ;
        RECT 54.435 177.575 55.615 177.745 ;
        RECT 53.075 176.965 53.245 177.425 ;
        RECT 54.435 177.355 54.765 177.575 ;
        RECT 53.515 177.175 54.765 177.355 ;
        RECT 54.935 176.965 55.105 177.405 ;
        RECT 55.275 177.160 55.615 177.575 ;
        RECT 56.245 177.135 56.940 177.765 ;
        RECT 57.145 176.965 57.455 177.765 ;
        RECT 57.625 177.615 57.795 178.645 ;
        RECT 58.070 178.515 58.825 178.765 ;
        RECT 58.995 178.590 59.325 178.835 ;
        RECT 59.930 178.715 60.245 179.515 ;
        RECT 60.510 179.160 61.590 179.330 ;
        RECT 58.070 178.480 58.840 178.515 ;
        RECT 58.070 178.470 58.855 178.480 ;
        RECT 57.965 178.455 58.860 178.470 ;
        RECT 57.965 178.440 58.880 178.455 ;
        RECT 57.965 178.430 58.900 178.440 ;
        RECT 57.965 178.420 58.925 178.430 ;
        RECT 57.965 178.390 58.995 178.420 ;
        RECT 57.965 178.360 59.015 178.390 ;
        RECT 57.965 178.330 59.035 178.360 ;
        RECT 57.965 178.305 59.065 178.330 ;
        RECT 57.965 178.270 59.100 178.305 ;
        RECT 57.965 178.265 59.130 178.270 ;
        RECT 57.965 177.870 58.195 178.265 ;
        RECT 58.740 178.260 59.130 178.265 ;
        RECT 58.765 178.250 59.130 178.260 ;
        RECT 58.780 178.245 59.130 178.250 ;
        RECT 58.795 178.240 59.130 178.245 ;
        RECT 59.495 178.240 59.755 178.690 ;
        RECT 60.510 178.545 60.680 179.160 ;
        RECT 58.795 178.235 59.755 178.240 ;
        RECT 58.805 178.225 59.755 178.235 ;
        RECT 58.815 178.220 59.755 178.225 ;
        RECT 58.825 178.210 59.755 178.220 ;
        RECT 58.830 178.200 59.755 178.210 ;
        RECT 58.835 178.195 59.755 178.200 ;
        RECT 58.845 178.180 59.755 178.195 ;
        RECT 58.850 178.165 59.755 178.180 ;
        RECT 58.860 178.140 59.755 178.165 ;
        RECT 58.365 177.670 58.695 178.095 ;
        RECT 57.625 177.135 57.885 177.615 ;
        RECT 58.055 176.965 58.305 177.505 ;
        RECT 58.475 177.185 58.695 177.670 ;
        RECT 58.865 178.070 59.755 178.140 ;
        RECT 58.865 177.345 59.035 178.070 ;
        RECT 59.205 177.515 59.755 177.900 ;
        RECT 59.925 177.535 60.195 178.545 ;
        RECT 60.365 178.375 60.680 178.545 ;
        RECT 60.365 177.705 60.535 178.375 ;
        RECT 60.850 178.205 61.085 178.885 ;
        RECT 61.255 178.375 61.590 179.160 ;
        RECT 62.685 178.375 63.025 179.345 ;
        RECT 63.195 178.375 63.365 179.515 ;
        RECT 63.635 178.715 63.885 179.515 ;
        RECT 64.530 178.545 64.860 179.345 ;
        RECT 65.160 178.715 65.490 179.515 ;
        RECT 65.660 178.545 65.990 179.345 ;
        RECT 63.555 178.375 65.990 178.545 ;
        RECT 66.365 178.425 69.875 179.515 ;
        RECT 60.705 177.875 61.085 178.205 ;
        RECT 61.255 177.875 61.590 178.205 ;
        RECT 62.685 177.765 62.860 178.375 ;
        RECT 63.555 178.125 63.725 178.375 ;
        RECT 63.030 177.955 63.725 178.125 ;
        RECT 63.900 177.955 64.320 178.155 ;
        RECT 64.490 177.955 64.820 178.155 ;
        RECT 64.990 177.955 65.320 178.155 ;
        RECT 60.365 177.535 61.590 177.705 ;
        RECT 58.865 177.175 59.755 177.345 ;
        RECT 59.995 176.965 60.325 177.365 ;
        RECT 60.495 177.265 60.665 177.535 ;
        RECT 60.835 176.965 61.165 177.365 ;
        RECT 61.335 177.265 61.590 177.535 ;
        RECT 62.685 177.135 63.025 177.765 ;
        RECT 63.195 176.965 63.445 177.765 ;
        RECT 63.635 177.615 64.860 177.785 ;
        RECT 63.635 177.135 63.965 177.615 ;
        RECT 64.135 176.965 64.360 177.425 ;
        RECT 64.530 177.135 64.860 177.615 ;
        RECT 65.490 177.745 65.660 178.375 ;
        RECT 65.845 177.955 66.195 178.205 ;
        RECT 65.490 177.135 65.990 177.745 ;
        RECT 66.365 177.735 68.015 178.255 ;
        RECT 68.185 177.905 69.875 178.425 ;
        RECT 70.055 178.375 70.385 179.515 ;
        RECT 70.915 178.545 71.245 179.330 ;
        RECT 70.565 178.375 71.245 178.545 ;
        RECT 71.435 178.545 71.765 179.330 ;
        RECT 71.435 178.375 72.115 178.545 ;
        RECT 72.295 178.375 72.625 179.515 ;
        RECT 72.805 178.425 76.315 179.515 ;
        RECT 76.485 178.425 77.695 179.515 ;
        RECT 70.045 177.955 70.395 178.205 ;
        RECT 70.565 177.775 70.735 178.375 ;
        RECT 70.905 177.955 71.255 178.205 ;
        RECT 71.425 177.955 71.775 178.205 ;
        RECT 71.945 177.775 72.115 178.375 ;
        RECT 72.285 177.955 72.635 178.205 ;
        RECT 66.365 176.965 69.875 177.735 ;
        RECT 70.055 176.965 70.325 177.775 ;
        RECT 70.495 177.135 70.825 177.775 ;
        RECT 70.995 176.965 71.235 177.775 ;
        RECT 71.445 176.965 71.685 177.775 ;
        RECT 71.855 177.135 72.185 177.775 ;
        RECT 72.355 176.965 72.625 177.775 ;
        RECT 72.805 177.735 74.455 178.255 ;
        RECT 74.625 177.905 76.315 178.425 ;
        RECT 72.805 176.965 76.315 177.735 ;
        RECT 76.485 177.715 77.005 178.255 ;
        RECT 77.175 177.885 77.695 178.425 ;
        RECT 77.865 178.350 78.155 179.515 ;
        RECT 78.325 179.080 83.670 179.515 ;
        RECT 83.845 179.080 89.190 179.515 ;
        RECT 76.485 176.965 77.695 177.715 ;
        RECT 77.865 176.965 78.155 177.690 ;
        RECT 79.910 177.510 80.250 178.340 ;
        RECT 81.730 177.830 82.080 179.080 ;
        RECT 85.430 177.510 85.770 178.340 ;
        RECT 87.250 177.830 87.600 179.080 ;
        RECT 89.365 178.425 90.575 179.515 ;
        RECT 89.365 177.715 89.885 178.255 ;
        RECT 90.055 177.885 90.575 178.425 ;
        RECT 90.745 178.425 91.955 179.515 ;
        RECT 90.745 177.885 91.265 178.425 ;
        RECT 91.435 177.715 91.955 178.255 ;
        RECT 78.325 176.965 83.670 177.510 ;
        RECT 83.845 176.965 89.190 177.510 ;
        RECT 89.365 176.965 90.575 177.715 ;
        RECT 90.745 176.965 91.955 177.715 ;
        RECT 13.380 176.795 92.040 176.965 ;
        RECT 13.465 176.045 14.675 176.795 ;
        RECT 14.845 176.250 20.190 176.795 ;
        RECT 20.830 176.290 21.165 176.795 ;
        RECT 13.465 175.505 13.985 176.045 ;
        RECT 14.155 175.335 14.675 175.875 ;
        RECT 16.430 175.420 16.770 176.250 ;
        RECT 21.335 176.225 21.575 176.600 ;
        RECT 21.855 176.465 22.025 176.610 ;
        RECT 21.855 176.270 22.230 176.465 ;
        RECT 22.590 176.300 22.985 176.795 ;
        RECT 13.465 174.245 14.675 175.335 ;
        RECT 18.250 174.680 18.600 175.930 ;
        RECT 20.885 175.265 21.185 176.115 ;
        RECT 21.355 176.075 21.575 176.225 ;
        RECT 21.355 175.745 21.890 176.075 ;
        RECT 22.060 175.935 22.230 176.270 ;
        RECT 23.155 176.105 23.395 176.625 ;
        RECT 23.585 176.250 28.930 176.795 ;
        RECT 29.105 176.250 34.450 176.795 ;
        RECT 21.355 175.095 21.590 175.745 ;
        RECT 22.060 175.575 23.045 175.935 ;
        RECT 20.915 174.865 21.590 175.095 ;
        RECT 21.760 175.555 23.045 175.575 ;
        RECT 21.760 175.405 22.620 175.555 ;
        RECT 14.845 174.245 20.190 174.680 ;
        RECT 20.915 174.435 21.085 174.865 ;
        RECT 21.255 174.245 21.585 174.695 ;
        RECT 21.760 174.460 22.045 175.405 ;
        RECT 23.220 175.300 23.395 176.105 ;
        RECT 25.170 175.420 25.510 176.250 ;
        RECT 22.220 174.925 22.915 175.235 ;
        RECT 22.225 174.245 22.910 174.715 ;
        RECT 23.090 174.515 23.395 175.300 ;
        RECT 26.990 174.680 27.340 175.930 ;
        RECT 30.690 175.420 31.030 176.250 ;
        RECT 34.625 176.025 38.135 176.795 ;
        RECT 39.225 176.070 39.515 176.795 ;
        RECT 39.685 176.025 43.195 176.795 ;
        RECT 43.365 176.045 44.575 176.795 ;
        RECT 32.510 174.680 32.860 175.930 ;
        RECT 34.625 175.505 36.275 176.025 ;
        RECT 36.445 175.335 38.135 175.855 ;
        RECT 39.685 175.505 41.335 176.025 ;
        RECT 23.585 174.245 28.930 174.680 ;
        RECT 29.105 174.245 34.450 174.680 ;
        RECT 34.625 174.245 38.135 175.335 ;
        RECT 39.225 174.245 39.515 175.410 ;
        RECT 41.505 175.335 43.195 175.855 ;
        RECT 43.365 175.505 43.885 176.045 ;
        RECT 44.765 175.985 45.005 176.795 ;
        RECT 45.175 175.985 45.505 176.625 ;
        RECT 45.675 175.985 45.945 176.795 ;
        RECT 46.125 176.250 51.470 176.795 ;
        RECT 51.645 176.250 56.990 176.795 ;
        RECT 57.165 176.250 62.510 176.795 ;
        RECT 44.055 175.335 44.575 175.875 ;
        RECT 44.745 175.555 45.095 175.805 ;
        RECT 45.265 175.385 45.435 175.985 ;
        RECT 45.605 175.555 45.955 175.805 ;
        RECT 47.710 175.420 48.050 176.250 ;
        RECT 39.685 174.245 43.195 175.335 ;
        RECT 43.365 174.245 44.575 175.335 ;
        RECT 44.755 175.215 45.435 175.385 ;
        RECT 44.755 174.430 45.085 175.215 ;
        RECT 45.615 174.245 45.945 175.385 ;
        RECT 49.530 174.680 49.880 175.930 ;
        RECT 53.230 175.420 53.570 176.250 ;
        RECT 55.050 174.680 55.400 175.930 ;
        RECT 58.750 175.420 59.090 176.250 ;
        RECT 62.685 176.025 64.355 176.795 ;
        RECT 64.985 176.070 65.275 176.795 ;
        RECT 65.445 176.025 68.035 176.795 ;
        RECT 60.570 174.680 60.920 175.930 ;
        RECT 62.685 175.505 63.435 176.025 ;
        RECT 63.605 175.335 64.355 175.855 ;
        RECT 65.445 175.505 66.655 176.025 ;
        RECT 68.265 175.975 68.475 176.795 ;
        RECT 68.645 175.995 68.975 176.625 ;
        RECT 46.125 174.245 51.470 174.680 ;
        RECT 51.645 174.245 56.990 174.680 ;
        RECT 57.165 174.245 62.510 174.680 ;
        RECT 62.685 174.245 64.355 175.335 ;
        RECT 64.985 174.245 65.275 175.410 ;
        RECT 66.825 175.335 68.035 175.855 ;
        RECT 68.645 175.395 68.895 175.995 ;
        RECT 69.145 175.975 69.375 176.795 ;
        RECT 70.525 175.985 70.765 176.795 ;
        RECT 70.935 175.985 71.265 176.625 ;
        RECT 71.435 175.985 71.705 176.795 ;
        RECT 71.895 175.985 72.165 176.795 ;
        RECT 72.335 175.985 72.665 176.625 ;
        RECT 72.835 175.985 73.075 176.795 ;
        RECT 73.265 175.995 73.960 176.625 ;
        RECT 74.165 175.995 74.475 176.795 ;
        RECT 74.645 176.250 79.990 176.795 ;
        RECT 80.165 176.250 85.510 176.795 ;
        RECT 69.065 175.555 69.395 175.805 ;
        RECT 70.505 175.555 70.855 175.805 ;
        RECT 65.445 174.245 68.035 175.335 ;
        RECT 68.265 174.245 68.475 175.385 ;
        RECT 68.645 174.415 68.975 175.395 ;
        RECT 71.025 175.385 71.195 175.985 ;
        RECT 71.365 175.555 71.715 175.805 ;
        RECT 71.885 175.555 72.235 175.805 ;
        RECT 72.405 175.385 72.575 175.985 ;
        RECT 73.785 175.945 73.960 175.995 ;
        RECT 72.745 175.555 73.095 175.805 ;
        RECT 73.285 175.555 73.620 175.805 ;
        RECT 73.790 175.395 73.960 175.945 ;
        RECT 74.130 175.555 74.465 175.825 ;
        RECT 76.230 175.420 76.570 176.250 ;
        RECT 69.145 174.245 69.375 175.385 ;
        RECT 70.515 175.215 71.195 175.385 ;
        RECT 70.515 174.430 70.845 175.215 ;
        RECT 71.375 174.245 71.705 175.385 ;
        RECT 71.895 174.245 72.225 175.385 ;
        RECT 72.405 175.215 73.085 175.385 ;
        RECT 72.755 174.430 73.085 175.215 ;
        RECT 73.265 174.245 73.525 175.385 ;
        RECT 73.695 174.415 74.025 175.395 ;
        RECT 74.195 174.245 74.475 175.385 ;
        RECT 78.050 174.680 78.400 175.930 ;
        RECT 81.750 175.420 82.090 176.250 ;
        RECT 85.685 176.025 89.195 176.795 ;
        RECT 89.365 176.045 90.575 176.795 ;
        RECT 90.745 176.045 91.955 176.795 ;
        RECT 100.630 176.790 106.370 176.800 ;
        RECT 83.570 174.680 83.920 175.930 ;
        RECT 85.685 175.505 87.335 176.025 ;
        RECT 87.505 175.335 89.195 175.855 ;
        RECT 89.365 175.505 89.885 176.045 ;
        RECT 90.055 175.335 90.575 175.875 ;
        RECT 74.645 174.245 79.990 174.680 ;
        RECT 80.165 174.245 85.510 174.680 ;
        RECT 85.685 174.245 89.195 175.335 ;
        RECT 89.365 174.245 90.575 175.335 ;
        RECT 90.745 175.335 91.265 175.875 ;
        RECT 91.435 175.505 91.955 176.045 ;
        RECT 100.140 176.630 106.370 176.790 ;
        RECT 90.745 174.245 91.955 175.335 ;
        RECT 100.140 174.370 100.810 176.630 ;
        RECT 101.480 176.060 105.520 176.230 ;
        RECT 101.140 175.000 101.310 176.000 ;
        RECT 105.690 175.000 105.860 176.000 ;
        RECT 101.480 174.770 105.520 174.940 ;
        RECT 106.200 174.370 106.370 176.630 ;
        RECT 13.380 174.075 92.040 174.245 ;
        RECT 100.140 174.200 106.370 174.370 ;
        RECT 13.465 172.985 14.675 174.075 ;
        RECT 14.845 173.640 20.190 174.075 ;
        RECT 20.365 173.640 25.710 174.075 ;
        RECT 13.465 172.275 13.985 172.815 ;
        RECT 14.155 172.445 14.675 172.985 ;
        RECT 13.465 171.525 14.675 172.275 ;
        RECT 16.430 172.070 16.770 172.900 ;
        RECT 18.250 172.390 18.600 173.640 ;
        RECT 21.950 172.070 22.290 172.900 ;
        RECT 23.770 172.390 24.120 173.640 ;
        RECT 26.345 172.910 26.635 174.075 ;
        RECT 26.805 172.985 29.395 174.075 ;
        RECT 30.025 173.520 30.630 174.075 ;
        RECT 30.805 173.565 31.285 173.905 ;
        RECT 31.455 173.530 31.710 174.075 ;
        RECT 30.025 173.420 30.640 173.520 ;
        RECT 30.455 173.395 30.640 173.420 ;
        RECT 26.805 172.295 28.015 172.815 ;
        RECT 28.185 172.465 29.395 172.985 ;
        RECT 30.025 172.800 30.285 173.250 ;
        RECT 30.455 173.150 30.785 173.395 ;
        RECT 30.955 173.075 31.710 173.325 ;
        RECT 31.880 173.205 32.155 173.905 ;
        RECT 30.940 173.040 31.710 173.075 ;
        RECT 30.925 173.030 31.710 173.040 ;
        RECT 30.920 173.015 31.815 173.030 ;
        RECT 30.900 173.000 31.815 173.015 ;
        RECT 30.880 172.990 31.815 173.000 ;
        RECT 30.855 172.980 31.815 172.990 ;
        RECT 30.785 172.950 31.815 172.980 ;
        RECT 30.765 172.920 31.815 172.950 ;
        RECT 30.745 172.890 31.815 172.920 ;
        RECT 30.715 172.865 31.815 172.890 ;
        RECT 30.680 172.830 31.815 172.865 ;
        RECT 30.650 172.825 31.815 172.830 ;
        RECT 30.650 172.820 31.040 172.825 ;
        RECT 30.650 172.810 31.015 172.820 ;
        RECT 30.650 172.805 31.000 172.810 ;
        RECT 30.650 172.800 30.985 172.805 ;
        RECT 30.025 172.795 30.985 172.800 ;
        RECT 30.025 172.785 30.975 172.795 ;
        RECT 30.025 172.780 30.965 172.785 ;
        RECT 30.025 172.770 30.955 172.780 ;
        RECT 30.025 172.760 30.950 172.770 ;
        RECT 30.025 172.755 30.945 172.760 ;
        RECT 30.025 172.740 30.935 172.755 ;
        RECT 30.025 172.725 30.930 172.740 ;
        RECT 30.025 172.700 30.920 172.725 ;
        RECT 30.025 172.630 30.915 172.700 ;
        RECT 14.845 171.525 20.190 172.070 ;
        RECT 20.365 171.525 25.710 172.070 ;
        RECT 26.345 171.525 26.635 172.250 ;
        RECT 26.805 171.525 29.395 172.295 ;
        RECT 30.025 172.075 30.575 172.460 ;
        RECT 30.745 171.905 30.915 172.630 ;
        RECT 30.025 171.735 30.915 171.905 ;
        RECT 31.085 172.230 31.415 172.655 ;
        RECT 31.585 172.430 31.815 172.825 ;
        RECT 31.085 171.745 31.305 172.230 ;
        RECT 31.985 172.175 32.155 173.205 ;
        RECT 31.475 171.525 31.725 172.065 ;
        RECT 31.895 171.695 32.155 172.175 ;
        RECT 32.325 173.205 32.600 173.905 ;
        RECT 32.770 173.530 33.025 174.075 ;
        RECT 33.195 173.565 33.675 173.905 ;
        RECT 33.850 173.520 34.455 174.075 ;
        RECT 33.840 173.420 34.455 173.520 ;
        RECT 33.840 173.395 34.025 173.420 ;
        RECT 32.325 172.175 32.495 173.205 ;
        RECT 32.770 173.075 33.525 173.325 ;
        RECT 33.695 173.150 34.025 173.395 ;
        RECT 32.770 173.040 33.540 173.075 ;
        RECT 32.770 173.030 33.555 173.040 ;
        RECT 32.665 173.015 33.560 173.030 ;
        RECT 32.665 173.000 33.580 173.015 ;
        RECT 32.665 172.990 33.600 173.000 ;
        RECT 32.665 172.980 33.625 172.990 ;
        RECT 32.665 172.950 33.695 172.980 ;
        RECT 32.665 172.920 33.715 172.950 ;
        RECT 32.665 172.890 33.735 172.920 ;
        RECT 32.665 172.865 33.765 172.890 ;
        RECT 32.665 172.830 33.800 172.865 ;
        RECT 32.665 172.825 33.830 172.830 ;
        RECT 32.665 172.430 32.895 172.825 ;
        RECT 33.440 172.820 33.830 172.825 ;
        RECT 33.465 172.810 33.830 172.820 ;
        RECT 33.480 172.805 33.830 172.810 ;
        RECT 33.495 172.800 33.830 172.805 ;
        RECT 34.195 172.800 34.455 173.250 ;
        RECT 34.625 172.985 37.215 174.075 ;
        RECT 38.095 173.345 38.390 174.075 ;
        RECT 38.560 173.175 38.820 173.900 ;
        RECT 38.990 173.345 39.250 174.075 ;
        RECT 39.420 173.175 39.680 173.900 ;
        RECT 39.850 173.345 40.110 174.075 ;
        RECT 40.280 173.175 40.540 173.900 ;
        RECT 40.710 173.345 40.970 174.075 ;
        RECT 41.140 173.175 41.400 173.900 ;
        RECT 33.495 172.795 34.455 172.800 ;
        RECT 33.505 172.785 34.455 172.795 ;
        RECT 33.515 172.780 34.455 172.785 ;
        RECT 33.525 172.770 34.455 172.780 ;
        RECT 33.530 172.760 34.455 172.770 ;
        RECT 33.535 172.755 34.455 172.760 ;
        RECT 33.545 172.740 34.455 172.755 ;
        RECT 33.550 172.725 34.455 172.740 ;
        RECT 33.560 172.700 34.455 172.725 ;
        RECT 33.065 172.230 33.395 172.655 ;
        RECT 33.145 172.205 33.395 172.230 ;
        RECT 32.325 171.695 32.585 172.175 ;
        RECT 32.755 171.525 33.005 172.065 ;
        RECT 33.175 171.745 33.395 172.205 ;
        RECT 33.565 172.630 34.455 172.700 ;
        RECT 33.565 171.905 33.735 172.630 ;
        RECT 33.905 172.075 34.455 172.460 ;
        RECT 34.625 172.295 35.835 172.815 ;
        RECT 36.005 172.465 37.215 172.985 ;
        RECT 38.090 172.935 41.400 173.175 ;
        RECT 41.570 172.965 41.830 174.075 ;
        RECT 38.090 172.345 39.060 172.935 ;
        RECT 42.000 172.765 42.250 173.900 ;
        RECT 42.430 172.965 42.725 174.075 ;
        RECT 42.905 173.205 43.180 173.905 ;
        RECT 43.350 173.530 43.605 174.075 ;
        RECT 43.775 173.565 44.255 173.905 ;
        RECT 44.430 173.520 45.035 174.075 ;
        RECT 44.420 173.420 45.035 173.520 ;
        RECT 44.420 173.395 44.605 173.420 ;
        RECT 39.230 172.515 42.250 172.765 ;
        RECT 33.565 171.735 34.455 171.905 ;
        RECT 34.625 171.525 37.215 172.295 ;
        RECT 38.090 172.175 41.400 172.345 ;
        RECT 38.090 171.525 38.390 172.005 ;
        RECT 38.560 171.720 38.820 172.175 ;
        RECT 38.990 171.525 39.250 172.005 ;
        RECT 39.420 171.720 39.680 172.175 ;
        RECT 39.850 171.525 40.110 172.005 ;
        RECT 40.280 171.720 40.540 172.175 ;
        RECT 40.710 171.525 40.970 172.005 ;
        RECT 41.140 171.720 41.400 172.175 ;
        RECT 41.570 171.525 41.830 172.050 ;
        RECT 42.000 171.705 42.250 172.515 ;
        RECT 42.420 172.155 42.735 172.765 ;
        RECT 42.905 172.175 43.075 173.205 ;
        RECT 43.350 173.075 44.105 173.325 ;
        RECT 44.275 173.150 44.605 173.395 ;
        RECT 43.350 173.040 44.120 173.075 ;
        RECT 43.350 173.030 44.135 173.040 ;
        RECT 43.245 173.015 44.140 173.030 ;
        RECT 43.245 173.000 44.160 173.015 ;
        RECT 43.245 172.990 44.180 173.000 ;
        RECT 43.245 172.980 44.205 172.990 ;
        RECT 43.245 172.950 44.275 172.980 ;
        RECT 43.245 172.920 44.295 172.950 ;
        RECT 43.245 172.890 44.315 172.920 ;
        RECT 43.245 172.865 44.345 172.890 ;
        RECT 43.245 172.830 44.380 172.865 ;
        RECT 43.245 172.825 44.410 172.830 ;
        RECT 43.245 172.430 43.475 172.825 ;
        RECT 44.020 172.820 44.410 172.825 ;
        RECT 44.045 172.810 44.410 172.820 ;
        RECT 44.060 172.805 44.410 172.810 ;
        RECT 44.075 172.800 44.410 172.805 ;
        RECT 44.775 172.800 45.035 173.250 ;
        RECT 44.075 172.795 45.035 172.800 ;
        RECT 44.085 172.785 45.035 172.795 ;
        RECT 44.095 172.780 45.035 172.785 ;
        RECT 44.105 172.770 45.035 172.780 ;
        RECT 44.110 172.760 45.035 172.770 ;
        RECT 44.115 172.755 45.035 172.760 ;
        RECT 44.125 172.740 45.035 172.755 ;
        RECT 44.130 172.725 45.035 172.740 ;
        RECT 44.140 172.700 45.035 172.725 ;
        RECT 43.645 172.230 43.975 172.655 ;
        RECT 42.430 171.525 42.675 171.985 ;
        RECT 42.905 171.695 43.165 172.175 ;
        RECT 43.335 171.525 43.585 172.065 ;
        RECT 43.755 171.745 43.975 172.230 ;
        RECT 44.145 172.630 45.035 172.700 ;
        RECT 45.205 173.205 45.480 173.905 ;
        RECT 45.650 173.530 45.905 174.075 ;
        RECT 46.075 173.565 46.555 173.905 ;
        RECT 46.730 173.520 47.335 174.075 ;
        RECT 46.720 173.420 47.335 173.520 ;
        RECT 47.515 173.465 47.845 173.895 ;
        RECT 48.025 173.635 48.220 174.075 ;
        RECT 48.390 173.465 48.720 173.895 ;
        RECT 46.720 173.395 46.905 173.420 ;
        RECT 44.145 171.905 44.315 172.630 ;
        RECT 44.485 172.075 45.035 172.460 ;
        RECT 45.205 172.175 45.375 173.205 ;
        RECT 45.650 173.075 46.405 173.325 ;
        RECT 46.575 173.150 46.905 173.395 ;
        RECT 47.515 173.295 48.720 173.465 ;
        RECT 45.650 173.040 46.420 173.075 ;
        RECT 45.650 173.030 46.435 173.040 ;
        RECT 45.545 173.015 46.440 173.030 ;
        RECT 45.545 173.000 46.460 173.015 ;
        RECT 45.545 172.990 46.480 173.000 ;
        RECT 45.545 172.980 46.505 172.990 ;
        RECT 45.545 172.950 46.575 172.980 ;
        RECT 45.545 172.920 46.595 172.950 ;
        RECT 45.545 172.890 46.615 172.920 ;
        RECT 45.545 172.865 46.645 172.890 ;
        RECT 45.545 172.830 46.680 172.865 ;
        RECT 45.545 172.825 46.710 172.830 ;
        RECT 45.545 172.430 45.775 172.825 ;
        RECT 46.320 172.820 46.710 172.825 ;
        RECT 46.345 172.810 46.710 172.820 ;
        RECT 46.360 172.805 46.710 172.810 ;
        RECT 46.375 172.800 46.710 172.805 ;
        RECT 47.075 172.800 47.335 173.250 ;
        RECT 47.515 172.965 48.410 173.295 ;
        RECT 48.890 173.125 49.165 173.895 ;
        RECT 46.375 172.795 47.335 172.800 ;
        RECT 46.385 172.785 47.335 172.795 ;
        RECT 46.395 172.780 47.335 172.785 ;
        RECT 46.405 172.770 47.335 172.780 ;
        RECT 46.410 172.760 47.335 172.770 ;
        RECT 48.580 172.935 49.165 173.125 ;
        RECT 49.345 172.985 51.935 174.075 ;
        RECT 46.415 172.755 47.335 172.760 ;
        RECT 46.425 172.740 47.335 172.755 ;
        RECT 46.430 172.725 47.335 172.740 ;
        RECT 46.440 172.700 47.335 172.725 ;
        RECT 45.945 172.230 46.275 172.655 ;
        RECT 44.145 171.735 45.035 171.905 ;
        RECT 45.205 171.695 45.465 172.175 ;
        RECT 45.635 171.525 45.885 172.065 ;
        RECT 46.055 171.745 46.275 172.230 ;
        RECT 46.445 172.630 47.335 172.700 ;
        RECT 46.445 171.905 46.615 172.630 ;
        RECT 46.785 172.075 47.335 172.460 ;
        RECT 47.520 172.435 47.815 172.765 ;
        RECT 47.995 172.435 48.410 172.765 ;
        RECT 46.445 171.735 47.335 171.905 ;
        RECT 47.515 171.525 47.815 172.255 ;
        RECT 47.995 171.815 48.225 172.435 ;
        RECT 48.580 172.265 48.755 172.935 ;
        RECT 48.425 172.085 48.755 172.265 ;
        RECT 48.925 172.115 49.165 172.765 ;
        RECT 49.345 172.295 50.555 172.815 ;
        RECT 50.725 172.465 51.935 172.985 ;
        RECT 52.105 172.910 52.395 174.075 ;
        RECT 52.565 173.105 52.835 173.875 ;
        RECT 53.005 173.295 53.335 174.075 ;
        RECT 53.540 173.470 53.725 173.875 ;
        RECT 53.895 173.650 54.230 174.075 ;
        RECT 54.410 173.650 54.745 174.075 ;
        RECT 54.915 173.470 55.100 173.875 ;
        RECT 53.540 173.295 54.205 173.470 ;
        RECT 52.565 172.935 53.695 173.105 ;
        RECT 48.425 171.705 48.650 172.085 ;
        RECT 48.820 171.525 49.150 171.915 ;
        RECT 49.345 171.525 51.935 172.295 ;
        RECT 52.105 171.525 52.395 172.250 ;
        RECT 52.565 172.025 52.735 172.935 ;
        RECT 52.905 172.185 53.265 172.765 ;
        RECT 53.445 172.435 53.695 172.935 ;
        RECT 53.865 172.265 54.205 173.295 ;
        RECT 53.520 172.095 54.205 172.265 ;
        RECT 54.435 173.295 55.100 173.470 ;
        RECT 55.305 173.295 55.635 174.075 ;
        RECT 54.435 172.265 54.775 173.295 ;
        RECT 55.805 173.105 56.075 173.875 ;
        RECT 54.945 172.935 56.075 173.105 ;
        RECT 56.245 172.985 57.455 174.075 ;
        RECT 54.945 172.435 55.195 172.935 ;
        RECT 54.435 172.095 55.120 172.265 ;
        RECT 55.375 172.185 55.735 172.765 ;
        RECT 52.565 171.695 52.825 172.025 ;
        RECT 53.035 171.525 53.310 172.005 ;
        RECT 53.520 171.695 53.725 172.095 ;
        RECT 53.895 171.525 54.230 171.925 ;
        RECT 54.410 171.525 54.745 171.925 ;
        RECT 54.915 171.695 55.120 172.095 ;
        RECT 55.905 172.025 56.075 172.935 ;
        RECT 55.330 171.525 55.605 172.005 ;
        RECT 55.815 171.695 56.075 172.025 ;
        RECT 56.245 172.275 56.765 172.815 ;
        RECT 56.935 172.445 57.455 172.985 ;
        RECT 57.635 172.935 57.965 174.075 ;
        RECT 58.495 173.105 58.825 173.890 ;
        RECT 58.145 172.935 58.825 173.105 ;
        RECT 59.005 173.225 59.265 173.905 ;
        RECT 59.435 173.295 59.685 174.075 ;
        RECT 59.935 173.525 60.185 173.905 ;
        RECT 60.355 173.695 60.710 174.075 ;
        RECT 61.715 173.685 62.050 173.905 ;
        RECT 61.315 173.525 61.545 173.565 ;
        RECT 59.935 173.325 61.545 173.525 ;
        RECT 59.935 173.315 60.770 173.325 ;
        RECT 61.360 173.235 61.545 173.325 ;
        RECT 57.625 172.515 57.975 172.765 ;
        RECT 58.145 172.335 58.315 172.935 ;
        RECT 58.485 172.515 58.835 172.765 ;
        RECT 56.245 171.525 57.455 172.275 ;
        RECT 57.635 171.525 57.905 172.335 ;
        RECT 58.075 171.695 58.405 172.335 ;
        RECT 58.575 171.525 58.815 172.335 ;
        RECT 59.005 172.025 59.175 173.225 ;
        RECT 60.875 173.125 61.205 173.155 ;
        RECT 59.405 173.065 61.205 173.125 ;
        RECT 61.795 173.065 62.050 173.685 ;
        RECT 62.725 173.615 62.940 174.075 ;
        RECT 63.110 173.445 63.440 173.905 ;
        RECT 59.345 172.955 62.050 173.065 ;
        RECT 59.345 172.920 59.545 172.955 ;
        RECT 59.345 172.345 59.515 172.920 ;
        RECT 60.875 172.895 62.050 172.955 ;
        RECT 62.270 173.275 63.440 173.445 ;
        RECT 63.610 173.275 63.860 174.075 ;
        RECT 59.745 172.480 60.155 172.785 ;
        RECT 60.325 172.515 60.655 172.725 ;
        RECT 59.345 172.225 59.615 172.345 ;
        RECT 59.345 172.180 60.190 172.225 ;
        RECT 59.435 172.055 60.190 172.180 ;
        RECT 60.445 172.115 60.655 172.515 ;
        RECT 60.900 172.515 61.375 172.725 ;
        RECT 61.565 172.515 62.055 172.715 ;
        RECT 60.900 172.115 61.120 172.515 ;
        RECT 59.005 171.695 59.265 172.025 ;
        RECT 60.020 171.905 60.190 172.055 ;
        RECT 59.435 171.525 59.765 171.885 ;
        RECT 60.020 171.695 61.320 171.905 ;
        RECT 61.595 171.525 62.050 172.290 ;
        RECT 62.270 171.985 62.640 173.275 ;
        RECT 64.070 173.105 64.350 173.265 ;
        RECT 63.015 172.935 64.350 173.105 ;
        RECT 64.525 172.985 66.195 174.075 ;
        RECT 63.015 172.765 63.185 172.935 ;
        RECT 62.810 172.515 63.185 172.765 ;
        RECT 63.355 172.515 63.830 172.755 ;
        RECT 64.000 172.515 64.350 172.755 ;
        RECT 63.015 172.345 63.185 172.515 ;
        RECT 63.015 172.175 64.350 172.345 ;
        RECT 62.270 171.695 63.020 171.985 ;
        RECT 63.530 171.525 63.860 171.985 ;
        RECT 64.080 171.965 64.350 172.175 ;
        RECT 64.525 172.295 65.275 172.815 ;
        RECT 65.445 172.465 66.195 172.985 ;
        RECT 66.825 173.645 67.165 173.905 ;
        RECT 64.525 171.525 66.195 172.295 ;
        RECT 66.825 172.245 67.085 173.645 ;
        RECT 67.335 173.275 67.665 174.075 ;
        RECT 68.130 173.105 68.380 173.905 ;
        RECT 68.565 173.355 68.895 174.075 ;
        RECT 69.115 173.105 69.365 173.905 ;
        RECT 69.535 173.695 69.870 174.075 ;
        RECT 67.275 172.935 69.465 173.105 ;
        RECT 67.275 172.765 67.590 172.935 ;
        RECT 67.260 172.515 67.590 172.765 ;
        RECT 66.825 171.735 67.165 172.245 ;
        RECT 67.335 171.525 67.605 172.325 ;
        RECT 67.785 171.795 68.065 172.765 ;
        RECT 68.245 171.795 68.545 172.765 ;
        RECT 68.725 171.800 69.075 172.765 ;
        RECT 69.295 172.025 69.465 172.935 ;
        RECT 69.635 172.205 69.875 173.515 ;
        RECT 70.045 173.355 70.505 173.905 ;
        RECT 70.695 173.355 71.025 174.075 ;
        RECT 69.295 171.695 69.790 172.025 ;
        RECT 70.045 171.985 70.295 173.355 ;
        RECT 71.225 173.185 71.525 173.735 ;
        RECT 71.695 173.405 71.975 174.075 ;
        RECT 72.350 173.695 72.685 174.075 ;
        RECT 70.585 173.015 71.525 173.185 ;
        RECT 70.585 172.765 70.755 173.015 ;
        RECT 71.895 172.765 72.160 173.125 ;
        RECT 70.465 172.435 70.755 172.765 ;
        RECT 70.925 172.515 71.265 172.765 ;
        RECT 71.485 172.515 72.160 172.765 ;
        RECT 70.585 172.345 70.755 172.435 ;
        RECT 70.585 172.155 71.975 172.345 ;
        RECT 72.345 172.205 72.585 173.515 ;
        RECT 72.855 173.105 73.105 173.905 ;
        RECT 73.325 173.355 73.655 174.075 ;
        RECT 73.840 173.105 74.090 173.905 ;
        RECT 74.555 173.275 74.885 174.075 ;
        RECT 75.055 173.645 75.395 173.905 ;
        RECT 72.755 172.935 74.945 173.105 ;
        RECT 70.045 171.695 70.605 171.985 ;
        RECT 70.775 171.525 71.025 171.985 ;
        RECT 71.645 171.795 71.975 172.155 ;
        RECT 72.755 172.025 72.925 172.935 ;
        RECT 74.630 172.765 74.945 172.935 ;
        RECT 72.430 171.695 72.925 172.025 ;
        RECT 73.145 171.800 73.495 172.765 ;
        RECT 73.675 171.795 73.975 172.765 ;
        RECT 74.155 171.795 74.435 172.765 ;
        RECT 74.630 172.515 74.960 172.765 ;
        RECT 74.615 171.525 74.885 172.325 ;
        RECT 75.135 172.245 75.395 173.645 ;
        RECT 75.055 171.735 75.395 172.245 ;
        RECT 75.600 173.285 76.135 173.905 ;
        RECT 75.600 172.265 75.915 173.285 ;
        RECT 76.305 173.275 76.635 174.075 ;
        RECT 77.120 173.105 77.510 173.280 ;
        RECT 76.085 172.935 77.510 173.105 ;
        RECT 76.085 172.435 76.255 172.935 ;
        RECT 75.600 171.695 76.215 172.265 ;
        RECT 76.505 172.205 76.770 172.765 ;
        RECT 76.940 172.035 77.110 172.935 ;
        RECT 77.865 172.910 78.155 174.075 ;
        RECT 78.415 173.405 78.585 173.905 ;
        RECT 78.755 173.575 79.085 174.075 ;
        RECT 78.415 173.235 79.080 173.405 ;
        RECT 77.280 172.205 77.635 172.765 ;
        RECT 78.330 172.415 78.680 173.065 ;
        RECT 76.385 171.525 76.600 172.035 ;
        RECT 76.830 171.705 77.110 172.035 ;
        RECT 77.290 171.525 77.530 172.035 ;
        RECT 77.865 171.525 78.155 172.250 ;
        RECT 78.850 172.245 79.080 173.235 ;
        RECT 78.415 172.075 79.080 172.245 ;
        RECT 78.415 171.785 78.585 172.075 ;
        RECT 78.755 171.525 79.085 171.905 ;
        RECT 79.255 171.785 79.440 173.905 ;
        RECT 79.680 173.615 79.945 174.075 ;
        RECT 80.115 173.480 80.365 173.905 ;
        RECT 80.575 173.630 81.680 173.800 ;
        RECT 80.060 173.350 80.365 173.480 ;
        RECT 79.610 172.155 79.890 173.105 ;
        RECT 80.060 172.245 80.230 173.350 ;
        RECT 80.400 172.565 80.640 173.160 ;
        RECT 80.810 173.095 81.340 173.460 ;
        RECT 80.810 172.395 80.980 173.095 ;
        RECT 81.510 173.015 81.680 173.630 ;
        RECT 81.850 173.275 82.020 174.075 ;
        RECT 82.190 173.575 82.440 173.905 ;
        RECT 82.665 173.605 83.550 173.775 ;
        RECT 81.510 172.925 82.020 173.015 ;
        RECT 80.060 172.115 80.285 172.245 ;
        RECT 80.455 172.175 80.980 172.395 ;
        RECT 81.150 172.755 82.020 172.925 ;
        RECT 79.695 171.525 79.945 171.985 ;
        RECT 80.115 171.975 80.285 172.115 ;
        RECT 81.150 171.975 81.320 172.755 ;
        RECT 81.850 172.685 82.020 172.755 ;
        RECT 81.530 172.505 81.730 172.535 ;
        RECT 82.190 172.505 82.360 173.575 ;
        RECT 82.530 172.685 82.720 173.405 ;
        RECT 81.530 172.205 82.360 172.505 ;
        RECT 82.890 172.475 83.210 173.435 ;
        RECT 80.115 171.805 80.450 171.975 ;
        RECT 80.645 171.805 81.320 171.975 ;
        RECT 81.640 171.525 82.010 172.025 ;
        RECT 82.190 171.975 82.360 172.205 ;
        RECT 82.745 172.145 83.210 172.475 ;
        RECT 83.380 172.765 83.550 173.605 ;
        RECT 83.730 173.575 84.045 174.075 ;
        RECT 84.275 173.345 84.615 173.905 ;
        RECT 83.720 172.970 84.615 173.345 ;
        RECT 84.785 173.065 84.955 174.075 ;
        RECT 84.425 172.765 84.615 172.970 ;
        RECT 85.125 173.015 85.455 173.860 ;
        RECT 85.125 172.935 85.515 173.015 ;
        RECT 85.685 172.985 89.195 174.075 ;
        RECT 89.365 172.985 90.575 174.075 ;
        RECT 85.300 172.885 85.515 172.935 ;
        RECT 83.380 172.435 84.255 172.765 ;
        RECT 84.425 172.435 85.175 172.765 ;
        RECT 83.380 171.975 83.550 172.435 ;
        RECT 84.425 172.265 84.625 172.435 ;
        RECT 85.345 172.305 85.515 172.885 ;
        RECT 85.290 172.265 85.515 172.305 ;
        RECT 82.190 171.805 82.595 171.975 ;
        RECT 82.765 171.805 83.550 171.975 ;
        RECT 83.825 171.525 84.035 172.055 ;
        RECT 84.295 171.740 84.625 172.265 ;
        RECT 85.135 172.180 85.515 172.265 ;
        RECT 85.685 172.295 87.335 172.815 ;
        RECT 87.505 172.465 89.195 172.985 ;
        RECT 84.795 171.525 84.965 172.135 ;
        RECT 85.135 171.745 85.465 172.180 ;
        RECT 85.685 171.525 89.195 172.295 ;
        RECT 89.365 172.275 89.885 172.815 ;
        RECT 90.055 172.445 90.575 172.985 ;
        RECT 90.745 172.985 91.955 174.075 ;
        RECT 90.745 172.445 91.265 172.985 ;
        RECT 91.435 172.275 91.955 172.815 ;
        RECT 89.365 171.525 90.575 172.275 ;
        RECT 90.745 171.525 91.955 172.275 ;
        RECT 13.380 171.355 92.040 171.525 ;
        RECT 13.465 170.605 14.675 171.355 ;
        RECT 14.845 170.810 20.190 171.355 ;
        RECT 13.465 170.065 13.985 170.605 ;
        RECT 14.155 169.895 14.675 170.435 ;
        RECT 16.430 169.980 16.770 170.810 ;
        RECT 20.365 170.585 22.035 171.355 ;
        RECT 22.295 170.805 22.465 171.095 ;
        RECT 22.635 170.975 22.965 171.355 ;
        RECT 22.295 170.635 22.960 170.805 ;
        RECT 13.465 168.805 14.675 169.895 ;
        RECT 18.250 169.240 18.600 170.490 ;
        RECT 20.365 170.065 21.115 170.585 ;
        RECT 21.285 169.895 22.035 170.415 ;
        RECT 14.845 168.805 20.190 169.240 ;
        RECT 20.365 168.805 22.035 169.895 ;
        RECT 22.210 169.815 22.560 170.465 ;
        RECT 22.730 169.645 22.960 170.635 ;
        RECT 22.295 169.475 22.960 169.645 ;
        RECT 22.295 168.975 22.465 169.475 ;
        RECT 22.635 168.805 22.965 169.305 ;
        RECT 23.135 168.975 23.320 171.095 ;
        RECT 23.575 170.895 23.825 171.355 ;
        RECT 23.995 170.905 24.330 171.075 ;
        RECT 24.525 170.905 25.200 171.075 ;
        RECT 23.995 170.765 24.165 170.905 ;
        RECT 23.490 169.775 23.770 170.725 ;
        RECT 23.940 170.635 24.165 170.765 ;
        RECT 23.940 169.530 24.110 170.635 ;
        RECT 24.335 170.485 24.860 170.705 ;
        RECT 24.280 169.720 24.520 170.315 ;
        RECT 24.690 169.785 24.860 170.485 ;
        RECT 25.030 170.125 25.200 170.905 ;
        RECT 25.520 170.855 25.890 171.355 ;
        RECT 26.070 170.905 26.475 171.075 ;
        RECT 26.645 170.905 27.430 171.075 ;
        RECT 26.070 170.675 26.240 170.905 ;
        RECT 25.410 170.375 26.240 170.675 ;
        RECT 26.625 170.405 27.090 170.735 ;
        RECT 25.410 170.345 25.610 170.375 ;
        RECT 25.730 170.125 25.900 170.195 ;
        RECT 25.030 169.955 25.900 170.125 ;
        RECT 25.390 169.865 25.900 169.955 ;
        RECT 23.940 169.400 24.245 169.530 ;
        RECT 24.690 169.420 25.220 169.785 ;
        RECT 23.560 168.805 23.825 169.265 ;
        RECT 23.995 168.975 24.245 169.400 ;
        RECT 25.390 169.250 25.560 169.865 ;
        RECT 24.455 169.080 25.560 169.250 ;
        RECT 25.730 168.805 25.900 169.605 ;
        RECT 26.070 169.305 26.240 170.375 ;
        RECT 26.410 169.475 26.600 170.195 ;
        RECT 26.770 169.445 27.090 170.405 ;
        RECT 27.260 170.445 27.430 170.905 ;
        RECT 27.705 170.825 27.915 171.355 ;
        RECT 28.175 170.615 28.505 171.140 ;
        RECT 28.675 170.745 28.845 171.355 ;
        RECT 29.015 170.700 29.345 171.135 ;
        RECT 29.015 170.615 29.395 170.700 ;
        RECT 28.305 170.445 28.505 170.615 ;
        RECT 29.170 170.575 29.395 170.615 ;
        RECT 27.260 170.115 28.135 170.445 ;
        RECT 28.305 170.115 29.055 170.445 ;
        RECT 26.070 168.975 26.320 169.305 ;
        RECT 27.260 169.275 27.430 170.115 ;
        RECT 28.305 169.910 28.495 170.115 ;
        RECT 29.225 169.995 29.395 170.575 ;
        RECT 29.565 170.555 29.875 171.355 ;
        RECT 30.080 170.555 30.775 171.185 ;
        RECT 31.035 170.805 31.205 171.095 ;
        RECT 31.375 170.975 31.705 171.355 ;
        RECT 31.035 170.635 31.700 170.805 ;
        RECT 29.575 170.115 29.910 170.385 ;
        RECT 29.180 169.945 29.395 169.995 ;
        RECT 30.080 169.955 30.250 170.555 ;
        RECT 30.420 170.115 30.755 170.365 ;
        RECT 27.600 169.535 28.495 169.910 ;
        RECT 29.005 169.865 29.395 169.945 ;
        RECT 26.545 169.105 27.430 169.275 ;
        RECT 27.610 168.805 27.925 169.305 ;
        RECT 28.155 168.975 28.495 169.535 ;
        RECT 28.665 168.805 28.835 169.815 ;
        RECT 29.005 169.020 29.335 169.865 ;
        RECT 29.565 168.805 29.845 169.945 ;
        RECT 30.015 168.975 30.345 169.955 ;
        RECT 30.515 168.805 30.775 169.945 ;
        RECT 30.950 169.815 31.300 170.465 ;
        RECT 31.470 169.645 31.700 170.635 ;
        RECT 31.035 169.475 31.700 169.645 ;
        RECT 31.035 168.975 31.205 169.475 ;
        RECT 31.375 168.805 31.705 169.305 ;
        RECT 31.875 168.975 32.060 171.095 ;
        RECT 32.315 170.895 32.565 171.355 ;
        RECT 32.735 170.905 33.070 171.075 ;
        RECT 33.265 170.905 33.940 171.075 ;
        RECT 32.735 170.765 32.905 170.905 ;
        RECT 32.230 169.775 32.510 170.725 ;
        RECT 32.680 170.635 32.905 170.765 ;
        RECT 32.680 169.530 32.850 170.635 ;
        RECT 33.075 170.485 33.600 170.705 ;
        RECT 33.020 169.720 33.260 170.315 ;
        RECT 33.430 169.785 33.600 170.485 ;
        RECT 33.770 170.125 33.940 170.905 ;
        RECT 34.260 170.855 34.630 171.355 ;
        RECT 34.810 170.905 35.215 171.075 ;
        RECT 35.385 170.905 36.170 171.075 ;
        RECT 34.810 170.675 34.980 170.905 ;
        RECT 34.150 170.375 34.980 170.675 ;
        RECT 35.365 170.405 35.830 170.735 ;
        RECT 34.150 170.345 34.350 170.375 ;
        RECT 34.470 170.125 34.640 170.195 ;
        RECT 33.770 169.955 34.640 170.125 ;
        RECT 34.130 169.865 34.640 169.955 ;
        RECT 32.680 169.400 32.985 169.530 ;
        RECT 33.430 169.420 33.960 169.785 ;
        RECT 32.300 168.805 32.565 169.265 ;
        RECT 32.735 168.975 32.985 169.400 ;
        RECT 34.130 169.250 34.300 169.865 ;
        RECT 33.195 169.080 34.300 169.250 ;
        RECT 34.470 168.805 34.640 169.605 ;
        RECT 34.810 169.305 34.980 170.375 ;
        RECT 35.150 169.475 35.340 170.195 ;
        RECT 35.510 169.445 35.830 170.405 ;
        RECT 36.000 170.445 36.170 170.905 ;
        RECT 36.445 170.825 36.655 171.355 ;
        RECT 36.915 170.615 37.245 171.140 ;
        RECT 37.415 170.745 37.585 171.355 ;
        RECT 37.755 170.700 38.085 171.135 ;
        RECT 37.755 170.615 38.135 170.700 ;
        RECT 39.225 170.630 39.515 171.355 ;
        RECT 39.770 170.965 41.780 171.185 ;
        RECT 37.045 170.445 37.245 170.615 ;
        RECT 37.910 170.575 38.135 170.615 ;
        RECT 36.000 170.115 36.875 170.445 ;
        RECT 37.045 170.115 37.795 170.445 ;
        RECT 34.810 168.975 35.060 169.305 ;
        RECT 36.000 169.275 36.170 170.115 ;
        RECT 37.045 169.910 37.235 170.115 ;
        RECT 37.965 169.995 38.135 170.575 ;
        RECT 37.920 169.945 38.135 169.995 ;
        RECT 39.685 170.535 41.360 170.795 ;
        RECT 41.530 170.715 41.780 170.965 ;
        RECT 41.950 170.885 42.120 171.355 ;
        RECT 42.290 170.715 42.620 171.185 ;
        RECT 42.790 170.885 42.960 171.355 ;
        RECT 43.130 170.715 43.460 171.185 ;
        RECT 41.530 170.535 43.460 170.715 ;
        RECT 43.635 170.535 43.910 171.355 ;
        RECT 44.080 170.715 44.410 171.185 ;
        RECT 44.580 170.885 44.750 171.355 ;
        RECT 44.920 170.715 45.250 171.185 ;
        RECT 45.420 170.885 45.590 171.355 ;
        RECT 45.760 170.715 46.090 171.185 ;
        RECT 46.260 170.885 46.430 171.355 ;
        RECT 46.600 170.715 46.930 171.185 ;
        RECT 47.100 170.885 47.370 171.355 ;
        RECT 47.560 170.965 49.570 171.135 ;
        RECT 44.080 170.705 47.030 170.715 ;
        RECT 47.560 170.705 47.810 170.965 ;
        RECT 49.895 170.805 50.065 171.095 ;
        RECT 50.235 170.975 50.565 171.355 ;
        RECT 44.080 170.535 47.810 170.705 ;
        RECT 47.980 170.535 49.635 170.795 ;
        RECT 49.895 170.635 50.560 170.805 ;
        RECT 39.685 169.995 39.920 170.535 ;
        RECT 40.090 170.165 41.455 170.365 ;
        RECT 41.775 170.165 44.990 170.365 ;
        RECT 45.160 170.165 47.030 170.365 ;
        RECT 47.200 170.165 49.245 170.365 ;
        RECT 41.285 169.995 41.455 170.165 ;
        RECT 45.160 169.995 45.330 170.165 ;
        RECT 47.200 169.995 47.370 170.165 ;
        RECT 49.415 169.995 49.635 170.535 ;
        RECT 36.340 169.535 37.235 169.910 ;
        RECT 37.745 169.865 38.135 169.945 ;
        RECT 35.285 169.105 36.170 169.275 ;
        RECT 36.350 168.805 36.665 169.305 ;
        RECT 36.895 168.975 37.235 169.535 ;
        RECT 37.405 168.805 37.575 169.815 ;
        RECT 37.745 169.020 38.075 169.865 ;
        RECT 39.225 168.805 39.515 169.970 ;
        RECT 39.685 169.825 40.900 169.995 ;
        RECT 41.285 169.825 45.330 169.995 ;
        RECT 45.500 169.825 47.370 169.995 ;
        RECT 39.685 168.975 40.060 169.825 ;
        RECT 40.650 169.655 40.900 169.825 ;
        RECT 47.560 169.775 49.635 169.995 ;
        RECT 49.810 169.815 50.160 170.465 ;
        RECT 47.560 169.655 47.850 169.775 ;
        RECT 40.230 168.805 40.480 169.605 ;
        RECT 40.650 169.435 43.420 169.655 ;
        RECT 40.650 168.975 40.900 169.435 ;
        RECT 41.070 168.805 41.320 169.265 ;
        RECT 41.490 168.975 41.740 169.435 ;
        RECT 41.910 168.805 42.160 169.265 ;
        RECT 42.330 168.975 42.580 169.435 ;
        RECT 42.750 168.805 43.000 169.265 ;
        RECT 43.170 168.975 43.420 169.435 ;
        RECT 43.635 169.435 45.590 169.655 ;
        RECT 43.635 168.975 43.950 169.435 ;
        RECT 44.120 168.805 44.370 169.265 ;
        RECT 44.540 168.975 44.790 169.435 ;
        RECT 44.960 168.805 45.210 169.265 ;
        RECT 45.380 169.225 45.590 169.435 ;
        RECT 45.760 169.395 47.850 169.655 ;
        RECT 45.380 168.975 47.350 169.225 ;
        RECT 47.560 168.975 47.850 169.395 ;
        RECT 48.020 168.805 48.270 169.605 ;
        RECT 48.440 168.975 48.690 169.775 ;
        RECT 48.860 168.805 49.110 169.605 ;
        RECT 49.280 168.975 49.635 169.775 ;
        RECT 50.330 169.645 50.560 170.635 ;
        RECT 49.895 169.475 50.560 169.645 ;
        RECT 49.895 168.975 50.065 169.475 ;
        RECT 50.235 168.805 50.565 169.305 ;
        RECT 50.735 168.975 50.920 171.095 ;
        RECT 51.175 170.895 51.425 171.355 ;
        RECT 51.595 170.905 51.930 171.075 ;
        RECT 52.125 170.905 52.800 171.075 ;
        RECT 51.595 170.765 51.765 170.905 ;
        RECT 51.090 169.775 51.370 170.725 ;
        RECT 51.540 170.635 51.765 170.765 ;
        RECT 51.540 169.530 51.710 170.635 ;
        RECT 51.935 170.485 52.460 170.705 ;
        RECT 51.880 169.720 52.120 170.315 ;
        RECT 52.290 169.785 52.460 170.485 ;
        RECT 52.630 170.125 52.800 170.905 ;
        RECT 53.120 170.855 53.490 171.355 ;
        RECT 53.670 170.905 54.075 171.075 ;
        RECT 54.245 170.905 55.030 171.075 ;
        RECT 53.670 170.675 53.840 170.905 ;
        RECT 53.010 170.375 53.840 170.675 ;
        RECT 54.225 170.405 54.690 170.735 ;
        RECT 53.010 170.345 53.210 170.375 ;
        RECT 53.330 170.125 53.500 170.195 ;
        RECT 52.630 169.955 53.500 170.125 ;
        RECT 52.990 169.865 53.500 169.955 ;
        RECT 51.540 169.400 51.845 169.530 ;
        RECT 52.290 169.420 52.820 169.785 ;
        RECT 51.160 168.805 51.425 169.265 ;
        RECT 51.595 168.975 51.845 169.400 ;
        RECT 52.990 169.250 53.160 169.865 ;
        RECT 52.055 169.080 53.160 169.250 ;
        RECT 53.330 168.805 53.500 169.605 ;
        RECT 53.670 169.305 53.840 170.375 ;
        RECT 54.010 169.475 54.200 170.195 ;
        RECT 54.370 169.445 54.690 170.405 ;
        RECT 54.860 170.445 55.030 170.905 ;
        RECT 55.305 170.825 55.515 171.355 ;
        RECT 55.775 170.615 56.105 171.140 ;
        RECT 56.275 170.745 56.445 171.355 ;
        RECT 56.615 170.700 56.945 171.135 ;
        RECT 57.165 170.745 57.505 171.160 ;
        RECT 57.675 170.915 57.845 171.355 ;
        RECT 58.035 170.965 59.295 171.145 ;
        RECT 58.035 170.745 58.365 170.965 ;
        RECT 56.615 170.615 56.995 170.700 ;
        RECT 55.905 170.445 56.105 170.615 ;
        RECT 56.770 170.575 56.995 170.615 ;
        RECT 57.165 170.615 58.365 170.745 ;
        RECT 58.535 170.615 58.885 170.795 ;
        RECT 57.165 170.575 58.195 170.615 ;
        RECT 54.860 170.115 55.735 170.445 ;
        RECT 55.905 170.115 56.655 170.445 ;
        RECT 53.670 168.975 53.920 169.305 ;
        RECT 54.860 169.275 55.030 170.115 ;
        RECT 55.905 169.910 56.095 170.115 ;
        RECT 56.825 169.995 56.995 170.575 ;
        RECT 57.165 170.165 57.625 170.365 ;
        RECT 57.795 170.195 58.160 170.365 ;
        RECT 57.795 169.995 57.975 170.195 ;
        RECT 58.375 170.025 58.545 170.445 ;
        RECT 56.780 169.945 56.995 169.995 ;
        RECT 55.200 169.535 56.095 169.910 ;
        RECT 56.605 169.865 56.995 169.945 ;
        RECT 54.145 169.105 55.030 169.275 ;
        RECT 55.210 168.805 55.525 169.305 ;
        RECT 55.755 168.975 56.095 169.535 ;
        RECT 56.265 168.805 56.435 169.815 ;
        RECT 56.605 169.020 56.935 169.865 ;
        RECT 57.165 168.805 57.485 169.985 ;
        RECT 57.655 169.825 57.975 169.995 ;
        RECT 57.655 169.035 57.855 169.825 ;
        RECT 58.145 169.775 58.545 170.025 ;
        RECT 58.715 169.605 58.885 170.615 ;
        RECT 58.045 169.395 58.885 169.605 ;
        RECT 59.055 169.450 59.295 170.775 ;
        RECT 60.390 170.515 60.650 171.355 ;
        RECT 60.825 170.610 61.080 171.185 ;
        RECT 61.250 170.975 61.580 171.355 ;
        RECT 61.795 170.805 61.965 171.185 ;
        RECT 61.250 170.635 61.965 170.805 ;
        RECT 58.045 168.975 58.545 169.395 ;
        RECT 59.035 168.805 59.245 169.265 ;
        RECT 60.390 168.805 60.650 169.955 ;
        RECT 60.825 169.880 60.995 170.610 ;
        RECT 61.250 170.445 61.420 170.635 ;
        RECT 62.225 170.585 64.815 171.355 ;
        RECT 64.985 170.630 65.275 171.355 ;
        RECT 65.445 170.615 65.785 171.185 ;
        RECT 65.980 170.690 66.150 171.355 ;
        RECT 66.430 171.015 66.650 171.060 ;
        RECT 66.425 170.845 66.650 171.015 ;
        RECT 66.820 170.875 67.265 171.045 ;
        RECT 66.430 170.705 66.650 170.845 ;
        RECT 61.165 170.115 61.420 170.445 ;
        RECT 61.250 169.905 61.420 170.115 ;
        RECT 61.700 170.085 62.055 170.455 ;
        RECT 62.225 170.065 63.435 170.585 ;
        RECT 60.825 168.975 61.080 169.880 ;
        RECT 61.250 169.735 61.965 169.905 ;
        RECT 63.605 169.895 64.815 170.415 ;
        RECT 61.250 168.805 61.580 169.565 ;
        RECT 61.795 168.975 61.965 169.735 ;
        RECT 62.225 168.805 64.815 169.895 ;
        RECT 64.985 168.805 65.275 169.970 ;
        RECT 65.445 169.645 65.620 170.615 ;
        RECT 66.430 170.535 66.925 170.705 ;
        RECT 65.790 169.995 65.960 170.445 ;
        RECT 66.130 170.165 66.580 170.365 ;
        RECT 66.750 170.340 66.925 170.535 ;
        RECT 67.095 170.085 67.265 170.875 ;
        RECT 67.435 170.750 67.685 171.120 ;
        RECT 67.515 170.365 67.685 170.750 ;
        RECT 67.855 170.715 68.105 171.120 ;
        RECT 68.275 170.885 68.445 171.355 ;
        RECT 68.615 170.715 68.955 171.120 ;
        RECT 67.855 170.535 68.955 170.715 ;
        RECT 69.125 170.585 70.795 171.355 ;
        RECT 71.015 170.700 71.345 171.135 ;
        RECT 71.515 170.745 71.685 171.355 ;
        RECT 70.965 170.615 71.345 170.700 ;
        RECT 71.855 170.615 72.185 171.140 ;
        RECT 72.445 170.825 72.655 171.355 ;
        RECT 72.930 170.905 73.715 171.075 ;
        RECT 73.885 170.905 74.290 171.075 ;
        RECT 67.515 170.195 67.710 170.365 ;
        RECT 65.790 169.825 66.185 169.995 ;
        RECT 67.095 169.945 67.370 170.085 ;
        RECT 65.445 168.975 65.705 169.645 ;
        RECT 66.015 169.555 66.185 169.825 ;
        RECT 66.355 169.725 67.370 169.945 ;
        RECT 67.540 169.945 67.710 170.195 ;
        RECT 67.880 170.115 68.440 170.365 ;
        RECT 67.540 169.555 68.095 169.945 ;
        RECT 66.015 169.385 68.095 169.555 ;
        RECT 65.875 168.805 66.205 169.205 ;
        RECT 67.075 168.805 67.475 169.205 ;
        RECT 67.765 169.150 68.095 169.385 ;
        RECT 68.265 169.015 68.440 170.115 ;
        RECT 68.610 169.795 68.955 170.365 ;
        RECT 69.125 170.065 69.875 170.585 ;
        RECT 70.965 170.575 71.190 170.615 ;
        RECT 70.045 169.895 70.795 170.415 ;
        RECT 68.610 168.805 68.955 169.625 ;
        RECT 69.125 168.805 70.795 169.895 ;
        RECT 70.965 169.995 71.135 170.575 ;
        RECT 71.855 170.445 72.055 170.615 ;
        RECT 72.930 170.445 73.100 170.905 ;
        RECT 71.305 170.115 72.055 170.445 ;
        RECT 72.225 170.115 73.100 170.445 ;
        RECT 70.965 169.945 71.180 169.995 ;
        RECT 70.965 169.865 71.355 169.945 ;
        RECT 71.025 169.020 71.355 169.865 ;
        RECT 71.865 169.910 72.055 170.115 ;
        RECT 71.525 168.805 71.695 169.815 ;
        RECT 71.865 169.535 72.760 169.910 ;
        RECT 71.865 168.975 72.205 169.535 ;
        RECT 72.435 168.805 72.750 169.305 ;
        RECT 72.930 169.275 73.100 170.115 ;
        RECT 73.270 170.405 73.735 170.735 ;
        RECT 74.120 170.675 74.290 170.905 ;
        RECT 74.470 170.855 74.840 171.355 ;
        RECT 75.160 170.905 75.835 171.075 ;
        RECT 76.030 170.905 76.365 171.075 ;
        RECT 73.270 169.445 73.590 170.405 ;
        RECT 74.120 170.375 74.950 170.675 ;
        RECT 73.760 169.475 73.950 170.195 ;
        RECT 74.120 169.305 74.290 170.375 ;
        RECT 74.750 170.345 74.950 170.375 ;
        RECT 74.460 170.125 74.630 170.195 ;
        RECT 75.160 170.125 75.330 170.905 ;
        RECT 76.195 170.765 76.365 170.905 ;
        RECT 76.535 170.895 76.785 171.355 ;
        RECT 74.460 169.955 75.330 170.125 ;
        RECT 75.500 170.485 76.025 170.705 ;
        RECT 76.195 170.635 76.420 170.765 ;
        RECT 74.460 169.865 74.970 169.955 ;
        RECT 72.930 169.105 73.815 169.275 ;
        RECT 74.040 168.975 74.290 169.305 ;
        RECT 74.460 168.805 74.630 169.605 ;
        RECT 74.800 169.250 74.970 169.865 ;
        RECT 75.500 169.785 75.670 170.485 ;
        RECT 75.140 169.420 75.670 169.785 ;
        RECT 75.840 169.720 76.080 170.315 ;
        RECT 76.250 169.530 76.420 170.635 ;
        RECT 76.590 169.775 76.870 170.725 ;
        RECT 76.115 169.400 76.420 169.530 ;
        RECT 74.800 169.080 75.905 169.250 ;
        RECT 76.115 168.975 76.365 169.400 ;
        RECT 76.535 168.805 76.800 169.265 ;
        RECT 77.040 168.975 77.225 171.095 ;
        RECT 77.395 170.975 77.725 171.355 ;
        RECT 77.895 170.805 78.065 171.095 ;
        RECT 78.325 170.810 83.670 171.355 ;
        RECT 83.845 170.810 89.190 171.355 ;
        RECT 77.400 170.635 78.065 170.805 ;
        RECT 77.400 169.645 77.630 170.635 ;
        RECT 77.800 169.815 78.150 170.465 ;
        RECT 79.910 169.980 80.250 170.810 ;
        RECT 77.400 169.475 78.065 169.645 ;
        RECT 77.395 168.805 77.725 169.305 ;
        RECT 77.895 168.975 78.065 169.475 ;
        RECT 81.730 169.240 82.080 170.490 ;
        RECT 85.430 169.980 85.770 170.810 ;
        RECT 89.365 170.605 90.575 171.355 ;
        RECT 90.745 170.605 91.955 171.355 ;
        RECT 87.250 169.240 87.600 170.490 ;
        RECT 89.365 170.065 89.885 170.605 ;
        RECT 90.055 169.895 90.575 170.435 ;
        RECT 78.325 168.805 83.670 169.240 ;
        RECT 83.845 168.805 89.190 169.240 ;
        RECT 89.365 168.805 90.575 169.895 ;
        RECT 90.745 169.895 91.265 170.435 ;
        RECT 91.435 170.065 91.955 170.605 ;
        RECT 100.140 170.940 100.810 174.200 ;
        RECT 101.480 173.630 105.520 173.800 ;
        RECT 101.140 171.570 101.310 173.570 ;
        RECT 105.690 171.570 105.860 173.570 ;
        RECT 101.480 171.340 105.520 171.510 ;
        RECT 106.200 170.940 106.370 174.200 ;
        RECT 100.140 170.770 106.370 170.940 ;
        RECT 90.745 168.805 91.955 169.895 ;
        RECT 13.380 168.635 92.040 168.805 ;
        RECT 13.465 167.545 14.675 168.635 ;
        RECT 14.845 168.200 20.190 168.635 ;
        RECT 13.465 166.835 13.985 167.375 ;
        RECT 14.155 167.005 14.675 167.545 ;
        RECT 13.465 166.085 14.675 166.835 ;
        RECT 16.430 166.630 16.770 167.460 ;
        RECT 18.250 166.950 18.600 168.200 ;
        RECT 20.365 167.545 22.035 168.635 ;
        RECT 20.365 166.855 21.115 167.375 ;
        RECT 21.285 167.025 22.035 167.545 ;
        RECT 22.665 167.765 22.940 168.465 ;
        RECT 23.150 168.090 23.365 168.635 ;
        RECT 23.535 168.125 24.010 168.465 ;
        RECT 24.180 168.130 24.795 168.635 ;
        RECT 24.180 167.955 24.375 168.130 ;
        RECT 14.845 166.085 20.190 166.630 ;
        RECT 20.365 166.085 22.035 166.855 ;
        RECT 22.665 166.735 22.835 167.765 ;
        RECT 23.110 167.595 23.825 167.890 ;
        RECT 24.045 167.765 24.375 167.955 ;
        RECT 24.545 167.595 24.795 167.960 ;
        RECT 23.005 167.425 24.795 167.595 ;
        RECT 23.005 166.995 23.235 167.425 ;
        RECT 22.665 166.255 22.925 166.735 ;
        RECT 23.405 166.725 23.815 167.245 ;
        RECT 23.095 166.085 23.425 166.545 ;
        RECT 23.615 166.305 23.815 166.725 ;
        RECT 23.985 166.570 24.240 167.425 ;
        RECT 25.035 167.245 25.205 168.465 ;
        RECT 25.455 168.125 25.715 168.635 ;
        RECT 24.410 166.995 25.205 167.245 ;
        RECT 25.375 167.075 25.715 167.955 ;
        RECT 26.345 167.470 26.635 168.635 ;
        RECT 24.955 166.905 25.205 166.995 ;
        RECT 23.985 166.305 24.775 166.570 ;
        RECT 24.955 166.485 25.285 166.905 ;
        RECT 25.455 166.085 25.715 166.905 ;
        RECT 26.345 166.085 26.635 166.810 ;
        RECT 26.815 166.265 27.075 168.455 ;
        RECT 27.245 167.905 27.585 168.635 ;
        RECT 27.765 167.725 28.035 168.455 ;
        RECT 27.265 167.505 28.035 167.725 ;
        RECT 28.215 167.745 28.445 168.455 ;
        RECT 28.615 167.925 28.945 168.635 ;
        RECT 29.115 167.745 29.375 168.455 ;
        RECT 29.735 167.835 29.990 168.635 ;
        RECT 28.215 167.505 29.375 167.745 ;
        RECT 30.160 167.665 30.490 168.465 ;
        RECT 30.660 167.835 30.830 168.635 ;
        RECT 31.000 167.665 31.330 168.465 ;
        RECT 31.500 167.835 31.670 168.635 ;
        RECT 31.840 167.665 32.170 168.465 ;
        RECT 32.340 167.835 32.510 168.635 ;
        RECT 32.680 167.665 33.010 168.465 ;
        RECT 33.180 167.835 33.480 168.635 ;
        RECT 27.265 166.835 27.555 167.505 ;
        RECT 29.565 167.495 33.535 167.665 ;
        RECT 33.705 167.545 35.375 168.635 ;
        RECT 27.735 167.015 28.200 167.325 ;
        RECT 28.380 167.015 28.905 167.325 ;
        RECT 27.265 166.635 28.495 166.835 ;
        RECT 27.335 166.085 28.005 166.455 ;
        RECT 28.185 166.265 28.495 166.635 ;
        RECT 28.675 166.375 28.905 167.015 ;
        RECT 29.085 166.995 29.385 167.325 ;
        RECT 29.565 166.905 29.910 167.495 ;
        RECT 30.160 167.075 33.015 167.325 ;
        RECT 33.215 166.905 33.535 167.495 ;
        RECT 29.085 166.085 29.375 166.815 ;
        RECT 29.565 166.715 33.535 166.905 ;
        RECT 33.705 166.855 34.455 167.375 ;
        RECT 34.625 167.025 35.375 167.545 ;
        RECT 35.730 167.665 36.120 167.840 ;
        RECT 36.605 167.835 36.935 168.635 ;
        RECT 37.105 167.845 37.640 168.465 ;
        RECT 35.730 167.495 37.155 167.665 ;
        RECT 29.735 166.085 29.990 166.545 ;
        RECT 30.160 166.255 30.490 166.715 ;
        RECT 30.660 166.085 30.830 166.545 ;
        RECT 31.000 166.255 31.330 166.715 ;
        RECT 31.500 166.085 31.670 166.545 ;
        RECT 31.840 166.255 32.170 166.715 ;
        RECT 32.340 166.085 32.510 166.545 ;
        RECT 32.680 166.255 33.010 166.715 ;
        RECT 33.180 166.085 33.485 166.545 ;
        RECT 33.705 166.085 35.375 166.855 ;
        RECT 35.605 166.765 35.960 167.325 ;
        RECT 36.130 166.595 36.300 167.495 ;
        RECT 36.470 166.765 36.735 167.325 ;
        RECT 36.985 166.995 37.155 167.495 ;
        RECT 37.325 166.825 37.640 167.845 ;
        RECT 37.890 167.495 38.185 168.635 ;
        RECT 38.445 167.665 38.775 168.465 ;
        RECT 38.945 167.835 39.115 168.635 ;
        RECT 39.285 167.665 39.615 168.465 ;
        RECT 39.785 167.835 39.955 168.635 ;
        RECT 40.125 167.685 40.455 168.465 ;
        RECT 40.625 168.175 40.795 168.635 ;
        RECT 41.155 167.965 41.325 168.465 ;
        RECT 41.495 168.135 41.825 168.635 ;
        RECT 41.155 167.795 41.820 167.965 ;
        RECT 40.125 167.665 40.895 167.685 ;
        RECT 38.445 167.495 40.895 167.665 ;
        RECT 37.865 167.075 40.375 167.325 ;
        RECT 40.545 166.905 40.895 167.495 ;
        RECT 41.070 166.975 41.420 167.625 ;
        RECT 35.710 166.085 35.950 166.595 ;
        RECT 36.130 166.265 36.410 166.595 ;
        RECT 36.640 166.085 36.855 166.595 ;
        RECT 37.025 166.255 37.640 166.825 ;
        RECT 38.525 166.725 40.895 166.905 ;
        RECT 41.590 166.805 41.820 167.795 ;
        RECT 37.890 166.085 38.155 166.545 ;
        RECT 38.525 166.255 38.695 166.725 ;
        RECT 38.945 166.085 39.115 166.545 ;
        RECT 39.365 166.255 39.535 166.725 ;
        RECT 39.785 166.085 39.955 166.545 ;
        RECT 40.205 166.255 40.375 166.725 ;
        RECT 41.155 166.635 41.820 166.805 ;
        RECT 40.545 166.085 40.795 166.550 ;
        RECT 41.155 166.345 41.325 166.635 ;
        RECT 41.495 166.085 41.825 166.465 ;
        RECT 41.995 166.345 42.180 168.465 ;
        RECT 42.420 168.175 42.685 168.635 ;
        RECT 42.855 168.040 43.105 168.465 ;
        RECT 43.315 168.190 44.420 168.360 ;
        RECT 42.800 167.910 43.105 168.040 ;
        RECT 42.350 166.715 42.630 167.665 ;
        RECT 42.800 166.805 42.970 167.910 ;
        RECT 43.140 167.125 43.380 167.720 ;
        RECT 43.550 167.655 44.080 168.020 ;
        RECT 43.550 166.955 43.720 167.655 ;
        RECT 44.250 167.575 44.420 168.190 ;
        RECT 44.590 167.835 44.760 168.635 ;
        RECT 44.930 168.135 45.180 168.465 ;
        RECT 45.405 168.165 46.290 168.335 ;
        RECT 44.250 167.485 44.760 167.575 ;
        RECT 42.800 166.675 43.025 166.805 ;
        RECT 43.195 166.735 43.720 166.955 ;
        RECT 43.890 167.315 44.760 167.485 ;
        RECT 42.435 166.085 42.685 166.545 ;
        RECT 42.855 166.535 43.025 166.675 ;
        RECT 43.890 166.535 44.060 167.315 ;
        RECT 44.590 167.245 44.760 167.315 ;
        RECT 44.270 167.065 44.470 167.095 ;
        RECT 44.930 167.065 45.100 168.135 ;
        RECT 45.270 167.245 45.460 167.965 ;
        RECT 44.270 166.765 45.100 167.065 ;
        RECT 45.630 167.035 45.950 167.995 ;
        RECT 42.855 166.365 43.190 166.535 ;
        RECT 43.385 166.365 44.060 166.535 ;
        RECT 44.380 166.085 44.750 166.585 ;
        RECT 44.930 166.535 45.100 166.765 ;
        RECT 45.485 166.705 45.950 167.035 ;
        RECT 46.120 167.325 46.290 168.165 ;
        RECT 46.470 168.135 46.785 168.635 ;
        RECT 47.015 167.905 47.355 168.465 ;
        RECT 46.460 167.530 47.355 167.905 ;
        RECT 47.525 167.625 47.695 168.635 ;
        RECT 47.165 167.325 47.355 167.530 ;
        RECT 47.865 167.575 48.195 168.420 ;
        RECT 48.630 167.665 48.960 168.465 ;
        RECT 49.130 167.835 49.460 168.635 ;
        RECT 49.760 167.665 50.090 168.465 ;
        RECT 50.735 167.835 50.985 168.635 ;
        RECT 47.865 167.495 48.255 167.575 ;
        RECT 48.630 167.495 51.065 167.665 ;
        RECT 51.255 167.495 51.425 168.635 ;
        RECT 51.595 167.495 51.935 168.465 ;
        RECT 48.040 167.445 48.255 167.495 ;
        RECT 46.120 166.995 46.995 167.325 ;
        RECT 47.165 166.995 47.915 167.325 ;
        RECT 46.120 166.535 46.290 166.995 ;
        RECT 47.165 166.825 47.365 166.995 ;
        RECT 48.085 166.865 48.255 167.445 ;
        RECT 48.425 167.075 48.775 167.325 ;
        RECT 48.960 166.865 49.130 167.495 ;
        RECT 49.300 167.075 49.630 167.275 ;
        RECT 49.800 167.075 50.130 167.275 ;
        RECT 50.300 167.075 50.720 167.275 ;
        RECT 50.895 167.245 51.065 167.495 ;
        RECT 50.895 167.075 51.590 167.245 ;
        RECT 48.030 166.825 48.255 166.865 ;
        RECT 44.930 166.365 45.335 166.535 ;
        RECT 45.505 166.365 46.290 166.535 ;
        RECT 46.565 166.085 46.775 166.615 ;
        RECT 47.035 166.300 47.365 166.825 ;
        RECT 47.875 166.740 48.255 166.825 ;
        RECT 47.535 166.085 47.705 166.695 ;
        RECT 47.875 166.305 48.205 166.740 ;
        RECT 48.630 166.255 49.130 166.865 ;
        RECT 49.760 166.735 50.985 166.905 ;
        RECT 51.760 166.885 51.935 167.495 ;
        RECT 52.105 167.470 52.395 168.635 ;
        RECT 52.565 167.495 52.845 168.635 ;
        RECT 53.015 167.485 53.345 168.465 ;
        RECT 53.515 167.495 53.775 168.635 ;
        RECT 53.985 167.495 54.215 168.635 ;
        RECT 54.385 167.485 54.715 168.465 ;
        RECT 54.885 167.495 55.095 168.635 ;
        RECT 55.415 168.015 55.585 168.445 ;
        RECT 55.755 168.185 56.085 168.635 ;
        RECT 55.415 167.785 56.090 168.015 ;
        RECT 52.575 167.055 52.910 167.325 ;
        RECT 53.080 166.885 53.250 167.485 ;
        RECT 53.420 167.075 53.755 167.325 ;
        RECT 53.965 167.075 54.295 167.325 ;
        RECT 49.760 166.255 50.090 166.735 ;
        RECT 50.260 166.085 50.485 166.545 ;
        RECT 50.655 166.255 50.985 166.735 ;
        RECT 51.175 166.085 51.425 166.885 ;
        RECT 51.595 166.255 51.935 166.885 ;
        RECT 52.105 166.085 52.395 166.810 ;
        RECT 52.565 166.085 52.875 166.885 ;
        RECT 53.080 166.255 53.775 166.885 ;
        RECT 53.985 166.085 54.215 166.905 ;
        RECT 54.465 166.885 54.715 167.485 ;
        RECT 54.385 166.255 54.715 166.885 ;
        RECT 54.885 166.085 55.095 166.905 ;
        RECT 55.385 166.765 55.685 167.615 ;
        RECT 55.855 167.135 56.090 167.785 ;
        RECT 56.260 167.475 56.545 168.420 ;
        RECT 56.725 168.165 57.410 168.635 ;
        RECT 56.720 167.645 57.415 167.955 ;
        RECT 57.590 167.580 57.895 168.365 ;
        RECT 56.260 167.325 57.120 167.475 ;
        RECT 57.685 167.445 57.895 167.580 ;
        RECT 58.095 167.525 58.390 168.635 ;
        RECT 56.260 167.305 57.545 167.325 ;
        RECT 55.855 166.805 56.390 167.135 ;
        RECT 56.560 166.945 57.545 167.305 ;
        RECT 55.855 166.655 56.075 166.805 ;
        RECT 55.330 166.085 55.665 166.590 ;
        RECT 55.835 166.280 56.075 166.655 ;
        RECT 56.560 166.610 56.730 166.945 ;
        RECT 57.720 166.775 57.895 167.445 ;
        RECT 58.570 167.325 58.820 168.460 ;
        RECT 58.990 167.525 59.250 168.635 ;
        RECT 59.420 167.735 59.680 168.460 ;
        RECT 59.850 167.905 60.110 168.635 ;
        RECT 60.280 167.735 60.540 168.460 ;
        RECT 60.710 167.905 60.970 168.635 ;
        RECT 61.140 167.735 61.400 168.460 ;
        RECT 61.570 167.905 61.830 168.635 ;
        RECT 62.000 167.735 62.260 168.460 ;
        RECT 62.430 167.905 62.725 168.635 ;
        RECT 63.145 167.785 63.525 168.465 ;
        RECT 64.115 167.785 64.285 168.635 ;
        RECT 64.455 167.955 64.785 168.465 ;
        RECT 64.955 168.125 65.125 168.635 ;
        RECT 65.295 167.955 65.695 168.465 ;
        RECT 64.455 167.785 65.695 167.955 ;
        RECT 59.420 167.495 62.730 167.735 ;
        RECT 56.355 166.415 56.730 166.610 ;
        RECT 56.355 166.270 56.525 166.415 ;
        RECT 57.090 166.085 57.485 166.580 ;
        RECT 57.655 166.255 57.895 166.775 ;
        RECT 58.085 166.715 58.400 167.325 ;
        RECT 58.570 167.075 61.590 167.325 ;
        RECT 58.145 166.085 58.390 166.545 ;
        RECT 58.570 166.265 58.820 167.075 ;
        RECT 61.760 166.905 62.730 167.495 ;
        RECT 59.420 166.735 62.730 166.905 ;
        RECT 63.145 166.825 63.315 167.785 ;
        RECT 63.485 167.445 64.790 167.615 ;
        RECT 65.875 167.535 66.195 168.465 ;
        RECT 66.365 167.545 68.035 168.635 ;
        RECT 63.485 166.995 63.730 167.445 ;
        RECT 63.900 167.075 64.450 167.275 ;
        RECT 64.620 167.245 64.790 167.445 ;
        RECT 65.565 167.365 66.195 167.535 ;
        RECT 64.620 167.075 64.995 167.245 ;
        RECT 65.165 166.825 65.395 167.325 ;
        RECT 58.990 166.085 59.250 166.610 ;
        RECT 59.420 166.280 59.680 166.735 ;
        RECT 59.850 166.085 60.110 166.565 ;
        RECT 60.280 166.280 60.540 166.735 ;
        RECT 60.710 166.085 60.970 166.565 ;
        RECT 61.140 166.280 61.400 166.735 ;
        RECT 61.570 166.085 61.830 166.565 ;
        RECT 62.000 166.280 62.260 166.735 ;
        RECT 63.145 166.655 65.395 166.825 ;
        RECT 62.430 166.085 62.730 166.565 ;
        RECT 63.195 166.085 63.525 166.475 ;
        RECT 63.695 166.335 63.865 166.655 ;
        RECT 65.565 166.485 65.735 167.365 ;
        RECT 64.035 166.085 64.365 166.475 ;
        RECT 64.780 166.315 65.735 166.485 ;
        RECT 65.905 166.085 66.195 166.920 ;
        RECT 66.365 166.855 67.115 167.375 ;
        RECT 67.285 167.025 68.035 167.545 ;
        RECT 68.710 167.495 69.005 168.635 ;
        RECT 69.265 167.665 69.595 168.465 ;
        RECT 69.765 167.835 69.935 168.635 ;
        RECT 70.105 167.665 70.435 168.465 ;
        RECT 70.605 167.835 70.775 168.635 ;
        RECT 70.945 167.685 71.275 168.465 ;
        RECT 71.445 168.175 71.615 168.635 ;
        RECT 71.885 167.765 72.160 168.465 ;
        RECT 72.330 168.090 72.585 168.635 ;
        RECT 72.755 168.125 73.235 168.465 ;
        RECT 73.410 168.080 74.015 168.635 ;
        RECT 73.400 167.980 74.015 168.080 ;
        RECT 73.400 167.955 73.585 167.980 ;
        RECT 70.945 167.665 71.715 167.685 ;
        RECT 69.265 167.495 71.715 167.665 ;
        RECT 68.685 167.075 71.195 167.325 ;
        RECT 71.365 166.905 71.715 167.495 ;
        RECT 66.365 166.085 68.035 166.855 ;
        RECT 69.345 166.725 71.715 166.905 ;
        RECT 71.885 166.735 72.055 167.765 ;
        RECT 72.330 167.635 73.085 167.885 ;
        RECT 73.255 167.710 73.585 167.955 ;
        RECT 72.330 167.600 73.100 167.635 ;
        RECT 72.330 167.590 73.115 167.600 ;
        RECT 72.225 167.575 73.120 167.590 ;
        RECT 72.225 167.560 73.140 167.575 ;
        RECT 72.225 167.550 73.160 167.560 ;
        RECT 72.225 167.540 73.185 167.550 ;
        RECT 72.225 167.510 73.255 167.540 ;
        RECT 72.225 167.480 73.275 167.510 ;
        RECT 72.225 167.450 73.295 167.480 ;
        RECT 72.225 167.425 73.325 167.450 ;
        RECT 72.225 167.390 73.360 167.425 ;
        RECT 72.225 167.385 73.390 167.390 ;
        RECT 72.225 166.990 72.455 167.385 ;
        RECT 73.000 167.380 73.390 167.385 ;
        RECT 73.025 167.370 73.390 167.380 ;
        RECT 73.040 167.365 73.390 167.370 ;
        RECT 73.055 167.360 73.390 167.365 ;
        RECT 73.755 167.360 74.015 167.810 ;
        RECT 74.185 167.545 77.695 168.635 ;
        RECT 73.055 167.355 74.015 167.360 ;
        RECT 73.065 167.345 74.015 167.355 ;
        RECT 73.075 167.340 74.015 167.345 ;
        RECT 73.085 167.330 74.015 167.340 ;
        RECT 73.090 167.320 74.015 167.330 ;
        RECT 73.095 167.315 74.015 167.320 ;
        RECT 73.105 167.300 74.015 167.315 ;
        RECT 73.110 167.285 74.015 167.300 ;
        RECT 73.120 167.260 74.015 167.285 ;
        RECT 72.625 166.790 72.955 167.215 ;
        RECT 72.705 166.765 72.955 166.790 ;
        RECT 68.710 166.085 68.975 166.545 ;
        RECT 69.345 166.255 69.515 166.725 ;
        RECT 69.765 166.085 69.935 166.545 ;
        RECT 70.185 166.255 70.355 166.725 ;
        RECT 70.605 166.085 70.775 166.545 ;
        RECT 71.025 166.255 71.195 166.725 ;
        RECT 71.365 166.085 71.615 166.550 ;
        RECT 71.885 166.255 72.145 166.735 ;
        RECT 72.315 166.085 72.565 166.625 ;
        RECT 72.735 166.305 72.955 166.765 ;
        RECT 73.125 167.190 74.015 167.260 ;
        RECT 73.125 166.465 73.295 167.190 ;
        RECT 73.465 166.635 74.015 167.020 ;
        RECT 74.185 166.855 75.835 167.375 ;
        RECT 76.005 167.025 77.695 167.545 ;
        RECT 77.865 167.470 78.155 168.635 ;
        RECT 78.325 168.200 83.670 168.635 ;
        RECT 83.845 168.200 89.190 168.635 ;
        RECT 73.125 166.295 74.015 166.465 ;
        RECT 74.185 166.085 77.695 166.855 ;
        RECT 77.865 166.085 78.155 166.810 ;
        RECT 79.910 166.630 80.250 167.460 ;
        RECT 81.730 166.950 82.080 168.200 ;
        RECT 85.430 166.630 85.770 167.460 ;
        RECT 87.250 166.950 87.600 168.200 ;
        RECT 89.365 167.545 90.575 168.635 ;
        RECT 89.365 166.835 89.885 167.375 ;
        RECT 90.055 167.005 90.575 167.545 ;
        RECT 90.745 167.545 91.955 168.635 ;
        RECT 90.745 167.005 91.265 167.545 ;
        RECT 100.140 167.510 100.810 170.770 ;
        RECT 101.480 170.200 105.520 170.370 ;
        RECT 101.140 168.140 101.310 170.140 ;
        RECT 105.690 168.140 105.860 170.140 ;
        RECT 101.480 167.910 105.520 168.080 ;
        RECT 106.200 167.510 106.370 170.770 ;
        RECT 100.140 167.500 106.370 167.510 ;
        RECT 107.960 176.770 117.790 176.810 ;
        RECT 140.540 176.790 146.280 176.800 ;
        RECT 107.960 176.640 118.590 176.770 ;
        RECT 120.510 176.740 126.250 176.750 ;
        RECT 107.960 174.380 108.130 176.640 ;
        RECT 108.855 176.070 116.895 176.240 ;
        RECT 108.470 175.010 108.640 176.010 ;
        RECT 117.110 175.010 117.280 176.010 ;
        RECT 108.855 174.780 116.895 174.950 ;
        RECT 117.620 174.380 118.590 176.640 ;
        RECT 107.960 174.210 118.590 174.380 ;
        RECT 107.960 170.950 108.130 174.210 ;
        RECT 108.855 173.640 116.895 173.810 ;
        RECT 108.470 171.580 108.640 173.580 ;
        RECT 117.110 171.580 117.280 173.580 ;
        RECT 108.855 171.350 116.895 171.520 ;
        RECT 117.620 170.950 118.590 174.210 ;
        RECT 107.960 170.780 118.590 170.950 ;
        RECT 107.960 167.520 108.130 170.780 ;
        RECT 108.855 170.210 116.895 170.380 ;
        RECT 108.470 168.150 108.640 170.150 ;
        RECT 117.110 168.150 117.280 170.150 ;
        RECT 108.855 167.920 116.895 168.090 ;
        RECT 117.620 167.520 118.590 170.780 ;
        RECT 100.140 167.400 106.380 167.500 ;
        RECT 91.435 166.835 91.955 167.375 ;
        RECT 78.325 166.085 83.670 166.630 ;
        RECT 83.845 166.085 89.190 166.630 ;
        RECT 89.365 166.085 90.575 166.835 ;
        RECT 90.745 166.085 91.955 166.835 ;
        RECT 100.130 166.840 106.380 167.400 ;
        RECT 100.130 166.820 105.300 166.840 ;
        RECT 100.130 166.750 104.120 166.820 ;
        RECT 13.380 165.915 92.040 166.085 ;
        RECT 13.465 165.165 14.675 165.915 ;
        RECT 14.845 165.370 20.190 165.915 ;
        RECT 13.465 164.625 13.985 165.165 ;
        RECT 14.155 164.455 14.675 164.995 ;
        RECT 16.430 164.540 16.770 165.370 ;
        RECT 20.365 165.145 23.875 165.915 ;
        RECT 24.210 165.405 24.450 165.915 ;
        RECT 24.630 165.405 24.910 165.735 ;
        RECT 25.140 165.405 25.355 165.915 ;
        RECT 13.465 163.365 14.675 164.455 ;
        RECT 18.250 163.800 18.600 165.050 ;
        RECT 20.365 164.625 22.015 165.145 ;
        RECT 22.185 164.455 23.875 164.975 ;
        RECT 24.105 164.675 24.460 165.235 ;
        RECT 24.630 164.505 24.800 165.405 ;
        RECT 24.970 164.675 25.235 165.235 ;
        RECT 25.525 165.175 26.140 165.745 ;
        RECT 25.485 164.505 25.655 165.005 ;
        RECT 14.845 163.365 20.190 163.800 ;
        RECT 20.365 163.365 23.875 164.455 ;
        RECT 24.230 164.335 25.655 164.505 ;
        RECT 24.230 164.160 24.620 164.335 ;
        RECT 25.105 163.365 25.435 164.165 ;
        RECT 25.825 164.155 26.140 165.175 ;
        RECT 25.605 163.535 26.140 164.155 ;
        RECT 26.345 165.195 26.685 165.705 ;
        RECT 26.345 163.795 26.605 165.195 ;
        RECT 26.855 165.115 27.125 165.915 ;
        RECT 26.780 164.675 27.110 164.925 ;
        RECT 27.305 164.675 27.585 165.645 ;
        RECT 27.765 164.675 28.065 165.645 ;
        RECT 28.245 164.675 28.595 165.640 ;
        RECT 28.815 165.415 29.310 165.745 ;
        RECT 29.810 165.435 30.110 165.915 ;
        RECT 26.795 164.505 27.110 164.675 ;
        RECT 28.815 164.505 28.985 165.415 ;
        RECT 30.280 165.265 30.540 165.720 ;
        RECT 30.710 165.435 30.970 165.915 ;
        RECT 31.140 165.265 31.400 165.720 ;
        RECT 31.570 165.435 31.830 165.915 ;
        RECT 32.000 165.265 32.260 165.720 ;
        RECT 32.430 165.435 32.690 165.915 ;
        RECT 32.860 165.265 33.120 165.720 ;
        RECT 33.290 165.390 33.550 165.915 ;
        RECT 26.795 164.335 28.985 164.505 ;
        RECT 26.345 163.535 26.685 163.795 ;
        RECT 26.855 163.365 27.185 164.165 ;
        RECT 27.650 163.535 27.900 164.335 ;
        RECT 28.085 163.365 28.415 164.085 ;
        RECT 28.635 163.535 28.885 164.335 ;
        RECT 29.155 163.925 29.395 165.235 ;
        RECT 29.810 165.095 33.120 165.265 ;
        RECT 29.810 164.505 30.780 165.095 ;
        RECT 33.720 164.925 33.970 165.735 ;
        RECT 34.150 165.455 34.395 165.915 ;
        RECT 30.950 164.675 33.970 164.925 ;
        RECT 34.140 164.675 34.455 165.285 ;
        RECT 29.810 164.265 33.120 164.505 ;
        RECT 29.055 163.365 29.390 163.745 ;
        RECT 29.815 163.365 30.110 164.095 ;
        RECT 30.280 163.540 30.540 164.265 ;
        RECT 30.710 163.365 30.970 164.095 ;
        RECT 31.140 163.540 31.400 164.265 ;
        RECT 31.570 163.365 31.830 164.095 ;
        RECT 32.000 163.540 32.260 164.265 ;
        RECT 32.430 163.365 32.690 164.095 ;
        RECT 32.860 163.540 33.120 164.265 ;
        RECT 33.290 163.365 33.550 164.475 ;
        RECT 33.720 163.540 33.970 164.675 ;
        RECT 34.150 163.365 34.445 164.475 ;
        RECT 34.635 163.545 34.895 165.735 ;
        RECT 35.155 165.545 35.825 165.915 ;
        RECT 36.005 165.365 36.315 165.735 ;
        RECT 35.085 165.165 36.315 165.365 ;
        RECT 35.085 164.495 35.375 165.165 ;
        RECT 36.495 164.985 36.725 165.625 ;
        RECT 36.905 165.185 37.195 165.915 ;
        RECT 37.385 165.145 39.055 165.915 ;
        RECT 39.225 165.190 39.515 165.915 ;
        RECT 39.685 165.370 45.030 165.915 ;
        RECT 45.205 165.370 50.550 165.915 ;
        RECT 50.725 165.370 56.070 165.915 ;
        RECT 35.555 164.675 36.020 164.985 ;
        RECT 36.200 164.675 36.725 164.985 ;
        RECT 36.905 164.675 37.205 165.005 ;
        RECT 37.385 164.625 38.135 165.145 ;
        RECT 35.085 164.275 35.855 164.495 ;
        RECT 35.065 163.365 35.405 164.095 ;
        RECT 35.585 163.545 35.855 164.275 ;
        RECT 36.035 164.255 37.195 164.495 ;
        RECT 38.305 164.455 39.055 164.975 ;
        RECT 41.270 164.540 41.610 165.370 ;
        RECT 36.035 163.545 36.265 164.255 ;
        RECT 36.435 163.365 36.765 164.075 ;
        RECT 36.935 163.545 37.195 164.255 ;
        RECT 37.385 163.365 39.055 164.455 ;
        RECT 39.225 163.365 39.515 164.530 ;
        RECT 43.090 163.800 43.440 165.050 ;
        RECT 46.790 164.540 47.130 165.370 ;
        RECT 48.610 163.800 48.960 165.050 ;
        RECT 52.310 164.540 52.650 165.370 ;
        RECT 56.245 165.145 57.915 165.915 ;
        RECT 58.255 165.455 58.510 165.915 ;
        RECT 58.680 165.285 59.010 165.745 ;
        RECT 59.180 165.455 59.350 165.915 ;
        RECT 59.520 165.285 59.850 165.745 ;
        RECT 60.020 165.455 60.190 165.915 ;
        RECT 60.360 165.285 60.690 165.745 ;
        RECT 60.860 165.455 61.030 165.915 ;
        RECT 61.200 165.285 61.530 165.745 ;
        RECT 61.700 165.455 62.005 165.915 ;
        RECT 54.130 163.800 54.480 165.050 ;
        RECT 56.245 164.625 56.995 165.145 ;
        RECT 58.085 165.095 62.055 165.285 ;
        RECT 62.690 165.265 62.960 165.475 ;
        RECT 63.180 165.455 63.510 165.915 ;
        RECT 64.020 165.455 64.770 165.745 ;
        RECT 62.690 165.095 64.025 165.265 ;
        RECT 57.165 164.455 57.915 164.975 ;
        RECT 39.685 163.365 45.030 163.800 ;
        RECT 45.205 163.365 50.550 163.800 ;
        RECT 50.725 163.365 56.070 163.800 ;
        RECT 56.245 163.365 57.915 164.455 ;
        RECT 58.085 164.505 58.430 165.095 ;
        RECT 58.680 164.895 61.535 164.925 ;
        RECT 58.605 164.725 61.535 164.895 ;
        RECT 58.680 164.675 61.535 164.725 ;
        RECT 61.735 164.505 62.055 165.095 ;
        RECT 63.855 164.925 64.025 165.095 ;
        RECT 62.690 164.685 63.040 164.925 ;
        RECT 63.210 164.685 63.685 164.925 ;
        RECT 63.855 164.675 64.230 164.925 ;
        RECT 63.855 164.505 64.025 164.675 ;
        RECT 58.085 164.335 62.055 164.505 ;
        RECT 62.690 164.335 64.025 164.505 ;
        RECT 58.255 163.365 58.510 164.165 ;
        RECT 58.680 163.535 59.010 164.335 ;
        RECT 59.180 163.365 59.350 164.165 ;
        RECT 59.520 163.535 59.850 164.335 ;
        RECT 60.020 163.365 60.190 164.165 ;
        RECT 60.360 163.535 60.690 164.335 ;
        RECT 60.860 163.365 61.030 164.165 ;
        RECT 61.200 163.535 61.530 164.335 ;
        RECT 62.690 164.175 62.970 164.335 ;
        RECT 64.400 164.165 64.770 165.455 ;
        RECT 64.985 165.190 65.275 165.915 ;
        RECT 65.445 165.415 65.745 165.745 ;
        RECT 65.915 165.435 66.190 165.915 ;
        RECT 61.700 163.365 62.000 164.165 ;
        RECT 63.180 163.365 63.430 164.165 ;
        RECT 63.600 163.995 64.770 164.165 ;
        RECT 63.600 163.535 63.930 163.995 ;
        RECT 64.100 163.365 64.315 163.825 ;
        RECT 64.985 163.365 65.275 164.530 ;
        RECT 65.445 164.505 65.615 165.415 ;
        RECT 66.370 165.265 66.665 165.655 ;
        RECT 66.835 165.435 67.090 165.915 ;
        RECT 67.265 165.265 67.525 165.655 ;
        RECT 67.695 165.435 67.975 165.915 ;
        RECT 68.725 165.455 68.970 165.915 ;
        RECT 65.785 164.675 66.135 165.245 ;
        RECT 66.370 165.095 68.020 165.265 ;
        RECT 66.305 164.755 67.445 164.925 ;
        RECT 66.305 164.505 66.475 164.755 ;
        RECT 67.615 164.585 68.020 165.095 ;
        RECT 68.665 164.675 68.980 165.285 ;
        RECT 69.150 164.925 69.400 165.735 ;
        RECT 69.570 165.390 69.830 165.915 ;
        RECT 70.000 165.265 70.260 165.720 ;
        RECT 70.430 165.435 70.690 165.915 ;
        RECT 70.860 165.265 71.120 165.720 ;
        RECT 71.290 165.435 71.550 165.915 ;
        RECT 71.720 165.265 71.980 165.720 ;
        RECT 72.150 165.435 72.410 165.915 ;
        RECT 72.580 165.265 72.840 165.720 ;
        RECT 73.010 165.435 73.310 165.915 ;
        RECT 73.725 165.370 79.070 165.915 ;
        RECT 79.245 165.370 84.590 165.915 ;
        RECT 84.765 165.370 90.110 165.915 ;
        RECT 70.000 165.095 73.310 165.265 ;
        RECT 69.150 164.675 72.170 164.925 ;
        RECT 65.445 164.335 66.475 164.505 ;
        RECT 67.265 164.415 68.020 164.585 ;
        RECT 65.445 163.535 65.755 164.335 ;
        RECT 67.265 164.165 67.525 164.415 ;
        RECT 65.925 163.365 66.235 164.165 ;
        RECT 66.405 163.995 67.525 164.165 ;
        RECT 66.405 163.535 66.665 163.995 ;
        RECT 66.835 163.365 67.090 163.825 ;
        RECT 67.265 163.535 67.525 163.995 ;
        RECT 67.695 163.365 67.980 164.235 ;
        RECT 68.675 163.365 68.970 164.475 ;
        RECT 69.150 163.540 69.400 164.675 ;
        RECT 72.340 164.505 73.310 165.095 ;
        RECT 75.310 164.540 75.650 165.370 ;
        RECT 69.570 163.365 69.830 164.475 ;
        RECT 70.000 164.265 73.310 164.505 ;
        RECT 70.000 163.540 70.260 164.265 ;
        RECT 70.430 163.365 70.690 164.095 ;
        RECT 70.860 163.540 71.120 164.265 ;
        RECT 71.290 163.365 71.550 164.095 ;
        RECT 71.720 163.540 71.980 164.265 ;
        RECT 72.150 163.365 72.410 164.095 ;
        RECT 72.580 163.540 72.840 164.265 ;
        RECT 73.010 163.365 73.305 164.095 ;
        RECT 77.130 163.800 77.480 165.050 ;
        RECT 80.830 164.540 81.170 165.370 ;
        RECT 82.650 163.800 83.000 165.050 ;
        RECT 86.350 164.540 86.690 165.370 ;
        RECT 90.745 165.165 91.955 165.915 ;
        RECT 100.130 165.480 102.050 166.750 ;
        RECT 103.560 166.740 104.120 166.750 ;
        RECT 103.790 165.650 104.120 166.740 ;
        RECT 104.490 166.270 105.530 166.440 ;
        RECT 104.490 165.830 105.530 166.000 ;
        RECT 105.700 165.970 105.870 166.300 ;
        RECT 103.950 165.430 104.120 165.650 ;
        RECT 106.210 165.430 106.380 166.840 ;
        RECT 103.950 165.260 106.380 165.430 ;
        RECT 107.960 167.350 118.590 167.520 ;
        RECT 120.020 176.580 126.250 176.740 ;
        RECT 120.020 174.320 120.690 176.580 ;
        RECT 121.360 176.010 125.400 176.180 ;
        RECT 121.020 174.950 121.190 175.950 ;
        RECT 125.570 174.950 125.740 175.950 ;
        RECT 121.360 174.720 125.400 174.890 ;
        RECT 126.080 174.320 126.250 176.580 ;
        RECT 120.020 174.150 126.250 174.320 ;
        RECT 120.020 170.890 120.690 174.150 ;
        RECT 121.360 173.580 125.400 173.750 ;
        RECT 121.020 171.520 121.190 173.520 ;
        RECT 125.570 171.520 125.740 173.520 ;
        RECT 121.360 171.290 125.400 171.460 ;
        RECT 126.080 170.890 126.250 174.150 ;
        RECT 120.020 170.720 126.250 170.890 ;
        RECT 120.020 167.460 120.690 170.720 ;
        RECT 121.360 170.150 125.400 170.320 ;
        RECT 121.020 168.090 121.190 170.090 ;
        RECT 125.570 168.090 125.740 170.090 ;
        RECT 121.360 167.860 125.400 168.030 ;
        RECT 126.080 167.460 126.250 170.720 ;
        RECT 120.020 167.450 126.250 167.460 ;
        RECT 127.840 176.720 137.670 176.760 ;
        RECT 127.840 176.590 138.470 176.720 ;
        RECT 127.840 174.330 128.010 176.590 ;
        RECT 128.735 176.020 136.775 176.190 ;
        RECT 128.350 174.960 128.520 175.960 ;
        RECT 136.990 174.960 137.160 175.960 ;
        RECT 128.735 174.730 136.775 174.900 ;
        RECT 137.500 174.330 138.470 176.590 ;
        RECT 127.840 174.160 138.470 174.330 ;
        RECT 127.840 170.900 128.010 174.160 ;
        RECT 128.735 173.590 136.775 173.760 ;
        RECT 128.350 171.530 128.520 173.530 ;
        RECT 136.990 171.530 137.160 173.530 ;
        RECT 128.735 171.300 136.775 171.470 ;
        RECT 137.500 170.900 138.470 174.160 ;
        RECT 127.840 170.730 138.470 170.900 ;
        RECT 127.840 167.470 128.010 170.730 ;
        RECT 128.735 170.160 136.775 170.330 ;
        RECT 128.350 168.100 128.520 170.100 ;
        RECT 136.990 168.100 137.160 170.100 ;
        RECT 128.735 167.870 136.775 168.040 ;
        RECT 137.500 167.470 138.470 170.730 ;
        RECT 120.020 167.350 126.260 167.450 ;
        RECT 88.170 163.800 88.520 165.050 ;
        RECT 90.745 164.455 91.265 164.995 ;
        RECT 91.435 164.625 91.955 165.165 ;
        RECT 107.960 165.090 108.130 167.350 ;
        RECT 108.855 166.780 116.895 166.950 ;
        RECT 108.470 165.720 108.640 166.720 ;
        RECT 117.110 165.720 117.280 166.720 ;
        RECT 108.855 165.490 116.895 165.660 ;
        RECT 117.620 165.090 118.590 167.350 ;
        RECT 120.010 166.790 126.260 167.350 ;
        RECT 120.010 166.770 125.180 166.790 ;
        RECT 120.010 166.700 124.000 166.770 ;
        RECT 120.010 165.430 121.930 166.700 ;
        RECT 123.440 166.690 124.000 166.700 ;
        RECT 123.670 165.600 124.000 166.690 ;
        RECT 124.370 166.220 125.410 166.390 ;
        RECT 124.370 165.780 125.410 165.950 ;
        RECT 125.580 165.920 125.750 166.250 ;
        RECT 123.830 165.380 124.000 165.600 ;
        RECT 126.090 165.380 126.260 166.790 ;
        RECT 123.830 165.210 126.260 165.380 ;
        RECT 127.840 167.300 138.470 167.470 ;
        RECT 140.050 176.630 146.280 176.790 ;
        RECT 140.050 174.370 140.720 176.630 ;
        RECT 141.390 176.060 145.430 176.230 ;
        RECT 141.050 175.000 141.220 176.000 ;
        RECT 145.600 175.000 145.770 176.000 ;
        RECT 141.390 174.770 145.430 174.940 ;
        RECT 146.110 174.370 146.280 176.630 ;
        RECT 140.050 174.200 146.280 174.370 ;
        RECT 140.050 170.940 140.720 174.200 ;
        RECT 141.390 173.630 145.430 173.800 ;
        RECT 141.050 171.570 141.220 173.570 ;
        RECT 145.600 171.570 145.770 173.570 ;
        RECT 141.390 171.340 145.430 171.510 ;
        RECT 146.110 170.940 146.280 174.200 ;
        RECT 140.050 170.770 146.280 170.940 ;
        RECT 140.050 167.510 140.720 170.770 ;
        RECT 141.390 170.200 145.430 170.370 ;
        RECT 141.050 168.140 141.220 170.140 ;
        RECT 145.600 168.140 145.770 170.140 ;
        RECT 141.390 167.910 145.430 168.080 ;
        RECT 146.110 167.510 146.280 170.770 ;
        RECT 140.050 167.500 146.280 167.510 ;
        RECT 147.870 176.770 157.700 176.810 ;
        RECT 147.870 176.640 158.500 176.770 ;
        RECT 147.870 174.380 148.040 176.640 ;
        RECT 148.765 176.070 156.805 176.240 ;
        RECT 148.380 175.010 148.550 176.010 ;
        RECT 157.020 175.010 157.190 176.010 ;
        RECT 148.765 174.780 156.805 174.950 ;
        RECT 157.530 174.380 158.500 176.640 ;
        RECT 147.870 174.210 158.500 174.380 ;
        RECT 147.870 170.950 148.040 174.210 ;
        RECT 148.765 173.640 156.805 173.810 ;
        RECT 148.380 171.580 148.550 173.580 ;
        RECT 157.020 171.580 157.190 173.580 ;
        RECT 148.765 171.350 156.805 171.520 ;
        RECT 157.530 170.950 158.500 174.210 ;
        RECT 147.870 170.780 158.500 170.950 ;
        RECT 147.870 167.520 148.040 170.780 ;
        RECT 148.765 170.210 156.805 170.380 ;
        RECT 148.380 168.150 148.550 170.150 ;
        RECT 157.020 168.150 157.190 170.150 ;
        RECT 148.765 167.920 156.805 168.090 ;
        RECT 157.530 167.520 158.500 170.780 ;
        RECT 140.050 167.400 146.290 167.500 ;
        RECT 107.960 165.060 118.590 165.090 ;
        RECT 107.930 164.950 118.590 165.060 ;
        RECT 127.840 165.040 128.010 167.300 ;
        RECT 128.735 166.730 136.775 166.900 ;
        RECT 128.350 165.670 128.520 166.670 ;
        RECT 136.990 165.670 137.160 166.670 ;
        RECT 128.735 165.440 136.775 165.610 ;
        RECT 137.500 165.040 138.470 167.300 ;
        RECT 140.040 166.840 146.290 167.400 ;
        RECT 140.040 166.820 145.210 166.840 ;
        RECT 140.040 166.750 144.030 166.820 ;
        RECT 140.040 165.480 141.960 166.750 ;
        RECT 143.470 166.740 144.030 166.750 ;
        RECT 143.700 165.650 144.030 166.740 ;
        RECT 144.400 166.270 145.440 166.440 ;
        RECT 144.400 165.830 145.440 166.000 ;
        RECT 145.610 165.970 145.780 166.300 ;
        RECT 143.860 165.430 144.030 165.650 ;
        RECT 146.120 165.430 146.290 166.840 ;
        RECT 143.860 165.260 146.290 165.430 ;
        RECT 147.870 167.350 158.500 167.520 ;
        RECT 147.870 165.090 148.040 167.350 ;
        RECT 148.765 166.780 156.805 166.950 ;
        RECT 148.380 165.720 148.550 166.720 ;
        RECT 157.020 165.720 157.190 166.720 ;
        RECT 148.765 165.490 156.805 165.660 ;
        RECT 157.530 165.090 158.500 167.350 ;
        RECT 147.870 165.060 158.500 165.090 ;
        RECT 127.840 165.010 138.470 165.040 ;
        RECT 106.180 164.900 118.590 164.950 ;
        RECT 127.810 164.900 138.470 165.010 ;
        RECT 147.840 164.950 158.500 165.060 ;
        RECT 146.090 164.900 158.500 164.950 ;
        RECT 101.840 164.730 118.590 164.900 ;
        RECT 126.060 164.850 138.470 164.900 ;
        RECT 73.725 163.365 79.070 163.800 ;
        RECT 79.245 163.365 84.590 163.800 ;
        RECT 84.765 163.365 90.110 163.800 ;
        RECT 90.745 163.365 91.955 164.455 ;
        RECT 13.380 163.195 92.040 163.365 ;
        RECT 101.840 163.320 102.010 164.730 ;
        RECT 102.380 164.160 105.420 164.330 ;
        RECT 102.380 163.720 105.420 163.890 ;
        RECT 105.635 163.860 105.805 164.190 ;
        RECT 106.140 163.970 118.590 164.730 ;
        RECT 121.720 164.680 138.470 164.850 ;
        RECT 106.140 163.960 118.480 163.970 ;
        RECT 106.140 163.950 112.020 163.960 ;
        RECT 106.140 163.930 106.710 163.950 ;
        RECT 107.930 163.940 112.020 163.950 ;
        RECT 106.150 163.320 106.320 163.930 ;
        RECT 13.465 162.105 14.675 163.195 ;
        RECT 14.845 162.760 20.190 163.195 ;
        RECT 20.365 162.760 25.710 163.195 ;
        RECT 13.465 161.395 13.985 161.935 ;
        RECT 14.155 161.565 14.675 162.105 ;
        RECT 13.465 160.645 14.675 161.395 ;
        RECT 16.430 161.190 16.770 162.020 ;
        RECT 18.250 161.510 18.600 162.760 ;
        RECT 21.950 161.190 22.290 162.020 ;
        RECT 23.770 161.510 24.120 162.760 ;
        RECT 26.345 162.030 26.635 163.195 ;
        RECT 26.805 162.685 27.065 163.195 ;
        RECT 26.805 161.635 27.145 162.515 ;
        RECT 27.315 161.805 27.485 163.025 ;
        RECT 27.725 162.690 28.340 163.195 ;
        RECT 27.725 162.155 27.975 162.520 ;
        RECT 28.145 162.515 28.340 162.690 ;
        RECT 28.510 162.685 28.985 163.025 ;
        RECT 29.155 162.650 29.370 163.195 ;
        RECT 28.145 162.325 28.475 162.515 ;
        RECT 28.695 162.155 29.410 162.450 ;
        RECT 29.580 162.325 29.855 163.025 ;
        RECT 27.725 161.985 29.515 162.155 ;
        RECT 27.315 161.555 28.110 161.805 ;
        RECT 27.315 161.465 27.565 161.555 ;
        RECT 14.845 160.645 20.190 161.190 ;
        RECT 20.365 160.645 25.710 161.190 ;
        RECT 26.345 160.645 26.635 161.370 ;
        RECT 26.805 160.645 27.065 161.465 ;
        RECT 27.235 161.045 27.565 161.465 ;
        RECT 28.280 161.130 28.535 161.985 ;
        RECT 27.745 160.865 28.535 161.130 ;
        RECT 28.705 161.285 29.115 161.805 ;
        RECT 29.285 161.555 29.515 161.985 ;
        RECT 29.685 161.295 29.855 162.325 ;
        RECT 30.210 162.225 30.600 162.400 ;
        RECT 31.085 162.395 31.415 163.195 ;
        RECT 31.585 162.405 32.120 163.025 ;
        RECT 30.210 162.055 31.635 162.225 ;
        RECT 30.085 161.325 30.440 161.885 ;
        RECT 28.705 160.865 28.905 161.285 ;
        RECT 29.095 160.645 29.425 161.105 ;
        RECT 29.595 160.815 29.855 161.295 ;
        RECT 30.610 161.155 30.780 162.055 ;
        RECT 30.950 161.325 31.215 161.885 ;
        RECT 31.465 161.555 31.635 162.055 ;
        RECT 31.805 161.385 32.120 162.405 ;
        RECT 32.940 162.185 33.240 163.025 ;
        RECT 33.435 162.355 33.685 163.195 ;
        RECT 34.275 162.605 35.080 163.025 ;
        RECT 33.855 162.435 35.420 162.605 ;
        RECT 33.855 162.185 34.025 162.435 ;
        RECT 32.940 162.015 34.025 162.185 ;
        RECT 32.785 161.555 33.115 161.845 ;
        RECT 33.285 161.385 33.455 162.015 ;
        RECT 34.195 161.885 34.515 162.265 ;
        RECT 34.705 162.175 35.080 162.265 ;
        RECT 34.685 162.005 35.080 162.175 ;
        RECT 35.250 162.185 35.420 162.435 ;
        RECT 35.590 162.355 35.920 163.195 ;
        RECT 36.090 162.435 36.755 163.025 ;
        RECT 35.250 162.015 36.170 162.185 ;
        RECT 33.625 161.635 33.955 161.845 ;
        RECT 34.135 161.635 34.515 161.885 ;
        RECT 34.705 161.845 35.080 162.005 ;
        RECT 36.000 161.845 36.170 162.015 ;
        RECT 34.705 161.635 35.190 161.845 ;
        RECT 35.380 161.635 35.830 161.845 ;
        RECT 36.000 161.635 36.335 161.845 ;
        RECT 36.505 161.465 36.755 162.435 ;
        RECT 30.190 160.645 30.430 161.155 ;
        RECT 30.610 160.825 30.890 161.155 ;
        RECT 31.120 160.645 31.335 161.155 ;
        RECT 31.505 160.815 32.120 161.385 ;
        RECT 32.945 161.205 33.455 161.385 ;
        RECT 33.860 161.295 35.560 161.465 ;
        RECT 33.860 161.205 34.245 161.295 ;
        RECT 32.945 160.815 33.275 161.205 ;
        RECT 33.445 160.865 34.630 161.035 ;
        RECT 34.890 160.645 35.060 161.115 ;
        RECT 35.230 160.830 35.560 161.295 ;
        RECT 35.730 160.645 35.900 161.465 ;
        RECT 36.070 160.825 36.755 161.465 ;
        RECT 36.925 161.590 37.205 163.025 ;
        RECT 37.375 162.420 38.085 163.195 ;
        RECT 38.255 162.250 38.585 163.025 ;
        RECT 37.435 162.035 38.585 162.250 ;
        RECT 36.925 160.815 37.265 161.590 ;
        RECT 37.435 161.465 37.720 162.035 ;
        RECT 37.905 161.635 38.375 161.865 ;
        RECT 38.780 161.835 38.995 162.950 ;
        RECT 39.175 162.475 39.505 163.195 ;
        RECT 40.625 162.685 40.925 163.195 ;
        RECT 41.095 162.685 41.475 162.855 ;
        RECT 42.055 162.685 42.685 163.195 ;
        RECT 41.095 162.515 41.265 162.685 ;
        RECT 42.855 162.515 43.185 163.025 ;
        RECT 43.355 162.685 43.655 163.195 ;
        RECT 40.605 162.315 41.265 162.515 ;
        RECT 41.435 162.345 43.655 162.515 ;
        RECT 39.285 161.835 39.515 162.175 ;
        RECT 38.545 161.655 38.995 161.835 ;
        RECT 38.545 161.635 38.875 161.655 ;
        RECT 39.185 161.635 39.515 161.835 ;
        RECT 37.435 161.275 38.145 161.465 ;
        RECT 37.845 161.135 38.145 161.275 ;
        RECT 38.335 161.275 39.515 161.465 ;
        RECT 38.335 161.195 38.665 161.275 ;
        RECT 37.845 161.125 38.160 161.135 ;
        RECT 37.845 161.115 38.170 161.125 ;
        RECT 37.845 161.110 38.180 161.115 ;
        RECT 37.435 160.645 37.605 161.105 ;
        RECT 37.845 161.100 38.185 161.110 ;
        RECT 37.845 161.095 38.190 161.100 ;
        RECT 37.845 161.085 38.195 161.095 ;
        RECT 37.845 161.080 38.200 161.085 ;
        RECT 37.845 160.815 38.205 161.080 ;
        RECT 38.835 160.645 39.005 161.105 ;
        RECT 39.175 160.815 39.515 161.275 ;
        RECT 40.605 161.385 40.775 162.315 ;
        RECT 41.435 162.145 41.605 162.345 ;
        RECT 40.945 161.975 41.605 162.145 ;
        RECT 41.775 162.005 43.315 162.175 ;
        RECT 40.945 161.555 41.115 161.975 ;
        RECT 41.775 161.805 41.945 162.005 ;
        RECT 41.345 161.635 41.945 161.805 ;
        RECT 42.115 161.635 42.810 161.835 ;
        RECT 43.070 161.555 43.315 162.005 ;
        RECT 41.435 161.385 42.345 161.465 ;
        RECT 40.605 160.905 40.925 161.385 ;
        RECT 41.095 161.295 42.345 161.385 ;
        RECT 41.095 161.215 41.605 161.295 ;
        RECT 41.095 160.815 41.325 161.215 ;
        RECT 41.495 160.645 41.845 161.035 ;
        RECT 42.015 160.815 42.345 161.295 ;
        RECT 42.515 160.645 42.685 161.465 ;
        RECT 43.485 161.385 43.655 162.345 ;
        RECT 43.825 162.105 46.415 163.195 ;
        RECT 47.050 162.770 47.385 163.195 ;
        RECT 47.555 162.590 47.740 162.995 ;
        RECT 43.190 160.840 43.655 161.385 ;
        RECT 43.825 161.415 45.035 161.935 ;
        RECT 45.205 161.585 46.415 162.105 ;
        RECT 47.075 162.415 47.740 162.590 ;
        RECT 47.945 162.415 48.275 163.195 ;
        RECT 43.825 160.645 46.415 161.415 ;
        RECT 47.075 161.385 47.415 162.415 ;
        RECT 48.445 162.225 48.715 162.995 ;
        RECT 47.585 162.055 48.715 162.225 ;
        RECT 47.585 161.555 47.835 162.055 ;
        RECT 47.075 161.215 47.760 161.385 ;
        RECT 48.015 161.305 48.375 161.885 ;
        RECT 47.050 160.645 47.385 161.045 ;
        RECT 47.555 160.815 47.760 161.215 ;
        RECT 48.545 161.145 48.715 162.055 ;
        RECT 47.970 160.645 48.245 161.125 ;
        RECT 48.455 160.815 48.715 161.145 ;
        RECT 48.895 162.135 49.225 162.985 ;
        RECT 48.895 161.370 49.085 162.135 ;
        RECT 49.395 162.055 49.645 163.195 ;
        RECT 49.835 162.555 50.085 162.975 ;
        RECT 50.315 162.725 50.645 163.195 ;
        RECT 50.875 162.555 51.125 162.975 ;
        RECT 49.835 162.385 51.125 162.555 ;
        RECT 51.305 162.555 51.635 162.985 ;
        RECT 51.305 162.385 51.760 162.555 ;
        RECT 49.825 161.885 50.040 162.215 ;
        RECT 49.255 161.555 49.565 161.885 ;
        RECT 49.735 161.555 50.040 161.885 ;
        RECT 50.215 161.555 50.500 162.215 ;
        RECT 50.695 161.555 50.960 162.215 ;
        RECT 51.175 161.555 51.420 162.215 ;
        RECT 49.395 161.385 49.565 161.555 ;
        RECT 51.590 161.385 51.760 162.385 ;
        RECT 52.105 162.030 52.395 163.195 ;
        RECT 52.565 162.105 53.775 163.195 ;
        RECT 48.895 160.860 49.225 161.370 ;
        RECT 49.395 161.215 51.760 161.385 ;
        RECT 52.565 161.395 53.085 161.935 ;
        RECT 53.255 161.565 53.775 162.105 ;
        RECT 53.980 162.405 54.515 163.025 ;
        RECT 49.395 160.645 49.725 161.045 ;
        RECT 50.775 160.875 51.105 161.215 ;
        RECT 51.275 160.645 51.605 161.045 ;
        RECT 52.105 160.645 52.395 161.370 ;
        RECT 52.565 160.645 53.775 161.395 ;
        RECT 53.980 161.385 54.295 162.405 ;
        RECT 54.685 162.395 55.015 163.195 ;
        RECT 55.500 162.225 55.890 162.400 ;
        RECT 54.465 162.055 55.890 162.225 ;
        RECT 56.335 162.265 56.505 163.025 ;
        RECT 56.720 162.435 57.050 163.195 ;
        RECT 56.335 162.095 57.050 162.265 ;
        RECT 57.220 162.120 57.475 163.025 ;
        RECT 54.465 161.555 54.635 162.055 ;
        RECT 53.980 160.815 54.595 161.385 ;
        RECT 54.885 161.325 55.150 161.885 ;
        RECT 55.320 161.155 55.490 162.055 ;
        RECT 55.660 161.325 56.015 161.885 ;
        RECT 56.245 161.545 56.600 161.915 ;
        RECT 56.880 161.885 57.050 162.095 ;
        RECT 56.880 161.555 57.135 161.885 ;
        RECT 56.880 161.365 57.050 161.555 ;
        RECT 57.305 161.390 57.475 162.120 ;
        RECT 57.650 162.045 57.910 163.195 ;
        RECT 59.015 162.055 59.345 163.195 ;
        RECT 59.875 162.225 60.205 163.010 ;
        RECT 59.525 162.055 60.205 162.225 ;
        RECT 60.390 162.805 60.725 163.025 ;
        RECT 61.730 162.815 62.085 163.195 ;
        RECT 60.390 162.185 60.645 162.805 ;
        RECT 60.895 162.645 61.125 162.685 ;
        RECT 62.255 162.645 62.505 163.025 ;
        RECT 60.895 162.445 62.505 162.645 ;
        RECT 60.895 162.355 61.080 162.445 ;
        RECT 61.670 162.435 62.505 162.445 ;
        RECT 62.755 162.415 63.005 163.195 ;
        RECT 63.175 162.345 63.435 163.025 ;
        RECT 64.105 162.735 64.320 163.195 ;
        RECT 64.490 162.565 64.820 163.025 ;
        RECT 61.235 162.245 61.565 162.275 ;
        RECT 61.235 162.185 63.035 162.245 ;
        RECT 60.390 162.075 63.095 162.185 ;
        RECT 59.005 161.635 59.355 161.885 ;
        RECT 56.335 161.195 57.050 161.365 ;
        RECT 54.765 160.645 54.980 161.155 ;
        RECT 55.210 160.825 55.490 161.155 ;
        RECT 55.670 160.645 55.910 161.155 ;
        RECT 56.335 160.815 56.505 161.195 ;
        RECT 56.720 160.645 57.050 161.025 ;
        RECT 57.220 160.815 57.475 161.390 ;
        RECT 57.650 160.645 57.910 161.485 ;
        RECT 59.525 161.455 59.695 162.055 ;
        RECT 60.390 162.015 61.565 162.075 ;
        RECT 62.895 162.040 63.095 162.075 ;
        RECT 59.865 161.635 60.215 161.885 ;
        RECT 60.385 161.635 60.875 161.835 ;
        RECT 61.065 161.635 61.540 161.845 ;
        RECT 59.015 160.645 59.285 161.455 ;
        RECT 59.455 160.815 59.785 161.455 ;
        RECT 59.955 160.645 60.195 161.455 ;
        RECT 60.390 160.645 60.845 161.410 ;
        RECT 61.320 161.235 61.540 161.635 ;
        RECT 61.785 161.635 62.115 161.845 ;
        RECT 61.785 161.235 61.995 161.635 ;
        RECT 62.285 161.600 62.695 161.905 ;
        RECT 62.925 161.465 63.095 162.040 ;
        RECT 62.825 161.345 63.095 161.465 ;
        RECT 62.250 161.300 63.095 161.345 ;
        RECT 62.250 161.175 63.005 161.300 ;
        RECT 62.250 161.025 62.420 161.175 ;
        RECT 63.265 161.155 63.435 162.345 ;
        RECT 63.205 161.145 63.435 161.155 ;
        RECT 61.120 160.815 62.420 161.025 ;
        RECT 62.675 160.645 63.005 161.005 ;
        RECT 63.175 160.815 63.435 161.145 ;
        RECT 63.650 162.395 64.820 162.565 ;
        RECT 64.990 162.395 65.240 163.195 ;
        RECT 63.650 161.105 64.020 162.395 ;
        RECT 65.450 162.225 65.730 162.385 ;
        RECT 64.395 162.055 65.730 162.225 ;
        RECT 65.905 162.105 67.575 163.195 ;
        RECT 64.395 161.885 64.565 162.055 ;
        RECT 64.190 161.635 64.565 161.885 ;
        RECT 64.735 161.635 65.210 161.875 ;
        RECT 65.380 161.635 65.730 161.875 ;
        RECT 64.395 161.465 64.565 161.635 ;
        RECT 64.395 161.295 65.730 161.465 ;
        RECT 63.650 160.815 64.400 161.105 ;
        RECT 64.910 160.645 65.240 161.105 ;
        RECT 65.460 161.085 65.730 161.295 ;
        RECT 65.905 161.415 66.655 161.935 ;
        RECT 66.825 161.585 67.575 162.105 ;
        RECT 67.745 162.345 68.125 163.025 ;
        RECT 68.715 162.345 68.885 163.195 ;
        RECT 69.055 162.515 69.385 163.025 ;
        RECT 69.555 162.685 69.725 163.195 ;
        RECT 69.895 162.515 70.295 163.025 ;
        RECT 69.055 162.345 70.295 162.515 ;
        RECT 65.905 160.645 67.575 161.415 ;
        RECT 67.745 161.385 67.915 162.345 ;
        RECT 68.085 162.005 69.390 162.175 ;
        RECT 70.475 162.095 70.795 163.025 ;
        RECT 71.050 162.575 71.225 163.025 ;
        RECT 71.395 162.755 71.725 163.195 ;
        RECT 72.030 162.605 72.200 163.025 ;
        RECT 72.435 162.785 73.105 163.195 ;
        RECT 73.320 162.605 73.490 163.025 ;
        RECT 73.690 162.785 74.020 163.195 ;
        RECT 71.050 162.405 71.680 162.575 ;
        RECT 68.085 161.555 68.330 162.005 ;
        RECT 68.500 161.635 69.050 161.835 ;
        RECT 69.220 161.805 69.390 162.005 ;
        RECT 70.165 161.925 70.795 162.095 ;
        RECT 69.220 161.635 69.595 161.805 ;
        RECT 69.765 161.385 69.995 161.885 ;
        RECT 67.745 161.215 69.995 161.385 ;
        RECT 67.795 160.645 68.125 161.035 ;
        RECT 68.295 160.895 68.465 161.215 ;
        RECT 70.165 161.045 70.335 161.925 ;
        RECT 70.965 161.555 71.330 162.235 ;
        RECT 71.510 161.885 71.680 162.405 ;
        RECT 72.030 162.435 74.045 162.605 ;
        RECT 71.510 161.555 71.860 161.885 ;
        RECT 68.635 160.645 68.965 161.035 ;
        RECT 69.380 160.875 70.335 161.045 ;
        RECT 70.505 160.645 70.795 161.480 ;
        RECT 71.510 161.385 71.680 161.555 ;
        RECT 71.050 161.215 71.680 161.385 ;
        RECT 71.050 160.815 71.225 161.215 ;
        RECT 72.030 161.145 72.200 162.435 ;
        RECT 71.395 160.645 71.725 161.025 ;
        RECT 71.970 160.815 72.200 161.145 ;
        RECT 72.400 160.980 72.680 162.255 ;
        RECT 72.905 161.835 73.175 162.255 ;
        RECT 72.865 161.665 73.175 161.835 ;
        RECT 72.905 160.980 73.175 161.665 ;
        RECT 73.365 161.225 73.705 162.255 ;
        RECT 73.875 161.885 74.045 162.435 ;
        RECT 74.215 162.055 74.475 163.025 ;
        RECT 74.645 162.105 77.235 163.195 ;
        RECT 73.875 161.555 74.135 161.885 ;
        RECT 74.305 161.365 74.475 162.055 ;
        RECT 73.635 160.645 73.965 161.025 ;
        RECT 74.135 160.900 74.475 161.365 ;
        RECT 74.645 161.415 75.855 161.935 ;
        RECT 76.025 161.585 77.235 162.105 ;
        RECT 77.865 162.030 78.155 163.195 ;
        RECT 78.325 162.760 83.670 163.195 ;
        RECT 83.845 162.760 89.190 163.195 ;
        RECT 74.135 160.855 74.470 160.900 ;
        RECT 74.645 160.645 77.235 161.415 ;
        RECT 77.865 160.645 78.155 161.370 ;
        RECT 79.910 161.190 80.250 162.020 ;
        RECT 81.730 161.510 82.080 162.760 ;
        RECT 85.430 161.190 85.770 162.020 ;
        RECT 87.250 161.510 87.600 162.760 ;
        RECT 89.365 162.105 90.575 163.195 ;
        RECT 89.365 161.395 89.885 161.935 ;
        RECT 90.055 161.565 90.575 162.105 ;
        RECT 90.745 162.105 91.955 163.195 ;
        RECT 101.840 163.150 106.320 163.320 ;
        RECT 121.720 163.270 121.890 164.680 ;
        RECT 122.260 164.110 125.300 164.280 ;
        RECT 122.260 163.670 125.300 163.840 ;
        RECT 125.515 163.810 125.685 164.140 ;
        RECT 126.020 163.920 138.470 164.680 ;
        RECT 141.750 164.730 158.500 164.900 ;
        RECT 126.020 163.910 138.360 163.920 ;
        RECT 126.020 163.900 131.900 163.910 ;
        RECT 126.020 163.880 126.590 163.900 ;
        RECT 127.810 163.890 131.900 163.900 ;
        RECT 126.030 163.270 126.200 163.880 ;
        RECT 121.720 163.100 126.200 163.270 ;
        RECT 141.750 163.320 141.920 164.730 ;
        RECT 142.290 164.160 145.330 164.330 ;
        RECT 142.290 163.720 145.330 163.890 ;
        RECT 145.545 163.860 145.715 164.190 ;
        RECT 146.050 163.970 158.500 164.730 ;
        RECT 146.050 163.960 158.390 163.970 ;
        RECT 146.050 163.950 151.930 163.960 ;
        RECT 146.050 163.930 146.620 163.950 ;
        RECT 147.840 163.940 151.930 163.950 ;
        RECT 146.060 163.320 146.230 163.930 ;
        RECT 141.750 163.150 146.230 163.320 ;
        RECT 90.745 161.565 91.265 162.105 ;
        RECT 91.435 161.395 91.955 161.935 ;
        RECT 100.630 161.790 106.370 161.800 ;
        RECT 78.325 160.645 83.670 161.190 ;
        RECT 83.845 160.645 89.190 161.190 ;
        RECT 89.365 160.645 90.575 161.395 ;
        RECT 90.745 160.645 91.955 161.395 ;
        RECT 100.140 161.630 106.370 161.790 ;
        RECT 13.380 160.475 92.040 160.645 ;
        RECT 13.465 159.725 14.675 160.475 ;
        RECT 14.845 159.930 20.190 160.475 ;
        RECT 13.465 159.185 13.985 159.725 ;
        RECT 14.155 159.015 14.675 159.555 ;
        RECT 16.430 159.100 16.770 159.930 ;
        RECT 20.365 159.705 23.875 160.475 ;
        RECT 24.555 159.820 24.885 160.255 ;
        RECT 25.055 159.865 25.225 160.475 ;
        RECT 24.505 159.735 24.885 159.820 ;
        RECT 25.395 159.735 25.725 160.260 ;
        RECT 25.985 159.945 26.195 160.475 ;
        RECT 26.470 160.025 27.255 160.195 ;
        RECT 27.425 160.025 27.830 160.195 ;
        RECT 13.465 157.925 14.675 159.015 ;
        RECT 18.250 158.360 18.600 159.610 ;
        RECT 20.365 159.185 22.015 159.705 ;
        RECT 24.505 159.695 24.730 159.735 ;
        RECT 22.185 159.015 23.875 159.535 ;
        RECT 14.845 157.925 20.190 158.360 ;
        RECT 20.365 157.925 23.875 159.015 ;
        RECT 24.505 159.115 24.675 159.695 ;
        RECT 25.395 159.565 25.595 159.735 ;
        RECT 26.470 159.565 26.640 160.025 ;
        RECT 24.845 159.235 25.595 159.565 ;
        RECT 25.765 159.235 26.640 159.565 ;
        RECT 24.505 159.065 24.720 159.115 ;
        RECT 24.505 158.985 24.895 159.065 ;
        RECT 24.565 158.140 24.895 158.985 ;
        RECT 25.405 159.030 25.595 159.235 ;
        RECT 25.065 157.925 25.235 158.935 ;
        RECT 25.405 158.655 26.300 159.030 ;
        RECT 25.405 158.095 25.745 158.655 ;
        RECT 25.975 157.925 26.290 158.425 ;
        RECT 26.470 158.395 26.640 159.235 ;
        RECT 26.810 159.525 27.275 159.855 ;
        RECT 27.660 159.795 27.830 160.025 ;
        RECT 28.010 159.975 28.380 160.475 ;
        RECT 28.700 160.025 29.375 160.195 ;
        RECT 29.570 160.025 29.905 160.195 ;
        RECT 26.810 158.565 27.130 159.525 ;
        RECT 27.660 159.495 28.490 159.795 ;
        RECT 27.300 158.595 27.490 159.315 ;
        RECT 27.660 158.425 27.830 159.495 ;
        RECT 28.290 159.465 28.490 159.495 ;
        RECT 28.000 159.245 28.170 159.315 ;
        RECT 28.700 159.245 28.870 160.025 ;
        RECT 29.735 159.885 29.905 160.025 ;
        RECT 30.075 160.015 30.325 160.475 ;
        RECT 28.000 159.075 28.870 159.245 ;
        RECT 29.040 159.605 29.565 159.825 ;
        RECT 29.735 159.755 29.960 159.885 ;
        RECT 28.000 158.985 28.510 159.075 ;
        RECT 26.470 158.225 27.355 158.395 ;
        RECT 27.580 158.095 27.830 158.425 ;
        RECT 28.000 157.925 28.170 158.725 ;
        RECT 28.340 158.370 28.510 158.985 ;
        RECT 29.040 158.905 29.210 159.605 ;
        RECT 28.680 158.540 29.210 158.905 ;
        RECT 29.380 158.840 29.620 159.435 ;
        RECT 29.790 158.650 29.960 159.755 ;
        RECT 30.130 158.895 30.410 159.845 ;
        RECT 29.655 158.520 29.960 158.650 ;
        RECT 28.340 158.200 29.445 158.370 ;
        RECT 29.655 158.095 29.905 158.520 ;
        RECT 30.075 157.925 30.340 158.385 ;
        RECT 30.580 158.095 30.765 160.215 ;
        RECT 30.935 160.095 31.265 160.475 ;
        RECT 31.435 159.925 31.605 160.215 ;
        RECT 30.940 159.755 31.605 159.925 ;
        RECT 30.940 158.765 31.170 159.755 ;
        RECT 31.340 158.935 31.690 159.585 ;
        RECT 32.785 159.530 33.125 160.305 ;
        RECT 33.295 160.015 33.465 160.475 ;
        RECT 33.705 160.040 34.065 160.305 ;
        RECT 33.705 160.035 34.060 160.040 ;
        RECT 33.705 160.025 34.055 160.035 ;
        RECT 33.705 160.020 34.050 160.025 ;
        RECT 33.705 160.010 34.045 160.020 ;
        RECT 34.695 160.015 34.865 160.475 ;
        RECT 33.705 160.005 34.040 160.010 ;
        RECT 33.705 159.995 34.030 160.005 ;
        RECT 33.705 159.985 34.020 159.995 ;
        RECT 33.705 159.845 34.005 159.985 ;
        RECT 33.295 159.655 34.005 159.845 ;
        RECT 34.195 159.845 34.525 159.925 ;
        RECT 35.035 159.845 35.375 160.305 ;
        RECT 34.195 159.655 35.375 159.845 ;
        RECT 35.545 159.705 37.215 160.475 ;
        RECT 30.940 158.595 31.605 158.765 ;
        RECT 30.935 157.925 31.265 158.425 ;
        RECT 31.435 158.095 31.605 158.595 ;
        RECT 32.785 158.095 33.065 159.530 ;
        RECT 33.295 159.085 33.580 159.655 ;
        RECT 33.765 159.255 34.235 159.485 ;
        RECT 34.405 159.465 34.735 159.485 ;
        RECT 34.405 159.285 34.855 159.465 ;
        RECT 35.045 159.285 35.375 159.485 ;
        RECT 33.295 158.870 34.445 159.085 ;
        RECT 33.235 157.925 33.945 158.700 ;
        RECT 34.115 158.095 34.445 158.870 ;
        RECT 34.640 158.170 34.855 159.285 ;
        RECT 35.145 158.945 35.375 159.285 ;
        RECT 35.545 159.185 36.295 159.705 ;
        RECT 37.845 159.675 38.155 160.475 ;
        RECT 38.360 159.675 39.055 160.305 ;
        RECT 39.225 159.750 39.515 160.475 ;
        RECT 40.235 159.925 40.405 160.215 ;
        RECT 40.575 160.095 40.905 160.475 ;
        RECT 40.235 159.755 40.900 159.925 ;
        RECT 36.465 159.015 37.215 159.535 ;
        RECT 37.855 159.235 38.190 159.505 ;
        RECT 38.360 159.075 38.530 159.675 ;
        RECT 38.700 159.235 39.035 159.485 ;
        RECT 35.035 157.925 35.365 158.645 ;
        RECT 35.545 157.925 37.215 159.015 ;
        RECT 37.845 157.925 38.125 159.065 ;
        RECT 38.295 158.095 38.625 159.075 ;
        RECT 38.795 157.925 39.055 159.065 ;
        RECT 39.225 157.925 39.515 159.090 ;
        RECT 40.150 158.935 40.500 159.585 ;
        RECT 40.670 158.765 40.900 159.755 ;
        RECT 40.235 158.595 40.900 158.765 ;
        RECT 40.235 158.095 40.405 158.595 ;
        RECT 40.575 157.925 40.905 158.425 ;
        RECT 41.075 158.095 41.260 160.215 ;
        RECT 41.515 160.015 41.765 160.475 ;
        RECT 41.935 160.025 42.270 160.195 ;
        RECT 42.465 160.025 43.140 160.195 ;
        RECT 41.935 159.885 42.105 160.025 ;
        RECT 41.430 158.895 41.710 159.845 ;
        RECT 41.880 159.755 42.105 159.885 ;
        RECT 41.880 158.650 42.050 159.755 ;
        RECT 42.275 159.605 42.800 159.825 ;
        RECT 42.220 158.840 42.460 159.435 ;
        RECT 42.630 158.905 42.800 159.605 ;
        RECT 42.970 159.245 43.140 160.025 ;
        RECT 43.460 159.975 43.830 160.475 ;
        RECT 44.010 160.025 44.415 160.195 ;
        RECT 44.585 160.025 45.370 160.195 ;
        RECT 44.010 159.795 44.180 160.025 ;
        RECT 43.350 159.495 44.180 159.795 ;
        RECT 44.565 159.525 45.030 159.855 ;
        RECT 43.350 159.465 43.550 159.495 ;
        RECT 43.670 159.245 43.840 159.315 ;
        RECT 42.970 159.075 43.840 159.245 ;
        RECT 43.330 158.985 43.840 159.075 ;
        RECT 41.880 158.520 42.185 158.650 ;
        RECT 42.630 158.540 43.160 158.905 ;
        RECT 41.500 157.925 41.765 158.385 ;
        RECT 41.935 158.095 42.185 158.520 ;
        RECT 43.330 158.370 43.500 158.985 ;
        RECT 42.395 158.200 43.500 158.370 ;
        RECT 43.670 157.925 43.840 158.725 ;
        RECT 44.010 158.425 44.180 159.495 ;
        RECT 44.350 158.595 44.540 159.315 ;
        RECT 44.710 158.565 45.030 159.525 ;
        RECT 45.200 159.565 45.370 160.025 ;
        RECT 45.645 159.945 45.855 160.475 ;
        RECT 46.115 159.735 46.445 160.260 ;
        RECT 46.615 159.865 46.785 160.475 ;
        RECT 46.955 159.820 47.285 160.255 ;
        RECT 47.595 159.925 47.765 160.215 ;
        RECT 47.935 160.095 48.265 160.475 ;
        RECT 46.955 159.735 47.335 159.820 ;
        RECT 47.595 159.755 48.260 159.925 ;
        RECT 46.245 159.565 46.445 159.735 ;
        RECT 47.110 159.695 47.335 159.735 ;
        RECT 45.200 159.235 46.075 159.565 ;
        RECT 46.245 159.235 46.995 159.565 ;
        RECT 44.010 158.095 44.260 158.425 ;
        RECT 45.200 158.395 45.370 159.235 ;
        RECT 46.245 159.030 46.435 159.235 ;
        RECT 47.165 159.115 47.335 159.695 ;
        RECT 47.120 159.065 47.335 159.115 ;
        RECT 45.540 158.655 46.435 159.030 ;
        RECT 46.945 158.985 47.335 159.065 ;
        RECT 44.485 158.225 45.370 158.395 ;
        RECT 45.550 157.925 45.865 158.425 ;
        RECT 46.095 158.095 46.435 158.655 ;
        RECT 46.605 157.925 46.775 158.935 ;
        RECT 46.945 158.140 47.275 158.985 ;
        RECT 47.510 158.935 47.860 159.585 ;
        RECT 48.030 158.765 48.260 159.755 ;
        RECT 47.595 158.595 48.260 158.765 ;
        RECT 47.595 158.095 47.765 158.595 ;
        RECT 47.935 157.925 48.265 158.425 ;
        RECT 48.435 158.095 48.620 160.215 ;
        RECT 48.875 160.015 49.125 160.475 ;
        RECT 49.295 160.025 49.630 160.195 ;
        RECT 49.825 160.025 50.500 160.195 ;
        RECT 49.295 159.885 49.465 160.025 ;
        RECT 48.790 158.895 49.070 159.845 ;
        RECT 49.240 159.755 49.465 159.885 ;
        RECT 49.240 158.650 49.410 159.755 ;
        RECT 49.635 159.605 50.160 159.825 ;
        RECT 49.580 158.840 49.820 159.435 ;
        RECT 49.990 158.905 50.160 159.605 ;
        RECT 50.330 159.245 50.500 160.025 ;
        RECT 50.820 159.975 51.190 160.475 ;
        RECT 51.370 160.025 51.775 160.195 ;
        RECT 51.945 160.025 52.730 160.195 ;
        RECT 51.370 159.795 51.540 160.025 ;
        RECT 50.710 159.495 51.540 159.795 ;
        RECT 51.925 159.525 52.390 159.855 ;
        RECT 50.710 159.465 50.910 159.495 ;
        RECT 51.030 159.245 51.200 159.315 ;
        RECT 50.330 159.075 51.200 159.245 ;
        RECT 50.690 158.985 51.200 159.075 ;
        RECT 49.240 158.520 49.545 158.650 ;
        RECT 49.990 158.540 50.520 158.905 ;
        RECT 48.860 157.925 49.125 158.385 ;
        RECT 49.295 158.095 49.545 158.520 ;
        RECT 50.690 158.370 50.860 158.985 ;
        RECT 49.755 158.200 50.860 158.370 ;
        RECT 51.030 157.925 51.200 158.725 ;
        RECT 51.370 158.425 51.540 159.495 ;
        RECT 51.710 158.595 51.900 159.315 ;
        RECT 52.070 158.565 52.390 159.525 ;
        RECT 52.560 159.565 52.730 160.025 ;
        RECT 53.005 159.945 53.215 160.475 ;
        RECT 53.475 159.735 53.805 160.260 ;
        RECT 53.975 159.865 54.145 160.475 ;
        RECT 54.315 159.820 54.645 160.255 ;
        RECT 54.315 159.735 54.695 159.820 ;
        RECT 53.605 159.565 53.805 159.735 ;
        RECT 54.470 159.695 54.695 159.735 ;
        RECT 52.560 159.235 53.435 159.565 ;
        RECT 53.605 159.235 54.355 159.565 ;
        RECT 51.370 158.095 51.620 158.425 ;
        RECT 52.560 158.395 52.730 159.235 ;
        RECT 53.605 159.030 53.795 159.235 ;
        RECT 54.525 159.115 54.695 159.695 ;
        RECT 54.865 159.725 56.075 160.475 ;
        RECT 54.865 159.185 55.385 159.725 ;
        RECT 54.480 159.065 54.695 159.115 ;
        RECT 52.900 158.655 53.795 159.030 ;
        RECT 54.305 158.985 54.695 159.065 ;
        RECT 55.555 159.015 56.075 159.555 ;
        RECT 51.845 158.225 52.730 158.395 ;
        RECT 52.910 157.925 53.225 158.425 ;
        RECT 53.455 158.095 53.795 158.655 ;
        RECT 53.965 157.925 54.135 158.935 ;
        RECT 54.305 158.140 54.635 158.985 ;
        RECT 54.865 157.925 56.075 159.015 ;
        RECT 56.245 159.530 56.585 160.305 ;
        RECT 56.755 160.015 56.925 160.475 ;
        RECT 57.165 160.040 57.525 160.305 ;
        RECT 57.165 160.035 57.520 160.040 ;
        RECT 57.165 160.025 57.515 160.035 ;
        RECT 57.165 160.020 57.510 160.025 ;
        RECT 57.165 160.010 57.505 160.020 ;
        RECT 58.155 160.015 58.325 160.475 ;
        RECT 57.165 160.005 57.500 160.010 ;
        RECT 57.165 159.995 57.490 160.005 ;
        RECT 57.165 159.985 57.480 159.995 ;
        RECT 57.165 159.845 57.465 159.985 ;
        RECT 56.755 159.655 57.465 159.845 ;
        RECT 57.655 159.845 57.985 159.925 ;
        RECT 58.495 159.845 58.835 160.305 ;
        RECT 59.005 159.930 64.350 160.475 ;
        RECT 57.655 159.655 58.835 159.845 ;
        RECT 56.245 158.095 56.525 159.530 ;
        RECT 56.755 159.085 57.040 159.655 ;
        RECT 57.225 159.255 57.695 159.485 ;
        RECT 57.865 159.465 58.195 159.485 ;
        RECT 57.865 159.285 58.315 159.465 ;
        RECT 58.505 159.285 58.835 159.485 ;
        RECT 56.755 158.870 57.905 159.085 ;
        RECT 56.695 157.925 57.405 158.700 ;
        RECT 57.575 158.095 57.905 158.870 ;
        RECT 58.100 158.170 58.315 159.285 ;
        RECT 58.605 158.945 58.835 159.285 ;
        RECT 60.590 159.100 60.930 159.930 ;
        RECT 64.985 159.750 65.275 160.475 ;
        RECT 65.445 159.930 70.790 160.475 ;
        RECT 58.495 157.925 58.825 158.645 ;
        RECT 62.410 158.360 62.760 159.610 ;
        RECT 67.030 159.100 67.370 159.930 ;
        RECT 70.965 159.705 72.635 160.475 ;
        RECT 73.355 159.925 73.525 160.215 ;
        RECT 73.695 160.095 74.025 160.475 ;
        RECT 73.355 159.755 74.020 159.925 ;
        RECT 59.005 157.925 64.350 158.360 ;
        RECT 64.985 157.925 65.275 159.090 ;
        RECT 68.850 158.360 69.200 159.610 ;
        RECT 70.965 159.185 71.715 159.705 ;
        RECT 71.885 159.015 72.635 159.535 ;
        RECT 65.445 157.925 70.790 158.360 ;
        RECT 70.965 157.925 72.635 159.015 ;
        RECT 73.270 158.935 73.620 159.585 ;
        RECT 73.790 158.765 74.020 159.755 ;
        RECT 73.355 158.595 74.020 158.765 ;
        RECT 73.355 158.095 73.525 158.595 ;
        RECT 73.695 157.925 74.025 158.425 ;
        RECT 74.195 158.095 74.380 160.215 ;
        RECT 74.635 160.015 74.885 160.475 ;
        RECT 75.055 160.025 75.390 160.195 ;
        RECT 75.585 160.025 76.260 160.195 ;
        RECT 75.055 159.885 75.225 160.025 ;
        RECT 74.550 158.895 74.830 159.845 ;
        RECT 75.000 159.755 75.225 159.885 ;
        RECT 75.000 158.650 75.170 159.755 ;
        RECT 75.395 159.605 75.920 159.825 ;
        RECT 75.340 158.840 75.580 159.435 ;
        RECT 75.750 158.905 75.920 159.605 ;
        RECT 76.090 159.245 76.260 160.025 ;
        RECT 76.580 159.975 76.950 160.475 ;
        RECT 77.130 160.025 77.535 160.195 ;
        RECT 77.705 160.025 78.490 160.195 ;
        RECT 77.130 159.795 77.300 160.025 ;
        RECT 76.470 159.495 77.300 159.795 ;
        RECT 77.685 159.525 78.150 159.855 ;
        RECT 76.470 159.465 76.670 159.495 ;
        RECT 76.790 159.245 76.960 159.315 ;
        RECT 76.090 159.075 76.960 159.245 ;
        RECT 76.450 158.985 76.960 159.075 ;
        RECT 75.000 158.520 75.305 158.650 ;
        RECT 75.750 158.540 76.280 158.905 ;
        RECT 74.620 157.925 74.885 158.385 ;
        RECT 75.055 158.095 75.305 158.520 ;
        RECT 76.450 158.370 76.620 158.985 ;
        RECT 75.515 158.200 76.620 158.370 ;
        RECT 76.790 157.925 76.960 158.725 ;
        RECT 77.130 158.425 77.300 159.495 ;
        RECT 77.470 158.595 77.660 159.315 ;
        RECT 77.830 158.565 78.150 159.525 ;
        RECT 78.320 159.565 78.490 160.025 ;
        RECT 78.765 159.945 78.975 160.475 ;
        RECT 79.235 159.735 79.565 160.260 ;
        RECT 79.735 159.865 79.905 160.475 ;
        RECT 80.075 159.820 80.405 160.255 ;
        RECT 80.625 159.930 85.970 160.475 ;
        RECT 80.075 159.735 80.455 159.820 ;
        RECT 79.365 159.565 79.565 159.735 ;
        RECT 80.230 159.695 80.455 159.735 ;
        RECT 78.320 159.235 79.195 159.565 ;
        RECT 79.365 159.235 80.115 159.565 ;
        RECT 77.130 158.095 77.380 158.425 ;
        RECT 78.320 158.395 78.490 159.235 ;
        RECT 79.365 159.030 79.555 159.235 ;
        RECT 80.285 159.115 80.455 159.695 ;
        RECT 80.240 159.065 80.455 159.115 ;
        RECT 82.210 159.100 82.550 159.930 ;
        RECT 86.145 159.705 89.655 160.475 ;
        RECT 90.745 159.725 91.955 160.475 ;
        RECT 78.660 158.655 79.555 159.030 ;
        RECT 80.065 158.985 80.455 159.065 ;
        RECT 77.605 158.225 78.490 158.395 ;
        RECT 78.670 157.925 78.985 158.425 ;
        RECT 79.215 158.095 79.555 158.655 ;
        RECT 79.725 157.925 79.895 158.935 ;
        RECT 80.065 158.140 80.395 158.985 ;
        RECT 84.030 158.360 84.380 159.610 ;
        RECT 86.145 159.185 87.795 159.705 ;
        RECT 87.965 159.015 89.655 159.535 ;
        RECT 80.625 157.925 85.970 158.360 ;
        RECT 86.145 157.925 89.655 159.015 ;
        RECT 90.745 159.015 91.265 159.555 ;
        RECT 91.435 159.185 91.955 159.725 ;
        RECT 100.140 159.370 100.810 161.630 ;
        RECT 101.480 161.060 105.520 161.230 ;
        RECT 101.140 160.000 101.310 161.000 ;
        RECT 105.690 160.000 105.860 161.000 ;
        RECT 101.480 159.770 105.520 159.940 ;
        RECT 106.200 159.370 106.370 161.630 ;
        RECT 100.140 159.200 106.370 159.370 ;
        RECT 90.745 157.925 91.955 159.015 ;
        RECT 13.380 157.755 92.040 157.925 ;
        RECT 13.465 156.665 14.675 157.755 ;
        RECT 14.845 157.320 20.190 157.755 ;
        RECT 20.365 157.320 25.710 157.755 ;
        RECT 13.465 155.955 13.985 156.495 ;
        RECT 14.155 156.125 14.675 156.665 ;
        RECT 13.465 155.205 14.675 155.955 ;
        RECT 16.430 155.750 16.770 156.580 ;
        RECT 18.250 156.070 18.600 157.320 ;
        RECT 21.950 155.750 22.290 156.580 ;
        RECT 23.770 156.070 24.120 157.320 ;
        RECT 26.345 156.590 26.635 157.755 ;
        RECT 26.805 156.615 27.065 157.755 ;
        RECT 27.235 156.605 27.565 157.585 ;
        RECT 27.735 156.615 28.015 157.755 ;
        RECT 28.185 156.665 31.695 157.755 ;
        RECT 31.865 156.665 33.075 157.755 ;
        RECT 26.825 156.195 27.160 156.445 ;
        RECT 27.330 156.005 27.500 156.605 ;
        RECT 27.670 156.175 28.005 156.445 ;
        RECT 14.845 155.205 20.190 155.750 ;
        RECT 20.365 155.205 25.710 155.750 ;
        RECT 26.345 155.205 26.635 155.930 ;
        RECT 26.805 155.375 27.500 156.005 ;
        RECT 27.705 155.205 28.015 156.005 ;
        RECT 28.185 155.975 29.835 156.495 ;
        RECT 30.005 156.145 31.695 156.665 ;
        RECT 28.185 155.205 31.695 155.975 ;
        RECT 31.865 155.955 32.385 156.495 ;
        RECT 32.555 156.125 33.075 156.665 ;
        RECT 33.245 157.035 33.705 157.585 ;
        RECT 33.895 157.035 34.225 157.755 ;
        RECT 31.865 155.205 33.075 155.955 ;
        RECT 33.245 155.665 33.495 157.035 ;
        RECT 34.425 156.865 34.725 157.415 ;
        RECT 34.895 157.085 35.175 157.755 ;
        RECT 33.785 156.695 34.725 156.865 ;
        RECT 33.785 156.445 33.955 156.695 ;
        RECT 35.095 156.445 35.360 156.805 ;
        RECT 35.545 156.665 39.055 157.755 ;
        RECT 39.225 156.665 40.435 157.755 ;
        RECT 33.665 156.115 33.955 156.445 ;
        RECT 34.125 156.195 34.465 156.445 ;
        RECT 34.685 156.195 35.360 156.445 ;
        RECT 33.785 156.025 33.955 156.115 ;
        RECT 33.785 155.835 35.175 156.025 ;
        RECT 33.245 155.375 33.805 155.665 ;
        RECT 33.975 155.205 34.225 155.665 ;
        RECT 34.845 155.475 35.175 155.835 ;
        RECT 35.545 155.975 37.195 156.495 ;
        RECT 37.365 156.145 39.055 156.665 ;
        RECT 35.545 155.205 39.055 155.975 ;
        RECT 39.225 155.955 39.745 156.495 ;
        RECT 39.915 156.125 40.435 156.665 ;
        RECT 40.605 156.615 40.865 157.585 ;
        RECT 41.060 157.345 41.390 157.755 ;
        RECT 41.590 157.165 41.760 157.585 ;
        RECT 41.975 157.345 42.645 157.755 ;
        RECT 42.880 157.165 43.050 157.585 ;
        RECT 43.355 157.315 43.685 157.755 ;
        RECT 41.035 156.995 43.050 157.165 ;
        RECT 43.855 157.135 44.030 157.585 ;
        RECT 39.225 155.205 40.435 155.955 ;
        RECT 40.605 155.925 40.775 156.615 ;
        RECT 41.035 156.445 41.205 156.995 ;
        RECT 40.945 156.115 41.205 156.445 ;
        RECT 40.605 155.460 40.945 155.925 ;
        RECT 41.375 155.785 41.715 156.815 ;
        RECT 41.905 155.715 42.175 156.815 ;
        RECT 40.610 155.415 40.945 155.460 ;
        RECT 41.115 155.205 41.445 155.585 ;
        RECT 41.905 155.545 42.215 155.715 ;
        RECT 41.905 155.540 42.175 155.545 ;
        RECT 42.400 155.540 42.680 156.815 ;
        RECT 42.880 155.705 43.050 156.995 ;
        RECT 43.400 156.965 44.030 157.135 ;
        RECT 43.400 156.445 43.570 156.965 ;
        RECT 43.220 156.115 43.570 156.445 ;
        RECT 43.750 156.115 44.115 156.795 ;
        RECT 44.285 156.665 45.495 157.755 ;
        RECT 45.750 157.135 45.925 157.585 ;
        RECT 46.095 157.315 46.425 157.755 ;
        RECT 46.730 157.165 46.900 157.585 ;
        RECT 47.135 157.345 47.805 157.755 ;
        RECT 48.020 157.165 48.190 157.585 ;
        RECT 48.390 157.345 48.720 157.755 ;
        RECT 45.750 156.965 46.380 157.135 ;
        RECT 43.400 155.945 43.570 156.115 ;
        RECT 44.285 155.955 44.805 156.495 ;
        RECT 44.975 156.125 45.495 156.665 ;
        RECT 45.665 156.115 46.030 156.795 ;
        RECT 46.210 156.445 46.380 156.965 ;
        RECT 46.730 156.995 48.745 157.165 ;
        RECT 46.210 156.115 46.560 156.445 ;
        RECT 43.400 155.775 44.030 155.945 ;
        RECT 42.880 155.375 43.110 155.705 ;
        RECT 43.355 155.205 43.685 155.585 ;
        RECT 43.855 155.375 44.030 155.775 ;
        RECT 44.285 155.205 45.495 155.955 ;
        RECT 46.210 155.945 46.380 156.115 ;
        RECT 45.750 155.775 46.380 155.945 ;
        RECT 45.750 155.375 45.925 155.775 ;
        RECT 46.730 155.705 46.900 156.995 ;
        RECT 46.095 155.205 46.425 155.585 ;
        RECT 46.670 155.375 46.900 155.705 ;
        RECT 47.100 155.540 47.380 156.815 ;
        RECT 47.605 155.715 47.875 156.815 ;
        RECT 48.065 155.785 48.405 156.815 ;
        RECT 48.575 156.445 48.745 156.995 ;
        RECT 48.915 156.615 49.175 157.585 ;
        RECT 49.345 156.665 51.935 157.755 ;
        RECT 48.575 156.115 48.835 156.445 ;
        RECT 49.005 155.925 49.175 156.615 ;
        RECT 47.565 155.545 47.875 155.715 ;
        RECT 47.605 155.540 47.875 155.545 ;
        RECT 48.335 155.205 48.665 155.585 ;
        RECT 48.835 155.460 49.175 155.925 ;
        RECT 49.345 155.975 50.555 156.495 ;
        RECT 50.725 156.145 51.935 156.665 ;
        RECT 52.105 156.590 52.395 157.755 ;
        RECT 52.565 156.665 54.235 157.755 ;
        RECT 52.565 155.975 53.315 156.495 ;
        RECT 53.485 156.145 54.235 156.665 ;
        RECT 54.405 156.915 54.665 157.585 ;
        RECT 54.835 157.355 55.165 157.755 ;
        RECT 56.035 157.355 56.435 157.755 ;
        RECT 56.725 157.175 57.055 157.410 ;
        RECT 54.975 157.005 57.055 157.175 ;
        RECT 48.835 155.415 49.170 155.460 ;
        RECT 49.345 155.205 51.935 155.975 ;
        RECT 52.105 155.205 52.395 155.930 ;
        RECT 52.565 155.205 54.235 155.975 ;
        RECT 54.405 155.945 54.580 156.915 ;
        RECT 54.975 156.735 55.145 157.005 ;
        RECT 54.750 156.565 55.145 156.735 ;
        RECT 55.315 156.615 56.330 156.835 ;
        RECT 54.750 156.115 54.920 156.565 ;
        RECT 56.055 156.475 56.330 156.615 ;
        RECT 56.500 156.615 57.055 157.005 ;
        RECT 55.090 156.195 55.540 156.395 ;
        RECT 55.710 156.025 55.885 156.220 ;
        RECT 54.405 155.375 54.745 155.945 ;
        RECT 54.940 155.205 55.110 155.870 ;
        RECT 55.390 155.855 55.885 156.025 ;
        RECT 55.390 155.715 55.610 155.855 ;
        RECT 55.385 155.545 55.610 155.715 ;
        RECT 56.055 155.685 56.225 156.475 ;
        RECT 56.500 156.365 56.670 156.615 ;
        RECT 57.225 156.445 57.400 157.545 ;
        RECT 57.570 156.935 57.915 157.755 ;
        RECT 56.475 156.195 56.670 156.365 ;
        RECT 56.840 156.195 57.400 156.445 ;
        RECT 57.570 156.195 57.915 156.765 ;
        RECT 58.085 156.615 58.360 157.585 ;
        RECT 58.570 156.955 58.850 157.755 ;
        RECT 59.020 157.415 61.070 157.535 ;
        RECT 59.020 157.245 61.075 157.415 ;
        RECT 59.020 156.905 60.650 157.075 ;
        RECT 59.020 156.785 59.190 156.905 ;
        RECT 58.530 156.615 59.190 156.785 ;
        RECT 56.475 155.810 56.645 156.195 ;
        RECT 55.390 155.500 55.610 155.545 ;
        RECT 55.780 155.515 56.225 155.685 ;
        RECT 56.395 155.440 56.645 155.810 ;
        RECT 56.815 155.845 57.915 156.025 ;
        RECT 56.815 155.440 57.065 155.845 ;
        RECT 57.235 155.205 57.405 155.675 ;
        RECT 57.575 155.440 57.915 155.845 ;
        RECT 58.085 155.880 58.255 156.615 ;
        RECT 58.530 156.445 58.700 156.615 ;
        RECT 58.425 156.115 58.700 156.445 ;
        RECT 58.870 156.115 59.250 156.445 ;
        RECT 59.420 156.115 60.160 156.735 ;
        RECT 60.330 156.615 60.650 156.905 ;
        RECT 60.845 156.445 61.085 157.040 ;
        RECT 61.255 156.680 61.595 157.755 ;
        RECT 61.770 156.805 62.035 157.575 ;
        RECT 62.205 157.035 62.535 157.755 ;
        RECT 62.725 157.215 62.985 157.575 ;
        RECT 63.155 157.385 63.485 157.755 ;
        RECT 63.655 157.215 63.915 157.575 ;
        RECT 62.725 156.985 63.915 157.215 ;
        RECT 64.485 156.805 64.775 157.575 ;
        RECT 65.005 157.245 65.305 157.755 ;
        RECT 65.475 157.245 65.855 157.415 ;
        RECT 66.435 157.245 67.065 157.755 ;
        RECT 65.475 157.075 65.645 157.245 ;
        RECT 67.235 157.075 67.565 157.585 ;
        RECT 67.735 157.245 68.035 157.755 ;
        RECT 68.225 157.245 68.525 157.755 ;
        RECT 68.695 157.245 69.075 157.415 ;
        RECT 69.655 157.245 70.285 157.755 ;
        RECT 68.695 157.075 68.865 157.245 ;
        RECT 70.455 157.075 70.785 157.585 ;
        RECT 70.955 157.245 71.255 157.755 ;
        RECT 60.430 156.115 61.085 156.445 ;
        RECT 58.530 155.945 58.700 156.115 ;
        RECT 58.085 155.535 58.360 155.880 ;
        RECT 58.530 155.775 60.115 155.945 ;
        RECT 58.550 155.205 58.930 155.605 ;
        RECT 59.100 155.425 59.270 155.775 ;
        RECT 59.440 155.205 59.770 155.605 ;
        RECT 59.945 155.425 60.115 155.775 ;
        RECT 60.315 155.205 60.645 155.705 ;
        RECT 60.840 155.425 61.085 156.115 ;
        RECT 61.255 155.875 61.595 156.445 ;
        RECT 61.255 155.205 61.595 155.705 ;
        RECT 61.770 155.385 62.105 156.805 ;
        RECT 62.280 156.625 64.775 156.805 ;
        RECT 64.985 156.875 65.645 157.075 ;
        RECT 65.815 156.905 68.035 157.075 ;
        RECT 62.280 155.935 62.505 156.625 ;
        RECT 62.705 156.115 62.985 156.445 ;
        RECT 63.165 156.115 63.740 156.445 ;
        RECT 63.920 156.115 64.355 156.445 ;
        RECT 64.535 156.115 64.805 156.445 ;
        RECT 64.985 155.945 65.155 156.875 ;
        RECT 65.815 156.705 65.985 156.905 ;
        RECT 65.325 156.535 65.985 156.705 ;
        RECT 66.155 156.565 67.695 156.735 ;
        RECT 65.325 156.115 65.495 156.535 ;
        RECT 66.155 156.365 66.325 156.565 ;
        RECT 65.725 156.195 66.325 156.365 ;
        RECT 66.495 156.195 67.190 156.395 ;
        RECT 67.450 156.115 67.695 156.565 ;
        RECT 65.815 155.945 66.725 156.025 ;
        RECT 62.280 155.745 64.765 155.935 ;
        RECT 62.285 155.205 63.030 155.575 ;
        RECT 63.595 155.385 63.850 155.745 ;
        RECT 64.030 155.205 64.360 155.575 ;
        RECT 64.540 155.385 64.765 155.745 ;
        RECT 64.985 155.465 65.305 155.945 ;
        RECT 65.475 155.855 66.725 155.945 ;
        RECT 65.475 155.775 65.985 155.855 ;
        RECT 65.475 155.375 65.705 155.775 ;
        RECT 65.875 155.205 66.225 155.595 ;
        RECT 66.395 155.375 66.725 155.855 ;
        RECT 66.895 155.205 67.065 156.025 ;
        RECT 67.865 155.945 68.035 156.905 ;
        RECT 67.570 155.400 68.035 155.945 ;
        RECT 68.205 156.875 68.865 157.075 ;
        RECT 69.035 156.905 71.255 157.075 ;
        RECT 68.205 155.945 68.375 156.875 ;
        RECT 69.035 156.705 69.205 156.905 ;
        RECT 68.545 156.535 69.205 156.705 ;
        RECT 69.375 156.565 70.915 156.735 ;
        RECT 68.545 156.115 68.715 156.535 ;
        RECT 69.375 156.365 69.545 156.565 ;
        RECT 68.945 156.195 69.545 156.365 ;
        RECT 69.715 156.195 70.410 156.395 ;
        RECT 70.670 156.115 70.915 156.565 ;
        RECT 69.035 155.945 69.945 156.025 ;
        RECT 68.205 155.465 68.525 155.945 ;
        RECT 68.695 155.855 69.945 155.945 ;
        RECT 68.695 155.775 69.205 155.855 ;
        RECT 68.695 155.375 68.925 155.775 ;
        RECT 69.095 155.205 69.445 155.595 ;
        RECT 69.615 155.375 69.945 155.855 ;
        RECT 70.115 155.205 70.285 156.025 ;
        RECT 71.085 155.945 71.255 156.905 ;
        RECT 71.895 156.615 72.225 157.755 ;
        RECT 72.755 156.785 73.085 157.570 ;
        RECT 73.350 157.135 73.525 157.585 ;
        RECT 73.695 157.315 74.025 157.755 ;
        RECT 74.330 157.165 74.500 157.585 ;
        RECT 74.735 157.345 75.405 157.755 ;
        RECT 75.620 157.165 75.790 157.585 ;
        RECT 75.990 157.345 76.320 157.755 ;
        RECT 73.350 156.965 73.980 157.135 ;
        RECT 72.405 156.615 73.085 156.785 ;
        RECT 71.885 156.195 72.235 156.445 ;
        RECT 72.405 156.015 72.575 156.615 ;
        RECT 72.745 156.195 73.095 156.445 ;
        RECT 73.265 156.115 73.630 156.795 ;
        RECT 73.810 156.445 73.980 156.965 ;
        RECT 74.330 156.995 76.345 157.165 ;
        RECT 73.810 156.115 74.160 156.445 ;
        RECT 70.790 155.400 71.255 155.945 ;
        RECT 71.895 155.205 72.165 156.015 ;
        RECT 72.335 155.375 72.665 156.015 ;
        RECT 72.835 155.205 73.075 156.015 ;
        RECT 73.810 155.945 73.980 156.115 ;
        RECT 73.350 155.775 73.980 155.945 ;
        RECT 73.350 155.375 73.525 155.775 ;
        RECT 74.330 155.705 74.500 156.995 ;
        RECT 73.695 155.205 74.025 155.585 ;
        RECT 74.270 155.375 74.500 155.705 ;
        RECT 74.700 155.540 74.980 156.815 ;
        RECT 75.205 156.395 75.475 156.815 ;
        RECT 75.165 156.225 75.475 156.395 ;
        RECT 75.205 155.540 75.475 156.225 ;
        RECT 75.665 155.785 76.005 156.815 ;
        RECT 76.175 156.445 76.345 156.995 ;
        RECT 76.515 156.615 76.775 157.585 ;
        RECT 76.175 156.115 76.435 156.445 ;
        RECT 76.605 155.925 76.775 156.615 ;
        RECT 77.865 156.590 78.155 157.755 ;
        RECT 78.415 157.085 78.585 157.585 ;
        RECT 78.755 157.255 79.085 157.755 ;
        RECT 78.415 156.915 79.080 157.085 ;
        RECT 78.330 156.095 78.680 156.745 ;
        RECT 75.935 155.205 76.265 155.585 ;
        RECT 76.435 155.460 76.775 155.925 ;
        RECT 76.435 155.415 76.770 155.460 ;
        RECT 77.865 155.205 78.155 155.930 ;
        RECT 78.850 155.925 79.080 156.915 ;
        RECT 78.415 155.755 79.080 155.925 ;
        RECT 78.415 155.465 78.585 155.755 ;
        RECT 78.755 155.205 79.085 155.585 ;
        RECT 79.255 155.465 79.440 157.585 ;
        RECT 79.680 157.295 79.945 157.755 ;
        RECT 80.115 157.160 80.365 157.585 ;
        RECT 80.575 157.310 81.680 157.480 ;
        RECT 80.060 157.030 80.365 157.160 ;
        RECT 79.610 155.835 79.890 156.785 ;
        RECT 80.060 155.925 80.230 157.030 ;
        RECT 80.400 156.245 80.640 156.840 ;
        RECT 80.810 156.775 81.340 157.140 ;
        RECT 80.810 156.075 80.980 156.775 ;
        RECT 81.510 156.695 81.680 157.310 ;
        RECT 81.850 156.955 82.020 157.755 ;
        RECT 82.190 157.255 82.440 157.585 ;
        RECT 82.665 157.285 83.550 157.455 ;
        RECT 81.510 156.605 82.020 156.695 ;
        RECT 80.060 155.795 80.285 155.925 ;
        RECT 80.455 155.855 80.980 156.075 ;
        RECT 81.150 156.435 82.020 156.605 ;
        RECT 79.695 155.205 79.945 155.665 ;
        RECT 80.115 155.655 80.285 155.795 ;
        RECT 81.150 155.655 81.320 156.435 ;
        RECT 81.850 156.365 82.020 156.435 ;
        RECT 81.530 156.185 81.730 156.215 ;
        RECT 82.190 156.185 82.360 157.255 ;
        RECT 82.530 156.365 82.720 157.085 ;
        RECT 81.530 155.885 82.360 156.185 ;
        RECT 82.890 156.155 83.210 157.115 ;
        RECT 80.115 155.485 80.450 155.655 ;
        RECT 80.645 155.485 81.320 155.655 ;
        RECT 81.640 155.205 82.010 155.705 ;
        RECT 82.190 155.655 82.360 155.885 ;
        RECT 82.745 155.825 83.210 156.155 ;
        RECT 83.380 156.445 83.550 157.285 ;
        RECT 83.730 157.255 84.045 157.755 ;
        RECT 84.275 157.025 84.615 157.585 ;
        RECT 83.720 156.650 84.615 157.025 ;
        RECT 84.785 156.745 84.955 157.755 ;
        RECT 84.425 156.445 84.615 156.650 ;
        RECT 85.125 156.695 85.455 157.540 ;
        RECT 85.125 156.615 85.515 156.695 ;
        RECT 85.685 156.665 89.195 157.755 ;
        RECT 89.365 156.665 90.575 157.755 ;
        RECT 85.300 156.565 85.515 156.615 ;
        RECT 83.380 156.115 84.255 156.445 ;
        RECT 84.425 156.115 85.175 156.445 ;
        RECT 83.380 155.655 83.550 156.115 ;
        RECT 84.425 155.945 84.625 156.115 ;
        RECT 85.345 155.985 85.515 156.565 ;
        RECT 85.290 155.945 85.515 155.985 ;
        RECT 82.190 155.485 82.595 155.655 ;
        RECT 82.765 155.485 83.550 155.655 ;
        RECT 83.825 155.205 84.035 155.735 ;
        RECT 84.295 155.420 84.625 155.945 ;
        RECT 85.135 155.860 85.515 155.945 ;
        RECT 85.685 155.975 87.335 156.495 ;
        RECT 87.505 156.145 89.195 156.665 ;
        RECT 84.795 155.205 84.965 155.815 ;
        RECT 85.135 155.425 85.465 155.860 ;
        RECT 85.685 155.205 89.195 155.975 ;
        RECT 89.365 155.955 89.885 156.495 ;
        RECT 90.055 156.125 90.575 156.665 ;
        RECT 90.745 156.665 91.955 157.755 ;
        RECT 90.745 156.125 91.265 156.665 ;
        RECT 91.435 155.955 91.955 156.495 ;
        RECT 89.365 155.205 90.575 155.955 ;
        RECT 90.745 155.205 91.955 155.955 ;
        RECT 100.140 155.940 100.810 159.200 ;
        RECT 101.480 158.630 105.520 158.800 ;
        RECT 101.140 156.570 101.310 158.570 ;
        RECT 105.690 156.570 105.860 158.570 ;
        RECT 101.480 156.340 105.520 156.510 ;
        RECT 106.200 155.940 106.370 159.200 ;
        RECT 100.140 155.770 106.370 155.940 ;
        RECT 13.380 155.035 92.040 155.205 ;
        RECT 13.465 154.285 14.675 155.035 ;
        RECT 14.845 154.490 20.190 155.035 ;
        RECT 13.465 153.745 13.985 154.285 ;
        RECT 14.155 153.575 14.675 154.115 ;
        RECT 16.430 153.660 16.770 154.490 ;
        RECT 20.365 154.265 22.035 155.035 ;
        RECT 22.665 154.655 23.555 154.825 ;
        RECT 13.465 152.485 14.675 153.575 ;
        RECT 18.250 152.920 18.600 154.170 ;
        RECT 20.365 153.745 21.115 154.265 ;
        RECT 22.665 154.100 23.215 154.485 ;
        RECT 21.285 153.575 22.035 154.095 ;
        RECT 23.385 153.930 23.555 154.655 ;
        RECT 14.845 152.485 20.190 152.920 ;
        RECT 20.365 152.485 22.035 153.575 ;
        RECT 22.665 153.860 23.555 153.930 ;
        RECT 23.725 154.355 23.945 154.815 ;
        RECT 24.115 154.495 24.365 155.035 ;
        RECT 24.535 154.385 24.795 154.865 ;
        RECT 23.725 154.330 23.975 154.355 ;
        RECT 23.725 153.905 24.055 154.330 ;
        RECT 22.665 153.835 23.560 153.860 ;
        RECT 22.665 153.820 23.570 153.835 ;
        RECT 22.665 153.805 23.575 153.820 ;
        RECT 22.665 153.800 23.585 153.805 ;
        RECT 22.665 153.790 23.590 153.800 ;
        RECT 22.665 153.780 23.595 153.790 ;
        RECT 22.665 153.775 23.605 153.780 ;
        RECT 22.665 153.765 23.615 153.775 ;
        RECT 22.665 153.760 23.625 153.765 ;
        RECT 22.665 153.310 22.925 153.760 ;
        RECT 23.290 153.755 23.625 153.760 ;
        RECT 23.290 153.750 23.640 153.755 ;
        RECT 23.290 153.740 23.655 153.750 ;
        RECT 23.290 153.735 23.680 153.740 ;
        RECT 24.225 153.735 24.455 154.130 ;
        RECT 23.290 153.730 24.455 153.735 ;
        RECT 23.320 153.695 24.455 153.730 ;
        RECT 23.355 153.670 24.455 153.695 ;
        RECT 23.385 153.640 24.455 153.670 ;
        RECT 23.405 153.610 24.455 153.640 ;
        RECT 23.425 153.580 24.455 153.610 ;
        RECT 23.495 153.570 24.455 153.580 ;
        RECT 23.520 153.560 24.455 153.570 ;
        RECT 23.540 153.545 24.455 153.560 ;
        RECT 23.560 153.530 24.455 153.545 ;
        RECT 23.565 153.520 24.350 153.530 ;
        RECT 23.580 153.485 24.350 153.520 ;
        RECT 23.095 153.165 23.425 153.410 ;
        RECT 23.595 153.235 24.350 153.485 ;
        RECT 24.625 153.355 24.795 154.385 ;
        RECT 23.095 153.140 23.280 153.165 ;
        RECT 22.665 153.040 23.280 153.140 ;
        RECT 22.665 152.485 23.270 153.040 ;
        RECT 23.445 152.655 23.925 152.995 ;
        RECT 24.095 152.485 24.350 153.030 ;
        RECT 24.520 152.655 24.795 153.355 ;
        RECT 25.000 154.295 25.615 154.865 ;
        RECT 25.785 154.525 26.000 155.035 ;
        RECT 26.230 154.525 26.510 154.855 ;
        RECT 26.690 154.525 26.930 155.035 ;
        RECT 25.000 153.275 25.315 154.295 ;
        RECT 25.485 153.625 25.655 154.125 ;
        RECT 25.905 153.795 26.170 154.355 ;
        RECT 26.340 153.625 26.510 154.525 ;
        RECT 27.355 154.485 27.525 154.775 ;
        RECT 27.695 154.655 28.025 155.035 ;
        RECT 26.680 153.795 27.035 154.355 ;
        RECT 27.355 154.315 28.020 154.485 ;
        RECT 25.485 153.455 26.910 153.625 ;
        RECT 27.270 153.495 27.620 154.145 ;
        RECT 25.000 152.655 25.535 153.275 ;
        RECT 25.705 152.485 26.035 153.285 ;
        RECT 26.520 153.280 26.910 153.455 ;
        RECT 27.790 153.325 28.020 154.315 ;
        RECT 27.355 153.155 28.020 153.325 ;
        RECT 27.355 152.655 27.525 153.155 ;
        RECT 27.695 152.485 28.025 152.985 ;
        RECT 28.195 152.655 28.380 154.775 ;
        RECT 28.635 154.575 28.885 155.035 ;
        RECT 29.055 154.585 29.390 154.755 ;
        RECT 29.585 154.585 30.260 154.755 ;
        RECT 29.055 154.445 29.225 154.585 ;
        RECT 28.550 153.455 28.830 154.405 ;
        RECT 29.000 154.315 29.225 154.445 ;
        RECT 29.000 153.210 29.170 154.315 ;
        RECT 29.395 154.165 29.920 154.385 ;
        RECT 29.340 153.400 29.580 153.995 ;
        RECT 29.750 153.465 29.920 154.165 ;
        RECT 30.090 153.805 30.260 154.585 ;
        RECT 30.580 154.535 30.950 155.035 ;
        RECT 31.130 154.585 31.535 154.755 ;
        RECT 31.705 154.585 32.490 154.755 ;
        RECT 31.130 154.355 31.300 154.585 ;
        RECT 30.470 154.055 31.300 154.355 ;
        RECT 31.685 154.085 32.150 154.415 ;
        RECT 30.470 154.025 30.670 154.055 ;
        RECT 30.790 153.805 30.960 153.875 ;
        RECT 30.090 153.635 30.960 153.805 ;
        RECT 30.450 153.545 30.960 153.635 ;
        RECT 29.000 153.080 29.305 153.210 ;
        RECT 29.750 153.100 30.280 153.465 ;
        RECT 28.620 152.485 28.885 152.945 ;
        RECT 29.055 152.655 29.305 153.080 ;
        RECT 30.450 152.930 30.620 153.545 ;
        RECT 29.515 152.760 30.620 152.930 ;
        RECT 30.790 152.485 30.960 153.285 ;
        RECT 31.130 152.985 31.300 154.055 ;
        RECT 31.470 153.155 31.660 153.875 ;
        RECT 31.830 153.125 32.150 154.085 ;
        RECT 32.320 154.125 32.490 154.585 ;
        RECT 32.765 154.505 32.975 155.035 ;
        RECT 33.235 154.295 33.565 154.820 ;
        RECT 33.735 154.425 33.905 155.035 ;
        RECT 34.075 154.380 34.405 154.815 ;
        RECT 34.075 154.295 34.455 154.380 ;
        RECT 33.365 154.125 33.565 154.295 ;
        RECT 34.230 154.255 34.455 154.295 ;
        RECT 32.320 153.795 33.195 154.125 ;
        RECT 33.365 153.795 34.115 154.125 ;
        RECT 31.130 152.655 31.380 152.985 ;
        RECT 32.320 152.955 32.490 153.795 ;
        RECT 33.365 153.590 33.555 153.795 ;
        RECT 34.285 153.675 34.455 154.255 ;
        RECT 34.625 154.265 38.135 155.035 ;
        RECT 39.225 154.310 39.515 155.035 ;
        RECT 39.685 154.490 45.030 155.035 ;
        RECT 34.625 153.745 36.275 154.265 ;
        RECT 34.240 153.625 34.455 153.675 ;
        RECT 32.660 153.215 33.555 153.590 ;
        RECT 34.065 153.545 34.455 153.625 ;
        RECT 36.445 153.575 38.135 154.095 ;
        RECT 41.270 153.660 41.610 154.490 ;
        RECT 45.205 154.265 48.715 155.035 ;
        RECT 48.885 154.285 50.095 155.035 ;
        RECT 31.605 152.785 32.490 152.955 ;
        RECT 32.670 152.485 32.985 152.985 ;
        RECT 33.215 152.655 33.555 153.215 ;
        RECT 33.725 152.485 33.895 153.495 ;
        RECT 34.065 152.700 34.395 153.545 ;
        RECT 34.625 152.485 38.135 153.575 ;
        RECT 39.225 152.485 39.515 153.650 ;
        RECT 43.090 152.920 43.440 154.170 ;
        RECT 45.205 153.745 46.855 154.265 ;
        RECT 47.025 153.575 48.715 154.095 ;
        RECT 48.885 153.745 49.405 154.285 ;
        RECT 50.285 154.225 50.525 155.035 ;
        RECT 50.695 154.225 51.025 154.865 ;
        RECT 51.195 154.225 51.465 155.035 ;
        RECT 51.645 154.295 52.085 154.855 ;
        RECT 52.255 154.295 52.705 155.035 ;
        RECT 52.875 154.465 53.045 154.865 ;
        RECT 53.215 154.635 53.635 155.035 ;
        RECT 53.805 154.465 54.035 154.865 ;
        RECT 52.875 154.295 54.035 154.465 ;
        RECT 54.205 154.295 54.695 154.865 ;
        RECT 54.875 154.535 55.205 155.035 ;
        RECT 55.405 154.465 55.575 154.815 ;
        RECT 55.775 154.635 56.105 155.035 ;
        RECT 56.275 154.465 56.445 154.815 ;
        RECT 56.615 154.635 56.995 155.035 ;
        RECT 49.575 153.575 50.095 154.115 ;
        RECT 50.265 153.795 50.615 154.045 ;
        RECT 50.785 153.625 50.955 154.225 ;
        RECT 51.125 153.795 51.475 154.045 ;
        RECT 39.685 152.485 45.030 152.920 ;
        RECT 45.205 152.485 48.715 153.575 ;
        RECT 48.885 152.485 50.095 153.575 ;
        RECT 50.275 153.455 50.955 153.625 ;
        RECT 50.275 152.670 50.605 153.455 ;
        RECT 51.135 152.485 51.465 153.625 ;
        RECT 51.645 153.285 51.955 154.295 ;
        RECT 52.125 153.675 52.295 154.125 ;
        RECT 52.465 153.845 52.855 154.125 ;
        RECT 53.040 153.795 53.285 154.125 ;
        RECT 52.125 153.505 52.915 153.675 ;
        RECT 51.645 152.655 52.085 153.285 ;
        RECT 52.260 152.485 52.575 153.335 ;
        RECT 52.745 152.825 52.915 153.505 ;
        RECT 53.085 152.995 53.285 153.795 ;
        RECT 53.485 152.995 53.735 154.125 ;
        RECT 53.950 153.795 54.355 154.125 ;
        RECT 54.525 153.625 54.695 154.295 ;
        RECT 54.870 153.795 55.220 154.365 ;
        RECT 55.405 154.295 57.015 154.465 ;
        RECT 57.185 154.360 57.455 154.705 ;
        RECT 56.845 154.125 57.015 154.295 ;
        RECT 55.390 153.675 56.100 154.125 ;
        RECT 56.270 153.795 56.675 154.125 ;
        RECT 56.845 153.795 57.115 154.125 ;
        RECT 53.925 153.455 54.695 153.625 ;
        RECT 53.925 152.825 54.175 153.455 ;
        RECT 54.870 153.335 55.190 153.625 ;
        RECT 55.385 153.505 56.100 153.675 ;
        RECT 56.845 153.625 57.015 153.795 ;
        RECT 57.285 153.625 57.455 154.360 ;
        RECT 57.625 154.265 61.135 155.035 ;
        RECT 62.230 154.360 62.505 154.705 ;
        RECT 62.695 154.635 63.075 155.035 ;
        RECT 63.245 154.465 63.415 154.815 ;
        RECT 63.585 154.635 63.915 155.035 ;
        RECT 64.085 154.465 64.340 154.815 ;
        RECT 57.625 153.745 59.275 154.265 ;
        RECT 56.290 153.455 57.015 153.625 ;
        RECT 56.290 153.335 56.460 153.455 ;
        RECT 52.745 152.655 54.175 152.825 ;
        RECT 54.355 152.485 54.685 153.285 ;
        RECT 54.870 153.165 56.460 153.335 ;
        RECT 54.870 152.705 56.525 152.995 ;
        RECT 56.695 152.485 56.975 153.285 ;
        RECT 57.185 152.655 57.455 153.625 ;
        RECT 59.445 153.575 61.135 154.095 ;
        RECT 57.625 152.485 61.135 153.575 ;
        RECT 62.230 153.625 62.400 154.360 ;
        RECT 62.675 154.295 64.340 154.465 ;
        RECT 64.985 154.310 65.275 155.035 ;
        RECT 66.370 154.360 66.645 154.705 ;
        RECT 66.835 154.635 67.215 155.035 ;
        RECT 67.385 154.465 67.555 154.815 ;
        RECT 67.725 154.635 68.055 155.035 ;
        RECT 68.225 154.465 68.480 154.815 ;
        RECT 62.675 154.125 62.845 154.295 ;
        RECT 62.570 153.795 62.845 154.125 ;
        RECT 63.015 153.795 63.840 154.125 ;
        RECT 64.010 153.795 64.355 154.125 ;
        RECT 62.675 153.625 62.845 153.795 ;
        RECT 62.230 152.655 62.505 153.625 ;
        RECT 62.675 153.455 63.335 153.625 ;
        RECT 63.645 153.505 63.840 153.795 ;
        RECT 63.165 153.335 63.335 153.455 ;
        RECT 64.010 153.335 64.335 153.625 ;
        RECT 62.715 152.485 62.995 153.285 ;
        RECT 63.165 153.165 64.335 153.335 ;
        RECT 63.165 152.705 64.355 152.995 ;
        RECT 64.985 152.485 65.275 153.650 ;
        RECT 66.370 153.625 66.540 154.360 ;
        RECT 66.815 154.295 68.480 154.465 ;
        RECT 69.585 154.315 69.925 154.825 ;
        RECT 66.815 154.125 66.985 154.295 ;
        RECT 66.710 153.795 66.985 154.125 ;
        RECT 67.155 153.795 67.980 154.125 ;
        RECT 68.150 153.795 68.495 154.125 ;
        RECT 66.815 153.625 66.985 153.795 ;
        RECT 66.370 152.655 66.645 153.625 ;
        RECT 66.815 153.455 67.475 153.625 ;
        RECT 67.785 153.505 67.980 153.795 ;
        RECT 67.305 153.335 67.475 153.455 ;
        RECT 68.150 153.335 68.475 153.625 ;
        RECT 66.855 152.485 67.135 153.285 ;
        RECT 67.305 153.165 68.475 153.335 ;
        RECT 67.305 152.705 68.495 152.995 ;
        RECT 69.585 152.915 69.845 154.315 ;
        RECT 70.095 154.235 70.365 155.035 ;
        RECT 70.020 153.795 70.350 154.045 ;
        RECT 70.545 153.795 70.825 154.765 ;
        RECT 71.005 153.795 71.305 154.765 ;
        RECT 71.485 153.795 71.835 154.760 ;
        RECT 72.055 154.535 72.550 154.865 ;
        RECT 70.035 153.625 70.350 153.795 ;
        RECT 72.055 153.625 72.225 154.535 ;
        RECT 70.035 153.455 72.225 153.625 ;
        RECT 69.585 152.655 69.925 152.915 ;
        RECT 70.095 152.485 70.425 153.285 ;
        RECT 70.890 152.655 71.140 153.455 ;
        RECT 71.325 152.485 71.655 153.205 ;
        RECT 71.875 152.655 72.125 153.455 ;
        RECT 72.395 153.045 72.635 154.355 ;
        RECT 72.805 154.265 74.475 155.035 ;
        RECT 74.645 154.385 74.905 154.865 ;
        RECT 75.075 154.495 75.325 155.035 ;
        RECT 72.805 153.745 73.555 154.265 ;
        RECT 73.725 153.575 74.475 154.095 ;
        RECT 72.295 152.485 72.630 152.865 ;
        RECT 72.805 152.485 74.475 153.575 ;
        RECT 74.645 153.355 74.815 154.385 ;
        RECT 75.495 154.355 75.715 154.815 ;
        RECT 75.465 154.330 75.715 154.355 ;
        RECT 74.985 153.735 75.215 154.130 ;
        RECT 75.385 153.905 75.715 154.330 ;
        RECT 75.885 154.655 76.775 154.825 ;
        RECT 75.885 153.930 76.055 154.655 ;
        RECT 76.225 154.100 76.775 154.485 ;
        RECT 76.955 154.305 77.255 155.035 ;
        RECT 77.435 154.125 77.665 154.745 ;
        RECT 77.865 154.475 78.090 154.855 ;
        RECT 78.260 154.645 78.590 155.035 ;
        RECT 78.785 154.490 84.130 155.035 ;
        RECT 84.305 154.490 89.650 155.035 ;
        RECT 77.865 154.295 78.195 154.475 ;
        RECT 75.885 153.860 76.775 153.930 ;
        RECT 75.880 153.835 76.775 153.860 ;
        RECT 75.870 153.820 76.775 153.835 ;
        RECT 75.865 153.805 76.775 153.820 ;
        RECT 75.855 153.800 76.775 153.805 ;
        RECT 75.850 153.790 76.775 153.800 ;
        RECT 76.960 153.795 77.255 154.125 ;
        RECT 77.435 153.795 77.850 154.125 ;
        RECT 75.845 153.780 76.775 153.790 ;
        RECT 75.835 153.775 76.775 153.780 ;
        RECT 75.825 153.765 76.775 153.775 ;
        RECT 75.815 153.760 76.775 153.765 ;
        RECT 75.815 153.755 76.150 153.760 ;
        RECT 75.800 153.750 76.150 153.755 ;
        RECT 75.785 153.740 76.150 153.750 ;
        RECT 75.760 153.735 76.150 153.740 ;
        RECT 74.985 153.730 76.150 153.735 ;
        RECT 74.985 153.695 76.120 153.730 ;
        RECT 74.985 153.670 76.085 153.695 ;
        RECT 74.985 153.640 76.055 153.670 ;
        RECT 74.985 153.610 76.035 153.640 ;
        RECT 74.985 153.580 76.015 153.610 ;
        RECT 74.985 153.570 75.945 153.580 ;
        RECT 74.985 153.560 75.920 153.570 ;
        RECT 74.985 153.545 75.900 153.560 ;
        RECT 74.985 153.530 75.880 153.545 ;
        RECT 75.090 153.520 75.875 153.530 ;
        RECT 75.090 153.485 75.860 153.520 ;
        RECT 74.645 152.655 74.920 153.355 ;
        RECT 75.090 153.235 75.845 153.485 ;
        RECT 76.015 153.165 76.345 153.410 ;
        RECT 76.515 153.310 76.775 153.760 ;
        RECT 78.020 153.625 78.195 154.295 ;
        RECT 78.365 153.795 78.605 154.445 ;
        RECT 80.370 153.660 80.710 154.490 ;
        RECT 76.160 153.140 76.345 153.165 ;
        RECT 76.955 153.265 77.850 153.595 ;
        RECT 78.020 153.435 78.605 153.625 ;
        RECT 76.160 153.040 76.775 153.140 ;
        RECT 75.090 152.485 75.345 153.030 ;
        RECT 75.515 152.655 75.995 152.995 ;
        RECT 76.170 152.485 76.775 153.040 ;
        RECT 76.955 153.095 78.160 153.265 ;
        RECT 76.955 152.665 77.285 153.095 ;
        RECT 77.465 152.485 77.660 152.925 ;
        RECT 77.830 152.665 78.160 153.095 ;
        RECT 78.330 152.665 78.605 153.435 ;
        RECT 82.190 152.920 82.540 154.170 ;
        RECT 85.890 153.660 86.230 154.490 ;
        RECT 90.745 154.285 91.955 155.035 ;
        RECT 87.710 152.920 88.060 154.170 ;
        RECT 90.745 153.575 91.265 154.115 ;
        RECT 91.435 153.745 91.955 154.285 ;
        RECT 78.785 152.485 84.130 152.920 ;
        RECT 84.305 152.485 89.650 152.920 ;
        RECT 90.745 152.485 91.955 153.575 ;
        RECT 100.140 152.510 100.810 155.770 ;
        RECT 101.480 155.200 105.520 155.370 ;
        RECT 101.140 153.140 101.310 155.140 ;
        RECT 105.690 153.140 105.860 155.140 ;
        RECT 101.480 152.910 105.520 153.080 ;
        RECT 106.200 152.510 106.370 155.770 ;
        RECT 100.140 152.500 106.370 152.510 ;
        RECT 107.960 161.770 117.790 161.810 ;
        RECT 120.510 161.790 126.250 161.800 ;
        RECT 107.960 161.640 118.590 161.770 ;
        RECT 107.960 159.380 108.130 161.640 ;
        RECT 108.855 161.070 116.895 161.240 ;
        RECT 108.470 160.010 108.640 161.010 ;
        RECT 117.110 160.010 117.280 161.010 ;
        RECT 108.855 159.780 116.895 159.950 ;
        RECT 117.620 159.380 118.590 161.640 ;
        RECT 107.960 159.210 118.590 159.380 ;
        RECT 107.960 155.950 108.130 159.210 ;
        RECT 108.855 158.640 116.895 158.810 ;
        RECT 108.470 156.580 108.640 158.580 ;
        RECT 117.110 156.580 117.280 158.580 ;
        RECT 108.855 156.350 116.895 156.520 ;
        RECT 117.620 155.950 118.590 159.210 ;
        RECT 107.960 155.780 118.590 155.950 ;
        RECT 107.960 152.520 108.130 155.780 ;
        RECT 108.855 155.210 116.895 155.380 ;
        RECT 108.470 153.150 108.640 155.150 ;
        RECT 117.110 153.150 117.280 155.150 ;
        RECT 108.855 152.920 116.895 153.090 ;
        RECT 117.620 152.520 118.590 155.780 ;
        RECT 13.380 152.315 92.040 152.485 ;
        RECT 100.140 152.400 106.380 152.500 ;
        RECT 13.465 151.225 14.675 152.315 ;
        RECT 14.845 151.225 18.355 152.315 ;
        RECT 19.075 151.645 19.245 152.145 ;
        RECT 19.415 151.815 19.745 152.315 ;
        RECT 19.075 151.475 19.740 151.645 ;
        RECT 13.465 150.515 13.985 151.055 ;
        RECT 14.155 150.685 14.675 151.225 ;
        RECT 14.845 150.535 16.495 151.055 ;
        RECT 16.665 150.705 18.355 151.225 ;
        RECT 18.990 150.655 19.340 151.305 ;
        RECT 13.465 149.765 14.675 150.515 ;
        RECT 14.845 149.765 18.355 150.535 ;
        RECT 19.510 150.485 19.740 151.475 ;
        RECT 19.075 150.315 19.740 150.485 ;
        RECT 19.075 150.025 19.245 150.315 ;
        RECT 19.415 149.765 19.745 150.145 ;
        RECT 19.915 150.025 20.100 152.145 ;
        RECT 20.340 151.855 20.605 152.315 ;
        RECT 20.775 151.720 21.025 152.145 ;
        RECT 21.235 151.870 22.340 152.040 ;
        RECT 20.720 151.590 21.025 151.720 ;
        RECT 20.270 150.395 20.550 151.345 ;
        RECT 20.720 150.485 20.890 151.590 ;
        RECT 21.060 150.805 21.300 151.400 ;
        RECT 21.470 151.335 22.000 151.700 ;
        RECT 21.470 150.635 21.640 151.335 ;
        RECT 22.170 151.255 22.340 151.870 ;
        RECT 22.510 151.515 22.680 152.315 ;
        RECT 22.850 151.815 23.100 152.145 ;
        RECT 23.325 151.845 24.210 152.015 ;
        RECT 22.170 151.165 22.680 151.255 ;
        RECT 20.720 150.355 20.945 150.485 ;
        RECT 21.115 150.415 21.640 150.635 ;
        RECT 21.810 150.995 22.680 151.165 ;
        RECT 20.355 149.765 20.605 150.225 ;
        RECT 20.775 150.215 20.945 150.355 ;
        RECT 21.810 150.215 21.980 150.995 ;
        RECT 22.510 150.925 22.680 150.995 ;
        RECT 22.190 150.745 22.390 150.775 ;
        RECT 22.850 150.745 23.020 151.815 ;
        RECT 23.190 150.925 23.380 151.645 ;
        RECT 22.190 150.445 23.020 150.745 ;
        RECT 23.550 150.715 23.870 151.675 ;
        RECT 20.775 150.045 21.110 150.215 ;
        RECT 21.305 150.045 21.980 150.215 ;
        RECT 22.300 149.765 22.670 150.265 ;
        RECT 22.850 150.215 23.020 150.445 ;
        RECT 23.405 150.385 23.870 150.715 ;
        RECT 24.040 151.005 24.210 151.845 ;
        RECT 24.390 151.815 24.705 152.315 ;
        RECT 24.935 151.585 25.275 152.145 ;
        RECT 24.380 151.210 25.275 151.585 ;
        RECT 25.445 151.305 25.615 152.315 ;
        RECT 25.085 151.005 25.275 151.210 ;
        RECT 25.785 151.255 26.115 152.100 ;
        RECT 25.785 151.175 26.175 151.255 ;
        RECT 25.960 151.125 26.175 151.175 ;
        RECT 26.345 151.150 26.635 152.315 ;
        RECT 24.040 150.675 24.915 151.005 ;
        RECT 25.085 150.675 25.835 151.005 ;
        RECT 24.040 150.215 24.210 150.675 ;
        RECT 25.085 150.505 25.285 150.675 ;
        RECT 26.005 150.545 26.175 151.125 ;
        RECT 25.950 150.505 26.175 150.545 ;
        RECT 22.850 150.045 23.255 150.215 ;
        RECT 23.425 150.045 24.210 150.215 ;
        RECT 24.485 149.765 24.695 150.295 ;
        RECT 24.955 149.980 25.285 150.505 ;
        RECT 25.795 150.420 26.175 150.505 ;
        RECT 25.455 149.765 25.625 150.375 ;
        RECT 25.795 149.985 26.125 150.420 ;
        RECT 26.345 149.765 26.635 150.490 ;
        RECT 26.815 149.945 27.075 152.135 ;
        RECT 27.245 151.585 27.585 152.315 ;
        RECT 27.765 151.405 28.035 152.135 ;
        RECT 27.265 151.185 28.035 151.405 ;
        RECT 28.215 151.425 28.445 152.135 ;
        RECT 28.615 151.605 28.945 152.315 ;
        RECT 29.115 151.425 29.375 152.135 ;
        RECT 28.215 151.185 29.375 151.425 ;
        RECT 29.565 151.225 32.155 152.315 ;
        RECT 27.265 150.515 27.555 151.185 ;
        RECT 27.735 150.695 28.200 151.005 ;
        RECT 28.380 150.695 28.905 151.005 ;
        RECT 27.265 150.315 28.495 150.515 ;
        RECT 27.335 149.765 28.005 150.135 ;
        RECT 28.185 149.945 28.495 150.315 ;
        RECT 28.675 150.055 28.905 150.695 ;
        RECT 29.085 150.675 29.385 151.005 ;
        RECT 29.565 150.535 30.775 151.055 ;
        RECT 30.945 150.705 32.155 151.225 ;
        RECT 32.415 151.305 32.585 152.145 ;
        RECT 32.755 151.975 33.925 152.145 ;
        RECT 32.755 151.475 33.085 151.975 ;
        RECT 33.595 151.935 33.925 151.975 ;
        RECT 34.115 151.895 34.470 152.315 ;
        RECT 33.255 151.715 33.485 151.805 ;
        RECT 34.640 151.715 34.890 152.145 ;
        RECT 33.255 151.475 34.890 151.715 ;
        RECT 35.060 151.555 35.390 152.315 ;
        RECT 35.560 151.475 35.815 152.145 ;
        RECT 32.415 151.135 35.475 151.305 ;
        RECT 32.330 150.755 32.680 150.965 ;
        RECT 32.850 150.755 33.295 150.955 ;
        RECT 33.465 150.755 33.940 150.955 ;
        RECT 29.085 149.765 29.375 150.495 ;
        RECT 29.565 149.765 32.155 150.535 ;
        RECT 32.415 150.415 33.480 150.585 ;
        RECT 32.415 149.935 32.585 150.415 ;
        RECT 32.755 149.765 33.085 150.245 ;
        RECT 33.310 150.185 33.480 150.415 ;
        RECT 33.660 150.355 33.940 150.755 ;
        RECT 34.210 150.755 34.540 150.955 ;
        RECT 34.710 150.785 35.085 150.955 ;
        RECT 34.710 150.755 35.075 150.785 ;
        RECT 34.210 150.355 34.495 150.755 ;
        RECT 35.305 150.585 35.475 151.135 ;
        RECT 34.675 150.415 35.475 150.585 ;
        RECT 34.675 150.185 34.845 150.415 ;
        RECT 35.645 150.345 35.815 151.475 ;
        RECT 36.005 151.225 37.215 152.315 ;
        RECT 37.885 151.855 38.100 152.315 ;
        RECT 38.270 151.685 38.600 152.145 ;
        RECT 35.630 150.275 35.815 150.345 ;
        RECT 35.605 150.265 35.815 150.275 ;
        RECT 33.310 149.935 34.845 150.185 ;
        RECT 35.015 149.765 35.345 150.245 ;
        RECT 35.560 149.935 35.815 150.265 ;
        RECT 36.005 150.515 36.525 151.055 ;
        RECT 36.695 150.685 37.215 151.225 ;
        RECT 37.430 151.515 38.600 151.685 ;
        RECT 38.770 151.515 39.020 152.315 ;
        RECT 36.005 149.765 37.215 150.515 ;
        RECT 37.430 150.225 37.800 151.515 ;
        RECT 39.230 151.345 39.510 151.505 ;
        RECT 38.175 151.175 39.510 151.345 ;
        RECT 40.145 151.465 40.525 152.145 ;
        RECT 41.115 151.465 41.285 152.315 ;
        RECT 41.455 151.635 41.785 152.145 ;
        RECT 41.955 151.805 42.125 152.315 ;
        RECT 42.295 151.635 42.695 152.145 ;
        RECT 41.455 151.465 42.695 151.635 ;
        RECT 38.175 151.005 38.345 151.175 ;
        RECT 37.970 150.755 38.345 151.005 ;
        RECT 38.515 150.755 38.990 150.995 ;
        RECT 39.160 150.755 39.510 150.995 ;
        RECT 38.175 150.585 38.345 150.755 ;
        RECT 38.175 150.415 39.510 150.585 ;
        RECT 37.430 149.935 38.180 150.225 ;
        RECT 38.690 149.765 39.020 150.225 ;
        RECT 39.240 150.205 39.510 150.415 ;
        RECT 40.145 150.505 40.315 151.465 ;
        RECT 40.485 151.125 41.790 151.295 ;
        RECT 42.875 151.215 43.195 152.145 ;
        RECT 43.365 151.225 44.575 152.315 ;
        RECT 44.745 151.805 45.045 152.315 ;
        RECT 45.215 151.635 45.545 152.145 ;
        RECT 45.715 151.805 46.345 152.315 ;
        RECT 46.925 151.805 47.305 151.975 ;
        RECT 47.475 151.805 47.775 152.315 ;
        RECT 47.135 151.635 47.305 151.805 ;
        RECT 40.485 150.675 40.730 151.125 ;
        RECT 40.900 150.755 41.450 150.955 ;
        RECT 41.620 150.925 41.790 151.125 ;
        RECT 42.565 151.045 43.195 151.215 ;
        RECT 41.620 150.755 41.995 150.925 ;
        RECT 42.165 150.505 42.395 151.005 ;
        RECT 40.145 150.335 42.395 150.505 ;
        RECT 40.195 149.765 40.525 150.155 ;
        RECT 40.695 150.015 40.865 150.335 ;
        RECT 42.565 150.165 42.735 151.045 ;
        RECT 41.035 149.765 41.365 150.155 ;
        RECT 41.780 149.995 42.735 150.165 ;
        RECT 42.905 149.765 43.195 150.600 ;
        RECT 43.365 150.515 43.885 151.055 ;
        RECT 44.055 150.685 44.575 151.225 ;
        RECT 44.745 151.465 46.965 151.635 ;
        RECT 43.365 149.765 44.575 150.515 ;
        RECT 44.745 150.505 44.915 151.465 ;
        RECT 45.085 151.125 46.625 151.295 ;
        RECT 45.085 150.675 45.330 151.125 ;
        RECT 45.590 150.755 46.285 150.955 ;
        RECT 46.455 150.925 46.625 151.125 ;
        RECT 46.795 151.265 46.965 151.465 ;
        RECT 47.135 151.435 47.795 151.635 ;
        RECT 46.795 151.095 47.455 151.265 ;
        RECT 46.455 150.755 47.055 150.925 ;
        RECT 47.285 150.675 47.455 151.095 ;
        RECT 44.745 149.960 45.210 150.505 ;
        RECT 45.715 149.765 45.885 150.585 ;
        RECT 46.055 150.505 46.965 150.585 ;
        RECT 47.625 150.505 47.795 151.435 ;
        RECT 47.965 151.225 49.175 152.315 ;
        RECT 49.350 151.805 51.005 152.095 ;
        RECT 46.055 150.415 47.305 150.505 ;
        RECT 46.055 149.935 46.385 150.415 ;
        RECT 46.795 150.335 47.305 150.415 ;
        RECT 46.555 149.765 46.905 150.155 ;
        RECT 47.075 149.935 47.305 150.335 ;
        RECT 47.475 150.025 47.795 150.505 ;
        RECT 47.965 150.515 48.485 151.055 ;
        RECT 48.655 150.685 49.175 151.225 ;
        RECT 49.350 151.465 50.940 151.635 ;
        RECT 51.175 151.515 51.455 152.315 ;
        RECT 49.350 151.175 49.670 151.465 ;
        RECT 50.770 151.345 50.940 151.465 ;
        RECT 47.965 149.765 49.175 150.515 ;
        RECT 49.350 150.435 49.700 151.005 ;
        RECT 49.870 150.675 50.580 151.295 ;
        RECT 50.770 151.175 51.495 151.345 ;
        RECT 51.665 151.175 51.935 152.145 ;
        RECT 51.325 151.005 51.495 151.175 ;
        RECT 50.750 150.675 51.155 151.005 ;
        RECT 51.325 150.675 51.595 151.005 ;
        RECT 51.325 150.505 51.495 150.675 ;
        RECT 49.885 150.335 51.495 150.505 ;
        RECT 51.765 150.440 51.935 151.175 ;
        RECT 52.105 151.150 52.395 152.315 ;
        RECT 52.570 151.345 52.865 152.315 ;
        RECT 53.435 151.955 53.765 152.315 ;
        RECT 53.935 151.955 55.915 152.145 ;
        RECT 53.035 151.785 53.255 151.870 ;
        RECT 53.935 151.785 54.115 151.955 ;
        RECT 56.095 151.875 56.365 152.315 ;
        RECT 56.915 151.955 57.245 152.315 ;
        RECT 57.760 151.955 58.090 152.315 ;
        RECT 58.600 151.955 58.935 152.315 ;
        RECT 59.835 151.955 60.165 152.315 ;
        RECT 53.035 151.615 54.115 151.785 ;
        RECT 54.285 151.705 55.950 151.785 ;
        RECT 56.525 151.705 60.160 151.785 ;
        RECT 53.035 151.540 53.255 151.615 ;
        RECT 54.285 151.535 60.160 151.705 ;
        RECT 53.445 151.195 56.110 151.365 ;
        RECT 53.445 151.010 53.890 151.195 ;
        RECT 52.880 150.755 53.890 151.010 ;
        RECT 54.185 150.755 55.660 151.025 ;
        RECT 55.830 150.675 56.110 151.195 ;
        RECT 56.740 151.195 59.480 151.365 ;
        RECT 56.740 151.090 57.455 151.195 ;
        RECT 56.280 150.675 57.455 151.090 ;
        RECT 57.850 150.755 58.920 151.025 ;
        RECT 59.310 150.675 59.480 151.195 ;
        RECT 59.650 151.020 60.160 151.535 ;
        RECT 60.475 151.305 60.645 152.145 ;
        RECT 60.815 151.975 61.985 152.145 ;
        RECT 60.815 151.475 61.145 151.975 ;
        RECT 61.655 151.935 61.985 151.975 ;
        RECT 62.175 151.895 62.530 152.315 ;
        RECT 61.315 151.715 61.545 151.805 ;
        RECT 62.700 151.715 62.950 152.145 ;
        RECT 61.315 151.475 62.950 151.715 ;
        RECT 63.120 151.555 63.450 152.315 ;
        RECT 63.620 151.475 63.875 152.145 ;
        RECT 60.475 151.135 63.535 151.305 ;
        RECT 52.635 150.545 54.275 150.585 ;
        RECT 49.355 149.765 49.685 150.265 ;
        RECT 49.885 149.985 50.055 150.335 ;
        RECT 50.255 149.765 50.585 150.165 ;
        RECT 50.755 149.985 50.925 150.335 ;
        RECT 51.095 149.765 51.475 150.165 ;
        RECT 51.665 150.095 51.935 150.440 ;
        RECT 52.105 149.765 52.395 150.490 ;
        RECT 52.635 150.475 55.610 150.545 ;
        RECT 59.650 150.505 59.830 151.020 ;
        RECT 60.390 150.755 60.740 150.965 ;
        RECT 60.910 150.755 61.355 150.955 ;
        RECT 61.525 150.755 62.000 150.955 ;
        RECT 52.635 150.375 56.315 150.475 ;
        RECT 52.635 150.305 53.720 150.375 ;
        RECT 54.255 150.305 56.315 150.375 ;
        RECT 56.485 150.315 58.650 150.495 ;
        RECT 59.045 150.335 59.830 150.505 ;
        RECT 60.475 150.415 61.540 150.585 ;
        RECT 52.635 150.215 52.835 150.305 ;
        RECT 53.005 149.765 53.335 150.125 ;
        RECT 53.505 150.105 53.720 150.305 ;
        RECT 53.945 149.765 54.115 150.205 ;
        RECT 56.085 150.135 56.315 150.305 ;
        RECT 54.725 149.765 55.055 150.125 ;
        RECT 55.585 149.765 55.915 150.125 ;
        RECT 56.085 149.935 57.400 150.135 ;
        RECT 59.045 150.130 59.215 150.335 ;
        RECT 59.990 150.160 60.160 150.275 ;
        RECT 57.760 149.950 59.215 150.130 ;
        RECT 59.460 149.990 60.160 150.160 ;
        RECT 60.475 149.935 60.645 150.415 ;
        RECT 60.815 149.765 61.145 150.245 ;
        RECT 61.370 150.185 61.540 150.415 ;
        RECT 61.720 150.355 62.000 150.755 ;
        RECT 62.270 150.755 62.600 150.955 ;
        RECT 62.770 150.755 63.135 150.955 ;
        RECT 62.270 150.355 62.555 150.755 ;
        RECT 63.365 150.585 63.535 151.135 ;
        RECT 62.735 150.415 63.535 150.585 ;
        RECT 62.735 150.185 62.905 150.415 ;
        RECT 63.705 150.345 63.875 151.475 ;
        RECT 64.065 151.175 64.325 152.315 ;
        RECT 64.495 151.165 64.825 152.145 ;
        RECT 64.995 151.175 65.275 152.315 ;
        RECT 65.445 151.880 70.790 152.315 ;
        RECT 64.085 150.755 64.420 151.005 ;
        RECT 64.590 150.565 64.760 151.165 ;
        RECT 64.930 150.735 65.265 151.005 ;
        RECT 63.690 150.275 63.875 150.345 ;
        RECT 63.665 150.265 63.875 150.275 ;
        RECT 61.370 149.935 62.905 150.185 ;
        RECT 63.075 149.765 63.405 150.245 ;
        RECT 63.620 149.935 63.875 150.265 ;
        RECT 64.065 149.935 64.760 150.565 ;
        RECT 64.965 149.765 65.275 150.565 ;
        RECT 67.030 150.310 67.370 151.140 ;
        RECT 68.850 150.630 69.200 151.880 ;
        RECT 70.965 151.225 73.555 152.315 ;
        RECT 70.965 150.535 72.175 151.055 ;
        RECT 72.345 150.705 73.555 151.225 ;
        RECT 73.735 151.175 74.065 152.315 ;
        RECT 74.595 151.345 74.925 152.130 ;
        RECT 74.245 151.175 74.925 151.345 ;
        RECT 75.115 151.345 75.445 152.130 ;
        RECT 75.115 151.175 75.795 151.345 ;
        RECT 75.975 151.175 76.305 152.315 ;
        RECT 76.485 151.225 77.695 152.315 ;
        RECT 73.725 150.755 74.075 151.005 ;
        RECT 74.245 150.575 74.415 151.175 ;
        RECT 74.585 150.755 74.935 151.005 ;
        RECT 75.105 150.755 75.455 151.005 ;
        RECT 75.625 150.575 75.795 151.175 ;
        RECT 75.965 150.755 76.315 151.005 ;
        RECT 65.445 149.765 70.790 150.310 ;
        RECT 70.965 149.765 73.555 150.535 ;
        RECT 73.735 149.765 74.005 150.575 ;
        RECT 74.175 149.935 74.505 150.575 ;
        RECT 74.675 149.765 74.915 150.575 ;
        RECT 75.125 149.765 75.365 150.575 ;
        RECT 75.535 149.935 75.865 150.575 ;
        RECT 76.035 149.765 76.305 150.575 ;
        RECT 76.485 150.515 77.005 151.055 ;
        RECT 77.175 150.685 77.695 151.225 ;
        RECT 77.865 151.150 78.155 152.315 ;
        RECT 78.325 151.880 83.670 152.315 ;
        RECT 83.845 151.880 89.190 152.315 ;
        RECT 76.485 149.765 77.695 150.515 ;
        RECT 77.865 149.765 78.155 150.490 ;
        RECT 79.910 150.310 80.250 151.140 ;
        RECT 81.730 150.630 82.080 151.880 ;
        RECT 85.430 150.310 85.770 151.140 ;
        RECT 87.250 150.630 87.600 151.880 ;
        RECT 89.365 151.225 90.575 152.315 ;
        RECT 89.365 150.515 89.885 151.055 ;
        RECT 90.055 150.685 90.575 151.225 ;
        RECT 90.745 151.225 91.955 152.315 ;
        RECT 100.130 151.840 106.380 152.400 ;
        RECT 100.130 151.820 105.300 151.840 ;
        RECT 100.130 151.750 104.120 151.820 ;
        RECT 90.745 150.685 91.265 151.225 ;
        RECT 91.435 150.515 91.955 151.055 ;
        RECT 78.325 149.765 83.670 150.310 ;
        RECT 83.845 149.765 89.190 150.310 ;
        RECT 89.365 149.765 90.575 150.515 ;
        RECT 90.745 149.765 91.955 150.515 ;
        RECT 100.130 150.480 102.050 151.750 ;
        RECT 103.560 151.740 104.120 151.750 ;
        RECT 103.790 150.650 104.120 151.740 ;
        RECT 104.490 151.270 105.530 151.440 ;
        RECT 104.490 150.830 105.530 151.000 ;
        RECT 105.700 150.970 105.870 151.300 ;
        RECT 103.950 150.430 104.120 150.650 ;
        RECT 106.210 150.430 106.380 151.840 ;
        RECT 103.950 150.260 106.380 150.430 ;
        RECT 107.960 152.350 118.590 152.520 ;
        RECT 120.020 161.630 126.250 161.790 ;
        RECT 120.020 159.370 120.690 161.630 ;
        RECT 121.360 161.060 125.400 161.230 ;
        RECT 121.020 160.000 121.190 161.000 ;
        RECT 125.570 160.000 125.740 161.000 ;
        RECT 121.360 159.770 125.400 159.940 ;
        RECT 126.080 159.370 126.250 161.630 ;
        RECT 120.020 159.200 126.250 159.370 ;
        RECT 120.020 155.940 120.690 159.200 ;
        RECT 121.360 158.630 125.400 158.800 ;
        RECT 121.020 156.570 121.190 158.570 ;
        RECT 125.570 156.570 125.740 158.570 ;
        RECT 121.360 156.340 125.400 156.510 ;
        RECT 126.080 155.940 126.250 159.200 ;
        RECT 120.020 155.770 126.250 155.940 ;
        RECT 120.020 152.510 120.690 155.770 ;
        RECT 121.360 155.200 125.400 155.370 ;
        RECT 121.020 153.140 121.190 155.140 ;
        RECT 125.570 153.140 125.740 155.140 ;
        RECT 121.360 152.910 125.400 153.080 ;
        RECT 126.080 152.510 126.250 155.770 ;
        RECT 120.020 152.500 126.250 152.510 ;
        RECT 127.840 161.770 137.670 161.810 ;
        RECT 127.840 161.640 138.470 161.770 ;
        RECT 140.590 161.740 146.330 161.750 ;
        RECT 127.840 159.380 128.010 161.640 ;
        RECT 128.735 161.070 136.775 161.240 ;
        RECT 128.350 160.010 128.520 161.010 ;
        RECT 136.990 160.010 137.160 161.010 ;
        RECT 128.735 159.780 136.775 159.950 ;
        RECT 137.500 159.380 138.470 161.640 ;
        RECT 127.840 159.210 138.470 159.380 ;
        RECT 127.840 155.950 128.010 159.210 ;
        RECT 128.735 158.640 136.775 158.810 ;
        RECT 128.350 156.580 128.520 158.580 ;
        RECT 136.990 156.580 137.160 158.580 ;
        RECT 128.735 156.350 136.775 156.520 ;
        RECT 137.500 155.950 138.470 159.210 ;
        RECT 127.840 155.780 138.470 155.950 ;
        RECT 127.840 152.520 128.010 155.780 ;
        RECT 128.735 155.210 136.775 155.380 ;
        RECT 128.350 153.150 128.520 155.150 ;
        RECT 136.990 153.150 137.160 155.150 ;
        RECT 128.735 152.920 136.775 153.090 ;
        RECT 137.500 152.520 138.470 155.780 ;
        RECT 120.020 152.400 126.260 152.500 ;
        RECT 107.960 150.090 108.130 152.350 ;
        RECT 108.855 151.780 116.895 151.950 ;
        RECT 108.470 150.720 108.640 151.720 ;
        RECT 117.110 150.720 117.280 151.720 ;
        RECT 108.855 150.490 116.895 150.660 ;
        RECT 117.620 150.090 118.590 152.350 ;
        RECT 120.010 151.840 126.260 152.400 ;
        RECT 120.010 151.820 125.180 151.840 ;
        RECT 120.010 151.750 124.000 151.820 ;
        RECT 120.010 150.480 121.930 151.750 ;
        RECT 123.440 151.740 124.000 151.750 ;
        RECT 123.670 150.650 124.000 151.740 ;
        RECT 124.370 151.270 125.410 151.440 ;
        RECT 124.370 150.830 125.410 151.000 ;
        RECT 125.580 150.970 125.750 151.300 ;
        RECT 123.830 150.430 124.000 150.650 ;
        RECT 126.090 150.430 126.260 151.840 ;
        RECT 123.830 150.260 126.260 150.430 ;
        RECT 127.840 152.350 138.470 152.520 ;
        RECT 140.100 161.580 146.330 161.740 ;
        RECT 140.100 159.320 140.770 161.580 ;
        RECT 141.440 161.010 145.480 161.180 ;
        RECT 141.100 159.950 141.270 160.950 ;
        RECT 145.650 159.950 145.820 160.950 ;
        RECT 141.440 159.720 145.480 159.890 ;
        RECT 146.160 159.320 146.330 161.580 ;
        RECT 140.100 159.150 146.330 159.320 ;
        RECT 140.100 155.890 140.770 159.150 ;
        RECT 141.440 158.580 145.480 158.750 ;
        RECT 141.100 156.520 141.270 158.520 ;
        RECT 145.650 156.520 145.820 158.520 ;
        RECT 141.440 156.290 145.480 156.460 ;
        RECT 146.160 155.890 146.330 159.150 ;
        RECT 140.100 155.720 146.330 155.890 ;
        RECT 140.100 152.460 140.770 155.720 ;
        RECT 141.440 155.150 145.480 155.320 ;
        RECT 141.100 153.090 141.270 155.090 ;
        RECT 145.650 153.090 145.820 155.090 ;
        RECT 141.440 152.860 145.480 153.030 ;
        RECT 146.160 152.460 146.330 155.720 ;
        RECT 140.100 152.450 146.330 152.460 ;
        RECT 147.920 161.720 157.750 161.760 ;
        RECT 147.920 161.590 158.550 161.720 ;
        RECT 147.920 159.330 148.090 161.590 ;
        RECT 148.815 161.020 156.855 161.190 ;
        RECT 148.430 159.960 148.600 160.960 ;
        RECT 157.070 159.960 157.240 160.960 ;
        RECT 148.815 159.730 156.855 159.900 ;
        RECT 157.580 159.330 158.550 161.590 ;
        RECT 147.920 159.160 158.550 159.330 ;
        RECT 147.920 155.900 148.090 159.160 ;
        RECT 148.815 158.590 156.855 158.760 ;
        RECT 148.430 156.530 148.600 158.530 ;
        RECT 157.070 156.530 157.240 158.530 ;
        RECT 148.815 156.300 156.855 156.470 ;
        RECT 157.580 155.900 158.550 159.160 ;
        RECT 147.920 155.730 158.550 155.900 ;
        RECT 147.920 152.470 148.090 155.730 ;
        RECT 148.815 155.160 156.855 155.330 ;
        RECT 148.430 153.100 148.600 155.100 ;
        RECT 157.070 153.100 157.240 155.100 ;
        RECT 148.815 152.870 156.855 153.040 ;
        RECT 157.580 152.470 158.550 155.730 ;
        RECT 140.100 152.350 146.340 152.450 ;
        RECT 107.960 150.060 118.590 150.090 ;
        RECT 127.840 150.090 128.010 152.350 ;
        RECT 128.735 151.780 136.775 151.950 ;
        RECT 128.350 150.720 128.520 151.720 ;
        RECT 136.990 150.720 137.160 151.720 ;
        RECT 128.735 150.490 136.775 150.660 ;
        RECT 137.500 150.090 138.470 152.350 ;
        RECT 140.090 151.790 146.340 152.350 ;
        RECT 140.090 151.770 145.260 151.790 ;
        RECT 140.090 151.700 144.080 151.770 ;
        RECT 140.090 150.430 142.010 151.700 ;
        RECT 143.520 151.690 144.080 151.700 ;
        RECT 143.750 150.600 144.080 151.690 ;
        RECT 144.450 151.220 145.490 151.390 ;
        RECT 144.450 150.780 145.490 150.950 ;
        RECT 145.660 150.920 145.830 151.250 ;
        RECT 143.910 150.380 144.080 150.600 ;
        RECT 146.170 150.380 146.340 151.790 ;
        RECT 143.910 150.210 146.340 150.380 ;
        RECT 147.920 152.300 158.550 152.470 ;
        RECT 127.840 150.060 138.470 150.090 ;
        RECT 107.930 149.950 118.590 150.060 ;
        RECT 127.810 149.950 138.470 150.060 ;
        RECT 147.920 150.040 148.090 152.300 ;
        RECT 148.815 151.730 156.855 151.900 ;
        RECT 148.430 150.670 148.600 151.670 ;
        RECT 157.070 150.670 157.240 151.670 ;
        RECT 148.815 150.440 156.855 150.610 ;
        RECT 157.580 150.040 158.550 152.300 ;
        RECT 147.920 150.010 158.550 150.040 ;
        RECT 106.180 149.900 118.590 149.950 ;
        RECT 126.060 149.900 138.470 149.950 ;
        RECT 147.890 149.900 158.550 150.010 ;
        RECT 13.380 149.595 92.040 149.765 ;
        RECT 101.840 149.730 118.590 149.900 ;
        RECT 13.465 148.845 14.675 149.595 ;
        RECT 14.845 149.050 20.190 149.595 ;
        RECT 13.465 148.305 13.985 148.845 ;
        RECT 14.155 148.135 14.675 148.675 ;
        RECT 16.430 148.220 16.770 149.050 ;
        RECT 20.365 148.945 20.625 149.425 ;
        RECT 20.795 149.135 21.125 149.595 ;
        RECT 21.315 148.955 21.515 149.375 ;
        RECT 13.465 147.045 14.675 148.135 ;
        RECT 18.250 147.480 18.600 148.730 ;
        RECT 20.365 147.915 20.535 148.945 ;
        RECT 20.705 148.255 20.935 148.685 ;
        RECT 21.105 148.435 21.515 148.955 ;
        RECT 21.685 149.110 22.475 149.375 ;
        RECT 21.685 148.255 21.940 149.110 ;
        RECT 22.655 148.775 22.985 149.195 ;
        RECT 23.155 148.775 23.415 149.595 ;
        RECT 24.045 148.945 24.305 149.425 ;
        RECT 24.475 149.055 24.725 149.595 ;
        RECT 22.655 148.685 22.905 148.775 ;
        RECT 22.110 148.435 22.905 148.685 ;
        RECT 20.705 148.085 22.495 148.255 ;
        RECT 14.845 147.045 20.190 147.480 ;
        RECT 20.365 147.215 20.640 147.915 ;
        RECT 20.810 147.790 21.525 148.085 ;
        RECT 21.745 147.725 22.075 147.915 ;
        RECT 20.850 147.045 21.065 147.590 ;
        RECT 21.235 147.215 21.710 147.555 ;
        RECT 21.880 147.550 22.075 147.725 ;
        RECT 22.245 147.720 22.495 148.085 ;
        RECT 21.880 147.045 22.495 147.550 ;
        RECT 22.735 147.215 22.905 148.435 ;
        RECT 23.075 147.725 23.415 148.605 ;
        RECT 24.045 147.915 24.215 148.945 ;
        RECT 24.895 148.890 25.115 149.375 ;
        RECT 24.385 148.295 24.615 148.690 ;
        RECT 24.785 148.465 25.115 148.890 ;
        RECT 25.285 149.215 26.175 149.385 ;
        RECT 25.285 148.490 25.455 149.215 ;
        RECT 26.345 149.050 31.690 149.595 ;
        RECT 25.625 148.660 26.175 149.045 ;
        RECT 25.285 148.420 26.175 148.490 ;
        RECT 25.280 148.395 26.175 148.420 ;
        RECT 25.270 148.380 26.175 148.395 ;
        RECT 25.265 148.365 26.175 148.380 ;
        RECT 25.255 148.360 26.175 148.365 ;
        RECT 25.250 148.350 26.175 148.360 ;
        RECT 25.245 148.340 26.175 148.350 ;
        RECT 25.235 148.335 26.175 148.340 ;
        RECT 25.225 148.325 26.175 148.335 ;
        RECT 25.215 148.320 26.175 148.325 ;
        RECT 25.215 148.315 25.550 148.320 ;
        RECT 25.200 148.310 25.550 148.315 ;
        RECT 25.185 148.300 25.550 148.310 ;
        RECT 25.160 148.295 25.550 148.300 ;
        RECT 24.385 148.290 25.550 148.295 ;
        RECT 24.385 148.255 25.520 148.290 ;
        RECT 24.385 148.230 25.485 148.255 ;
        RECT 24.385 148.200 25.455 148.230 ;
        RECT 24.385 148.170 25.435 148.200 ;
        RECT 24.385 148.140 25.415 148.170 ;
        RECT 24.385 148.130 25.345 148.140 ;
        RECT 24.385 148.120 25.320 148.130 ;
        RECT 24.385 148.105 25.300 148.120 ;
        RECT 24.385 148.090 25.280 148.105 ;
        RECT 24.490 148.080 25.275 148.090 ;
        RECT 24.490 148.045 25.260 148.080 ;
        RECT 23.155 147.045 23.415 147.555 ;
        RECT 24.045 147.215 24.320 147.915 ;
        RECT 24.490 147.795 25.245 148.045 ;
        RECT 25.415 147.725 25.745 147.970 ;
        RECT 25.915 147.870 26.175 148.320 ;
        RECT 27.930 148.220 28.270 149.050 ;
        RECT 31.865 148.945 32.205 149.425 ;
        RECT 32.570 149.115 32.900 149.425 ;
        RECT 33.070 149.115 33.320 149.595 ;
        RECT 32.730 148.945 32.900 149.115 ;
        RECT 33.490 148.945 33.820 149.425 ;
        RECT 33.990 149.115 34.240 149.595 ;
        RECT 34.410 148.945 34.740 149.425 ;
        RECT 31.865 148.775 32.560 148.945 ;
        RECT 32.730 148.775 34.740 148.945 ;
        RECT 35.085 148.825 38.595 149.595 ;
        RECT 39.225 148.870 39.515 149.595 ;
        RECT 39.735 148.940 40.065 149.375 ;
        RECT 40.235 148.985 40.405 149.595 ;
        RECT 39.685 148.855 40.065 148.940 ;
        RECT 40.575 148.855 40.905 149.380 ;
        RECT 41.165 149.065 41.375 149.595 ;
        RECT 41.650 149.145 42.435 149.315 ;
        RECT 42.605 149.145 43.010 149.315 ;
        RECT 25.560 147.700 25.745 147.725 ;
        RECT 25.560 147.600 26.175 147.700 ;
        RECT 24.490 147.045 24.745 147.590 ;
        RECT 24.915 147.215 25.395 147.555 ;
        RECT 25.570 147.045 26.175 147.600 ;
        RECT 29.750 147.480 30.100 148.730 ;
        RECT 31.885 148.405 32.220 148.605 ;
        RECT 26.345 147.045 31.690 147.480 ;
        RECT 31.865 147.045 32.125 148.235 ;
        RECT 32.390 148.195 32.560 148.775 ;
        RECT 32.770 148.435 33.100 148.605 ;
        RECT 32.295 147.215 32.625 148.195 ;
        RECT 32.795 147.325 33.100 148.435 ;
        RECT 33.280 148.435 33.610 148.605 ;
        RECT 33.280 147.325 33.600 148.435 ;
        RECT 33.780 148.265 34.110 148.605 ;
        RECT 34.280 148.355 34.860 148.605 ;
        RECT 35.085 148.305 36.735 148.825 ;
        RECT 39.685 148.815 39.910 148.855 ;
        RECT 33.770 147.325 34.110 148.265 ;
        RECT 34.410 147.045 34.740 148.185 ;
        RECT 36.905 148.135 38.595 148.655 ;
        RECT 39.685 148.235 39.855 148.815 ;
        RECT 40.575 148.685 40.775 148.855 ;
        RECT 41.650 148.685 41.820 149.145 ;
        RECT 40.025 148.355 40.775 148.685 ;
        RECT 40.945 148.355 41.820 148.685 ;
        RECT 35.085 147.045 38.595 148.135 ;
        RECT 39.225 147.045 39.515 148.210 ;
        RECT 39.685 148.185 39.900 148.235 ;
        RECT 39.685 148.105 40.075 148.185 ;
        RECT 39.745 147.260 40.075 148.105 ;
        RECT 40.585 148.150 40.775 148.355 ;
        RECT 40.245 147.045 40.415 148.055 ;
        RECT 40.585 147.775 41.480 148.150 ;
        RECT 40.585 147.215 40.925 147.775 ;
        RECT 41.155 147.045 41.470 147.545 ;
        RECT 41.650 147.515 41.820 148.355 ;
        RECT 41.990 148.645 42.455 148.975 ;
        RECT 42.840 148.915 43.010 149.145 ;
        RECT 43.190 149.095 43.560 149.595 ;
        RECT 43.880 149.145 44.555 149.315 ;
        RECT 44.750 149.145 45.085 149.315 ;
        RECT 41.990 147.685 42.310 148.645 ;
        RECT 42.840 148.615 43.670 148.915 ;
        RECT 42.480 147.715 42.670 148.435 ;
        RECT 42.840 147.545 43.010 148.615 ;
        RECT 43.470 148.585 43.670 148.615 ;
        RECT 43.180 148.365 43.350 148.435 ;
        RECT 43.880 148.365 44.050 149.145 ;
        RECT 44.915 149.005 45.085 149.145 ;
        RECT 45.255 149.135 45.505 149.595 ;
        RECT 43.180 148.195 44.050 148.365 ;
        RECT 44.220 148.725 44.745 148.945 ;
        RECT 44.915 148.875 45.140 149.005 ;
        RECT 43.180 148.105 43.690 148.195 ;
        RECT 41.650 147.345 42.535 147.515 ;
        RECT 42.760 147.215 43.010 147.545 ;
        RECT 43.180 147.045 43.350 147.845 ;
        RECT 43.520 147.490 43.690 148.105 ;
        RECT 44.220 148.025 44.390 148.725 ;
        RECT 43.860 147.660 44.390 148.025 ;
        RECT 44.560 147.960 44.800 148.555 ;
        RECT 44.970 147.770 45.140 148.875 ;
        RECT 45.310 148.015 45.590 148.965 ;
        RECT 44.835 147.640 45.140 147.770 ;
        RECT 43.520 147.320 44.625 147.490 ;
        RECT 44.835 147.215 45.085 147.640 ;
        RECT 45.255 147.045 45.520 147.505 ;
        RECT 45.760 147.215 45.945 149.335 ;
        RECT 46.115 149.215 46.445 149.595 ;
        RECT 46.615 149.045 46.785 149.335 ;
        RECT 46.120 148.875 46.785 149.045 ;
        RECT 46.120 147.885 46.350 148.875 ;
        RECT 47.045 148.825 48.715 149.595 ;
        RECT 49.365 148.865 49.655 149.595 ;
        RECT 46.520 148.055 46.870 148.705 ;
        RECT 47.045 148.305 47.795 148.825 ;
        RECT 47.965 148.135 48.715 148.655 ;
        RECT 49.355 148.355 49.655 148.685 ;
        RECT 49.835 148.665 50.065 149.305 ;
        RECT 50.245 149.045 50.555 149.415 ;
        RECT 50.735 149.225 51.405 149.595 ;
        RECT 50.245 148.845 51.475 149.045 ;
        RECT 49.835 148.355 50.360 148.665 ;
        RECT 50.540 148.355 51.005 148.665 ;
        RECT 51.185 148.175 51.475 148.845 ;
        RECT 46.120 147.715 46.785 147.885 ;
        RECT 46.115 147.045 46.445 147.545 ;
        RECT 46.615 147.215 46.785 147.715 ;
        RECT 47.045 147.045 48.715 148.135 ;
        RECT 49.365 147.935 50.525 148.175 ;
        RECT 49.365 147.225 49.625 147.935 ;
        RECT 49.795 147.045 50.125 147.755 ;
        RECT 50.295 147.225 50.525 147.935 ;
        RECT 50.705 147.955 51.475 148.175 ;
        RECT 50.705 147.225 50.975 147.955 ;
        RECT 51.155 147.045 51.495 147.775 ;
        RECT 51.665 147.225 51.925 149.415 ;
        RECT 52.105 149.050 57.450 149.595 ;
        RECT 53.690 148.220 54.030 149.050 ;
        RECT 57.625 148.845 58.835 149.595 ;
        RECT 59.170 149.085 59.410 149.595 ;
        RECT 59.590 149.085 59.870 149.415 ;
        RECT 60.100 149.085 60.315 149.595 ;
        RECT 55.510 147.480 55.860 148.730 ;
        RECT 57.625 148.305 58.145 148.845 ;
        RECT 58.315 148.135 58.835 148.675 ;
        RECT 59.065 148.355 59.420 148.915 ;
        RECT 59.590 148.185 59.760 149.085 ;
        RECT 59.930 148.355 60.195 148.915 ;
        RECT 60.485 148.855 61.100 149.425 ;
        RECT 60.445 148.185 60.615 148.685 ;
        RECT 52.105 147.045 57.450 147.480 ;
        RECT 57.625 147.045 58.835 148.135 ;
        RECT 59.190 148.015 60.615 148.185 ;
        RECT 59.190 147.840 59.580 148.015 ;
        RECT 60.065 147.045 60.395 147.845 ;
        RECT 60.785 147.835 61.100 148.855 ;
        RECT 60.565 147.215 61.100 147.835 ;
        RECT 61.305 148.795 61.645 149.425 ;
        RECT 61.815 148.795 62.065 149.595 ;
        RECT 62.255 148.945 62.585 149.425 ;
        RECT 62.755 149.135 62.980 149.595 ;
        RECT 63.150 148.945 63.480 149.425 ;
        RECT 61.305 148.185 61.480 148.795 ;
        RECT 62.255 148.775 63.480 148.945 ;
        RECT 64.110 148.815 64.610 149.425 ;
        RECT 64.985 148.870 65.275 149.595 ;
        RECT 61.650 148.435 62.345 148.605 ;
        RECT 62.175 148.185 62.345 148.435 ;
        RECT 62.520 148.405 62.940 148.605 ;
        RECT 63.110 148.405 63.440 148.605 ;
        RECT 63.610 148.405 63.940 148.605 ;
        RECT 64.110 148.185 64.280 148.815 ;
        RECT 65.445 148.795 65.785 149.425 ;
        RECT 65.955 148.795 66.205 149.595 ;
        RECT 66.395 148.945 66.725 149.425 ;
        RECT 66.895 149.135 67.120 149.595 ;
        RECT 67.290 148.945 67.620 149.425 ;
        RECT 65.445 148.745 65.675 148.795 ;
        RECT 66.395 148.775 67.620 148.945 ;
        RECT 68.250 148.815 68.750 149.425 ;
        RECT 69.170 149.135 69.920 149.425 ;
        RECT 70.430 149.135 70.760 149.595 ;
        RECT 64.465 148.355 64.815 148.605 ;
        RECT 61.305 147.215 61.645 148.185 ;
        RECT 61.815 147.045 61.985 148.185 ;
        RECT 62.175 148.015 64.610 148.185 ;
        RECT 62.255 147.045 62.505 147.845 ;
        RECT 63.150 147.215 63.480 148.015 ;
        RECT 63.780 147.045 64.110 147.845 ;
        RECT 64.280 147.215 64.610 148.015 ;
        RECT 64.985 147.045 65.275 148.210 ;
        RECT 65.445 148.185 65.620 148.745 ;
        RECT 65.790 148.435 66.485 148.605 ;
        RECT 66.315 148.185 66.485 148.435 ;
        RECT 66.660 148.405 67.080 148.605 ;
        RECT 67.250 148.405 67.580 148.605 ;
        RECT 67.750 148.405 68.080 148.605 ;
        RECT 68.250 148.185 68.420 148.815 ;
        RECT 68.605 148.355 68.955 148.605 ;
        RECT 65.445 147.215 65.785 148.185 ;
        RECT 65.955 147.045 66.125 148.185 ;
        RECT 66.315 148.015 68.750 148.185 ;
        RECT 66.395 147.045 66.645 147.845 ;
        RECT 67.290 147.215 67.620 148.015 ;
        RECT 67.920 147.045 68.250 147.845 ;
        RECT 68.420 147.215 68.750 148.015 ;
        RECT 69.170 147.845 69.540 149.135 ;
        RECT 70.980 148.945 71.250 149.155 ;
        RECT 69.915 148.775 71.250 148.945 ;
        RECT 71.510 149.025 71.685 149.425 ;
        RECT 71.855 149.215 72.185 149.595 ;
        RECT 72.430 149.095 72.660 149.425 ;
        RECT 71.510 148.855 72.140 149.025 ;
        RECT 69.915 148.605 70.085 148.775 ;
        RECT 71.970 148.685 72.140 148.855 ;
        RECT 69.710 148.355 70.085 148.605 ;
        RECT 70.255 148.365 70.730 148.605 ;
        RECT 70.900 148.365 71.250 148.605 ;
        RECT 69.915 148.185 70.085 148.355 ;
        RECT 69.915 148.015 71.250 148.185 ;
        RECT 70.970 147.855 71.250 148.015 ;
        RECT 71.425 148.005 71.790 148.685 ;
        RECT 71.970 148.355 72.320 148.685 ;
        RECT 69.170 147.675 70.340 147.845 ;
        RECT 69.625 147.045 69.840 147.505 ;
        RECT 70.010 147.215 70.340 147.675 ;
        RECT 70.510 147.045 70.760 147.845 ;
        RECT 71.970 147.835 72.140 148.355 ;
        RECT 71.510 147.665 72.140 147.835 ;
        RECT 72.490 147.805 72.660 149.095 ;
        RECT 72.860 147.985 73.140 149.260 ;
        RECT 73.365 149.255 73.635 149.260 ;
        RECT 73.325 149.085 73.635 149.255 ;
        RECT 74.095 149.215 74.425 149.595 ;
        RECT 74.595 149.340 74.930 149.385 ;
        RECT 73.365 147.985 73.635 149.085 ;
        RECT 73.825 147.985 74.165 149.015 ;
        RECT 74.595 148.875 74.935 149.340 ;
        RECT 75.195 149.045 75.365 149.335 ;
        RECT 75.535 149.215 75.865 149.595 ;
        RECT 75.195 148.875 75.860 149.045 ;
        RECT 74.335 148.355 74.595 148.685 ;
        RECT 74.335 147.805 74.505 148.355 ;
        RECT 74.765 148.185 74.935 148.875 ;
        RECT 71.510 147.215 71.685 147.665 ;
        RECT 72.490 147.635 74.505 147.805 ;
        RECT 71.855 147.045 72.185 147.485 ;
        RECT 72.490 147.215 72.660 147.635 ;
        RECT 72.895 147.045 73.565 147.455 ;
        RECT 73.780 147.215 73.950 147.635 ;
        RECT 74.150 147.045 74.480 147.455 ;
        RECT 74.675 147.215 74.935 148.185 ;
        RECT 75.110 148.055 75.460 148.705 ;
        RECT 75.630 147.885 75.860 148.875 ;
        RECT 75.195 147.715 75.860 147.885 ;
        RECT 75.195 147.215 75.365 147.715 ;
        RECT 75.535 147.045 75.865 147.545 ;
        RECT 76.035 147.215 76.220 149.335 ;
        RECT 76.475 149.135 76.725 149.595 ;
        RECT 76.895 149.145 77.230 149.315 ;
        RECT 77.425 149.145 78.100 149.315 ;
        RECT 76.895 149.005 77.065 149.145 ;
        RECT 76.390 148.015 76.670 148.965 ;
        RECT 76.840 148.875 77.065 149.005 ;
        RECT 76.840 147.770 77.010 148.875 ;
        RECT 77.235 148.725 77.760 148.945 ;
        RECT 77.180 147.960 77.420 148.555 ;
        RECT 77.590 148.025 77.760 148.725 ;
        RECT 77.930 148.365 78.100 149.145 ;
        RECT 78.420 149.095 78.790 149.595 ;
        RECT 78.970 149.145 79.375 149.315 ;
        RECT 79.545 149.145 80.330 149.315 ;
        RECT 78.970 148.915 79.140 149.145 ;
        RECT 78.310 148.615 79.140 148.915 ;
        RECT 79.525 148.645 79.990 148.975 ;
        RECT 78.310 148.585 78.510 148.615 ;
        RECT 78.630 148.365 78.800 148.435 ;
        RECT 77.930 148.195 78.800 148.365 ;
        RECT 78.290 148.105 78.800 148.195 ;
        RECT 76.840 147.640 77.145 147.770 ;
        RECT 77.590 147.660 78.120 148.025 ;
        RECT 76.460 147.045 76.725 147.505 ;
        RECT 76.895 147.215 77.145 147.640 ;
        RECT 78.290 147.490 78.460 148.105 ;
        RECT 77.355 147.320 78.460 147.490 ;
        RECT 78.630 147.045 78.800 147.845 ;
        RECT 78.970 147.545 79.140 148.615 ;
        RECT 79.310 147.715 79.500 148.435 ;
        RECT 79.670 147.685 79.990 148.645 ;
        RECT 80.160 148.685 80.330 149.145 ;
        RECT 80.605 149.065 80.815 149.595 ;
        RECT 81.075 148.855 81.405 149.380 ;
        RECT 81.575 148.985 81.745 149.595 ;
        RECT 81.915 148.940 82.245 149.375 ;
        RECT 82.465 149.050 87.810 149.595 ;
        RECT 81.915 148.855 82.295 148.940 ;
        RECT 81.205 148.685 81.405 148.855 ;
        RECT 82.070 148.815 82.295 148.855 ;
        RECT 80.160 148.355 81.035 148.685 ;
        RECT 81.205 148.355 81.955 148.685 ;
        RECT 78.970 147.215 79.220 147.545 ;
        RECT 80.160 147.515 80.330 148.355 ;
        RECT 81.205 148.150 81.395 148.355 ;
        RECT 82.125 148.235 82.295 148.815 ;
        RECT 82.080 148.185 82.295 148.235 ;
        RECT 84.050 148.220 84.390 149.050 ;
        RECT 87.985 148.825 90.575 149.595 ;
        RECT 90.745 148.845 91.955 149.595 ;
        RECT 80.500 147.775 81.395 148.150 ;
        RECT 81.905 148.105 82.295 148.185 ;
        RECT 79.445 147.345 80.330 147.515 ;
        RECT 80.510 147.045 80.825 147.545 ;
        RECT 81.055 147.215 81.395 147.775 ;
        RECT 81.565 147.045 81.735 148.055 ;
        RECT 81.905 147.260 82.235 148.105 ;
        RECT 85.870 147.480 86.220 148.730 ;
        RECT 87.985 148.305 89.195 148.825 ;
        RECT 89.365 148.135 90.575 148.655 ;
        RECT 82.465 147.045 87.810 147.480 ;
        RECT 87.985 147.045 90.575 148.135 ;
        RECT 90.745 148.135 91.265 148.675 ;
        RECT 91.435 148.305 91.955 148.845 ;
        RECT 101.840 148.320 102.010 149.730 ;
        RECT 102.380 149.160 105.420 149.330 ;
        RECT 102.380 148.720 105.420 148.890 ;
        RECT 105.635 148.860 105.805 149.190 ;
        RECT 106.140 148.970 118.590 149.730 ;
        RECT 121.720 149.730 138.470 149.900 ;
        RECT 146.140 149.850 158.550 149.900 ;
        RECT 106.140 148.960 118.480 148.970 ;
        RECT 106.140 148.950 112.020 148.960 ;
        RECT 106.140 148.930 106.710 148.950 ;
        RECT 107.930 148.940 112.020 148.950 ;
        RECT 106.150 148.320 106.320 148.930 ;
        RECT 101.840 148.150 106.320 148.320 ;
        RECT 121.720 148.320 121.890 149.730 ;
        RECT 122.260 149.160 125.300 149.330 ;
        RECT 122.260 148.720 125.300 148.890 ;
        RECT 125.515 148.860 125.685 149.190 ;
        RECT 126.020 148.970 138.470 149.730 ;
        RECT 141.800 149.680 158.550 149.850 ;
        RECT 126.020 148.960 138.360 148.970 ;
        RECT 126.020 148.950 131.900 148.960 ;
        RECT 126.020 148.930 126.590 148.950 ;
        RECT 127.810 148.940 131.900 148.950 ;
        RECT 126.030 148.320 126.200 148.930 ;
        RECT 121.720 148.150 126.200 148.320 ;
        RECT 141.800 148.270 141.970 149.680 ;
        RECT 142.340 149.110 145.380 149.280 ;
        RECT 142.340 148.670 145.380 148.840 ;
        RECT 145.595 148.810 145.765 149.140 ;
        RECT 146.100 148.920 158.550 149.680 ;
        RECT 146.100 148.910 158.440 148.920 ;
        RECT 146.100 148.900 151.980 148.910 ;
        RECT 146.100 148.880 146.670 148.900 ;
        RECT 147.890 148.890 151.980 148.900 ;
        RECT 146.110 148.270 146.280 148.880 ;
        RECT 90.745 147.045 91.955 148.135 ;
        RECT 141.800 148.100 146.280 148.270 ;
        RECT 13.380 146.875 92.040 147.045 ;
        RECT 13.465 145.785 14.675 146.875 ;
        RECT 14.845 146.440 20.190 146.875 ;
        RECT 20.365 146.440 25.710 146.875 ;
        RECT 13.465 145.075 13.985 145.615 ;
        RECT 14.155 145.245 14.675 145.785 ;
        RECT 13.465 144.325 14.675 145.075 ;
        RECT 16.430 144.870 16.770 145.700 ;
        RECT 18.250 145.190 18.600 146.440 ;
        RECT 21.950 144.870 22.290 145.700 ;
        RECT 23.770 145.190 24.120 146.440 ;
        RECT 26.345 145.710 26.635 146.875 ;
        RECT 26.805 145.785 28.015 146.875 ;
        RECT 26.805 145.075 27.325 145.615 ;
        RECT 27.495 145.245 28.015 145.785 ;
        RECT 28.185 145.735 28.465 146.875 ;
        RECT 28.635 145.725 28.965 146.705 ;
        RECT 29.135 145.735 29.395 146.875 ;
        RECT 28.195 145.295 28.530 145.565 ;
        RECT 28.700 145.125 28.870 145.725 ;
        RECT 29.040 145.315 29.375 145.565 ;
        RECT 14.845 144.325 20.190 144.870 ;
        RECT 20.365 144.325 25.710 144.870 ;
        RECT 26.345 144.325 26.635 145.050 ;
        RECT 26.805 144.325 28.015 145.075 ;
        RECT 28.185 144.325 28.495 145.125 ;
        RECT 28.700 144.495 29.395 145.125 ;
        RECT 30.495 144.505 30.755 146.695 ;
        RECT 30.925 146.145 31.265 146.875 ;
        RECT 31.445 145.965 31.715 146.695 ;
        RECT 30.945 145.745 31.715 145.965 ;
        RECT 31.895 145.985 32.125 146.695 ;
        RECT 32.295 146.165 32.625 146.875 ;
        RECT 32.795 145.985 33.055 146.695 ;
        RECT 33.360 146.245 33.645 146.705 ;
        RECT 33.815 146.415 34.085 146.875 ;
        RECT 33.360 146.025 34.315 146.245 ;
        RECT 31.895 145.745 33.055 145.985 ;
        RECT 30.945 145.075 31.235 145.745 ;
        RECT 31.415 145.255 31.880 145.565 ;
        RECT 32.060 145.255 32.585 145.565 ;
        RECT 30.945 144.875 32.175 145.075 ;
        RECT 31.015 144.325 31.685 144.695 ;
        RECT 31.865 144.505 32.175 144.875 ;
        RECT 32.355 144.615 32.585 145.255 ;
        RECT 32.765 145.235 33.065 145.565 ;
        RECT 33.245 145.295 33.935 145.855 ;
        RECT 34.105 145.125 34.315 146.025 ;
        RECT 32.765 144.325 33.055 145.055 ;
        RECT 33.360 144.955 34.315 145.125 ;
        RECT 34.485 145.855 34.885 146.705 ;
        RECT 35.075 146.245 35.355 146.705 ;
        RECT 35.875 146.415 36.200 146.875 ;
        RECT 35.075 146.025 36.200 146.245 ;
        RECT 34.485 145.295 35.580 145.855 ;
        RECT 35.750 145.565 36.200 146.025 ;
        RECT 36.370 145.735 36.755 146.705 ;
        RECT 37.110 145.905 37.500 146.080 ;
        RECT 37.985 146.075 38.315 146.875 ;
        RECT 38.485 146.085 39.020 146.705 ;
        RECT 37.110 145.735 38.535 145.905 ;
        RECT 33.360 144.495 33.645 144.955 ;
        RECT 33.815 144.325 34.085 144.785 ;
        RECT 34.485 144.495 34.885 145.295 ;
        RECT 35.750 145.235 36.305 145.565 ;
        RECT 35.750 145.125 36.200 145.235 ;
        RECT 35.075 144.955 36.200 145.125 ;
        RECT 36.475 145.065 36.755 145.735 ;
        RECT 35.075 144.495 35.355 144.955 ;
        RECT 35.875 144.325 36.200 144.785 ;
        RECT 36.370 144.495 36.755 145.065 ;
        RECT 36.985 145.005 37.340 145.565 ;
        RECT 37.510 144.835 37.680 145.735 ;
        RECT 37.850 145.005 38.115 145.565 ;
        RECT 38.365 145.235 38.535 145.735 ;
        RECT 38.705 145.065 39.020 146.085 ;
        RECT 39.265 145.735 39.495 146.875 ;
        RECT 39.665 145.725 39.995 146.705 ;
        RECT 40.165 145.735 40.375 146.875 ;
        RECT 40.690 146.255 40.865 146.705 ;
        RECT 41.035 146.435 41.365 146.875 ;
        RECT 41.670 146.285 41.840 146.705 ;
        RECT 42.075 146.465 42.745 146.875 ;
        RECT 42.960 146.285 43.130 146.705 ;
        RECT 43.330 146.465 43.660 146.875 ;
        RECT 40.690 146.085 41.320 146.255 ;
        RECT 39.245 145.315 39.575 145.565 ;
        RECT 37.090 144.325 37.330 144.835 ;
        RECT 37.510 144.505 37.790 144.835 ;
        RECT 38.020 144.325 38.235 144.835 ;
        RECT 38.405 144.495 39.020 145.065 ;
        RECT 39.265 144.325 39.495 145.145 ;
        RECT 39.745 145.125 39.995 145.725 ;
        RECT 40.605 145.235 40.970 145.915 ;
        RECT 41.150 145.565 41.320 146.085 ;
        RECT 41.670 146.115 43.685 146.285 ;
        RECT 41.150 145.235 41.500 145.565 ;
        RECT 39.665 144.495 39.995 145.125 ;
        RECT 40.165 144.325 40.375 145.145 ;
        RECT 41.150 145.065 41.320 145.235 ;
        RECT 40.690 144.895 41.320 145.065 ;
        RECT 40.690 144.495 40.865 144.895 ;
        RECT 41.670 144.825 41.840 146.115 ;
        RECT 41.035 144.325 41.365 144.705 ;
        RECT 41.610 144.495 41.840 144.825 ;
        RECT 42.040 144.660 42.320 145.935 ;
        RECT 42.545 145.855 42.815 145.935 ;
        RECT 42.505 145.685 42.815 145.855 ;
        RECT 42.545 144.660 42.815 145.685 ;
        RECT 43.005 144.905 43.345 145.935 ;
        RECT 43.515 145.565 43.685 146.115 ;
        RECT 43.855 145.735 44.115 146.705 ;
        RECT 44.285 146.440 49.630 146.875 ;
        RECT 43.515 145.235 43.775 145.565 ;
        RECT 43.945 145.045 44.115 145.735 ;
        RECT 43.275 144.325 43.605 144.705 ;
        RECT 43.775 144.580 44.115 145.045 ;
        RECT 45.870 144.870 46.210 145.700 ;
        RECT 47.690 145.190 48.040 146.440 ;
        RECT 49.805 145.785 51.475 146.875 ;
        RECT 49.805 145.095 50.555 145.615 ;
        RECT 50.725 145.265 51.475 145.785 ;
        RECT 52.105 145.710 52.395 146.875 ;
        RECT 52.565 146.440 57.910 146.875 ;
        RECT 43.775 144.535 44.110 144.580 ;
        RECT 44.285 144.325 49.630 144.870 ;
        RECT 49.805 144.325 51.475 145.095 ;
        RECT 52.105 144.325 52.395 145.050 ;
        RECT 54.150 144.870 54.490 145.700 ;
        RECT 55.970 145.190 56.320 146.440 ;
        RECT 58.745 146.205 59.025 146.875 ;
        RECT 59.195 145.985 59.495 146.535 ;
        RECT 59.695 146.155 60.025 146.875 ;
        RECT 60.215 146.155 60.675 146.705 ;
        RECT 58.560 145.565 58.825 145.925 ;
        RECT 59.195 145.815 60.135 145.985 ;
        RECT 59.965 145.565 60.135 145.815 ;
        RECT 58.560 145.315 59.235 145.565 ;
        RECT 59.455 145.315 59.795 145.565 ;
        RECT 59.965 145.235 60.255 145.565 ;
        RECT 59.965 145.145 60.135 145.235 ;
        RECT 58.745 144.955 60.135 145.145 ;
        RECT 52.565 144.325 57.910 144.870 ;
        RECT 58.745 144.595 59.075 144.955 ;
        RECT 60.425 144.785 60.675 146.155 ;
        RECT 60.845 145.735 61.105 146.875 ;
        RECT 61.345 146.365 62.960 146.695 ;
        RECT 61.355 145.565 61.525 146.125 ;
        RECT 61.785 146.025 62.960 146.195 ;
        RECT 63.130 146.075 63.410 146.875 ;
        RECT 61.785 145.735 62.115 146.025 ;
        RECT 62.790 145.905 62.960 146.025 ;
        RECT 62.285 145.565 62.530 145.855 ;
        RECT 62.790 145.735 63.450 145.905 ;
        RECT 63.620 145.735 63.895 146.705 ;
        RECT 64.165 146.415 64.335 146.875 ;
        RECT 64.505 145.925 64.835 146.705 ;
        RECT 65.005 146.075 65.175 146.875 ;
        RECT 63.280 145.565 63.450 145.735 ;
        RECT 60.850 145.315 61.185 145.565 ;
        RECT 61.355 145.235 62.070 145.565 ;
        RECT 62.285 145.235 63.110 145.565 ;
        RECT 63.280 145.235 63.555 145.565 ;
        RECT 61.355 145.145 61.605 145.235 ;
        RECT 59.695 144.325 59.945 144.785 ;
        RECT 60.115 144.495 60.675 144.785 ;
        RECT 60.845 144.325 61.105 145.145 ;
        RECT 61.275 144.725 61.605 145.145 ;
        RECT 63.280 145.065 63.450 145.235 ;
        RECT 61.785 144.895 63.450 145.065 ;
        RECT 63.725 145.000 63.895 145.735 ;
        RECT 61.785 144.495 62.045 144.895 ;
        RECT 62.215 144.325 62.545 144.725 ;
        RECT 62.715 144.545 62.885 144.895 ;
        RECT 63.055 144.325 63.430 144.725 ;
        RECT 63.620 144.655 63.895 145.000 ;
        RECT 64.065 145.905 64.835 145.925 ;
        RECT 65.345 145.905 65.675 146.705 ;
        RECT 65.845 146.075 66.015 146.875 ;
        RECT 66.185 145.905 66.515 146.705 ;
        RECT 64.065 145.735 66.515 145.905 ;
        RECT 66.775 145.735 67.070 146.875 ;
        RECT 67.295 145.765 67.590 146.875 ;
        RECT 64.065 145.145 64.415 145.735 ;
        RECT 67.770 145.565 68.020 146.700 ;
        RECT 68.190 145.765 68.450 146.875 ;
        RECT 68.620 145.975 68.880 146.700 ;
        RECT 69.050 146.145 69.310 146.875 ;
        RECT 69.480 145.975 69.740 146.700 ;
        RECT 69.910 146.145 70.170 146.875 ;
        RECT 70.340 145.975 70.600 146.700 ;
        RECT 70.770 146.145 71.030 146.875 ;
        RECT 71.200 145.975 71.460 146.700 ;
        RECT 71.630 146.145 71.925 146.875 ;
        RECT 68.620 145.735 71.930 145.975 ;
        RECT 64.585 145.315 67.095 145.565 ;
        RECT 64.065 144.965 66.435 145.145 ;
        RECT 64.165 144.325 64.415 144.790 ;
        RECT 64.585 144.495 64.755 144.965 ;
        RECT 65.005 144.325 65.175 144.785 ;
        RECT 65.425 144.495 65.595 144.965 ;
        RECT 65.845 144.325 66.015 144.785 ;
        RECT 66.265 144.495 66.435 144.965 ;
        RECT 67.285 144.955 67.600 145.565 ;
        RECT 67.770 145.315 70.790 145.565 ;
        RECT 66.805 144.325 67.070 144.785 ;
        RECT 67.345 144.325 67.590 144.785 ;
        RECT 67.770 144.505 68.020 145.315 ;
        RECT 70.960 145.145 71.930 145.735 ;
        RECT 68.620 144.975 71.930 145.145 ;
        RECT 68.190 144.325 68.450 144.850 ;
        RECT 68.620 144.520 68.880 144.975 ;
        RECT 69.050 144.325 69.310 144.805 ;
        RECT 69.480 144.520 69.740 144.975 ;
        RECT 69.910 144.325 70.170 144.805 ;
        RECT 70.340 144.520 70.600 144.975 ;
        RECT 70.770 144.325 71.030 144.805 ;
        RECT 71.200 144.520 71.460 144.975 ;
        RECT 71.630 144.325 71.930 144.805 ;
        RECT 72.345 144.495 72.605 146.705 ;
        RECT 72.775 146.495 73.105 146.875 ;
        RECT 73.530 146.325 73.700 146.705 ;
        RECT 73.960 146.495 74.290 146.875 ;
        RECT 74.485 146.325 74.655 146.705 ;
        RECT 74.865 146.495 75.195 146.875 ;
        RECT 75.445 146.325 75.635 146.705 ;
        RECT 75.875 146.495 76.205 146.875 ;
        RECT 76.515 146.375 76.775 146.705 ;
        RECT 72.775 146.155 74.725 146.325 ;
        RECT 72.775 145.235 72.945 146.155 ;
        RECT 73.315 145.565 73.510 145.875 ;
        RECT 73.780 145.565 73.965 145.875 ;
        RECT 73.255 145.235 73.510 145.565 ;
        RECT 73.735 145.235 73.965 145.565 ;
        RECT 72.775 144.325 73.105 144.705 ;
        RECT 73.315 144.660 73.510 145.235 ;
        RECT 73.780 144.655 73.965 145.235 ;
        RECT 74.215 144.665 74.385 145.565 ;
        RECT 74.555 145.165 74.725 146.155 ;
        RECT 74.895 146.155 75.635 146.325 ;
        RECT 74.895 145.645 75.065 146.155 ;
        RECT 75.235 145.815 75.815 145.985 ;
        RECT 76.085 145.865 76.435 146.195 ;
        RECT 75.645 145.695 75.815 145.815 ;
        RECT 76.605 145.695 76.775 146.375 ;
        RECT 77.865 145.710 78.155 146.875 ;
        RECT 78.325 145.800 78.595 146.705 ;
        RECT 78.765 146.115 79.095 146.875 ;
        RECT 79.275 145.945 79.445 146.705 ;
        RECT 79.705 146.440 85.050 146.875 ;
        RECT 85.225 146.440 90.570 146.875 ;
        RECT 74.895 145.475 75.465 145.645 ;
        RECT 75.645 145.525 76.775 145.695 ;
        RECT 74.555 144.835 75.105 145.165 ;
        RECT 75.295 144.995 75.465 145.475 ;
        RECT 75.635 145.185 76.255 145.355 ;
        RECT 76.045 145.005 76.255 145.185 ;
        RECT 75.295 144.665 75.695 144.995 ;
        RECT 76.605 144.825 76.775 145.525 ;
        RECT 74.215 144.495 75.695 144.665 ;
        RECT 75.875 144.325 76.205 144.705 ;
        RECT 76.515 144.495 76.775 144.825 ;
        RECT 77.865 144.325 78.155 145.050 ;
        RECT 78.325 145.000 78.495 145.800 ;
        RECT 78.780 145.775 79.445 145.945 ;
        RECT 78.780 145.630 78.950 145.775 ;
        RECT 78.665 145.300 78.950 145.630 ;
        RECT 78.780 145.045 78.950 145.300 ;
        RECT 79.185 145.225 79.515 145.595 ;
        RECT 78.325 144.495 78.585 145.000 ;
        RECT 78.780 144.875 79.445 145.045 ;
        RECT 78.765 144.325 79.095 144.705 ;
        RECT 79.275 144.495 79.445 144.875 ;
        RECT 81.290 144.870 81.630 145.700 ;
        RECT 83.110 145.190 83.460 146.440 ;
        RECT 86.810 144.870 87.150 145.700 ;
        RECT 88.630 145.190 88.980 146.440 ;
        RECT 90.745 145.785 91.955 146.875 ;
        RECT 100.630 146.740 106.370 146.750 ;
        RECT 100.140 146.580 106.370 146.740 ;
        RECT 90.745 145.245 91.265 145.785 ;
        RECT 91.435 145.075 91.955 145.615 ;
        RECT 79.705 144.325 85.050 144.870 ;
        RECT 85.225 144.325 90.570 144.870 ;
        RECT 90.745 144.325 91.955 145.075 ;
        RECT 13.380 144.155 92.040 144.325 ;
        RECT 100.140 144.320 100.810 146.580 ;
        RECT 101.480 146.010 105.520 146.180 ;
        RECT 101.140 144.950 101.310 145.950 ;
        RECT 105.690 144.950 105.860 145.950 ;
        RECT 101.480 144.720 105.520 144.890 ;
        RECT 106.200 144.320 106.370 146.580 ;
        RECT 13.465 143.405 14.675 144.155 ;
        RECT 14.845 143.610 20.190 144.155 ;
        RECT 13.465 142.865 13.985 143.405 ;
        RECT 14.155 142.695 14.675 143.235 ;
        RECT 16.430 142.780 16.770 143.610 ;
        RECT 20.365 143.385 22.955 144.155 ;
        RECT 23.125 143.695 23.685 143.985 ;
        RECT 23.855 143.695 24.105 144.155 ;
        RECT 13.465 141.605 14.675 142.695 ;
        RECT 18.250 142.040 18.600 143.290 ;
        RECT 20.365 142.865 21.575 143.385 ;
        RECT 21.745 142.695 22.955 143.215 ;
        RECT 14.845 141.605 20.190 142.040 ;
        RECT 20.365 141.605 22.955 142.695 ;
        RECT 23.125 142.325 23.375 143.695 ;
        RECT 24.725 143.525 25.055 143.885 ;
        RECT 25.590 143.645 25.830 144.155 ;
        RECT 26.010 143.645 26.290 143.975 ;
        RECT 26.520 143.645 26.735 144.155 ;
        RECT 23.665 143.335 25.055 143.525 ;
        RECT 23.665 143.245 23.835 143.335 ;
        RECT 23.545 142.915 23.835 143.245 ;
        RECT 24.005 142.915 24.345 143.165 ;
        RECT 24.565 142.915 25.240 143.165 ;
        RECT 25.485 142.915 25.840 143.475 ;
        RECT 23.665 142.665 23.835 142.915 ;
        RECT 23.665 142.495 24.605 142.665 ;
        RECT 24.975 142.555 25.240 142.915 ;
        RECT 26.010 142.745 26.180 143.645 ;
        RECT 26.350 142.915 26.615 143.475 ;
        RECT 26.905 143.415 27.520 143.985 ;
        RECT 27.725 143.655 28.065 144.155 ;
        RECT 26.865 142.745 27.035 143.245 ;
        RECT 25.610 142.575 27.035 142.745 ;
        RECT 23.125 141.775 23.585 142.325 ;
        RECT 23.775 141.605 24.105 142.325 ;
        RECT 24.305 141.945 24.605 142.495 ;
        RECT 25.610 142.400 26.000 142.575 ;
        RECT 24.775 141.605 25.055 142.275 ;
        RECT 26.485 141.605 26.815 142.405 ;
        RECT 27.205 142.395 27.520 143.415 ;
        RECT 27.725 142.915 28.065 143.485 ;
        RECT 28.235 143.245 28.480 143.935 ;
        RECT 28.675 143.655 29.005 144.155 ;
        RECT 29.205 143.585 29.375 143.935 ;
        RECT 29.550 143.755 29.880 144.155 ;
        RECT 30.050 143.585 30.220 143.935 ;
        RECT 30.390 143.755 30.770 144.155 ;
        RECT 29.205 143.415 30.790 143.585 ;
        RECT 30.960 143.480 31.235 143.825 ;
        RECT 31.465 143.695 31.710 144.155 ;
        RECT 30.620 143.245 30.790 143.415 ;
        RECT 28.235 142.915 28.890 143.245 ;
        RECT 26.985 141.775 27.520 142.395 ;
        RECT 27.725 141.605 28.065 142.680 ;
        RECT 28.235 142.320 28.475 142.915 ;
        RECT 28.670 142.455 28.990 142.745 ;
        RECT 29.160 142.625 29.900 143.245 ;
        RECT 30.070 142.915 30.450 143.245 ;
        RECT 30.620 142.915 30.895 143.245 ;
        RECT 30.620 142.745 30.790 142.915 ;
        RECT 31.065 142.745 31.235 143.480 ;
        RECT 31.405 142.915 31.720 143.525 ;
        RECT 31.890 143.165 32.140 143.975 ;
        RECT 32.310 143.630 32.570 144.155 ;
        RECT 32.740 143.505 33.000 143.960 ;
        RECT 33.170 143.675 33.430 144.155 ;
        RECT 33.600 143.505 33.860 143.960 ;
        RECT 34.030 143.675 34.290 144.155 ;
        RECT 34.460 143.505 34.720 143.960 ;
        RECT 34.890 143.675 35.150 144.155 ;
        RECT 35.320 143.505 35.580 143.960 ;
        RECT 35.750 143.675 36.050 144.155 ;
        RECT 36.745 143.525 37.125 143.975 ;
        RECT 32.740 143.335 36.050 143.505 ;
        RECT 31.890 142.915 34.910 143.165 ;
        RECT 30.130 142.575 30.790 142.745 ;
        RECT 30.130 142.455 30.300 142.575 ;
        RECT 28.670 142.285 30.300 142.455 ;
        RECT 28.245 141.945 30.300 142.115 ;
        RECT 28.250 141.825 30.300 141.945 ;
        RECT 30.470 141.605 30.750 142.405 ;
        RECT 30.960 141.775 31.235 142.745 ;
        RECT 31.415 141.605 31.710 142.715 ;
        RECT 31.890 141.780 32.140 142.915 ;
        RECT 35.080 142.745 36.050 143.335 ;
        RECT 32.310 141.605 32.570 142.715 ;
        RECT 32.740 142.505 36.050 142.745 ;
        RECT 36.485 142.575 36.715 143.265 ;
        RECT 36.895 143.075 37.125 143.525 ;
        RECT 37.305 143.375 37.535 144.155 ;
        RECT 37.715 143.445 38.145 143.975 ;
        RECT 37.715 143.195 37.960 143.445 ;
        RECT 38.325 143.245 38.535 143.865 ;
        RECT 38.705 143.425 39.035 144.155 ;
        RECT 39.225 143.430 39.515 144.155 ;
        RECT 39.695 143.665 40.025 144.155 ;
        RECT 40.195 143.560 40.815 143.985 ;
        RECT 32.740 141.780 33.000 142.505 ;
        RECT 33.170 141.605 33.430 142.335 ;
        RECT 33.600 141.780 33.860 142.505 ;
        RECT 34.030 141.605 34.290 142.335 ;
        RECT 34.460 141.780 34.720 142.505 ;
        RECT 34.890 141.605 35.150 142.335 ;
        RECT 35.320 141.780 35.580 142.505 ;
        RECT 36.895 142.395 37.235 143.075 ;
        RECT 35.750 141.605 36.045 142.335 ;
        RECT 36.475 142.195 37.235 142.395 ;
        RECT 37.425 142.895 37.960 143.195 ;
        RECT 38.140 142.895 38.535 143.245 ;
        RECT 38.730 142.895 39.020 143.245 ;
        RECT 39.685 142.915 40.025 143.495 ;
        RECT 40.195 143.225 40.555 143.560 ;
        RECT 41.275 143.465 41.605 144.155 ;
        RECT 42.445 143.480 42.705 143.985 ;
        RECT 42.885 143.775 43.215 144.155 ;
        RECT 43.395 143.605 43.565 143.985 ;
        RECT 40.195 142.945 41.615 143.225 ;
        RECT 36.475 141.805 36.735 142.195 ;
        RECT 36.905 141.605 37.235 142.015 ;
        RECT 37.425 141.785 37.755 142.895 ;
        RECT 37.925 142.515 38.965 142.715 ;
        RECT 37.925 141.785 38.115 142.515 ;
        RECT 38.285 141.605 38.615 142.335 ;
        RECT 38.795 141.785 38.965 142.515 ;
        RECT 39.225 141.605 39.515 142.770 ;
        RECT 39.695 141.605 40.025 142.745 ;
        RECT 40.195 141.775 40.555 142.945 ;
        RECT 40.755 141.605 41.085 142.775 ;
        RECT 41.285 141.775 41.615 142.945 ;
        RECT 41.815 141.605 42.145 142.775 ;
        RECT 42.445 142.680 42.615 143.480 ;
        RECT 42.900 143.435 43.565 143.605 ;
        RECT 42.900 143.180 43.070 143.435 ;
        RECT 44.755 143.345 45.025 144.155 ;
        RECT 45.195 143.345 45.525 143.985 ;
        RECT 45.695 143.345 45.935 144.155 ;
        RECT 46.125 143.385 47.795 144.155 ;
        RECT 42.785 142.850 43.070 143.180 ;
        RECT 43.305 142.885 43.635 143.255 ;
        RECT 44.745 142.915 45.095 143.165 ;
        RECT 42.900 142.705 43.070 142.850 ;
        RECT 45.265 142.745 45.435 143.345 ;
        RECT 45.605 142.915 45.955 143.165 ;
        RECT 46.125 142.865 46.875 143.385 ;
        RECT 48.435 143.345 48.705 144.155 ;
        RECT 48.875 143.345 49.205 143.985 ;
        RECT 49.375 143.345 49.615 144.155 ;
        RECT 49.810 143.755 50.145 144.155 ;
        RECT 50.315 143.585 50.520 143.985 ;
        RECT 50.730 143.675 51.005 144.155 ;
        RECT 51.215 143.655 51.475 143.985 ;
        RECT 49.835 143.415 50.520 143.585 ;
        RECT 42.445 141.775 42.715 142.680 ;
        RECT 42.900 142.535 43.565 142.705 ;
        RECT 42.885 141.605 43.215 142.365 ;
        RECT 43.395 141.775 43.565 142.535 ;
        RECT 44.755 141.605 45.085 142.745 ;
        RECT 45.265 142.575 45.945 142.745 ;
        RECT 47.045 142.695 47.795 143.215 ;
        RECT 48.425 142.915 48.775 143.165 ;
        RECT 48.945 142.745 49.115 143.345 ;
        RECT 49.285 142.915 49.635 143.165 ;
        RECT 45.615 141.790 45.945 142.575 ;
        RECT 46.125 141.605 47.795 142.695 ;
        RECT 48.435 141.605 48.765 142.745 ;
        RECT 48.945 142.575 49.625 142.745 ;
        RECT 49.295 141.790 49.625 142.575 ;
        RECT 49.835 142.385 50.175 143.415 ;
        RECT 50.345 142.745 50.595 143.245 ;
        RECT 50.775 142.915 51.135 143.495 ;
        RECT 51.305 142.745 51.475 143.655 ;
        RECT 51.695 143.500 52.025 143.935 ;
        RECT 52.195 143.545 52.365 144.155 ;
        RECT 50.345 142.575 51.475 142.745 ;
        RECT 51.645 143.415 52.025 143.500 ;
        RECT 52.535 143.415 52.865 143.940 ;
        RECT 53.125 143.625 53.335 144.155 ;
        RECT 53.610 143.705 54.395 143.875 ;
        RECT 54.565 143.705 54.970 143.875 ;
        RECT 51.645 143.375 51.870 143.415 ;
        RECT 51.645 142.795 51.815 143.375 ;
        RECT 52.535 143.245 52.735 143.415 ;
        RECT 53.610 143.245 53.780 143.705 ;
        RECT 51.985 142.915 52.735 143.245 ;
        RECT 52.905 142.915 53.780 143.245 ;
        RECT 51.645 142.745 51.860 142.795 ;
        RECT 51.645 142.665 52.035 142.745 ;
        RECT 49.835 142.210 50.500 142.385 ;
        RECT 49.810 141.605 50.145 142.030 ;
        RECT 50.315 141.805 50.500 142.210 ;
        RECT 50.705 141.605 51.035 142.385 ;
        RECT 51.205 141.805 51.475 142.575 ;
        RECT 51.705 141.820 52.035 142.665 ;
        RECT 52.545 142.710 52.735 142.915 ;
        RECT 52.205 141.605 52.375 142.615 ;
        RECT 52.545 142.335 53.440 142.710 ;
        RECT 52.545 141.775 52.885 142.335 ;
        RECT 53.115 141.605 53.430 142.105 ;
        RECT 53.610 142.075 53.780 142.915 ;
        RECT 53.950 143.205 54.415 143.535 ;
        RECT 54.800 143.475 54.970 143.705 ;
        RECT 55.150 143.655 55.520 144.155 ;
        RECT 55.840 143.705 56.515 143.875 ;
        RECT 56.710 143.705 57.045 143.875 ;
        RECT 53.950 142.245 54.270 143.205 ;
        RECT 54.800 143.175 55.630 143.475 ;
        RECT 54.440 142.275 54.630 142.995 ;
        RECT 54.800 142.105 54.970 143.175 ;
        RECT 55.430 143.145 55.630 143.175 ;
        RECT 55.140 142.925 55.310 142.995 ;
        RECT 55.840 142.925 56.010 143.705 ;
        RECT 56.875 143.565 57.045 143.705 ;
        RECT 57.215 143.695 57.465 144.155 ;
        RECT 55.140 142.755 56.010 142.925 ;
        RECT 56.180 143.285 56.705 143.505 ;
        RECT 56.875 143.435 57.100 143.565 ;
        RECT 55.140 142.665 55.650 142.755 ;
        RECT 53.610 141.905 54.495 142.075 ;
        RECT 54.720 141.775 54.970 142.105 ;
        RECT 55.140 141.605 55.310 142.405 ;
        RECT 55.480 142.050 55.650 142.665 ;
        RECT 56.180 142.585 56.350 143.285 ;
        RECT 55.820 142.220 56.350 142.585 ;
        RECT 56.520 142.520 56.760 143.115 ;
        RECT 56.930 142.330 57.100 143.435 ;
        RECT 57.270 142.575 57.550 143.525 ;
        RECT 56.795 142.200 57.100 142.330 ;
        RECT 55.480 141.880 56.585 142.050 ;
        RECT 56.795 141.775 57.045 142.200 ;
        RECT 57.215 141.605 57.480 142.065 ;
        RECT 57.720 141.775 57.905 143.895 ;
        RECT 58.075 143.775 58.405 144.155 ;
        RECT 58.575 143.605 58.745 143.895 ;
        RECT 58.080 143.435 58.745 143.605 ;
        RECT 58.080 142.445 58.310 143.435 ;
        RECT 58.480 142.615 58.830 143.265 ;
        RECT 58.080 142.275 58.745 142.445 ;
        RECT 58.075 141.605 58.405 142.105 ;
        RECT 58.575 141.775 58.745 142.275 ;
        RECT 59.925 141.775 60.205 143.875 ;
        RECT 60.435 143.695 60.605 144.155 ;
        RECT 60.875 143.765 62.125 143.945 ;
        RECT 61.260 143.525 61.625 143.595 ;
        RECT 60.375 143.345 61.625 143.525 ;
        RECT 61.795 143.545 62.125 143.765 ;
        RECT 62.295 143.715 62.465 144.155 ;
        RECT 62.635 143.545 62.975 143.960 ;
        RECT 61.795 143.375 62.975 143.545 ;
        RECT 63.145 143.385 64.815 144.155 ;
        RECT 64.985 143.430 65.275 144.155 ;
        RECT 60.375 142.745 60.650 143.345 ;
        RECT 60.820 142.915 61.175 143.165 ;
        RECT 61.370 143.135 61.835 143.165 ;
        RECT 61.365 142.965 61.835 143.135 ;
        RECT 61.370 142.915 61.835 142.965 ;
        RECT 62.005 142.915 62.335 143.165 ;
        RECT 62.510 142.965 62.975 143.165 ;
        RECT 62.155 142.795 62.335 142.915 ;
        RECT 63.145 142.865 63.895 143.385 ;
        RECT 60.375 142.535 61.985 142.745 ;
        RECT 62.155 142.625 62.485 142.795 ;
        RECT 61.575 142.435 61.985 142.535 ;
        RECT 60.395 141.605 61.180 142.365 ;
        RECT 61.575 141.775 61.960 142.435 ;
        RECT 62.285 141.835 62.485 142.625 ;
        RECT 62.655 141.605 62.975 142.785 ;
        RECT 64.065 142.695 64.815 143.215 ;
        RECT 65.445 143.210 65.785 143.985 ;
        RECT 65.955 143.695 66.125 144.155 ;
        RECT 66.365 143.720 66.725 143.985 ;
        RECT 66.365 143.715 66.720 143.720 ;
        RECT 66.365 143.705 66.715 143.715 ;
        RECT 66.365 143.700 66.710 143.705 ;
        RECT 66.365 143.690 66.705 143.700 ;
        RECT 67.355 143.695 67.525 144.155 ;
        RECT 66.365 143.685 66.700 143.690 ;
        RECT 66.365 143.675 66.690 143.685 ;
        RECT 66.365 143.665 66.680 143.675 ;
        RECT 66.365 143.525 66.665 143.665 ;
        RECT 65.955 143.335 66.665 143.525 ;
        RECT 66.855 143.525 67.185 143.605 ;
        RECT 67.695 143.525 68.035 143.985 ;
        RECT 66.855 143.335 68.035 143.525 ;
        RECT 68.205 143.385 69.875 144.155 ;
        RECT 70.135 143.605 70.305 143.895 ;
        RECT 70.475 143.775 70.805 144.155 ;
        RECT 70.135 143.435 70.800 143.605 ;
        RECT 63.145 141.605 64.815 142.695 ;
        RECT 64.985 141.605 65.275 142.770 ;
        RECT 65.445 141.775 65.725 143.210 ;
        RECT 65.955 142.765 66.240 143.335 ;
        RECT 66.425 142.935 66.895 143.165 ;
        RECT 67.065 143.145 67.395 143.165 ;
        RECT 67.065 142.965 67.515 143.145 ;
        RECT 67.705 142.965 68.035 143.165 ;
        RECT 65.955 142.550 67.105 142.765 ;
        RECT 65.895 141.605 66.605 142.380 ;
        RECT 66.775 141.775 67.105 142.550 ;
        RECT 67.300 141.850 67.515 142.965 ;
        RECT 67.805 142.625 68.035 142.965 ;
        RECT 68.205 142.865 68.955 143.385 ;
        RECT 69.125 142.695 69.875 143.215 ;
        RECT 67.695 141.605 68.025 142.325 ;
        RECT 68.205 141.605 69.875 142.695 ;
        RECT 70.050 142.615 70.400 143.265 ;
        RECT 70.570 142.445 70.800 143.435 ;
        RECT 70.135 142.275 70.800 142.445 ;
        RECT 70.135 141.775 70.305 142.275 ;
        RECT 70.475 141.605 70.805 142.105 ;
        RECT 70.975 141.775 71.160 143.895 ;
        RECT 71.415 143.695 71.665 144.155 ;
        RECT 71.835 143.705 72.170 143.875 ;
        RECT 72.365 143.705 73.040 143.875 ;
        RECT 71.835 143.565 72.005 143.705 ;
        RECT 71.330 142.575 71.610 143.525 ;
        RECT 71.780 143.435 72.005 143.565 ;
        RECT 71.780 142.330 71.950 143.435 ;
        RECT 72.175 143.285 72.700 143.505 ;
        RECT 72.120 142.520 72.360 143.115 ;
        RECT 72.530 142.585 72.700 143.285 ;
        RECT 72.870 142.925 73.040 143.705 ;
        RECT 73.360 143.655 73.730 144.155 ;
        RECT 73.910 143.705 74.315 143.875 ;
        RECT 74.485 143.705 75.270 143.875 ;
        RECT 73.910 143.475 74.080 143.705 ;
        RECT 73.250 143.175 74.080 143.475 ;
        RECT 74.465 143.205 74.930 143.535 ;
        RECT 73.250 143.145 73.450 143.175 ;
        RECT 73.570 142.925 73.740 142.995 ;
        RECT 72.870 142.755 73.740 142.925 ;
        RECT 73.230 142.665 73.740 142.755 ;
        RECT 71.780 142.200 72.085 142.330 ;
        RECT 72.530 142.220 73.060 142.585 ;
        RECT 71.400 141.605 71.665 142.065 ;
        RECT 71.835 141.775 72.085 142.200 ;
        RECT 73.230 142.050 73.400 142.665 ;
        RECT 72.295 141.880 73.400 142.050 ;
        RECT 73.570 141.605 73.740 142.405 ;
        RECT 73.910 142.105 74.080 143.175 ;
        RECT 74.250 142.275 74.440 142.995 ;
        RECT 74.610 142.245 74.930 143.205 ;
        RECT 75.100 143.245 75.270 143.705 ;
        RECT 75.545 143.625 75.755 144.155 ;
        RECT 76.015 143.415 76.345 143.940 ;
        RECT 76.515 143.545 76.685 144.155 ;
        RECT 76.855 143.500 77.185 143.935 ;
        RECT 77.405 143.610 82.750 144.155 ;
        RECT 82.925 143.610 88.270 144.155 ;
        RECT 76.855 143.415 77.235 143.500 ;
        RECT 76.145 143.245 76.345 143.415 ;
        RECT 77.010 143.375 77.235 143.415 ;
        RECT 75.100 142.915 75.975 143.245 ;
        RECT 76.145 142.915 76.895 143.245 ;
        RECT 73.910 141.775 74.160 142.105 ;
        RECT 75.100 142.075 75.270 142.915 ;
        RECT 76.145 142.710 76.335 142.915 ;
        RECT 77.065 142.795 77.235 143.375 ;
        RECT 77.020 142.745 77.235 142.795 ;
        RECT 78.990 142.780 79.330 143.610 ;
        RECT 75.440 142.335 76.335 142.710 ;
        RECT 76.845 142.665 77.235 142.745 ;
        RECT 74.385 141.905 75.270 142.075 ;
        RECT 75.450 141.605 75.765 142.105 ;
        RECT 75.995 141.775 76.335 142.335 ;
        RECT 76.505 141.605 76.675 142.615 ;
        RECT 76.845 141.820 77.175 142.665 ;
        RECT 80.810 142.040 81.160 143.290 ;
        RECT 84.510 142.780 84.850 143.610 ;
        RECT 88.445 143.385 90.115 144.155 ;
        RECT 90.745 143.405 91.955 144.155 ;
        RECT 86.330 142.040 86.680 143.290 ;
        RECT 88.445 142.865 89.195 143.385 ;
        RECT 89.365 142.695 90.115 143.215 ;
        RECT 77.405 141.605 82.750 142.040 ;
        RECT 82.925 141.605 88.270 142.040 ;
        RECT 88.445 141.605 90.115 142.695 ;
        RECT 90.745 142.695 91.265 143.235 ;
        RECT 91.435 142.865 91.955 143.405 ;
        RECT 100.140 144.150 106.370 144.320 ;
        RECT 90.745 141.605 91.955 142.695 ;
        RECT 13.380 141.435 92.040 141.605 ;
        RECT 13.465 140.345 14.675 141.435 ;
        RECT 14.845 140.345 18.355 141.435 ;
        RECT 19.075 140.765 19.245 141.265 ;
        RECT 19.415 140.935 19.745 141.435 ;
        RECT 19.075 140.595 19.740 140.765 ;
        RECT 13.465 139.635 13.985 140.175 ;
        RECT 14.155 139.805 14.675 140.345 ;
        RECT 14.845 139.655 16.495 140.175 ;
        RECT 16.665 139.825 18.355 140.345 ;
        RECT 18.990 139.775 19.340 140.425 ;
        RECT 13.465 138.885 14.675 139.635 ;
        RECT 14.845 138.885 18.355 139.655 ;
        RECT 19.510 139.605 19.740 140.595 ;
        RECT 19.075 139.435 19.740 139.605 ;
        RECT 19.075 139.145 19.245 139.435 ;
        RECT 19.415 138.885 19.745 139.265 ;
        RECT 19.915 139.145 20.100 141.265 ;
        RECT 20.340 140.975 20.605 141.435 ;
        RECT 20.775 140.840 21.025 141.265 ;
        RECT 21.235 140.990 22.340 141.160 ;
        RECT 20.720 140.710 21.025 140.840 ;
        RECT 20.270 139.515 20.550 140.465 ;
        RECT 20.720 139.605 20.890 140.710 ;
        RECT 21.060 139.925 21.300 140.520 ;
        RECT 21.470 140.455 22.000 140.820 ;
        RECT 21.470 139.755 21.640 140.455 ;
        RECT 22.170 140.375 22.340 140.990 ;
        RECT 22.510 140.635 22.680 141.435 ;
        RECT 22.850 140.935 23.100 141.265 ;
        RECT 23.325 140.965 24.210 141.135 ;
        RECT 22.170 140.285 22.680 140.375 ;
        RECT 20.720 139.475 20.945 139.605 ;
        RECT 21.115 139.535 21.640 139.755 ;
        RECT 21.810 140.115 22.680 140.285 ;
        RECT 20.355 138.885 20.605 139.345 ;
        RECT 20.775 139.335 20.945 139.475 ;
        RECT 21.810 139.335 21.980 140.115 ;
        RECT 22.510 140.045 22.680 140.115 ;
        RECT 22.190 139.865 22.390 139.895 ;
        RECT 22.850 139.865 23.020 140.935 ;
        RECT 23.190 140.045 23.380 140.765 ;
        RECT 22.190 139.565 23.020 139.865 ;
        RECT 23.550 139.835 23.870 140.795 ;
        RECT 20.775 139.165 21.110 139.335 ;
        RECT 21.305 139.165 21.980 139.335 ;
        RECT 22.300 138.885 22.670 139.385 ;
        RECT 22.850 139.335 23.020 139.565 ;
        RECT 23.405 139.505 23.870 139.835 ;
        RECT 24.040 140.125 24.210 140.965 ;
        RECT 24.390 140.935 24.705 141.435 ;
        RECT 24.935 140.705 25.275 141.265 ;
        RECT 24.380 140.330 25.275 140.705 ;
        RECT 25.445 140.425 25.615 141.435 ;
        RECT 25.085 140.125 25.275 140.330 ;
        RECT 25.785 140.375 26.115 141.220 ;
        RECT 25.785 140.295 26.175 140.375 ;
        RECT 25.960 140.245 26.175 140.295 ;
        RECT 26.345 140.270 26.635 141.435 ;
        RECT 27.265 140.465 27.535 141.235 ;
        RECT 27.705 140.655 28.035 141.435 ;
        RECT 28.240 140.830 28.425 141.235 ;
        RECT 28.595 141.010 28.930 141.435 ;
        RECT 28.240 140.655 28.905 140.830 ;
        RECT 27.265 140.295 28.395 140.465 ;
        RECT 24.040 139.795 24.915 140.125 ;
        RECT 25.085 139.795 25.835 140.125 ;
        RECT 24.040 139.335 24.210 139.795 ;
        RECT 25.085 139.625 25.285 139.795 ;
        RECT 26.005 139.665 26.175 140.245 ;
        RECT 25.950 139.625 26.175 139.665 ;
        RECT 22.850 139.165 23.255 139.335 ;
        RECT 23.425 139.165 24.210 139.335 ;
        RECT 24.485 138.885 24.695 139.415 ;
        RECT 24.955 139.100 25.285 139.625 ;
        RECT 25.795 139.540 26.175 139.625 ;
        RECT 25.455 138.885 25.625 139.495 ;
        RECT 25.795 139.105 26.125 139.540 ;
        RECT 26.345 138.885 26.635 139.610 ;
        RECT 27.265 139.385 27.435 140.295 ;
        RECT 27.605 139.545 27.965 140.125 ;
        RECT 28.145 139.795 28.395 140.295 ;
        RECT 28.565 139.625 28.905 140.655 ;
        RECT 29.165 140.375 29.495 141.220 ;
        RECT 29.665 140.425 29.835 141.435 ;
        RECT 30.005 140.705 30.345 141.265 ;
        RECT 30.575 140.935 30.890 141.435 ;
        RECT 31.070 140.965 31.955 141.135 ;
        RECT 28.220 139.455 28.905 139.625 ;
        RECT 29.105 140.295 29.495 140.375 ;
        RECT 30.005 140.330 30.900 140.705 ;
        RECT 29.105 140.245 29.320 140.295 ;
        RECT 29.105 139.665 29.275 140.245 ;
        RECT 30.005 140.125 30.195 140.330 ;
        RECT 31.070 140.125 31.240 140.965 ;
        RECT 32.180 140.935 32.430 141.265 ;
        RECT 29.445 139.795 30.195 140.125 ;
        RECT 30.365 139.795 31.240 140.125 ;
        RECT 29.105 139.625 29.330 139.665 ;
        RECT 29.995 139.625 30.195 139.795 ;
        RECT 29.105 139.540 29.485 139.625 ;
        RECT 27.265 139.055 27.525 139.385 ;
        RECT 27.735 138.885 28.010 139.365 ;
        RECT 28.220 139.055 28.425 139.455 ;
        RECT 28.595 138.885 28.930 139.285 ;
        RECT 29.155 139.105 29.485 139.540 ;
        RECT 29.655 138.885 29.825 139.495 ;
        RECT 29.995 139.100 30.325 139.625 ;
        RECT 30.585 138.885 30.795 139.415 ;
        RECT 31.070 139.335 31.240 139.795 ;
        RECT 31.410 139.835 31.730 140.795 ;
        RECT 31.900 140.045 32.090 140.765 ;
        RECT 32.260 139.865 32.430 140.935 ;
        RECT 32.600 140.635 32.770 141.435 ;
        RECT 32.940 140.990 34.045 141.160 ;
        RECT 32.940 140.375 33.110 140.990 ;
        RECT 34.255 140.840 34.505 141.265 ;
        RECT 34.675 140.975 34.940 141.435 ;
        RECT 33.280 140.455 33.810 140.820 ;
        RECT 34.255 140.710 34.560 140.840 ;
        RECT 32.600 140.285 33.110 140.375 ;
        RECT 32.600 140.115 33.470 140.285 ;
        RECT 32.600 140.045 32.770 140.115 ;
        RECT 32.890 139.865 33.090 139.895 ;
        RECT 31.410 139.505 31.875 139.835 ;
        RECT 32.260 139.565 33.090 139.865 ;
        RECT 32.260 139.335 32.430 139.565 ;
        RECT 31.070 139.165 31.855 139.335 ;
        RECT 32.025 139.165 32.430 139.335 ;
        RECT 32.610 138.885 32.980 139.385 ;
        RECT 33.300 139.335 33.470 140.115 ;
        RECT 33.640 139.755 33.810 140.455 ;
        RECT 33.980 139.925 34.220 140.520 ;
        RECT 33.640 139.535 34.165 139.755 ;
        RECT 34.390 139.605 34.560 140.710 ;
        RECT 34.335 139.475 34.560 139.605 ;
        RECT 34.730 139.515 35.010 140.465 ;
        RECT 34.335 139.335 34.505 139.475 ;
        RECT 33.300 139.165 33.975 139.335 ;
        RECT 34.170 139.165 34.505 139.335 ;
        RECT 34.675 138.885 34.925 139.345 ;
        RECT 35.180 139.145 35.365 141.265 ;
        RECT 35.535 140.935 35.865 141.435 ;
        RECT 36.035 140.765 36.205 141.265 ;
        RECT 35.540 140.595 36.205 140.765 ;
        RECT 35.540 139.605 35.770 140.595 ;
        RECT 35.940 139.775 36.290 140.425 ;
        RECT 36.465 140.295 36.850 141.265 ;
        RECT 37.020 140.975 37.345 141.435 ;
        RECT 37.865 140.805 38.145 141.265 ;
        RECT 37.020 140.585 38.145 140.805 ;
        RECT 36.465 139.625 36.745 140.295 ;
        RECT 37.020 140.125 37.470 140.585 ;
        RECT 38.335 140.415 38.735 141.265 ;
        RECT 39.135 140.975 39.405 141.435 ;
        RECT 39.575 140.805 39.860 141.265 ;
        RECT 36.915 139.795 37.470 140.125 ;
        RECT 37.640 139.855 38.735 140.415 ;
        RECT 37.020 139.685 37.470 139.795 ;
        RECT 35.540 139.435 36.205 139.605 ;
        RECT 35.535 138.885 35.865 139.265 ;
        RECT 36.035 139.145 36.205 139.435 ;
        RECT 36.465 139.055 36.850 139.625 ;
        RECT 37.020 139.515 38.145 139.685 ;
        RECT 37.020 138.885 37.345 139.345 ;
        RECT 37.865 139.055 38.145 139.515 ;
        RECT 38.335 139.055 38.735 139.855 ;
        RECT 38.905 140.585 39.860 140.805 ;
        RECT 38.905 139.685 39.115 140.585 ;
        RECT 39.285 139.855 39.975 140.415 ;
        RECT 40.145 140.345 41.815 141.435 ;
        RECT 42.075 140.765 42.245 141.265 ;
        RECT 42.415 140.935 42.745 141.435 ;
        RECT 42.075 140.595 42.740 140.765 ;
        RECT 38.905 139.515 39.860 139.685 ;
        RECT 39.135 138.885 39.405 139.345 ;
        RECT 39.575 139.055 39.860 139.515 ;
        RECT 40.145 139.655 40.895 140.175 ;
        RECT 41.065 139.825 41.815 140.345 ;
        RECT 41.990 139.775 42.340 140.425 ;
        RECT 40.145 138.885 41.815 139.655 ;
        RECT 42.510 139.605 42.740 140.595 ;
        RECT 42.075 139.435 42.740 139.605 ;
        RECT 42.075 139.145 42.245 139.435 ;
        RECT 42.415 138.885 42.745 139.265 ;
        RECT 42.915 139.145 43.100 141.265 ;
        RECT 43.340 140.975 43.605 141.435 ;
        RECT 43.775 140.840 44.025 141.265 ;
        RECT 44.235 140.990 45.340 141.160 ;
        RECT 43.720 140.710 44.025 140.840 ;
        RECT 43.270 139.515 43.550 140.465 ;
        RECT 43.720 139.605 43.890 140.710 ;
        RECT 44.060 139.925 44.300 140.520 ;
        RECT 44.470 140.455 45.000 140.820 ;
        RECT 44.470 139.755 44.640 140.455 ;
        RECT 45.170 140.375 45.340 140.990 ;
        RECT 45.510 140.635 45.680 141.435 ;
        RECT 45.850 140.935 46.100 141.265 ;
        RECT 46.325 140.965 47.210 141.135 ;
        RECT 45.170 140.285 45.680 140.375 ;
        RECT 43.720 139.475 43.945 139.605 ;
        RECT 44.115 139.535 44.640 139.755 ;
        RECT 44.810 140.115 45.680 140.285 ;
        RECT 43.355 138.885 43.605 139.345 ;
        RECT 43.775 139.335 43.945 139.475 ;
        RECT 44.810 139.335 44.980 140.115 ;
        RECT 45.510 140.045 45.680 140.115 ;
        RECT 45.190 139.865 45.390 139.895 ;
        RECT 45.850 139.865 46.020 140.935 ;
        RECT 46.190 140.045 46.380 140.765 ;
        RECT 45.190 139.565 46.020 139.865 ;
        RECT 46.550 139.835 46.870 140.795 ;
        RECT 43.775 139.165 44.110 139.335 ;
        RECT 44.305 139.165 44.980 139.335 ;
        RECT 45.300 138.885 45.670 139.385 ;
        RECT 45.850 139.335 46.020 139.565 ;
        RECT 46.405 139.505 46.870 139.835 ;
        RECT 47.040 140.125 47.210 140.965 ;
        RECT 47.390 140.935 47.705 141.435 ;
        RECT 47.935 140.705 48.275 141.265 ;
        RECT 47.380 140.330 48.275 140.705 ;
        RECT 48.445 140.425 48.615 141.435 ;
        RECT 48.085 140.125 48.275 140.330 ;
        RECT 48.785 140.375 49.115 141.220 ;
        RECT 49.805 140.880 50.410 141.435 ;
        RECT 50.585 140.925 51.065 141.265 ;
        RECT 51.235 140.890 51.490 141.435 ;
        RECT 49.805 140.780 50.420 140.880 ;
        RECT 50.235 140.755 50.420 140.780 ;
        RECT 48.785 140.295 49.175 140.375 ;
        RECT 48.960 140.245 49.175 140.295 ;
        RECT 47.040 139.795 47.915 140.125 ;
        RECT 48.085 139.795 48.835 140.125 ;
        RECT 47.040 139.335 47.210 139.795 ;
        RECT 48.085 139.625 48.285 139.795 ;
        RECT 49.005 139.665 49.175 140.245 ;
        RECT 49.805 140.160 50.065 140.610 ;
        RECT 50.235 140.510 50.565 140.755 ;
        RECT 50.735 140.435 51.490 140.685 ;
        RECT 51.660 140.565 51.935 141.265 ;
        RECT 50.720 140.400 51.490 140.435 ;
        RECT 50.705 140.390 51.490 140.400 ;
        RECT 50.700 140.375 51.595 140.390 ;
        RECT 50.680 140.360 51.595 140.375 ;
        RECT 50.660 140.350 51.595 140.360 ;
        RECT 50.635 140.340 51.595 140.350 ;
        RECT 50.565 140.310 51.595 140.340 ;
        RECT 50.545 140.280 51.595 140.310 ;
        RECT 50.525 140.250 51.595 140.280 ;
        RECT 50.495 140.225 51.595 140.250 ;
        RECT 50.460 140.190 51.595 140.225 ;
        RECT 50.430 140.185 51.595 140.190 ;
        RECT 50.430 140.180 50.820 140.185 ;
        RECT 50.430 140.170 50.795 140.180 ;
        RECT 50.430 140.165 50.780 140.170 ;
        RECT 50.430 140.160 50.765 140.165 ;
        RECT 49.805 140.155 50.765 140.160 ;
        RECT 49.805 140.145 50.755 140.155 ;
        RECT 49.805 140.140 50.745 140.145 ;
        RECT 49.805 140.130 50.735 140.140 ;
        RECT 49.805 140.120 50.730 140.130 ;
        RECT 49.805 140.115 50.725 140.120 ;
        RECT 49.805 140.100 50.715 140.115 ;
        RECT 49.805 140.085 50.710 140.100 ;
        RECT 49.805 140.060 50.700 140.085 ;
        RECT 49.805 139.990 50.695 140.060 ;
        RECT 48.950 139.625 49.175 139.665 ;
        RECT 45.850 139.165 46.255 139.335 ;
        RECT 46.425 139.165 47.210 139.335 ;
        RECT 47.485 138.885 47.695 139.415 ;
        RECT 47.955 139.100 48.285 139.625 ;
        RECT 48.795 139.540 49.175 139.625 ;
        RECT 48.455 138.885 48.625 139.495 ;
        RECT 48.795 139.105 49.125 139.540 ;
        RECT 49.805 139.435 50.355 139.820 ;
        RECT 50.525 139.265 50.695 139.990 ;
        RECT 49.805 139.095 50.695 139.265 ;
        RECT 50.865 139.590 51.195 140.015 ;
        RECT 51.365 139.790 51.595 140.185 ;
        RECT 50.865 139.565 51.115 139.590 ;
        RECT 50.865 139.105 51.085 139.565 ;
        RECT 51.765 139.535 51.935 140.565 ;
        RECT 52.105 140.270 52.395 141.435 ;
        RECT 52.650 140.815 52.825 141.265 ;
        RECT 52.995 140.995 53.325 141.435 ;
        RECT 53.630 140.845 53.800 141.265 ;
        RECT 54.035 141.025 54.705 141.435 ;
        RECT 54.920 140.845 55.090 141.265 ;
        RECT 55.290 141.025 55.620 141.435 ;
        RECT 52.650 140.645 53.280 140.815 ;
        RECT 52.565 139.795 52.930 140.475 ;
        RECT 53.110 140.125 53.280 140.645 ;
        RECT 53.630 140.675 55.645 140.845 ;
        RECT 53.110 139.795 53.460 140.125 ;
        RECT 53.110 139.625 53.280 139.795 ;
        RECT 51.255 138.885 51.505 139.425 ;
        RECT 51.675 139.055 51.935 139.535 ;
        RECT 52.105 138.885 52.395 139.610 ;
        RECT 52.650 139.455 53.280 139.625 ;
        RECT 52.650 139.055 52.825 139.455 ;
        RECT 53.630 139.385 53.800 140.675 ;
        RECT 52.995 138.885 53.325 139.265 ;
        RECT 53.570 139.055 53.800 139.385 ;
        RECT 54.000 139.220 54.280 140.495 ;
        RECT 54.505 139.395 54.775 140.495 ;
        RECT 54.965 139.465 55.305 140.495 ;
        RECT 55.475 140.125 55.645 140.675 ;
        RECT 55.815 140.295 56.075 141.265 ;
        RECT 56.255 140.485 56.530 141.255 ;
        RECT 56.700 140.825 57.030 141.255 ;
        RECT 57.200 140.995 57.395 141.435 ;
        RECT 57.575 140.825 57.905 141.255 ;
        RECT 56.700 140.655 57.905 140.825 ;
        RECT 58.335 140.705 58.630 141.435 ;
        RECT 56.255 140.295 56.840 140.485 ;
        RECT 57.010 140.325 57.905 140.655 ;
        RECT 58.800 140.535 59.060 141.260 ;
        RECT 59.230 140.705 59.490 141.435 ;
        RECT 59.660 140.535 59.920 141.260 ;
        RECT 60.090 140.705 60.350 141.435 ;
        RECT 60.520 140.535 60.780 141.260 ;
        RECT 60.950 140.705 61.210 141.435 ;
        RECT 61.380 140.535 61.640 141.260 ;
        RECT 55.475 139.795 55.735 140.125 ;
        RECT 55.905 139.605 56.075 140.295 ;
        RECT 54.465 139.225 54.775 139.395 ;
        RECT 54.505 139.220 54.775 139.225 ;
        RECT 55.235 138.885 55.565 139.265 ;
        RECT 55.735 139.140 56.075 139.605 ;
        RECT 56.255 139.475 56.495 140.125 ;
        RECT 56.665 139.625 56.840 140.295 ;
        RECT 58.330 140.295 61.640 140.535 ;
        RECT 61.810 140.325 62.070 141.435 ;
        RECT 57.010 139.795 57.425 140.125 ;
        RECT 57.605 139.795 57.900 140.125 ;
        RECT 56.665 139.445 56.995 139.625 ;
        RECT 55.735 139.095 56.070 139.140 ;
        RECT 56.270 138.885 56.600 139.275 ;
        RECT 56.770 139.065 56.995 139.445 ;
        RECT 57.195 139.175 57.425 139.795 ;
        RECT 58.330 139.705 59.300 140.295 ;
        RECT 62.240 140.125 62.490 141.260 ;
        RECT 62.670 140.325 62.965 141.435 ;
        RECT 63.145 140.345 64.355 141.435 ;
        RECT 59.470 139.875 62.490 140.125 ;
        RECT 57.605 138.885 57.905 139.615 ;
        RECT 58.330 139.535 61.640 139.705 ;
        RECT 58.330 138.885 58.630 139.365 ;
        RECT 58.800 139.080 59.060 139.535 ;
        RECT 59.230 138.885 59.490 139.365 ;
        RECT 59.660 139.080 59.920 139.535 ;
        RECT 60.090 138.885 60.350 139.365 ;
        RECT 60.520 139.080 60.780 139.535 ;
        RECT 60.950 138.885 61.210 139.365 ;
        RECT 61.380 139.080 61.640 139.535 ;
        RECT 61.810 138.885 62.070 139.410 ;
        RECT 62.240 139.065 62.490 139.875 ;
        RECT 62.660 139.515 62.975 140.125 ;
        RECT 63.145 139.635 63.665 140.175 ;
        RECT 63.835 139.805 64.355 140.345 ;
        RECT 64.525 141.005 64.865 141.265 ;
        RECT 62.670 138.885 62.915 139.345 ;
        RECT 63.145 138.885 64.355 139.635 ;
        RECT 64.525 139.605 64.785 141.005 ;
        RECT 65.035 140.635 65.365 141.435 ;
        RECT 65.830 140.465 66.080 141.265 ;
        RECT 66.265 140.715 66.595 141.435 ;
        RECT 66.815 140.465 67.065 141.265 ;
        RECT 67.235 141.055 67.570 141.435 ;
        RECT 67.745 141.000 73.090 141.435 ;
        RECT 64.975 140.295 67.165 140.465 ;
        RECT 64.975 140.125 65.290 140.295 ;
        RECT 64.960 139.875 65.290 140.125 ;
        RECT 64.525 139.095 64.865 139.605 ;
        RECT 65.035 138.885 65.305 139.685 ;
        RECT 65.485 139.155 65.765 140.125 ;
        RECT 65.945 139.155 66.245 140.125 ;
        RECT 66.425 139.160 66.775 140.125 ;
        RECT 66.995 139.385 67.165 140.295 ;
        RECT 67.335 139.565 67.575 140.875 ;
        RECT 69.330 139.430 69.670 140.260 ;
        RECT 71.150 139.750 71.500 141.000 ;
        RECT 73.265 140.345 76.775 141.435 ;
        RECT 73.265 139.655 74.915 140.175 ;
        RECT 75.085 139.825 76.775 140.345 ;
        RECT 77.865 140.270 78.155 141.435 ;
        RECT 78.325 141.000 83.670 141.435 ;
        RECT 83.845 141.000 89.190 141.435 ;
        RECT 66.995 139.055 67.490 139.385 ;
        RECT 67.745 138.885 73.090 139.430 ;
        RECT 73.265 138.885 76.775 139.655 ;
        RECT 77.865 138.885 78.155 139.610 ;
        RECT 79.910 139.430 80.250 140.260 ;
        RECT 81.730 139.750 82.080 141.000 ;
        RECT 85.430 139.430 85.770 140.260 ;
        RECT 87.250 139.750 87.600 141.000 ;
        RECT 89.365 140.345 90.575 141.435 ;
        RECT 89.365 139.635 89.885 140.175 ;
        RECT 90.055 139.805 90.575 140.345 ;
        RECT 90.745 140.345 91.955 141.435 ;
        RECT 100.140 140.890 100.810 144.150 ;
        RECT 101.480 143.580 105.520 143.750 ;
        RECT 101.140 141.520 101.310 143.520 ;
        RECT 105.690 141.520 105.860 143.520 ;
        RECT 101.480 141.290 105.520 141.460 ;
        RECT 106.200 140.890 106.370 144.150 ;
        RECT 100.140 140.720 106.370 140.890 ;
        RECT 90.745 139.805 91.265 140.345 ;
        RECT 91.435 139.635 91.955 140.175 ;
        RECT 78.325 138.885 83.670 139.430 ;
        RECT 83.845 138.885 89.190 139.430 ;
        RECT 89.365 138.885 90.575 139.635 ;
        RECT 90.745 138.885 91.955 139.635 ;
        RECT 13.380 138.715 92.040 138.885 ;
        RECT 13.465 137.965 14.675 138.715 ;
        RECT 13.465 137.425 13.985 137.965 ;
        RECT 14.850 137.875 15.110 138.715 ;
        RECT 15.285 137.970 15.540 138.545 ;
        RECT 15.710 138.335 16.040 138.715 ;
        RECT 16.255 138.165 16.425 138.545 ;
        RECT 15.710 137.995 16.425 138.165 ;
        RECT 14.155 137.255 14.675 137.795 ;
        RECT 13.465 136.165 14.675 137.255 ;
        RECT 14.850 136.165 15.110 137.315 ;
        RECT 15.285 137.240 15.455 137.970 ;
        RECT 15.710 137.805 15.880 137.995 ;
        RECT 16.685 137.945 20.195 138.715 ;
        RECT 21.285 138.065 21.545 138.545 ;
        RECT 21.715 138.255 22.045 138.715 ;
        RECT 22.235 138.075 22.435 138.495 ;
        RECT 15.625 137.475 15.880 137.805 ;
        RECT 15.710 137.265 15.880 137.475 ;
        RECT 16.160 137.445 16.515 137.815 ;
        RECT 16.685 137.425 18.335 137.945 ;
        RECT 15.285 136.335 15.540 137.240 ;
        RECT 15.710 137.095 16.425 137.265 ;
        RECT 18.505 137.255 20.195 137.775 ;
        RECT 15.710 136.165 16.040 136.925 ;
        RECT 16.255 136.335 16.425 137.095 ;
        RECT 16.685 136.165 20.195 137.255 ;
        RECT 21.285 137.035 21.455 138.065 ;
        RECT 21.625 137.375 21.855 137.805 ;
        RECT 22.025 137.555 22.435 138.075 ;
        RECT 22.605 138.230 23.395 138.495 ;
        RECT 22.605 137.375 22.860 138.230 ;
        RECT 23.575 137.895 23.905 138.315 ;
        RECT 24.075 137.895 24.335 138.715 ;
        RECT 24.505 137.965 25.715 138.715 ;
        RECT 26.050 138.205 26.290 138.715 ;
        RECT 26.470 138.205 26.750 138.535 ;
        RECT 26.980 138.205 27.195 138.715 ;
        RECT 23.575 137.805 23.825 137.895 ;
        RECT 23.030 137.555 23.825 137.805 ;
        RECT 21.625 137.205 23.415 137.375 ;
        RECT 21.285 136.335 21.560 137.035 ;
        RECT 21.730 136.910 22.445 137.205 ;
        RECT 22.665 136.845 22.995 137.035 ;
        RECT 21.770 136.165 21.985 136.710 ;
        RECT 22.155 136.335 22.630 136.675 ;
        RECT 22.800 136.670 22.995 136.845 ;
        RECT 23.165 136.840 23.415 137.205 ;
        RECT 22.800 136.165 23.415 136.670 ;
        RECT 23.655 136.335 23.825 137.555 ;
        RECT 23.995 136.845 24.335 137.725 ;
        RECT 24.505 137.425 25.025 137.965 ;
        RECT 25.195 137.255 25.715 137.795 ;
        RECT 25.945 137.475 26.300 138.035 ;
        RECT 26.470 137.305 26.640 138.205 ;
        RECT 26.810 137.475 27.075 138.035 ;
        RECT 27.365 137.975 27.980 138.545 ;
        RECT 28.185 138.335 29.075 138.505 ;
        RECT 27.325 137.305 27.495 137.805 ;
        RECT 24.075 136.165 24.335 136.675 ;
        RECT 24.505 136.165 25.715 137.255 ;
        RECT 26.070 137.135 27.495 137.305 ;
        RECT 26.070 136.960 26.460 137.135 ;
        RECT 26.945 136.165 27.275 136.965 ;
        RECT 27.665 136.955 27.980 137.975 ;
        RECT 28.185 137.780 28.735 138.165 ;
        RECT 28.905 137.610 29.075 138.335 ;
        RECT 28.185 137.540 29.075 137.610 ;
        RECT 29.245 138.010 29.465 138.495 ;
        RECT 29.635 138.175 29.885 138.715 ;
        RECT 30.055 138.065 30.315 138.545 ;
        RECT 29.245 137.585 29.575 138.010 ;
        RECT 28.185 137.515 29.080 137.540 ;
        RECT 28.185 137.500 29.090 137.515 ;
        RECT 28.185 137.485 29.095 137.500 ;
        RECT 28.185 137.480 29.105 137.485 ;
        RECT 28.185 137.470 29.110 137.480 ;
        RECT 28.185 137.460 29.115 137.470 ;
        RECT 28.185 137.455 29.125 137.460 ;
        RECT 28.185 137.445 29.135 137.455 ;
        RECT 28.185 137.440 29.145 137.445 ;
        RECT 28.185 136.990 28.445 137.440 ;
        RECT 28.810 137.435 29.145 137.440 ;
        RECT 28.810 137.430 29.160 137.435 ;
        RECT 28.810 137.420 29.175 137.430 ;
        RECT 28.810 137.415 29.200 137.420 ;
        RECT 29.745 137.415 29.975 137.810 ;
        RECT 28.810 137.410 29.975 137.415 ;
        RECT 28.840 137.375 29.975 137.410 ;
        RECT 28.875 137.350 29.975 137.375 ;
        RECT 28.905 137.320 29.975 137.350 ;
        RECT 28.925 137.290 29.975 137.320 ;
        RECT 28.945 137.260 29.975 137.290 ;
        RECT 29.015 137.250 29.975 137.260 ;
        RECT 29.040 137.240 29.975 137.250 ;
        RECT 29.060 137.225 29.975 137.240 ;
        RECT 29.080 137.210 29.975 137.225 ;
        RECT 29.085 137.200 29.870 137.210 ;
        RECT 29.100 137.165 29.870 137.200 ;
        RECT 27.445 136.335 27.980 136.955 ;
        RECT 28.615 136.845 28.945 137.090 ;
        RECT 29.115 136.915 29.870 137.165 ;
        RECT 30.145 137.035 30.315 138.065 ;
        RECT 30.575 138.165 30.745 138.455 ;
        RECT 30.915 138.335 31.245 138.715 ;
        RECT 30.575 137.995 31.240 138.165 ;
        RECT 30.490 137.175 30.840 137.825 ;
        RECT 28.615 136.820 28.800 136.845 ;
        RECT 28.185 136.720 28.800 136.820 ;
        RECT 28.185 136.165 28.790 136.720 ;
        RECT 28.965 136.335 29.445 136.675 ;
        RECT 29.615 136.165 29.870 136.710 ;
        RECT 30.040 136.335 30.315 137.035 ;
        RECT 31.010 137.005 31.240 137.995 ;
        RECT 30.575 136.835 31.240 137.005 ;
        RECT 30.575 136.335 30.745 136.835 ;
        RECT 30.915 136.165 31.245 136.665 ;
        RECT 31.415 136.335 31.600 138.455 ;
        RECT 31.855 138.255 32.105 138.715 ;
        RECT 32.275 138.265 32.610 138.435 ;
        RECT 32.805 138.265 33.480 138.435 ;
        RECT 32.275 138.125 32.445 138.265 ;
        RECT 31.770 137.135 32.050 138.085 ;
        RECT 32.220 137.995 32.445 138.125 ;
        RECT 32.220 136.890 32.390 137.995 ;
        RECT 32.615 137.845 33.140 138.065 ;
        RECT 32.560 137.080 32.800 137.675 ;
        RECT 32.970 137.145 33.140 137.845 ;
        RECT 33.310 137.485 33.480 138.265 ;
        RECT 33.800 138.215 34.170 138.715 ;
        RECT 34.350 138.265 34.755 138.435 ;
        RECT 34.925 138.265 35.710 138.435 ;
        RECT 34.350 138.035 34.520 138.265 ;
        RECT 33.690 137.735 34.520 138.035 ;
        RECT 34.905 137.765 35.370 138.095 ;
        RECT 33.690 137.705 33.890 137.735 ;
        RECT 34.010 137.485 34.180 137.555 ;
        RECT 33.310 137.315 34.180 137.485 ;
        RECT 33.670 137.225 34.180 137.315 ;
        RECT 32.220 136.760 32.525 136.890 ;
        RECT 32.970 136.780 33.500 137.145 ;
        RECT 31.840 136.165 32.105 136.625 ;
        RECT 32.275 136.335 32.525 136.760 ;
        RECT 33.670 136.610 33.840 137.225 ;
        RECT 32.735 136.440 33.840 136.610 ;
        RECT 34.010 136.165 34.180 136.965 ;
        RECT 34.350 136.665 34.520 137.735 ;
        RECT 34.690 136.835 34.880 137.555 ;
        RECT 35.050 136.805 35.370 137.765 ;
        RECT 35.540 137.805 35.710 138.265 ;
        RECT 35.985 138.185 36.195 138.715 ;
        RECT 36.455 137.975 36.785 138.500 ;
        RECT 36.955 138.105 37.125 138.715 ;
        RECT 37.295 138.060 37.625 138.495 ;
        RECT 37.295 137.975 37.675 138.060 ;
        RECT 36.585 137.805 36.785 137.975 ;
        RECT 37.450 137.935 37.675 137.975 ;
        RECT 35.540 137.475 36.415 137.805 ;
        RECT 36.585 137.475 37.335 137.805 ;
        RECT 34.350 136.335 34.600 136.665 ;
        RECT 35.540 136.635 35.710 137.475 ;
        RECT 36.585 137.270 36.775 137.475 ;
        RECT 37.505 137.355 37.675 137.935 ;
        RECT 37.845 137.965 39.055 138.715 ;
        RECT 39.225 137.990 39.515 138.715 ;
        RECT 40.665 138.255 40.910 138.715 ;
        RECT 37.845 137.425 38.365 137.965 ;
        RECT 37.460 137.305 37.675 137.355 ;
        RECT 35.880 136.895 36.775 137.270 ;
        RECT 37.285 137.225 37.675 137.305 ;
        RECT 38.535 137.255 39.055 137.795 ;
        RECT 40.605 137.475 40.920 138.085 ;
        RECT 41.090 137.725 41.340 138.535 ;
        RECT 41.510 138.190 41.770 138.715 ;
        RECT 41.940 138.065 42.200 138.520 ;
        RECT 42.370 138.235 42.630 138.715 ;
        RECT 42.800 138.065 43.060 138.520 ;
        RECT 43.230 138.235 43.490 138.715 ;
        RECT 43.660 138.065 43.920 138.520 ;
        RECT 44.090 138.235 44.350 138.715 ;
        RECT 44.520 138.065 44.780 138.520 ;
        RECT 44.950 138.235 45.250 138.715 ;
        RECT 45.670 138.460 46.005 138.505 ;
        RECT 41.940 137.895 45.250 138.065 ;
        RECT 41.090 137.475 44.110 137.725 ;
        RECT 34.825 136.465 35.710 136.635 ;
        RECT 35.890 136.165 36.205 136.665 ;
        RECT 36.435 136.335 36.775 136.895 ;
        RECT 36.945 136.165 37.115 137.175 ;
        RECT 37.285 136.380 37.615 137.225 ;
        RECT 37.845 136.165 39.055 137.255 ;
        RECT 39.225 136.165 39.515 137.330 ;
        RECT 40.615 136.165 40.910 137.275 ;
        RECT 41.090 136.340 41.340 137.475 ;
        RECT 44.280 137.305 45.250 137.895 ;
        RECT 41.510 136.165 41.770 137.275 ;
        RECT 41.940 137.065 45.250 137.305 ;
        RECT 45.665 137.995 46.005 138.460 ;
        RECT 46.175 138.335 46.505 138.715 ;
        RECT 46.965 138.375 47.235 138.380 ;
        RECT 46.965 138.205 47.275 138.375 ;
        RECT 45.665 137.305 45.835 137.995 ;
        RECT 46.005 137.475 46.265 137.805 ;
        RECT 41.940 136.340 42.200 137.065 ;
        RECT 42.370 136.165 42.630 136.895 ;
        RECT 42.800 136.340 43.060 137.065 ;
        RECT 43.230 136.165 43.490 136.895 ;
        RECT 43.660 136.340 43.920 137.065 ;
        RECT 44.090 136.165 44.350 136.895 ;
        RECT 44.520 136.340 44.780 137.065 ;
        RECT 44.950 136.165 45.245 136.895 ;
        RECT 45.665 136.335 45.925 137.305 ;
        RECT 46.095 136.925 46.265 137.475 ;
        RECT 46.435 137.105 46.775 138.135 ;
        RECT 46.965 137.105 47.235 138.205 ;
        RECT 47.460 137.105 47.740 138.380 ;
        RECT 47.940 138.215 48.170 138.545 ;
        RECT 48.415 138.335 48.745 138.715 ;
        RECT 47.940 136.925 48.110 138.215 ;
        RECT 48.915 138.145 49.090 138.545 ;
        RECT 48.460 137.975 49.090 138.145 ;
        RECT 49.345 137.995 49.685 138.505 ;
        RECT 48.460 137.805 48.630 137.975 ;
        RECT 48.280 137.475 48.630 137.805 ;
        RECT 46.095 136.755 48.110 136.925 ;
        RECT 48.460 136.955 48.630 137.475 ;
        RECT 48.810 137.125 49.175 137.805 ;
        RECT 48.460 136.785 49.090 136.955 ;
        RECT 46.120 136.165 46.450 136.575 ;
        RECT 46.650 136.335 46.820 136.755 ;
        RECT 47.035 136.165 47.705 136.575 ;
        RECT 47.940 136.335 48.110 136.755 ;
        RECT 48.415 136.165 48.745 136.605 ;
        RECT 48.915 136.335 49.090 136.785 ;
        RECT 49.345 136.595 49.605 137.995 ;
        RECT 49.855 137.915 50.125 138.715 ;
        RECT 49.780 137.475 50.110 137.725 ;
        RECT 50.305 137.475 50.585 138.445 ;
        RECT 50.765 137.475 51.065 138.445 ;
        RECT 51.245 137.475 51.595 138.440 ;
        RECT 51.815 138.215 52.310 138.545 ;
        RECT 49.795 137.305 50.110 137.475 ;
        RECT 51.815 137.305 51.985 138.215 ;
        RECT 49.795 137.135 51.985 137.305 ;
        RECT 49.345 136.335 49.685 136.595 ;
        RECT 49.855 136.165 50.185 136.965 ;
        RECT 50.650 136.335 50.900 137.135 ;
        RECT 51.085 136.165 51.415 136.885 ;
        RECT 51.635 136.335 51.885 137.135 ;
        RECT 52.155 136.725 52.395 138.035 ;
        RECT 52.575 137.905 52.845 138.715 ;
        RECT 53.015 137.905 53.345 138.545 ;
        RECT 53.515 137.905 53.755 138.715 ;
        RECT 53.945 137.945 57.455 138.715 ;
        RECT 58.130 138.255 58.395 138.715 ;
        RECT 58.765 138.075 58.935 138.545 ;
        RECT 59.185 138.255 59.355 138.715 ;
        RECT 59.605 138.075 59.775 138.545 ;
        RECT 60.025 138.255 60.195 138.715 ;
        RECT 60.445 138.075 60.615 138.545 ;
        RECT 60.785 138.250 61.035 138.715 ;
        RECT 52.565 137.475 52.915 137.725 ;
        RECT 53.085 137.305 53.255 137.905 ;
        RECT 53.425 137.475 53.775 137.725 ;
        RECT 53.945 137.425 55.595 137.945 ;
        RECT 58.765 137.895 61.135 138.075 ;
        RECT 52.055 136.165 52.390 136.545 ;
        RECT 52.575 136.165 52.905 137.305 ;
        RECT 53.085 137.135 53.765 137.305 ;
        RECT 55.765 137.255 57.455 137.775 ;
        RECT 58.105 137.475 60.615 137.725 ;
        RECT 60.785 137.305 61.135 137.895 ;
        RECT 61.305 137.945 64.815 138.715 ;
        RECT 64.985 137.990 65.275 138.715 ;
        RECT 65.445 137.945 67.115 138.715 ;
        RECT 61.305 137.425 62.955 137.945 ;
        RECT 53.435 136.350 53.765 137.135 ;
        RECT 53.945 136.165 57.455 137.255 ;
        RECT 58.130 136.165 58.425 137.305 ;
        RECT 58.685 137.135 61.135 137.305 ;
        RECT 63.125 137.255 64.815 137.775 ;
        RECT 65.445 137.425 66.195 137.945 ;
        RECT 67.295 137.905 67.565 138.715 ;
        RECT 67.735 137.905 68.065 138.545 ;
        RECT 68.235 137.905 68.475 138.715 ;
        RECT 68.665 137.965 69.875 138.715 ;
        RECT 70.130 138.145 70.305 138.545 ;
        RECT 70.475 138.335 70.805 138.715 ;
        RECT 71.050 138.215 71.280 138.545 ;
        RECT 70.130 137.975 70.760 138.145 ;
        RECT 58.685 136.335 59.015 137.135 ;
        RECT 59.185 136.165 59.355 136.965 ;
        RECT 59.525 136.335 59.855 137.135 ;
        RECT 60.365 137.115 61.135 137.135 ;
        RECT 60.025 136.165 60.195 136.965 ;
        RECT 60.365 136.335 60.695 137.115 ;
        RECT 60.865 136.165 61.035 136.625 ;
        RECT 61.305 136.165 64.815 137.255 ;
        RECT 64.985 136.165 65.275 137.330 ;
        RECT 66.365 137.255 67.115 137.775 ;
        RECT 67.285 137.475 67.635 137.725 ;
        RECT 67.805 137.305 67.975 137.905 ;
        RECT 68.145 137.475 68.495 137.725 ;
        RECT 68.665 137.425 69.185 137.965 ;
        RECT 70.590 137.805 70.760 137.975 ;
        RECT 65.445 136.165 67.115 137.255 ;
        RECT 67.295 136.165 67.625 137.305 ;
        RECT 67.805 137.135 68.485 137.305 ;
        RECT 69.355 137.255 69.875 137.795 ;
        RECT 68.155 136.350 68.485 137.135 ;
        RECT 68.665 136.165 69.875 137.255 ;
        RECT 70.045 137.125 70.410 137.805 ;
        RECT 70.590 137.475 70.940 137.805 ;
        RECT 70.590 136.955 70.760 137.475 ;
        RECT 70.130 136.785 70.760 136.955 ;
        RECT 71.110 136.925 71.280 138.215 ;
        RECT 71.480 137.105 71.760 138.380 ;
        RECT 71.985 138.375 72.255 138.380 ;
        RECT 71.945 138.205 72.255 138.375 ;
        RECT 72.715 138.335 73.045 138.715 ;
        RECT 73.215 138.460 73.550 138.505 ;
        RECT 71.985 137.105 72.255 138.205 ;
        RECT 72.445 137.105 72.785 138.135 ;
        RECT 73.215 137.995 73.555 138.460 ;
        RECT 73.775 138.060 74.105 138.495 ;
        RECT 74.275 138.105 74.445 138.715 ;
        RECT 72.955 137.475 73.215 137.805 ;
        RECT 72.955 136.925 73.125 137.475 ;
        RECT 73.385 137.305 73.555 137.995 ;
        RECT 70.130 136.335 70.305 136.785 ;
        RECT 71.110 136.755 73.125 136.925 ;
        RECT 70.475 136.165 70.805 136.605 ;
        RECT 71.110 136.335 71.280 136.755 ;
        RECT 71.515 136.165 72.185 136.575 ;
        RECT 72.400 136.335 72.570 136.755 ;
        RECT 72.770 136.165 73.100 136.575 ;
        RECT 73.295 136.335 73.555 137.305 ;
        RECT 73.725 137.975 74.105 138.060 ;
        RECT 74.615 137.975 74.945 138.500 ;
        RECT 75.205 138.185 75.415 138.715 ;
        RECT 75.690 138.265 76.475 138.435 ;
        RECT 76.645 138.265 77.050 138.435 ;
        RECT 73.725 137.935 73.950 137.975 ;
        RECT 73.725 137.355 73.895 137.935 ;
        RECT 74.615 137.805 74.815 137.975 ;
        RECT 75.690 137.805 75.860 138.265 ;
        RECT 74.065 137.475 74.815 137.805 ;
        RECT 74.985 137.475 75.860 137.805 ;
        RECT 73.725 137.305 73.940 137.355 ;
        RECT 73.725 137.225 74.115 137.305 ;
        RECT 73.785 136.380 74.115 137.225 ;
        RECT 74.625 137.270 74.815 137.475 ;
        RECT 74.285 136.165 74.455 137.175 ;
        RECT 74.625 136.895 75.520 137.270 ;
        RECT 74.625 136.335 74.965 136.895 ;
        RECT 75.195 136.165 75.510 136.665 ;
        RECT 75.690 136.635 75.860 137.475 ;
        RECT 76.030 137.765 76.495 138.095 ;
        RECT 76.880 138.035 77.050 138.265 ;
        RECT 77.230 138.215 77.600 138.715 ;
        RECT 77.920 138.265 78.595 138.435 ;
        RECT 78.790 138.265 79.125 138.435 ;
        RECT 76.030 136.805 76.350 137.765 ;
        RECT 76.880 137.735 77.710 138.035 ;
        RECT 76.520 136.835 76.710 137.555 ;
        RECT 76.880 136.665 77.050 137.735 ;
        RECT 77.510 137.705 77.710 137.735 ;
        RECT 77.220 137.485 77.390 137.555 ;
        RECT 77.920 137.485 78.090 138.265 ;
        RECT 78.955 138.125 79.125 138.265 ;
        RECT 79.295 138.255 79.545 138.715 ;
        RECT 77.220 137.315 78.090 137.485 ;
        RECT 78.260 137.845 78.785 138.065 ;
        RECT 78.955 137.995 79.180 138.125 ;
        RECT 77.220 137.225 77.730 137.315 ;
        RECT 75.690 136.465 76.575 136.635 ;
        RECT 76.800 136.335 77.050 136.665 ;
        RECT 77.220 136.165 77.390 136.965 ;
        RECT 77.560 136.610 77.730 137.225 ;
        RECT 78.260 137.145 78.430 137.845 ;
        RECT 77.900 136.780 78.430 137.145 ;
        RECT 78.600 137.080 78.840 137.675 ;
        RECT 79.010 136.890 79.180 137.995 ;
        RECT 79.350 137.135 79.630 138.085 ;
        RECT 78.875 136.760 79.180 136.890 ;
        RECT 77.560 136.440 78.665 136.610 ;
        RECT 78.875 136.335 79.125 136.760 ;
        RECT 79.295 136.165 79.560 136.625 ;
        RECT 79.800 136.335 79.985 138.455 ;
        RECT 80.155 138.335 80.485 138.715 ;
        RECT 80.655 138.165 80.825 138.455 ;
        RECT 81.085 138.170 86.430 138.715 ;
        RECT 80.160 137.995 80.825 138.165 ;
        RECT 80.160 137.005 80.390 137.995 ;
        RECT 80.560 137.175 80.910 137.825 ;
        RECT 82.670 137.340 83.010 138.170 ;
        RECT 86.605 137.945 90.115 138.715 ;
        RECT 90.745 137.965 91.955 138.715 ;
        RECT 80.160 136.835 80.825 137.005 ;
        RECT 80.155 136.165 80.485 136.665 ;
        RECT 80.655 136.335 80.825 136.835 ;
        RECT 84.490 136.600 84.840 137.850 ;
        RECT 86.605 137.425 88.255 137.945 ;
        RECT 88.425 137.255 90.115 137.775 ;
        RECT 81.085 136.165 86.430 136.600 ;
        RECT 86.605 136.165 90.115 137.255 ;
        RECT 90.745 137.255 91.265 137.795 ;
        RECT 91.435 137.425 91.955 137.965 ;
        RECT 100.140 137.460 100.810 140.720 ;
        RECT 101.480 140.150 105.520 140.320 ;
        RECT 101.140 138.090 101.310 140.090 ;
        RECT 105.690 138.090 105.860 140.090 ;
        RECT 101.480 137.860 105.520 138.030 ;
        RECT 106.200 137.460 106.370 140.720 ;
        RECT 100.140 137.450 106.370 137.460 ;
        RECT 107.960 146.720 117.790 146.760 ;
        RECT 120.510 146.740 126.250 146.750 ;
        RECT 107.960 146.590 118.590 146.720 ;
        RECT 107.960 144.330 108.130 146.590 ;
        RECT 108.855 146.020 116.895 146.190 ;
        RECT 108.470 144.960 108.640 145.960 ;
        RECT 117.110 144.960 117.280 145.960 ;
        RECT 108.855 144.730 116.895 144.900 ;
        RECT 117.620 144.330 118.590 146.590 ;
        RECT 107.960 144.160 118.590 144.330 ;
        RECT 107.960 140.900 108.130 144.160 ;
        RECT 108.855 143.590 116.895 143.760 ;
        RECT 108.470 141.530 108.640 143.530 ;
        RECT 117.110 141.530 117.280 143.530 ;
        RECT 108.855 141.300 116.895 141.470 ;
        RECT 117.620 140.900 118.590 144.160 ;
        RECT 107.960 140.730 118.590 140.900 ;
        RECT 107.960 137.470 108.130 140.730 ;
        RECT 108.855 140.160 116.895 140.330 ;
        RECT 108.470 138.100 108.640 140.100 ;
        RECT 117.110 138.100 117.280 140.100 ;
        RECT 108.855 137.870 116.895 138.040 ;
        RECT 117.620 137.470 118.590 140.730 ;
        RECT 100.140 137.350 106.380 137.450 ;
        RECT 90.745 136.165 91.955 137.255 ;
        RECT 100.130 136.790 106.380 137.350 ;
        RECT 100.130 136.770 105.300 136.790 ;
        RECT 100.130 136.700 104.120 136.770 ;
        RECT 13.380 135.995 92.040 136.165 ;
        RECT 13.465 134.905 14.675 135.995 ;
        RECT 14.845 135.560 20.190 135.995 ;
        RECT 20.365 135.560 25.710 135.995 ;
        RECT 13.465 134.195 13.985 134.735 ;
        RECT 14.155 134.365 14.675 134.905 ;
        RECT 13.465 133.445 14.675 134.195 ;
        RECT 16.430 133.990 16.770 134.820 ;
        RECT 18.250 134.310 18.600 135.560 ;
        RECT 21.950 133.990 22.290 134.820 ;
        RECT 23.770 134.310 24.120 135.560 ;
        RECT 26.345 134.830 26.635 135.995 ;
        RECT 26.805 134.905 30.315 135.995 ;
        RECT 26.805 134.215 28.455 134.735 ;
        RECT 28.625 134.385 30.315 134.905 ;
        RECT 31.415 134.855 31.745 135.995 ;
        RECT 14.845 133.445 20.190 133.990 ;
        RECT 20.365 133.445 25.710 133.990 ;
        RECT 26.345 133.445 26.635 134.170 ;
        RECT 26.805 133.445 30.315 134.215 ;
        RECT 31.405 134.105 31.745 134.685 ;
        RECT 31.915 134.655 32.275 135.825 ;
        RECT 32.475 134.825 32.805 135.995 ;
        RECT 33.005 134.655 33.335 135.825 ;
        RECT 33.535 134.825 33.865 135.995 ;
        RECT 34.175 135.045 34.450 135.815 ;
        RECT 34.620 135.385 34.950 135.815 ;
        RECT 35.120 135.555 35.315 135.995 ;
        RECT 35.495 135.385 35.825 135.815 ;
        RECT 34.620 135.215 35.825 135.385 ;
        RECT 34.175 134.855 34.760 135.045 ;
        RECT 34.930 134.885 35.825 135.215 ;
        RECT 36.005 134.905 37.675 135.995 ;
        RECT 38.395 135.325 38.565 135.825 ;
        RECT 38.735 135.495 39.065 135.995 ;
        RECT 38.395 135.155 39.060 135.325 ;
        RECT 31.915 134.375 33.335 134.655 ;
        RECT 31.915 134.040 32.275 134.375 ;
        RECT 31.415 133.445 31.745 133.935 ;
        RECT 31.915 133.615 32.535 134.040 ;
        RECT 32.995 133.445 33.325 134.135 ;
        RECT 34.175 134.035 34.415 134.685 ;
        RECT 34.585 134.185 34.760 134.855 ;
        RECT 34.930 134.355 35.345 134.685 ;
        RECT 35.525 134.355 35.820 134.685 ;
        RECT 34.585 134.005 34.915 134.185 ;
        RECT 34.190 133.445 34.520 133.835 ;
        RECT 34.690 133.625 34.915 134.005 ;
        RECT 35.115 133.735 35.345 134.355 ;
        RECT 36.005 134.215 36.755 134.735 ;
        RECT 36.925 134.385 37.675 134.905 ;
        RECT 38.310 134.335 38.660 134.985 ;
        RECT 35.525 133.445 35.825 134.175 ;
        RECT 36.005 133.445 37.675 134.215 ;
        RECT 38.830 134.165 39.060 135.155 ;
        RECT 38.395 133.995 39.060 134.165 ;
        RECT 38.395 133.705 38.565 133.995 ;
        RECT 38.735 133.445 39.065 133.825 ;
        RECT 39.235 133.705 39.420 135.825 ;
        RECT 39.660 135.535 39.925 135.995 ;
        RECT 40.095 135.400 40.345 135.825 ;
        RECT 40.555 135.550 41.660 135.720 ;
        RECT 40.040 135.270 40.345 135.400 ;
        RECT 39.590 134.075 39.870 135.025 ;
        RECT 40.040 134.165 40.210 135.270 ;
        RECT 40.380 134.485 40.620 135.080 ;
        RECT 40.790 135.015 41.320 135.380 ;
        RECT 40.790 134.315 40.960 135.015 ;
        RECT 41.490 134.935 41.660 135.550 ;
        RECT 41.830 135.195 42.000 135.995 ;
        RECT 42.170 135.495 42.420 135.825 ;
        RECT 42.645 135.525 43.530 135.695 ;
        RECT 41.490 134.845 42.000 134.935 ;
        RECT 40.040 134.035 40.265 134.165 ;
        RECT 40.435 134.095 40.960 134.315 ;
        RECT 41.130 134.675 42.000 134.845 ;
        RECT 39.675 133.445 39.925 133.905 ;
        RECT 40.095 133.895 40.265 134.035 ;
        RECT 41.130 133.895 41.300 134.675 ;
        RECT 41.830 134.605 42.000 134.675 ;
        RECT 41.510 134.425 41.710 134.455 ;
        RECT 42.170 134.425 42.340 135.495 ;
        RECT 42.510 134.605 42.700 135.325 ;
        RECT 41.510 134.125 42.340 134.425 ;
        RECT 42.870 134.395 43.190 135.355 ;
        RECT 40.095 133.725 40.430 133.895 ;
        RECT 40.625 133.725 41.300 133.895 ;
        RECT 41.620 133.445 41.990 133.945 ;
        RECT 42.170 133.895 42.340 134.125 ;
        RECT 42.725 134.065 43.190 134.395 ;
        RECT 43.360 134.685 43.530 135.525 ;
        RECT 43.710 135.495 44.025 135.995 ;
        RECT 44.255 135.265 44.595 135.825 ;
        RECT 43.700 134.890 44.595 135.265 ;
        RECT 44.765 134.985 44.935 135.995 ;
        RECT 44.405 134.685 44.595 134.890 ;
        RECT 45.105 134.935 45.435 135.780 ;
        RECT 45.665 135.560 51.010 135.995 ;
        RECT 45.105 134.855 45.495 134.935 ;
        RECT 45.280 134.805 45.495 134.855 ;
        RECT 43.360 134.355 44.235 134.685 ;
        RECT 44.405 134.355 45.155 134.685 ;
        RECT 43.360 133.895 43.530 134.355 ;
        RECT 44.405 134.185 44.605 134.355 ;
        RECT 45.325 134.225 45.495 134.805 ;
        RECT 45.270 134.185 45.495 134.225 ;
        RECT 42.170 133.725 42.575 133.895 ;
        RECT 42.745 133.725 43.530 133.895 ;
        RECT 43.805 133.445 44.015 133.975 ;
        RECT 44.275 133.660 44.605 134.185 ;
        RECT 45.115 134.100 45.495 134.185 ;
        RECT 44.775 133.445 44.945 134.055 ;
        RECT 45.115 133.665 45.445 134.100 ;
        RECT 47.250 133.990 47.590 134.820 ;
        RECT 49.070 134.310 49.420 135.560 ;
        RECT 52.105 134.830 52.395 135.995 ;
        RECT 52.570 135.570 52.905 135.995 ;
        RECT 53.075 135.390 53.260 135.795 ;
        RECT 52.595 135.215 53.260 135.390 ;
        RECT 53.465 135.215 53.795 135.995 ;
        RECT 52.595 134.185 52.935 135.215 ;
        RECT 53.965 135.025 54.235 135.795 ;
        RECT 53.105 134.855 54.235 135.025 ;
        RECT 54.405 134.905 57.915 135.995 ;
        RECT 58.170 135.375 58.345 135.825 ;
        RECT 58.515 135.555 58.845 135.995 ;
        RECT 59.150 135.405 59.320 135.825 ;
        RECT 59.555 135.585 60.225 135.995 ;
        RECT 60.440 135.405 60.610 135.825 ;
        RECT 60.810 135.585 61.140 135.995 ;
        RECT 58.170 135.205 58.800 135.375 ;
        RECT 53.105 134.355 53.355 134.855 ;
        RECT 45.665 133.445 51.010 133.990 ;
        RECT 52.105 133.445 52.395 134.170 ;
        RECT 52.595 134.015 53.280 134.185 ;
        RECT 53.535 134.105 53.895 134.685 ;
        RECT 52.570 133.445 52.905 133.845 ;
        RECT 53.075 133.615 53.280 134.015 ;
        RECT 54.065 133.945 54.235 134.855 ;
        RECT 53.490 133.445 53.765 133.925 ;
        RECT 53.975 133.615 54.235 133.945 ;
        RECT 54.405 134.215 56.055 134.735 ;
        RECT 56.225 134.385 57.915 134.905 ;
        RECT 58.085 134.355 58.450 135.035 ;
        RECT 58.630 134.685 58.800 135.205 ;
        RECT 59.150 135.235 61.165 135.405 ;
        RECT 58.630 134.355 58.980 134.685 ;
        RECT 54.405 133.445 57.915 134.215 ;
        RECT 58.630 134.185 58.800 134.355 ;
        RECT 58.170 134.015 58.800 134.185 ;
        RECT 58.170 133.615 58.345 134.015 ;
        RECT 59.150 133.945 59.320 135.235 ;
        RECT 58.515 133.445 58.845 133.825 ;
        RECT 59.090 133.615 59.320 133.945 ;
        RECT 59.520 133.780 59.800 135.055 ;
        RECT 60.025 134.975 60.295 135.055 ;
        RECT 59.985 134.805 60.295 134.975 ;
        RECT 60.025 133.780 60.295 134.805 ;
        RECT 60.485 134.025 60.825 135.055 ;
        RECT 60.995 134.685 61.165 135.235 ;
        RECT 61.335 134.855 61.595 135.825 ;
        RECT 61.775 134.855 62.105 135.995 ;
        RECT 62.635 135.025 62.965 135.810 ;
        RECT 62.285 134.855 62.965 135.025 ;
        RECT 63.615 134.855 63.945 135.995 ;
        RECT 64.475 135.025 64.805 135.810 ;
        RECT 64.125 134.855 64.805 135.025 ;
        RECT 65.905 135.125 66.180 135.825 ;
        RECT 66.350 135.450 66.605 135.995 ;
        RECT 66.775 135.485 67.255 135.825 ;
        RECT 67.430 135.440 68.035 135.995 ;
        RECT 67.420 135.340 68.035 135.440 ;
        RECT 67.420 135.315 67.605 135.340 ;
        RECT 60.995 134.355 61.255 134.685 ;
        RECT 61.425 134.165 61.595 134.855 ;
        RECT 61.765 134.435 62.115 134.685 ;
        RECT 62.285 134.255 62.455 134.855 ;
        RECT 62.625 134.435 62.975 134.685 ;
        RECT 63.605 134.435 63.955 134.685 ;
        RECT 64.125 134.255 64.295 134.855 ;
        RECT 64.465 134.435 64.815 134.685 ;
        RECT 60.755 133.445 61.085 133.825 ;
        RECT 61.255 133.700 61.595 134.165 ;
        RECT 61.255 133.655 61.590 133.700 ;
        RECT 61.775 133.445 62.045 134.255 ;
        RECT 62.215 133.615 62.545 134.255 ;
        RECT 62.715 133.445 62.955 134.255 ;
        RECT 63.615 133.445 63.885 134.255 ;
        RECT 64.055 133.615 64.385 134.255 ;
        RECT 64.555 133.445 64.795 134.255 ;
        RECT 65.905 134.095 66.075 135.125 ;
        RECT 66.350 134.995 67.105 135.245 ;
        RECT 67.275 135.070 67.605 135.315 ;
        RECT 66.350 134.960 67.120 134.995 ;
        RECT 66.350 134.950 67.135 134.960 ;
        RECT 66.245 134.935 67.140 134.950 ;
        RECT 66.245 134.920 67.160 134.935 ;
        RECT 66.245 134.910 67.180 134.920 ;
        RECT 66.245 134.900 67.205 134.910 ;
        RECT 66.245 134.870 67.275 134.900 ;
        RECT 66.245 134.840 67.295 134.870 ;
        RECT 66.245 134.810 67.315 134.840 ;
        RECT 66.245 134.785 67.345 134.810 ;
        RECT 66.245 134.750 67.380 134.785 ;
        RECT 66.245 134.745 67.410 134.750 ;
        RECT 66.245 134.350 66.475 134.745 ;
        RECT 67.020 134.740 67.410 134.745 ;
        RECT 67.045 134.730 67.410 134.740 ;
        RECT 67.060 134.725 67.410 134.730 ;
        RECT 67.075 134.720 67.410 134.725 ;
        RECT 67.775 134.720 68.035 135.170 ;
        RECT 68.215 135.045 68.490 135.815 ;
        RECT 68.660 135.385 68.990 135.815 ;
        RECT 69.160 135.555 69.355 135.995 ;
        RECT 69.535 135.385 69.865 135.815 ;
        RECT 68.660 135.215 69.865 135.385 ;
        RECT 68.215 134.855 68.800 135.045 ;
        RECT 68.970 134.885 69.865 135.215 ;
        RECT 70.965 135.145 71.345 135.825 ;
        RECT 71.935 135.145 72.105 135.995 ;
        RECT 72.275 135.315 72.605 135.825 ;
        RECT 72.775 135.485 72.945 135.995 ;
        RECT 73.115 135.315 73.515 135.825 ;
        RECT 72.275 135.145 73.515 135.315 ;
        RECT 67.075 134.715 68.035 134.720 ;
        RECT 67.085 134.705 68.035 134.715 ;
        RECT 67.095 134.700 68.035 134.705 ;
        RECT 67.105 134.690 68.035 134.700 ;
        RECT 67.110 134.680 68.035 134.690 ;
        RECT 67.115 134.675 68.035 134.680 ;
        RECT 67.125 134.660 68.035 134.675 ;
        RECT 67.130 134.645 68.035 134.660 ;
        RECT 67.140 134.620 68.035 134.645 ;
        RECT 66.645 134.150 66.975 134.575 ;
        RECT 65.905 133.615 66.165 134.095 ;
        RECT 66.335 133.445 66.585 133.985 ;
        RECT 66.755 133.665 66.975 134.150 ;
        RECT 67.145 134.550 68.035 134.620 ;
        RECT 67.145 133.825 67.315 134.550 ;
        RECT 67.485 133.995 68.035 134.380 ;
        RECT 68.215 134.035 68.455 134.685 ;
        RECT 68.625 134.185 68.800 134.855 ;
        RECT 68.970 134.355 69.385 134.685 ;
        RECT 69.565 134.355 69.860 134.685 ;
        RECT 68.625 134.005 68.955 134.185 ;
        RECT 67.145 133.655 68.035 133.825 ;
        RECT 68.230 133.445 68.560 133.835 ;
        RECT 68.730 133.625 68.955 134.005 ;
        RECT 69.155 133.735 69.385 134.355 ;
        RECT 70.965 134.185 71.135 135.145 ;
        RECT 71.305 134.805 72.610 134.975 ;
        RECT 73.695 134.895 74.015 135.825 ;
        RECT 74.185 134.905 77.695 135.995 ;
        RECT 71.305 134.355 71.550 134.805 ;
        RECT 71.720 134.435 72.270 134.635 ;
        RECT 72.440 134.605 72.610 134.805 ;
        RECT 73.385 134.725 74.015 134.895 ;
        RECT 72.440 134.435 72.815 134.605 ;
        RECT 72.985 134.185 73.215 134.685 ;
        RECT 69.565 133.445 69.865 134.175 ;
        RECT 70.965 134.015 73.215 134.185 ;
        RECT 71.015 133.445 71.345 133.835 ;
        RECT 71.515 133.695 71.685 134.015 ;
        RECT 73.385 133.845 73.555 134.725 ;
        RECT 71.855 133.445 72.185 133.835 ;
        RECT 72.600 133.675 73.555 133.845 ;
        RECT 73.725 133.445 74.015 134.280 ;
        RECT 74.185 134.215 75.835 134.735 ;
        RECT 76.005 134.385 77.695 134.905 ;
        RECT 77.865 134.830 78.155 135.995 ;
        RECT 78.325 135.560 83.670 135.995 ;
        RECT 83.845 135.560 89.190 135.995 ;
        RECT 74.185 133.445 77.695 134.215 ;
        RECT 77.865 133.445 78.155 134.170 ;
        RECT 79.910 133.990 80.250 134.820 ;
        RECT 81.730 134.310 82.080 135.560 ;
        RECT 85.430 133.990 85.770 134.820 ;
        RECT 87.250 134.310 87.600 135.560 ;
        RECT 89.365 134.905 90.575 135.995 ;
        RECT 89.365 134.195 89.885 134.735 ;
        RECT 90.055 134.365 90.575 134.905 ;
        RECT 90.745 134.905 91.955 135.995 ;
        RECT 100.130 135.430 102.050 136.700 ;
        RECT 103.560 136.690 104.120 136.700 ;
        RECT 103.790 135.600 104.120 136.690 ;
        RECT 104.490 136.220 105.530 136.390 ;
        RECT 104.490 135.780 105.530 135.950 ;
        RECT 105.700 135.920 105.870 136.250 ;
        RECT 103.950 135.380 104.120 135.600 ;
        RECT 106.210 135.380 106.380 136.790 ;
        RECT 103.950 135.210 106.380 135.380 ;
        RECT 107.960 137.300 118.590 137.470 ;
        RECT 120.020 146.580 126.250 146.740 ;
        RECT 120.020 144.320 120.690 146.580 ;
        RECT 121.360 146.010 125.400 146.180 ;
        RECT 121.020 144.950 121.190 145.950 ;
        RECT 125.570 144.950 125.740 145.950 ;
        RECT 121.360 144.720 125.400 144.890 ;
        RECT 126.080 144.320 126.250 146.580 ;
        RECT 120.020 144.150 126.250 144.320 ;
        RECT 120.020 140.890 120.690 144.150 ;
        RECT 121.360 143.580 125.400 143.750 ;
        RECT 121.020 141.520 121.190 143.520 ;
        RECT 125.570 141.520 125.740 143.520 ;
        RECT 121.360 141.290 125.400 141.460 ;
        RECT 126.080 140.890 126.250 144.150 ;
        RECT 120.020 140.720 126.250 140.890 ;
        RECT 120.020 137.460 120.690 140.720 ;
        RECT 121.360 140.150 125.400 140.320 ;
        RECT 121.020 138.090 121.190 140.090 ;
        RECT 125.570 138.090 125.740 140.090 ;
        RECT 121.360 137.860 125.400 138.030 ;
        RECT 126.080 137.460 126.250 140.720 ;
        RECT 120.020 137.450 126.250 137.460 ;
        RECT 127.840 146.720 137.670 146.760 ;
        RECT 140.540 146.740 146.280 146.750 ;
        RECT 127.840 146.590 138.470 146.720 ;
        RECT 127.840 144.330 128.010 146.590 ;
        RECT 128.735 146.020 136.775 146.190 ;
        RECT 128.350 144.960 128.520 145.960 ;
        RECT 136.990 144.960 137.160 145.960 ;
        RECT 128.735 144.730 136.775 144.900 ;
        RECT 137.500 144.330 138.470 146.590 ;
        RECT 127.840 144.160 138.470 144.330 ;
        RECT 127.840 140.900 128.010 144.160 ;
        RECT 128.735 143.590 136.775 143.760 ;
        RECT 128.350 141.530 128.520 143.530 ;
        RECT 136.990 141.530 137.160 143.530 ;
        RECT 128.735 141.300 136.775 141.470 ;
        RECT 137.500 140.900 138.470 144.160 ;
        RECT 127.840 140.730 138.470 140.900 ;
        RECT 127.840 137.470 128.010 140.730 ;
        RECT 128.735 140.160 136.775 140.330 ;
        RECT 128.350 138.100 128.520 140.100 ;
        RECT 136.990 138.100 137.160 140.100 ;
        RECT 128.735 137.870 136.775 138.040 ;
        RECT 137.500 137.470 138.470 140.730 ;
        RECT 120.020 137.350 126.260 137.450 ;
        RECT 107.960 135.040 108.130 137.300 ;
        RECT 108.855 136.730 116.895 136.900 ;
        RECT 108.470 135.670 108.640 136.670 ;
        RECT 117.110 135.670 117.280 136.670 ;
        RECT 108.855 135.440 116.895 135.610 ;
        RECT 117.620 135.040 118.590 137.300 ;
        RECT 120.010 136.790 126.260 137.350 ;
        RECT 120.010 136.770 125.180 136.790 ;
        RECT 120.010 136.700 124.000 136.770 ;
        RECT 120.010 135.430 121.930 136.700 ;
        RECT 123.440 136.690 124.000 136.700 ;
        RECT 123.670 135.600 124.000 136.690 ;
        RECT 124.370 136.220 125.410 136.390 ;
        RECT 124.370 135.780 125.410 135.950 ;
        RECT 125.580 135.920 125.750 136.250 ;
        RECT 123.830 135.380 124.000 135.600 ;
        RECT 126.090 135.380 126.260 136.790 ;
        RECT 123.830 135.210 126.260 135.380 ;
        RECT 127.840 137.300 138.470 137.470 ;
        RECT 140.050 146.580 146.280 146.740 ;
        RECT 140.050 144.320 140.720 146.580 ;
        RECT 141.390 146.010 145.430 146.180 ;
        RECT 141.050 144.950 141.220 145.950 ;
        RECT 145.600 144.950 145.770 145.950 ;
        RECT 141.390 144.720 145.430 144.890 ;
        RECT 146.110 144.320 146.280 146.580 ;
        RECT 140.050 144.150 146.280 144.320 ;
        RECT 140.050 140.890 140.720 144.150 ;
        RECT 141.390 143.580 145.430 143.750 ;
        RECT 141.050 141.520 141.220 143.520 ;
        RECT 145.600 141.520 145.770 143.520 ;
        RECT 141.390 141.290 145.430 141.460 ;
        RECT 146.110 140.890 146.280 144.150 ;
        RECT 140.050 140.720 146.280 140.890 ;
        RECT 140.050 137.460 140.720 140.720 ;
        RECT 141.390 140.150 145.430 140.320 ;
        RECT 141.050 138.090 141.220 140.090 ;
        RECT 145.600 138.090 145.770 140.090 ;
        RECT 141.390 137.860 145.430 138.030 ;
        RECT 146.110 137.460 146.280 140.720 ;
        RECT 140.050 137.450 146.280 137.460 ;
        RECT 147.870 146.720 157.700 146.760 ;
        RECT 147.870 146.590 158.500 146.720 ;
        RECT 147.870 144.330 148.040 146.590 ;
        RECT 148.765 146.020 156.805 146.190 ;
        RECT 148.380 144.960 148.550 145.960 ;
        RECT 157.020 144.960 157.190 145.960 ;
        RECT 148.765 144.730 156.805 144.900 ;
        RECT 157.530 144.330 158.500 146.590 ;
        RECT 147.870 144.160 158.500 144.330 ;
        RECT 147.870 140.900 148.040 144.160 ;
        RECT 148.765 143.590 156.805 143.760 ;
        RECT 148.380 141.530 148.550 143.530 ;
        RECT 157.020 141.530 157.190 143.530 ;
        RECT 148.765 141.300 156.805 141.470 ;
        RECT 157.530 140.900 158.500 144.160 ;
        RECT 147.870 140.730 158.500 140.900 ;
        RECT 147.870 137.470 148.040 140.730 ;
        RECT 148.765 140.160 156.805 140.330 ;
        RECT 148.380 138.100 148.550 140.100 ;
        RECT 157.020 138.100 157.190 140.100 ;
        RECT 148.765 137.870 156.805 138.040 ;
        RECT 157.530 137.470 158.500 140.730 ;
        RECT 140.050 137.350 146.290 137.450 ;
        RECT 107.960 135.010 118.590 135.040 ;
        RECT 127.840 135.040 128.010 137.300 ;
        RECT 128.735 136.730 136.775 136.900 ;
        RECT 128.350 135.670 128.520 136.670 ;
        RECT 136.990 135.670 137.160 136.670 ;
        RECT 128.735 135.440 136.775 135.610 ;
        RECT 137.500 135.040 138.470 137.300 ;
        RECT 140.040 136.790 146.290 137.350 ;
        RECT 140.040 136.770 145.210 136.790 ;
        RECT 140.040 136.700 144.030 136.770 ;
        RECT 140.040 135.430 141.960 136.700 ;
        RECT 143.470 136.690 144.030 136.700 ;
        RECT 143.700 135.600 144.030 136.690 ;
        RECT 144.400 136.220 145.440 136.390 ;
        RECT 144.400 135.780 145.440 135.950 ;
        RECT 145.610 135.920 145.780 136.250 ;
        RECT 143.860 135.380 144.030 135.600 ;
        RECT 146.120 135.380 146.290 136.790 ;
        RECT 143.860 135.210 146.290 135.380 ;
        RECT 147.870 137.300 158.500 137.470 ;
        RECT 127.840 135.010 138.470 135.040 ;
        RECT 147.870 135.040 148.040 137.300 ;
        RECT 148.765 136.730 156.805 136.900 ;
        RECT 148.380 135.670 148.550 136.670 ;
        RECT 157.020 135.670 157.190 136.670 ;
        RECT 148.765 135.440 156.805 135.610 ;
        RECT 157.530 135.040 158.500 137.300 ;
        RECT 147.870 135.010 158.500 135.040 ;
        RECT 90.745 134.365 91.265 134.905 ;
        RECT 107.930 134.900 118.590 135.010 ;
        RECT 127.810 134.900 138.470 135.010 ;
        RECT 147.840 134.900 158.500 135.010 ;
        RECT 106.180 134.850 118.590 134.900 ;
        RECT 126.060 134.850 138.470 134.900 ;
        RECT 146.090 134.850 158.500 134.900 ;
        RECT 91.435 134.195 91.955 134.735 ;
        RECT 78.325 133.445 83.670 133.990 ;
        RECT 83.845 133.445 89.190 133.990 ;
        RECT 89.365 133.445 90.575 134.195 ;
        RECT 90.745 133.445 91.955 134.195 ;
        RECT 101.840 134.680 118.590 134.850 ;
        RECT 13.380 133.275 92.040 133.445 ;
        RECT 13.465 132.525 14.675 133.275 ;
        RECT 14.845 132.730 20.190 133.275 ;
        RECT 20.365 132.730 25.710 133.275 ;
        RECT 13.465 131.985 13.985 132.525 ;
        RECT 14.155 131.815 14.675 132.355 ;
        RECT 16.430 131.900 16.770 132.730 ;
        RECT 13.465 130.725 14.675 131.815 ;
        RECT 18.250 131.160 18.600 132.410 ;
        RECT 21.950 131.900 22.290 132.730 ;
        RECT 25.885 132.525 27.095 133.275 ;
        RECT 27.265 132.625 27.525 133.105 ;
        RECT 27.695 132.815 28.025 133.275 ;
        RECT 28.215 132.635 28.415 133.055 ;
        RECT 23.770 131.160 24.120 132.410 ;
        RECT 25.885 131.985 26.405 132.525 ;
        RECT 26.575 131.815 27.095 132.355 ;
        RECT 14.845 130.725 20.190 131.160 ;
        RECT 20.365 130.725 25.710 131.160 ;
        RECT 25.885 130.725 27.095 131.815 ;
        RECT 27.265 131.595 27.435 132.625 ;
        RECT 27.605 131.935 27.835 132.365 ;
        RECT 28.005 132.115 28.415 132.635 ;
        RECT 28.585 132.790 29.375 133.055 ;
        RECT 28.585 131.935 28.840 132.790 ;
        RECT 29.555 132.455 29.885 132.875 ;
        RECT 30.055 132.455 30.315 133.275 ;
        RECT 31.060 132.645 31.345 133.105 ;
        RECT 31.515 132.815 31.785 133.275 ;
        RECT 31.060 132.475 32.015 132.645 ;
        RECT 29.555 132.365 29.805 132.455 ;
        RECT 29.010 132.115 29.805 132.365 ;
        RECT 27.605 131.765 29.395 131.935 ;
        RECT 27.265 130.895 27.540 131.595 ;
        RECT 27.710 131.470 28.425 131.765 ;
        RECT 28.645 131.405 28.975 131.595 ;
        RECT 27.750 130.725 27.965 131.270 ;
        RECT 28.135 130.895 28.610 131.235 ;
        RECT 28.780 131.230 28.975 131.405 ;
        RECT 29.145 131.400 29.395 131.765 ;
        RECT 28.780 130.725 29.395 131.230 ;
        RECT 29.635 130.895 29.805 132.115 ;
        RECT 29.975 131.405 30.315 132.285 ;
        RECT 30.945 131.745 31.635 132.305 ;
        RECT 31.805 131.575 32.015 132.475 ;
        RECT 31.060 131.355 32.015 131.575 ;
        RECT 32.185 132.305 32.585 133.105 ;
        RECT 32.775 132.645 33.055 133.105 ;
        RECT 33.575 132.815 33.900 133.275 ;
        RECT 32.775 132.475 33.900 132.645 ;
        RECT 34.070 132.535 34.455 133.105 ;
        RECT 33.450 132.365 33.900 132.475 ;
        RECT 32.185 131.745 33.280 132.305 ;
        RECT 33.450 132.035 34.005 132.365 ;
        RECT 30.055 130.725 30.315 131.235 ;
        RECT 31.060 130.895 31.345 131.355 ;
        RECT 31.515 130.725 31.785 131.185 ;
        RECT 32.185 130.895 32.585 131.745 ;
        RECT 33.450 131.575 33.900 132.035 ;
        RECT 34.175 131.865 34.455 132.535 ;
        RECT 35.660 132.645 35.945 133.105 ;
        RECT 36.115 132.815 36.385 133.275 ;
        RECT 35.660 132.475 36.615 132.645 ;
        RECT 32.775 131.355 33.900 131.575 ;
        RECT 32.775 130.895 33.055 131.355 ;
        RECT 33.575 130.725 33.900 131.185 ;
        RECT 34.070 130.895 34.455 131.865 ;
        RECT 35.545 131.745 36.235 132.305 ;
        RECT 36.405 131.575 36.615 132.475 ;
        RECT 35.660 131.355 36.615 131.575 ;
        RECT 36.785 132.305 37.185 133.105 ;
        RECT 37.375 132.645 37.655 133.105 ;
        RECT 38.175 132.815 38.500 133.275 ;
        RECT 37.375 132.475 38.500 132.645 ;
        RECT 38.670 132.535 39.055 133.105 ;
        RECT 39.225 132.550 39.515 133.275 ;
        RECT 39.710 132.885 40.040 133.275 ;
        RECT 40.210 132.715 40.435 133.095 ;
        RECT 38.050 132.365 38.500 132.475 ;
        RECT 36.785 131.745 37.880 132.305 ;
        RECT 38.050 132.035 38.605 132.365 ;
        RECT 35.660 130.895 35.945 131.355 ;
        RECT 36.115 130.725 36.385 131.185 ;
        RECT 36.785 130.895 37.185 131.745 ;
        RECT 38.050 131.575 38.500 132.035 ;
        RECT 38.775 131.865 39.055 132.535 ;
        RECT 39.695 132.035 39.935 132.685 ;
        RECT 40.105 132.535 40.435 132.715 ;
        RECT 37.375 131.355 38.500 131.575 ;
        RECT 37.375 130.895 37.655 131.355 ;
        RECT 38.175 130.725 38.500 131.185 ;
        RECT 38.670 130.895 39.055 131.865 ;
        RECT 39.225 130.725 39.515 131.890 ;
        RECT 40.105 131.865 40.280 132.535 ;
        RECT 40.635 132.365 40.865 132.985 ;
        RECT 41.045 132.545 41.345 133.275 ;
        RECT 41.525 132.525 42.735 133.275 ;
        RECT 42.905 132.535 43.290 133.105 ;
        RECT 43.460 132.815 43.785 133.275 ;
        RECT 44.305 132.645 44.585 133.105 ;
        RECT 40.450 132.035 40.865 132.365 ;
        RECT 41.045 132.035 41.340 132.365 ;
        RECT 41.525 131.985 42.045 132.525 ;
        RECT 39.695 131.675 40.280 131.865 ;
        RECT 39.695 130.905 39.970 131.675 ;
        RECT 40.450 131.505 41.345 131.835 ;
        RECT 42.215 131.815 42.735 132.355 ;
        RECT 40.140 131.335 41.345 131.505 ;
        RECT 40.140 130.905 40.470 131.335 ;
        RECT 40.640 130.725 40.835 131.165 ;
        RECT 41.015 130.905 41.345 131.335 ;
        RECT 41.525 130.725 42.735 131.815 ;
        RECT 42.905 131.865 43.185 132.535 ;
        RECT 43.460 132.475 44.585 132.645 ;
        RECT 43.460 132.365 43.910 132.475 ;
        RECT 43.355 132.035 43.910 132.365 ;
        RECT 44.775 132.305 45.175 133.105 ;
        RECT 45.575 132.815 45.845 133.275 ;
        RECT 46.015 132.645 46.300 133.105 ;
        RECT 42.905 130.895 43.290 131.865 ;
        RECT 43.460 131.575 43.910 132.035 ;
        RECT 44.080 131.745 45.175 132.305 ;
        RECT 43.460 131.355 44.585 131.575 ;
        RECT 43.460 130.725 43.785 131.185 ;
        RECT 44.305 130.895 44.585 131.355 ;
        RECT 44.775 130.895 45.175 131.745 ;
        RECT 45.345 132.475 46.300 132.645 ;
        RECT 46.585 132.475 47.280 133.105 ;
        RECT 47.485 132.475 47.795 133.275 ;
        RECT 48.935 132.885 49.265 133.275 ;
        RECT 49.435 132.705 49.605 133.025 ;
        RECT 49.775 132.885 50.105 133.275 ;
        RECT 50.520 132.875 51.475 133.045 ;
        RECT 48.885 132.535 51.135 132.705 ;
        RECT 45.345 131.575 45.555 132.475 ;
        RECT 45.725 131.745 46.415 132.305 ;
        RECT 46.605 132.035 46.940 132.285 ;
        RECT 47.110 131.875 47.280 132.475 ;
        RECT 47.450 132.035 47.785 132.305 ;
        RECT 45.345 131.355 46.300 131.575 ;
        RECT 45.575 130.725 45.845 131.185 ;
        RECT 46.015 130.895 46.300 131.355 ;
        RECT 46.585 130.725 46.845 131.865 ;
        RECT 47.015 130.895 47.345 131.875 ;
        RECT 47.515 130.725 47.795 131.865 ;
        RECT 48.885 131.575 49.055 132.535 ;
        RECT 49.225 131.915 49.470 132.365 ;
        RECT 49.640 132.085 50.190 132.285 ;
        RECT 50.360 132.115 50.735 132.285 ;
        RECT 50.360 131.915 50.530 132.115 ;
        RECT 50.905 132.035 51.135 132.535 ;
        RECT 49.225 131.745 50.530 131.915 ;
        RECT 51.305 131.995 51.475 132.875 ;
        RECT 51.645 132.440 51.935 133.275 ;
        RECT 52.190 132.705 52.365 133.105 ;
        RECT 52.535 132.895 52.865 133.275 ;
        RECT 53.110 132.775 53.340 133.105 ;
        RECT 52.190 132.535 52.820 132.705 ;
        RECT 52.650 132.365 52.820 132.535 ;
        RECT 51.305 131.825 51.935 131.995 ;
        RECT 48.885 130.895 49.265 131.575 ;
        RECT 49.855 130.725 50.025 131.575 ;
        RECT 50.195 131.405 51.435 131.575 ;
        RECT 50.195 130.895 50.525 131.405 ;
        RECT 50.695 130.725 50.865 131.235 ;
        RECT 51.035 130.895 51.435 131.405 ;
        RECT 51.615 130.895 51.935 131.825 ;
        RECT 52.105 131.685 52.470 132.365 ;
        RECT 52.650 132.035 53.000 132.365 ;
        RECT 52.650 131.515 52.820 132.035 ;
        RECT 52.190 131.345 52.820 131.515 ;
        RECT 53.170 131.485 53.340 132.775 ;
        RECT 53.540 131.665 53.820 132.940 ;
        RECT 54.045 132.935 54.315 132.940 ;
        RECT 54.005 132.765 54.315 132.935 ;
        RECT 54.775 132.895 55.105 133.275 ;
        RECT 55.275 133.020 55.610 133.065 ;
        RECT 54.045 131.665 54.315 132.765 ;
        RECT 54.505 131.665 54.845 132.695 ;
        RECT 55.275 132.555 55.615 133.020 ;
        RECT 55.015 132.035 55.275 132.365 ;
        RECT 55.015 131.485 55.185 132.035 ;
        RECT 55.445 131.865 55.615 132.555 ;
        RECT 55.785 132.505 57.455 133.275 ;
        RECT 57.715 132.725 57.885 133.015 ;
        RECT 58.055 132.895 58.385 133.275 ;
        RECT 57.715 132.555 58.380 132.725 ;
        RECT 55.785 131.985 56.535 132.505 ;
        RECT 52.190 130.895 52.365 131.345 ;
        RECT 53.170 131.315 55.185 131.485 ;
        RECT 52.535 130.725 52.865 131.165 ;
        RECT 53.170 130.895 53.340 131.315 ;
        RECT 53.575 130.725 54.245 131.135 ;
        RECT 54.460 130.895 54.630 131.315 ;
        RECT 54.830 130.725 55.160 131.135 ;
        RECT 55.355 130.895 55.615 131.865 ;
        RECT 56.705 131.815 57.455 132.335 ;
        RECT 55.785 130.725 57.455 131.815 ;
        RECT 57.630 131.735 57.980 132.385 ;
        RECT 58.150 131.565 58.380 132.555 ;
        RECT 57.715 131.395 58.380 131.565 ;
        RECT 57.715 130.895 57.885 131.395 ;
        RECT 58.055 130.725 58.385 131.225 ;
        RECT 58.555 130.895 58.740 133.015 ;
        RECT 58.995 132.815 59.245 133.275 ;
        RECT 59.415 132.825 59.750 132.995 ;
        RECT 59.945 132.825 60.620 132.995 ;
        RECT 59.415 132.685 59.585 132.825 ;
        RECT 58.910 131.695 59.190 132.645 ;
        RECT 59.360 132.555 59.585 132.685 ;
        RECT 59.360 131.450 59.530 132.555 ;
        RECT 59.755 132.405 60.280 132.625 ;
        RECT 59.700 131.640 59.940 132.235 ;
        RECT 60.110 131.705 60.280 132.405 ;
        RECT 60.450 132.045 60.620 132.825 ;
        RECT 60.940 132.775 61.310 133.275 ;
        RECT 61.490 132.825 61.895 132.995 ;
        RECT 62.065 132.825 62.850 132.995 ;
        RECT 61.490 132.595 61.660 132.825 ;
        RECT 60.830 132.295 61.660 132.595 ;
        RECT 62.045 132.325 62.510 132.655 ;
        RECT 60.830 132.265 61.030 132.295 ;
        RECT 61.150 132.045 61.320 132.115 ;
        RECT 60.450 131.875 61.320 132.045 ;
        RECT 60.810 131.785 61.320 131.875 ;
        RECT 59.360 131.320 59.665 131.450 ;
        RECT 60.110 131.340 60.640 131.705 ;
        RECT 58.980 130.725 59.245 131.185 ;
        RECT 59.415 130.895 59.665 131.320 ;
        RECT 60.810 131.170 60.980 131.785 ;
        RECT 59.875 131.000 60.980 131.170 ;
        RECT 61.150 130.725 61.320 131.525 ;
        RECT 61.490 131.225 61.660 132.295 ;
        RECT 61.830 131.395 62.020 132.115 ;
        RECT 62.190 131.365 62.510 132.325 ;
        RECT 62.680 132.365 62.850 132.825 ;
        RECT 63.125 132.745 63.335 133.275 ;
        RECT 63.595 132.535 63.925 133.060 ;
        RECT 64.095 132.665 64.265 133.275 ;
        RECT 64.435 132.620 64.765 133.055 ;
        RECT 64.435 132.535 64.815 132.620 ;
        RECT 64.985 132.550 65.275 133.275 ;
        RECT 66.455 132.725 66.625 133.015 ;
        RECT 66.795 132.895 67.125 133.275 ;
        RECT 66.455 132.555 67.120 132.725 ;
        RECT 63.725 132.365 63.925 132.535 ;
        RECT 64.590 132.495 64.815 132.535 ;
        RECT 62.680 132.035 63.555 132.365 ;
        RECT 63.725 132.035 64.475 132.365 ;
        RECT 61.490 130.895 61.740 131.225 ;
        RECT 62.680 131.195 62.850 132.035 ;
        RECT 63.725 131.830 63.915 132.035 ;
        RECT 64.645 131.915 64.815 132.495 ;
        RECT 64.600 131.865 64.815 131.915 ;
        RECT 63.020 131.455 63.915 131.830 ;
        RECT 64.425 131.785 64.815 131.865 ;
        RECT 61.965 131.025 62.850 131.195 ;
        RECT 63.030 130.725 63.345 131.225 ;
        RECT 63.575 130.895 63.915 131.455 ;
        RECT 64.085 130.725 64.255 131.735 ;
        RECT 64.425 130.940 64.755 131.785 ;
        RECT 64.985 130.725 65.275 131.890 ;
        RECT 66.370 131.735 66.720 132.385 ;
        RECT 66.890 131.565 67.120 132.555 ;
        RECT 66.455 131.395 67.120 131.565 ;
        RECT 66.455 130.895 66.625 131.395 ;
        RECT 66.795 130.725 67.125 131.225 ;
        RECT 67.295 130.895 67.480 133.015 ;
        RECT 67.735 132.815 67.985 133.275 ;
        RECT 68.155 132.825 68.490 132.995 ;
        RECT 68.685 132.825 69.360 132.995 ;
        RECT 68.155 132.685 68.325 132.825 ;
        RECT 67.650 131.695 67.930 132.645 ;
        RECT 68.100 132.555 68.325 132.685 ;
        RECT 68.100 131.450 68.270 132.555 ;
        RECT 68.495 132.405 69.020 132.625 ;
        RECT 68.440 131.640 68.680 132.235 ;
        RECT 68.850 131.705 69.020 132.405 ;
        RECT 69.190 132.045 69.360 132.825 ;
        RECT 69.680 132.775 70.050 133.275 ;
        RECT 70.230 132.825 70.635 132.995 ;
        RECT 70.805 132.825 71.590 132.995 ;
        RECT 70.230 132.595 70.400 132.825 ;
        RECT 69.570 132.295 70.400 132.595 ;
        RECT 70.785 132.325 71.250 132.655 ;
        RECT 69.570 132.265 69.770 132.295 ;
        RECT 69.890 132.045 70.060 132.115 ;
        RECT 69.190 131.875 70.060 132.045 ;
        RECT 69.550 131.785 70.060 131.875 ;
        RECT 68.100 131.320 68.405 131.450 ;
        RECT 68.850 131.340 69.380 131.705 ;
        RECT 67.720 130.725 67.985 131.185 ;
        RECT 68.155 130.895 68.405 131.320 ;
        RECT 69.550 131.170 69.720 131.785 ;
        RECT 68.615 131.000 69.720 131.170 ;
        RECT 69.890 130.725 70.060 131.525 ;
        RECT 70.230 131.225 70.400 132.295 ;
        RECT 70.570 131.395 70.760 132.115 ;
        RECT 70.930 131.365 71.250 132.325 ;
        RECT 71.420 132.365 71.590 132.825 ;
        RECT 71.865 132.745 72.075 133.275 ;
        RECT 72.335 132.535 72.665 133.060 ;
        RECT 72.835 132.665 73.005 133.275 ;
        RECT 73.175 132.620 73.505 133.055 ;
        RECT 73.725 132.730 79.070 133.275 ;
        RECT 79.245 132.730 84.590 133.275 ;
        RECT 84.765 132.730 90.110 133.275 ;
        RECT 73.175 132.535 73.555 132.620 ;
        RECT 72.465 132.365 72.665 132.535 ;
        RECT 73.330 132.495 73.555 132.535 ;
        RECT 71.420 132.035 72.295 132.365 ;
        RECT 72.465 132.035 73.215 132.365 ;
        RECT 70.230 130.895 70.480 131.225 ;
        RECT 71.420 131.195 71.590 132.035 ;
        RECT 72.465 131.830 72.655 132.035 ;
        RECT 73.385 131.915 73.555 132.495 ;
        RECT 73.340 131.865 73.555 131.915 ;
        RECT 75.310 131.900 75.650 132.730 ;
        RECT 71.760 131.455 72.655 131.830 ;
        RECT 73.165 131.785 73.555 131.865 ;
        RECT 70.705 131.025 71.590 131.195 ;
        RECT 71.770 130.725 72.085 131.225 ;
        RECT 72.315 130.895 72.655 131.455 ;
        RECT 72.825 130.725 72.995 131.735 ;
        RECT 73.165 130.940 73.495 131.785 ;
        RECT 77.130 131.160 77.480 132.410 ;
        RECT 80.830 131.900 81.170 132.730 ;
        RECT 82.650 131.160 83.000 132.410 ;
        RECT 86.350 131.900 86.690 132.730 ;
        RECT 90.745 132.525 91.955 133.275 ;
        RECT 101.840 133.270 102.010 134.680 ;
        RECT 102.380 134.110 105.420 134.280 ;
        RECT 102.380 133.670 105.420 133.840 ;
        RECT 105.635 133.810 105.805 134.140 ;
        RECT 106.140 133.920 118.590 134.680 ;
        RECT 121.720 134.680 138.470 134.850 ;
        RECT 106.140 133.910 118.480 133.920 ;
        RECT 106.140 133.900 112.020 133.910 ;
        RECT 106.140 133.880 106.710 133.900 ;
        RECT 107.930 133.890 112.020 133.900 ;
        RECT 106.150 133.270 106.320 133.880 ;
        RECT 101.840 133.100 106.320 133.270 ;
        RECT 121.720 133.270 121.890 134.680 ;
        RECT 122.260 134.110 125.300 134.280 ;
        RECT 122.260 133.670 125.300 133.840 ;
        RECT 125.515 133.810 125.685 134.140 ;
        RECT 126.020 133.920 138.470 134.680 ;
        RECT 141.750 134.680 158.500 134.850 ;
        RECT 126.020 133.910 138.360 133.920 ;
        RECT 126.020 133.900 131.900 133.910 ;
        RECT 126.020 133.880 126.590 133.900 ;
        RECT 127.810 133.890 131.900 133.900 ;
        RECT 126.030 133.270 126.200 133.880 ;
        RECT 121.720 133.100 126.200 133.270 ;
        RECT 141.750 133.270 141.920 134.680 ;
        RECT 142.290 134.110 145.330 134.280 ;
        RECT 142.290 133.670 145.330 133.840 ;
        RECT 145.545 133.810 145.715 134.140 ;
        RECT 146.050 133.920 158.500 134.680 ;
        RECT 146.050 133.910 158.390 133.920 ;
        RECT 146.050 133.900 151.930 133.910 ;
        RECT 146.050 133.880 146.620 133.900 ;
        RECT 147.840 133.890 151.930 133.900 ;
        RECT 146.060 133.270 146.230 133.880 ;
        RECT 141.750 133.100 146.230 133.270 ;
        RECT 88.170 131.160 88.520 132.410 ;
        RECT 90.745 131.815 91.265 132.355 ;
        RECT 91.435 131.985 91.955 132.525 ;
        RECT 73.725 130.725 79.070 131.160 ;
        RECT 79.245 130.725 84.590 131.160 ;
        RECT 84.765 130.725 90.110 131.160 ;
        RECT 90.745 130.725 91.955 131.815 ;
        RECT 120.510 131.800 126.250 131.810 ;
        RECT 100.630 131.740 106.370 131.750 ;
        RECT 100.140 131.580 106.370 131.740 ;
        RECT 13.380 130.555 92.040 130.725 ;
        RECT 13.465 129.465 14.675 130.555 ;
        RECT 14.845 130.120 20.190 130.555 ;
        RECT 20.365 130.120 25.710 130.555 ;
        RECT 13.465 128.755 13.985 129.295 ;
        RECT 14.155 128.925 14.675 129.465 ;
        RECT 13.465 128.005 14.675 128.755 ;
        RECT 16.430 128.550 16.770 129.380 ;
        RECT 18.250 128.870 18.600 130.120 ;
        RECT 21.950 128.550 22.290 129.380 ;
        RECT 23.770 128.870 24.120 130.120 ;
        RECT 26.345 129.390 26.635 130.555 ;
        RECT 26.865 129.495 27.195 130.340 ;
        RECT 27.365 129.545 27.535 130.555 ;
        RECT 27.705 129.825 28.045 130.385 ;
        RECT 28.275 130.055 28.590 130.555 ;
        RECT 28.770 130.085 29.655 130.255 ;
        RECT 26.805 129.415 27.195 129.495 ;
        RECT 27.705 129.450 28.600 129.825 ;
        RECT 26.805 129.365 27.020 129.415 ;
        RECT 26.805 128.785 26.975 129.365 ;
        RECT 27.705 129.245 27.895 129.450 ;
        RECT 28.770 129.245 28.940 130.085 ;
        RECT 29.880 130.055 30.130 130.385 ;
        RECT 27.145 128.915 27.895 129.245 ;
        RECT 28.065 128.915 28.940 129.245 ;
        RECT 26.805 128.745 27.030 128.785 ;
        RECT 27.695 128.745 27.895 128.915 ;
        RECT 14.845 128.005 20.190 128.550 ;
        RECT 20.365 128.005 25.710 128.550 ;
        RECT 26.345 128.005 26.635 128.730 ;
        RECT 26.805 128.660 27.185 128.745 ;
        RECT 26.855 128.225 27.185 128.660 ;
        RECT 27.355 128.005 27.525 128.615 ;
        RECT 27.695 128.220 28.025 128.745 ;
        RECT 28.285 128.005 28.495 128.535 ;
        RECT 28.770 128.455 28.940 128.915 ;
        RECT 29.110 128.955 29.430 129.915 ;
        RECT 29.600 129.165 29.790 129.885 ;
        RECT 29.960 128.985 30.130 130.055 ;
        RECT 30.300 129.755 30.470 130.555 ;
        RECT 30.640 130.110 31.745 130.280 ;
        RECT 30.640 129.495 30.810 130.110 ;
        RECT 31.955 129.960 32.205 130.385 ;
        RECT 32.375 130.095 32.640 130.555 ;
        RECT 30.980 129.575 31.510 129.940 ;
        RECT 31.955 129.830 32.260 129.960 ;
        RECT 30.300 129.405 30.810 129.495 ;
        RECT 30.300 129.235 31.170 129.405 ;
        RECT 30.300 129.165 30.470 129.235 ;
        RECT 30.590 128.985 30.790 129.015 ;
        RECT 29.110 128.625 29.575 128.955 ;
        RECT 29.960 128.685 30.790 128.985 ;
        RECT 29.960 128.455 30.130 128.685 ;
        RECT 28.770 128.285 29.555 128.455 ;
        RECT 29.725 128.285 30.130 128.455 ;
        RECT 30.310 128.005 30.680 128.505 ;
        RECT 31.000 128.455 31.170 129.235 ;
        RECT 31.340 128.875 31.510 129.575 ;
        RECT 31.680 129.045 31.920 129.640 ;
        RECT 31.340 128.655 31.865 128.875 ;
        RECT 32.090 128.725 32.260 129.830 ;
        RECT 32.035 128.595 32.260 128.725 ;
        RECT 32.430 128.635 32.710 129.585 ;
        RECT 32.035 128.455 32.205 128.595 ;
        RECT 31.000 128.285 31.675 128.455 ;
        RECT 31.870 128.285 32.205 128.455 ;
        RECT 32.375 128.005 32.625 128.465 ;
        RECT 32.880 128.265 33.065 130.385 ;
        RECT 33.235 130.055 33.565 130.555 ;
        RECT 33.735 129.885 33.905 130.385 ;
        RECT 33.240 129.715 33.905 129.885 ;
        RECT 34.200 129.765 34.735 130.385 ;
        RECT 33.240 128.725 33.470 129.715 ;
        RECT 33.640 128.895 33.990 129.545 ;
        RECT 34.200 128.745 34.515 129.765 ;
        RECT 34.905 129.755 35.235 130.555 ;
        RECT 36.555 129.885 36.725 130.385 ;
        RECT 36.895 130.055 37.225 130.555 ;
        RECT 35.720 129.585 36.110 129.760 ;
        RECT 36.555 129.715 37.220 129.885 ;
        RECT 34.685 129.415 36.110 129.585 ;
        RECT 34.685 128.915 34.855 129.415 ;
        RECT 33.240 128.555 33.905 128.725 ;
        RECT 33.235 128.005 33.565 128.385 ;
        RECT 33.735 128.265 33.905 128.555 ;
        RECT 34.200 128.175 34.815 128.745 ;
        RECT 35.105 128.685 35.370 129.245 ;
        RECT 35.540 128.515 35.710 129.415 ;
        RECT 35.880 128.685 36.235 129.245 ;
        RECT 36.470 128.895 36.820 129.545 ;
        RECT 36.990 128.725 37.220 129.715 ;
        RECT 36.555 128.555 37.220 128.725 ;
        RECT 34.985 128.005 35.200 128.515 ;
        RECT 35.430 128.185 35.710 128.515 ;
        RECT 35.890 128.005 36.130 128.515 ;
        RECT 36.555 128.265 36.725 128.555 ;
        RECT 36.895 128.005 37.225 128.385 ;
        RECT 37.395 128.265 37.580 130.385 ;
        RECT 37.820 130.095 38.085 130.555 ;
        RECT 38.255 129.960 38.505 130.385 ;
        RECT 38.715 130.110 39.820 130.280 ;
        RECT 38.200 129.830 38.505 129.960 ;
        RECT 37.750 128.635 38.030 129.585 ;
        RECT 38.200 128.725 38.370 129.830 ;
        RECT 38.540 129.045 38.780 129.640 ;
        RECT 38.950 129.575 39.480 129.940 ;
        RECT 38.950 128.875 39.120 129.575 ;
        RECT 39.650 129.495 39.820 130.110 ;
        RECT 39.990 129.755 40.160 130.555 ;
        RECT 40.330 130.055 40.580 130.385 ;
        RECT 40.805 130.085 41.690 130.255 ;
        RECT 39.650 129.405 40.160 129.495 ;
        RECT 38.200 128.595 38.425 128.725 ;
        RECT 38.595 128.655 39.120 128.875 ;
        RECT 39.290 129.235 40.160 129.405 ;
        RECT 37.835 128.005 38.085 128.465 ;
        RECT 38.255 128.455 38.425 128.595 ;
        RECT 39.290 128.455 39.460 129.235 ;
        RECT 39.990 129.165 40.160 129.235 ;
        RECT 39.670 128.985 39.870 129.015 ;
        RECT 40.330 128.985 40.500 130.055 ;
        RECT 40.670 129.165 40.860 129.885 ;
        RECT 39.670 128.685 40.500 128.985 ;
        RECT 41.030 128.955 41.350 129.915 ;
        RECT 38.255 128.285 38.590 128.455 ;
        RECT 38.785 128.285 39.460 128.455 ;
        RECT 39.780 128.005 40.150 128.505 ;
        RECT 40.330 128.455 40.500 128.685 ;
        RECT 40.885 128.625 41.350 128.955 ;
        RECT 41.520 129.245 41.690 130.085 ;
        RECT 41.870 130.055 42.185 130.555 ;
        RECT 42.415 129.825 42.755 130.385 ;
        RECT 41.860 129.450 42.755 129.825 ;
        RECT 42.925 129.545 43.095 130.555 ;
        RECT 42.565 129.245 42.755 129.450 ;
        RECT 43.265 129.495 43.595 130.340 ;
        RECT 43.905 129.925 44.085 130.385 ;
        RECT 44.255 130.095 44.505 130.555 ;
        RECT 44.675 130.175 45.005 130.345 ;
        RECT 45.175 130.290 45.430 130.385 ;
        RECT 44.675 129.925 44.845 130.175 ;
        RECT 45.175 130.120 46.315 130.290 ;
        RECT 46.575 130.155 46.905 130.555 ;
        RECT 45.175 129.985 45.430 130.120 ;
        RECT 43.905 129.755 44.845 129.925 ;
        RECT 45.020 129.815 45.430 129.985 ;
        RECT 46.145 129.895 46.315 130.120 ;
        RECT 43.265 129.415 43.655 129.495 ;
        RECT 43.440 129.365 43.655 129.415 ;
        RECT 41.520 128.915 42.395 129.245 ;
        RECT 42.565 128.915 43.315 129.245 ;
        RECT 41.520 128.455 41.690 128.915 ;
        RECT 42.565 128.745 42.765 128.915 ;
        RECT 43.485 128.785 43.655 129.365 ;
        RECT 43.430 128.745 43.655 128.785 ;
        RECT 40.330 128.285 40.735 128.455 ;
        RECT 40.905 128.285 41.690 128.455 ;
        RECT 41.965 128.005 42.175 128.535 ;
        RECT 42.435 128.220 42.765 128.745 ;
        RECT 43.275 128.660 43.655 128.745 ;
        RECT 43.880 128.685 44.140 129.575 ;
        RECT 44.340 129.275 44.820 129.575 ;
        RECT 44.340 128.685 44.600 129.275 ;
        RECT 45.020 128.790 45.190 129.815 ;
        RECT 45.710 129.635 45.880 129.825 ;
        RECT 46.145 129.725 46.905 129.895 ;
        RECT 42.935 128.005 43.105 128.615 ;
        RECT 43.275 128.225 43.605 128.660 ;
        RECT 44.840 128.620 45.190 128.790 ;
        RECT 45.360 129.465 45.880 129.635 ;
        RECT 45.360 128.745 45.530 129.465 ;
        RECT 45.720 128.915 46.010 129.295 ;
        RECT 46.180 128.915 46.510 129.535 ;
        RECT 46.735 129.245 46.905 129.725 ;
        RECT 47.075 129.445 47.335 130.385 ;
        RECT 46.735 128.915 46.990 129.245 ;
        RECT 43.865 128.005 44.265 128.515 ;
        RECT 44.840 128.175 45.010 128.620 ;
        RECT 45.360 128.575 46.240 128.745 ;
        RECT 47.160 128.730 47.335 129.445 ;
        RECT 45.180 128.005 45.900 128.405 ;
        RECT 46.070 128.175 46.240 128.575 ;
        RECT 46.475 128.005 46.905 128.450 ;
        RECT 47.075 128.175 47.335 128.730 ;
        RECT 47.505 129.415 47.890 130.385 ;
        RECT 48.060 130.095 48.385 130.555 ;
        RECT 48.905 129.925 49.185 130.385 ;
        RECT 48.060 129.705 49.185 129.925 ;
        RECT 47.505 128.745 47.785 129.415 ;
        RECT 48.060 129.245 48.510 129.705 ;
        RECT 49.375 129.535 49.775 130.385 ;
        RECT 50.175 130.095 50.445 130.555 ;
        RECT 50.615 129.925 50.900 130.385 ;
        RECT 47.955 128.915 48.510 129.245 ;
        RECT 48.680 128.975 49.775 129.535 ;
        RECT 48.060 128.805 48.510 128.915 ;
        RECT 47.505 128.175 47.890 128.745 ;
        RECT 48.060 128.635 49.185 128.805 ;
        RECT 48.060 128.005 48.385 128.465 ;
        RECT 48.905 128.175 49.185 128.635 ;
        RECT 49.375 128.175 49.775 128.975 ;
        RECT 49.945 129.705 50.900 129.925 ;
        RECT 49.945 128.805 50.155 129.705 ;
        RECT 50.325 128.975 51.015 129.535 ;
        RECT 52.105 129.390 52.395 130.555 ;
        RECT 52.565 129.415 52.825 130.555 ;
        RECT 52.995 129.405 53.325 130.385 ;
        RECT 53.495 129.415 53.775 130.555 ;
        RECT 54.035 129.885 54.205 130.385 ;
        RECT 54.375 130.055 54.705 130.555 ;
        RECT 54.035 129.715 54.700 129.885 ;
        RECT 52.585 128.995 52.920 129.245 ;
        RECT 53.090 128.805 53.260 129.405 ;
        RECT 53.430 128.975 53.765 129.245 ;
        RECT 53.950 128.895 54.300 129.545 ;
        RECT 49.945 128.635 50.900 128.805 ;
        RECT 50.175 128.005 50.445 128.465 ;
        RECT 50.615 128.175 50.900 128.635 ;
        RECT 52.105 128.005 52.395 128.730 ;
        RECT 52.565 128.175 53.260 128.805 ;
        RECT 53.465 128.005 53.775 128.805 ;
        RECT 54.470 128.725 54.700 129.715 ;
        RECT 54.035 128.555 54.700 128.725 ;
        RECT 54.035 128.265 54.205 128.555 ;
        RECT 54.375 128.005 54.705 128.385 ;
        RECT 54.875 128.265 55.060 130.385 ;
        RECT 55.300 130.095 55.565 130.555 ;
        RECT 55.735 129.960 55.985 130.385 ;
        RECT 56.195 130.110 57.300 130.280 ;
        RECT 55.680 129.830 55.985 129.960 ;
        RECT 55.230 128.635 55.510 129.585 ;
        RECT 55.680 128.725 55.850 129.830 ;
        RECT 56.020 129.045 56.260 129.640 ;
        RECT 56.430 129.575 56.960 129.940 ;
        RECT 56.430 128.875 56.600 129.575 ;
        RECT 57.130 129.495 57.300 130.110 ;
        RECT 57.470 129.755 57.640 130.555 ;
        RECT 57.810 130.055 58.060 130.385 ;
        RECT 58.285 130.085 59.170 130.255 ;
        RECT 57.130 129.405 57.640 129.495 ;
        RECT 55.680 128.595 55.905 128.725 ;
        RECT 56.075 128.655 56.600 128.875 ;
        RECT 56.770 129.235 57.640 129.405 ;
        RECT 55.315 128.005 55.565 128.465 ;
        RECT 55.735 128.455 55.905 128.595 ;
        RECT 56.770 128.455 56.940 129.235 ;
        RECT 57.470 129.165 57.640 129.235 ;
        RECT 57.150 128.985 57.350 129.015 ;
        RECT 57.810 128.985 57.980 130.055 ;
        RECT 58.150 129.165 58.340 129.885 ;
        RECT 57.150 128.685 57.980 128.985 ;
        RECT 58.510 128.955 58.830 129.915 ;
        RECT 55.735 128.285 56.070 128.455 ;
        RECT 56.265 128.285 56.940 128.455 ;
        RECT 57.260 128.005 57.630 128.505 ;
        RECT 57.810 128.455 57.980 128.685 ;
        RECT 58.365 128.625 58.830 128.955 ;
        RECT 59.000 129.245 59.170 130.085 ;
        RECT 59.350 130.055 59.665 130.555 ;
        RECT 59.895 129.825 60.235 130.385 ;
        RECT 59.340 129.450 60.235 129.825 ;
        RECT 60.405 129.545 60.575 130.555 ;
        RECT 60.045 129.245 60.235 129.450 ;
        RECT 60.745 129.495 61.075 130.340 ;
        RECT 60.745 129.415 61.135 129.495 ;
        RECT 61.305 129.465 64.815 130.555 ;
        RECT 65.530 129.935 65.705 130.385 ;
        RECT 65.875 130.115 66.205 130.555 ;
        RECT 66.510 129.965 66.680 130.385 ;
        RECT 66.915 130.145 67.585 130.555 ;
        RECT 67.800 129.965 67.970 130.385 ;
        RECT 68.170 130.145 68.500 130.555 ;
        RECT 65.530 129.765 66.160 129.935 ;
        RECT 60.920 129.365 61.135 129.415 ;
        RECT 59.000 128.915 59.875 129.245 ;
        RECT 60.045 128.915 60.795 129.245 ;
        RECT 59.000 128.455 59.170 128.915 ;
        RECT 60.045 128.745 60.245 128.915 ;
        RECT 60.965 128.785 61.135 129.365 ;
        RECT 60.910 128.745 61.135 128.785 ;
        RECT 57.810 128.285 58.215 128.455 ;
        RECT 58.385 128.285 59.170 128.455 ;
        RECT 59.445 128.005 59.655 128.535 ;
        RECT 59.915 128.220 60.245 128.745 ;
        RECT 60.755 128.660 61.135 128.745 ;
        RECT 61.305 128.775 62.955 129.295 ;
        RECT 63.125 128.945 64.815 129.465 ;
        RECT 65.445 128.915 65.810 129.595 ;
        RECT 65.990 129.245 66.160 129.765 ;
        RECT 66.510 129.795 68.525 129.965 ;
        RECT 65.990 128.915 66.340 129.245 ;
        RECT 60.415 128.005 60.585 128.615 ;
        RECT 60.755 128.225 61.085 128.660 ;
        RECT 61.305 128.005 64.815 128.775 ;
        RECT 65.990 128.745 66.160 128.915 ;
        RECT 65.530 128.575 66.160 128.745 ;
        RECT 65.530 128.175 65.705 128.575 ;
        RECT 66.510 128.505 66.680 129.795 ;
        RECT 65.875 128.005 66.205 128.385 ;
        RECT 66.450 128.175 66.680 128.505 ;
        RECT 66.880 128.340 67.160 129.615 ;
        RECT 67.385 128.515 67.655 129.615 ;
        RECT 67.845 128.585 68.185 129.615 ;
        RECT 68.355 129.245 68.525 129.795 ;
        RECT 68.695 129.415 68.955 130.385 ;
        RECT 69.125 130.120 74.470 130.555 ;
        RECT 68.355 128.915 68.615 129.245 ;
        RECT 68.785 128.725 68.955 129.415 ;
        RECT 67.345 128.345 67.655 128.515 ;
        RECT 67.385 128.340 67.655 128.345 ;
        RECT 68.115 128.005 68.445 128.385 ;
        RECT 68.615 128.260 68.955 128.725 ;
        RECT 70.710 128.550 71.050 129.380 ;
        RECT 72.530 128.870 72.880 130.120 ;
        RECT 74.645 129.465 77.235 130.555 ;
        RECT 74.645 128.775 75.855 129.295 ;
        RECT 76.025 128.945 77.235 129.465 ;
        RECT 77.865 129.390 78.155 130.555 ;
        RECT 78.325 130.120 83.670 130.555 ;
        RECT 83.845 130.120 89.190 130.555 ;
        RECT 68.615 128.215 68.950 128.260 ;
        RECT 69.125 128.005 74.470 128.550 ;
        RECT 74.645 128.005 77.235 128.775 ;
        RECT 77.865 128.005 78.155 128.730 ;
        RECT 79.910 128.550 80.250 129.380 ;
        RECT 81.730 128.870 82.080 130.120 ;
        RECT 85.430 128.550 85.770 129.380 ;
        RECT 87.250 128.870 87.600 130.120 ;
        RECT 89.365 129.465 90.575 130.555 ;
        RECT 89.365 128.755 89.885 129.295 ;
        RECT 90.055 128.925 90.575 129.465 ;
        RECT 90.745 129.465 91.955 130.555 ;
        RECT 90.745 128.925 91.265 129.465 ;
        RECT 100.140 129.320 100.810 131.580 ;
        RECT 101.480 131.010 105.520 131.180 ;
        RECT 101.140 129.950 101.310 130.950 ;
        RECT 105.690 129.950 105.860 130.950 ;
        RECT 101.480 129.720 105.520 129.890 ;
        RECT 106.200 129.320 106.370 131.580 ;
        RECT 91.435 128.755 91.955 129.295 ;
        RECT 78.325 128.005 83.670 128.550 ;
        RECT 83.845 128.005 89.190 128.550 ;
        RECT 89.365 128.005 90.575 128.755 ;
        RECT 90.745 128.005 91.955 128.755 ;
        RECT 100.140 129.150 106.370 129.320 ;
        RECT 13.380 127.835 92.040 128.005 ;
        RECT 13.465 127.085 14.675 127.835 ;
        RECT 14.845 127.290 20.190 127.835 ;
        RECT 20.365 127.290 25.710 127.835 ;
        RECT 13.465 126.545 13.985 127.085 ;
        RECT 14.155 126.375 14.675 126.915 ;
        RECT 16.430 126.460 16.770 127.290 ;
        RECT 13.465 125.285 14.675 126.375 ;
        RECT 18.250 125.720 18.600 126.970 ;
        RECT 21.950 126.460 22.290 127.290 ;
        RECT 25.885 127.065 28.475 127.835 ;
        RECT 28.695 127.180 29.025 127.615 ;
        RECT 29.195 127.225 29.365 127.835 ;
        RECT 28.645 127.095 29.025 127.180 ;
        RECT 29.535 127.095 29.865 127.620 ;
        RECT 30.125 127.305 30.335 127.835 ;
        RECT 30.610 127.385 31.395 127.555 ;
        RECT 31.565 127.385 31.970 127.555 ;
        RECT 23.770 125.720 24.120 126.970 ;
        RECT 25.885 126.545 27.095 127.065 ;
        RECT 28.645 127.055 28.870 127.095 ;
        RECT 27.265 126.375 28.475 126.895 ;
        RECT 14.845 125.285 20.190 125.720 ;
        RECT 20.365 125.285 25.710 125.720 ;
        RECT 25.885 125.285 28.475 126.375 ;
        RECT 28.645 126.475 28.815 127.055 ;
        RECT 29.535 126.925 29.735 127.095 ;
        RECT 30.610 126.925 30.780 127.385 ;
        RECT 28.985 126.595 29.735 126.925 ;
        RECT 29.905 126.595 30.780 126.925 ;
        RECT 28.645 126.425 28.860 126.475 ;
        RECT 28.645 126.345 29.035 126.425 ;
        RECT 28.705 125.500 29.035 126.345 ;
        RECT 29.545 126.390 29.735 126.595 ;
        RECT 29.205 125.285 29.375 126.295 ;
        RECT 29.545 126.015 30.440 126.390 ;
        RECT 29.545 125.455 29.885 126.015 ;
        RECT 30.115 125.285 30.430 125.785 ;
        RECT 30.610 125.755 30.780 126.595 ;
        RECT 30.950 126.885 31.415 127.215 ;
        RECT 31.800 127.155 31.970 127.385 ;
        RECT 32.150 127.335 32.520 127.835 ;
        RECT 32.840 127.385 33.515 127.555 ;
        RECT 33.710 127.385 34.045 127.555 ;
        RECT 30.950 125.925 31.270 126.885 ;
        RECT 31.800 126.855 32.630 127.155 ;
        RECT 31.440 125.955 31.630 126.675 ;
        RECT 31.800 125.785 31.970 126.855 ;
        RECT 32.430 126.825 32.630 126.855 ;
        RECT 32.140 126.605 32.310 126.675 ;
        RECT 32.840 126.605 33.010 127.385 ;
        RECT 33.875 127.245 34.045 127.385 ;
        RECT 34.215 127.375 34.465 127.835 ;
        RECT 32.140 126.435 33.010 126.605 ;
        RECT 33.180 126.965 33.705 127.185 ;
        RECT 33.875 127.115 34.100 127.245 ;
        RECT 32.140 126.345 32.650 126.435 ;
        RECT 30.610 125.585 31.495 125.755 ;
        RECT 31.720 125.455 31.970 125.785 ;
        RECT 32.140 125.285 32.310 126.085 ;
        RECT 32.480 125.730 32.650 126.345 ;
        RECT 33.180 126.265 33.350 126.965 ;
        RECT 32.820 125.900 33.350 126.265 ;
        RECT 33.520 126.200 33.760 126.795 ;
        RECT 33.930 126.010 34.100 127.115 ;
        RECT 34.270 126.255 34.550 127.205 ;
        RECT 33.795 125.880 34.100 126.010 ;
        RECT 32.480 125.560 33.585 125.730 ;
        RECT 33.795 125.455 34.045 125.880 ;
        RECT 34.215 125.285 34.480 125.745 ;
        RECT 34.720 125.455 34.905 127.575 ;
        RECT 35.075 127.455 35.405 127.835 ;
        RECT 35.575 127.285 35.745 127.575 ;
        RECT 35.080 127.115 35.745 127.285 ;
        RECT 35.080 126.125 35.310 127.115 ;
        RECT 36.005 127.095 36.325 127.575 ;
        RECT 36.495 127.265 36.725 127.665 ;
        RECT 36.895 127.445 37.245 127.835 ;
        RECT 36.495 127.185 37.005 127.265 ;
        RECT 37.415 127.185 37.745 127.665 ;
        RECT 36.495 127.095 37.745 127.185 ;
        RECT 35.480 126.295 35.830 126.945 ;
        RECT 36.005 126.165 36.175 127.095 ;
        RECT 36.835 127.015 37.745 127.095 ;
        RECT 37.915 127.015 38.085 127.835 ;
        RECT 38.590 127.095 39.055 127.640 ;
        RECT 39.225 127.110 39.515 127.835 ;
        RECT 40.720 127.205 41.005 127.665 ;
        RECT 41.175 127.375 41.445 127.835 ;
        RECT 36.345 126.505 36.515 126.925 ;
        RECT 36.745 126.675 37.345 126.845 ;
        RECT 36.345 126.335 37.005 126.505 ;
        RECT 35.080 125.955 35.745 126.125 ;
        RECT 36.005 125.965 36.665 126.165 ;
        RECT 36.835 126.135 37.005 126.335 ;
        RECT 37.175 126.475 37.345 126.675 ;
        RECT 37.515 126.645 38.210 126.845 ;
        RECT 38.470 126.475 38.715 126.925 ;
        RECT 37.175 126.305 38.715 126.475 ;
        RECT 38.885 126.135 39.055 127.095 ;
        RECT 40.720 127.035 41.675 127.205 ;
        RECT 36.835 125.965 39.055 126.135 ;
        RECT 35.075 125.285 35.405 125.785 ;
        RECT 35.575 125.455 35.745 125.955 ;
        RECT 36.495 125.795 36.665 125.965 ;
        RECT 36.025 125.285 36.325 125.795 ;
        RECT 36.495 125.625 36.875 125.795 ;
        RECT 37.455 125.285 38.085 125.795 ;
        RECT 38.255 125.455 38.585 125.965 ;
        RECT 38.755 125.285 39.055 125.795 ;
        RECT 39.225 125.285 39.515 126.450 ;
        RECT 40.605 126.305 41.295 126.865 ;
        RECT 41.465 126.135 41.675 127.035 ;
        RECT 40.720 125.915 41.675 126.135 ;
        RECT 41.845 126.865 42.245 127.665 ;
        RECT 42.435 127.205 42.715 127.665 ;
        RECT 43.235 127.375 43.560 127.835 ;
        RECT 42.435 127.035 43.560 127.205 ;
        RECT 43.730 127.095 44.115 127.665 ;
        RECT 44.325 127.325 44.725 127.835 ;
        RECT 45.300 127.220 45.470 127.665 ;
        RECT 45.640 127.435 46.360 127.835 ;
        RECT 46.530 127.265 46.700 127.665 ;
        RECT 46.935 127.390 47.365 127.835 ;
        RECT 43.110 126.925 43.560 127.035 ;
        RECT 41.845 126.305 42.940 126.865 ;
        RECT 43.110 126.595 43.665 126.925 ;
        RECT 40.720 125.455 41.005 125.915 ;
        RECT 41.175 125.285 41.445 125.745 ;
        RECT 41.845 125.455 42.245 126.305 ;
        RECT 43.110 126.135 43.560 126.595 ;
        RECT 43.835 126.425 44.115 127.095 ;
        RECT 42.435 125.915 43.560 126.135 ;
        RECT 42.435 125.455 42.715 125.915 ;
        RECT 43.235 125.285 43.560 125.745 ;
        RECT 43.730 125.455 44.115 126.425 ;
        RECT 44.340 126.265 44.600 127.155 ;
        RECT 44.800 126.565 45.060 127.155 ;
        RECT 45.300 127.050 45.650 127.220 ;
        RECT 44.800 126.265 45.280 126.565 ;
        RECT 44.365 125.915 45.305 126.085 ;
        RECT 44.365 125.455 44.545 125.915 ;
        RECT 44.715 125.285 44.965 125.745 ;
        RECT 45.135 125.665 45.305 125.915 ;
        RECT 45.480 126.025 45.650 127.050 ;
        RECT 45.820 127.095 46.700 127.265 ;
        RECT 47.535 127.110 47.795 127.665 ;
        RECT 48.055 127.285 48.225 127.575 ;
        RECT 48.395 127.455 48.725 127.835 ;
        RECT 48.055 127.115 48.720 127.285 ;
        RECT 45.820 126.375 45.990 127.095 ;
        RECT 46.180 126.545 46.470 126.925 ;
        RECT 45.820 126.205 46.340 126.375 ;
        RECT 46.640 126.305 46.970 126.925 ;
        RECT 47.195 126.595 47.450 126.925 ;
        RECT 45.480 125.855 45.890 126.025 ;
        RECT 46.170 126.015 46.340 126.205 ;
        RECT 47.195 126.115 47.365 126.595 ;
        RECT 47.620 126.395 47.795 127.110 ;
        RECT 45.635 125.720 45.890 125.855 ;
        RECT 46.605 125.945 47.365 126.115 ;
        RECT 46.605 125.720 46.775 125.945 ;
        RECT 45.135 125.495 45.465 125.665 ;
        RECT 45.635 125.550 46.775 125.720 ;
        RECT 45.635 125.455 45.890 125.550 ;
        RECT 47.035 125.285 47.365 125.685 ;
        RECT 47.535 125.455 47.795 126.395 ;
        RECT 47.970 126.295 48.320 126.945 ;
        RECT 48.490 126.125 48.720 127.115 ;
        RECT 48.055 125.955 48.720 126.125 ;
        RECT 48.055 125.455 48.225 125.955 ;
        RECT 48.395 125.285 48.725 125.785 ;
        RECT 48.895 125.455 49.080 127.575 ;
        RECT 49.335 127.375 49.585 127.835 ;
        RECT 49.755 127.385 50.090 127.555 ;
        RECT 50.285 127.385 50.960 127.555 ;
        RECT 49.755 127.245 49.925 127.385 ;
        RECT 49.250 126.255 49.530 127.205 ;
        RECT 49.700 127.115 49.925 127.245 ;
        RECT 49.700 126.010 49.870 127.115 ;
        RECT 50.095 126.965 50.620 127.185 ;
        RECT 50.040 126.200 50.280 126.795 ;
        RECT 50.450 126.265 50.620 126.965 ;
        RECT 50.790 126.605 50.960 127.385 ;
        RECT 51.280 127.335 51.650 127.835 ;
        RECT 51.830 127.385 52.235 127.555 ;
        RECT 52.405 127.385 53.190 127.555 ;
        RECT 51.830 127.155 52.000 127.385 ;
        RECT 51.170 126.855 52.000 127.155 ;
        RECT 52.385 126.885 52.850 127.215 ;
        RECT 51.170 126.825 51.370 126.855 ;
        RECT 51.490 126.605 51.660 126.675 ;
        RECT 50.790 126.435 51.660 126.605 ;
        RECT 51.150 126.345 51.660 126.435 ;
        RECT 49.700 125.880 50.005 126.010 ;
        RECT 50.450 125.900 50.980 126.265 ;
        RECT 49.320 125.285 49.585 125.745 ;
        RECT 49.755 125.455 50.005 125.880 ;
        RECT 51.150 125.730 51.320 126.345 ;
        RECT 50.215 125.560 51.320 125.730 ;
        RECT 51.490 125.285 51.660 126.085 ;
        RECT 51.830 125.785 52.000 126.855 ;
        RECT 52.170 125.955 52.360 126.675 ;
        RECT 52.530 125.925 52.850 126.885 ;
        RECT 53.020 126.925 53.190 127.385 ;
        RECT 53.465 127.305 53.675 127.835 ;
        RECT 53.935 127.095 54.265 127.620 ;
        RECT 54.435 127.225 54.605 127.835 ;
        RECT 54.775 127.180 55.105 127.615 ;
        RECT 55.325 127.290 60.670 127.835 ;
        RECT 54.775 127.095 55.155 127.180 ;
        RECT 54.065 126.925 54.265 127.095 ;
        RECT 54.930 127.055 55.155 127.095 ;
        RECT 53.020 126.595 53.895 126.925 ;
        RECT 54.065 126.595 54.815 126.925 ;
        RECT 51.830 125.455 52.080 125.785 ;
        RECT 53.020 125.755 53.190 126.595 ;
        RECT 54.065 126.390 54.255 126.595 ;
        RECT 54.985 126.475 55.155 127.055 ;
        RECT 54.940 126.425 55.155 126.475 ;
        RECT 56.910 126.460 57.250 127.290 ;
        RECT 60.845 127.065 64.355 127.835 ;
        RECT 64.985 127.110 65.275 127.835 ;
        RECT 65.445 127.290 70.790 127.835 ;
        RECT 70.965 127.290 76.310 127.835 ;
        RECT 76.485 127.290 81.830 127.835 ;
        RECT 82.005 127.290 87.350 127.835 ;
        RECT 53.360 126.015 54.255 126.390 ;
        RECT 54.765 126.345 55.155 126.425 ;
        RECT 52.305 125.585 53.190 125.755 ;
        RECT 53.370 125.285 53.685 125.785 ;
        RECT 53.915 125.455 54.255 126.015 ;
        RECT 54.425 125.285 54.595 126.295 ;
        RECT 54.765 125.500 55.095 126.345 ;
        RECT 58.730 125.720 59.080 126.970 ;
        RECT 60.845 126.545 62.495 127.065 ;
        RECT 62.665 126.375 64.355 126.895 ;
        RECT 67.030 126.460 67.370 127.290 ;
        RECT 55.325 125.285 60.670 125.720 ;
        RECT 60.845 125.285 64.355 126.375 ;
        RECT 64.985 125.285 65.275 126.450 ;
        RECT 68.850 125.720 69.200 126.970 ;
        RECT 72.550 126.460 72.890 127.290 ;
        RECT 74.370 125.720 74.720 126.970 ;
        RECT 78.070 126.460 78.410 127.290 ;
        RECT 79.890 125.720 80.240 126.970 ;
        RECT 83.590 126.460 83.930 127.290 ;
        RECT 87.525 127.065 90.115 127.835 ;
        RECT 90.745 127.085 91.955 127.835 ;
        RECT 85.410 125.720 85.760 126.970 ;
        RECT 87.525 126.545 88.735 127.065 ;
        RECT 88.905 126.375 90.115 126.895 ;
        RECT 65.445 125.285 70.790 125.720 ;
        RECT 70.965 125.285 76.310 125.720 ;
        RECT 76.485 125.285 81.830 125.720 ;
        RECT 82.005 125.285 87.350 125.720 ;
        RECT 87.525 125.285 90.115 126.375 ;
        RECT 90.745 126.375 91.265 126.915 ;
        RECT 91.435 126.545 91.955 127.085 ;
        RECT 90.745 125.285 91.955 126.375 ;
        RECT 100.140 125.890 100.810 129.150 ;
        RECT 101.480 128.580 105.520 128.750 ;
        RECT 101.140 126.520 101.310 128.520 ;
        RECT 105.690 126.520 105.860 128.520 ;
        RECT 101.480 126.290 105.520 126.460 ;
        RECT 106.200 125.890 106.370 129.150 ;
        RECT 100.140 125.720 106.370 125.890 ;
        RECT 13.380 125.115 92.040 125.285 ;
        RECT 13.465 124.025 14.675 125.115 ;
        RECT 14.845 124.680 20.190 125.115 ;
        RECT 20.365 124.680 25.710 125.115 ;
        RECT 13.465 123.315 13.985 123.855 ;
        RECT 14.155 123.485 14.675 124.025 ;
        RECT 13.465 122.565 14.675 123.315 ;
        RECT 16.430 123.110 16.770 123.940 ;
        RECT 18.250 123.430 18.600 124.680 ;
        RECT 21.950 123.110 22.290 123.940 ;
        RECT 23.770 123.430 24.120 124.680 ;
        RECT 26.345 123.950 26.635 125.115 ;
        RECT 26.805 124.025 28.015 125.115 ;
        RECT 28.300 124.485 28.585 124.945 ;
        RECT 28.755 124.655 29.025 125.115 ;
        RECT 28.300 124.265 29.255 124.485 ;
        RECT 26.805 123.315 27.325 123.855 ;
        RECT 27.495 123.485 28.015 124.025 ;
        RECT 28.185 123.535 28.875 124.095 ;
        RECT 29.045 123.365 29.255 124.265 ;
        RECT 14.845 122.565 20.190 123.110 ;
        RECT 20.365 122.565 25.710 123.110 ;
        RECT 26.345 122.565 26.635 123.290 ;
        RECT 26.805 122.565 28.015 123.315 ;
        RECT 28.300 123.195 29.255 123.365 ;
        RECT 29.425 124.095 29.825 124.945 ;
        RECT 30.015 124.485 30.295 124.945 ;
        RECT 30.815 124.655 31.140 125.115 ;
        RECT 30.015 124.265 31.140 124.485 ;
        RECT 29.425 123.535 30.520 124.095 ;
        RECT 30.690 123.805 31.140 124.265 ;
        RECT 31.310 123.975 31.695 124.945 ;
        RECT 31.865 124.025 34.455 125.115 ;
        RECT 28.300 122.735 28.585 123.195 ;
        RECT 28.755 122.565 29.025 123.025 ;
        RECT 29.425 122.735 29.825 123.535 ;
        RECT 30.690 123.475 31.245 123.805 ;
        RECT 30.690 123.365 31.140 123.475 ;
        RECT 30.015 123.195 31.140 123.365 ;
        RECT 31.415 123.305 31.695 123.975 ;
        RECT 30.015 122.735 30.295 123.195 ;
        RECT 30.815 122.565 31.140 123.025 ;
        RECT 31.310 122.735 31.695 123.305 ;
        RECT 31.865 123.335 33.075 123.855 ;
        RECT 33.245 123.505 34.455 124.025 ;
        RECT 35.085 123.550 35.435 124.945 ;
        RECT 35.605 124.315 36.010 125.115 ;
        RECT 36.180 124.775 37.715 124.945 ;
        RECT 36.180 124.145 36.350 124.775 ;
        RECT 35.605 123.975 36.350 124.145 ;
        RECT 31.865 122.565 34.455 123.335 ;
        RECT 35.085 122.735 35.355 123.550 ;
        RECT 35.605 123.475 35.775 123.975 ;
        RECT 36.520 123.805 36.790 124.550 ;
        RECT 35.945 123.475 36.280 123.805 ;
        RECT 36.450 123.475 36.790 123.805 ;
        RECT 36.980 123.805 37.215 124.550 ;
        RECT 37.385 124.145 37.715 124.775 ;
        RECT 37.900 124.315 38.135 125.115 ;
        RECT 38.305 124.145 38.595 124.945 ;
        RECT 37.385 123.975 38.595 124.145 ;
        RECT 38.765 124.525 39.465 124.945 ;
        RECT 39.665 124.755 39.995 125.115 ;
        RECT 40.165 124.525 40.495 124.925 ;
        RECT 38.765 124.295 40.495 124.525 ;
        RECT 36.980 123.475 37.270 123.805 ;
        RECT 37.440 123.475 37.840 123.805 ;
        RECT 38.010 123.305 38.180 123.975 ;
        RECT 38.350 123.475 38.595 123.805 ;
        RECT 38.765 123.325 38.970 124.295 ;
        RECT 39.140 123.555 39.470 124.095 ;
        RECT 39.645 123.805 39.970 124.095 ;
        RECT 40.165 124.075 40.495 124.295 ;
        RECT 40.665 123.805 40.835 124.775 ;
        RECT 41.015 124.055 41.345 125.115 ;
        RECT 41.615 124.445 41.785 124.945 ;
        RECT 41.955 124.615 42.285 125.115 ;
        RECT 41.615 124.275 42.280 124.445 ;
        RECT 39.645 123.475 40.140 123.805 ;
        RECT 40.460 123.475 40.835 123.805 ;
        RECT 41.045 123.475 41.355 123.805 ;
        RECT 41.530 123.455 41.880 124.105 ;
        RECT 35.525 122.565 36.195 123.305 ;
        RECT 36.365 123.135 37.760 123.305 ;
        RECT 36.365 122.790 36.660 123.135 ;
        RECT 36.840 122.565 37.215 122.965 ;
        RECT 37.430 122.790 37.760 123.135 ;
        RECT 38.010 122.735 38.595 123.305 ;
        RECT 38.765 122.735 39.475 123.325 ;
        RECT 39.985 123.095 41.345 123.305 ;
        RECT 42.050 123.285 42.280 124.275 ;
        RECT 39.985 122.735 40.315 123.095 ;
        RECT 40.515 122.565 40.845 122.925 ;
        RECT 41.015 122.735 41.345 123.095 ;
        RECT 41.615 123.115 42.280 123.285 ;
        RECT 41.615 122.825 41.785 123.115 ;
        RECT 41.955 122.565 42.285 122.945 ;
        RECT 42.455 122.825 42.640 124.945 ;
        RECT 42.880 124.655 43.145 125.115 ;
        RECT 43.315 124.520 43.565 124.945 ;
        RECT 43.775 124.670 44.880 124.840 ;
        RECT 43.260 124.390 43.565 124.520 ;
        RECT 42.810 123.195 43.090 124.145 ;
        RECT 43.260 123.285 43.430 124.390 ;
        RECT 43.600 123.605 43.840 124.200 ;
        RECT 44.010 124.135 44.540 124.500 ;
        RECT 44.010 123.435 44.180 124.135 ;
        RECT 44.710 124.055 44.880 124.670 ;
        RECT 45.050 124.315 45.220 125.115 ;
        RECT 45.390 124.615 45.640 124.945 ;
        RECT 45.865 124.645 46.750 124.815 ;
        RECT 44.710 123.965 45.220 124.055 ;
        RECT 43.260 123.155 43.485 123.285 ;
        RECT 43.655 123.215 44.180 123.435 ;
        RECT 44.350 123.795 45.220 123.965 ;
        RECT 42.895 122.565 43.145 123.025 ;
        RECT 43.315 123.015 43.485 123.155 ;
        RECT 44.350 123.015 44.520 123.795 ;
        RECT 45.050 123.725 45.220 123.795 ;
        RECT 44.730 123.545 44.930 123.575 ;
        RECT 45.390 123.545 45.560 124.615 ;
        RECT 45.730 123.725 45.920 124.445 ;
        RECT 44.730 123.245 45.560 123.545 ;
        RECT 46.090 123.515 46.410 124.475 ;
        RECT 43.315 122.845 43.650 123.015 ;
        RECT 43.845 122.845 44.520 123.015 ;
        RECT 44.840 122.565 45.210 123.065 ;
        RECT 45.390 123.015 45.560 123.245 ;
        RECT 45.945 123.185 46.410 123.515 ;
        RECT 46.580 123.805 46.750 124.645 ;
        RECT 46.930 124.615 47.245 125.115 ;
        RECT 47.475 124.385 47.815 124.945 ;
        RECT 46.920 124.010 47.815 124.385 ;
        RECT 47.985 124.105 48.155 125.115 ;
        RECT 47.625 123.805 47.815 124.010 ;
        RECT 48.325 124.055 48.655 124.900 ;
        RECT 48.885 124.605 50.075 124.895 ;
        RECT 48.905 124.265 50.075 124.435 ;
        RECT 50.245 124.315 50.525 125.115 ;
        RECT 48.325 123.975 48.715 124.055 ;
        RECT 48.905 123.975 49.230 124.265 ;
        RECT 49.905 124.145 50.075 124.265 ;
        RECT 48.500 123.925 48.715 123.975 ;
        RECT 46.580 123.475 47.455 123.805 ;
        RECT 47.625 123.475 48.375 123.805 ;
        RECT 46.580 123.015 46.750 123.475 ;
        RECT 47.625 123.305 47.825 123.475 ;
        RECT 48.545 123.345 48.715 123.925 ;
        RECT 49.400 123.805 49.595 124.095 ;
        RECT 49.905 123.975 50.565 124.145 ;
        RECT 50.735 123.975 51.010 124.945 ;
        RECT 50.395 123.805 50.565 123.975 ;
        RECT 48.885 123.475 49.230 123.805 ;
        RECT 49.400 123.475 50.225 123.805 ;
        RECT 50.395 123.475 50.670 123.805 ;
        RECT 48.490 123.305 48.715 123.345 ;
        RECT 50.395 123.305 50.565 123.475 ;
        RECT 45.390 122.845 45.795 123.015 ;
        RECT 45.965 122.845 46.750 123.015 ;
        RECT 47.025 122.565 47.235 123.095 ;
        RECT 47.495 122.780 47.825 123.305 ;
        RECT 48.335 123.220 48.715 123.305 ;
        RECT 47.995 122.565 48.165 123.175 ;
        RECT 48.335 122.785 48.665 123.220 ;
        RECT 48.900 123.135 50.565 123.305 ;
        RECT 50.840 123.240 51.010 123.975 ;
        RECT 52.105 123.950 52.395 125.115 ;
        RECT 52.565 124.145 52.875 124.945 ;
        RECT 53.045 124.315 53.355 125.115 ;
        RECT 53.525 124.485 53.785 124.945 ;
        RECT 53.955 124.655 54.210 125.115 ;
        RECT 54.385 124.485 54.645 124.945 ;
        RECT 53.525 124.315 54.645 124.485 ;
        RECT 54.005 124.265 54.175 124.315 ;
        RECT 52.565 123.975 53.595 124.145 ;
        RECT 48.900 122.785 49.155 123.135 ;
        RECT 49.325 122.565 49.655 122.965 ;
        RECT 49.825 122.785 49.995 123.135 ;
        RECT 50.165 122.565 50.545 122.965 ;
        RECT 50.735 122.895 51.010 123.240 ;
        RECT 52.105 122.565 52.395 123.290 ;
        RECT 52.565 123.065 52.735 123.975 ;
        RECT 52.905 123.235 53.255 123.805 ;
        RECT 53.425 123.725 53.595 123.975 ;
        RECT 54.385 124.065 54.645 124.315 ;
        RECT 54.815 124.245 55.100 125.115 ;
        RECT 54.385 123.895 55.140 124.065 ;
        RECT 55.325 124.025 56.995 125.115 ;
        RECT 53.425 123.555 54.565 123.725 ;
        RECT 54.735 123.385 55.140 123.895 ;
        RECT 53.490 123.215 55.140 123.385 ;
        RECT 55.325 123.335 56.075 123.855 ;
        RECT 56.245 123.505 56.995 124.025 ;
        RECT 57.165 123.975 57.550 124.945 ;
        RECT 57.720 124.655 58.045 125.115 ;
        RECT 58.565 124.485 58.845 124.945 ;
        RECT 57.720 124.265 58.845 124.485 ;
        RECT 52.565 122.735 52.865 123.065 ;
        RECT 53.035 122.565 53.310 123.045 ;
        RECT 53.490 122.825 53.785 123.215 ;
        RECT 53.955 122.565 54.210 123.045 ;
        RECT 54.385 122.825 54.645 123.215 ;
        RECT 54.815 122.565 55.095 123.045 ;
        RECT 55.325 122.565 56.995 123.335 ;
        RECT 57.165 123.305 57.445 123.975 ;
        RECT 57.720 123.805 58.170 124.265 ;
        RECT 59.035 124.095 59.435 124.945 ;
        RECT 59.835 124.655 60.105 125.115 ;
        RECT 60.275 124.485 60.560 124.945 ;
        RECT 57.615 123.475 58.170 123.805 ;
        RECT 58.340 123.535 59.435 124.095 ;
        RECT 57.720 123.365 58.170 123.475 ;
        RECT 57.165 122.735 57.550 123.305 ;
        RECT 57.720 123.195 58.845 123.365 ;
        RECT 57.720 122.565 58.045 123.025 ;
        RECT 58.565 122.735 58.845 123.195 ;
        RECT 59.035 122.735 59.435 123.535 ;
        RECT 59.605 124.265 60.560 124.485 ;
        RECT 59.605 123.365 59.815 124.265 ;
        RECT 59.985 123.535 60.675 124.095 ;
        RECT 60.845 124.025 62.515 125.115 ;
        RECT 59.605 123.195 60.560 123.365 ;
        RECT 59.835 122.565 60.105 123.025 ;
        RECT 60.275 122.735 60.560 123.195 ;
        RECT 60.845 123.335 61.595 123.855 ;
        RECT 61.765 123.505 62.515 124.025 ;
        RECT 62.685 123.975 63.070 124.945 ;
        RECT 63.240 124.655 63.565 125.115 ;
        RECT 64.085 124.485 64.365 124.945 ;
        RECT 63.240 124.265 64.365 124.485 ;
        RECT 60.845 122.565 62.515 123.335 ;
        RECT 62.685 123.305 62.965 123.975 ;
        RECT 63.240 123.805 63.690 124.265 ;
        RECT 64.555 124.095 64.955 124.945 ;
        RECT 65.355 124.655 65.625 125.115 ;
        RECT 65.795 124.485 66.080 124.945 ;
        RECT 63.135 123.475 63.690 123.805 ;
        RECT 63.860 123.535 64.955 124.095 ;
        RECT 63.240 123.365 63.690 123.475 ;
        RECT 62.685 122.735 63.070 123.305 ;
        RECT 63.240 123.195 64.365 123.365 ;
        RECT 63.240 122.565 63.565 123.025 ;
        RECT 64.085 122.735 64.365 123.195 ;
        RECT 64.555 122.735 64.955 123.535 ;
        RECT 65.125 124.265 66.080 124.485 ;
        RECT 65.125 123.365 65.335 124.265 ;
        RECT 65.505 123.535 66.195 124.095 ;
        RECT 66.365 123.975 66.705 124.945 ;
        RECT 66.875 123.975 67.045 125.115 ;
        RECT 67.315 124.315 67.565 125.115 ;
        RECT 68.210 124.145 68.540 124.945 ;
        RECT 68.840 124.315 69.170 125.115 ;
        RECT 69.340 124.145 69.670 124.945 ;
        RECT 70.045 124.680 75.390 125.115 ;
        RECT 67.235 123.975 69.670 124.145 ;
        RECT 66.365 123.925 66.595 123.975 ;
        RECT 66.365 123.365 66.540 123.925 ;
        RECT 67.235 123.725 67.405 123.975 ;
        RECT 66.710 123.555 67.405 123.725 ;
        RECT 67.580 123.555 68.000 123.755 ;
        RECT 68.170 123.555 68.500 123.755 ;
        RECT 68.670 123.555 69.000 123.755 ;
        RECT 65.125 123.195 66.080 123.365 ;
        RECT 65.355 122.565 65.625 123.025 ;
        RECT 65.795 122.735 66.080 123.195 ;
        RECT 66.365 122.735 66.705 123.365 ;
        RECT 66.875 122.565 67.125 123.365 ;
        RECT 67.315 123.215 68.540 123.385 ;
        RECT 67.315 122.735 67.645 123.215 ;
        RECT 67.815 122.565 68.040 123.025 ;
        RECT 68.210 122.735 68.540 123.215 ;
        RECT 69.170 123.345 69.340 123.975 ;
        RECT 69.525 123.555 69.875 123.805 ;
        RECT 69.170 122.735 69.670 123.345 ;
        RECT 71.630 123.110 71.970 123.940 ;
        RECT 73.450 123.430 73.800 124.680 ;
        RECT 75.565 124.025 77.235 125.115 ;
        RECT 75.565 123.335 76.315 123.855 ;
        RECT 76.485 123.505 77.235 124.025 ;
        RECT 77.865 123.950 78.155 125.115 ;
        RECT 78.325 124.680 83.670 125.115 ;
        RECT 83.845 124.680 89.190 125.115 ;
        RECT 70.045 122.565 75.390 123.110 ;
        RECT 75.565 122.565 77.235 123.335 ;
        RECT 77.865 122.565 78.155 123.290 ;
        RECT 79.910 123.110 80.250 123.940 ;
        RECT 81.730 123.430 82.080 124.680 ;
        RECT 85.430 123.110 85.770 123.940 ;
        RECT 87.250 123.430 87.600 124.680 ;
        RECT 89.365 124.025 90.575 125.115 ;
        RECT 89.365 123.315 89.885 123.855 ;
        RECT 90.055 123.485 90.575 124.025 ;
        RECT 90.745 124.025 91.955 125.115 ;
        RECT 90.745 123.485 91.265 124.025 ;
        RECT 91.435 123.315 91.955 123.855 ;
        RECT 78.325 122.565 83.670 123.110 ;
        RECT 83.845 122.565 89.190 123.110 ;
        RECT 89.365 122.565 90.575 123.315 ;
        RECT 90.745 122.565 91.955 123.315 ;
        RECT 13.380 122.395 92.040 122.565 ;
        RECT 100.140 122.460 100.810 125.720 ;
        RECT 101.480 125.150 105.520 125.320 ;
        RECT 101.140 123.090 101.310 125.090 ;
        RECT 105.690 123.090 105.860 125.090 ;
        RECT 101.480 122.860 105.520 123.030 ;
        RECT 106.200 122.460 106.370 125.720 ;
        RECT 100.140 122.450 106.370 122.460 ;
        RECT 107.960 131.720 117.790 131.760 ;
        RECT 107.960 131.590 118.590 131.720 ;
        RECT 107.960 129.330 108.130 131.590 ;
        RECT 108.855 131.020 116.895 131.190 ;
        RECT 108.470 129.960 108.640 130.960 ;
        RECT 117.110 129.960 117.280 130.960 ;
        RECT 108.855 129.730 116.895 129.900 ;
        RECT 117.620 129.330 118.590 131.590 ;
        RECT 107.960 129.160 118.590 129.330 ;
        RECT 107.960 125.900 108.130 129.160 ;
        RECT 108.855 128.590 116.895 128.760 ;
        RECT 108.470 126.530 108.640 128.530 ;
        RECT 117.110 126.530 117.280 128.530 ;
        RECT 108.855 126.300 116.895 126.470 ;
        RECT 117.620 125.900 118.590 129.160 ;
        RECT 107.960 125.730 118.590 125.900 ;
        RECT 107.960 122.470 108.130 125.730 ;
        RECT 108.855 125.160 116.895 125.330 ;
        RECT 108.470 123.100 108.640 125.100 ;
        RECT 117.110 123.100 117.280 125.100 ;
        RECT 108.855 122.870 116.895 123.040 ;
        RECT 117.620 122.470 118.590 125.730 ;
        RECT 13.465 121.645 14.675 122.395 ;
        RECT 14.845 121.850 20.190 122.395 ;
        RECT 13.465 121.105 13.985 121.645 ;
        RECT 14.155 120.935 14.675 121.475 ;
        RECT 16.430 121.020 16.770 121.850 ;
        RECT 20.365 121.625 22.955 122.395 ;
        RECT 23.215 121.845 23.385 122.135 ;
        RECT 23.555 122.015 23.885 122.395 ;
        RECT 23.215 121.675 23.880 121.845 ;
        RECT 13.465 119.845 14.675 120.935 ;
        RECT 18.250 120.280 18.600 121.530 ;
        RECT 20.365 121.105 21.575 121.625 ;
        RECT 21.745 120.935 22.955 121.455 ;
        RECT 14.845 119.845 20.190 120.280 ;
        RECT 20.365 119.845 22.955 120.935 ;
        RECT 23.130 120.855 23.480 121.505 ;
        RECT 23.650 120.685 23.880 121.675 ;
        RECT 23.215 120.515 23.880 120.685 ;
        RECT 23.215 120.015 23.385 120.515 ;
        RECT 23.555 119.845 23.885 120.345 ;
        RECT 24.055 120.015 24.240 122.135 ;
        RECT 24.495 121.935 24.745 122.395 ;
        RECT 24.915 121.945 25.250 122.115 ;
        RECT 25.445 121.945 26.120 122.115 ;
        RECT 24.915 121.805 25.085 121.945 ;
        RECT 24.410 120.815 24.690 121.765 ;
        RECT 24.860 121.675 25.085 121.805 ;
        RECT 24.860 120.570 25.030 121.675 ;
        RECT 25.255 121.525 25.780 121.745 ;
        RECT 25.200 120.760 25.440 121.355 ;
        RECT 25.610 120.825 25.780 121.525 ;
        RECT 25.950 121.165 26.120 121.945 ;
        RECT 26.440 121.895 26.810 122.395 ;
        RECT 26.990 121.945 27.395 122.115 ;
        RECT 27.565 121.945 28.350 122.115 ;
        RECT 26.990 121.715 27.160 121.945 ;
        RECT 26.330 121.415 27.160 121.715 ;
        RECT 27.545 121.445 28.010 121.775 ;
        RECT 26.330 121.385 26.530 121.415 ;
        RECT 26.650 121.165 26.820 121.235 ;
        RECT 25.950 120.995 26.820 121.165 ;
        RECT 26.310 120.905 26.820 120.995 ;
        RECT 24.860 120.440 25.165 120.570 ;
        RECT 25.610 120.460 26.140 120.825 ;
        RECT 24.480 119.845 24.745 120.305 ;
        RECT 24.915 120.015 25.165 120.440 ;
        RECT 26.310 120.290 26.480 120.905 ;
        RECT 25.375 120.120 26.480 120.290 ;
        RECT 26.650 119.845 26.820 120.645 ;
        RECT 26.990 120.345 27.160 121.415 ;
        RECT 27.330 120.515 27.520 121.235 ;
        RECT 27.690 120.485 28.010 121.445 ;
        RECT 28.180 121.485 28.350 121.945 ;
        RECT 28.625 121.865 28.835 122.395 ;
        RECT 29.095 121.655 29.425 122.180 ;
        RECT 29.595 121.785 29.765 122.395 ;
        RECT 29.935 121.740 30.265 122.175 ;
        RECT 30.485 121.850 35.830 122.395 ;
        RECT 29.935 121.655 30.315 121.740 ;
        RECT 29.225 121.485 29.425 121.655 ;
        RECT 30.090 121.615 30.315 121.655 ;
        RECT 28.180 121.155 29.055 121.485 ;
        RECT 29.225 121.155 29.975 121.485 ;
        RECT 26.990 120.015 27.240 120.345 ;
        RECT 28.180 120.315 28.350 121.155 ;
        RECT 29.225 120.950 29.415 121.155 ;
        RECT 30.145 121.035 30.315 121.615 ;
        RECT 30.100 120.985 30.315 121.035 ;
        RECT 32.070 121.020 32.410 121.850 ;
        RECT 36.005 121.625 38.595 122.395 ;
        RECT 39.225 121.670 39.515 122.395 ;
        RECT 39.685 121.850 45.030 122.395 ;
        RECT 28.520 120.575 29.415 120.950 ;
        RECT 29.925 120.905 30.315 120.985 ;
        RECT 27.465 120.145 28.350 120.315 ;
        RECT 28.530 119.845 28.845 120.345 ;
        RECT 29.075 120.015 29.415 120.575 ;
        RECT 29.585 119.845 29.755 120.855 ;
        RECT 29.925 120.060 30.255 120.905 ;
        RECT 33.890 120.280 34.240 121.530 ;
        RECT 36.005 121.105 37.215 121.625 ;
        RECT 37.385 120.935 38.595 121.455 ;
        RECT 41.270 121.020 41.610 121.850 ;
        RECT 45.240 121.655 45.855 122.225 ;
        RECT 46.025 121.885 46.240 122.395 ;
        RECT 46.470 121.885 46.750 122.215 ;
        RECT 46.930 121.885 47.170 122.395 ;
        RECT 30.485 119.845 35.830 120.280 ;
        RECT 36.005 119.845 38.595 120.935 ;
        RECT 39.225 119.845 39.515 121.010 ;
        RECT 43.090 120.280 43.440 121.530 ;
        RECT 45.240 120.635 45.555 121.655 ;
        RECT 45.725 120.985 45.895 121.485 ;
        RECT 46.145 121.155 46.410 121.715 ;
        RECT 46.580 120.985 46.750 121.885 ;
        RECT 46.920 121.155 47.275 121.715 ;
        RECT 47.565 121.575 47.775 122.395 ;
        RECT 47.945 121.595 48.275 122.225 ;
        RECT 47.945 120.995 48.195 121.595 ;
        RECT 48.445 121.575 48.675 122.395 ;
        RECT 48.895 121.585 49.165 122.395 ;
        RECT 49.335 121.585 49.665 122.225 ;
        RECT 49.835 121.585 50.075 122.395 ;
        RECT 50.265 121.625 53.775 122.395 ;
        RECT 53.945 121.645 55.155 122.395 ;
        RECT 55.415 121.845 55.585 122.135 ;
        RECT 55.755 122.015 56.085 122.395 ;
        RECT 55.415 121.675 56.080 121.845 ;
        RECT 48.365 121.155 48.695 121.405 ;
        RECT 48.885 121.155 49.235 121.405 ;
        RECT 45.725 120.815 47.150 120.985 ;
        RECT 39.685 119.845 45.030 120.280 ;
        RECT 45.240 120.015 45.775 120.635 ;
        RECT 45.945 119.845 46.275 120.645 ;
        RECT 46.760 120.640 47.150 120.815 ;
        RECT 47.565 119.845 47.775 120.985 ;
        RECT 47.945 120.015 48.275 120.995 ;
        RECT 49.405 120.985 49.575 121.585 ;
        RECT 49.745 121.155 50.095 121.405 ;
        RECT 50.265 121.105 51.915 121.625 ;
        RECT 48.445 119.845 48.675 120.985 ;
        RECT 48.895 119.845 49.225 120.985 ;
        RECT 49.405 120.815 50.085 120.985 ;
        RECT 52.085 120.935 53.775 121.455 ;
        RECT 53.945 121.105 54.465 121.645 ;
        RECT 54.635 120.935 55.155 121.475 ;
        RECT 49.755 120.030 50.085 120.815 ;
        RECT 50.265 119.845 53.775 120.935 ;
        RECT 53.945 119.845 55.155 120.935 ;
        RECT 55.330 120.855 55.680 121.505 ;
        RECT 55.850 120.685 56.080 121.675 ;
        RECT 55.415 120.515 56.080 120.685 ;
        RECT 55.415 120.015 55.585 120.515 ;
        RECT 55.755 119.845 56.085 120.345 ;
        RECT 56.255 120.015 56.440 122.135 ;
        RECT 56.695 121.935 56.945 122.395 ;
        RECT 57.115 121.945 57.450 122.115 ;
        RECT 57.645 121.945 58.320 122.115 ;
        RECT 57.115 121.805 57.285 121.945 ;
        RECT 56.610 120.815 56.890 121.765 ;
        RECT 57.060 121.675 57.285 121.805 ;
        RECT 57.060 120.570 57.230 121.675 ;
        RECT 57.455 121.525 57.980 121.745 ;
        RECT 57.400 120.760 57.640 121.355 ;
        RECT 57.810 120.825 57.980 121.525 ;
        RECT 58.150 121.165 58.320 121.945 ;
        RECT 58.640 121.895 59.010 122.395 ;
        RECT 59.190 121.945 59.595 122.115 ;
        RECT 59.765 121.945 60.550 122.115 ;
        RECT 59.190 121.715 59.360 121.945 ;
        RECT 58.530 121.415 59.360 121.715 ;
        RECT 59.745 121.445 60.210 121.775 ;
        RECT 58.530 121.385 58.730 121.415 ;
        RECT 58.850 121.165 59.020 121.235 ;
        RECT 58.150 120.995 59.020 121.165 ;
        RECT 58.510 120.905 59.020 120.995 ;
        RECT 57.060 120.440 57.365 120.570 ;
        RECT 57.810 120.460 58.340 120.825 ;
        RECT 56.680 119.845 56.945 120.305 ;
        RECT 57.115 120.015 57.365 120.440 ;
        RECT 58.510 120.290 58.680 120.905 ;
        RECT 57.575 120.120 58.680 120.290 ;
        RECT 58.850 119.845 59.020 120.645 ;
        RECT 59.190 120.345 59.360 121.415 ;
        RECT 59.530 120.515 59.720 121.235 ;
        RECT 59.890 120.485 60.210 121.445 ;
        RECT 60.380 121.485 60.550 121.945 ;
        RECT 60.825 121.865 61.035 122.395 ;
        RECT 61.295 121.655 61.625 122.180 ;
        RECT 61.795 121.785 61.965 122.395 ;
        RECT 62.135 121.740 62.465 122.175 ;
        RECT 62.135 121.655 62.515 121.740 ;
        RECT 61.425 121.485 61.625 121.655 ;
        RECT 62.290 121.615 62.515 121.655 ;
        RECT 60.380 121.155 61.255 121.485 ;
        RECT 61.425 121.155 62.175 121.485 ;
        RECT 59.190 120.015 59.440 120.345 ;
        RECT 60.380 120.315 60.550 121.155 ;
        RECT 61.425 120.950 61.615 121.155 ;
        RECT 62.345 121.035 62.515 121.615 ;
        RECT 62.705 121.585 62.945 122.395 ;
        RECT 63.115 121.585 63.445 122.225 ;
        RECT 63.615 121.585 63.885 122.395 ;
        RECT 64.985 121.670 65.275 122.395 ;
        RECT 65.445 121.625 67.115 122.395 ;
        RECT 67.335 121.740 67.665 122.175 ;
        RECT 67.835 121.785 68.005 122.395 ;
        RECT 67.285 121.655 67.665 121.740 ;
        RECT 68.175 121.655 68.505 122.180 ;
        RECT 68.765 121.865 68.975 122.395 ;
        RECT 69.250 121.945 70.035 122.115 ;
        RECT 70.205 121.945 70.610 122.115 ;
        RECT 62.685 121.155 63.035 121.405 ;
        RECT 62.300 120.985 62.515 121.035 ;
        RECT 63.205 120.985 63.375 121.585 ;
        RECT 63.545 121.155 63.895 121.405 ;
        RECT 65.445 121.105 66.195 121.625 ;
        RECT 67.285 121.615 67.510 121.655 ;
        RECT 60.720 120.575 61.615 120.950 ;
        RECT 62.125 120.905 62.515 120.985 ;
        RECT 59.665 120.145 60.550 120.315 ;
        RECT 60.730 119.845 61.045 120.345 ;
        RECT 61.275 120.015 61.615 120.575 ;
        RECT 61.785 119.845 61.955 120.855 ;
        RECT 62.125 120.060 62.455 120.905 ;
        RECT 62.695 120.815 63.375 120.985 ;
        RECT 62.695 120.030 63.025 120.815 ;
        RECT 63.555 119.845 63.885 120.985 ;
        RECT 64.985 119.845 65.275 121.010 ;
        RECT 66.365 120.935 67.115 121.455 ;
        RECT 65.445 119.845 67.115 120.935 ;
        RECT 67.285 121.035 67.455 121.615 ;
        RECT 68.175 121.485 68.375 121.655 ;
        RECT 69.250 121.485 69.420 121.945 ;
        RECT 67.625 121.155 68.375 121.485 ;
        RECT 68.545 121.155 69.420 121.485 ;
        RECT 67.285 120.985 67.500 121.035 ;
        RECT 67.285 120.905 67.675 120.985 ;
        RECT 67.345 120.060 67.675 120.905 ;
        RECT 68.185 120.950 68.375 121.155 ;
        RECT 67.845 119.845 68.015 120.855 ;
        RECT 68.185 120.575 69.080 120.950 ;
        RECT 68.185 120.015 68.525 120.575 ;
        RECT 68.755 119.845 69.070 120.345 ;
        RECT 69.250 120.315 69.420 121.155 ;
        RECT 69.590 121.445 70.055 121.775 ;
        RECT 70.440 121.715 70.610 121.945 ;
        RECT 70.790 121.895 71.160 122.395 ;
        RECT 71.480 121.945 72.155 122.115 ;
        RECT 72.350 121.945 72.685 122.115 ;
        RECT 69.590 120.485 69.910 121.445 ;
        RECT 70.440 121.415 71.270 121.715 ;
        RECT 70.080 120.515 70.270 121.235 ;
        RECT 70.440 120.345 70.610 121.415 ;
        RECT 71.070 121.385 71.270 121.415 ;
        RECT 70.780 121.165 70.950 121.235 ;
        RECT 71.480 121.165 71.650 121.945 ;
        RECT 72.515 121.805 72.685 121.945 ;
        RECT 72.855 121.935 73.105 122.395 ;
        RECT 70.780 120.995 71.650 121.165 ;
        RECT 71.820 121.525 72.345 121.745 ;
        RECT 72.515 121.675 72.740 121.805 ;
        RECT 70.780 120.905 71.290 120.995 ;
        RECT 69.250 120.145 70.135 120.315 ;
        RECT 70.360 120.015 70.610 120.345 ;
        RECT 70.780 119.845 70.950 120.645 ;
        RECT 71.120 120.290 71.290 120.905 ;
        RECT 71.820 120.825 71.990 121.525 ;
        RECT 71.460 120.460 71.990 120.825 ;
        RECT 72.160 120.760 72.400 121.355 ;
        RECT 72.570 120.570 72.740 121.675 ;
        RECT 72.910 120.815 73.190 121.765 ;
        RECT 72.435 120.440 72.740 120.570 ;
        RECT 71.120 120.120 72.225 120.290 ;
        RECT 72.435 120.015 72.685 120.440 ;
        RECT 72.855 119.845 73.120 120.305 ;
        RECT 73.360 120.015 73.545 122.135 ;
        RECT 73.715 122.015 74.045 122.395 ;
        RECT 74.215 121.845 74.385 122.135 ;
        RECT 74.645 121.850 79.990 122.395 ;
        RECT 80.165 121.850 85.510 122.395 ;
        RECT 73.720 121.675 74.385 121.845 ;
        RECT 73.720 120.685 73.950 121.675 ;
        RECT 74.120 120.855 74.470 121.505 ;
        RECT 76.230 121.020 76.570 121.850 ;
        RECT 73.720 120.515 74.385 120.685 ;
        RECT 73.715 119.845 74.045 120.345 ;
        RECT 74.215 120.015 74.385 120.515 ;
        RECT 78.050 120.280 78.400 121.530 ;
        RECT 81.750 121.020 82.090 121.850 ;
        RECT 85.685 121.625 89.195 122.395 ;
        RECT 89.365 121.645 90.575 122.395 ;
        RECT 90.745 121.645 91.955 122.395 ;
        RECT 100.140 122.350 106.380 122.450 ;
        RECT 83.570 120.280 83.920 121.530 ;
        RECT 85.685 121.105 87.335 121.625 ;
        RECT 87.505 120.935 89.195 121.455 ;
        RECT 89.365 121.105 89.885 121.645 ;
        RECT 90.055 120.935 90.575 121.475 ;
        RECT 74.645 119.845 79.990 120.280 ;
        RECT 80.165 119.845 85.510 120.280 ;
        RECT 85.685 119.845 89.195 120.935 ;
        RECT 89.365 119.845 90.575 120.935 ;
        RECT 90.745 120.935 91.265 121.475 ;
        RECT 91.435 121.105 91.955 121.645 ;
        RECT 100.130 121.790 106.380 122.350 ;
        RECT 100.130 121.770 105.300 121.790 ;
        RECT 100.130 121.700 104.120 121.770 ;
        RECT 90.745 119.845 91.955 120.935 ;
        RECT 100.130 120.430 102.050 121.700 ;
        RECT 103.560 121.690 104.120 121.700 ;
        RECT 103.790 120.600 104.120 121.690 ;
        RECT 104.490 121.220 105.530 121.390 ;
        RECT 104.490 120.780 105.530 120.950 ;
        RECT 105.700 120.920 105.870 121.250 ;
        RECT 103.950 120.380 104.120 120.600 ;
        RECT 106.210 120.380 106.380 121.790 ;
        RECT 103.950 120.210 106.380 120.380 ;
        RECT 107.960 122.300 118.590 122.470 ;
        RECT 120.020 131.640 126.250 131.800 ;
        RECT 120.020 129.380 120.690 131.640 ;
        RECT 121.360 131.070 125.400 131.240 ;
        RECT 121.020 130.010 121.190 131.010 ;
        RECT 125.570 130.010 125.740 131.010 ;
        RECT 121.360 129.780 125.400 129.950 ;
        RECT 126.080 129.380 126.250 131.640 ;
        RECT 120.020 129.210 126.250 129.380 ;
        RECT 120.020 125.950 120.690 129.210 ;
        RECT 121.360 128.640 125.400 128.810 ;
        RECT 121.020 126.580 121.190 128.580 ;
        RECT 125.570 126.580 125.740 128.580 ;
        RECT 121.360 126.350 125.400 126.520 ;
        RECT 126.080 125.950 126.250 129.210 ;
        RECT 120.020 125.780 126.250 125.950 ;
        RECT 120.020 122.520 120.690 125.780 ;
        RECT 121.360 125.210 125.400 125.380 ;
        RECT 121.020 123.150 121.190 125.150 ;
        RECT 125.570 123.150 125.740 125.150 ;
        RECT 121.360 122.920 125.400 123.090 ;
        RECT 126.080 122.520 126.250 125.780 ;
        RECT 120.020 122.510 126.250 122.520 ;
        RECT 127.840 131.780 137.670 131.820 ;
        RECT 140.540 131.800 146.280 131.810 ;
        RECT 127.840 131.650 138.470 131.780 ;
        RECT 127.840 129.390 128.010 131.650 ;
        RECT 128.735 131.080 136.775 131.250 ;
        RECT 128.350 130.020 128.520 131.020 ;
        RECT 136.990 130.020 137.160 131.020 ;
        RECT 128.735 129.790 136.775 129.960 ;
        RECT 137.500 129.390 138.470 131.650 ;
        RECT 127.840 129.220 138.470 129.390 ;
        RECT 127.840 125.960 128.010 129.220 ;
        RECT 128.735 128.650 136.775 128.820 ;
        RECT 128.350 126.590 128.520 128.590 ;
        RECT 136.990 126.590 137.160 128.590 ;
        RECT 128.735 126.360 136.775 126.530 ;
        RECT 137.500 125.960 138.470 129.220 ;
        RECT 127.840 125.790 138.470 125.960 ;
        RECT 127.840 122.530 128.010 125.790 ;
        RECT 128.735 125.220 136.775 125.390 ;
        RECT 128.350 123.160 128.520 125.160 ;
        RECT 136.990 123.160 137.160 125.160 ;
        RECT 128.735 122.930 136.775 123.100 ;
        RECT 137.500 122.530 138.470 125.790 ;
        RECT 120.020 122.410 126.260 122.510 ;
        RECT 107.960 120.040 108.130 122.300 ;
        RECT 108.855 121.730 116.895 121.900 ;
        RECT 108.470 120.670 108.640 121.670 ;
        RECT 117.110 120.670 117.280 121.670 ;
        RECT 108.855 120.440 116.895 120.610 ;
        RECT 117.620 120.040 118.590 122.300 ;
        RECT 120.010 121.850 126.260 122.410 ;
        RECT 120.010 121.830 125.180 121.850 ;
        RECT 120.010 121.760 124.000 121.830 ;
        RECT 120.010 120.490 121.930 121.760 ;
        RECT 123.440 121.750 124.000 121.760 ;
        RECT 123.670 120.660 124.000 121.750 ;
        RECT 124.370 121.280 125.410 121.450 ;
        RECT 124.370 120.840 125.410 121.010 ;
        RECT 125.580 120.980 125.750 121.310 ;
        RECT 123.830 120.440 124.000 120.660 ;
        RECT 126.090 120.440 126.260 121.850 ;
        RECT 123.830 120.270 126.260 120.440 ;
        RECT 127.840 122.360 138.470 122.530 ;
        RECT 140.050 131.640 146.280 131.800 ;
        RECT 140.050 129.380 140.720 131.640 ;
        RECT 141.390 131.070 145.430 131.240 ;
        RECT 141.050 130.010 141.220 131.010 ;
        RECT 145.600 130.010 145.770 131.010 ;
        RECT 141.390 129.780 145.430 129.950 ;
        RECT 146.110 129.380 146.280 131.640 ;
        RECT 140.050 129.210 146.280 129.380 ;
        RECT 140.050 125.950 140.720 129.210 ;
        RECT 141.390 128.640 145.430 128.810 ;
        RECT 141.050 126.580 141.220 128.580 ;
        RECT 145.600 126.580 145.770 128.580 ;
        RECT 141.390 126.350 145.430 126.520 ;
        RECT 146.110 125.950 146.280 129.210 ;
        RECT 140.050 125.780 146.280 125.950 ;
        RECT 140.050 122.520 140.720 125.780 ;
        RECT 141.390 125.210 145.430 125.380 ;
        RECT 141.050 123.150 141.220 125.150 ;
        RECT 145.600 123.150 145.770 125.150 ;
        RECT 141.390 122.920 145.430 123.090 ;
        RECT 146.110 122.520 146.280 125.780 ;
        RECT 140.050 122.510 146.280 122.520 ;
        RECT 147.870 131.780 157.700 131.820 ;
        RECT 147.870 131.650 158.500 131.780 ;
        RECT 147.870 129.390 148.040 131.650 ;
        RECT 148.765 131.080 156.805 131.250 ;
        RECT 148.380 130.020 148.550 131.020 ;
        RECT 157.020 130.020 157.190 131.020 ;
        RECT 148.765 129.790 156.805 129.960 ;
        RECT 157.530 129.390 158.500 131.650 ;
        RECT 147.870 129.220 158.500 129.390 ;
        RECT 147.870 125.960 148.040 129.220 ;
        RECT 148.765 128.650 156.805 128.820 ;
        RECT 148.380 126.590 148.550 128.590 ;
        RECT 157.020 126.590 157.190 128.590 ;
        RECT 148.765 126.360 156.805 126.530 ;
        RECT 157.530 125.960 158.500 129.220 ;
        RECT 147.870 125.790 158.500 125.960 ;
        RECT 147.870 122.530 148.040 125.790 ;
        RECT 148.765 125.220 156.805 125.390 ;
        RECT 148.380 123.160 148.550 125.160 ;
        RECT 157.020 123.160 157.190 125.160 ;
        RECT 148.765 122.930 156.805 123.100 ;
        RECT 157.530 122.530 158.500 125.790 ;
        RECT 140.050 122.410 146.290 122.510 ;
        RECT 127.840 120.100 128.010 122.360 ;
        RECT 128.735 121.790 136.775 121.960 ;
        RECT 128.350 120.730 128.520 121.730 ;
        RECT 136.990 120.730 137.160 121.730 ;
        RECT 128.735 120.500 136.775 120.670 ;
        RECT 137.500 120.100 138.470 122.360 ;
        RECT 140.040 121.850 146.290 122.410 ;
        RECT 140.040 121.830 145.210 121.850 ;
        RECT 140.040 121.760 144.030 121.830 ;
        RECT 140.040 120.490 141.960 121.760 ;
        RECT 143.470 121.750 144.030 121.760 ;
        RECT 143.700 120.660 144.030 121.750 ;
        RECT 144.400 121.280 145.440 121.450 ;
        RECT 144.400 120.840 145.440 121.010 ;
        RECT 145.610 120.980 145.780 121.310 ;
        RECT 143.860 120.440 144.030 120.660 ;
        RECT 146.120 120.440 146.290 121.850 ;
        RECT 143.860 120.270 146.290 120.440 ;
        RECT 147.870 122.360 158.500 122.530 ;
        RECT 127.840 120.070 138.470 120.100 ;
        RECT 147.870 120.100 148.040 122.360 ;
        RECT 148.765 121.790 156.805 121.960 ;
        RECT 148.380 120.730 148.550 121.730 ;
        RECT 157.020 120.730 157.190 121.730 ;
        RECT 148.765 120.500 156.805 120.670 ;
        RECT 157.530 120.100 158.500 122.360 ;
        RECT 147.870 120.070 158.500 120.100 ;
        RECT 107.960 120.010 118.590 120.040 ;
        RECT 107.930 119.900 118.590 120.010 ;
        RECT 127.810 119.960 138.470 120.070 ;
        RECT 147.840 119.960 158.500 120.070 ;
        RECT 126.060 119.910 138.470 119.960 ;
        RECT 146.090 119.910 158.500 119.960 ;
        RECT 106.180 119.850 118.590 119.900 ;
        RECT 13.380 119.675 92.040 119.845 ;
        RECT 101.840 119.680 118.590 119.850 ;
        RECT 13.465 118.585 14.675 119.675 ;
        RECT 14.845 118.585 16.055 119.675 ;
        RECT 16.285 118.615 16.615 119.460 ;
        RECT 16.785 118.665 16.955 119.675 ;
        RECT 17.125 118.945 17.465 119.505 ;
        RECT 17.695 119.175 18.010 119.675 ;
        RECT 18.190 119.205 19.075 119.375 ;
        RECT 13.465 117.875 13.985 118.415 ;
        RECT 14.155 118.045 14.675 118.585 ;
        RECT 14.845 117.875 15.365 118.415 ;
        RECT 15.535 118.045 16.055 118.585 ;
        RECT 16.225 118.535 16.615 118.615 ;
        RECT 17.125 118.570 18.020 118.945 ;
        RECT 16.225 118.485 16.440 118.535 ;
        RECT 16.225 117.905 16.395 118.485 ;
        RECT 17.125 118.365 17.315 118.570 ;
        RECT 18.190 118.365 18.360 119.205 ;
        RECT 19.300 119.175 19.550 119.505 ;
        RECT 16.565 118.035 17.315 118.365 ;
        RECT 17.485 118.035 18.360 118.365 ;
        RECT 13.465 117.125 14.675 117.875 ;
        RECT 14.845 117.125 16.055 117.875 ;
        RECT 16.225 117.865 16.450 117.905 ;
        RECT 17.115 117.865 17.315 118.035 ;
        RECT 16.225 117.780 16.605 117.865 ;
        RECT 16.275 117.345 16.605 117.780 ;
        RECT 16.775 117.125 16.945 117.735 ;
        RECT 17.115 117.340 17.445 117.865 ;
        RECT 17.705 117.125 17.915 117.655 ;
        RECT 18.190 117.575 18.360 118.035 ;
        RECT 18.530 118.075 18.850 119.035 ;
        RECT 19.020 118.285 19.210 119.005 ;
        RECT 19.380 118.105 19.550 119.175 ;
        RECT 19.720 118.875 19.890 119.675 ;
        RECT 20.060 119.230 21.165 119.400 ;
        RECT 20.060 118.615 20.230 119.230 ;
        RECT 21.375 119.080 21.625 119.505 ;
        RECT 21.795 119.215 22.060 119.675 ;
        RECT 20.400 118.695 20.930 119.060 ;
        RECT 21.375 118.950 21.680 119.080 ;
        RECT 19.720 118.525 20.230 118.615 ;
        RECT 19.720 118.355 20.590 118.525 ;
        RECT 19.720 118.285 19.890 118.355 ;
        RECT 20.010 118.105 20.210 118.135 ;
        RECT 18.530 117.745 18.995 118.075 ;
        RECT 19.380 117.805 20.210 118.105 ;
        RECT 19.380 117.575 19.550 117.805 ;
        RECT 18.190 117.405 18.975 117.575 ;
        RECT 19.145 117.405 19.550 117.575 ;
        RECT 19.730 117.125 20.100 117.625 ;
        RECT 20.420 117.575 20.590 118.355 ;
        RECT 20.760 117.995 20.930 118.695 ;
        RECT 21.100 118.165 21.340 118.760 ;
        RECT 20.760 117.775 21.285 117.995 ;
        RECT 21.510 117.845 21.680 118.950 ;
        RECT 21.455 117.715 21.680 117.845 ;
        RECT 21.850 117.755 22.130 118.705 ;
        RECT 21.455 117.575 21.625 117.715 ;
        RECT 20.420 117.405 21.095 117.575 ;
        RECT 21.290 117.405 21.625 117.575 ;
        RECT 21.795 117.125 22.045 117.585 ;
        RECT 22.300 117.385 22.485 119.505 ;
        RECT 22.655 119.175 22.985 119.675 ;
        RECT 23.155 119.005 23.325 119.505 ;
        RECT 22.660 118.835 23.325 119.005 ;
        RECT 22.660 117.845 22.890 118.835 ;
        RECT 23.060 118.015 23.410 118.665 ;
        RECT 23.585 118.070 23.865 119.505 ;
        RECT 24.035 118.900 24.745 119.675 ;
        RECT 24.915 118.730 25.245 119.505 ;
        RECT 24.095 118.515 25.245 118.730 ;
        RECT 22.660 117.675 23.325 117.845 ;
        RECT 22.655 117.125 22.985 117.505 ;
        RECT 23.155 117.385 23.325 117.675 ;
        RECT 23.585 117.295 23.925 118.070 ;
        RECT 24.095 117.945 24.380 118.515 ;
        RECT 24.565 118.115 25.035 118.345 ;
        RECT 25.440 118.315 25.655 119.430 ;
        RECT 25.835 118.955 26.165 119.675 ;
        RECT 25.945 118.315 26.175 118.655 ;
        RECT 26.345 118.510 26.635 119.675 ;
        RECT 26.895 119.005 27.065 119.505 ;
        RECT 27.235 119.175 27.565 119.675 ;
        RECT 26.895 118.835 27.560 119.005 ;
        RECT 25.205 118.135 25.655 118.315 ;
        RECT 25.205 118.115 25.535 118.135 ;
        RECT 25.845 118.115 26.175 118.315 ;
        RECT 26.810 118.015 27.160 118.665 ;
        RECT 24.095 117.755 24.805 117.945 ;
        RECT 24.505 117.615 24.805 117.755 ;
        RECT 24.995 117.755 26.175 117.945 ;
        RECT 24.995 117.675 25.325 117.755 ;
        RECT 24.505 117.605 24.820 117.615 ;
        RECT 24.505 117.595 24.830 117.605 ;
        RECT 24.505 117.590 24.840 117.595 ;
        RECT 24.095 117.125 24.265 117.585 ;
        RECT 24.505 117.580 24.845 117.590 ;
        RECT 24.505 117.575 24.850 117.580 ;
        RECT 24.505 117.565 24.855 117.575 ;
        RECT 24.505 117.560 24.860 117.565 ;
        RECT 24.505 117.295 24.865 117.560 ;
        RECT 25.495 117.125 25.665 117.585 ;
        RECT 25.835 117.295 26.175 117.755 ;
        RECT 26.345 117.125 26.635 117.850 ;
        RECT 27.330 117.845 27.560 118.835 ;
        RECT 26.895 117.675 27.560 117.845 ;
        RECT 26.895 117.385 27.065 117.675 ;
        RECT 27.235 117.125 27.565 117.505 ;
        RECT 27.735 117.385 27.920 119.505 ;
        RECT 28.160 119.215 28.425 119.675 ;
        RECT 28.595 119.080 28.845 119.505 ;
        RECT 29.055 119.230 30.160 119.400 ;
        RECT 28.540 118.950 28.845 119.080 ;
        RECT 28.090 117.755 28.370 118.705 ;
        RECT 28.540 117.845 28.710 118.950 ;
        RECT 28.880 118.165 29.120 118.760 ;
        RECT 29.290 118.695 29.820 119.060 ;
        RECT 29.290 117.995 29.460 118.695 ;
        RECT 29.990 118.615 30.160 119.230 ;
        RECT 30.330 118.875 30.500 119.675 ;
        RECT 30.670 119.175 30.920 119.505 ;
        RECT 31.145 119.205 32.030 119.375 ;
        RECT 29.990 118.525 30.500 118.615 ;
        RECT 28.540 117.715 28.765 117.845 ;
        RECT 28.935 117.775 29.460 117.995 ;
        RECT 29.630 118.355 30.500 118.525 ;
        RECT 28.175 117.125 28.425 117.585 ;
        RECT 28.595 117.575 28.765 117.715 ;
        RECT 29.630 117.575 29.800 118.355 ;
        RECT 30.330 118.285 30.500 118.355 ;
        RECT 30.010 118.105 30.210 118.135 ;
        RECT 30.670 118.105 30.840 119.175 ;
        RECT 31.010 118.285 31.200 119.005 ;
        RECT 30.010 117.805 30.840 118.105 ;
        RECT 31.370 118.075 31.690 119.035 ;
        RECT 28.595 117.405 28.930 117.575 ;
        RECT 29.125 117.405 29.800 117.575 ;
        RECT 30.120 117.125 30.490 117.625 ;
        RECT 30.670 117.575 30.840 117.805 ;
        RECT 31.225 117.745 31.690 118.075 ;
        RECT 31.860 118.365 32.030 119.205 ;
        RECT 32.210 119.175 32.525 119.675 ;
        RECT 32.755 118.945 33.095 119.505 ;
        RECT 32.200 118.570 33.095 118.945 ;
        RECT 33.265 118.665 33.435 119.675 ;
        RECT 32.905 118.365 33.095 118.570 ;
        RECT 33.605 118.615 33.935 119.460 ;
        RECT 33.605 118.535 33.995 118.615 ;
        RECT 33.780 118.485 33.995 118.535 ;
        RECT 31.860 118.035 32.735 118.365 ;
        RECT 32.905 118.035 33.655 118.365 ;
        RECT 31.860 117.575 32.030 118.035 ;
        RECT 32.905 117.865 33.105 118.035 ;
        RECT 33.825 117.905 33.995 118.485 ;
        RECT 33.770 117.865 33.995 117.905 ;
        RECT 30.670 117.405 31.075 117.575 ;
        RECT 31.245 117.405 32.030 117.575 ;
        RECT 32.305 117.125 32.515 117.655 ;
        RECT 32.775 117.340 33.105 117.865 ;
        RECT 33.615 117.780 33.995 117.865 ;
        RECT 34.165 118.535 34.550 119.505 ;
        RECT 34.720 119.215 35.045 119.675 ;
        RECT 35.565 119.045 35.845 119.505 ;
        RECT 34.720 118.825 35.845 119.045 ;
        RECT 34.165 117.865 34.445 118.535 ;
        RECT 34.720 118.365 35.170 118.825 ;
        RECT 36.035 118.655 36.435 119.505 ;
        RECT 36.835 119.215 37.105 119.675 ;
        RECT 37.275 119.045 37.560 119.505 ;
        RECT 34.615 118.035 35.170 118.365 ;
        RECT 35.340 118.095 36.435 118.655 ;
        RECT 34.720 117.925 35.170 118.035 ;
        RECT 33.275 117.125 33.445 117.735 ;
        RECT 33.615 117.345 33.945 117.780 ;
        RECT 34.165 117.295 34.550 117.865 ;
        RECT 34.720 117.755 35.845 117.925 ;
        RECT 34.720 117.125 35.045 117.585 ;
        RECT 35.565 117.295 35.845 117.755 ;
        RECT 36.035 117.295 36.435 118.095 ;
        RECT 36.605 118.825 37.560 119.045 ;
        RECT 36.605 117.925 36.815 118.825 ;
        RECT 36.985 118.095 37.675 118.655 ;
        RECT 38.305 118.535 38.690 119.505 ;
        RECT 38.860 119.215 39.185 119.675 ;
        RECT 39.705 119.045 39.985 119.505 ;
        RECT 38.860 118.825 39.985 119.045 ;
        RECT 36.605 117.755 37.560 117.925 ;
        RECT 36.835 117.125 37.105 117.585 ;
        RECT 37.275 117.295 37.560 117.755 ;
        RECT 38.305 117.865 38.585 118.535 ;
        RECT 38.860 118.365 39.310 118.825 ;
        RECT 40.175 118.655 40.575 119.505 ;
        RECT 40.975 119.215 41.245 119.675 ;
        RECT 41.415 119.045 41.700 119.505 ;
        RECT 41.985 119.240 47.330 119.675 ;
        RECT 38.755 118.035 39.310 118.365 ;
        RECT 39.480 118.095 40.575 118.655 ;
        RECT 38.860 117.925 39.310 118.035 ;
        RECT 38.305 117.295 38.690 117.865 ;
        RECT 38.860 117.755 39.985 117.925 ;
        RECT 38.860 117.125 39.185 117.585 ;
        RECT 39.705 117.295 39.985 117.755 ;
        RECT 40.175 117.295 40.575 118.095 ;
        RECT 40.745 118.825 41.700 119.045 ;
        RECT 40.745 117.925 40.955 118.825 ;
        RECT 41.125 118.095 41.815 118.655 ;
        RECT 40.745 117.755 41.700 117.925 ;
        RECT 40.975 117.125 41.245 117.585 ;
        RECT 41.415 117.295 41.700 117.755 ;
        RECT 43.570 117.670 43.910 118.500 ;
        RECT 45.390 117.990 45.740 119.240 ;
        RECT 47.505 118.585 51.015 119.675 ;
        RECT 47.505 117.895 49.155 118.415 ;
        RECT 49.325 118.065 51.015 118.585 ;
        RECT 52.105 118.510 52.395 119.675 ;
        RECT 52.655 119.005 52.825 119.505 ;
        RECT 52.995 119.175 53.325 119.675 ;
        RECT 52.655 118.835 53.320 119.005 ;
        RECT 52.570 118.015 52.920 118.665 ;
        RECT 41.985 117.125 47.330 117.670 ;
        RECT 47.505 117.125 51.015 117.895 ;
        RECT 52.105 117.125 52.395 117.850 ;
        RECT 53.090 117.845 53.320 118.835 ;
        RECT 52.655 117.675 53.320 117.845 ;
        RECT 52.655 117.385 52.825 117.675 ;
        RECT 52.995 117.125 53.325 117.505 ;
        RECT 53.495 117.385 53.680 119.505 ;
        RECT 53.920 119.215 54.185 119.675 ;
        RECT 54.355 119.080 54.605 119.505 ;
        RECT 54.815 119.230 55.920 119.400 ;
        RECT 54.300 118.950 54.605 119.080 ;
        RECT 53.850 117.755 54.130 118.705 ;
        RECT 54.300 117.845 54.470 118.950 ;
        RECT 54.640 118.165 54.880 118.760 ;
        RECT 55.050 118.695 55.580 119.060 ;
        RECT 55.050 117.995 55.220 118.695 ;
        RECT 55.750 118.615 55.920 119.230 ;
        RECT 56.090 118.875 56.260 119.675 ;
        RECT 56.430 119.175 56.680 119.505 ;
        RECT 56.905 119.205 57.790 119.375 ;
        RECT 55.750 118.525 56.260 118.615 ;
        RECT 54.300 117.715 54.525 117.845 ;
        RECT 54.695 117.775 55.220 117.995 ;
        RECT 55.390 118.355 56.260 118.525 ;
        RECT 53.935 117.125 54.185 117.585 ;
        RECT 54.355 117.575 54.525 117.715 ;
        RECT 55.390 117.575 55.560 118.355 ;
        RECT 56.090 118.285 56.260 118.355 ;
        RECT 55.770 118.105 55.970 118.135 ;
        RECT 56.430 118.105 56.600 119.175 ;
        RECT 56.770 118.285 56.960 119.005 ;
        RECT 55.770 117.805 56.600 118.105 ;
        RECT 57.130 118.075 57.450 119.035 ;
        RECT 54.355 117.405 54.690 117.575 ;
        RECT 54.885 117.405 55.560 117.575 ;
        RECT 55.880 117.125 56.250 117.625 ;
        RECT 56.430 117.575 56.600 117.805 ;
        RECT 56.985 117.745 57.450 118.075 ;
        RECT 57.620 118.365 57.790 119.205 ;
        RECT 57.970 119.175 58.285 119.675 ;
        RECT 58.515 118.945 58.855 119.505 ;
        RECT 57.960 118.570 58.855 118.945 ;
        RECT 59.025 118.665 59.195 119.675 ;
        RECT 58.665 118.365 58.855 118.570 ;
        RECT 59.365 118.615 59.695 119.460 ;
        RECT 60.475 119.005 60.645 119.505 ;
        RECT 60.815 119.175 61.145 119.675 ;
        RECT 60.475 118.835 61.140 119.005 ;
        RECT 59.365 118.535 59.755 118.615 ;
        RECT 59.540 118.485 59.755 118.535 ;
        RECT 57.620 118.035 58.495 118.365 ;
        RECT 58.665 118.035 59.415 118.365 ;
        RECT 57.620 117.575 57.790 118.035 ;
        RECT 58.665 117.865 58.865 118.035 ;
        RECT 59.585 117.905 59.755 118.485 ;
        RECT 60.390 118.015 60.740 118.665 ;
        RECT 59.530 117.865 59.755 117.905 ;
        RECT 56.430 117.405 56.835 117.575 ;
        RECT 57.005 117.405 57.790 117.575 ;
        RECT 58.065 117.125 58.275 117.655 ;
        RECT 58.535 117.340 58.865 117.865 ;
        RECT 59.375 117.780 59.755 117.865 ;
        RECT 60.910 117.845 61.140 118.835 ;
        RECT 59.035 117.125 59.205 117.735 ;
        RECT 59.375 117.345 59.705 117.780 ;
        RECT 60.475 117.675 61.140 117.845 ;
        RECT 60.475 117.385 60.645 117.675 ;
        RECT 60.815 117.125 61.145 117.505 ;
        RECT 61.315 117.385 61.500 119.505 ;
        RECT 61.740 119.215 62.005 119.675 ;
        RECT 62.175 119.080 62.425 119.505 ;
        RECT 62.635 119.230 63.740 119.400 ;
        RECT 62.120 118.950 62.425 119.080 ;
        RECT 61.670 117.755 61.950 118.705 ;
        RECT 62.120 117.845 62.290 118.950 ;
        RECT 62.460 118.165 62.700 118.760 ;
        RECT 62.870 118.695 63.400 119.060 ;
        RECT 62.870 117.995 63.040 118.695 ;
        RECT 63.570 118.615 63.740 119.230 ;
        RECT 63.910 118.875 64.080 119.675 ;
        RECT 64.250 119.175 64.500 119.505 ;
        RECT 64.725 119.205 65.610 119.375 ;
        RECT 63.570 118.525 64.080 118.615 ;
        RECT 62.120 117.715 62.345 117.845 ;
        RECT 62.515 117.775 63.040 117.995 ;
        RECT 63.210 118.355 64.080 118.525 ;
        RECT 61.755 117.125 62.005 117.585 ;
        RECT 62.175 117.575 62.345 117.715 ;
        RECT 63.210 117.575 63.380 118.355 ;
        RECT 63.910 118.285 64.080 118.355 ;
        RECT 63.590 118.105 63.790 118.135 ;
        RECT 64.250 118.105 64.420 119.175 ;
        RECT 64.590 118.285 64.780 119.005 ;
        RECT 63.590 117.805 64.420 118.105 ;
        RECT 64.950 118.075 65.270 119.035 ;
        RECT 62.175 117.405 62.510 117.575 ;
        RECT 62.705 117.405 63.380 117.575 ;
        RECT 63.700 117.125 64.070 117.625 ;
        RECT 64.250 117.575 64.420 117.805 ;
        RECT 64.805 117.745 65.270 118.075 ;
        RECT 65.440 118.365 65.610 119.205 ;
        RECT 65.790 119.175 66.105 119.675 ;
        RECT 66.335 118.945 66.675 119.505 ;
        RECT 65.780 118.570 66.675 118.945 ;
        RECT 66.845 118.665 67.015 119.675 ;
        RECT 66.485 118.365 66.675 118.570 ;
        RECT 67.185 118.615 67.515 119.460 ;
        RECT 67.185 118.535 67.575 118.615 ;
        RECT 67.360 118.485 67.575 118.535 ;
        RECT 65.440 118.035 66.315 118.365 ;
        RECT 66.485 118.035 67.235 118.365 ;
        RECT 65.440 117.575 65.610 118.035 ;
        RECT 66.485 117.865 66.685 118.035 ;
        RECT 67.405 117.905 67.575 118.485 ;
        RECT 67.350 117.865 67.575 117.905 ;
        RECT 64.250 117.405 64.655 117.575 ;
        RECT 64.825 117.405 65.610 117.575 ;
        RECT 65.885 117.125 66.095 117.655 ;
        RECT 66.355 117.340 66.685 117.865 ;
        RECT 67.195 117.780 67.575 117.865 ;
        RECT 67.745 118.535 68.130 119.505 ;
        RECT 68.300 119.215 68.625 119.675 ;
        RECT 69.145 119.045 69.425 119.505 ;
        RECT 68.300 118.825 69.425 119.045 ;
        RECT 67.745 117.865 68.025 118.535 ;
        RECT 68.300 118.365 68.750 118.825 ;
        RECT 69.615 118.655 70.015 119.505 ;
        RECT 70.415 119.215 70.685 119.675 ;
        RECT 70.855 119.045 71.140 119.505 ;
        RECT 68.195 118.035 68.750 118.365 ;
        RECT 68.920 118.095 70.015 118.655 ;
        RECT 68.300 117.925 68.750 118.035 ;
        RECT 66.855 117.125 67.025 117.735 ;
        RECT 67.195 117.345 67.525 117.780 ;
        RECT 67.745 117.295 68.130 117.865 ;
        RECT 68.300 117.755 69.425 117.925 ;
        RECT 68.300 117.125 68.625 117.585 ;
        RECT 69.145 117.295 69.425 117.755 ;
        RECT 69.615 117.295 70.015 118.095 ;
        RECT 70.185 118.825 71.140 119.045 ;
        RECT 71.430 119.285 71.765 119.505 ;
        RECT 72.770 119.295 73.125 119.675 ;
        RECT 70.185 117.925 70.395 118.825 ;
        RECT 71.430 118.665 71.685 119.285 ;
        RECT 71.935 119.125 72.165 119.165 ;
        RECT 73.295 119.125 73.545 119.505 ;
        RECT 71.935 118.925 73.545 119.125 ;
        RECT 71.935 118.835 72.120 118.925 ;
        RECT 72.710 118.915 73.545 118.925 ;
        RECT 73.795 118.895 74.045 119.675 ;
        RECT 74.215 118.825 74.475 119.505 ;
        RECT 72.275 118.725 72.605 118.755 ;
        RECT 72.275 118.665 74.075 118.725 ;
        RECT 70.565 118.095 71.255 118.655 ;
        RECT 71.430 118.555 74.135 118.665 ;
        RECT 71.430 118.495 72.605 118.555 ;
        RECT 73.935 118.520 74.135 118.555 ;
        RECT 71.425 118.115 71.915 118.315 ;
        RECT 72.105 118.115 72.580 118.325 ;
        RECT 70.185 117.755 71.140 117.925 ;
        RECT 70.415 117.125 70.685 117.585 ;
        RECT 70.855 117.295 71.140 117.755 ;
        RECT 71.430 117.125 71.885 117.890 ;
        RECT 72.360 117.715 72.580 118.115 ;
        RECT 72.825 118.115 73.155 118.325 ;
        RECT 72.825 117.715 73.035 118.115 ;
        RECT 73.325 118.080 73.735 118.385 ;
        RECT 73.965 117.945 74.135 118.520 ;
        RECT 73.865 117.825 74.135 117.945 ;
        RECT 73.290 117.780 74.135 117.825 ;
        RECT 73.290 117.655 74.045 117.780 ;
        RECT 73.290 117.505 73.460 117.655 ;
        RECT 74.305 117.625 74.475 118.825 ;
        RECT 74.645 118.585 77.235 119.675 ;
        RECT 72.160 117.295 73.460 117.505 ;
        RECT 73.715 117.125 74.045 117.485 ;
        RECT 74.215 117.295 74.475 117.625 ;
        RECT 74.645 117.895 75.855 118.415 ;
        RECT 76.025 118.065 77.235 118.585 ;
        RECT 77.865 118.510 78.155 119.675 ;
        RECT 78.325 119.240 83.670 119.675 ;
        RECT 83.845 119.240 89.190 119.675 ;
        RECT 74.645 117.125 77.235 117.895 ;
        RECT 77.865 117.125 78.155 117.850 ;
        RECT 79.910 117.670 80.250 118.500 ;
        RECT 81.730 117.990 82.080 119.240 ;
        RECT 85.430 117.670 85.770 118.500 ;
        RECT 87.250 117.990 87.600 119.240 ;
        RECT 89.365 118.585 90.575 119.675 ;
        RECT 89.365 117.875 89.885 118.415 ;
        RECT 90.055 118.045 90.575 118.585 ;
        RECT 90.745 118.585 91.955 119.675 ;
        RECT 90.745 118.045 91.265 118.585 ;
        RECT 91.435 117.875 91.955 118.415 ;
        RECT 101.840 118.270 102.010 119.680 ;
        RECT 102.380 119.110 105.420 119.280 ;
        RECT 102.380 118.670 105.420 118.840 ;
        RECT 105.635 118.810 105.805 119.140 ;
        RECT 106.140 118.920 118.590 119.680 ;
        RECT 121.720 119.740 138.470 119.910 ;
        RECT 106.140 118.910 118.480 118.920 ;
        RECT 106.140 118.900 112.020 118.910 ;
        RECT 106.140 118.880 106.710 118.900 ;
        RECT 107.930 118.890 112.020 118.900 ;
        RECT 106.150 118.270 106.320 118.880 ;
        RECT 101.840 118.100 106.320 118.270 ;
        RECT 121.720 118.330 121.890 119.740 ;
        RECT 122.260 119.170 125.300 119.340 ;
        RECT 122.260 118.730 125.300 118.900 ;
        RECT 125.515 118.870 125.685 119.200 ;
        RECT 126.020 118.980 138.470 119.740 ;
        RECT 141.750 119.740 158.500 119.910 ;
        RECT 126.020 118.970 138.360 118.980 ;
        RECT 126.020 118.960 131.900 118.970 ;
        RECT 126.020 118.940 126.590 118.960 ;
        RECT 127.810 118.950 131.900 118.960 ;
        RECT 126.030 118.330 126.200 118.940 ;
        RECT 121.720 118.160 126.200 118.330 ;
        RECT 141.750 118.330 141.920 119.740 ;
        RECT 142.290 119.170 145.330 119.340 ;
        RECT 142.290 118.730 145.330 118.900 ;
        RECT 145.545 118.870 145.715 119.200 ;
        RECT 146.050 118.980 158.500 119.740 ;
        RECT 146.050 118.970 158.390 118.980 ;
        RECT 146.050 118.960 151.930 118.970 ;
        RECT 146.050 118.940 146.620 118.960 ;
        RECT 147.840 118.950 151.930 118.960 ;
        RECT 146.060 118.330 146.230 118.940 ;
        RECT 141.750 118.160 146.230 118.330 ;
        RECT 78.325 117.125 83.670 117.670 ;
        RECT 83.845 117.125 89.190 117.670 ;
        RECT 89.365 117.125 90.575 117.875 ;
        RECT 90.745 117.125 91.955 117.875 ;
        RECT 13.380 116.955 92.040 117.125 ;
        RECT 13.465 116.205 14.675 116.955 ;
        RECT 14.845 116.455 15.105 116.785 ;
        RECT 15.315 116.475 15.590 116.955 ;
        RECT 13.465 115.665 13.985 116.205 ;
        RECT 14.155 115.495 14.675 116.035 ;
        RECT 13.465 114.405 14.675 115.495 ;
        RECT 14.845 115.545 15.015 116.455 ;
        RECT 15.800 116.385 16.005 116.785 ;
        RECT 16.175 116.555 16.510 116.955 ;
        RECT 16.685 116.410 22.030 116.955 ;
        RECT 15.185 115.715 15.545 116.295 ;
        RECT 15.800 116.215 16.485 116.385 ;
        RECT 15.725 115.545 15.975 116.045 ;
        RECT 14.845 115.375 15.975 115.545 ;
        RECT 14.845 114.605 15.115 115.375 ;
        RECT 16.145 115.185 16.485 116.215 ;
        RECT 18.270 115.580 18.610 116.410 ;
        RECT 22.205 116.185 23.875 116.955 ;
        RECT 24.070 116.565 24.400 116.955 ;
        RECT 24.570 116.395 24.795 116.775 ;
        RECT 15.285 114.405 15.615 115.185 ;
        RECT 15.820 115.010 16.485 115.185 ;
        RECT 15.820 114.605 16.005 115.010 ;
        RECT 20.090 114.840 20.440 116.090 ;
        RECT 22.205 115.665 22.955 116.185 ;
        RECT 23.125 115.495 23.875 116.015 ;
        RECT 24.055 115.715 24.295 116.365 ;
        RECT 24.465 116.215 24.795 116.395 ;
        RECT 24.465 115.545 24.640 116.215 ;
        RECT 24.995 116.045 25.225 116.665 ;
        RECT 25.405 116.225 25.705 116.955 ;
        RECT 25.885 116.305 26.145 116.785 ;
        RECT 26.315 116.415 26.565 116.955 ;
        RECT 24.810 115.715 25.225 116.045 ;
        RECT 25.405 115.715 25.700 116.045 ;
        RECT 16.175 114.405 16.510 114.830 ;
        RECT 16.685 114.405 22.030 114.840 ;
        RECT 22.205 114.405 23.875 115.495 ;
        RECT 24.055 115.355 24.640 115.545 ;
        RECT 24.055 114.585 24.330 115.355 ;
        RECT 24.810 115.185 25.705 115.515 ;
        RECT 24.500 115.015 25.705 115.185 ;
        RECT 24.500 114.585 24.830 115.015 ;
        RECT 25.000 114.405 25.195 114.845 ;
        RECT 25.375 114.585 25.705 115.015 ;
        RECT 25.885 115.275 26.055 116.305 ;
        RECT 26.735 116.250 26.955 116.735 ;
        RECT 26.225 115.655 26.455 116.050 ;
        RECT 26.625 115.825 26.955 116.250 ;
        RECT 27.125 116.575 28.015 116.745 ;
        RECT 27.125 115.850 27.295 116.575 ;
        RECT 27.465 116.020 28.015 116.405 ;
        RECT 28.185 116.215 28.570 116.785 ;
        RECT 28.740 116.495 29.065 116.955 ;
        RECT 29.585 116.325 29.865 116.785 ;
        RECT 27.125 115.780 28.015 115.850 ;
        RECT 27.120 115.755 28.015 115.780 ;
        RECT 27.110 115.740 28.015 115.755 ;
        RECT 27.105 115.725 28.015 115.740 ;
        RECT 27.095 115.720 28.015 115.725 ;
        RECT 27.090 115.710 28.015 115.720 ;
        RECT 27.085 115.700 28.015 115.710 ;
        RECT 27.075 115.695 28.015 115.700 ;
        RECT 27.065 115.685 28.015 115.695 ;
        RECT 27.055 115.680 28.015 115.685 ;
        RECT 27.055 115.675 27.390 115.680 ;
        RECT 27.040 115.670 27.390 115.675 ;
        RECT 27.025 115.660 27.390 115.670 ;
        RECT 27.000 115.655 27.390 115.660 ;
        RECT 26.225 115.650 27.390 115.655 ;
        RECT 26.225 115.615 27.360 115.650 ;
        RECT 26.225 115.590 27.325 115.615 ;
        RECT 26.225 115.560 27.295 115.590 ;
        RECT 26.225 115.530 27.275 115.560 ;
        RECT 26.225 115.500 27.255 115.530 ;
        RECT 26.225 115.490 27.185 115.500 ;
        RECT 26.225 115.480 27.160 115.490 ;
        RECT 26.225 115.465 27.140 115.480 ;
        RECT 26.225 115.450 27.120 115.465 ;
        RECT 26.330 115.440 27.115 115.450 ;
        RECT 26.330 115.405 27.100 115.440 ;
        RECT 25.885 114.575 26.160 115.275 ;
        RECT 26.330 115.155 27.085 115.405 ;
        RECT 27.255 115.085 27.585 115.330 ;
        RECT 27.755 115.230 28.015 115.680 ;
        RECT 28.185 115.545 28.465 116.215 ;
        RECT 28.740 116.155 29.865 116.325 ;
        RECT 28.740 116.045 29.190 116.155 ;
        RECT 28.635 115.715 29.190 116.045 ;
        RECT 30.055 115.985 30.455 116.785 ;
        RECT 30.855 116.495 31.125 116.955 ;
        RECT 31.295 116.325 31.580 116.785 ;
        RECT 27.400 115.060 27.585 115.085 ;
        RECT 27.400 114.960 28.015 115.060 ;
        RECT 26.330 114.405 26.585 114.950 ;
        RECT 26.755 114.575 27.235 114.915 ;
        RECT 27.410 114.405 28.015 114.960 ;
        RECT 28.185 114.575 28.570 115.545 ;
        RECT 28.740 115.255 29.190 115.715 ;
        RECT 29.360 115.425 30.455 115.985 ;
        RECT 28.740 115.035 29.865 115.255 ;
        RECT 28.740 114.405 29.065 114.865 ;
        RECT 29.585 114.575 29.865 115.035 ;
        RECT 30.055 114.575 30.455 115.425 ;
        RECT 30.625 116.155 31.580 116.325 ;
        RECT 30.625 115.255 30.835 116.155 ;
        RECT 31.885 116.145 32.125 116.955 ;
        RECT 32.295 116.145 32.625 116.785 ;
        RECT 32.795 116.145 33.065 116.955 ;
        RECT 33.245 116.185 35.835 116.955 ;
        RECT 36.015 116.230 36.345 116.740 ;
        RECT 36.515 116.555 36.845 116.955 ;
        RECT 37.895 116.385 38.225 116.725 ;
        RECT 38.395 116.555 38.725 116.955 ;
        RECT 31.005 115.425 31.695 115.985 ;
        RECT 31.865 115.715 32.215 115.965 ;
        RECT 32.385 115.545 32.555 116.145 ;
        RECT 32.725 115.715 33.075 115.965 ;
        RECT 33.245 115.665 34.455 116.185 ;
        RECT 31.875 115.375 32.555 115.545 ;
        RECT 30.625 115.035 31.580 115.255 ;
        RECT 30.855 114.405 31.125 114.865 ;
        RECT 31.295 114.575 31.580 115.035 ;
        RECT 31.875 114.590 32.205 115.375 ;
        RECT 32.735 114.405 33.065 115.545 ;
        RECT 34.625 115.495 35.835 116.015 ;
        RECT 33.245 114.405 35.835 115.495 ;
        RECT 36.015 115.465 36.205 116.230 ;
        RECT 36.515 116.215 38.880 116.385 ;
        RECT 39.225 116.230 39.515 116.955 ;
        RECT 36.515 116.045 36.685 116.215 ;
        RECT 36.375 115.715 36.685 116.045 ;
        RECT 36.855 115.715 37.160 116.045 ;
        RECT 36.015 114.615 36.345 115.465 ;
        RECT 36.515 114.405 36.765 115.545 ;
        RECT 36.945 115.385 37.160 115.715 ;
        RECT 37.335 115.385 37.620 116.045 ;
        RECT 37.815 115.385 38.080 116.045 ;
        RECT 38.295 115.385 38.540 116.045 ;
        RECT 38.710 115.215 38.880 116.215 ;
        RECT 40.145 116.155 40.840 116.785 ;
        RECT 41.045 116.155 41.355 116.955 ;
        RECT 41.640 116.325 41.925 116.785 ;
        RECT 42.095 116.495 42.365 116.955 ;
        RECT 41.640 116.155 42.595 116.325 ;
        RECT 40.165 115.715 40.500 115.965 ;
        RECT 36.955 115.045 38.245 115.215 ;
        RECT 36.955 114.625 37.205 115.045 ;
        RECT 37.435 114.405 37.765 114.875 ;
        RECT 37.995 114.625 38.245 115.045 ;
        RECT 38.425 115.045 38.880 115.215 ;
        RECT 38.425 114.615 38.755 115.045 ;
        RECT 39.225 114.405 39.515 115.570 ;
        RECT 40.670 115.555 40.840 116.155 ;
        RECT 41.010 115.715 41.345 115.985 ;
        RECT 40.145 114.405 40.405 115.545 ;
        RECT 40.575 114.575 40.905 115.555 ;
        RECT 41.075 114.405 41.355 115.545 ;
        RECT 41.525 115.425 42.215 115.985 ;
        RECT 42.385 115.255 42.595 116.155 ;
        RECT 41.640 115.035 42.595 115.255 ;
        RECT 42.765 115.985 43.165 116.785 ;
        RECT 43.355 116.325 43.635 116.785 ;
        RECT 44.155 116.495 44.480 116.955 ;
        RECT 43.355 116.155 44.480 116.325 ;
        RECT 44.650 116.215 45.035 116.785 ;
        RECT 44.030 116.045 44.480 116.155 ;
        RECT 42.765 115.425 43.860 115.985 ;
        RECT 44.030 115.715 44.585 116.045 ;
        RECT 41.640 114.575 41.925 115.035 ;
        RECT 42.095 114.405 42.365 114.865 ;
        RECT 42.765 114.575 43.165 115.425 ;
        RECT 44.030 115.255 44.480 115.715 ;
        RECT 44.755 115.545 45.035 116.215 ;
        RECT 45.205 116.155 45.515 116.955 ;
        RECT 45.720 116.155 46.415 116.785 ;
        RECT 46.585 116.215 46.970 116.785 ;
        RECT 47.140 116.495 47.465 116.955 ;
        RECT 47.985 116.325 48.265 116.785 ;
        RECT 45.215 115.715 45.550 115.985 ;
        RECT 45.720 115.555 45.890 116.155 ;
        RECT 46.060 115.715 46.395 115.965 ;
        RECT 43.355 115.035 44.480 115.255 ;
        RECT 43.355 114.575 43.635 115.035 ;
        RECT 44.155 114.405 44.480 114.865 ;
        RECT 44.650 114.575 45.035 115.545 ;
        RECT 45.205 114.405 45.485 115.545 ;
        RECT 45.655 114.575 45.985 115.555 ;
        RECT 46.585 115.545 46.865 116.215 ;
        RECT 47.140 116.155 48.265 116.325 ;
        RECT 47.140 116.045 47.590 116.155 ;
        RECT 47.035 115.715 47.590 116.045 ;
        RECT 48.455 115.985 48.855 116.785 ;
        RECT 49.255 116.495 49.525 116.955 ;
        RECT 49.695 116.325 49.980 116.785 ;
        RECT 46.155 114.405 46.415 115.545 ;
        RECT 46.585 114.575 46.970 115.545 ;
        RECT 47.140 115.255 47.590 115.715 ;
        RECT 47.760 115.425 48.855 115.985 ;
        RECT 47.140 115.035 48.265 115.255 ;
        RECT 47.140 114.405 47.465 114.865 ;
        RECT 47.985 114.575 48.265 115.035 ;
        RECT 48.455 114.575 48.855 115.425 ;
        RECT 49.025 116.155 49.980 116.325 ;
        RECT 50.355 116.405 50.525 116.695 ;
        RECT 50.695 116.575 51.025 116.955 ;
        RECT 50.355 116.235 51.020 116.405 ;
        RECT 49.025 115.255 49.235 116.155 ;
        RECT 49.405 115.425 50.095 115.985 ;
        RECT 50.270 115.415 50.620 116.065 ;
        RECT 49.025 115.035 49.980 115.255 ;
        RECT 50.790 115.245 51.020 116.235 ;
        RECT 49.255 114.405 49.525 114.865 ;
        RECT 49.695 114.575 49.980 115.035 ;
        RECT 50.355 115.075 51.020 115.245 ;
        RECT 50.355 114.575 50.525 115.075 ;
        RECT 50.695 114.405 51.025 114.905 ;
        RECT 51.195 114.575 51.380 116.695 ;
        RECT 51.635 116.495 51.885 116.955 ;
        RECT 52.055 116.505 52.390 116.675 ;
        RECT 52.585 116.505 53.260 116.675 ;
        RECT 52.055 116.365 52.225 116.505 ;
        RECT 51.550 115.375 51.830 116.325 ;
        RECT 52.000 116.235 52.225 116.365 ;
        RECT 52.000 115.130 52.170 116.235 ;
        RECT 52.395 116.085 52.920 116.305 ;
        RECT 52.340 115.320 52.580 115.915 ;
        RECT 52.750 115.385 52.920 116.085 ;
        RECT 53.090 115.725 53.260 116.505 ;
        RECT 53.580 116.455 53.950 116.955 ;
        RECT 54.130 116.505 54.535 116.675 ;
        RECT 54.705 116.505 55.490 116.675 ;
        RECT 54.130 116.275 54.300 116.505 ;
        RECT 53.470 115.975 54.300 116.275 ;
        RECT 54.685 116.005 55.150 116.335 ;
        RECT 53.470 115.945 53.670 115.975 ;
        RECT 53.790 115.725 53.960 115.795 ;
        RECT 53.090 115.555 53.960 115.725 ;
        RECT 53.450 115.465 53.960 115.555 ;
        RECT 52.000 115.000 52.305 115.130 ;
        RECT 52.750 115.020 53.280 115.385 ;
        RECT 51.620 114.405 51.885 114.865 ;
        RECT 52.055 114.575 52.305 115.000 ;
        RECT 53.450 114.850 53.620 115.465 ;
        RECT 52.515 114.680 53.620 114.850 ;
        RECT 53.790 114.405 53.960 115.205 ;
        RECT 54.130 114.905 54.300 115.975 ;
        RECT 54.470 115.075 54.660 115.795 ;
        RECT 54.830 115.045 55.150 116.005 ;
        RECT 55.320 116.045 55.490 116.505 ;
        RECT 55.765 116.425 55.975 116.955 ;
        RECT 56.235 116.215 56.565 116.740 ;
        RECT 56.735 116.345 56.905 116.955 ;
        RECT 57.075 116.300 57.405 116.735 ;
        RECT 57.625 116.410 62.970 116.955 ;
        RECT 57.075 116.215 57.455 116.300 ;
        RECT 56.365 116.045 56.565 116.215 ;
        RECT 57.230 116.175 57.455 116.215 ;
        RECT 55.320 115.715 56.195 116.045 ;
        RECT 56.365 115.715 57.115 116.045 ;
        RECT 54.130 114.575 54.380 114.905 ;
        RECT 55.320 114.875 55.490 115.715 ;
        RECT 56.365 115.510 56.555 115.715 ;
        RECT 57.285 115.595 57.455 116.175 ;
        RECT 57.240 115.545 57.455 115.595 ;
        RECT 59.210 115.580 59.550 116.410 ;
        RECT 63.145 116.185 64.815 116.955 ;
        RECT 64.985 116.230 65.275 116.955 ;
        RECT 55.660 115.135 56.555 115.510 ;
        RECT 57.065 115.465 57.455 115.545 ;
        RECT 54.605 114.705 55.490 114.875 ;
        RECT 55.670 114.405 55.985 114.905 ;
        RECT 56.215 114.575 56.555 115.135 ;
        RECT 56.725 114.405 56.895 115.415 ;
        RECT 57.065 114.620 57.395 115.465 ;
        RECT 61.030 114.840 61.380 116.090 ;
        RECT 63.145 115.665 63.895 116.185 ;
        RECT 65.905 116.155 66.600 116.785 ;
        RECT 66.805 116.155 67.115 116.955 ;
        RECT 67.285 116.205 68.495 116.955 ;
        RECT 64.065 115.495 64.815 116.015 ;
        RECT 65.925 115.715 66.260 115.965 ;
        RECT 57.625 114.405 62.970 114.840 ;
        RECT 63.145 114.405 64.815 115.495 ;
        RECT 64.985 114.405 65.275 115.570 ;
        RECT 66.430 115.555 66.600 116.155 ;
        RECT 66.770 115.715 67.105 115.985 ;
        RECT 67.285 115.665 67.805 116.205 ;
        RECT 68.685 116.145 68.925 116.955 ;
        RECT 69.095 116.145 69.425 116.785 ;
        RECT 69.595 116.145 69.865 116.955 ;
        RECT 70.045 116.185 71.715 116.955 ;
        RECT 72.350 116.450 72.685 116.955 ;
        RECT 72.855 116.385 73.095 116.760 ;
        RECT 73.375 116.625 73.545 116.770 ;
        RECT 73.375 116.430 73.750 116.625 ;
        RECT 74.110 116.460 74.505 116.955 ;
        RECT 65.905 114.405 66.165 115.545 ;
        RECT 66.335 114.575 66.665 115.555 ;
        RECT 66.835 114.405 67.115 115.545 ;
        RECT 67.975 115.495 68.495 116.035 ;
        RECT 68.665 115.715 69.015 115.965 ;
        RECT 69.185 115.545 69.355 116.145 ;
        RECT 69.525 115.715 69.875 115.965 ;
        RECT 70.045 115.665 70.795 116.185 ;
        RECT 67.285 114.405 68.495 115.495 ;
        RECT 68.675 115.375 69.355 115.545 ;
        RECT 68.675 114.590 69.005 115.375 ;
        RECT 69.535 114.405 69.865 115.545 ;
        RECT 70.965 115.495 71.715 116.015 ;
        RECT 70.045 114.405 71.715 115.495 ;
        RECT 72.405 115.425 72.705 116.275 ;
        RECT 72.875 116.235 73.095 116.385 ;
        RECT 72.875 115.905 73.410 116.235 ;
        RECT 73.580 116.095 73.750 116.430 ;
        RECT 74.675 116.265 74.915 116.785 ;
        RECT 75.105 116.410 80.450 116.955 ;
        RECT 80.625 116.410 85.970 116.955 ;
        RECT 72.875 115.255 73.110 115.905 ;
        RECT 73.580 115.735 74.565 116.095 ;
        RECT 72.435 115.025 73.110 115.255 ;
        RECT 73.280 115.715 74.565 115.735 ;
        RECT 73.280 115.565 74.140 115.715 ;
        RECT 72.435 114.595 72.605 115.025 ;
        RECT 72.775 114.405 73.105 114.855 ;
        RECT 73.280 114.620 73.565 115.565 ;
        RECT 74.740 115.460 74.915 116.265 ;
        RECT 76.690 115.580 77.030 116.410 ;
        RECT 73.740 115.085 74.435 115.395 ;
        RECT 73.745 114.405 74.430 114.875 ;
        RECT 74.610 114.675 74.915 115.460 ;
        RECT 78.510 114.840 78.860 116.090 ;
        RECT 82.210 115.580 82.550 116.410 ;
        RECT 86.145 116.185 88.735 116.955 ;
        RECT 88.995 116.405 89.165 116.785 ;
        RECT 89.380 116.575 89.710 116.955 ;
        RECT 88.995 116.235 89.710 116.405 ;
        RECT 84.030 114.840 84.380 116.090 ;
        RECT 86.145 115.665 87.355 116.185 ;
        RECT 87.525 115.495 88.735 116.015 ;
        RECT 88.905 115.685 89.260 116.055 ;
        RECT 89.540 116.045 89.710 116.235 ;
        RECT 89.880 116.210 90.135 116.785 ;
        RECT 89.540 115.715 89.795 116.045 ;
        RECT 89.540 115.505 89.710 115.715 ;
        RECT 75.105 114.405 80.450 114.840 ;
        RECT 80.625 114.405 85.970 114.840 ;
        RECT 86.145 114.405 88.735 115.495 ;
        RECT 88.995 115.335 89.710 115.505 ;
        RECT 89.965 115.480 90.135 116.210 ;
        RECT 90.310 116.115 90.570 116.955 ;
        RECT 90.745 116.205 91.955 116.955 ;
        RECT 100.580 116.800 106.320 116.810 ;
        RECT 88.995 114.575 89.165 115.335 ;
        RECT 89.380 114.405 89.710 115.165 ;
        RECT 89.880 114.575 90.135 115.480 ;
        RECT 90.310 114.405 90.570 115.555 ;
        RECT 90.745 115.495 91.265 116.035 ;
        RECT 91.435 115.665 91.955 116.205 ;
        RECT 100.090 116.640 106.320 116.800 ;
        RECT 90.745 114.405 91.955 115.495 ;
        RECT 13.380 114.235 92.040 114.405 ;
        RECT 100.090 114.380 100.760 116.640 ;
        RECT 101.430 116.070 105.470 116.240 ;
        RECT 101.090 115.010 101.260 116.010 ;
        RECT 105.640 115.010 105.810 116.010 ;
        RECT 101.430 114.780 105.470 114.950 ;
        RECT 106.150 114.380 106.320 116.640 ;
        RECT 13.465 113.145 14.675 114.235 ;
        RECT 14.845 113.640 15.280 114.065 ;
        RECT 15.450 113.810 15.835 114.235 ;
        RECT 14.845 113.470 15.835 113.640 ;
        RECT 13.465 112.435 13.985 112.975 ;
        RECT 14.155 112.605 14.675 113.145 ;
        RECT 14.845 112.595 15.330 113.300 ;
        RECT 15.500 112.925 15.835 113.470 ;
        RECT 16.005 113.275 16.430 114.065 ;
        RECT 16.600 113.640 16.875 114.065 ;
        RECT 17.045 113.810 17.430 114.235 ;
        RECT 16.600 113.445 17.430 113.640 ;
        RECT 16.005 113.095 16.910 113.275 ;
        RECT 15.500 112.595 15.910 112.925 ;
        RECT 16.080 112.595 16.910 113.095 ;
        RECT 17.080 112.925 17.430 113.445 ;
        RECT 17.600 113.275 17.845 114.065 ;
        RECT 18.035 113.640 18.290 114.065 ;
        RECT 18.460 113.810 18.845 114.235 ;
        RECT 18.035 113.445 18.845 113.640 ;
        RECT 17.600 113.095 18.325 113.275 ;
        RECT 17.080 112.595 17.505 112.925 ;
        RECT 17.675 112.595 18.325 113.095 ;
        RECT 18.495 112.925 18.845 113.445 ;
        RECT 19.015 113.095 19.275 114.065 ;
        RECT 18.495 112.595 18.920 112.925 ;
        RECT 13.465 111.685 14.675 112.435 ;
        RECT 15.500 112.425 15.835 112.595 ;
        RECT 16.080 112.425 16.430 112.595 ;
        RECT 17.080 112.425 17.430 112.595 ;
        RECT 17.675 112.425 17.845 112.595 ;
        RECT 18.495 112.425 18.845 112.595 ;
        RECT 19.090 112.425 19.275 113.095 ;
        RECT 14.845 112.255 15.835 112.425 ;
        RECT 14.845 111.855 15.280 112.255 ;
        RECT 15.450 111.685 15.835 112.085 ;
        RECT 16.005 111.855 16.430 112.425 ;
        RECT 16.620 112.255 17.430 112.425 ;
        RECT 16.620 111.855 16.875 112.255 ;
        RECT 17.045 111.685 17.430 112.085 ;
        RECT 17.600 111.855 17.845 112.425 ;
        RECT 18.035 112.255 18.845 112.425 ;
        RECT 18.035 111.855 18.290 112.255 ;
        RECT 18.460 111.685 18.845 112.085 ;
        RECT 19.015 111.855 19.275 112.425 ;
        RECT 19.445 113.095 19.830 114.065 ;
        RECT 20.000 113.775 20.325 114.235 ;
        RECT 20.845 113.605 21.125 114.065 ;
        RECT 20.000 113.385 21.125 113.605 ;
        RECT 19.445 112.425 19.725 113.095 ;
        RECT 20.000 112.925 20.450 113.385 ;
        RECT 21.315 113.215 21.715 114.065 ;
        RECT 22.115 113.775 22.385 114.235 ;
        RECT 22.555 113.605 22.840 114.065 ;
        RECT 19.895 112.595 20.450 112.925 ;
        RECT 20.620 112.655 21.715 113.215 ;
        RECT 20.000 112.485 20.450 112.595 ;
        RECT 19.445 111.855 19.830 112.425 ;
        RECT 20.000 112.315 21.125 112.485 ;
        RECT 20.000 111.685 20.325 112.145 ;
        RECT 20.845 111.855 21.125 112.315 ;
        RECT 21.315 111.855 21.715 112.655 ;
        RECT 21.885 113.385 22.840 113.605 ;
        RECT 21.885 112.485 22.095 113.385 ;
        RECT 22.265 112.655 22.955 113.215 ;
        RECT 23.125 113.145 25.715 114.235 ;
        RECT 21.885 112.315 22.840 112.485 ;
        RECT 22.115 111.685 22.385 112.145 ;
        RECT 22.555 111.855 22.840 112.315 ;
        RECT 23.125 112.455 24.335 112.975 ;
        RECT 24.505 112.625 25.715 113.145 ;
        RECT 26.345 113.070 26.635 114.235 ;
        RECT 26.805 113.800 32.150 114.235 ;
        RECT 23.125 111.685 25.715 112.455 ;
        RECT 26.345 111.685 26.635 112.410 ;
        RECT 28.390 112.230 28.730 113.060 ;
        RECT 30.210 112.550 30.560 113.800 ;
        RECT 32.325 113.145 33.995 114.235 ;
        RECT 34.715 113.565 34.885 114.065 ;
        RECT 35.055 113.735 35.385 114.235 ;
        RECT 34.715 113.395 35.380 113.565 ;
        RECT 32.325 112.455 33.075 112.975 ;
        RECT 33.245 112.625 33.995 113.145 ;
        RECT 34.630 112.575 34.980 113.225 ;
        RECT 26.805 111.685 32.150 112.230 ;
        RECT 32.325 111.685 33.995 112.455 ;
        RECT 35.150 112.405 35.380 113.395 ;
        RECT 34.715 112.235 35.380 112.405 ;
        RECT 34.715 111.945 34.885 112.235 ;
        RECT 35.055 111.685 35.385 112.065 ;
        RECT 35.555 111.945 35.740 114.065 ;
        RECT 35.980 113.775 36.245 114.235 ;
        RECT 36.415 113.640 36.665 114.065 ;
        RECT 36.875 113.790 37.980 113.960 ;
        RECT 36.360 113.510 36.665 113.640 ;
        RECT 35.910 112.315 36.190 113.265 ;
        RECT 36.360 112.405 36.530 113.510 ;
        RECT 36.700 112.725 36.940 113.320 ;
        RECT 37.110 113.255 37.640 113.620 ;
        RECT 37.110 112.555 37.280 113.255 ;
        RECT 37.810 113.175 37.980 113.790 ;
        RECT 38.150 113.435 38.320 114.235 ;
        RECT 38.490 113.735 38.740 114.065 ;
        RECT 38.965 113.765 39.850 113.935 ;
        RECT 37.810 113.085 38.320 113.175 ;
        RECT 36.360 112.275 36.585 112.405 ;
        RECT 36.755 112.335 37.280 112.555 ;
        RECT 37.450 112.915 38.320 113.085 ;
        RECT 35.995 111.685 36.245 112.145 ;
        RECT 36.415 112.135 36.585 112.275 ;
        RECT 37.450 112.135 37.620 112.915 ;
        RECT 38.150 112.845 38.320 112.915 ;
        RECT 37.830 112.665 38.030 112.695 ;
        RECT 38.490 112.665 38.660 113.735 ;
        RECT 38.830 112.845 39.020 113.565 ;
        RECT 37.830 112.365 38.660 112.665 ;
        RECT 39.190 112.635 39.510 113.595 ;
        RECT 36.415 111.965 36.750 112.135 ;
        RECT 36.945 111.965 37.620 112.135 ;
        RECT 37.940 111.685 38.310 112.185 ;
        RECT 38.490 112.135 38.660 112.365 ;
        RECT 39.045 112.305 39.510 112.635 ;
        RECT 39.680 112.925 39.850 113.765 ;
        RECT 40.030 113.735 40.345 114.235 ;
        RECT 40.575 113.505 40.915 114.065 ;
        RECT 40.020 113.130 40.915 113.505 ;
        RECT 41.085 113.225 41.255 114.235 ;
        RECT 40.725 112.925 40.915 113.130 ;
        RECT 41.425 113.175 41.755 114.020 ;
        RECT 41.425 113.095 41.815 113.175 ;
        RECT 41.600 113.045 41.815 113.095 ;
        RECT 39.680 112.595 40.555 112.925 ;
        RECT 40.725 112.595 41.475 112.925 ;
        RECT 39.680 112.135 39.850 112.595 ;
        RECT 40.725 112.425 40.925 112.595 ;
        RECT 41.645 112.465 41.815 113.045 ;
        RECT 41.590 112.425 41.815 112.465 ;
        RECT 38.490 111.965 38.895 112.135 ;
        RECT 39.065 111.965 39.850 112.135 ;
        RECT 40.125 111.685 40.335 112.215 ;
        RECT 40.595 111.900 40.925 112.425 ;
        RECT 41.435 112.340 41.815 112.425 ;
        RECT 41.095 111.685 41.265 112.295 ;
        RECT 41.435 111.905 41.765 112.340 ;
        RECT 41.995 111.865 42.255 114.055 ;
        RECT 42.425 113.505 42.765 114.235 ;
        RECT 42.945 113.325 43.215 114.055 ;
        RECT 42.445 113.105 43.215 113.325 ;
        RECT 43.395 113.345 43.625 114.055 ;
        RECT 43.795 113.525 44.125 114.235 ;
        RECT 44.295 113.345 44.555 114.055 ;
        RECT 44.835 113.565 45.005 114.065 ;
        RECT 45.175 113.735 45.505 114.235 ;
        RECT 44.835 113.395 45.500 113.565 ;
        RECT 43.395 113.105 44.555 113.345 ;
        RECT 42.445 112.435 42.735 113.105 ;
        RECT 42.915 112.615 43.380 112.925 ;
        RECT 43.560 112.615 44.085 112.925 ;
        RECT 42.445 112.235 43.675 112.435 ;
        RECT 42.515 111.685 43.185 112.055 ;
        RECT 43.365 111.865 43.675 112.235 ;
        RECT 43.855 111.975 44.085 112.615 ;
        RECT 44.265 112.595 44.565 112.925 ;
        RECT 44.750 112.575 45.100 113.225 ;
        RECT 44.265 111.685 44.555 112.415 ;
        RECT 45.270 112.405 45.500 113.395 ;
        RECT 44.835 112.235 45.500 112.405 ;
        RECT 44.835 111.945 45.005 112.235 ;
        RECT 45.175 111.685 45.505 112.065 ;
        RECT 45.675 111.945 45.860 114.065 ;
        RECT 46.100 113.775 46.365 114.235 ;
        RECT 46.535 113.640 46.785 114.065 ;
        RECT 46.995 113.790 48.100 113.960 ;
        RECT 46.480 113.510 46.785 113.640 ;
        RECT 46.030 112.315 46.310 113.265 ;
        RECT 46.480 112.405 46.650 113.510 ;
        RECT 46.820 112.725 47.060 113.320 ;
        RECT 47.230 113.255 47.760 113.620 ;
        RECT 47.230 112.555 47.400 113.255 ;
        RECT 47.930 113.175 48.100 113.790 ;
        RECT 48.270 113.435 48.440 114.235 ;
        RECT 48.610 113.735 48.860 114.065 ;
        RECT 49.085 113.765 49.970 113.935 ;
        RECT 47.930 113.085 48.440 113.175 ;
        RECT 46.480 112.275 46.705 112.405 ;
        RECT 46.875 112.335 47.400 112.555 ;
        RECT 47.570 112.915 48.440 113.085 ;
        RECT 46.115 111.685 46.365 112.145 ;
        RECT 46.535 112.135 46.705 112.275 ;
        RECT 47.570 112.135 47.740 112.915 ;
        RECT 48.270 112.845 48.440 112.915 ;
        RECT 47.950 112.665 48.150 112.695 ;
        RECT 48.610 112.665 48.780 113.735 ;
        RECT 48.950 112.845 49.140 113.565 ;
        RECT 47.950 112.365 48.780 112.665 ;
        RECT 49.310 112.635 49.630 113.595 ;
        RECT 46.535 111.965 46.870 112.135 ;
        RECT 47.065 111.965 47.740 112.135 ;
        RECT 48.060 111.685 48.430 112.185 ;
        RECT 48.610 112.135 48.780 112.365 ;
        RECT 49.165 112.305 49.630 112.635 ;
        RECT 49.800 112.925 49.970 113.765 ;
        RECT 50.150 113.735 50.465 114.235 ;
        RECT 50.695 113.505 51.035 114.065 ;
        RECT 50.140 113.130 51.035 113.505 ;
        RECT 51.205 113.225 51.375 114.235 ;
        RECT 50.845 112.925 51.035 113.130 ;
        RECT 51.545 113.175 51.875 114.020 ;
        RECT 51.545 113.095 51.935 113.175 ;
        RECT 51.720 113.045 51.935 113.095 ;
        RECT 52.105 113.070 52.395 114.235 ;
        RECT 52.565 113.145 55.155 114.235 ;
        RECT 55.325 113.725 55.585 114.235 ;
        RECT 49.800 112.595 50.675 112.925 ;
        RECT 50.845 112.595 51.595 112.925 ;
        RECT 49.800 112.135 49.970 112.595 ;
        RECT 50.845 112.425 51.045 112.595 ;
        RECT 51.765 112.465 51.935 113.045 ;
        RECT 51.710 112.425 51.935 112.465 ;
        RECT 48.610 111.965 49.015 112.135 ;
        RECT 49.185 111.965 49.970 112.135 ;
        RECT 50.245 111.685 50.455 112.215 ;
        RECT 50.715 111.900 51.045 112.425 ;
        RECT 51.555 112.340 51.935 112.425 ;
        RECT 52.565 112.455 53.775 112.975 ;
        RECT 53.945 112.625 55.155 113.145 ;
        RECT 55.325 112.675 55.665 113.555 ;
        RECT 55.835 112.845 56.005 114.065 ;
        RECT 56.245 113.730 56.860 114.235 ;
        RECT 56.245 113.195 56.495 113.560 ;
        RECT 56.665 113.555 56.860 113.730 ;
        RECT 57.030 113.725 57.505 114.065 ;
        RECT 57.675 113.690 57.890 114.235 ;
        RECT 56.665 113.365 56.995 113.555 ;
        RECT 57.215 113.195 57.930 113.490 ;
        RECT 58.100 113.365 58.375 114.065 ;
        RECT 58.635 113.565 58.805 114.065 ;
        RECT 58.975 113.735 59.305 114.235 ;
        RECT 58.635 113.395 59.300 113.565 ;
        RECT 56.245 113.025 58.035 113.195 ;
        RECT 55.835 112.595 56.630 112.845 ;
        RECT 55.835 112.505 56.085 112.595 ;
        RECT 51.215 111.685 51.385 112.295 ;
        RECT 51.555 111.905 51.885 112.340 ;
        RECT 52.105 111.685 52.395 112.410 ;
        RECT 52.565 111.685 55.155 112.455 ;
        RECT 55.325 111.685 55.585 112.505 ;
        RECT 55.755 112.085 56.085 112.505 ;
        RECT 56.800 112.170 57.055 113.025 ;
        RECT 56.265 111.905 57.055 112.170 ;
        RECT 57.225 112.325 57.635 112.845 ;
        RECT 57.805 112.595 58.035 113.025 ;
        RECT 58.205 112.335 58.375 113.365 ;
        RECT 58.550 112.575 58.900 113.225 ;
        RECT 59.070 112.405 59.300 113.395 ;
        RECT 57.225 111.905 57.425 112.325 ;
        RECT 57.615 111.685 57.945 112.145 ;
        RECT 58.115 111.855 58.375 112.335 ;
        RECT 58.635 112.235 59.300 112.405 ;
        RECT 58.635 111.945 58.805 112.235 ;
        RECT 58.975 111.685 59.305 112.065 ;
        RECT 59.475 111.945 59.660 114.065 ;
        RECT 59.900 113.775 60.165 114.235 ;
        RECT 60.335 113.640 60.585 114.065 ;
        RECT 60.795 113.790 61.900 113.960 ;
        RECT 60.280 113.510 60.585 113.640 ;
        RECT 59.830 112.315 60.110 113.265 ;
        RECT 60.280 112.405 60.450 113.510 ;
        RECT 60.620 112.725 60.860 113.320 ;
        RECT 61.030 113.255 61.560 113.620 ;
        RECT 61.030 112.555 61.200 113.255 ;
        RECT 61.730 113.175 61.900 113.790 ;
        RECT 62.070 113.435 62.240 114.235 ;
        RECT 62.410 113.735 62.660 114.065 ;
        RECT 62.885 113.765 63.770 113.935 ;
        RECT 61.730 113.085 62.240 113.175 ;
        RECT 60.280 112.275 60.505 112.405 ;
        RECT 60.675 112.335 61.200 112.555 ;
        RECT 61.370 112.915 62.240 113.085 ;
        RECT 59.915 111.685 60.165 112.145 ;
        RECT 60.335 112.135 60.505 112.275 ;
        RECT 61.370 112.135 61.540 112.915 ;
        RECT 62.070 112.845 62.240 112.915 ;
        RECT 61.750 112.665 61.950 112.695 ;
        RECT 62.410 112.665 62.580 113.735 ;
        RECT 62.750 112.845 62.940 113.565 ;
        RECT 61.750 112.365 62.580 112.665 ;
        RECT 63.110 112.635 63.430 113.595 ;
        RECT 60.335 111.965 60.670 112.135 ;
        RECT 60.865 111.965 61.540 112.135 ;
        RECT 61.860 111.685 62.230 112.185 ;
        RECT 62.410 112.135 62.580 112.365 ;
        RECT 62.965 112.305 63.430 112.635 ;
        RECT 63.600 112.925 63.770 113.765 ;
        RECT 63.950 113.735 64.265 114.235 ;
        RECT 64.495 113.505 64.835 114.065 ;
        RECT 63.940 113.130 64.835 113.505 ;
        RECT 65.005 113.225 65.175 114.235 ;
        RECT 64.645 112.925 64.835 113.130 ;
        RECT 65.345 113.175 65.675 114.020 ;
        RECT 65.915 113.265 66.245 114.050 ;
        RECT 65.345 113.095 65.735 113.175 ;
        RECT 65.915 113.095 66.595 113.265 ;
        RECT 66.775 113.095 67.105 114.235 ;
        RECT 67.285 113.145 68.495 114.235 ;
        RECT 65.520 113.045 65.735 113.095 ;
        RECT 63.600 112.595 64.475 112.925 ;
        RECT 64.645 112.595 65.395 112.925 ;
        RECT 63.600 112.135 63.770 112.595 ;
        RECT 64.645 112.425 64.845 112.595 ;
        RECT 65.565 112.465 65.735 113.045 ;
        RECT 65.905 112.675 66.255 112.925 ;
        RECT 66.425 112.495 66.595 113.095 ;
        RECT 66.765 112.675 67.115 112.925 ;
        RECT 65.510 112.425 65.735 112.465 ;
        RECT 62.410 111.965 62.815 112.135 ;
        RECT 62.985 111.965 63.770 112.135 ;
        RECT 64.045 111.685 64.255 112.215 ;
        RECT 64.515 111.900 64.845 112.425 ;
        RECT 65.355 112.340 65.735 112.425 ;
        RECT 65.015 111.685 65.185 112.295 ;
        RECT 65.355 111.905 65.685 112.340 ;
        RECT 65.925 111.685 66.165 112.495 ;
        RECT 66.335 111.855 66.665 112.495 ;
        RECT 66.835 111.685 67.105 112.495 ;
        RECT 67.285 112.435 67.805 112.975 ;
        RECT 67.975 112.605 68.495 113.145 ;
        RECT 68.725 113.095 68.935 114.235 ;
        RECT 69.105 113.085 69.435 114.065 ;
        RECT 69.605 113.095 69.835 114.235 ;
        RECT 70.105 113.175 70.435 114.020 ;
        RECT 70.605 113.225 70.775 114.235 ;
        RECT 70.945 113.505 71.285 114.065 ;
        RECT 71.515 113.735 71.830 114.235 ;
        RECT 72.010 113.765 72.895 113.935 ;
        RECT 70.045 113.095 70.435 113.175 ;
        RECT 70.945 113.130 71.840 113.505 ;
        RECT 67.285 111.685 68.495 112.435 ;
        RECT 68.725 111.685 68.935 112.505 ;
        RECT 69.105 112.485 69.355 113.085 ;
        RECT 70.045 113.045 70.260 113.095 ;
        RECT 69.525 112.675 69.855 112.925 ;
        RECT 69.105 111.855 69.435 112.485 ;
        RECT 69.605 111.685 69.835 112.505 ;
        RECT 70.045 112.465 70.215 113.045 ;
        RECT 70.945 112.925 71.135 113.130 ;
        RECT 72.010 112.925 72.180 113.765 ;
        RECT 73.120 113.735 73.370 114.065 ;
        RECT 70.385 112.595 71.135 112.925 ;
        RECT 71.305 112.595 72.180 112.925 ;
        RECT 70.045 112.425 70.270 112.465 ;
        RECT 70.935 112.425 71.135 112.595 ;
        RECT 70.045 112.340 70.425 112.425 ;
        RECT 70.095 111.905 70.425 112.340 ;
        RECT 70.595 111.685 70.765 112.295 ;
        RECT 70.935 111.900 71.265 112.425 ;
        RECT 71.525 111.685 71.735 112.215 ;
        RECT 72.010 112.135 72.180 112.595 ;
        RECT 72.350 112.635 72.670 113.595 ;
        RECT 72.840 112.845 73.030 113.565 ;
        RECT 73.200 112.665 73.370 113.735 ;
        RECT 73.540 113.435 73.710 114.235 ;
        RECT 73.880 113.790 74.985 113.960 ;
        RECT 73.880 113.175 74.050 113.790 ;
        RECT 75.195 113.640 75.445 114.065 ;
        RECT 75.615 113.775 75.880 114.235 ;
        RECT 74.220 113.255 74.750 113.620 ;
        RECT 75.195 113.510 75.500 113.640 ;
        RECT 73.540 113.085 74.050 113.175 ;
        RECT 73.540 112.915 74.410 113.085 ;
        RECT 73.540 112.845 73.710 112.915 ;
        RECT 73.830 112.665 74.030 112.695 ;
        RECT 72.350 112.305 72.815 112.635 ;
        RECT 73.200 112.365 74.030 112.665 ;
        RECT 73.200 112.135 73.370 112.365 ;
        RECT 72.010 111.965 72.795 112.135 ;
        RECT 72.965 111.965 73.370 112.135 ;
        RECT 73.550 111.685 73.920 112.185 ;
        RECT 74.240 112.135 74.410 112.915 ;
        RECT 74.580 112.555 74.750 113.255 ;
        RECT 74.920 112.725 75.160 113.320 ;
        RECT 74.580 112.335 75.105 112.555 ;
        RECT 75.330 112.405 75.500 113.510 ;
        RECT 75.275 112.275 75.500 112.405 ;
        RECT 75.670 112.315 75.950 113.265 ;
        RECT 75.275 112.135 75.445 112.275 ;
        RECT 74.240 111.965 74.915 112.135 ;
        RECT 75.110 111.965 75.445 112.135 ;
        RECT 75.615 111.685 75.865 112.145 ;
        RECT 76.120 111.945 76.305 114.065 ;
        RECT 76.475 113.735 76.805 114.235 ;
        RECT 76.975 113.565 77.145 114.065 ;
        RECT 76.480 113.395 77.145 113.565 ;
        RECT 76.480 112.405 76.710 113.395 ;
        RECT 76.880 112.575 77.230 113.225 ;
        RECT 77.865 113.070 78.155 114.235 ;
        RECT 78.325 113.800 83.670 114.235 ;
        RECT 76.480 112.235 77.145 112.405 ;
        RECT 76.475 111.685 76.805 112.065 ;
        RECT 76.975 111.945 77.145 112.235 ;
        RECT 77.865 111.685 78.155 112.410 ;
        RECT 79.910 112.230 80.250 113.060 ;
        RECT 81.730 112.550 82.080 113.800 ;
        RECT 83.845 113.145 87.355 114.235 ;
        RECT 83.845 112.455 85.495 112.975 ;
        RECT 85.665 112.625 87.355 113.145 ;
        RECT 87.615 113.305 87.785 114.065 ;
        RECT 87.965 113.475 88.295 114.235 ;
        RECT 87.615 113.135 88.280 113.305 ;
        RECT 88.465 113.160 88.735 114.065 ;
        RECT 88.110 112.990 88.280 113.135 ;
        RECT 87.545 112.585 87.875 112.955 ;
        RECT 88.110 112.660 88.395 112.990 ;
        RECT 78.325 111.685 83.670 112.230 ;
        RECT 83.845 111.685 87.355 112.455 ;
        RECT 88.110 112.405 88.280 112.660 ;
        RECT 87.615 112.235 88.280 112.405 ;
        RECT 88.565 112.360 88.735 113.160 ;
        RECT 88.995 113.305 89.165 114.065 ;
        RECT 89.380 113.475 89.710 114.235 ;
        RECT 88.995 113.135 89.710 113.305 ;
        RECT 89.880 113.160 90.135 114.065 ;
        RECT 88.905 112.585 89.260 112.955 ;
        RECT 89.540 112.925 89.710 113.135 ;
        RECT 89.540 112.595 89.795 112.925 ;
        RECT 89.540 112.405 89.710 112.595 ;
        RECT 89.965 112.430 90.135 113.160 ;
        RECT 90.310 113.085 90.570 114.235 ;
        RECT 90.745 113.145 91.955 114.235 ;
        RECT 100.090 114.210 106.320 114.380 ;
        RECT 90.745 112.605 91.265 113.145 ;
        RECT 87.615 111.855 87.785 112.235 ;
        RECT 87.965 111.685 88.295 112.065 ;
        RECT 88.475 111.855 88.735 112.360 ;
        RECT 88.995 112.235 89.710 112.405 ;
        RECT 88.995 111.855 89.165 112.235 ;
        RECT 89.380 111.685 89.710 112.065 ;
        RECT 89.880 111.855 90.135 112.430 ;
        RECT 90.310 111.685 90.570 112.525 ;
        RECT 91.435 112.435 91.955 112.975 ;
        RECT 90.745 111.685 91.955 112.435 ;
        RECT 13.380 111.515 92.040 111.685 ;
        RECT 13.465 110.765 14.675 111.515 ;
        RECT 14.845 110.765 16.055 111.515 ;
        RECT 16.230 110.985 16.520 111.335 ;
        RECT 16.715 111.155 17.045 111.515 ;
        RECT 17.215 110.985 17.445 111.290 ;
        RECT 16.230 110.815 17.445 110.985 ;
        RECT 13.465 110.225 13.985 110.765 ;
        RECT 14.155 110.055 14.675 110.595 ;
        RECT 14.845 110.225 15.365 110.765 ;
        RECT 17.635 110.645 17.805 111.210 ;
        RECT 18.180 110.885 18.465 111.345 ;
        RECT 18.635 111.055 18.905 111.515 ;
        RECT 18.180 110.715 19.135 110.885 ;
        RECT 15.535 110.055 16.055 110.595 ;
        RECT 16.290 110.495 16.550 110.605 ;
        RECT 16.285 110.325 16.550 110.495 ;
        RECT 16.290 110.275 16.550 110.325 ;
        RECT 16.730 110.275 17.115 110.605 ;
        RECT 17.285 110.475 17.805 110.645 ;
        RECT 13.465 108.965 14.675 110.055 ;
        RECT 14.845 108.965 16.055 110.055 ;
        RECT 16.230 108.965 16.550 110.105 ;
        RECT 16.730 109.225 16.925 110.275 ;
        RECT 17.285 110.095 17.455 110.475 ;
        RECT 17.105 109.815 17.455 110.095 ;
        RECT 17.645 109.945 17.890 110.305 ;
        RECT 18.065 109.985 18.755 110.545 ;
        RECT 18.925 109.815 19.135 110.715 ;
        RECT 17.105 109.135 17.435 109.815 ;
        RECT 17.635 108.965 17.890 109.765 ;
        RECT 18.180 109.595 19.135 109.815 ;
        RECT 19.305 110.545 19.705 111.345 ;
        RECT 19.895 110.885 20.175 111.345 ;
        RECT 20.695 111.055 21.020 111.515 ;
        RECT 19.895 110.715 21.020 110.885 ;
        RECT 21.190 110.775 21.575 111.345 ;
        RECT 21.835 110.965 22.005 111.255 ;
        RECT 22.175 111.135 22.505 111.515 ;
        RECT 21.835 110.795 22.500 110.965 ;
        RECT 20.570 110.605 21.020 110.715 ;
        RECT 19.305 109.985 20.400 110.545 ;
        RECT 20.570 110.275 21.125 110.605 ;
        RECT 18.180 109.135 18.465 109.595 ;
        RECT 18.635 108.965 18.905 109.425 ;
        RECT 19.305 109.135 19.705 109.985 ;
        RECT 20.570 109.815 21.020 110.275 ;
        RECT 21.295 110.105 21.575 110.775 ;
        RECT 19.895 109.595 21.020 109.815 ;
        RECT 19.895 109.135 20.175 109.595 ;
        RECT 20.695 108.965 21.020 109.425 ;
        RECT 21.190 109.135 21.575 110.105 ;
        RECT 21.750 109.975 22.100 110.625 ;
        RECT 22.270 109.805 22.500 110.795 ;
        RECT 21.835 109.635 22.500 109.805 ;
        RECT 21.835 109.135 22.005 109.635 ;
        RECT 22.175 108.965 22.505 109.465 ;
        RECT 22.675 109.135 22.860 111.255 ;
        RECT 23.115 111.055 23.365 111.515 ;
        RECT 23.535 111.065 23.870 111.235 ;
        RECT 24.065 111.065 24.740 111.235 ;
        RECT 23.535 110.925 23.705 111.065 ;
        RECT 23.030 109.935 23.310 110.885 ;
        RECT 23.480 110.795 23.705 110.925 ;
        RECT 23.480 109.690 23.650 110.795 ;
        RECT 23.875 110.645 24.400 110.865 ;
        RECT 23.820 109.880 24.060 110.475 ;
        RECT 24.230 109.945 24.400 110.645 ;
        RECT 24.570 110.285 24.740 111.065 ;
        RECT 25.060 111.015 25.430 111.515 ;
        RECT 25.610 111.065 26.015 111.235 ;
        RECT 26.185 111.065 26.970 111.235 ;
        RECT 25.610 110.835 25.780 111.065 ;
        RECT 24.950 110.535 25.780 110.835 ;
        RECT 26.165 110.565 26.630 110.895 ;
        RECT 24.950 110.505 25.150 110.535 ;
        RECT 25.270 110.285 25.440 110.355 ;
        RECT 24.570 110.115 25.440 110.285 ;
        RECT 24.930 110.025 25.440 110.115 ;
        RECT 23.480 109.560 23.785 109.690 ;
        RECT 24.230 109.580 24.760 109.945 ;
        RECT 23.100 108.965 23.365 109.425 ;
        RECT 23.535 109.135 23.785 109.560 ;
        RECT 24.930 109.410 25.100 110.025 ;
        RECT 23.995 109.240 25.100 109.410 ;
        RECT 25.270 108.965 25.440 109.765 ;
        RECT 25.610 109.465 25.780 110.535 ;
        RECT 25.950 109.635 26.140 110.355 ;
        RECT 26.310 109.605 26.630 110.565 ;
        RECT 26.800 110.605 26.970 111.065 ;
        RECT 27.245 110.985 27.455 111.515 ;
        RECT 27.715 110.775 28.045 111.300 ;
        RECT 28.215 110.905 28.385 111.515 ;
        RECT 28.555 110.860 28.885 111.295 ;
        RECT 28.555 110.775 28.935 110.860 ;
        RECT 27.845 110.605 28.045 110.775 ;
        RECT 28.710 110.735 28.935 110.775 ;
        RECT 26.800 110.275 27.675 110.605 ;
        RECT 27.845 110.275 28.595 110.605 ;
        RECT 25.610 109.135 25.860 109.465 ;
        RECT 26.800 109.435 26.970 110.275 ;
        RECT 27.845 110.070 28.035 110.275 ;
        RECT 28.765 110.155 28.935 110.735 ;
        RECT 29.125 110.705 29.365 111.515 ;
        RECT 29.535 110.705 29.865 111.345 ;
        RECT 30.035 110.705 30.305 111.515 ;
        RECT 31.495 110.965 31.665 111.255 ;
        RECT 31.835 111.135 32.165 111.515 ;
        RECT 31.495 110.795 32.160 110.965 ;
        RECT 29.105 110.275 29.455 110.525 ;
        RECT 28.720 110.105 28.935 110.155 ;
        RECT 29.625 110.105 29.795 110.705 ;
        RECT 29.965 110.275 30.315 110.525 ;
        RECT 27.140 109.695 28.035 110.070 ;
        RECT 28.545 110.025 28.935 110.105 ;
        RECT 26.085 109.265 26.970 109.435 ;
        RECT 27.150 108.965 27.465 109.465 ;
        RECT 27.695 109.135 28.035 109.695 ;
        RECT 28.205 108.965 28.375 109.975 ;
        RECT 28.545 109.180 28.875 110.025 ;
        RECT 29.115 109.935 29.795 110.105 ;
        RECT 29.115 109.150 29.445 109.935 ;
        RECT 29.975 108.965 30.305 110.105 ;
        RECT 31.410 109.975 31.760 110.625 ;
        RECT 31.930 109.805 32.160 110.795 ;
        RECT 31.495 109.635 32.160 109.805 ;
        RECT 31.495 109.135 31.665 109.635 ;
        RECT 31.835 108.965 32.165 109.465 ;
        RECT 32.335 109.135 32.520 111.255 ;
        RECT 32.775 111.055 33.025 111.515 ;
        RECT 33.195 111.065 33.530 111.235 ;
        RECT 33.725 111.065 34.400 111.235 ;
        RECT 33.195 110.925 33.365 111.065 ;
        RECT 32.690 109.935 32.970 110.885 ;
        RECT 33.140 110.795 33.365 110.925 ;
        RECT 33.140 109.690 33.310 110.795 ;
        RECT 33.535 110.645 34.060 110.865 ;
        RECT 33.480 109.880 33.720 110.475 ;
        RECT 33.890 109.945 34.060 110.645 ;
        RECT 34.230 110.285 34.400 111.065 ;
        RECT 34.720 111.015 35.090 111.515 ;
        RECT 35.270 111.065 35.675 111.235 ;
        RECT 35.845 111.065 36.630 111.235 ;
        RECT 35.270 110.835 35.440 111.065 ;
        RECT 34.610 110.535 35.440 110.835 ;
        RECT 35.825 110.565 36.290 110.895 ;
        RECT 34.610 110.505 34.810 110.535 ;
        RECT 34.930 110.285 35.100 110.355 ;
        RECT 34.230 110.115 35.100 110.285 ;
        RECT 34.590 110.025 35.100 110.115 ;
        RECT 33.140 109.560 33.445 109.690 ;
        RECT 33.890 109.580 34.420 109.945 ;
        RECT 32.760 108.965 33.025 109.425 ;
        RECT 33.195 109.135 33.445 109.560 ;
        RECT 34.590 109.410 34.760 110.025 ;
        RECT 33.655 109.240 34.760 109.410 ;
        RECT 34.930 108.965 35.100 109.765 ;
        RECT 35.270 109.465 35.440 110.535 ;
        RECT 35.610 109.635 35.800 110.355 ;
        RECT 35.970 109.605 36.290 110.565 ;
        RECT 36.460 110.605 36.630 111.065 ;
        RECT 36.905 110.985 37.115 111.515 ;
        RECT 37.375 110.775 37.705 111.300 ;
        RECT 37.875 110.905 38.045 111.515 ;
        RECT 38.215 110.860 38.545 111.295 ;
        RECT 38.215 110.775 38.595 110.860 ;
        RECT 39.225 110.790 39.515 111.515 ;
        RECT 39.700 110.945 39.955 111.295 ;
        RECT 40.125 111.115 40.455 111.515 ;
        RECT 40.625 110.945 40.795 111.295 ;
        RECT 40.965 111.115 41.345 111.515 ;
        RECT 39.700 110.775 41.365 110.945 ;
        RECT 41.535 110.840 41.810 111.185 ;
        RECT 42.610 111.005 42.850 111.515 ;
        RECT 43.030 111.005 43.310 111.335 ;
        RECT 43.540 111.005 43.755 111.515 ;
        RECT 37.505 110.605 37.705 110.775 ;
        RECT 38.370 110.735 38.595 110.775 ;
        RECT 36.460 110.275 37.335 110.605 ;
        RECT 37.505 110.275 38.255 110.605 ;
        RECT 35.270 109.135 35.520 109.465 ;
        RECT 36.460 109.435 36.630 110.275 ;
        RECT 37.505 110.070 37.695 110.275 ;
        RECT 38.425 110.155 38.595 110.735 ;
        RECT 41.195 110.605 41.365 110.775 ;
        RECT 39.685 110.275 40.030 110.605 ;
        RECT 40.200 110.275 41.025 110.605 ;
        RECT 41.195 110.275 41.470 110.605 ;
        RECT 38.380 110.105 38.595 110.155 ;
        RECT 36.800 109.695 37.695 110.070 ;
        RECT 38.205 110.025 38.595 110.105 ;
        RECT 35.745 109.265 36.630 109.435 ;
        RECT 36.810 108.965 37.125 109.465 ;
        RECT 37.355 109.135 37.695 109.695 ;
        RECT 37.865 108.965 38.035 109.975 ;
        RECT 38.205 109.180 38.535 110.025 ;
        RECT 39.225 108.965 39.515 110.130 ;
        RECT 39.705 109.815 40.030 110.105 ;
        RECT 40.200 109.985 40.395 110.275 ;
        RECT 41.195 110.105 41.365 110.275 ;
        RECT 41.640 110.105 41.810 110.840 ;
        RECT 42.505 110.275 42.860 110.835 ;
        RECT 43.030 110.105 43.200 111.005 ;
        RECT 43.370 110.275 43.635 110.835 ;
        RECT 43.925 110.775 44.540 111.345 ;
        RECT 44.750 110.985 45.040 111.335 ;
        RECT 45.235 111.155 45.565 111.515 ;
        RECT 45.735 110.985 45.965 111.290 ;
        RECT 44.750 110.815 45.965 110.985 ;
        RECT 46.155 111.175 46.325 111.210 ;
        RECT 46.155 111.005 46.355 111.175 ;
        RECT 43.885 110.105 44.055 110.605 ;
        RECT 40.705 109.935 41.365 110.105 ;
        RECT 40.705 109.815 40.875 109.935 ;
        RECT 39.705 109.645 40.875 109.815 ;
        RECT 39.685 109.185 40.875 109.475 ;
        RECT 41.045 108.965 41.325 109.765 ;
        RECT 41.535 109.135 41.810 110.105 ;
        RECT 42.630 109.935 44.055 110.105 ;
        RECT 42.630 109.760 43.020 109.935 ;
        RECT 43.505 108.965 43.835 109.765 ;
        RECT 44.225 109.755 44.540 110.775 ;
        RECT 46.155 110.645 46.325 111.005 ;
        RECT 46.625 110.695 46.855 111.515 ;
        RECT 47.025 110.715 47.355 111.345 ;
        RECT 44.810 110.495 45.070 110.605 ;
        RECT 44.805 110.325 45.070 110.495 ;
        RECT 44.810 110.275 45.070 110.325 ;
        RECT 45.250 110.275 45.635 110.605 ;
        RECT 45.805 110.475 46.325 110.645 ;
        RECT 44.005 109.135 44.540 109.755 ;
        RECT 44.750 108.965 45.070 110.105 ;
        RECT 45.250 109.225 45.445 110.275 ;
        RECT 45.805 110.095 45.975 110.475 ;
        RECT 45.625 109.815 45.975 110.095 ;
        RECT 46.165 109.945 46.410 110.305 ;
        RECT 46.605 110.275 46.935 110.525 ;
        RECT 47.105 110.115 47.355 110.715 ;
        RECT 47.525 110.695 47.735 111.515 ;
        RECT 47.965 110.970 53.310 111.515 ;
        RECT 49.550 110.140 49.890 110.970 ;
        RECT 53.485 110.745 55.155 111.515 ;
        RECT 55.790 110.945 56.110 111.345 ;
        RECT 45.625 109.135 45.955 109.815 ;
        RECT 46.155 108.965 46.410 109.765 ;
        RECT 46.625 108.965 46.855 110.105 ;
        RECT 47.025 109.135 47.355 110.115 ;
        RECT 47.525 108.965 47.735 110.105 ;
        RECT 51.370 109.400 51.720 110.650 ;
        RECT 53.485 110.225 54.235 110.745 ;
        RECT 54.405 110.055 55.155 110.575 ;
        RECT 47.965 108.965 53.310 109.400 ;
        RECT 53.485 108.965 55.155 110.055 ;
        RECT 55.790 110.155 55.960 110.945 ;
        RECT 56.280 110.695 56.590 111.515 ;
        RECT 56.760 110.885 57.090 111.345 ;
        RECT 57.260 111.055 57.510 111.515 ;
        RECT 57.700 111.135 59.750 111.345 ;
        RECT 57.700 110.885 58.450 110.965 ;
        RECT 56.760 110.695 58.450 110.885 ;
        RECT 58.620 110.695 58.790 111.135 ;
        RECT 58.960 110.695 59.750 110.965 ;
        RECT 56.130 110.325 56.480 110.525 ;
        RECT 56.760 110.325 57.440 110.525 ;
        RECT 57.650 110.325 58.840 110.525 ;
        RECT 59.020 110.155 59.350 110.525 ;
        RECT 55.790 109.985 59.350 110.155 ;
        RECT 55.790 109.535 55.960 109.985 ;
        RECT 59.550 109.815 59.750 110.695 ;
        RECT 59.925 110.745 61.595 111.515 ;
        RECT 62.225 110.885 62.565 111.345 ;
        RECT 62.735 111.055 62.905 111.515 ;
        RECT 63.535 111.080 63.895 111.345 ;
        RECT 63.540 111.075 63.895 111.080 ;
        RECT 63.545 111.065 63.895 111.075 ;
        RECT 63.550 111.060 63.895 111.065 ;
        RECT 63.555 111.050 63.895 111.060 ;
        RECT 64.135 111.055 64.305 111.515 ;
        RECT 63.560 111.045 63.895 111.050 ;
        RECT 63.570 111.035 63.895 111.045 ;
        RECT 63.580 111.025 63.895 111.035 ;
        RECT 63.075 110.885 63.405 110.965 ;
        RECT 59.925 110.225 60.675 110.745 ;
        RECT 62.225 110.695 63.405 110.885 ;
        RECT 63.595 110.885 63.895 111.025 ;
        RECT 63.595 110.695 64.305 110.885 ;
        RECT 60.845 110.055 61.595 110.575 ;
        RECT 55.790 109.135 56.110 109.535 ;
        RECT 56.280 108.965 56.590 109.765 ;
        RECT 56.760 109.645 59.750 109.815 ;
        RECT 56.760 109.595 57.930 109.645 ;
        RECT 56.760 109.135 57.090 109.595 ;
        RECT 57.260 108.965 57.430 109.425 ;
        RECT 57.600 109.135 57.930 109.595 ;
        RECT 58.960 109.595 59.750 109.645 ;
        RECT 58.100 108.965 58.350 109.425 ;
        RECT 58.540 108.965 58.790 109.425 ;
        RECT 58.960 109.135 59.210 109.595 ;
        RECT 59.460 108.965 59.750 109.425 ;
        RECT 59.925 108.965 61.595 110.055 ;
        RECT 62.225 110.325 62.555 110.525 ;
        RECT 62.865 110.505 63.195 110.525 ;
        RECT 62.745 110.325 63.195 110.505 ;
        RECT 62.225 109.985 62.455 110.325 ;
        RECT 62.235 108.965 62.565 109.685 ;
        RECT 62.745 109.210 62.960 110.325 ;
        RECT 63.365 110.295 63.835 110.525 ;
        RECT 64.020 110.125 64.305 110.695 ;
        RECT 64.475 110.570 64.815 111.345 ;
        RECT 64.985 110.790 65.275 111.515 ;
        RECT 65.530 110.945 65.705 111.345 ;
        RECT 65.875 111.135 66.205 111.515 ;
        RECT 66.450 111.015 66.680 111.345 ;
        RECT 65.530 110.775 66.160 110.945 ;
        RECT 65.990 110.605 66.160 110.775 ;
        RECT 63.155 109.910 64.305 110.125 ;
        RECT 63.155 109.135 63.485 109.910 ;
        RECT 63.655 108.965 64.365 109.740 ;
        RECT 64.535 109.135 64.815 110.570 ;
        RECT 64.985 108.965 65.275 110.130 ;
        RECT 65.445 109.925 65.810 110.605 ;
        RECT 65.990 110.275 66.340 110.605 ;
        RECT 65.990 109.755 66.160 110.275 ;
        RECT 65.530 109.585 66.160 109.755 ;
        RECT 66.510 109.725 66.680 111.015 ;
        RECT 66.880 109.905 67.160 111.180 ;
        RECT 67.385 111.175 67.655 111.180 ;
        RECT 67.345 111.005 67.655 111.175 ;
        RECT 68.115 111.135 68.445 111.515 ;
        RECT 68.615 111.260 68.950 111.305 ;
        RECT 67.385 109.905 67.655 111.005 ;
        RECT 67.845 109.905 68.185 110.935 ;
        RECT 68.615 110.795 68.955 111.260 ;
        RECT 68.355 110.275 68.615 110.605 ;
        RECT 68.355 109.725 68.525 110.275 ;
        RECT 68.785 110.105 68.955 110.795 ;
        RECT 65.530 109.135 65.705 109.585 ;
        RECT 66.510 109.555 68.525 109.725 ;
        RECT 65.875 108.965 66.205 109.405 ;
        RECT 66.510 109.135 66.680 109.555 ;
        RECT 66.915 108.965 67.585 109.375 ;
        RECT 67.800 109.135 67.970 109.555 ;
        RECT 68.170 108.965 68.500 109.375 ;
        RECT 68.695 109.135 68.955 110.105 ;
        RECT 70.045 110.775 70.430 111.345 ;
        RECT 70.600 111.055 70.925 111.515 ;
        RECT 71.445 110.885 71.725 111.345 ;
        RECT 70.045 110.105 70.325 110.775 ;
        RECT 70.600 110.715 71.725 110.885 ;
        RECT 70.600 110.605 71.050 110.715 ;
        RECT 70.495 110.275 71.050 110.605 ;
        RECT 71.915 110.545 72.315 111.345 ;
        RECT 72.715 111.055 72.985 111.515 ;
        RECT 73.155 110.885 73.440 111.345 ;
        RECT 73.725 111.125 74.985 111.305 ;
        RECT 70.045 109.135 70.430 110.105 ;
        RECT 70.600 109.815 71.050 110.275 ;
        RECT 71.220 109.985 72.315 110.545 ;
        RECT 70.600 109.595 71.725 109.815 ;
        RECT 70.600 108.965 70.925 109.425 ;
        RECT 71.445 109.135 71.725 109.595 ;
        RECT 71.915 109.135 72.315 109.985 ;
        RECT 72.485 110.715 73.440 110.885 ;
        RECT 72.485 109.815 72.695 110.715 ;
        RECT 72.865 109.985 73.555 110.545 ;
        RECT 72.485 109.595 73.440 109.815 ;
        RECT 73.725 109.610 73.965 110.935 ;
        RECT 74.135 110.775 74.485 110.955 ;
        RECT 74.655 110.905 74.985 111.125 ;
        RECT 75.175 111.075 75.345 111.515 ;
        RECT 75.515 110.905 75.855 111.320 ;
        RECT 74.655 110.775 75.855 110.905 ;
        RECT 74.135 109.765 74.305 110.775 ;
        RECT 74.825 110.735 75.855 110.775 ;
        RECT 76.025 110.745 79.535 111.515 ;
        RECT 79.795 110.965 79.965 111.255 ;
        RECT 80.135 111.135 80.465 111.515 ;
        RECT 79.795 110.795 80.460 110.965 ;
        RECT 74.475 110.185 74.645 110.605 ;
        RECT 74.860 110.355 75.225 110.525 ;
        RECT 74.475 109.935 74.875 110.185 ;
        RECT 75.045 110.155 75.225 110.355 ;
        RECT 75.395 110.325 75.855 110.525 ;
        RECT 76.025 110.225 77.675 110.745 ;
        RECT 75.045 109.985 75.365 110.155 ;
        RECT 72.715 108.965 72.985 109.425 ;
        RECT 73.155 109.135 73.440 109.595 ;
        RECT 74.135 109.555 74.975 109.765 ;
        RECT 73.775 108.965 73.985 109.425 ;
        RECT 74.475 109.135 74.975 109.555 ;
        RECT 75.165 109.195 75.365 109.985 ;
        RECT 75.535 108.965 75.855 110.145 ;
        RECT 77.845 110.055 79.535 110.575 ;
        RECT 76.025 108.965 79.535 110.055 ;
        RECT 79.710 109.975 80.060 110.625 ;
        RECT 80.230 109.805 80.460 110.795 ;
        RECT 79.795 109.635 80.460 109.805 ;
        RECT 79.795 109.135 79.965 109.635 ;
        RECT 80.135 108.965 80.465 109.465 ;
        RECT 80.635 109.135 80.820 111.255 ;
        RECT 81.075 111.055 81.325 111.515 ;
        RECT 81.495 111.065 81.830 111.235 ;
        RECT 82.025 111.065 82.700 111.235 ;
        RECT 81.495 110.925 81.665 111.065 ;
        RECT 80.990 109.935 81.270 110.885 ;
        RECT 81.440 110.795 81.665 110.925 ;
        RECT 81.440 109.690 81.610 110.795 ;
        RECT 81.835 110.645 82.360 110.865 ;
        RECT 81.780 109.880 82.020 110.475 ;
        RECT 82.190 109.945 82.360 110.645 ;
        RECT 82.530 110.285 82.700 111.065 ;
        RECT 83.020 111.015 83.390 111.515 ;
        RECT 83.570 111.065 83.975 111.235 ;
        RECT 84.145 111.065 84.930 111.235 ;
        RECT 83.570 110.835 83.740 111.065 ;
        RECT 82.910 110.535 83.740 110.835 ;
        RECT 84.125 110.565 84.590 110.895 ;
        RECT 82.910 110.505 83.110 110.535 ;
        RECT 83.230 110.285 83.400 110.355 ;
        RECT 82.530 110.115 83.400 110.285 ;
        RECT 82.890 110.025 83.400 110.115 ;
        RECT 81.440 109.560 81.745 109.690 ;
        RECT 82.190 109.580 82.720 109.945 ;
        RECT 81.060 108.965 81.325 109.425 ;
        RECT 81.495 109.135 81.745 109.560 ;
        RECT 82.890 109.410 83.060 110.025 ;
        RECT 81.955 109.240 83.060 109.410 ;
        RECT 83.230 108.965 83.400 109.765 ;
        RECT 83.570 109.465 83.740 110.535 ;
        RECT 83.910 109.635 84.100 110.355 ;
        RECT 84.270 109.605 84.590 110.565 ;
        RECT 84.760 110.605 84.930 111.065 ;
        RECT 85.205 110.985 85.415 111.515 ;
        RECT 85.675 110.775 86.005 111.300 ;
        RECT 86.175 110.905 86.345 111.515 ;
        RECT 86.515 110.860 86.845 111.295 ;
        RECT 86.515 110.775 86.895 110.860 ;
        RECT 85.805 110.605 86.005 110.775 ;
        RECT 86.670 110.735 86.895 110.775 ;
        RECT 84.760 110.275 85.635 110.605 ;
        RECT 85.805 110.275 86.555 110.605 ;
        RECT 83.570 109.135 83.820 109.465 ;
        RECT 84.760 109.435 84.930 110.275 ;
        RECT 85.805 110.070 85.995 110.275 ;
        RECT 86.725 110.155 86.895 110.735 ;
        RECT 86.680 110.105 86.895 110.155 ;
        RECT 85.100 109.695 85.995 110.070 ;
        RECT 86.505 110.025 86.895 110.105 ;
        RECT 87.065 110.775 87.450 111.345 ;
        RECT 87.620 111.055 87.945 111.515 ;
        RECT 88.465 110.885 88.745 111.345 ;
        RECT 87.065 110.105 87.345 110.775 ;
        RECT 87.620 110.715 88.745 110.885 ;
        RECT 87.620 110.605 88.070 110.715 ;
        RECT 87.515 110.275 88.070 110.605 ;
        RECT 88.935 110.545 89.335 111.345 ;
        RECT 89.735 111.055 90.005 111.515 ;
        RECT 90.175 110.885 90.460 111.345 ;
        RECT 84.045 109.265 84.930 109.435 ;
        RECT 85.110 108.965 85.425 109.465 ;
        RECT 85.655 109.135 85.995 109.695 ;
        RECT 86.165 108.965 86.335 109.975 ;
        RECT 86.505 109.180 86.835 110.025 ;
        RECT 87.065 109.135 87.450 110.105 ;
        RECT 87.620 109.815 88.070 110.275 ;
        RECT 88.240 109.985 89.335 110.545 ;
        RECT 87.620 109.595 88.745 109.815 ;
        RECT 87.620 108.965 87.945 109.425 ;
        RECT 88.465 109.135 88.745 109.595 ;
        RECT 88.935 109.135 89.335 109.985 ;
        RECT 89.505 110.715 90.460 110.885 ;
        RECT 90.745 110.765 91.955 111.515 ;
        RECT 89.505 109.815 89.715 110.715 ;
        RECT 89.885 109.985 90.575 110.545 ;
        RECT 90.745 110.055 91.265 110.595 ;
        RECT 91.435 110.225 91.955 110.765 ;
        RECT 100.090 110.950 100.760 114.210 ;
        RECT 101.430 113.640 105.470 113.810 ;
        RECT 101.090 111.580 101.260 113.580 ;
        RECT 105.640 111.580 105.810 113.580 ;
        RECT 101.430 111.350 105.470 111.520 ;
        RECT 106.150 110.950 106.320 114.210 ;
        RECT 100.090 110.780 106.320 110.950 ;
        RECT 89.505 109.595 90.460 109.815 ;
        RECT 89.735 108.965 90.005 109.425 ;
        RECT 90.175 109.135 90.460 109.595 ;
        RECT 90.745 108.965 91.955 110.055 ;
        RECT 13.380 108.795 92.040 108.965 ;
        RECT 13.465 107.705 14.675 108.795 ;
        RECT 14.935 108.125 15.105 108.625 ;
        RECT 15.275 108.295 15.605 108.795 ;
        RECT 14.935 107.955 15.600 108.125 ;
        RECT 13.465 106.995 13.985 107.535 ;
        RECT 14.155 107.165 14.675 107.705 ;
        RECT 14.850 107.135 15.200 107.785 ;
        RECT 13.465 106.245 14.675 106.995 ;
        RECT 15.370 106.965 15.600 107.955 ;
        RECT 14.935 106.795 15.600 106.965 ;
        RECT 14.935 106.505 15.105 106.795 ;
        RECT 15.275 106.245 15.605 106.625 ;
        RECT 15.775 106.505 15.960 108.625 ;
        RECT 16.200 108.335 16.465 108.795 ;
        RECT 16.635 108.200 16.885 108.625 ;
        RECT 17.095 108.350 18.200 108.520 ;
        RECT 16.580 108.070 16.885 108.200 ;
        RECT 16.130 106.875 16.410 107.825 ;
        RECT 16.580 106.965 16.750 108.070 ;
        RECT 16.920 107.285 17.160 107.880 ;
        RECT 17.330 107.815 17.860 108.180 ;
        RECT 17.330 107.115 17.500 107.815 ;
        RECT 18.030 107.735 18.200 108.350 ;
        RECT 18.370 107.995 18.540 108.795 ;
        RECT 18.710 108.295 18.960 108.625 ;
        RECT 19.185 108.325 20.070 108.495 ;
        RECT 18.030 107.645 18.540 107.735 ;
        RECT 16.580 106.835 16.805 106.965 ;
        RECT 16.975 106.895 17.500 107.115 ;
        RECT 17.670 107.475 18.540 107.645 ;
        RECT 16.215 106.245 16.465 106.705 ;
        RECT 16.635 106.695 16.805 106.835 ;
        RECT 17.670 106.695 17.840 107.475 ;
        RECT 18.370 107.405 18.540 107.475 ;
        RECT 18.050 107.225 18.250 107.255 ;
        RECT 18.710 107.225 18.880 108.295 ;
        RECT 19.050 107.405 19.240 108.125 ;
        RECT 18.050 106.925 18.880 107.225 ;
        RECT 19.410 107.195 19.730 108.155 ;
        RECT 16.635 106.525 16.970 106.695 ;
        RECT 17.165 106.525 17.840 106.695 ;
        RECT 18.160 106.245 18.530 106.745 ;
        RECT 18.710 106.695 18.880 106.925 ;
        RECT 19.265 106.865 19.730 107.195 ;
        RECT 19.900 107.485 20.070 108.325 ;
        RECT 20.250 108.295 20.565 108.795 ;
        RECT 20.795 108.065 21.135 108.625 ;
        RECT 20.240 107.690 21.135 108.065 ;
        RECT 21.305 107.785 21.475 108.795 ;
        RECT 20.945 107.485 21.135 107.690 ;
        RECT 21.645 107.735 21.975 108.580 ;
        RECT 21.645 107.655 22.035 107.735 ;
        RECT 22.210 107.655 22.530 108.795 ;
        RECT 21.820 107.605 22.035 107.655 ;
        RECT 19.900 107.155 20.775 107.485 ;
        RECT 20.945 107.155 21.695 107.485 ;
        RECT 19.900 106.695 20.070 107.155 ;
        RECT 20.945 106.985 21.145 107.155 ;
        RECT 21.865 107.025 22.035 107.605 ;
        RECT 22.710 107.485 22.905 108.535 ;
        RECT 23.085 107.945 23.415 108.625 ;
        RECT 23.615 107.995 23.870 108.795 ;
        RECT 24.080 108.005 24.615 108.625 ;
        RECT 23.085 107.665 23.435 107.945 ;
        RECT 22.270 107.435 22.530 107.485 ;
        RECT 22.265 107.265 22.530 107.435 ;
        RECT 22.270 107.155 22.530 107.265 ;
        RECT 22.710 107.155 23.095 107.485 ;
        RECT 23.265 107.285 23.435 107.665 ;
        RECT 23.625 107.455 23.870 107.815 ;
        RECT 23.265 107.115 23.785 107.285 ;
        RECT 21.810 106.985 22.035 107.025 ;
        RECT 18.710 106.525 19.115 106.695 ;
        RECT 19.285 106.525 20.070 106.695 ;
        RECT 20.345 106.245 20.555 106.775 ;
        RECT 20.815 106.460 21.145 106.985 ;
        RECT 21.655 106.900 22.035 106.985 ;
        RECT 21.315 106.245 21.485 106.855 ;
        RECT 21.655 106.465 21.985 106.900 ;
        RECT 22.210 106.775 23.425 106.945 ;
        RECT 22.210 106.425 22.500 106.775 ;
        RECT 22.695 106.245 23.025 106.605 ;
        RECT 23.195 106.470 23.425 106.775 ;
        RECT 23.615 106.550 23.785 107.115 ;
        RECT 24.080 106.985 24.395 108.005 ;
        RECT 24.785 107.995 25.115 108.795 ;
        RECT 25.600 107.825 25.990 108.000 ;
        RECT 24.565 107.655 25.990 107.825 ;
        RECT 24.565 107.155 24.735 107.655 ;
        RECT 24.080 106.415 24.695 106.985 ;
        RECT 24.985 106.925 25.250 107.485 ;
        RECT 25.420 106.755 25.590 107.655 ;
        RECT 26.345 107.630 26.635 108.795 ;
        RECT 27.725 108.285 28.925 108.525 ;
        RECT 29.105 108.370 29.435 108.795 ;
        RECT 29.950 108.370 30.310 108.795 ;
        RECT 30.515 108.200 30.775 108.380 ;
        RECT 29.140 108.115 30.775 108.200 ;
        RECT 27.725 107.655 28.030 108.085 ;
        RECT 28.200 108.030 30.775 108.115 ;
        RECT 28.200 107.945 29.310 108.030 ;
        RECT 30.095 107.970 30.775 108.030 ;
        RECT 25.760 106.925 26.115 107.485 ;
        RECT 27.725 106.985 27.895 107.655 ;
        RECT 28.200 107.485 28.370 107.945 ;
        RECT 28.070 107.155 28.370 107.485 ;
        RECT 28.630 107.235 29.165 107.775 ;
        RECT 29.530 107.655 29.925 107.860 ;
        RECT 29.415 107.095 29.585 107.485 ;
        RECT 29.265 107.065 29.585 107.095 ;
        RECT 28.700 106.985 29.585 107.065 ;
        RECT 24.865 106.245 25.080 106.755 ;
        RECT 25.310 106.425 25.590 106.755 ;
        RECT 25.770 106.245 26.010 106.755 ;
        RECT 26.345 106.245 26.635 106.970 ;
        RECT 27.725 106.925 29.585 106.985 ;
        RECT 27.725 106.895 29.435 106.925 ;
        RECT 27.725 106.815 28.870 106.895 ;
        RECT 27.725 106.765 28.030 106.815 ;
        RECT 27.775 106.465 28.030 106.765 ;
        RECT 28.200 106.245 28.530 106.645 ;
        RECT 28.700 106.465 28.870 106.815 ;
        RECT 29.755 106.755 29.925 107.655 ;
        RECT 30.095 107.065 30.265 107.970 ;
        RECT 30.435 107.235 30.775 107.800 ;
        RECT 30.950 107.655 31.225 108.625 ;
        RECT 31.435 107.995 31.715 108.795 ;
        RECT 31.885 108.285 33.075 108.575 ;
        RECT 31.885 107.945 33.055 108.115 ;
        RECT 31.885 107.825 32.055 107.945 ;
        RECT 31.395 107.655 32.055 107.825 ;
        RECT 30.095 106.895 30.775 107.065 ;
        RECT 29.170 106.245 29.340 106.725 ;
        RECT 29.575 106.425 29.925 106.755 ;
        RECT 30.095 106.245 30.265 106.725 ;
        RECT 30.515 106.450 30.775 106.895 ;
        RECT 30.950 106.920 31.120 107.655 ;
        RECT 31.395 107.485 31.565 107.655 ;
        RECT 32.365 107.485 32.560 107.775 ;
        RECT 32.730 107.655 33.055 107.945 ;
        RECT 33.245 107.705 34.915 108.795 ;
        RECT 31.290 107.155 31.565 107.485 ;
        RECT 31.735 107.155 32.560 107.485 ;
        RECT 32.730 107.155 33.075 107.485 ;
        RECT 31.395 106.985 31.565 107.155 ;
        RECT 33.245 107.015 33.995 107.535 ;
        RECT 34.165 107.185 34.915 107.705 ;
        RECT 35.545 107.655 35.825 108.795 ;
        RECT 35.995 107.645 36.325 108.625 ;
        RECT 36.495 107.655 36.755 108.795 ;
        RECT 36.925 107.655 37.200 108.625 ;
        RECT 37.410 107.995 37.690 108.795 ;
        RECT 37.860 108.285 39.475 108.615 ;
        RECT 37.860 107.945 39.035 108.115 ;
        RECT 37.860 107.825 38.030 107.945 ;
        RECT 37.370 107.655 38.030 107.825 ;
        RECT 35.555 107.215 35.890 107.485 ;
        RECT 36.060 107.045 36.230 107.645 ;
        RECT 36.400 107.235 36.735 107.485 ;
        RECT 30.950 106.575 31.225 106.920 ;
        RECT 31.395 106.815 33.060 106.985 ;
        RECT 31.415 106.245 31.795 106.645 ;
        RECT 31.965 106.465 32.135 106.815 ;
        RECT 32.305 106.245 32.635 106.645 ;
        RECT 32.805 106.465 33.060 106.815 ;
        RECT 33.245 106.245 34.915 107.015 ;
        RECT 35.545 106.245 35.855 107.045 ;
        RECT 36.060 106.415 36.755 107.045 ;
        RECT 36.925 106.920 37.095 107.655 ;
        RECT 37.370 107.485 37.540 107.655 ;
        RECT 38.290 107.485 38.535 107.775 ;
        RECT 38.705 107.655 39.035 107.945 ;
        RECT 39.295 107.485 39.465 108.045 ;
        RECT 39.715 107.655 39.975 108.795 ;
        RECT 40.145 107.655 40.530 108.625 ;
        RECT 40.700 108.335 41.025 108.795 ;
        RECT 41.545 108.165 41.825 108.625 ;
        RECT 40.700 107.945 41.825 108.165 ;
        RECT 37.265 107.155 37.540 107.485 ;
        RECT 37.710 107.155 38.535 107.485 ;
        RECT 38.750 107.155 39.465 107.485 ;
        RECT 39.635 107.235 39.970 107.485 ;
        RECT 37.370 106.985 37.540 107.155 ;
        RECT 39.215 107.065 39.465 107.155 ;
        RECT 36.925 106.575 37.200 106.920 ;
        RECT 37.370 106.815 39.035 106.985 ;
        RECT 37.390 106.245 37.765 106.645 ;
        RECT 37.935 106.465 38.105 106.815 ;
        RECT 38.275 106.245 38.605 106.645 ;
        RECT 38.775 106.415 39.035 106.815 ;
        RECT 39.215 106.645 39.545 107.065 ;
        RECT 39.715 106.245 39.975 107.065 ;
        RECT 40.145 106.985 40.425 107.655 ;
        RECT 40.700 107.485 41.150 107.945 ;
        RECT 42.015 107.775 42.415 108.625 ;
        RECT 42.815 108.335 43.085 108.795 ;
        RECT 43.255 108.165 43.540 108.625 ;
        RECT 40.595 107.155 41.150 107.485 ;
        RECT 41.320 107.215 42.415 107.775 ;
        RECT 40.700 107.045 41.150 107.155 ;
        RECT 40.145 106.415 40.530 106.985 ;
        RECT 40.700 106.875 41.825 107.045 ;
        RECT 40.700 106.245 41.025 106.705 ;
        RECT 41.545 106.415 41.825 106.875 ;
        RECT 42.015 106.415 42.415 107.215 ;
        RECT 42.585 107.945 43.540 108.165 ;
        RECT 44.025 108.125 44.305 108.795 ;
        RECT 42.585 107.045 42.795 107.945 ;
        RECT 44.475 107.905 44.775 108.455 ;
        RECT 44.975 108.075 45.305 108.795 ;
        RECT 45.495 108.075 45.955 108.625 ;
        RECT 42.965 107.215 43.655 107.775 ;
        RECT 43.840 107.485 44.105 107.845 ;
        RECT 44.475 107.735 45.415 107.905 ;
        RECT 45.245 107.485 45.415 107.735 ;
        RECT 43.840 107.235 44.515 107.485 ;
        RECT 44.735 107.235 45.075 107.485 ;
        RECT 45.245 107.155 45.535 107.485 ;
        RECT 45.245 107.065 45.415 107.155 ;
        RECT 42.585 106.875 43.540 107.045 ;
        RECT 42.815 106.245 43.085 106.705 ;
        RECT 43.255 106.415 43.540 106.875 ;
        RECT 44.025 106.875 45.415 107.065 ;
        RECT 44.025 106.515 44.355 106.875 ;
        RECT 45.705 106.705 45.955 108.075 ;
        RECT 46.125 107.705 49.635 108.795 ;
        RECT 49.805 108.240 50.410 108.795 ;
        RECT 50.585 108.285 51.065 108.625 ;
        RECT 51.235 108.250 51.490 108.795 ;
        RECT 49.805 108.140 50.420 108.240 ;
        RECT 50.235 108.115 50.420 108.140 ;
        RECT 44.975 106.245 45.225 106.705 ;
        RECT 45.395 106.415 45.955 106.705 ;
        RECT 46.125 107.015 47.775 107.535 ;
        RECT 47.945 107.185 49.635 107.705 ;
        RECT 49.805 107.520 50.065 107.970 ;
        RECT 50.235 107.870 50.565 108.115 ;
        RECT 50.735 107.795 51.490 108.045 ;
        RECT 51.660 107.925 51.935 108.625 ;
        RECT 50.720 107.760 51.490 107.795 ;
        RECT 50.705 107.750 51.490 107.760 ;
        RECT 50.700 107.735 51.595 107.750 ;
        RECT 50.680 107.720 51.595 107.735 ;
        RECT 50.660 107.710 51.595 107.720 ;
        RECT 50.635 107.700 51.595 107.710 ;
        RECT 50.565 107.670 51.595 107.700 ;
        RECT 50.545 107.640 51.595 107.670 ;
        RECT 50.525 107.610 51.595 107.640 ;
        RECT 50.495 107.585 51.595 107.610 ;
        RECT 50.460 107.550 51.595 107.585 ;
        RECT 50.430 107.545 51.595 107.550 ;
        RECT 50.430 107.540 50.820 107.545 ;
        RECT 50.430 107.530 50.795 107.540 ;
        RECT 50.430 107.525 50.780 107.530 ;
        RECT 50.430 107.520 50.765 107.525 ;
        RECT 49.805 107.515 50.765 107.520 ;
        RECT 49.805 107.505 50.755 107.515 ;
        RECT 49.805 107.500 50.745 107.505 ;
        RECT 49.805 107.490 50.735 107.500 ;
        RECT 49.805 107.480 50.730 107.490 ;
        RECT 49.805 107.475 50.725 107.480 ;
        RECT 49.805 107.460 50.715 107.475 ;
        RECT 49.805 107.445 50.710 107.460 ;
        RECT 49.805 107.420 50.700 107.445 ;
        RECT 49.805 107.350 50.695 107.420 ;
        RECT 46.125 106.245 49.635 107.015 ;
        RECT 49.805 106.795 50.355 107.180 ;
        RECT 50.525 106.625 50.695 107.350 ;
        RECT 49.805 106.455 50.695 106.625 ;
        RECT 50.865 106.950 51.195 107.375 ;
        RECT 51.365 107.150 51.595 107.545 ;
        RECT 50.865 106.465 51.085 106.950 ;
        RECT 51.765 106.895 51.935 107.925 ;
        RECT 52.105 107.630 52.395 108.795 ;
        RECT 52.575 107.985 52.870 108.795 ;
        RECT 53.050 107.485 53.295 108.625 ;
        RECT 53.470 107.985 53.730 108.795 ;
        RECT 54.330 108.790 60.605 108.795 ;
        RECT 53.910 107.485 54.160 108.620 ;
        RECT 54.330 107.995 54.590 108.790 ;
        RECT 54.760 107.895 55.020 108.620 ;
        RECT 55.190 108.065 55.450 108.790 ;
        RECT 55.620 107.895 55.880 108.620 ;
        RECT 56.050 108.065 56.310 108.790 ;
        RECT 56.480 107.895 56.740 108.620 ;
        RECT 56.910 108.065 57.170 108.790 ;
        RECT 57.340 107.895 57.600 108.620 ;
        RECT 57.770 108.065 58.015 108.790 ;
        RECT 58.185 107.895 58.445 108.620 ;
        RECT 58.630 108.065 58.875 108.790 ;
        RECT 59.045 107.895 59.305 108.620 ;
        RECT 59.490 108.065 59.735 108.790 ;
        RECT 59.905 107.895 60.165 108.620 ;
        RECT 60.350 108.065 60.605 108.790 ;
        RECT 54.760 107.880 60.165 107.895 ;
        RECT 60.775 107.880 61.065 108.620 ;
        RECT 61.235 108.050 61.505 108.795 ;
        RECT 54.760 107.655 61.505 107.880 ;
        RECT 61.765 107.705 65.275 108.795 ;
        RECT 51.255 106.245 51.505 106.785 ;
        RECT 51.675 106.415 51.935 106.895 ;
        RECT 52.105 106.245 52.395 106.970 ;
        RECT 52.565 106.925 52.880 107.485 ;
        RECT 53.050 107.235 60.170 107.485 ;
        RECT 52.565 106.245 52.870 106.755 ;
        RECT 53.050 106.425 53.300 107.235 ;
        RECT 53.470 106.245 53.730 106.770 ;
        RECT 53.910 106.425 54.160 107.235 ;
        RECT 60.340 107.065 61.505 107.655 ;
        RECT 54.760 106.895 61.505 107.065 ;
        RECT 61.765 107.015 63.415 107.535 ;
        RECT 63.585 107.185 65.275 107.705 ;
        RECT 66.405 107.655 66.635 108.795 ;
        RECT 66.805 107.645 67.135 108.625 ;
        RECT 67.305 107.655 67.515 108.795 ;
        RECT 67.745 107.705 68.955 108.795 ;
        RECT 66.385 107.235 66.715 107.485 ;
        RECT 54.330 106.245 54.590 106.805 ;
        RECT 54.760 106.440 55.020 106.895 ;
        RECT 55.190 106.245 55.450 106.725 ;
        RECT 55.620 106.440 55.880 106.895 ;
        RECT 56.050 106.245 56.310 106.725 ;
        RECT 56.480 106.440 56.740 106.895 ;
        RECT 56.910 106.245 57.155 106.725 ;
        RECT 57.325 106.440 57.600 106.895 ;
        RECT 57.770 106.245 58.015 106.725 ;
        RECT 58.185 106.440 58.445 106.895 ;
        RECT 58.625 106.245 58.875 106.725 ;
        RECT 59.045 106.440 59.305 106.895 ;
        RECT 59.485 106.245 59.735 106.725 ;
        RECT 59.905 106.440 60.165 106.895 ;
        RECT 60.345 106.245 60.605 106.725 ;
        RECT 60.775 106.440 61.035 106.895 ;
        RECT 61.205 106.245 61.505 106.725 ;
        RECT 61.765 106.245 65.275 107.015 ;
        RECT 66.405 106.245 66.635 107.065 ;
        RECT 66.885 107.045 67.135 107.645 ;
        RECT 66.805 106.415 67.135 107.045 ;
        RECT 67.305 106.245 67.515 107.065 ;
        RECT 67.745 106.995 68.265 107.535 ;
        RECT 68.435 107.165 68.955 107.705 ;
        RECT 69.125 107.925 69.400 108.625 ;
        RECT 69.610 108.250 69.825 108.795 ;
        RECT 69.995 108.285 70.470 108.625 ;
        RECT 70.640 108.290 71.255 108.795 ;
        RECT 70.640 108.115 70.835 108.290 ;
        RECT 67.745 106.245 68.955 106.995 ;
        RECT 69.125 106.895 69.295 107.925 ;
        RECT 69.570 107.755 70.285 108.050 ;
        RECT 70.505 107.925 70.835 108.115 ;
        RECT 71.005 107.755 71.255 108.120 ;
        RECT 69.465 107.585 71.255 107.755 ;
        RECT 69.465 107.155 69.695 107.585 ;
        RECT 69.125 106.415 69.385 106.895 ;
        RECT 69.865 106.885 70.275 107.405 ;
        RECT 69.555 106.245 69.885 106.705 ;
        RECT 70.075 106.465 70.275 106.885 ;
        RECT 70.445 106.730 70.700 107.585 ;
        RECT 71.495 107.405 71.665 108.625 ;
        RECT 71.915 108.285 72.175 108.795 ;
        RECT 72.345 108.285 73.535 108.575 ;
        RECT 70.870 107.155 71.665 107.405 ;
        RECT 71.835 107.235 72.175 108.115 ;
        RECT 72.365 107.945 73.535 108.115 ;
        RECT 73.705 107.995 73.985 108.795 ;
        RECT 72.365 107.655 72.690 107.945 ;
        RECT 73.365 107.825 73.535 107.945 ;
        RECT 72.860 107.485 73.055 107.775 ;
        RECT 73.365 107.655 74.025 107.825 ;
        RECT 74.195 107.655 74.470 108.625 ;
        RECT 74.645 107.655 74.905 108.795 ;
        RECT 75.075 107.825 75.405 108.625 ;
        RECT 75.575 107.995 75.745 108.795 ;
        RECT 75.915 107.825 76.245 108.625 ;
        RECT 76.415 107.995 76.670 108.795 ;
        RECT 75.075 107.655 76.775 107.825 ;
        RECT 73.855 107.485 74.025 107.655 ;
        RECT 72.345 107.155 72.690 107.485 ;
        RECT 72.860 107.155 73.685 107.485 ;
        RECT 73.855 107.155 74.130 107.485 ;
        RECT 71.415 107.065 71.665 107.155 ;
        RECT 70.445 106.465 71.235 106.730 ;
        RECT 71.415 106.645 71.745 107.065 ;
        RECT 71.915 106.245 72.175 107.065 ;
        RECT 73.855 106.985 74.025 107.155 ;
        RECT 72.360 106.815 74.025 106.985 ;
        RECT 74.300 106.920 74.470 107.655 ;
        RECT 74.645 107.235 75.405 107.485 ;
        RECT 75.575 107.235 76.325 107.485 ;
        RECT 76.495 107.065 76.775 107.655 ;
        RECT 77.865 107.630 78.155 108.795 ;
        RECT 78.820 107.995 79.070 108.795 ;
        RECT 79.240 108.165 79.570 108.625 ;
        RECT 79.740 108.335 79.955 108.795 ;
        RECT 79.240 107.995 80.410 108.165 ;
        RECT 78.330 107.825 78.610 107.985 ;
        RECT 78.330 107.655 79.665 107.825 ;
        RECT 79.495 107.485 79.665 107.655 ;
        RECT 78.330 107.235 78.680 107.475 ;
        RECT 78.850 107.235 79.325 107.475 ;
        RECT 79.495 107.235 79.870 107.485 ;
        RECT 79.495 107.065 79.665 107.235 ;
        RECT 72.360 106.465 72.615 106.815 ;
        RECT 72.785 106.245 73.115 106.645 ;
        RECT 73.285 106.465 73.455 106.815 ;
        RECT 73.625 106.245 74.005 106.645 ;
        RECT 74.195 106.575 74.470 106.920 ;
        RECT 74.645 106.875 75.745 107.045 ;
        RECT 74.645 106.415 74.985 106.875 ;
        RECT 75.155 106.245 75.325 106.705 ;
        RECT 75.495 106.625 75.745 106.875 ;
        RECT 75.915 106.815 76.775 107.065 ;
        RECT 76.335 106.625 76.665 106.645 ;
        RECT 75.495 106.415 76.665 106.625 ;
        RECT 77.865 106.245 78.155 106.970 ;
        RECT 78.330 106.895 79.665 107.065 ;
        RECT 78.330 106.685 78.600 106.895 ;
        RECT 80.040 106.705 80.410 107.995 ;
        RECT 80.625 107.705 81.835 108.795 ;
        RECT 78.820 106.245 79.150 106.705 ;
        RECT 79.660 106.415 80.410 106.705 ;
        RECT 80.625 106.995 81.145 107.535 ;
        RECT 81.315 107.165 81.835 107.705 ;
        RECT 82.010 107.655 82.345 108.625 ;
        RECT 82.515 107.655 82.685 108.795 ;
        RECT 82.855 108.455 84.885 108.625 ;
        RECT 80.625 106.245 81.835 106.995 ;
        RECT 82.010 106.985 82.180 107.655 ;
        RECT 82.855 107.485 83.025 108.455 ;
        RECT 82.350 107.155 82.605 107.485 ;
        RECT 82.830 107.155 83.025 107.485 ;
        RECT 83.195 108.115 84.320 108.285 ;
        RECT 82.435 106.985 82.605 107.155 ;
        RECT 83.195 106.985 83.365 108.115 ;
        RECT 82.010 106.415 82.265 106.985 ;
        RECT 82.435 106.815 83.365 106.985 ;
        RECT 83.535 107.775 84.545 107.945 ;
        RECT 83.535 106.975 83.705 107.775 ;
        RECT 83.910 107.435 84.185 107.575 ;
        RECT 83.905 107.265 84.185 107.435 ;
        RECT 83.190 106.780 83.365 106.815 ;
        RECT 82.435 106.245 82.765 106.645 ;
        RECT 83.190 106.415 83.720 106.780 ;
        RECT 83.910 106.415 84.185 107.265 ;
        RECT 84.355 106.415 84.545 107.775 ;
        RECT 84.715 107.790 84.885 108.455 ;
        RECT 85.055 108.035 85.225 108.795 ;
        RECT 85.460 108.035 85.975 108.445 ;
        RECT 84.715 107.600 85.465 107.790 ;
        RECT 85.635 107.225 85.975 108.035 ;
        RECT 86.145 107.705 87.355 108.795 ;
        RECT 84.745 107.055 85.975 107.225 ;
        RECT 84.725 106.245 85.235 106.780 ;
        RECT 85.455 106.450 85.700 107.055 ;
        RECT 86.145 106.995 86.665 107.535 ;
        RECT 86.835 107.165 87.355 107.705 ;
        RECT 87.615 107.865 87.785 108.625 ;
        RECT 87.965 108.035 88.295 108.795 ;
        RECT 87.615 107.695 88.280 107.865 ;
        RECT 88.465 107.720 88.735 108.625 ;
        RECT 88.110 107.550 88.280 107.695 ;
        RECT 87.545 107.145 87.875 107.515 ;
        RECT 88.110 107.220 88.395 107.550 ;
        RECT 86.145 106.245 87.355 106.995 ;
        RECT 88.110 106.965 88.280 107.220 ;
        RECT 87.615 106.795 88.280 106.965 ;
        RECT 88.565 106.920 88.735 107.720 ;
        RECT 88.905 107.705 90.575 108.795 ;
        RECT 87.615 106.415 87.785 106.795 ;
        RECT 87.965 106.245 88.295 106.625 ;
        RECT 88.475 106.415 88.735 106.920 ;
        RECT 88.905 107.015 89.655 107.535 ;
        RECT 89.825 107.185 90.575 107.705 ;
        RECT 90.745 107.705 91.955 108.795 ;
        RECT 90.745 107.165 91.265 107.705 ;
        RECT 88.905 106.245 90.575 107.015 ;
        RECT 91.435 106.995 91.955 107.535 ;
        RECT 100.090 107.520 100.760 110.780 ;
        RECT 101.430 110.210 105.470 110.380 ;
        RECT 101.090 108.150 101.260 110.150 ;
        RECT 105.640 108.150 105.810 110.150 ;
        RECT 101.430 107.920 105.470 108.090 ;
        RECT 106.150 107.520 106.320 110.780 ;
        RECT 100.090 107.510 106.320 107.520 ;
        RECT 107.910 116.780 117.740 116.820 ;
        RECT 120.510 116.800 126.250 116.810 ;
        RECT 107.910 116.650 118.540 116.780 ;
        RECT 107.910 114.390 108.080 116.650 ;
        RECT 108.805 116.080 116.845 116.250 ;
        RECT 108.420 115.020 108.590 116.020 ;
        RECT 117.060 115.020 117.230 116.020 ;
        RECT 108.805 114.790 116.845 114.960 ;
        RECT 117.570 114.390 118.540 116.650 ;
        RECT 107.910 114.220 118.540 114.390 ;
        RECT 107.910 110.960 108.080 114.220 ;
        RECT 108.805 113.650 116.845 113.820 ;
        RECT 108.420 111.590 108.590 113.590 ;
        RECT 117.060 111.590 117.230 113.590 ;
        RECT 108.805 111.360 116.845 111.530 ;
        RECT 117.570 110.960 118.540 114.220 ;
        RECT 107.910 110.790 118.540 110.960 ;
        RECT 107.910 107.530 108.080 110.790 ;
        RECT 108.805 110.220 116.845 110.390 ;
        RECT 108.420 108.160 108.590 110.160 ;
        RECT 117.060 108.160 117.230 110.160 ;
        RECT 108.805 107.930 116.845 108.100 ;
        RECT 117.570 107.530 118.540 110.790 ;
        RECT 100.090 107.410 106.330 107.510 ;
        RECT 90.745 106.245 91.955 106.995 ;
        RECT 100.080 106.850 106.330 107.410 ;
        RECT 100.080 106.830 105.250 106.850 ;
        RECT 100.080 106.760 104.070 106.830 ;
        RECT 13.380 106.075 92.040 106.245 ;
        RECT 13.465 105.325 14.675 106.075 ;
        RECT 15.310 105.600 15.645 105.860 ;
        RECT 15.815 105.675 16.145 106.075 ;
        RECT 16.315 105.675 17.930 105.845 ;
        RECT 13.465 104.785 13.985 105.325 ;
        RECT 14.155 104.615 14.675 105.155 ;
        RECT 13.465 103.525 14.675 104.615 ;
        RECT 15.310 104.245 15.565 105.600 ;
        RECT 16.315 105.505 16.485 105.675 ;
        RECT 15.925 105.335 16.485 105.505 ;
        RECT 16.750 105.395 17.020 105.495 ;
        RECT 17.210 105.395 17.500 105.495 ;
        RECT 15.925 105.165 16.095 105.335 ;
        RECT 16.745 105.225 17.020 105.395 ;
        RECT 17.205 105.225 17.500 105.395 ;
        RECT 15.790 104.835 16.095 105.165 ;
        RECT 16.290 105.055 16.540 105.165 ;
        RECT 16.285 104.885 16.540 105.055 ;
        RECT 16.290 104.835 16.540 104.885 ;
        RECT 16.750 104.835 17.020 105.225 ;
        RECT 17.210 104.835 17.500 105.225 ;
        RECT 17.670 104.835 18.090 105.500 ;
        RECT 18.475 105.355 18.805 106.075 ;
        RECT 18.990 105.235 19.250 106.075 ;
        RECT 19.425 105.330 19.680 105.905 ;
        RECT 19.850 105.695 20.180 106.075 ;
        RECT 20.395 105.525 20.565 105.905 ;
        RECT 19.850 105.355 20.565 105.525 ;
        RECT 18.400 105.055 18.750 105.165 ;
        RECT 18.400 104.885 18.755 105.055 ;
        RECT 18.400 104.835 18.750 104.885 ;
        RECT 15.925 104.665 16.095 104.835 ;
        RECT 15.925 104.495 18.295 104.665 ;
        RECT 18.545 104.545 18.750 104.835 ;
        RECT 15.310 103.735 15.645 104.245 ;
        RECT 15.895 103.525 16.225 104.325 ;
        RECT 16.470 104.115 17.895 104.285 ;
        RECT 16.470 103.695 16.755 104.115 ;
        RECT 17.010 103.525 17.340 103.945 ;
        RECT 17.565 103.865 17.895 104.115 ;
        RECT 18.125 104.035 18.295 104.495 ;
        RECT 18.555 103.865 18.725 104.365 ;
        RECT 17.565 103.695 18.725 103.865 ;
        RECT 18.990 103.525 19.250 104.675 ;
        RECT 19.425 104.600 19.595 105.330 ;
        RECT 19.850 105.165 20.020 105.355 ;
        RECT 21.745 105.275 22.055 106.075 ;
        RECT 22.260 105.275 22.955 105.905 ;
        RECT 23.215 105.525 23.385 105.905 ;
        RECT 23.565 105.695 23.895 106.075 ;
        RECT 23.215 105.355 23.880 105.525 ;
        RECT 24.075 105.400 24.335 105.905 ;
        RECT 25.055 105.735 25.225 105.770 ;
        RECT 25.025 105.565 25.225 105.735 ;
        RECT 19.765 104.835 20.020 105.165 ;
        RECT 19.850 104.625 20.020 104.835 ;
        RECT 20.300 104.805 20.655 105.175 ;
        RECT 21.755 104.835 22.090 105.105 ;
        RECT 22.260 104.715 22.430 105.275 ;
        RECT 22.600 104.835 22.935 105.085 ;
        RECT 23.145 104.805 23.485 105.175 ;
        RECT 23.710 105.100 23.880 105.355 ;
        RECT 23.710 104.770 23.985 105.100 ;
        RECT 22.260 104.675 22.435 104.715 ;
        RECT 19.425 103.695 19.680 104.600 ;
        RECT 19.850 104.455 20.565 104.625 ;
        RECT 19.850 103.525 20.180 104.285 ;
        RECT 20.395 103.695 20.565 104.455 ;
        RECT 21.745 103.525 22.025 104.665 ;
        RECT 22.195 103.695 22.525 104.675 ;
        RECT 22.695 103.525 22.955 104.665 ;
        RECT 23.710 104.625 23.880 104.770 ;
        RECT 23.205 104.455 23.880 104.625 ;
        RECT 24.155 104.600 24.335 105.400 ;
        RECT 25.055 105.205 25.225 105.565 ;
        RECT 25.415 105.545 25.645 105.850 ;
        RECT 25.815 105.715 26.145 106.075 ;
        RECT 26.340 105.545 26.630 105.895 ;
        RECT 25.415 105.375 26.630 105.545 ;
        RECT 26.805 105.325 28.015 106.075 ;
        RECT 28.185 105.335 28.570 105.905 ;
        RECT 28.740 105.615 29.065 106.075 ;
        RECT 29.585 105.445 29.865 105.905 ;
        RECT 25.055 105.035 25.575 105.205 ;
        RECT 23.205 103.695 23.385 104.455 ;
        RECT 23.565 103.525 23.895 104.285 ;
        RECT 24.065 103.695 24.335 104.600 ;
        RECT 24.970 104.505 25.215 104.865 ;
        RECT 25.405 104.655 25.575 105.035 ;
        RECT 25.745 104.835 26.130 105.165 ;
        RECT 26.310 105.055 26.570 105.165 ;
        RECT 26.310 104.885 26.575 105.055 ;
        RECT 26.310 104.835 26.570 104.885 ;
        RECT 25.405 104.375 25.755 104.655 ;
        RECT 24.970 103.525 25.225 104.325 ;
        RECT 25.425 103.695 25.755 104.375 ;
        RECT 25.935 103.785 26.130 104.835 ;
        RECT 26.805 104.785 27.325 105.325 ;
        RECT 26.310 103.525 26.630 104.665 ;
        RECT 27.495 104.615 28.015 105.155 ;
        RECT 26.805 103.525 28.015 104.615 ;
        RECT 28.185 104.665 28.465 105.335 ;
        RECT 28.740 105.275 29.865 105.445 ;
        RECT 28.740 105.165 29.190 105.275 ;
        RECT 28.635 104.835 29.190 105.165 ;
        RECT 30.055 105.105 30.455 105.905 ;
        RECT 30.855 105.615 31.125 106.075 ;
        RECT 31.295 105.445 31.580 105.905 ;
        RECT 28.185 103.695 28.570 104.665 ;
        RECT 28.740 104.375 29.190 104.835 ;
        RECT 29.360 104.545 30.455 105.105 ;
        RECT 28.740 104.155 29.865 104.375 ;
        RECT 28.740 103.525 29.065 103.985 ;
        RECT 29.585 103.695 29.865 104.155 ;
        RECT 30.055 103.695 30.455 104.545 ;
        RECT 30.625 105.275 31.580 105.445 ;
        RECT 31.955 105.525 32.125 105.815 ;
        RECT 32.295 105.695 32.625 106.075 ;
        RECT 31.955 105.355 32.620 105.525 ;
        RECT 30.625 104.375 30.835 105.275 ;
        RECT 31.005 104.545 31.695 105.105 ;
        RECT 31.870 104.535 32.220 105.185 ;
        RECT 30.625 104.155 31.580 104.375 ;
        RECT 32.390 104.365 32.620 105.355 ;
        RECT 30.855 103.525 31.125 103.985 ;
        RECT 31.295 103.695 31.580 104.155 ;
        RECT 31.955 104.195 32.620 104.365 ;
        RECT 31.955 103.695 32.125 104.195 ;
        RECT 32.295 103.525 32.625 104.025 ;
        RECT 32.795 103.695 32.980 105.815 ;
        RECT 33.235 105.615 33.485 106.075 ;
        RECT 33.655 105.625 33.990 105.795 ;
        RECT 34.185 105.625 34.860 105.795 ;
        RECT 33.655 105.485 33.825 105.625 ;
        RECT 33.150 104.495 33.430 105.445 ;
        RECT 33.600 105.355 33.825 105.485 ;
        RECT 33.600 104.250 33.770 105.355 ;
        RECT 33.995 105.205 34.520 105.425 ;
        RECT 33.940 104.440 34.180 105.035 ;
        RECT 34.350 104.505 34.520 105.205 ;
        RECT 34.690 104.845 34.860 105.625 ;
        RECT 35.180 105.575 35.550 106.075 ;
        RECT 35.730 105.625 36.135 105.795 ;
        RECT 36.305 105.625 37.090 105.795 ;
        RECT 35.730 105.395 35.900 105.625 ;
        RECT 35.070 105.095 35.900 105.395 ;
        RECT 36.285 105.125 36.750 105.455 ;
        RECT 35.070 105.065 35.270 105.095 ;
        RECT 35.390 104.845 35.560 104.915 ;
        RECT 34.690 104.675 35.560 104.845 ;
        RECT 35.050 104.585 35.560 104.675 ;
        RECT 33.600 104.120 33.905 104.250 ;
        RECT 34.350 104.140 34.880 104.505 ;
        RECT 33.220 103.525 33.485 103.985 ;
        RECT 33.655 103.695 33.905 104.120 ;
        RECT 35.050 103.970 35.220 104.585 ;
        RECT 34.115 103.800 35.220 103.970 ;
        RECT 35.390 103.525 35.560 104.325 ;
        RECT 35.730 104.025 35.900 105.095 ;
        RECT 36.070 104.195 36.260 104.915 ;
        RECT 36.430 104.165 36.750 105.125 ;
        RECT 36.920 105.165 37.090 105.625 ;
        RECT 37.365 105.545 37.575 106.075 ;
        RECT 37.835 105.335 38.165 105.860 ;
        RECT 38.335 105.465 38.505 106.075 ;
        RECT 38.675 105.420 39.005 105.855 ;
        RECT 38.675 105.335 39.055 105.420 ;
        RECT 39.225 105.350 39.515 106.075 ;
        RECT 39.705 105.345 39.995 106.075 ;
        RECT 37.965 105.165 38.165 105.335 ;
        RECT 38.830 105.295 39.055 105.335 ;
        RECT 36.920 104.835 37.795 105.165 ;
        RECT 37.965 104.835 38.715 105.165 ;
        RECT 35.730 103.695 35.980 104.025 ;
        RECT 36.920 103.995 37.090 104.835 ;
        RECT 37.965 104.630 38.155 104.835 ;
        RECT 38.885 104.715 39.055 105.295 ;
        RECT 39.695 104.835 39.995 105.165 ;
        RECT 40.175 105.145 40.405 105.785 ;
        RECT 40.585 105.525 40.895 105.895 ;
        RECT 41.075 105.705 41.745 106.075 ;
        RECT 40.585 105.325 41.815 105.525 ;
        RECT 40.175 104.835 40.700 105.145 ;
        RECT 40.880 104.835 41.345 105.145 ;
        RECT 38.840 104.665 39.055 104.715 ;
        RECT 37.260 104.255 38.155 104.630 ;
        RECT 38.665 104.585 39.055 104.665 ;
        RECT 36.205 103.825 37.090 103.995 ;
        RECT 37.270 103.525 37.585 104.025 ;
        RECT 37.815 103.695 38.155 104.255 ;
        RECT 38.325 103.525 38.495 104.535 ;
        RECT 38.665 103.740 38.995 104.585 ;
        RECT 39.225 103.525 39.515 104.690 ;
        RECT 41.525 104.655 41.815 105.325 ;
        RECT 39.705 104.415 40.865 104.655 ;
        RECT 39.705 103.705 39.965 104.415 ;
        RECT 40.135 103.525 40.465 104.235 ;
        RECT 40.635 103.705 40.865 104.415 ;
        RECT 41.045 104.435 41.815 104.655 ;
        RECT 41.045 103.705 41.315 104.435 ;
        RECT 41.495 103.525 41.835 104.255 ;
        RECT 42.005 103.705 42.265 105.895 ;
        RECT 42.455 105.265 42.725 106.075 ;
        RECT 42.895 105.265 43.225 105.905 ;
        RECT 43.395 105.265 43.635 106.075 ;
        RECT 43.915 105.525 44.085 105.815 ;
        RECT 44.255 105.695 44.585 106.075 ;
        RECT 43.915 105.355 44.580 105.525 ;
        RECT 42.445 104.835 42.795 105.085 ;
        RECT 42.965 104.665 43.135 105.265 ;
        RECT 43.305 104.835 43.655 105.085 ;
        RECT 42.455 103.525 42.785 104.665 ;
        RECT 42.965 104.495 43.645 104.665 ;
        RECT 43.830 104.535 44.180 105.185 ;
        RECT 43.315 103.710 43.645 104.495 ;
        RECT 44.350 104.365 44.580 105.355 ;
        RECT 43.915 104.195 44.580 104.365 ;
        RECT 43.915 103.695 44.085 104.195 ;
        RECT 44.255 103.525 44.585 104.025 ;
        RECT 44.755 103.695 44.940 105.815 ;
        RECT 45.195 105.615 45.445 106.075 ;
        RECT 45.615 105.625 45.950 105.795 ;
        RECT 46.145 105.625 46.820 105.795 ;
        RECT 45.615 105.485 45.785 105.625 ;
        RECT 45.110 104.495 45.390 105.445 ;
        RECT 45.560 105.355 45.785 105.485 ;
        RECT 45.560 104.250 45.730 105.355 ;
        RECT 45.955 105.205 46.480 105.425 ;
        RECT 45.900 104.440 46.140 105.035 ;
        RECT 46.310 104.505 46.480 105.205 ;
        RECT 46.650 104.845 46.820 105.625 ;
        RECT 47.140 105.575 47.510 106.075 ;
        RECT 47.690 105.625 48.095 105.795 ;
        RECT 48.265 105.625 49.050 105.795 ;
        RECT 47.690 105.395 47.860 105.625 ;
        RECT 47.030 105.095 47.860 105.395 ;
        RECT 48.245 105.125 48.710 105.455 ;
        RECT 47.030 105.065 47.230 105.095 ;
        RECT 47.350 104.845 47.520 104.915 ;
        RECT 46.650 104.675 47.520 104.845 ;
        RECT 47.010 104.585 47.520 104.675 ;
        RECT 45.560 104.120 45.865 104.250 ;
        RECT 46.310 104.140 46.840 104.505 ;
        RECT 45.180 103.525 45.445 103.985 ;
        RECT 45.615 103.695 45.865 104.120 ;
        RECT 47.010 103.970 47.180 104.585 ;
        RECT 46.075 103.800 47.180 103.970 ;
        RECT 47.350 103.525 47.520 104.325 ;
        RECT 47.690 104.025 47.860 105.095 ;
        RECT 48.030 104.195 48.220 104.915 ;
        RECT 48.390 104.165 48.710 105.125 ;
        RECT 48.880 105.165 49.050 105.625 ;
        RECT 49.325 105.545 49.535 106.075 ;
        RECT 49.795 105.335 50.125 105.860 ;
        RECT 50.295 105.465 50.465 106.075 ;
        RECT 50.635 105.420 50.965 105.855 ;
        RECT 50.635 105.335 51.015 105.420 ;
        RECT 49.925 105.165 50.125 105.335 ;
        RECT 50.790 105.295 51.015 105.335 ;
        RECT 48.880 104.835 49.755 105.165 ;
        RECT 49.925 104.835 50.675 105.165 ;
        RECT 47.690 103.695 47.940 104.025 ;
        RECT 48.880 103.995 49.050 104.835 ;
        RECT 49.925 104.630 50.115 104.835 ;
        RECT 50.845 104.715 51.015 105.295 ;
        RECT 50.800 104.665 51.015 104.715 ;
        RECT 49.220 104.255 50.115 104.630 ;
        RECT 50.625 104.585 51.015 104.665 ;
        RECT 52.105 105.335 52.490 105.905 ;
        RECT 52.660 105.615 52.985 106.075 ;
        RECT 53.505 105.445 53.785 105.905 ;
        RECT 52.105 104.665 52.385 105.335 ;
        RECT 52.660 105.275 53.785 105.445 ;
        RECT 52.660 105.165 53.110 105.275 ;
        RECT 52.555 104.835 53.110 105.165 ;
        RECT 53.975 105.105 54.375 105.905 ;
        RECT 54.775 105.615 55.045 106.075 ;
        RECT 55.215 105.445 55.500 105.905 ;
        RECT 56.245 105.695 57.135 105.865 ;
        RECT 48.165 103.825 49.050 103.995 ;
        RECT 49.230 103.525 49.545 104.025 ;
        RECT 49.775 103.695 50.115 104.255 ;
        RECT 50.285 103.525 50.455 104.535 ;
        RECT 50.625 103.740 50.955 104.585 ;
        RECT 52.105 103.695 52.490 104.665 ;
        RECT 52.660 104.375 53.110 104.835 ;
        RECT 53.280 104.545 54.375 105.105 ;
        RECT 52.660 104.155 53.785 104.375 ;
        RECT 52.660 103.525 52.985 103.985 ;
        RECT 53.505 103.695 53.785 104.155 ;
        RECT 53.975 103.695 54.375 104.545 ;
        RECT 54.545 105.275 55.500 105.445 ;
        RECT 54.545 104.375 54.755 105.275 ;
        RECT 56.245 105.140 56.795 105.525 ;
        RECT 54.925 104.545 55.615 105.105 ;
        RECT 56.965 104.970 57.135 105.695 ;
        RECT 56.245 104.900 57.135 104.970 ;
        RECT 57.305 105.370 57.525 105.855 ;
        RECT 57.695 105.535 57.945 106.075 ;
        RECT 58.115 105.425 58.375 105.905 ;
        RECT 57.305 104.945 57.635 105.370 ;
        RECT 56.245 104.875 57.140 104.900 ;
        RECT 56.245 104.860 57.150 104.875 ;
        RECT 56.245 104.845 57.155 104.860 ;
        RECT 56.245 104.840 57.165 104.845 ;
        RECT 56.245 104.830 57.170 104.840 ;
        RECT 56.245 104.820 57.175 104.830 ;
        RECT 56.245 104.815 57.185 104.820 ;
        RECT 56.245 104.805 57.195 104.815 ;
        RECT 56.245 104.800 57.205 104.805 ;
        RECT 54.545 104.155 55.500 104.375 ;
        RECT 56.245 104.350 56.505 104.800 ;
        RECT 56.870 104.795 57.205 104.800 ;
        RECT 56.870 104.790 57.220 104.795 ;
        RECT 56.870 104.780 57.235 104.790 ;
        RECT 56.870 104.775 57.260 104.780 ;
        RECT 57.805 104.775 58.035 105.170 ;
        RECT 56.870 104.770 58.035 104.775 ;
        RECT 56.900 104.735 58.035 104.770 ;
        RECT 56.935 104.710 58.035 104.735 ;
        RECT 56.965 104.680 58.035 104.710 ;
        RECT 56.985 104.650 58.035 104.680 ;
        RECT 57.005 104.620 58.035 104.650 ;
        RECT 57.075 104.610 58.035 104.620 ;
        RECT 57.100 104.600 58.035 104.610 ;
        RECT 57.120 104.585 58.035 104.600 ;
        RECT 57.140 104.570 58.035 104.585 ;
        RECT 57.145 104.560 57.930 104.570 ;
        RECT 57.160 104.525 57.930 104.560 ;
        RECT 56.675 104.205 57.005 104.450 ;
        RECT 57.175 104.275 57.930 104.525 ;
        RECT 58.205 104.395 58.375 105.425 ;
        RECT 58.660 105.445 58.945 105.905 ;
        RECT 59.115 105.615 59.385 106.075 ;
        RECT 58.660 105.275 59.615 105.445 ;
        RECT 58.545 104.545 59.235 105.105 ;
        RECT 56.675 104.180 56.860 104.205 ;
        RECT 54.775 103.525 55.045 103.985 ;
        RECT 55.215 103.695 55.500 104.155 ;
        RECT 56.245 104.080 56.860 104.180 ;
        RECT 56.245 103.525 56.850 104.080 ;
        RECT 57.025 103.695 57.505 104.035 ;
        RECT 57.675 103.525 57.930 104.070 ;
        RECT 58.100 103.695 58.375 104.395 ;
        RECT 59.405 104.375 59.615 105.275 ;
        RECT 58.660 104.155 59.615 104.375 ;
        RECT 59.785 105.105 60.185 105.905 ;
        RECT 60.375 105.445 60.655 105.905 ;
        RECT 61.175 105.615 61.500 106.075 ;
        RECT 60.375 105.275 61.500 105.445 ;
        RECT 61.670 105.335 62.055 105.905 ;
        RECT 61.050 105.165 61.500 105.275 ;
        RECT 59.785 104.545 60.880 105.105 ;
        RECT 61.050 104.835 61.605 105.165 ;
        RECT 58.660 103.695 58.945 104.155 ;
        RECT 59.115 103.525 59.385 103.985 ;
        RECT 59.785 103.695 60.185 104.545 ;
        RECT 61.050 104.375 61.500 104.835 ;
        RECT 61.775 104.665 62.055 105.335 ;
        RECT 62.225 105.305 64.815 106.075 ;
        RECT 64.985 105.350 65.275 106.075 ;
        RECT 65.450 105.545 65.740 105.895 ;
        RECT 65.935 105.715 66.265 106.075 ;
        RECT 66.435 105.545 66.665 105.850 ;
        RECT 65.450 105.375 66.665 105.545 ;
        RECT 62.225 104.785 63.435 105.305 ;
        RECT 66.855 105.205 67.025 105.770 ;
        RECT 67.285 105.530 72.630 106.075 ;
        RECT 73.285 105.565 73.525 106.075 ;
        RECT 73.695 105.565 73.985 105.905 ;
        RECT 74.215 105.565 74.530 106.075 ;
        RECT 60.375 104.155 61.500 104.375 ;
        RECT 60.375 103.695 60.655 104.155 ;
        RECT 61.175 103.525 61.500 103.985 ;
        RECT 61.670 103.695 62.055 104.665 ;
        RECT 63.605 104.615 64.815 105.135 ;
        RECT 65.510 105.055 65.770 105.165 ;
        RECT 65.505 104.885 65.770 105.055 ;
        RECT 65.510 104.835 65.770 104.885 ;
        RECT 65.950 104.835 66.335 105.165 ;
        RECT 66.505 105.035 67.025 105.205 ;
        RECT 62.225 103.525 64.815 104.615 ;
        RECT 64.985 103.525 65.275 104.690 ;
        RECT 65.450 103.525 65.770 104.665 ;
        RECT 65.950 103.785 66.145 104.835 ;
        RECT 66.505 104.655 66.675 105.035 ;
        RECT 66.325 104.375 66.675 104.655 ;
        RECT 66.865 104.505 67.110 104.865 ;
        RECT 68.870 104.700 69.210 105.530 ;
        RECT 66.325 103.695 66.655 104.375 ;
        RECT 66.855 103.525 67.110 104.325 ;
        RECT 70.690 103.960 71.040 105.210 ;
        RECT 73.330 105.055 73.525 105.395 ;
        RECT 73.325 104.885 73.525 105.055 ;
        RECT 73.330 104.835 73.525 104.885 ;
        RECT 73.695 104.665 73.875 105.565 ;
        RECT 74.700 105.505 74.870 105.775 ;
        RECT 75.040 105.675 75.370 106.075 ;
        RECT 74.045 104.835 74.455 105.395 ;
        RECT 74.700 105.335 75.395 105.505 ;
        RECT 74.625 104.665 74.795 105.165 ;
        RECT 73.335 104.495 74.795 104.665 ;
        RECT 73.335 104.320 73.695 104.495 ;
        RECT 74.965 104.325 75.395 105.335 ;
        RECT 75.770 105.295 76.270 105.905 ;
        RECT 75.565 104.835 75.915 105.085 ;
        RECT 76.100 104.665 76.270 105.295 ;
        RECT 76.900 105.425 77.230 105.905 ;
        RECT 77.400 105.615 77.625 106.075 ;
        RECT 77.795 105.425 78.125 105.905 ;
        RECT 76.900 105.255 78.125 105.425 ;
        RECT 78.315 105.275 78.565 106.075 ;
        RECT 78.735 105.275 79.075 105.905 ;
        RECT 76.440 104.885 76.770 105.085 ;
        RECT 76.940 104.885 77.270 105.085 ;
        RECT 77.440 104.885 77.860 105.085 ;
        RECT 78.035 104.915 78.730 105.085 ;
        RECT 78.035 104.665 78.205 104.915 ;
        RECT 78.900 104.665 79.075 105.275 ;
        RECT 79.250 105.235 79.510 106.075 ;
        RECT 79.685 105.330 79.940 105.905 ;
        RECT 80.110 105.695 80.440 106.075 ;
        RECT 80.655 105.525 80.825 105.905 ;
        RECT 80.110 105.355 80.825 105.525 ;
        RECT 67.285 103.525 72.630 103.960 ;
        RECT 74.280 103.525 74.450 104.325 ;
        RECT 74.620 104.155 75.395 104.325 ;
        RECT 75.770 104.495 78.205 104.665 ;
        RECT 74.620 103.695 74.950 104.155 ;
        RECT 75.120 103.525 75.290 103.985 ;
        RECT 75.770 103.695 76.100 104.495 ;
        RECT 76.270 103.525 76.600 104.325 ;
        RECT 76.900 103.695 77.230 104.495 ;
        RECT 77.875 103.525 78.125 104.325 ;
        RECT 78.395 103.525 78.565 104.665 ;
        RECT 78.735 103.695 79.075 104.665 ;
        RECT 79.250 103.525 79.510 104.675 ;
        RECT 79.685 104.600 79.855 105.330 ;
        RECT 80.110 105.165 80.280 105.355 ;
        RECT 81.085 105.305 84.595 106.075 ;
        RECT 84.765 105.325 85.975 106.075 ;
        RECT 86.145 105.335 86.530 105.905 ;
        RECT 86.700 105.615 87.025 106.075 ;
        RECT 87.545 105.445 87.825 105.905 ;
        RECT 80.025 104.835 80.280 105.165 ;
        RECT 80.110 104.625 80.280 104.835 ;
        RECT 80.560 104.805 80.915 105.175 ;
        RECT 81.085 104.785 82.735 105.305 ;
        RECT 79.685 103.695 79.940 104.600 ;
        RECT 80.110 104.455 80.825 104.625 ;
        RECT 82.905 104.615 84.595 105.135 ;
        RECT 84.765 104.785 85.285 105.325 ;
        RECT 85.455 104.615 85.975 105.155 ;
        RECT 80.110 103.525 80.440 104.285 ;
        RECT 80.655 103.695 80.825 104.455 ;
        RECT 81.085 103.525 84.595 104.615 ;
        RECT 84.765 103.525 85.975 104.615 ;
        RECT 86.145 104.665 86.425 105.335 ;
        RECT 86.700 105.275 87.825 105.445 ;
        RECT 86.700 105.165 87.150 105.275 ;
        RECT 86.595 104.835 87.150 105.165 ;
        RECT 88.015 105.105 88.415 105.905 ;
        RECT 88.815 105.615 89.085 106.075 ;
        RECT 89.255 105.445 89.540 105.905 ;
        RECT 86.145 103.695 86.530 104.665 ;
        RECT 86.700 104.375 87.150 104.835 ;
        RECT 87.320 104.545 88.415 105.105 ;
        RECT 86.700 104.155 87.825 104.375 ;
        RECT 86.700 103.525 87.025 103.985 ;
        RECT 87.545 103.695 87.825 104.155 ;
        RECT 88.015 103.695 88.415 104.545 ;
        RECT 88.585 105.275 89.540 105.445 ;
        RECT 90.745 105.325 91.955 106.075 ;
        RECT 100.080 105.490 102.000 106.760 ;
        RECT 103.510 106.750 104.070 106.760 ;
        RECT 103.740 105.660 104.070 106.750 ;
        RECT 104.440 106.280 105.480 106.450 ;
        RECT 104.440 105.840 105.480 106.010 ;
        RECT 105.650 105.980 105.820 106.310 ;
        RECT 88.585 104.375 88.795 105.275 ;
        RECT 88.965 104.545 89.655 105.105 ;
        RECT 90.745 104.615 91.265 105.155 ;
        RECT 91.435 104.785 91.955 105.325 ;
        RECT 103.900 105.440 104.070 105.660 ;
        RECT 106.160 105.440 106.330 106.850 ;
        RECT 103.900 105.270 106.330 105.440 ;
        RECT 107.910 107.360 118.540 107.530 ;
        RECT 120.020 116.640 126.250 116.800 ;
        RECT 120.020 114.380 120.690 116.640 ;
        RECT 121.360 116.070 125.400 116.240 ;
        RECT 121.020 115.010 121.190 116.010 ;
        RECT 125.570 115.010 125.740 116.010 ;
        RECT 121.360 114.780 125.400 114.950 ;
        RECT 126.080 114.380 126.250 116.640 ;
        RECT 120.020 114.210 126.250 114.380 ;
        RECT 120.020 110.950 120.690 114.210 ;
        RECT 121.360 113.640 125.400 113.810 ;
        RECT 121.020 111.580 121.190 113.580 ;
        RECT 125.570 111.580 125.740 113.580 ;
        RECT 121.360 111.350 125.400 111.520 ;
        RECT 126.080 110.950 126.250 114.210 ;
        RECT 120.020 110.780 126.250 110.950 ;
        RECT 120.020 107.520 120.690 110.780 ;
        RECT 121.360 110.210 125.400 110.380 ;
        RECT 121.020 108.150 121.190 110.150 ;
        RECT 125.570 108.150 125.740 110.150 ;
        RECT 121.360 107.920 125.400 108.090 ;
        RECT 126.080 107.520 126.250 110.780 ;
        RECT 120.020 107.510 126.250 107.520 ;
        RECT 127.840 116.780 137.670 116.820 ;
        RECT 140.540 116.800 146.280 116.810 ;
        RECT 127.840 116.650 138.470 116.780 ;
        RECT 127.840 114.390 128.010 116.650 ;
        RECT 128.735 116.080 136.775 116.250 ;
        RECT 128.350 115.020 128.520 116.020 ;
        RECT 136.990 115.020 137.160 116.020 ;
        RECT 128.735 114.790 136.775 114.960 ;
        RECT 137.500 114.390 138.470 116.650 ;
        RECT 127.840 114.220 138.470 114.390 ;
        RECT 127.840 110.960 128.010 114.220 ;
        RECT 128.735 113.650 136.775 113.820 ;
        RECT 128.350 111.590 128.520 113.590 ;
        RECT 136.990 111.590 137.160 113.590 ;
        RECT 128.735 111.360 136.775 111.530 ;
        RECT 137.500 110.960 138.470 114.220 ;
        RECT 127.840 110.790 138.470 110.960 ;
        RECT 127.840 107.530 128.010 110.790 ;
        RECT 128.735 110.220 136.775 110.390 ;
        RECT 128.350 108.160 128.520 110.160 ;
        RECT 136.990 108.160 137.160 110.160 ;
        RECT 128.735 107.930 136.775 108.100 ;
        RECT 137.500 107.530 138.470 110.790 ;
        RECT 120.020 107.410 126.260 107.510 ;
        RECT 107.910 105.100 108.080 107.360 ;
        RECT 108.805 106.790 116.845 106.960 ;
        RECT 108.420 105.730 108.590 106.730 ;
        RECT 117.060 105.730 117.230 106.730 ;
        RECT 108.805 105.500 116.845 105.670 ;
        RECT 117.570 105.100 118.540 107.360 ;
        RECT 120.010 106.850 126.260 107.410 ;
        RECT 120.010 106.830 125.180 106.850 ;
        RECT 120.010 106.760 124.000 106.830 ;
        RECT 120.010 106.250 121.930 106.760 ;
        RECT 123.440 106.750 124.000 106.760 ;
        RECT 107.910 105.070 118.540 105.100 ;
        RECT 107.880 104.960 118.540 105.070 ;
        RECT 106.130 104.910 118.540 104.960 ;
        RECT 101.790 104.740 118.540 104.910 ;
        RECT 88.585 104.155 89.540 104.375 ;
        RECT 88.815 103.525 89.085 103.985 ;
        RECT 89.255 103.695 89.540 104.155 ;
        RECT 90.745 103.525 91.955 104.615 ;
        RECT 13.380 103.355 92.040 103.525 ;
        RECT 13.465 102.265 14.675 103.355 ;
        RECT 13.465 101.555 13.985 102.095 ;
        RECT 14.155 101.725 14.675 102.265 ;
        RECT 14.845 102.385 15.115 103.155 ;
        RECT 15.285 102.575 15.615 103.355 ;
        RECT 15.820 102.750 16.005 103.155 ;
        RECT 16.175 102.930 16.510 103.355 ;
        RECT 15.820 102.575 16.485 102.750 ;
        RECT 14.845 102.215 15.975 102.385 ;
        RECT 13.465 100.805 14.675 101.555 ;
        RECT 14.845 101.305 15.015 102.215 ;
        RECT 15.185 101.465 15.545 102.045 ;
        RECT 15.725 101.715 15.975 102.215 ;
        RECT 16.145 101.545 16.485 102.575 ;
        RECT 17.605 102.215 17.885 103.355 ;
        RECT 18.055 102.205 18.385 103.185 ;
        RECT 18.555 102.215 18.815 103.355 ;
        RECT 19.100 102.725 19.385 103.185 ;
        RECT 19.555 102.895 19.825 103.355 ;
        RECT 19.100 102.505 20.055 102.725 ;
        RECT 17.615 101.775 17.950 102.045 ;
        RECT 18.120 101.605 18.290 102.205 ;
        RECT 18.460 101.795 18.795 102.045 ;
        RECT 18.985 101.775 19.675 102.335 ;
        RECT 19.845 101.605 20.055 102.505 ;
        RECT 15.800 101.375 16.485 101.545 ;
        RECT 14.845 100.975 15.105 101.305 ;
        RECT 15.315 100.805 15.590 101.285 ;
        RECT 15.800 100.975 16.005 101.375 ;
        RECT 16.175 100.805 16.510 101.205 ;
        RECT 17.605 100.805 17.915 101.605 ;
        RECT 18.120 100.975 18.815 101.605 ;
        RECT 19.100 101.435 20.055 101.605 ;
        RECT 20.225 102.335 20.625 103.185 ;
        RECT 20.815 102.725 21.095 103.185 ;
        RECT 21.615 102.895 21.940 103.355 ;
        RECT 20.815 102.505 21.940 102.725 ;
        RECT 20.225 101.775 21.320 102.335 ;
        RECT 21.490 102.045 21.940 102.505 ;
        RECT 22.110 102.215 22.495 103.185 ;
        RECT 23.125 102.845 23.425 103.355 ;
        RECT 23.595 102.675 23.925 103.185 ;
        RECT 24.095 102.845 24.725 103.355 ;
        RECT 25.305 102.845 25.685 103.015 ;
        RECT 25.855 102.845 26.155 103.355 ;
        RECT 25.515 102.675 25.685 102.845 ;
        RECT 19.100 100.975 19.385 101.435 ;
        RECT 19.555 100.805 19.825 101.265 ;
        RECT 20.225 100.975 20.625 101.775 ;
        RECT 21.490 101.715 22.045 102.045 ;
        RECT 21.490 101.605 21.940 101.715 ;
        RECT 20.815 101.435 21.940 101.605 ;
        RECT 22.215 101.545 22.495 102.215 ;
        RECT 20.815 100.975 21.095 101.435 ;
        RECT 21.615 100.805 21.940 101.265 ;
        RECT 22.110 100.975 22.495 101.545 ;
        RECT 23.125 102.505 25.345 102.675 ;
        RECT 23.125 101.545 23.295 102.505 ;
        RECT 23.465 102.165 25.005 102.335 ;
        RECT 23.465 101.715 23.710 102.165 ;
        RECT 23.970 101.795 24.665 101.995 ;
        RECT 24.835 101.965 25.005 102.165 ;
        RECT 25.175 102.305 25.345 102.505 ;
        RECT 25.515 102.475 26.175 102.675 ;
        RECT 25.175 102.135 25.835 102.305 ;
        RECT 24.835 101.795 25.435 101.965 ;
        RECT 25.665 101.715 25.835 102.135 ;
        RECT 23.125 101.000 23.590 101.545 ;
        RECT 24.095 100.805 24.265 101.625 ;
        RECT 24.435 101.545 25.345 101.625 ;
        RECT 26.005 101.545 26.175 102.475 ;
        RECT 26.345 102.190 26.635 103.355 ;
        RECT 26.895 102.685 27.065 103.185 ;
        RECT 27.235 102.855 27.565 103.355 ;
        RECT 26.895 102.515 27.560 102.685 ;
        RECT 26.810 101.695 27.160 102.345 ;
        RECT 24.435 101.455 25.685 101.545 ;
        RECT 24.435 100.975 24.765 101.455 ;
        RECT 25.175 101.375 25.685 101.455 ;
        RECT 24.935 100.805 25.285 101.195 ;
        RECT 25.455 100.975 25.685 101.375 ;
        RECT 25.855 101.065 26.175 101.545 ;
        RECT 26.345 100.805 26.635 101.530 ;
        RECT 27.330 101.525 27.560 102.515 ;
        RECT 26.895 101.355 27.560 101.525 ;
        RECT 26.895 101.065 27.065 101.355 ;
        RECT 27.235 100.805 27.565 101.185 ;
        RECT 27.735 101.065 27.920 103.185 ;
        RECT 28.160 102.895 28.425 103.355 ;
        RECT 28.595 102.760 28.845 103.185 ;
        RECT 29.055 102.910 30.160 103.080 ;
        RECT 28.540 102.630 28.845 102.760 ;
        RECT 28.090 101.435 28.370 102.385 ;
        RECT 28.540 101.525 28.710 102.630 ;
        RECT 28.880 101.845 29.120 102.440 ;
        RECT 29.290 102.375 29.820 102.740 ;
        RECT 29.290 101.675 29.460 102.375 ;
        RECT 29.990 102.295 30.160 102.910 ;
        RECT 30.330 102.555 30.500 103.355 ;
        RECT 30.670 102.855 30.920 103.185 ;
        RECT 31.145 102.885 32.030 103.055 ;
        RECT 29.990 102.205 30.500 102.295 ;
        RECT 28.540 101.395 28.765 101.525 ;
        RECT 28.935 101.455 29.460 101.675 ;
        RECT 29.630 102.035 30.500 102.205 ;
        RECT 28.175 100.805 28.425 101.265 ;
        RECT 28.595 101.255 28.765 101.395 ;
        RECT 29.630 101.255 29.800 102.035 ;
        RECT 30.330 101.965 30.500 102.035 ;
        RECT 30.010 101.785 30.210 101.815 ;
        RECT 30.670 101.785 30.840 102.855 ;
        RECT 31.010 101.965 31.200 102.685 ;
        RECT 30.010 101.485 30.840 101.785 ;
        RECT 31.370 101.755 31.690 102.715 ;
        RECT 28.595 101.085 28.930 101.255 ;
        RECT 29.125 101.085 29.800 101.255 ;
        RECT 30.120 100.805 30.490 101.305 ;
        RECT 30.670 101.255 30.840 101.485 ;
        RECT 31.225 101.425 31.690 101.755 ;
        RECT 31.860 102.045 32.030 102.885 ;
        RECT 32.210 102.855 32.525 103.355 ;
        RECT 32.755 102.625 33.095 103.185 ;
        RECT 32.200 102.250 33.095 102.625 ;
        RECT 33.265 102.345 33.435 103.355 ;
        RECT 32.905 102.045 33.095 102.250 ;
        RECT 33.605 102.295 33.935 103.140 ;
        RECT 33.605 102.215 33.995 102.295 ;
        RECT 34.165 102.265 37.675 103.355 ;
        RECT 33.780 102.165 33.995 102.215 ;
        RECT 31.860 101.715 32.735 102.045 ;
        RECT 32.905 101.715 33.655 102.045 ;
        RECT 31.860 101.255 32.030 101.715 ;
        RECT 32.905 101.545 33.105 101.715 ;
        RECT 33.825 101.585 33.995 102.165 ;
        RECT 33.770 101.545 33.995 101.585 ;
        RECT 30.670 101.085 31.075 101.255 ;
        RECT 31.245 101.085 32.030 101.255 ;
        RECT 32.305 100.805 32.515 101.335 ;
        RECT 32.775 101.020 33.105 101.545 ;
        RECT 33.615 101.460 33.995 101.545 ;
        RECT 34.165 101.575 35.815 102.095 ;
        RECT 35.985 101.745 37.675 102.265 ;
        RECT 38.305 102.215 38.565 103.355 ;
        RECT 38.735 102.205 39.065 103.185 ;
        RECT 39.235 102.215 39.515 103.355 ;
        RECT 40.150 102.405 40.415 103.175 ;
        RECT 40.585 102.635 40.915 103.355 ;
        RECT 41.105 102.815 41.365 103.175 ;
        RECT 41.535 102.985 41.865 103.355 ;
        RECT 42.035 102.815 42.295 103.175 ;
        RECT 41.105 102.585 42.295 102.815 ;
        RECT 42.865 102.405 43.155 103.175 ;
        RECT 38.325 101.795 38.660 102.045 ;
        RECT 38.830 101.605 39.000 102.205 ;
        RECT 39.170 101.775 39.505 102.045 ;
        RECT 33.275 100.805 33.445 101.415 ;
        RECT 33.615 101.025 33.945 101.460 ;
        RECT 34.165 100.805 37.675 101.575 ;
        RECT 38.305 100.975 39.000 101.605 ;
        RECT 39.205 100.805 39.515 101.605 ;
        RECT 40.150 100.985 40.485 102.405 ;
        RECT 40.660 102.225 43.155 102.405 ;
        RECT 40.660 101.535 40.885 102.225 ;
        RECT 43.365 102.215 43.655 103.355 ;
        RECT 44.450 103.015 45.815 103.185 ;
        RECT 44.450 102.805 44.780 103.015 ;
        RECT 43.825 102.555 44.780 102.805 ;
        RECT 41.085 101.715 41.365 102.045 ;
        RECT 41.545 101.715 42.120 102.045 ;
        RECT 42.300 101.715 42.735 102.045 ;
        RECT 42.915 101.715 43.185 102.045 ;
        RECT 43.365 101.715 43.640 102.045 ;
        RECT 43.825 101.545 43.995 102.555 ;
        RECT 44.165 101.715 44.520 102.380 ;
        RECT 44.705 101.715 44.980 102.380 ;
        RECT 45.150 102.045 45.475 102.845 ;
        RECT 45.645 102.385 45.815 103.015 ;
        RECT 45.985 102.555 46.275 103.355 ;
        RECT 45.645 102.215 46.320 102.385 ;
        RECT 46.490 102.215 46.875 103.175 ;
        RECT 47.045 102.265 50.555 103.355 ;
        RECT 46.150 102.045 46.320 102.215 ;
        RECT 45.150 101.715 45.495 102.045 ;
        RECT 45.705 101.795 45.955 102.045 ;
        RECT 46.150 101.795 46.515 102.045 ;
        RECT 45.785 101.715 45.955 101.795 ;
        RECT 46.325 101.715 46.515 101.795 ;
        RECT 46.700 101.545 46.875 102.215 ;
        RECT 40.660 101.345 43.145 101.535 ;
        RECT 40.665 100.805 41.410 101.175 ;
        RECT 41.975 100.985 42.230 101.345 ;
        RECT 42.410 100.805 42.740 101.175 ;
        RECT 42.920 100.985 43.145 101.345 ;
        RECT 43.365 101.185 43.655 101.455 ;
        RECT 43.825 101.355 44.250 101.545 ;
        RECT 44.420 101.375 45.820 101.545 ;
        RECT 44.420 101.185 44.750 101.375 ;
        RECT 43.365 100.975 44.750 101.185 ;
        RECT 44.985 100.805 45.315 101.205 ;
        RECT 45.490 100.975 45.820 101.375 ;
        RECT 46.025 100.805 46.195 101.365 ;
        RECT 46.365 100.975 46.875 101.545 ;
        RECT 47.045 101.575 48.695 102.095 ;
        RECT 48.865 101.745 50.555 102.265 ;
        RECT 50.785 102.215 50.995 103.355 ;
        RECT 51.165 102.205 51.495 103.185 ;
        RECT 51.665 102.215 51.895 103.355 ;
        RECT 47.045 100.805 50.555 101.575 ;
        RECT 50.785 100.805 50.995 101.625 ;
        RECT 51.165 101.605 51.415 102.205 ;
        RECT 52.105 102.190 52.395 103.355 ;
        RECT 53.545 102.295 53.875 103.140 ;
        RECT 54.045 102.345 54.215 103.355 ;
        RECT 54.385 102.625 54.725 103.185 ;
        RECT 54.955 102.855 55.270 103.355 ;
        RECT 55.450 102.885 56.335 103.055 ;
        RECT 53.485 102.215 53.875 102.295 ;
        RECT 54.385 102.250 55.280 102.625 ;
        RECT 53.485 102.165 53.700 102.215 ;
        RECT 51.585 101.795 51.915 102.045 ;
        RECT 51.165 100.975 51.495 101.605 ;
        RECT 51.665 100.805 51.895 101.625 ;
        RECT 53.485 101.585 53.655 102.165 ;
        RECT 54.385 102.045 54.575 102.250 ;
        RECT 55.450 102.045 55.620 102.885 ;
        RECT 56.560 102.855 56.810 103.185 ;
        RECT 53.825 101.715 54.575 102.045 ;
        RECT 54.745 101.715 55.620 102.045 ;
        RECT 53.485 101.545 53.710 101.585 ;
        RECT 54.375 101.545 54.575 101.715 ;
        RECT 52.105 100.805 52.395 101.530 ;
        RECT 53.485 101.460 53.865 101.545 ;
        RECT 53.535 101.025 53.865 101.460 ;
        RECT 54.035 100.805 54.205 101.415 ;
        RECT 54.375 101.020 54.705 101.545 ;
        RECT 54.965 100.805 55.175 101.335 ;
        RECT 55.450 101.255 55.620 101.715 ;
        RECT 55.790 101.755 56.110 102.715 ;
        RECT 56.280 101.965 56.470 102.685 ;
        RECT 56.640 101.785 56.810 102.855 ;
        RECT 56.980 102.555 57.150 103.355 ;
        RECT 57.320 102.910 58.425 103.080 ;
        RECT 57.320 102.295 57.490 102.910 ;
        RECT 58.635 102.760 58.885 103.185 ;
        RECT 59.055 102.895 59.320 103.355 ;
        RECT 57.660 102.375 58.190 102.740 ;
        RECT 58.635 102.630 58.940 102.760 ;
        RECT 56.980 102.205 57.490 102.295 ;
        RECT 56.980 102.035 57.850 102.205 ;
        RECT 56.980 101.965 57.150 102.035 ;
        RECT 57.270 101.785 57.470 101.815 ;
        RECT 55.790 101.425 56.255 101.755 ;
        RECT 56.640 101.485 57.470 101.785 ;
        RECT 56.640 101.255 56.810 101.485 ;
        RECT 55.450 101.085 56.235 101.255 ;
        RECT 56.405 101.085 56.810 101.255 ;
        RECT 56.990 100.805 57.360 101.305 ;
        RECT 57.680 101.255 57.850 102.035 ;
        RECT 58.020 101.675 58.190 102.375 ;
        RECT 58.360 101.845 58.600 102.440 ;
        RECT 58.020 101.455 58.545 101.675 ;
        RECT 58.770 101.525 58.940 102.630 ;
        RECT 58.715 101.395 58.940 101.525 ;
        RECT 59.110 101.435 59.390 102.385 ;
        RECT 58.715 101.255 58.885 101.395 ;
        RECT 57.680 101.085 58.355 101.255 ;
        RECT 58.550 101.085 58.885 101.255 ;
        RECT 59.055 100.805 59.305 101.265 ;
        RECT 59.560 101.065 59.745 103.185 ;
        RECT 59.915 102.855 60.245 103.355 ;
        RECT 60.415 102.685 60.585 103.185 ;
        RECT 59.920 102.515 60.585 102.685 ;
        RECT 59.920 101.525 60.150 102.515 ;
        RECT 60.320 101.695 60.670 102.345 ;
        RECT 60.850 102.215 61.185 103.185 ;
        RECT 61.355 102.215 61.525 103.355 ;
        RECT 61.695 103.015 63.725 103.185 ;
        RECT 60.850 101.545 61.020 102.215 ;
        RECT 61.695 102.045 61.865 103.015 ;
        RECT 61.190 101.715 61.445 102.045 ;
        RECT 61.670 101.715 61.865 102.045 ;
        RECT 62.035 102.675 63.160 102.845 ;
        RECT 61.275 101.545 61.445 101.715 ;
        RECT 62.035 101.545 62.205 102.675 ;
        RECT 59.920 101.355 60.585 101.525 ;
        RECT 59.915 100.805 60.245 101.185 ;
        RECT 60.415 101.065 60.585 101.355 ;
        RECT 60.850 100.975 61.105 101.545 ;
        RECT 61.275 101.375 62.205 101.545 ;
        RECT 62.375 102.335 63.385 102.505 ;
        RECT 62.375 101.535 62.545 102.335 ;
        RECT 62.750 101.655 63.025 102.135 ;
        RECT 62.745 101.485 63.025 101.655 ;
        RECT 62.030 101.340 62.205 101.375 ;
        RECT 61.275 100.805 61.605 101.205 ;
        RECT 62.030 100.975 62.560 101.340 ;
        RECT 62.750 100.975 63.025 101.485 ;
        RECT 63.195 100.975 63.385 102.335 ;
        RECT 63.555 102.350 63.725 103.015 ;
        RECT 63.895 102.595 64.065 103.355 ;
        RECT 64.300 102.595 64.815 103.005 ;
        RECT 63.555 102.160 64.305 102.350 ;
        RECT 64.475 101.785 64.815 102.595 ;
        RECT 65.075 102.425 65.245 103.185 ;
        RECT 65.460 102.595 65.790 103.355 ;
        RECT 65.075 102.255 65.790 102.425 ;
        RECT 65.960 102.280 66.215 103.185 ;
        RECT 63.585 101.615 64.815 101.785 ;
        RECT 64.985 101.705 65.340 102.075 ;
        RECT 65.620 102.045 65.790 102.255 ;
        RECT 65.620 101.715 65.875 102.045 ;
        RECT 63.565 100.805 64.075 101.340 ;
        RECT 64.295 101.010 64.540 101.615 ;
        RECT 65.620 101.525 65.790 101.715 ;
        RECT 66.045 101.550 66.215 102.280 ;
        RECT 66.390 102.205 66.650 103.355 ;
        RECT 66.835 102.385 67.165 103.170 ;
        RECT 66.835 102.215 67.515 102.385 ;
        RECT 67.695 102.215 68.025 103.355 ;
        RECT 68.205 102.265 71.715 103.355 ;
        RECT 66.825 101.795 67.175 102.045 ;
        RECT 65.075 101.355 65.790 101.525 ;
        RECT 65.075 100.975 65.245 101.355 ;
        RECT 65.460 100.805 65.790 101.185 ;
        RECT 65.960 100.975 66.215 101.550 ;
        RECT 66.390 100.805 66.650 101.645 ;
        RECT 67.345 101.615 67.515 102.215 ;
        RECT 67.685 101.795 68.035 102.045 ;
        RECT 66.845 100.805 67.085 101.615 ;
        RECT 67.255 100.975 67.585 101.615 ;
        RECT 67.755 100.805 68.025 101.615 ;
        RECT 68.205 101.575 69.855 102.095 ;
        RECT 70.025 101.745 71.715 102.265 ;
        RECT 72.805 102.215 73.065 103.355 ;
        RECT 73.235 102.205 73.565 103.185 ;
        RECT 73.735 102.215 74.015 103.355 ;
        RECT 73.325 102.165 73.500 102.205 ;
        RECT 74.185 102.175 74.505 103.355 ;
        RECT 74.675 102.335 74.875 103.125 ;
        RECT 75.200 102.525 75.585 103.185 ;
        RECT 75.980 102.595 76.765 103.355 ;
        RECT 75.175 102.425 75.585 102.525 ;
        RECT 74.675 102.165 75.005 102.335 ;
        RECT 75.175 102.215 76.785 102.425 ;
        RECT 72.825 101.795 73.160 102.045 ;
        RECT 73.330 101.605 73.500 102.165 ;
        RECT 74.825 102.045 75.005 102.165 ;
        RECT 73.670 101.775 74.005 102.045 ;
        RECT 74.185 101.795 74.650 101.995 ;
        RECT 74.825 101.795 75.155 102.045 ;
        RECT 75.325 101.995 75.790 102.045 ;
        RECT 75.325 101.825 75.795 101.995 ;
        RECT 75.325 101.795 75.790 101.825 ;
        RECT 75.985 101.795 76.340 102.045 ;
        RECT 76.510 101.615 76.785 102.215 ;
        RECT 68.205 100.805 71.715 101.575 ;
        RECT 72.805 100.975 73.500 101.605 ;
        RECT 73.705 100.805 74.015 101.605 ;
        RECT 74.185 101.415 75.365 101.585 ;
        RECT 74.185 101.000 74.525 101.415 ;
        RECT 74.695 100.805 74.865 101.245 ;
        RECT 75.035 101.195 75.365 101.415 ;
        RECT 75.535 101.435 76.785 101.615 ;
        RECT 75.535 101.365 75.900 101.435 ;
        RECT 75.035 101.015 76.285 101.195 ;
        RECT 76.555 100.805 76.725 101.265 ;
        RECT 76.955 101.085 77.235 103.185 ;
        RECT 77.865 102.190 78.155 103.355 ;
        RECT 78.325 102.265 79.995 103.355 ;
        RECT 80.715 102.685 80.885 103.185 ;
        RECT 81.055 102.855 81.385 103.355 ;
        RECT 80.715 102.515 81.380 102.685 ;
        RECT 78.325 101.575 79.075 102.095 ;
        RECT 79.245 101.745 79.995 102.265 ;
        RECT 80.630 101.695 80.980 102.345 ;
        RECT 77.865 100.805 78.155 101.530 ;
        RECT 78.325 100.805 79.995 101.575 ;
        RECT 81.150 101.525 81.380 102.515 ;
        RECT 80.715 101.355 81.380 101.525 ;
        RECT 80.715 101.065 80.885 101.355 ;
        RECT 81.055 100.805 81.385 101.185 ;
        RECT 81.555 101.065 81.740 103.185 ;
        RECT 81.980 102.895 82.245 103.355 ;
        RECT 82.415 102.760 82.665 103.185 ;
        RECT 82.875 102.910 83.980 103.080 ;
        RECT 82.360 102.630 82.665 102.760 ;
        RECT 81.910 101.435 82.190 102.385 ;
        RECT 82.360 101.525 82.530 102.630 ;
        RECT 82.700 101.845 82.940 102.440 ;
        RECT 83.110 102.375 83.640 102.740 ;
        RECT 83.110 101.675 83.280 102.375 ;
        RECT 83.810 102.295 83.980 102.910 ;
        RECT 84.150 102.555 84.320 103.355 ;
        RECT 84.490 102.855 84.740 103.185 ;
        RECT 84.965 102.885 85.850 103.055 ;
        RECT 83.810 102.205 84.320 102.295 ;
        RECT 82.360 101.395 82.585 101.525 ;
        RECT 82.755 101.455 83.280 101.675 ;
        RECT 83.450 102.035 84.320 102.205 ;
        RECT 81.995 100.805 82.245 101.265 ;
        RECT 82.415 101.255 82.585 101.395 ;
        RECT 83.450 101.255 83.620 102.035 ;
        RECT 84.150 101.965 84.320 102.035 ;
        RECT 83.830 101.785 84.030 101.815 ;
        RECT 84.490 101.785 84.660 102.855 ;
        RECT 84.830 101.965 85.020 102.685 ;
        RECT 83.830 101.485 84.660 101.785 ;
        RECT 85.190 101.755 85.510 102.715 ;
        RECT 82.415 101.085 82.750 101.255 ;
        RECT 82.945 101.085 83.620 101.255 ;
        RECT 83.940 100.805 84.310 101.305 ;
        RECT 84.490 101.255 84.660 101.485 ;
        RECT 85.045 101.425 85.510 101.755 ;
        RECT 85.680 102.045 85.850 102.885 ;
        RECT 86.030 102.855 86.345 103.355 ;
        RECT 86.575 102.625 86.915 103.185 ;
        RECT 86.020 102.250 86.915 102.625 ;
        RECT 87.085 102.345 87.255 103.355 ;
        RECT 86.725 102.045 86.915 102.250 ;
        RECT 87.425 102.295 87.755 103.140 ;
        RECT 87.425 102.215 87.815 102.295 ;
        RECT 87.985 102.265 90.575 103.355 ;
        RECT 87.600 102.165 87.815 102.215 ;
        RECT 85.680 101.715 86.555 102.045 ;
        RECT 86.725 101.715 87.475 102.045 ;
        RECT 85.680 101.255 85.850 101.715 ;
        RECT 86.725 101.545 86.925 101.715 ;
        RECT 87.645 101.585 87.815 102.165 ;
        RECT 87.590 101.545 87.815 101.585 ;
        RECT 84.490 101.085 84.895 101.255 ;
        RECT 85.065 101.085 85.850 101.255 ;
        RECT 86.125 100.805 86.335 101.335 ;
        RECT 86.595 101.020 86.925 101.545 ;
        RECT 87.435 101.460 87.815 101.545 ;
        RECT 87.985 101.575 89.195 102.095 ;
        RECT 89.365 101.745 90.575 102.265 ;
        RECT 90.745 102.265 91.955 103.355 ;
        RECT 101.790 103.330 101.960 104.740 ;
        RECT 102.330 104.170 105.370 104.340 ;
        RECT 102.330 103.730 105.370 103.900 ;
        RECT 105.585 103.870 105.755 104.200 ;
        RECT 106.090 103.980 118.540 104.740 ;
        RECT 120.000 105.490 121.930 106.250 ;
        RECT 123.670 105.660 124.000 106.750 ;
        RECT 124.370 106.280 125.410 106.450 ;
        RECT 124.370 105.840 125.410 106.010 ;
        RECT 125.580 105.980 125.750 106.310 ;
        RECT 106.090 103.970 118.430 103.980 ;
        RECT 106.090 103.960 111.970 103.970 ;
        RECT 106.090 103.940 106.660 103.960 ;
        RECT 107.880 103.950 111.970 103.960 ;
        RECT 106.100 103.330 106.270 103.940 ;
        RECT 101.790 103.160 106.270 103.330 ;
        RECT 120.000 102.740 120.960 105.490 ;
        RECT 123.830 105.440 124.000 105.660 ;
        RECT 126.090 105.440 126.260 106.850 ;
        RECT 123.830 105.270 126.260 105.440 ;
        RECT 127.840 107.360 138.470 107.530 ;
        RECT 140.050 116.640 146.280 116.800 ;
        RECT 140.050 114.380 140.720 116.640 ;
        RECT 141.390 116.070 145.430 116.240 ;
        RECT 141.050 115.010 141.220 116.010 ;
        RECT 145.600 115.010 145.770 116.010 ;
        RECT 141.390 114.780 145.430 114.950 ;
        RECT 146.110 114.380 146.280 116.640 ;
        RECT 140.050 114.210 146.280 114.380 ;
        RECT 140.050 110.950 140.720 114.210 ;
        RECT 141.390 113.640 145.430 113.810 ;
        RECT 141.050 111.580 141.220 113.580 ;
        RECT 145.600 111.580 145.770 113.580 ;
        RECT 141.390 111.350 145.430 111.520 ;
        RECT 146.110 110.950 146.280 114.210 ;
        RECT 140.050 110.780 146.280 110.950 ;
        RECT 140.050 107.520 140.720 110.780 ;
        RECT 141.390 110.210 145.430 110.380 ;
        RECT 141.050 108.150 141.220 110.150 ;
        RECT 145.600 108.150 145.770 110.150 ;
        RECT 141.390 107.920 145.430 108.090 ;
        RECT 146.110 107.520 146.280 110.780 ;
        RECT 140.050 107.510 146.280 107.520 ;
        RECT 147.870 116.780 157.700 116.820 ;
        RECT 147.870 116.650 158.500 116.780 ;
        RECT 147.870 114.390 148.040 116.650 ;
        RECT 148.765 116.080 156.805 116.250 ;
        RECT 148.380 115.020 148.550 116.020 ;
        RECT 157.020 115.020 157.190 116.020 ;
        RECT 148.765 114.790 156.805 114.960 ;
        RECT 157.530 114.390 158.500 116.650 ;
        RECT 147.870 114.220 158.500 114.390 ;
        RECT 147.870 110.960 148.040 114.220 ;
        RECT 148.765 113.650 156.805 113.820 ;
        RECT 148.380 111.590 148.550 113.590 ;
        RECT 157.020 111.590 157.190 113.590 ;
        RECT 148.765 111.360 156.805 111.530 ;
        RECT 157.530 110.960 158.500 114.220 ;
        RECT 147.870 110.790 158.500 110.960 ;
        RECT 147.870 107.530 148.040 110.790 ;
        RECT 148.765 110.220 156.805 110.390 ;
        RECT 148.380 108.160 148.550 110.160 ;
        RECT 157.020 108.160 157.190 110.160 ;
        RECT 148.765 107.930 156.805 108.100 ;
        RECT 157.530 107.530 158.500 110.790 ;
        RECT 140.050 107.410 146.290 107.510 ;
        RECT 127.840 105.100 128.010 107.360 ;
        RECT 128.735 106.790 136.775 106.960 ;
        RECT 128.350 105.730 128.520 106.730 ;
        RECT 136.990 105.730 137.160 106.730 ;
        RECT 128.735 105.500 136.775 105.670 ;
        RECT 137.500 105.100 138.470 107.360 ;
        RECT 140.040 106.850 146.290 107.410 ;
        RECT 140.040 106.830 145.210 106.850 ;
        RECT 140.040 106.760 144.030 106.830 ;
        RECT 140.040 105.490 141.960 106.760 ;
        RECT 143.470 106.750 144.030 106.760 ;
        RECT 143.700 105.660 144.030 106.750 ;
        RECT 144.400 106.280 145.440 106.450 ;
        RECT 144.400 105.840 145.440 106.010 ;
        RECT 145.610 105.980 145.780 106.310 ;
        RECT 143.860 105.440 144.030 105.660 ;
        RECT 146.120 105.440 146.290 106.850 ;
        RECT 143.860 105.270 146.290 105.440 ;
        RECT 147.870 107.360 158.500 107.530 ;
        RECT 127.840 105.070 138.470 105.100 ;
        RECT 147.870 105.100 148.040 107.360 ;
        RECT 148.765 106.790 156.805 106.960 ;
        RECT 148.380 105.730 148.550 106.730 ;
        RECT 157.020 105.730 157.190 106.730 ;
        RECT 148.765 105.500 156.805 105.670 ;
        RECT 157.530 105.100 158.500 107.360 ;
        RECT 147.870 105.070 158.500 105.100 ;
        RECT 127.810 104.960 138.470 105.070 ;
        RECT 147.840 104.960 158.500 105.070 ;
        RECT 126.060 104.910 138.470 104.960 ;
        RECT 146.090 104.910 158.500 104.960 ;
        RECT 121.720 104.740 138.470 104.910 ;
        RECT 121.720 103.330 121.890 104.740 ;
        RECT 122.260 104.170 125.300 104.340 ;
        RECT 122.260 103.730 125.300 103.900 ;
        RECT 125.515 103.870 125.685 104.200 ;
        RECT 126.020 103.980 138.470 104.740 ;
        RECT 141.750 104.740 158.500 104.910 ;
        RECT 126.020 103.970 138.360 103.980 ;
        RECT 126.020 103.960 131.900 103.970 ;
        RECT 126.020 103.940 126.590 103.960 ;
        RECT 127.810 103.950 131.900 103.960 ;
        RECT 126.030 103.330 126.200 103.940 ;
        RECT 121.720 103.160 126.200 103.330 ;
        RECT 141.750 103.330 141.920 104.740 ;
        RECT 142.290 104.170 145.330 104.340 ;
        RECT 142.290 103.730 145.330 103.900 ;
        RECT 145.545 103.870 145.715 104.200 ;
        RECT 146.050 103.980 158.500 104.740 ;
        RECT 146.050 103.970 158.390 103.980 ;
        RECT 146.050 103.960 151.930 103.970 ;
        RECT 146.050 103.940 146.620 103.960 ;
        RECT 147.840 103.950 151.930 103.960 ;
        RECT 146.060 103.330 146.230 103.940 ;
        RECT 141.750 103.160 146.230 103.330 ;
        RECT 120.000 102.570 158.300 102.740 ;
        RECT 90.745 101.725 91.265 102.265 ;
        RECT 87.095 100.805 87.265 101.415 ;
        RECT 87.435 101.025 87.765 101.460 ;
        RECT 87.985 100.805 90.575 101.575 ;
        RECT 91.435 101.555 91.955 102.095 ;
        RECT 120.000 101.720 134.620 102.570 ;
        RECT 120.000 101.650 120.960 101.720 ;
        RECT 90.745 100.805 91.955 101.555 ;
        RECT 13.380 100.635 92.040 100.805 ;
        RECT 13.465 99.885 14.675 100.635 ;
        RECT 14.935 100.085 15.105 100.375 ;
        RECT 15.275 100.255 15.605 100.635 ;
        RECT 14.935 99.915 15.600 100.085 ;
        RECT 13.465 99.345 13.985 99.885 ;
        RECT 14.155 99.175 14.675 99.715 ;
        RECT 13.465 98.085 14.675 99.175 ;
        RECT 14.850 99.095 15.200 99.745 ;
        RECT 15.370 98.925 15.600 99.915 ;
        RECT 14.935 98.755 15.600 98.925 ;
        RECT 14.935 98.255 15.105 98.755 ;
        RECT 15.275 98.085 15.605 98.585 ;
        RECT 15.775 98.255 15.960 100.375 ;
        RECT 16.215 100.175 16.465 100.635 ;
        RECT 16.635 100.185 16.970 100.355 ;
        RECT 17.165 100.185 17.840 100.355 ;
        RECT 16.635 100.045 16.805 100.185 ;
        RECT 16.130 99.055 16.410 100.005 ;
        RECT 16.580 99.915 16.805 100.045 ;
        RECT 16.580 98.810 16.750 99.915 ;
        RECT 16.975 99.765 17.500 99.985 ;
        RECT 16.920 99.000 17.160 99.595 ;
        RECT 17.330 99.065 17.500 99.765 ;
        RECT 17.670 99.405 17.840 100.185 ;
        RECT 18.160 100.135 18.530 100.635 ;
        RECT 18.710 100.185 19.115 100.355 ;
        RECT 19.285 100.185 20.070 100.355 ;
        RECT 18.710 99.955 18.880 100.185 ;
        RECT 18.050 99.655 18.880 99.955 ;
        RECT 19.265 99.685 19.730 100.015 ;
        RECT 18.050 99.625 18.250 99.655 ;
        RECT 18.370 99.405 18.540 99.475 ;
        RECT 17.670 99.235 18.540 99.405 ;
        RECT 18.030 99.145 18.540 99.235 ;
        RECT 16.580 98.680 16.885 98.810 ;
        RECT 17.330 98.700 17.860 99.065 ;
        RECT 16.200 98.085 16.465 98.545 ;
        RECT 16.635 98.255 16.885 98.680 ;
        RECT 18.030 98.530 18.200 99.145 ;
        RECT 17.095 98.360 18.200 98.530 ;
        RECT 18.370 98.085 18.540 98.885 ;
        RECT 18.710 98.585 18.880 99.655 ;
        RECT 19.050 98.755 19.240 99.475 ;
        RECT 19.410 98.725 19.730 99.685 ;
        RECT 19.900 99.725 20.070 100.185 ;
        RECT 20.345 100.105 20.555 100.635 ;
        RECT 20.815 99.895 21.145 100.420 ;
        RECT 21.315 100.025 21.485 100.635 ;
        RECT 21.655 99.980 21.985 100.415 ;
        RECT 22.210 100.380 22.545 100.425 ;
        RECT 21.655 99.895 22.035 99.980 ;
        RECT 20.945 99.725 21.145 99.895 ;
        RECT 21.810 99.855 22.035 99.895 ;
        RECT 19.900 99.395 20.775 99.725 ;
        RECT 20.945 99.395 21.695 99.725 ;
        RECT 18.710 98.255 18.960 98.585 ;
        RECT 19.900 98.555 20.070 99.395 ;
        RECT 20.945 99.190 21.135 99.395 ;
        RECT 21.865 99.275 22.035 99.855 ;
        RECT 21.820 99.225 22.035 99.275 ;
        RECT 20.240 98.815 21.135 99.190 ;
        RECT 21.645 99.145 22.035 99.225 ;
        RECT 22.205 99.915 22.545 100.380 ;
        RECT 22.715 100.255 23.045 100.635 ;
        RECT 23.505 100.295 23.775 100.300 ;
        RECT 23.505 100.125 23.815 100.295 ;
        RECT 22.205 99.225 22.375 99.915 ;
        RECT 22.545 99.395 22.805 99.725 ;
        RECT 19.185 98.385 20.070 98.555 ;
        RECT 20.250 98.085 20.565 98.585 ;
        RECT 20.795 98.255 21.135 98.815 ;
        RECT 21.305 98.085 21.475 99.095 ;
        RECT 21.645 98.300 21.975 99.145 ;
        RECT 22.205 98.255 22.465 99.225 ;
        RECT 22.635 98.845 22.805 99.395 ;
        RECT 22.975 99.025 23.315 100.055 ;
        RECT 23.505 99.025 23.775 100.125 ;
        RECT 24.000 99.025 24.280 100.300 ;
        RECT 24.480 100.135 24.710 100.465 ;
        RECT 24.955 100.255 25.285 100.635 ;
        RECT 24.480 98.845 24.650 100.135 ;
        RECT 25.455 100.065 25.630 100.465 ;
        RECT 25.000 99.895 25.630 100.065 ;
        RECT 25.000 99.725 25.170 99.895 ;
        RECT 25.885 99.835 26.195 100.635 ;
        RECT 26.400 99.835 27.095 100.465 ;
        RECT 27.265 100.090 32.610 100.635 ;
        RECT 32.785 100.090 38.130 100.635 ;
        RECT 26.400 99.785 26.575 99.835 ;
        RECT 24.820 99.395 25.170 99.725 ;
        RECT 22.635 98.675 24.650 98.845 ;
        RECT 25.000 98.875 25.170 99.395 ;
        RECT 25.350 99.045 25.715 99.725 ;
        RECT 25.895 99.395 26.230 99.665 ;
        RECT 26.400 99.235 26.570 99.785 ;
        RECT 26.740 99.395 27.075 99.645 ;
        RECT 28.850 99.260 29.190 100.090 ;
        RECT 25.000 98.705 25.630 98.875 ;
        RECT 22.660 98.085 22.990 98.495 ;
        RECT 23.190 98.255 23.360 98.675 ;
        RECT 23.575 98.085 24.245 98.495 ;
        RECT 24.480 98.255 24.650 98.675 ;
        RECT 24.955 98.085 25.285 98.525 ;
        RECT 25.455 98.255 25.630 98.705 ;
        RECT 25.885 98.085 26.165 99.225 ;
        RECT 26.335 98.255 26.665 99.235 ;
        RECT 26.835 98.085 27.095 99.225 ;
        RECT 30.670 98.520 31.020 99.770 ;
        RECT 34.370 99.260 34.710 100.090 ;
        RECT 39.225 99.910 39.515 100.635 ;
        RECT 39.685 99.865 42.275 100.635 ;
        RECT 42.910 99.895 43.165 100.465 ;
        RECT 43.335 100.235 43.665 100.635 ;
        RECT 44.090 100.100 44.620 100.465 ;
        RECT 44.810 100.295 45.085 100.465 ;
        RECT 44.805 100.125 45.085 100.295 ;
        RECT 44.090 100.065 44.265 100.100 ;
        RECT 43.335 99.895 44.265 100.065 ;
        RECT 36.190 98.520 36.540 99.770 ;
        RECT 39.685 99.345 40.895 99.865 ;
        RECT 27.265 98.085 32.610 98.520 ;
        RECT 32.785 98.085 38.130 98.520 ;
        RECT 39.225 98.085 39.515 99.250 ;
        RECT 41.065 99.175 42.275 99.695 ;
        RECT 39.685 98.085 42.275 99.175 ;
        RECT 42.910 99.225 43.080 99.895 ;
        RECT 43.335 99.725 43.505 99.895 ;
        RECT 43.250 99.395 43.505 99.725 ;
        RECT 43.730 99.395 43.925 99.725 ;
        RECT 42.910 98.255 43.245 99.225 ;
        RECT 43.415 98.085 43.585 99.225 ;
        RECT 43.755 98.425 43.925 99.395 ;
        RECT 44.095 98.765 44.265 99.895 ;
        RECT 44.435 99.105 44.605 99.905 ;
        RECT 44.810 99.305 45.085 100.125 ;
        RECT 45.255 99.105 45.445 100.465 ;
        RECT 45.625 100.100 46.135 100.635 ;
        RECT 46.355 99.825 46.600 100.430 ;
        RECT 47.135 100.085 47.305 100.375 ;
        RECT 47.475 100.255 47.805 100.635 ;
        RECT 47.135 99.915 47.800 100.085 ;
        RECT 45.645 99.655 46.875 99.825 ;
        RECT 44.435 98.935 45.445 99.105 ;
        RECT 45.615 99.090 46.365 99.280 ;
        RECT 44.095 98.595 45.220 98.765 ;
        RECT 45.615 98.425 45.785 99.090 ;
        RECT 46.535 98.845 46.875 99.655 ;
        RECT 47.050 99.095 47.400 99.745 ;
        RECT 47.570 98.925 47.800 99.915 ;
        RECT 43.755 98.255 45.785 98.425 ;
        RECT 45.955 98.085 46.125 98.845 ;
        RECT 46.360 98.435 46.875 98.845 ;
        RECT 47.135 98.755 47.800 98.925 ;
        RECT 47.135 98.255 47.305 98.755 ;
        RECT 47.475 98.085 47.805 98.585 ;
        RECT 47.975 98.255 48.160 100.375 ;
        RECT 48.415 100.175 48.665 100.635 ;
        RECT 48.835 100.185 49.170 100.355 ;
        RECT 49.365 100.185 50.040 100.355 ;
        RECT 48.835 100.045 49.005 100.185 ;
        RECT 48.330 99.055 48.610 100.005 ;
        RECT 48.780 99.915 49.005 100.045 ;
        RECT 48.780 98.810 48.950 99.915 ;
        RECT 49.175 99.765 49.700 99.985 ;
        RECT 49.120 99.000 49.360 99.595 ;
        RECT 49.530 99.065 49.700 99.765 ;
        RECT 49.870 99.405 50.040 100.185 ;
        RECT 50.360 100.135 50.730 100.635 ;
        RECT 50.910 100.185 51.315 100.355 ;
        RECT 51.485 100.185 52.270 100.355 ;
        RECT 50.910 99.955 51.080 100.185 ;
        RECT 50.250 99.655 51.080 99.955 ;
        RECT 51.465 99.685 51.930 100.015 ;
        RECT 50.250 99.625 50.450 99.655 ;
        RECT 50.570 99.405 50.740 99.475 ;
        RECT 49.870 99.235 50.740 99.405 ;
        RECT 50.230 99.145 50.740 99.235 ;
        RECT 48.780 98.680 49.085 98.810 ;
        RECT 49.530 98.700 50.060 99.065 ;
        RECT 48.400 98.085 48.665 98.545 ;
        RECT 48.835 98.255 49.085 98.680 ;
        RECT 50.230 98.530 50.400 99.145 ;
        RECT 49.295 98.360 50.400 98.530 ;
        RECT 50.570 98.085 50.740 98.885 ;
        RECT 50.910 98.585 51.080 99.655 ;
        RECT 51.250 98.755 51.440 99.475 ;
        RECT 51.610 98.725 51.930 99.685 ;
        RECT 52.100 99.725 52.270 100.185 ;
        RECT 52.545 100.105 52.755 100.635 ;
        RECT 53.015 99.895 53.345 100.420 ;
        RECT 53.515 100.025 53.685 100.635 ;
        RECT 53.855 99.980 54.185 100.415 ;
        RECT 54.590 100.155 54.760 100.635 ;
        RECT 54.930 99.985 55.260 100.455 ;
        RECT 55.430 100.155 55.600 100.635 ;
        RECT 55.770 99.985 56.100 100.455 ;
        RECT 53.855 99.895 54.235 99.980 ;
        RECT 53.145 99.725 53.345 99.895 ;
        RECT 54.010 99.855 54.235 99.895 ;
        RECT 52.100 99.395 52.975 99.725 ;
        RECT 53.145 99.395 53.895 99.725 ;
        RECT 50.910 98.255 51.160 98.585 ;
        RECT 52.100 98.555 52.270 99.395 ;
        RECT 53.145 99.190 53.335 99.395 ;
        RECT 54.065 99.275 54.235 99.855 ;
        RECT 54.020 99.225 54.235 99.275 ;
        RECT 52.440 98.815 53.335 99.190 ;
        RECT 53.845 99.145 54.235 99.225 ;
        RECT 54.405 99.815 56.100 99.985 ;
        RECT 56.310 99.895 56.480 100.635 ;
        RECT 56.695 99.895 57.025 100.430 ;
        RECT 57.195 100.125 57.435 100.635 ;
        RECT 57.715 100.085 57.885 100.375 ;
        RECT 58.055 100.255 58.385 100.635 ;
        RECT 54.405 99.225 54.750 99.815 ;
        RECT 54.920 99.475 56.130 99.645 ;
        RECT 55.925 99.225 56.130 99.475 ;
        RECT 56.300 99.395 56.675 99.725 ;
        RECT 56.845 99.225 57.025 99.895 ;
        RECT 57.195 99.395 57.450 99.955 ;
        RECT 57.715 99.915 58.380 100.085 ;
        RECT 51.385 98.385 52.270 98.555 ;
        RECT 52.450 98.085 52.765 98.585 ;
        RECT 52.995 98.255 53.335 98.815 ;
        RECT 53.505 98.085 53.675 99.095 ;
        RECT 53.845 98.300 54.175 99.145 ;
        RECT 54.405 99.055 55.260 99.225 ;
        RECT 55.925 99.055 57.385 99.225 ;
        RECT 57.630 99.095 57.980 99.745 ;
        RECT 54.930 98.885 55.260 99.055 ;
        RECT 54.590 98.085 54.760 98.885 ;
        RECT 54.930 98.715 56.100 98.885 ;
        RECT 54.930 98.255 55.260 98.715 ;
        RECT 55.430 98.085 55.600 98.545 ;
        RECT 55.770 98.255 56.100 98.715 ;
        RECT 56.310 98.085 56.480 98.885 ;
        RECT 57.025 98.255 57.385 99.055 ;
        RECT 58.150 98.925 58.380 99.915 ;
        RECT 57.715 98.755 58.380 98.925 ;
        RECT 57.715 98.255 57.885 98.755 ;
        RECT 58.055 98.085 58.385 98.585 ;
        RECT 58.555 98.255 58.740 100.375 ;
        RECT 58.995 100.175 59.245 100.635 ;
        RECT 59.415 100.185 59.750 100.355 ;
        RECT 59.945 100.185 60.620 100.355 ;
        RECT 59.415 100.045 59.585 100.185 ;
        RECT 58.910 99.055 59.190 100.005 ;
        RECT 59.360 99.915 59.585 100.045 ;
        RECT 59.360 98.810 59.530 99.915 ;
        RECT 59.755 99.765 60.280 99.985 ;
        RECT 59.700 99.000 59.940 99.595 ;
        RECT 60.110 99.065 60.280 99.765 ;
        RECT 60.450 99.405 60.620 100.185 ;
        RECT 60.940 100.135 61.310 100.635 ;
        RECT 61.490 100.185 61.895 100.355 ;
        RECT 62.065 100.185 62.850 100.355 ;
        RECT 61.490 99.955 61.660 100.185 ;
        RECT 60.830 99.655 61.660 99.955 ;
        RECT 62.045 99.685 62.510 100.015 ;
        RECT 60.830 99.625 61.030 99.655 ;
        RECT 61.150 99.405 61.320 99.475 ;
        RECT 60.450 99.235 61.320 99.405 ;
        RECT 60.810 99.145 61.320 99.235 ;
        RECT 59.360 98.680 59.665 98.810 ;
        RECT 60.110 98.700 60.640 99.065 ;
        RECT 58.980 98.085 59.245 98.545 ;
        RECT 59.415 98.255 59.665 98.680 ;
        RECT 60.810 98.530 60.980 99.145 ;
        RECT 59.875 98.360 60.980 98.530 ;
        RECT 61.150 98.085 61.320 98.885 ;
        RECT 61.490 98.585 61.660 99.655 ;
        RECT 61.830 98.755 62.020 99.475 ;
        RECT 62.190 98.725 62.510 99.685 ;
        RECT 62.680 99.725 62.850 100.185 ;
        RECT 63.125 100.105 63.335 100.635 ;
        RECT 63.595 99.895 63.925 100.420 ;
        RECT 64.095 100.025 64.265 100.635 ;
        RECT 64.435 99.980 64.765 100.415 ;
        RECT 64.435 99.895 64.815 99.980 ;
        RECT 64.985 99.910 65.275 100.635 ;
        RECT 63.725 99.725 63.925 99.895 ;
        RECT 64.590 99.855 64.815 99.895 ;
        RECT 62.680 99.395 63.555 99.725 ;
        RECT 63.725 99.395 64.475 99.725 ;
        RECT 61.490 98.255 61.740 98.585 ;
        RECT 62.680 98.555 62.850 99.395 ;
        RECT 63.725 99.190 63.915 99.395 ;
        RECT 64.645 99.275 64.815 99.855 ;
        RECT 64.600 99.225 64.815 99.275 ;
        RECT 65.450 99.895 65.705 100.465 ;
        RECT 65.875 100.235 66.205 100.635 ;
        RECT 66.630 100.100 67.160 100.465 ;
        RECT 66.630 100.065 66.805 100.100 ;
        RECT 65.875 99.895 66.805 100.065 ;
        RECT 63.020 98.815 63.915 99.190 ;
        RECT 64.425 99.145 64.815 99.225 ;
        RECT 61.965 98.385 62.850 98.555 ;
        RECT 63.030 98.085 63.345 98.585 ;
        RECT 63.575 98.255 63.915 98.815 ;
        RECT 64.085 98.085 64.255 99.095 ;
        RECT 64.425 98.300 64.755 99.145 ;
        RECT 64.985 98.085 65.275 99.250 ;
        RECT 65.450 99.225 65.620 99.895 ;
        RECT 65.875 99.725 66.045 99.895 ;
        RECT 65.790 99.395 66.045 99.725 ;
        RECT 66.270 99.395 66.465 99.725 ;
        RECT 65.450 98.255 65.785 99.225 ;
        RECT 65.955 98.085 66.125 99.225 ;
        RECT 66.295 98.425 66.465 99.395 ;
        RECT 66.635 98.765 66.805 99.895 ;
        RECT 66.975 99.105 67.145 99.905 ;
        RECT 67.350 99.615 67.625 100.465 ;
        RECT 67.345 99.445 67.625 99.615 ;
        RECT 67.350 99.305 67.625 99.445 ;
        RECT 67.795 99.105 67.985 100.465 ;
        RECT 68.165 100.100 68.675 100.635 ;
        RECT 68.895 99.825 69.140 100.430 ;
        RECT 69.585 99.865 71.255 100.635 ;
        RECT 71.885 99.895 72.375 100.465 ;
        RECT 72.545 100.065 72.775 100.465 ;
        RECT 72.945 100.235 73.365 100.635 ;
        RECT 73.535 100.065 73.705 100.465 ;
        RECT 72.545 99.895 73.705 100.065 ;
        RECT 73.875 99.895 74.325 100.635 ;
        RECT 74.495 99.895 74.935 100.455 ;
        RECT 75.155 100.165 75.445 100.635 ;
        RECT 75.615 99.995 75.945 100.465 ;
        RECT 76.115 100.165 76.285 100.635 ;
        RECT 76.455 99.995 76.785 100.465 ;
        RECT 75.615 99.985 76.785 99.995 ;
        RECT 68.185 99.655 69.415 99.825 ;
        RECT 66.975 98.935 67.985 99.105 ;
        RECT 68.155 99.090 68.905 99.280 ;
        RECT 66.635 98.595 67.760 98.765 ;
        RECT 68.155 98.425 68.325 99.090 ;
        RECT 69.075 98.845 69.415 99.655 ;
        RECT 69.585 99.345 70.335 99.865 ;
        RECT 70.505 99.175 71.255 99.695 ;
        RECT 66.295 98.255 68.325 98.425 ;
        RECT 68.495 98.085 68.665 98.845 ;
        RECT 68.900 98.435 69.415 98.845 ;
        RECT 69.585 98.085 71.255 99.175 ;
        RECT 71.885 99.225 72.055 99.895 ;
        RECT 72.225 99.395 72.630 99.725 ;
        RECT 71.885 99.055 72.655 99.225 ;
        RECT 71.895 98.085 72.225 98.885 ;
        RECT 72.405 98.425 72.655 99.055 ;
        RECT 72.845 98.595 73.095 99.725 ;
        RECT 73.295 99.395 73.540 99.725 ;
        RECT 73.725 99.445 74.115 99.725 ;
        RECT 73.295 98.595 73.495 99.395 ;
        RECT 74.285 99.275 74.455 99.725 ;
        RECT 73.665 99.105 74.455 99.275 ;
        RECT 73.665 98.425 73.835 99.105 ;
        RECT 72.405 98.255 73.835 98.425 ;
        RECT 74.005 98.085 74.320 98.935 ;
        RECT 74.625 98.885 74.935 99.895 ;
        RECT 75.185 99.815 76.785 99.985 ;
        RECT 76.955 99.815 77.230 100.635 ;
        RECT 77.410 99.960 77.685 100.305 ;
        RECT 77.875 100.235 78.255 100.635 ;
        RECT 78.425 100.065 78.595 100.415 ;
        RECT 78.765 100.235 79.095 100.635 ;
        RECT 79.265 100.065 79.520 100.415 ;
        RECT 79.725 100.125 79.965 100.635 ;
        RECT 80.135 100.125 80.425 100.465 ;
        RECT 80.655 100.125 80.970 100.635 ;
        RECT 75.185 99.275 75.400 99.815 ;
        RECT 75.570 99.445 76.340 99.645 ;
        RECT 76.510 99.445 77.230 99.645 ;
        RECT 75.185 99.055 75.945 99.275 ;
        RECT 74.495 98.255 74.935 98.885 ;
        RECT 75.145 98.425 75.445 98.885 ;
        RECT 75.615 98.595 75.945 99.055 ;
        RECT 76.115 99.055 77.230 99.265 ;
        RECT 76.115 98.425 76.285 99.055 ;
        RECT 75.145 98.255 76.285 98.425 ;
        RECT 76.455 98.085 76.785 98.885 ;
        RECT 76.955 98.255 77.230 99.055 ;
        RECT 77.410 99.225 77.580 99.960 ;
        RECT 77.855 99.895 79.520 100.065 ;
        RECT 77.855 99.725 78.025 99.895 ;
        RECT 77.750 99.395 78.025 99.725 ;
        RECT 78.195 99.395 79.020 99.725 ;
        RECT 79.190 99.395 79.535 99.725 ;
        RECT 79.770 99.615 79.965 99.955 ;
        RECT 79.765 99.445 79.965 99.615 ;
        RECT 79.770 99.395 79.965 99.445 ;
        RECT 77.855 99.225 78.025 99.395 ;
        RECT 77.410 98.255 77.685 99.225 ;
        RECT 77.855 99.055 78.515 99.225 ;
        RECT 78.825 99.105 79.020 99.395 ;
        RECT 80.135 99.225 80.315 100.125 ;
        RECT 81.140 100.065 81.310 100.335 ;
        RECT 81.480 100.235 81.810 100.635 ;
        RECT 80.485 99.395 80.895 99.955 ;
        RECT 81.140 99.895 81.835 100.065 ;
        RECT 81.065 99.225 81.235 99.725 ;
        RECT 78.345 98.935 78.515 99.055 ;
        RECT 79.190 98.935 79.515 99.225 ;
        RECT 77.895 98.085 78.175 98.885 ;
        RECT 78.345 98.765 79.515 98.935 ;
        RECT 79.775 99.055 81.235 99.225 ;
        RECT 79.775 98.880 80.135 99.055 ;
        RECT 81.405 98.885 81.835 99.895 ;
        RECT 78.345 98.305 79.535 98.595 ;
        RECT 80.720 98.085 80.890 98.885 ;
        RECT 81.060 98.715 81.835 98.885 ;
        RECT 82.470 99.895 82.725 100.465 ;
        RECT 82.895 100.235 83.225 100.635 ;
        RECT 83.650 100.100 84.180 100.465 ;
        RECT 84.370 100.295 84.645 100.465 ;
        RECT 84.365 100.125 84.645 100.295 ;
        RECT 83.650 100.065 83.825 100.100 ;
        RECT 82.895 99.895 83.825 100.065 ;
        RECT 82.470 99.225 82.640 99.895 ;
        RECT 82.895 99.725 83.065 99.895 ;
        RECT 82.810 99.395 83.065 99.725 ;
        RECT 83.290 99.395 83.485 99.725 ;
        RECT 81.060 98.255 81.390 98.715 ;
        RECT 81.560 98.085 81.730 98.545 ;
        RECT 82.470 98.255 82.805 99.225 ;
        RECT 82.975 98.085 83.145 99.225 ;
        RECT 83.315 98.425 83.485 99.395 ;
        RECT 83.655 98.765 83.825 99.895 ;
        RECT 83.995 99.105 84.165 99.905 ;
        RECT 84.370 99.305 84.645 100.125 ;
        RECT 84.815 99.105 85.005 100.465 ;
        RECT 85.185 100.100 85.695 100.635 ;
        RECT 85.915 99.825 86.160 100.430 ;
        RECT 86.605 99.865 90.115 100.635 ;
        RECT 90.745 99.885 91.955 100.635 ;
        RECT 100.030 100.395 112.740 101.005 ;
        RECT 85.205 99.655 86.435 99.825 ;
        RECT 83.995 98.935 85.005 99.105 ;
        RECT 85.175 99.090 85.925 99.280 ;
        RECT 83.655 98.595 84.780 98.765 ;
        RECT 85.175 98.425 85.345 99.090 ;
        RECT 86.095 98.845 86.435 99.655 ;
        RECT 86.605 99.345 88.255 99.865 ;
        RECT 88.425 99.175 90.115 99.695 ;
        RECT 83.315 98.255 85.345 98.425 ;
        RECT 85.515 98.085 85.685 98.845 ;
        RECT 85.920 98.435 86.435 98.845 ;
        RECT 86.605 98.085 90.115 99.175 ;
        RECT 90.745 99.175 91.265 99.715 ;
        RECT 91.435 99.345 91.955 99.885 ;
        RECT 99.980 100.195 112.790 100.395 ;
        RECT 90.745 98.085 91.955 99.175 ;
        RECT 13.380 97.915 92.040 98.085 ;
        RECT 13.465 96.825 14.675 97.915 ;
        RECT 14.845 96.825 18.355 97.915 ;
        RECT 13.465 96.115 13.985 96.655 ;
        RECT 14.155 96.285 14.675 96.825 ;
        RECT 14.845 96.135 16.495 96.655 ;
        RECT 16.665 96.305 18.355 96.825 ;
        RECT 18.530 96.775 18.850 97.915 ;
        RECT 19.030 96.605 19.225 97.655 ;
        RECT 19.405 97.065 19.735 97.745 ;
        RECT 19.935 97.115 20.190 97.915 ;
        RECT 19.405 96.785 19.755 97.065 ;
        RECT 18.590 96.555 18.850 96.605 ;
        RECT 18.585 96.385 18.850 96.555 ;
        RECT 18.590 96.275 18.850 96.385 ;
        RECT 19.030 96.275 19.415 96.605 ;
        RECT 19.585 96.405 19.755 96.785 ;
        RECT 19.945 96.575 20.190 96.935 ;
        RECT 20.365 96.775 20.750 97.745 ;
        RECT 20.920 97.455 21.245 97.915 ;
        RECT 21.765 97.285 22.045 97.745 ;
        RECT 20.920 97.065 22.045 97.285 ;
        RECT 19.585 96.235 20.105 96.405 ;
        RECT 13.465 95.365 14.675 96.115 ;
        RECT 14.845 95.365 18.355 96.135 ;
        RECT 18.530 95.895 19.745 96.065 ;
        RECT 18.530 95.545 18.820 95.895 ;
        RECT 19.015 95.365 19.345 95.725 ;
        RECT 19.515 95.590 19.745 95.895 ;
        RECT 19.935 95.670 20.105 96.235 ;
        RECT 20.365 96.105 20.645 96.775 ;
        RECT 20.920 96.605 21.370 97.065 ;
        RECT 22.235 96.895 22.635 97.745 ;
        RECT 23.035 97.455 23.305 97.915 ;
        RECT 23.475 97.285 23.760 97.745 ;
        RECT 20.815 96.275 21.370 96.605 ;
        RECT 21.540 96.335 22.635 96.895 ;
        RECT 20.920 96.165 21.370 96.275 ;
        RECT 20.365 95.535 20.750 96.105 ;
        RECT 20.920 95.995 22.045 96.165 ;
        RECT 20.920 95.365 21.245 95.825 ;
        RECT 21.765 95.535 22.045 95.995 ;
        RECT 22.235 95.535 22.635 96.335 ;
        RECT 22.805 97.065 23.760 97.285 ;
        RECT 22.805 96.165 23.015 97.065 ;
        RECT 23.185 96.335 23.875 96.895 ;
        RECT 24.045 96.825 25.715 97.915 ;
        RECT 22.805 95.995 23.760 96.165 ;
        RECT 23.035 95.365 23.305 95.825 ;
        RECT 23.475 95.535 23.760 95.995 ;
        RECT 24.045 96.135 24.795 96.655 ;
        RECT 24.965 96.305 25.715 96.825 ;
        RECT 26.345 96.750 26.635 97.915 ;
        RECT 26.805 97.480 32.150 97.915 ;
        RECT 24.045 95.365 25.715 96.135 ;
        RECT 26.345 95.365 26.635 96.090 ;
        RECT 28.390 95.910 28.730 96.740 ;
        RECT 30.210 96.230 30.560 97.480 ;
        RECT 32.325 96.825 33.995 97.915 ;
        RECT 34.255 97.245 34.425 97.745 ;
        RECT 34.595 97.415 34.925 97.915 ;
        RECT 34.255 97.075 34.920 97.245 ;
        RECT 32.325 96.135 33.075 96.655 ;
        RECT 33.245 96.305 33.995 96.825 ;
        RECT 34.170 96.255 34.520 96.905 ;
        RECT 26.805 95.365 32.150 95.910 ;
        RECT 32.325 95.365 33.995 96.135 ;
        RECT 34.690 96.085 34.920 97.075 ;
        RECT 34.255 95.915 34.920 96.085 ;
        RECT 34.255 95.625 34.425 95.915 ;
        RECT 34.595 95.365 34.925 95.745 ;
        RECT 35.095 95.625 35.280 97.745 ;
        RECT 35.520 97.455 35.785 97.915 ;
        RECT 35.955 97.320 36.205 97.745 ;
        RECT 36.415 97.470 37.520 97.640 ;
        RECT 35.900 97.190 36.205 97.320 ;
        RECT 35.450 95.995 35.730 96.945 ;
        RECT 35.900 96.085 36.070 97.190 ;
        RECT 36.240 96.405 36.480 97.000 ;
        RECT 36.650 96.935 37.180 97.300 ;
        RECT 36.650 96.235 36.820 96.935 ;
        RECT 37.350 96.855 37.520 97.470 ;
        RECT 37.690 97.115 37.860 97.915 ;
        RECT 38.030 97.415 38.280 97.745 ;
        RECT 38.505 97.445 39.390 97.615 ;
        RECT 37.350 96.765 37.860 96.855 ;
        RECT 35.900 95.955 36.125 96.085 ;
        RECT 36.295 96.015 36.820 96.235 ;
        RECT 36.990 96.595 37.860 96.765 ;
        RECT 35.535 95.365 35.785 95.825 ;
        RECT 35.955 95.815 36.125 95.955 ;
        RECT 36.990 95.815 37.160 96.595 ;
        RECT 37.690 96.525 37.860 96.595 ;
        RECT 37.370 96.345 37.570 96.375 ;
        RECT 38.030 96.345 38.200 97.415 ;
        RECT 38.370 96.525 38.560 97.245 ;
        RECT 37.370 96.045 38.200 96.345 ;
        RECT 38.730 96.315 39.050 97.275 ;
        RECT 35.955 95.645 36.290 95.815 ;
        RECT 36.485 95.645 37.160 95.815 ;
        RECT 37.480 95.365 37.850 95.865 ;
        RECT 38.030 95.815 38.200 96.045 ;
        RECT 38.585 95.985 39.050 96.315 ;
        RECT 39.220 96.605 39.390 97.445 ;
        RECT 39.570 97.415 39.885 97.915 ;
        RECT 40.115 97.185 40.455 97.745 ;
        RECT 39.560 96.810 40.455 97.185 ;
        RECT 40.625 96.905 40.795 97.915 ;
        RECT 40.265 96.605 40.455 96.810 ;
        RECT 40.965 96.855 41.295 97.700 ;
        RECT 40.965 96.775 41.355 96.855 ;
        RECT 41.140 96.725 41.355 96.775 ;
        RECT 39.220 96.275 40.095 96.605 ;
        RECT 40.265 96.275 41.015 96.605 ;
        RECT 39.220 95.815 39.390 96.275 ;
        RECT 40.265 96.105 40.465 96.275 ;
        RECT 41.185 96.145 41.355 96.725 ;
        RECT 41.130 96.105 41.355 96.145 ;
        RECT 38.030 95.645 38.435 95.815 ;
        RECT 38.605 95.645 39.390 95.815 ;
        RECT 39.665 95.365 39.875 95.895 ;
        RECT 40.135 95.580 40.465 96.105 ;
        RECT 40.975 96.020 41.355 96.105 ;
        RECT 41.525 96.775 41.910 97.745 ;
        RECT 42.080 97.455 42.405 97.915 ;
        RECT 42.925 97.285 43.205 97.745 ;
        RECT 42.080 97.065 43.205 97.285 ;
        RECT 41.525 96.105 41.805 96.775 ;
        RECT 42.080 96.605 42.530 97.065 ;
        RECT 43.395 96.895 43.795 97.745 ;
        RECT 44.195 97.455 44.465 97.915 ;
        RECT 44.635 97.285 44.920 97.745 ;
        RECT 41.975 96.275 42.530 96.605 ;
        RECT 42.700 96.335 43.795 96.895 ;
        RECT 42.080 96.165 42.530 96.275 ;
        RECT 40.635 95.365 40.805 95.975 ;
        RECT 40.975 95.585 41.305 96.020 ;
        RECT 41.525 95.535 41.910 96.105 ;
        RECT 42.080 95.995 43.205 96.165 ;
        RECT 42.080 95.365 42.405 95.825 ;
        RECT 42.925 95.535 43.205 95.995 ;
        RECT 43.395 95.535 43.795 96.335 ;
        RECT 43.965 97.065 44.920 97.285 ;
        RECT 43.965 96.165 44.175 97.065 ;
        RECT 44.345 96.335 45.035 96.895 ;
        RECT 45.205 96.825 47.795 97.915 ;
        RECT 43.965 95.995 44.920 96.165 ;
        RECT 44.195 95.365 44.465 95.825 ;
        RECT 44.635 95.535 44.920 95.995 ;
        RECT 45.205 96.135 46.415 96.655 ;
        RECT 46.585 96.305 47.795 96.825 ;
        RECT 47.970 96.775 48.305 97.745 ;
        RECT 48.475 96.775 48.645 97.915 ;
        RECT 48.815 97.575 50.845 97.745 ;
        RECT 45.205 95.365 47.795 96.135 ;
        RECT 47.970 96.105 48.140 96.775 ;
        RECT 48.815 96.605 48.985 97.575 ;
        RECT 48.310 96.275 48.565 96.605 ;
        RECT 48.790 96.275 48.985 96.605 ;
        RECT 49.155 97.235 50.280 97.405 ;
        RECT 48.395 96.105 48.565 96.275 ;
        RECT 49.155 96.105 49.325 97.235 ;
        RECT 47.970 95.535 48.225 96.105 ;
        RECT 48.395 95.935 49.325 96.105 ;
        RECT 49.495 96.895 50.505 97.065 ;
        RECT 49.495 96.095 49.665 96.895 ;
        RECT 49.870 96.215 50.145 96.695 ;
        RECT 49.865 96.045 50.145 96.215 ;
        RECT 49.150 95.900 49.325 95.935 ;
        RECT 48.395 95.365 48.725 95.765 ;
        RECT 49.150 95.535 49.680 95.900 ;
        RECT 49.870 95.535 50.145 96.045 ;
        RECT 50.315 95.535 50.505 96.895 ;
        RECT 50.675 96.910 50.845 97.575 ;
        RECT 51.015 97.155 51.185 97.915 ;
        RECT 51.420 97.155 51.935 97.565 ;
        RECT 50.675 96.720 51.425 96.910 ;
        RECT 51.595 96.345 51.935 97.155 ;
        RECT 52.105 96.750 52.395 97.915 ;
        RECT 52.570 96.775 52.905 97.745 ;
        RECT 53.075 96.775 53.245 97.915 ;
        RECT 53.415 97.575 55.445 97.745 ;
        RECT 50.705 96.175 51.935 96.345 ;
        RECT 50.685 95.365 51.195 95.900 ;
        RECT 51.415 95.570 51.660 96.175 ;
        RECT 52.570 96.105 52.740 96.775 ;
        RECT 53.415 96.605 53.585 97.575 ;
        RECT 52.910 96.275 53.165 96.605 ;
        RECT 53.390 96.275 53.585 96.605 ;
        RECT 53.755 97.235 54.880 97.405 ;
        RECT 52.995 96.105 53.165 96.275 ;
        RECT 53.755 96.105 53.925 97.235 ;
        RECT 52.105 95.365 52.395 96.090 ;
        RECT 52.570 95.535 52.825 96.105 ;
        RECT 52.995 95.935 53.925 96.105 ;
        RECT 54.095 96.895 55.105 97.065 ;
        RECT 54.095 96.095 54.265 96.895 ;
        RECT 54.470 96.555 54.745 96.695 ;
        RECT 54.465 96.385 54.745 96.555 ;
        RECT 53.750 95.900 53.925 95.935 ;
        RECT 52.995 95.365 53.325 95.765 ;
        RECT 53.750 95.535 54.280 95.900 ;
        RECT 54.470 95.535 54.745 96.385 ;
        RECT 54.915 95.535 55.105 96.895 ;
        RECT 55.275 96.910 55.445 97.575 ;
        RECT 55.615 97.155 55.785 97.915 ;
        RECT 56.020 97.155 56.535 97.565 ;
        RECT 55.275 96.720 56.025 96.910 ;
        RECT 56.195 96.345 56.535 97.155 ;
        RECT 56.705 96.825 60.215 97.915 ;
        RECT 60.385 96.825 61.595 97.915 ;
        RECT 61.880 97.285 62.165 97.745 ;
        RECT 62.335 97.455 62.605 97.915 ;
        RECT 61.880 97.065 62.835 97.285 ;
        RECT 55.305 96.175 56.535 96.345 ;
        RECT 55.285 95.365 55.795 95.900 ;
        RECT 56.015 95.570 56.260 96.175 ;
        RECT 56.705 96.135 58.355 96.655 ;
        RECT 58.525 96.305 60.215 96.825 ;
        RECT 56.705 95.365 60.215 96.135 ;
        RECT 60.385 96.115 60.905 96.655 ;
        RECT 61.075 96.285 61.595 96.825 ;
        RECT 61.765 96.335 62.455 96.895 ;
        RECT 62.625 96.165 62.835 97.065 ;
        RECT 60.385 95.365 61.595 96.115 ;
        RECT 61.880 95.995 62.835 96.165 ;
        RECT 63.005 96.895 63.405 97.745 ;
        RECT 63.595 97.285 63.875 97.745 ;
        RECT 64.395 97.455 64.720 97.915 ;
        RECT 63.595 97.065 64.720 97.285 ;
        RECT 63.005 96.335 64.100 96.895 ;
        RECT 64.270 96.605 64.720 97.065 ;
        RECT 64.890 96.775 65.275 97.745 ;
        RECT 65.445 96.825 67.115 97.915 ;
        RECT 61.880 95.535 62.165 95.995 ;
        RECT 62.335 95.365 62.605 95.825 ;
        RECT 63.005 95.535 63.405 96.335 ;
        RECT 64.270 96.275 64.825 96.605 ;
        RECT 64.270 96.165 64.720 96.275 ;
        RECT 63.595 95.995 64.720 96.165 ;
        RECT 64.995 96.105 65.275 96.775 ;
        RECT 63.595 95.535 63.875 95.995 ;
        RECT 64.395 95.365 64.720 95.825 ;
        RECT 64.890 95.535 65.275 96.105 ;
        RECT 65.445 96.135 66.195 96.655 ;
        RECT 66.365 96.305 67.115 96.825 ;
        RECT 67.285 97.045 67.560 97.745 ;
        RECT 67.730 97.370 67.985 97.915 ;
        RECT 68.155 97.405 68.635 97.745 ;
        RECT 68.810 97.360 69.415 97.915 ;
        RECT 68.800 97.260 69.415 97.360 ;
        RECT 68.800 97.235 68.985 97.260 ;
        RECT 65.445 95.365 67.115 96.135 ;
        RECT 67.285 96.015 67.455 97.045 ;
        RECT 67.730 96.915 68.485 97.165 ;
        RECT 68.655 96.990 68.985 97.235 ;
        RECT 67.730 96.880 68.500 96.915 ;
        RECT 67.730 96.870 68.515 96.880 ;
        RECT 67.625 96.855 68.520 96.870 ;
        RECT 67.625 96.840 68.540 96.855 ;
        RECT 67.625 96.830 68.560 96.840 ;
        RECT 67.625 96.820 68.585 96.830 ;
        RECT 67.625 96.790 68.655 96.820 ;
        RECT 67.625 96.760 68.675 96.790 ;
        RECT 67.625 96.730 68.695 96.760 ;
        RECT 67.625 96.705 68.725 96.730 ;
        RECT 67.625 96.670 68.760 96.705 ;
        RECT 67.625 96.665 68.790 96.670 ;
        RECT 67.625 96.270 67.855 96.665 ;
        RECT 68.400 96.660 68.790 96.665 ;
        RECT 68.425 96.650 68.790 96.660 ;
        RECT 68.440 96.645 68.790 96.650 ;
        RECT 68.455 96.640 68.790 96.645 ;
        RECT 69.155 96.640 69.415 97.090 ;
        RECT 69.595 96.945 69.925 97.730 ;
        RECT 69.595 96.775 70.275 96.945 ;
        RECT 70.455 96.775 70.785 97.915 ;
        RECT 70.965 96.825 73.555 97.915 ;
        RECT 74.185 97.405 75.375 97.695 ;
        RECT 68.455 96.635 69.415 96.640 ;
        RECT 68.465 96.625 69.415 96.635 ;
        RECT 68.475 96.620 69.415 96.625 ;
        RECT 68.485 96.610 69.415 96.620 ;
        RECT 68.490 96.600 69.415 96.610 ;
        RECT 68.495 96.595 69.415 96.600 ;
        RECT 68.505 96.580 69.415 96.595 ;
        RECT 68.510 96.565 69.415 96.580 ;
        RECT 68.520 96.540 69.415 96.565 ;
        RECT 68.025 96.070 68.355 96.495 ;
        RECT 67.285 95.535 67.545 96.015 ;
        RECT 67.715 95.365 67.965 95.905 ;
        RECT 68.135 95.585 68.355 96.070 ;
        RECT 68.525 96.470 69.415 96.540 ;
        RECT 68.525 95.745 68.695 96.470 ;
        RECT 69.585 96.355 69.935 96.605 ;
        RECT 68.865 95.915 69.415 96.300 ;
        RECT 70.105 96.175 70.275 96.775 ;
        RECT 70.445 96.355 70.795 96.605 ;
        RECT 68.525 95.575 69.415 95.745 ;
        RECT 69.605 95.365 69.845 96.175 ;
        RECT 70.015 95.535 70.345 96.175 ;
        RECT 70.515 95.365 70.785 96.175 ;
        RECT 70.965 96.135 72.175 96.655 ;
        RECT 72.345 96.305 73.555 96.825 ;
        RECT 74.205 97.065 75.375 97.235 ;
        RECT 75.545 97.115 75.825 97.915 ;
        RECT 74.205 96.775 74.530 97.065 ;
        RECT 75.205 96.945 75.375 97.065 ;
        RECT 74.700 96.605 74.895 96.895 ;
        RECT 75.205 96.775 75.865 96.945 ;
        RECT 76.035 96.775 76.310 97.745 ;
        RECT 76.485 96.825 77.695 97.915 ;
        RECT 75.695 96.605 75.865 96.775 ;
        RECT 74.185 96.275 74.530 96.605 ;
        RECT 74.700 96.275 75.525 96.605 ;
        RECT 75.695 96.275 75.970 96.605 ;
        RECT 70.965 95.365 73.555 96.135 ;
        RECT 75.695 96.105 75.865 96.275 ;
        RECT 74.200 95.935 75.865 96.105 ;
        RECT 76.140 96.040 76.310 96.775 ;
        RECT 74.200 95.585 74.455 95.935 ;
        RECT 74.625 95.365 74.955 95.765 ;
        RECT 75.125 95.585 75.295 95.935 ;
        RECT 75.465 95.365 75.845 95.765 ;
        RECT 76.035 95.695 76.310 96.040 ;
        RECT 76.485 96.115 77.005 96.655 ;
        RECT 77.175 96.285 77.695 96.825 ;
        RECT 77.865 96.750 78.155 97.915 ;
        RECT 79.245 97.155 79.760 97.565 ;
        RECT 79.995 97.155 80.165 97.915 ;
        RECT 80.335 97.575 82.365 97.745 ;
        RECT 79.245 96.345 79.585 97.155 ;
        RECT 80.335 96.910 80.505 97.575 ;
        RECT 80.900 97.235 82.025 97.405 ;
        RECT 79.755 96.720 80.505 96.910 ;
        RECT 80.675 96.895 81.685 97.065 ;
        RECT 79.245 96.175 80.475 96.345 ;
        RECT 76.485 95.365 77.695 96.115 ;
        RECT 77.865 95.365 78.155 96.090 ;
        RECT 79.520 95.570 79.765 96.175 ;
        RECT 79.985 95.365 80.495 95.900 ;
        RECT 80.675 95.535 80.865 96.895 ;
        RECT 81.035 95.875 81.310 96.695 ;
        RECT 81.515 96.095 81.685 96.895 ;
        RECT 81.855 96.105 82.025 97.235 ;
        RECT 82.195 96.605 82.365 97.575 ;
        RECT 82.535 96.775 82.705 97.915 ;
        RECT 82.875 96.775 83.210 97.745 ;
        RECT 83.385 97.480 88.730 97.915 ;
        RECT 82.195 96.275 82.390 96.605 ;
        RECT 82.615 96.275 82.870 96.605 ;
        RECT 82.615 96.105 82.785 96.275 ;
        RECT 83.040 96.105 83.210 96.775 ;
        RECT 81.855 95.935 82.785 96.105 ;
        RECT 81.855 95.900 82.030 95.935 ;
        RECT 81.035 95.705 81.315 95.875 ;
        RECT 81.035 95.535 81.310 95.705 ;
        RECT 81.500 95.535 82.030 95.900 ;
        RECT 82.455 95.365 82.785 95.765 ;
        RECT 82.955 95.535 83.210 96.105 ;
        RECT 84.970 95.910 85.310 96.740 ;
        RECT 86.790 96.230 87.140 97.480 ;
        RECT 88.905 96.825 90.575 97.915 ;
        RECT 88.905 96.135 89.655 96.655 ;
        RECT 89.825 96.305 90.575 96.825 ;
        RECT 90.745 96.825 91.955 97.915 ;
        RECT 90.745 96.285 91.265 96.825 ;
        RECT 83.385 95.365 88.730 95.910 ;
        RECT 88.905 95.365 90.575 96.135 ;
        RECT 91.435 96.115 91.955 96.655 ;
        RECT 90.745 95.365 91.955 96.115 ;
        RECT 13.380 95.195 92.040 95.365 ;
        RECT 13.465 94.445 14.675 95.195 ;
        RECT 14.845 94.445 16.055 95.195 ;
        RECT 16.230 94.455 16.485 95.025 ;
        RECT 16.655 94.795 16.985 95.195 ;
        RECT 17.410 94.660 17.940 95.025 ;
        RECT 17.410 94.625 17.585 94.660 ;
        RECT 16.655 94.455 17.585 94.625 ;
        RECT 13.465 93.905 13.985 94.445 ;
        RECT 14.155 93.735 14.675 94.275 ;
        RECT 14.845 93.905 15.365 94.445 ;
        RECT 15.535 93.735 16.055 94.275 ;
        RECT 13.465 92.645 14.675 93.735 ;
        RECT 14.845 92.645 16.055 93.735 ;
        RECT 16.230 93.785 16.400 94.455 ;
        RECT 16.655 94.285 16.825 94.455 ;
        RECT 16.570 93.955 16.825 94.285 ;
        RECT 17.050 93.955 17.245 94.285 ;
        RECT 16.230 92.815 16.565 93.785 ;
        RECT 16.735 92.645 16.905 93.785 ;
        RECT 17.075 92.985 17.245 93.955 ;
        RECT 17.415 93.325 17.585 94.455 ;
        RECT 17.755 93.665 17.925 94.465 ;
        RECT 18.130 94.175 18.405 95.025 ;
        RECT 18.125 94.005 18.405 94.175 ;
        RECT 18.130 93.865 18.405 94.005 ;
        RECT 18.575 93.665 18.765 95.025 ;
        RECT 18.945 94.660 19.455 95.195 ;
        RECT 19.675 94.385 19.920 94.990 ;
        RECT 20.845 94.625 21.100 94.975 ;
        RECT 21.270 94.795 21.600 95.195 ;
        RECT 21.770 94.625 21.940 94.975 ;
        RECT 22.110 94.795 22.490 95.195 ;
        RECT 20.845 94.455 22.510 94.625 ;
        RECT 22.680 94.520 22.955 94.865 ;
        RECT 18.965 94.215 20.195 94.385 ;
        RECT 22.340 94.285 22.510 94.455 ;
        RECT 17.755 93.495 18.765 93.665 ;
        RECT 18.935 93.650 19.685 93.840 ;
        RECT 17.415 93.155 18.540 93.325 ;
        RECT 18.935 92.985 19.105 93.650 ;
        RECT 19.855 93.405 20.195 94.215 ;
        RECT 20.825 93.955 21.175 94.285 ;
        RECT 21.345 93.955 22.170 94.285 ;
        RECT 22.340 93.955 22.615 94.285 ;
        RECT 17.075 92.815 19.105 92.985 ;
        RECT 19.275 92.645 19.445 93.405 ;
        RECT 19.680 92.995 20.195 93.405 ;
        RECT 20.845 93.495 21.175 93.785 ;
        RECT 21.345 93.665 21.570 93.955 ;
        RECT 22.340 93.785 22.510 93.955 ;
        RECT 22.785 93.785 22.955 94.520 ;
        RECT 23.125 94.365 23.415 95.195 ;
        RECT 23.585 94.425 26.175 95.195 ;
        RECT 26.435 94.645 26.605 94.935 ;
        RECT 26.775 94.815 27.105 95.195 ;
        RECT 26.435 94.475 27.100 94.645 ;
        RECT 23.585 93.905 24.795 94.425 ;
        RECT 21.840 93.615 22.510 93.785 ;
        RECT 21.840 93.495 22.010 93.615 ;
        RECT 20.845 93.325 22.010 93.495 ;
        RECT 20.825 92.865 22.020 93.155 ;
        RECT 22.190 92.645 22.470 93.445 ;
        RECT 22.680 92.815 22.955 93.785 ;
        RECT 23.125 92.645 23.415 93.850 ;
        RECT 24.965 93.735 26.175 94.255 ;
        RECT 23.585 92.645 26.175 93.735 ;
        RECT 26.350 93.655 26.700 94.305 ;
        RECT 26.870 93.485 27.100 94.475 ;
        RECT 26.435 93.315 27.100 93.485 ;
        RECT 26.435 92.815 26.605 93.315 ;
        RECT 26.775 92.645 27.105 93.145 ;
        RECT 27.275 92.815 27.460 94.935 ;
        RECT 27.715 94.735 27.965 95.195 ;
        RECT 28.135 94.745 28.470 94.915 ;
        RECT 28.665 94.745 29.340 94.915 ;
        RECT 28.135 94.605 28.305 94.745 ;
        RECT 27.630 93.615 27.910 94.565 ;
        RECT 28.080 94.475 28.305 94.605 ;
        RECT 28.080 93.370 28.250 94.475 ;
        RECT 28.475 94.325 29.000 94.545 ;
        RECT 28.420 93.560 28.660 94.155 ;
        RECT 28.830 93.625 29.000 94.325 ;
        RECT 29.170 93.965 29.340 94.745 ;
        RECT 29.660 94.695 30.030 95.195 ;
        RECT 30.210 94.745 30.615 94.915 ;
        RECT 30.785 94.745 31.570 94.915 ;
        RECT 30.210 94.515 30.380 94.745 ;
        RECT 29.550 94.215 30.380 94.515 ;
        RECT 30.765 94.245 31.230 94.575 ;
        RECT 29.550 94.185 29.750 94.215 ;
        RECT 29.870 93.965 30.040 94.035 ;
        RECT 29.170 93.795 30.040 93.965 ;
        RECT 29.530 93.705 30.040 93.795 ;
        RECT 28.080 93.240 28.385 93.370 ;
        RECT 28.830 93.260 29.360 93.625 ;
        RECT 27.700 92.645 27.965 93.105 ;
        RECT 28.135 92.815 28.385 93.240 ;
        RECT 29.530 93.090 29.700 93.705 ;
        RECT 28.595 92.920 29.700 93.090 ;
        RECT 29.870 92.645 30.040 93.445 ;
        RECT 30.210 93.145 30.380 94.215 ;
        RECT 30.550 93.315 30.740 94.035 ;
        RECT 30.910 93.285 31.230 94.245 ;
        RECT 31.400 94.285 31.570 94.745 ;
        RECT 31.845 94.665 32.055 95.195 ;
        RECT 32.315 94.455 32.645 94.980 ;
        RECT 32.815 94.585 32.985 95.195 ;
        RECT 33.155 94.540 33.485 94.975 ;
        RECT 33.655 94.680 33.825 95.195 ;
        RECT 33.155 94.455 33.535 94.540 ;
        RECT 32.445 94.285 32.645 94.455 ;
        RECT 33.310 94.415 33.535 94.455 ;
        RECT 31.400 93.955 32.275 94.285 ;
        RECT 32.445 93.955 33.195 94.285 ;
        RECT 30.210 92.815 30.460 93.145 ;
        RECT 31.400 93.115 31.570 93.955 ;
        RECT 32.445 93.750 32.635 93.955 ;
        RECT 33.365 93.835 33.535 94.415 ;
        RECT 33.320 93.785 33.535 93.835 ;
        RECT 31.740 93.375 32.635 93.750 ;
        RECT 33.145 93.705 33.535 93.785 ;
        RECT 35.090 94.455 35.345 95.025 ;
        RECT 35.515 94.795 35.845 95.195 ;
        RECT 36.270 94.660 36.800 95.025 ;
        RECT 36.990 94.855 37.265 95.025 ;
        RECT 36.985 94.685 37.265 94.855 ;
        RECT 36.270 94.625 36.445 94.660 ;
        RECT 35.515 94.455 36.445 94.625 ;
        RECT 35.090 93.785 35.260 94.455 ;
        RECT 35.515 94.285 35.685 94.455 ;
        RECT 35.430 93.955 35.685 94.285 ;
        RECT 35.910 93.955 36.105 94.285 ;
        RECT 30.685 92.945 31.570 93.115 ;
        RECT 31.750 92.645 32.065 93.145 ;
        RECT 32.295 92.815 32.635 93.375 ;
        RECT 32.805 92.645 32.975 93.655 ;
        RECT 33.145 92.860 33.475 93.705 ;
        RECT 33.645 92.645 33.815 93.560 ;
        RECT 35.090 92.815 35.425 93.785 ;
        RECT 35.595 92.645 35.765 93.785 ;
        RECT 35.935 92.985 36.105 93.955 ;
        RECT 36.275 93.325 36.445 94.455 ;
        RECT 36.615 93.665 36.785 94.465 ;
        RECT 36.990 93.865 37.265 94.685 ;
        RECT 37.435 93.665 37.625 95.025 ;
        RECT 37.805 94.660 38.315 95.195 ;
        RECT 38.535 94.385 38.780 94.990 ;
        RECT 39.225 94.470 39.515 95.195 ;
        RECT 40.150 94.455 40.405 95.025 ;
        RECT 40.575 94.795 40.905 95.195 ;
        RECT 41.330 94.660 41.860 95.025 ;
        RECT 41.330 94.625 41.505 94.660 ;
        RECT 40.575 94.455 41.505 94.625 ;
        RECT 37.825 94.215 39.055 94.385 ;
        RECT 36.615 93.495 37.625 93.665 ;
        RECT 37.795 93.650 38.545 93.840 ;
        RECT 36.275 93.155 37.400 93.325 ;
        RECT 37.795 92.985 37.965 93.650 ;
        RECT 38.715 93.405 39.055 94.215 ;
        RECT 35.935 92.815 37.965 92.985 ;
        RECT 38.135 92.645 38.305 93.405 ;
        RECT 38.540 92.995 39.055 93.405 ;
        RECT 39.225 92.645 39.515 93.810 ;
        RECT 40.150 93.785 40.320 94.455 ;
        RECT 40.575 94.285 40.745 94.455 ;
        RECT 40.490 93.955 40.745 94.285 ;
        RECT 40.970 93.955 41.165 94.285 ;
        RECT 40.150 92.815 40.485 93.785 ;
        RECT 40.655 92.645 40.825 93.785 ;
        RECT 40.995 92.985 41.165 93.955 ;
        RECT 41.335 93.325 41.505 94.455 ;
        RECT 41.675 93.665 41.845 94.465 ;
        RECT 42.050 94.175 42.325 95.025 ;
        RECT 42.045 94.005 42.325 94.175 ;
        RECT 42.050 93.865 42.325 94.005 ;
        RECT 42.495 93.665 42.685 95.025 ;
        RECT 42.865 94.660 43.375 95.195 ;
        RECT 43.595 94.385 43.840 94.990 ;
        RECT 44.285 94.815 45.175 94.985 ;
        RECT 42.885 94.215 44.115 94.385 ;
        RECT 44.285 94.260 44.835 94.645 ;
        RECT 41.675 93.495 42.685 93.665 ;
        RECT 42.855 93.650 43.605 93.840 ;
        RECT 41.335 93.155 42.460 93.325 ;
        RECT 42.855 92.985 43.025 93.650 ;
        RECT 43.775 93.405 44.115 94.215 ;
        RECT 45.005 94.090 45.175 94.815 ;
        RECT 44.285 94.020 45.175 94.090 ;
        RECT 45.345 94.490 45.565 94.975 ;
        RECT 45.735 94.655 45.985 95.195 ;
        RECT 46.155 94.545 46.415 95.025 ;
        RECT 46.585 94.650 51.930 95.195 ;
        RECT 45.345 94.065 45.675 94.490 ;
        RECT 44.285 93.995 45.180 94.020 ;
        RECT 44.285 93.980 45.190 93.995 ;
        RECT 44.285 93.965 45.195 93.980 ;
        RECT 44.285 93.960 45.205 93.965 ;
        RECT 44.285 93.950 45.210 93.960 ;
        RECT 44.285 93.940 45.215 93.950 ;
        RECT 44.285 93.935 45.225 93.940 ;
        RECT 44.285 93.925 45.235 93.935 ;
        RECT 44.285 93.920 45.245 93.925 ;
        RECT 44.285 93.470 44.545 93.920 ;
        RECT 44.910 93.915 45.245 93.920 ;
        RECT 44.910 93.910 45.260 93.915 ;
        RECT 44.910 93.900 45.275 93.910 ;
        RECT 44.910 93.895 45.300 93.900 ;
        RECT 45.845 93.895 46.075 94.290 ;
        RECT 44.910 93.890 46.075 93.895 ;
        RECT 44.940 93.855 46.075 93.890 ;
        RECT 44.975 93.830 46.075 93.855 ;
        RECT 45.005 93.800 46.075 93.830 ;
        RECT 45.025 93.770 46.075 93.800 ;
        RECT 45.045 93.740 46.075 93.770 ;
        RECT 45.115 93.730 46.075 93.740 ;
        RECT 45.140 93.720 46.075 93.730 ;
        RECT 45.160 93.705 46.075 93.720 ;
        RECT 45.180 93.690 46.075 93.705 ;
        RECT 45.185 93.680 45.970 93.690 ;
        RECT 45.200 93.645 45.970 93.680 ;
        RECT 40.995 92.815 43.025 92.985 ;
        RECT 43.195 92.645 43.365 93.405 ;
        RECT 43.600 92.995 44.115 93.405 ;
        RECT 44.715 93.325 45.045 93.570 ;
        RECT 45.215 93.395 45.970 93.645 ;
        RECT 46.245 93.515 46.415 94.545 ;
        RECT 48.170 93.820 48.510 94.650 ;
        RECT 52.105 94.425 54.695 95.195 ;
        RECT 55.375 94.540 55.705 94.975 ;
        RECT 55.875 94.585 56.045 95.195 ;
        RECT 55.325 94.455 55.705 94.540 ;
        RECT 56.215 94.455 56.545 94.980 ;
        RECT 56.805 94.665 57.015 95.195 ;
        RECT 57.290 94.745 58.075 94.915 ;
        RECT 58.245 94.745 58.650 94.915 ;
        RECT 44.715 93.300 44.900 93.325 ;
        RECT 44.285 93.200 44.900 93.300 ;
        RECT 44.285 92.645 44.890 93.200 ;
        RECT 45.065 92.815 45.545 93.155 ;
        RECT 45.715 92.645 45.970 93.190 ;
        RECT 46.140 92.815 46.415 93.515 ;
        RECT 49.990 93.080 50.340 94.330 ;
        RECT 52.105 93.905 53.315 94.425 ;
        RECT 55.325 94.415 55.550 94.455 ;
        RECT 53.485 93.735 54.695 94.255 ;
        RECT 46.585 92.645 51.930 93.080 ;
        RECT 52.105 92.645 54.695 93.735 ;
        RECT 55.325 93.835 55.495 94.415 ;
        RECT 56.215 94.285 56.415 94.455 ;
        RECT 57.290 94.285 57.460 94.745 ;
        RECT 55.665 93.955 56.415 94.285 ;
        RECT 56.585 93.955 57.460 94.285 ;
        RECT 55.325 93.785 55.540 93.835 ;
        RECT 55.325 93.705 55.715 93.785 ;
        RECT 55.385 92.860 55.715 93.705 ;
        RECT 56.225 93.750 56.415 93.955 ;
        RECT 55.885 92.645 56.055 93.655 ;
        RECT 56.225 93.375 57.120 93.750 ;
        RECT 56.225 92.815 56.565 93.375 ;
        RECT 56.795 92.645 57.110 93.145 ;
        RECT 57.290 93.115 57.460 93.955 ;
        RECT 57.630 94.245 58.095 94.575 ;
        RECT 58.480 94.515 58.650 94.745 ;
        RECT 58.830 94.695 59.200 95.195 ;
        RECT 59.520 94.745 60.195 94.915 ;
        RECT 60.390 94.745 60.725 94.915 ;
        RECT 57.630 93.285 57.950 94.245 ;
        RECT 58.480 94.215 59.310 94.515 ;
        RECT 58.120 93.315 58.310 94.035 ;
        RECT 58.480 93.145 58.650 94.215 ;
        RECT 59.110 94.185 59.310 94.215 ;
        RECT 58.820 93.965 58.990 94.035 ;
        RECT 59.520 93.965 59.690 94.745 ;
        RECT 60.555 94.605 60.725 94.745 ;
        RECT 60.895 94.735 61.145 95.195 ;
        RECT 58.820 93.795 59.690 93.965 ;
        RECT 59.860 94.325 60.385 94.545 ;
        RECT 60.555 94.475 60.780 94.605 ;
        RECT 58.820 93.705 59.330 93.795 ;
        RECT 57.290 92.945 58.175 93.115 ;
        RECT 58.400 92.815 58.650 93.145 ;
        RECT 58.820 92.645 58.990 93.445 ;
        RECT 59.160 93.090 59.330 93.705 ;
        RECT 59.860 93.625 60.030 94.325 ;
        RECT 59.500 93.260 60.030 93.625 ;
        RECT 60.200 93.560 60.440 94.155 ;
        RECT 60.610 93.370 60.780 94.475 ;
        RECT 60.950 93.615 61.230 94.565 ;
        RECT 60.475 93.240 60.780 93.370 ;
        RECT 59.160 92.920 60.265 93.090 ;
        RECT 60.475 92.815 60.725 93.240 ;
        RECT 60.895 92.645 61.160 93.105 ;
        RECT 61.400 92.815 61.585 94.935 ;
        RECT 61.755 94.815 62.085 95.195 ;
        RECT 62.255 94.645 62.425 94.935 ;
        RECT 61.760 94.475 62.425 94.645 ;
        RECT 61.760 93.485 61.990 94.475 ;
        RECT 62.685 94.425 64.355 95.195 ;
        RECT 64.985 94.470 65.275 95.195 ;
        RECT 65.445 94.695 65.705 95.025 ;
        RECT 65.875 94.835 66.205 95.195 ;
        RECT 66.460 94.815 67.760 95.025 ;
        RECT 65.445 94.685 65.675 94.695 ;
        RECT 62.160 93.655 62.510 94.305 ;
        RECT 62.685 93.905 63.435 94.425 ;
        RECT 63.605 93.735 64.355 94.255 ;
        RECT 61.760 93.315 62.425 93.485 ;
        RECT 61.755 92.645 62.085 93.145 ;
        RECT 62.255 92.815 62.425 93.315 ;
        RECT 62.685 92.645 64.355 93.735 ;
        RECT 64.985 92.645 65.275 93.810 ;
        RECT 65.445 93.495 65.615 94.685 ;
        RECT 66.460 94.665 66.630 94.815 ;
        RECT 65.875 94.540 66.630 94.665 ;
        RECT 65.785 94.495 66.630 94.540 ;
        RECT 65.785 94.375 66.055 94.495 ;
        RECT 65.785 93.800 65.955 94.375 ;
        RECT 66.185 93.935 66.595 94.240 ;
        RECT 66.885 94.205 67.095 94.605 ;
        RECT 66.765 93.995 67.095 94.205 ;
        RECT 67.340 94.205 67.560 94.605 ;
        RECT 68.035 94.430 68.490 95.195 ;
        RECT 67.340 93.995 67.815 94.205 ;
        RECT 68.005 94.005 68.495 94.205 ;
        RECT 65.785 93.765 65.985 93.800 ;
        RECT 67.315 93.765 68.490 93.825 ;
        RECT 65.785 93.655 68.490 93.765 ;
        RECT 65.845 93.595 67.645 93.655 ;
        RECT 67.315 93.565 67.645 93.595 ;
        RECT 65.445 92.815 65.705 93.495 ;
        RECT 65.875 92.645 66.125 93.425 ;
        RECT 66.375 93.395 67.210 93.405 ;
        RECT 67.800 93.395 67.985 93.485 ;
        RECT 66.375 93.195 67.985 93.395 ;
        RECT 66.375 92.815 66.625 93.195 ;
        RECT 67.755 93.155 67.985 93.195 ;
        RECT 68.235 93.035 68.490 93.655 ;
        RECT 66.795 92.645 67.150 93.025 ;
        RECT 68.155 92.815 68.490 93.035 ;
        RECT 69.130 93.595 69.465 95.015 ;
        RECT 69.645 94.825 70.390 95.195 ;
        RECT 70.955 94.655 71.210 95.015 ;
        RECT 71.390 94.825 71.720 95.195 ;
        RECT 71.900 94.655 72.125 95.015 ;
        RECT 69.640 94.465 72.125 94.655 ;
        RECT 69.640 93.775 69.865 94.465 ;
        RECT 72.345 94.425 74.015 95.195 ;
        RECT 74.200 94.625 74.455 94.975 ;
        RECT 74.625 94.795 74.955 95.195 ;
        RECT 75.125 94.625 75.295 94.975 ;
        RECT 75.465 94.795 75.845 95.195 ;
        RECT 74.200 94.455 75.865 94.625 ;
        RECT 76.035 94.520 76.310 94.865 ;
        RECT 76.650 94.685 76.890 95.195 ;
        RECT 77.070 94.685 77.350 95.015 ;
        RECT 77.580 94.685 77.795 95.195 ;
        RECT 70.065 93.955 70.345 94.285 ;
        RECT 70.525 93.955 71.100 94.285 ;
        RECT 71.280 93.955 71.715 94.285 ;
        RECT 71.895 93.955 72.165 94.285 ;
        RECT 72.345 93.905 73.095 94.425 ;
        RECT 75.695 94.285 75.865 94.455 ;
        RECT 69.640 93.595 72.135 93.775 ;
        RECT 73.265 93.735 74.015 94.255 ;
        RECT 74.185 93.955 74.530 94.285 ;
        RECT 74.700 93.955 75.525 94.285 ;
        RECT 75.695 93.955 75.970 94.285 ;
        RECT 69.130 92.825 69.395 93.595 ;
        RECT 69.565 92.645 69.895 93.365 ;
        RECT 70.085 93.185 71.275 93.415 ;
        RECT 70.085 92.825 70.345 93.185 ;
        RECT 70.515 92.645 70.845 93.015 ;
        RECT 71.015 92.825 71.275 93.185 ;
        RECT 71.845 92.825 72.135 93.595 ;
        RECT 72.345 92.645 74.015 93.735 ;
        RECT 74.205 93.495 74.530 93.785 ;
        RECT 74.700 93.665 74.895 93.955 ;
        RECT 75.695 93.785 75.865 93.955 ;
        RECT 76.140 93.785 76.310 94.520 ;
        RECT 76.545 93.955 76.900 94.515 ;
        RECT 77.070 93.785 77.240 94.685 ;
        RECT 77.410 93.955 77.675 94.515 ;
        RECT 77.965 94.455 78.580 95.025 ;
        RECT 77.925 93.785 78.095 94.285 ;
        RECT 75.205 93.615 75.865 93.785 ;
        RECT 75.205 93.495 75.375 93.615 ;
        RECT 74.205 93.325 75.375 93.495 ;
        RECT 74.185 92.865 75.375 93.155 ;
        RECT 75.545 92.645 75.825 93.445 ;
        RECT 76.035 92.815 76.310 93.785 ;
        RECT 76.670 93.615 78.095 93.785 ;
        RECT 76.670 93.440 77.060 93.615 ;
        RECT 77.545 92.645 77.875 93.445 ;
        RECT 78.265 93.435 78.580 94.455 ;
        RECT 79.710 94.430 80.165 95.195 ;
        RECT 80.440 94.815 81.740 95.025 ;
        RECT 81.995 94.835 82.325 95.195 ;
        RECT 81.570 94.665 81.740 94.815 ;
        RECT 82.495 94.695 82.755 95.025 ;
        RECT 82.525 94.685 82.755 94.695 ;
        RECT 80.640 94.205 80.860 94.605 ;
        RECT 79.705 94.005 80.195 94.205 ;
        RECT 80.385 93.995 80.860 94.205 ;
        RECT 81.105 94.205 81.315 94.605 ;
        RECT 81.570 94.540 82.325 94.665 ;
        RECT 81.570 94.495 82.415 94.540 ;
        RECT 82.145 94.375 82.415 94.495 ;
        RECT 81.105 93.995 81.435 94.205 ;
        RECT 81.605 93.935 82.015 94.240 ;
        RECT 78.045 92.815 78.580 93.435 ;
        RECT 79.710 93.765 80.885 93.825 ;
        RECT 82.245 93.800 82.415 94.375 ;
        RECT 82.215 93.765 82.415 93.800 ;
        RECT 79.710 93.655 82.415 93.765 ;
        RECT 79.710 93.035 79.965 93.655 ;
        RECT 80.555 93.595 82.355 93.655 ;
        RECT 80.555 93.565 80.885 93.595 ;
        RECT 82.585 93.495 82.755 94.685 ;
        RECT 82.925 94.650 88.270 95.195 ;
        RECT 84.510 93.820 84.850 94.650 ;
        RECT 88.445 94.425 90.115 95.195 ;
        RECT 90.745 94.445 91.955 95.195 ;
        RECT 80.215 93.395 80.400 93.485 ;
        RECT 80.990 93.395 81.825 93.405 ;
        RECT 80.215 93.195 81.825 93.395 ;
        RECT 80.215 93.155 80.445 93.195 ;
        RECT 79.710 92.815 80.045 93.035 ;
        RECT 81.050 92.645 81.405 93.025 ;
        RECT 81.575 92.815 81.825 93.195 ;
        RECT 82.075 92.645 82.325 93.425 ;
        RECT 82.495 92.815 82.755 93.495 ;
        RECT 86.330 93.080 86.680 94.330 ;
        RECT 88.445 93.905 89.195 94.425 ;
        RECT 89.365 93.735 90.115 94.255 ;
        RECT 82.925 92.645 88.270 93.080 ;
        RECT 88.445 92.645 90.115 93.735 ;
        RECT 90.745 93.735 91.265 94.275 ;
        RECT 91.435 93.905 91.955 94.445 ;
        RECT 90.745 92.645 91.955 93.735 ;
        RECT 99.980 93.085 100.150 100.195 ;
        RECT 100.550 93.815 100.720 99.855 ;
        RECT 100.990 93.815 101.160 99.855 ;
        RECT 100.690 93.430 101.020 93.600 ;
        RECT 101.560 93.085 101.730 100.195 ;
        RECT 102.130 93.815 102.300 99.855 ;
        RECT 102.570 93.815 102.740 99.855 ;
        RECT 102.270 93.430 102.600 93.600 ;
        RECT 103.140 93.085 103.310 100.195 ;
        RECT 103.710 93.815 103.880 99.855 ;
        RECT 104.150 93.815 104.320 99.855 ;
        RECT 103.850 93.430 104.180 93.600 ;
        RECT 104.720 93.085 104.890 100.195 ;
        RECT 105.290 93.815 105.460 99.855 ;
        RECT 105.730 93.815 105.900 99.855 ;
        RECT 105.430 93.430 105.760 93.600 ;
        RECT 106.300 93.085 106.470 100.195 ;
        RECT 106.870 93.815 107.040 99.855 ;
        RECT 107.310 93.815 107.480 99.855 ;
        RECT 107.010 93.430 107.340 93.600 ;
        RECT 107.880 93.085 108.050 100.195 ;
        RECT 108.450 93.815 108.620 99.855 ;
        RECT 108.890 93.815 109.060 99.855 ;
        RECT 108.590 93.430 108.920 93.600 ;
        RECT 109.460 93.085 109.630 100.195 ;
        RECT 110.030 93.815 110.200 99.855 ;
        RECT 110.470 93.815 110.640 99.855 ;
        RECT 110.170 93.430 110.500 93.600 ;
        RECT 111.040 93.085 111.210 100.195 ;
        RECT 111.610 93.815 111.780 99.855 ;
        RECT 112.050 93.815 112.220 99.855 ;
        RECT 111.750 93.430 112.080 93.600 ;
        RECT 112.620 93.085 112.790 100.195 ;
        RECT 134.450 96.750 134.620 101.720 ;
        RECT 135.100 99.930 135.450 102.090 ;
        RECT 135.100 97.230 135.450 99.390 ;
        RECT 135.930 96.750 136.100 102.570 ;
        RECT 136.580 99.930 136.930 102.090 ;
        RECT 136.580 97.230 136.930 99.390 ;
        RECT 137.410 96.750 137.580 102.570 ;
        RECT 138.060 99.930 138.410 102.090 ;
        RECT 138.060 97.230 138.410 99.390 ;
        RECT 138.890 96.750 139.060 102.570 ;
        RECT 139.540 99.930 139.890 102.090 ;
        RECT 139.540 97.230 139.890 99.390 ;
        RECT 140.370 96.750 140.540 102.570 ;
        RECT 141.020 99.930 141.370 102.090 ;
        RECT 141.020 97.230 141.370 99.390 ;
        RECT 141.850 96.750 142.020 102.570 ;
        RECT 142.500 99.930 142.850 102.090 ;
        RECT 142.500 97.230 142.850 99.390 ;
        RECT 143.330 96.750 143.500 102.570 ;
        RECT 143.980 99.930 144.330 102.090 ;
        RECT 143.980 97.230 144.330 99.390 ;
        RECT 144.810 96.750 144.980 102.570 ;
        RECT 145.460 99.930 145.810 102.090 ;
        RECT 145.460 97.230 145.810 99.390 ;
        RECT 146.290 96.750 146.460 102.570 ;
        RECT 146.940 99.930 147.290 102.090 ;
        RECT 146.940 97.230 147.290 99.390 ;
        RECT 147.770 96.750 147.940 102.570 ;
        RECT 148.420 99.930 148.770 102.090 ;
        RECT 148.420 97.230 148.770 99.390 ;
        RECT 149.250 96.750 149.420 102.570 ;
        RECT 149.900 99.930 150.250 102.090 ;
        RECT 149.900 97.230 150.250 99.390 ;
        RECT 150.730 96.750 150.900 102.570 ;
        RECT 151.380 99.930 151.730 102.090 ;
        RECT 151.380 97.230 151.730 99.390 ;
        RECT 152.210 96.750 152.380 102.570 ;
        RECT 152.860 99.930 153.210 102.090 ;
        RECT 152.860 97.230 153.210 99.390 ;
        RECT 153.690 96.750 153.860 102.570 ;
        RECT 154.340 99.930 154.690 102.090 ;
        RECT 154.340 97.230 154.690 99.390 ;
        RECT 155.170 96.750 155.340 102.570 ;
        RECT 155.820 99.930 156.170 102.090 ;
        RECT 155.820 97.230 156.170 99.390 ;
        RECT 156.650 96.750 156.820 102.570 ;
        RECT 157.300 99.930 157.650 102.090 ;
        RECT 157.300 97.230 157.650 99.390 ;
        RECT 158.130 96.750 158.300 102.570 ;
        RECT 134.450 96.580 158.300 96.750 ;
        RECT 99.980 92.915 112.790 93.085 ;
        RECT 117.630 93.120 130.430 93.230 ;
        RECT 13.380 92.475 92.040 92.645 ;
        RECT 13.465 91.385 14.675 92.475 ;
        RECT 14.935 91.805 15.105 92.305 ;
        RECT 15.275 91.975 15.605 92.475 ;
        RECT 14.935 91.635 15.600 91.805 ;
        RECT 13.465 90.675 13.985 91.215 ;
        RECT 14.155 90.845 14.675 91.385 ;
        RECT 14.850 90.815 15.200 91.465 ;
        RECT 13.465 89.925 14.675 90.675 ;
        RECT 15.370 90.645 15.600 91.635 ;
        RECT 14.935 90.475 15.600 90.645 ;
        RECT 14.935 90.185 15.105 90.475 ;
        RECT 15.275 89.925 15.605 90.305 ;
        RECT 15.775 90.185 15.960 92.305 ;
        RECT 16.200 92.015 16.465 92.475 ;
        RECT 16.635 91.880 16.885 92.305 ;
        RECT 17.095 92.030 18.200 92.200 ;
        RECT 16.580 91.750 16.885 91.880 ;
        RECT 16.130 90.555 16.410 91.505 ;
        RECT 16.580 90.645 16.750 91.750 ;
        RECT 16.920 90.965 17.160 91.560 ;
        RECT 17.330 91.495 17.860 91.860 ;
        RECT 17.330 90.795 17.500 91.495 ;
        RECT 18.030 91.415 18.200 92.030 ;
        RECT 18.370 91.675 18.540 92.475 ;
        RECT 18.710 91.975 18.960 92.305 ;
        RECT 19.185 92.005 20.070 92.175 ;
        RECT 18.030 91.325 18.540 91.415 ;
        RECT 16.580 90.515 16.805 90.645 ;
        RECT 16.975 90.575 17.500 90.795 ;
        RECT 17.670 91.155 18.540 91.325 ;
        RECT 16.215 89.925 16.465 90.385 ;
        RECT 16.635 90.375 16.805 90.515 ;
        RECT 17.670 90.375 17.840 91.155 ;
        RECT 18.370 91.085 18.540 91.155 ;
        RECT 18.050 90.905 18.250 90.935 ;
        RECT 18.710 90.905 18.880 91.975 ;
        RECT 19.050 91.085 19.240 91.805 ;
        RECT 18.050 90.605 18.880 90.905 ;
        RECT 19.410 90.875 19.730 91.835 ;
        RECT 16.635 90.205 16.970 90.375 ;
        RECT 17.165 90.205 17.840 90.375 ;
        RECT 18.160 89.925 18.530 90.425 ;
        RECT 18.710 90.375 18.880 90.605 ;
        RECT 19.265 90.545 19.730 90.875 ;
        RECT 19.900 91.165 20.070 92.005 ;
        RECT 20.250 91.975 20.565 92.475 ;
        RECT 20.795 91.745 21.135 92.305 ;
        RECT 20.240 91.370 21.135 91.745 ;
        RECT 21.305 91.465 21.475 92.475 ;
        RECT 20.945 91.165 21.135 91.370 ;
        RECT 21.645 91.415 21.975 92.260 ;
        RECT 22.145 91.560 22.315 92.475 ;
        RECT 23.585 91.920 24.190 92.475 ;
        RECT 24.365 91.965 24.845 92.305 ;
        RECT 25.015 91.930 25.270 92.475 ;
        RECT 23.585 91.820 24.200 91.920 ;
        RECT 24.015 91.795 24.200 91.820 ;
        RECT 21.645 91.335 22.035 91.415 ;
        RECT 21.820 91.285 22.035 91.335 ;
        RECT 19.900 90.835 20.775 91.165 ;
        RECT 20.945 90.835 21.695 91.165 ;
        RECT 19.900 90.375 20.070 90.835 ;
        RECT 20.945 90.665 21.145 90.835 ;
        RECT 21.865 90.705 22.035 91.285 ;
        RECT 23.585 91.200 23.845 91.650 ;
        RECT 24.015 91.550 24.345 91.795 ;
        RECT 24.515 91.475 25.270 91.725 ;
        RECT 25.440 91.605 25.715 92.305 ;
        RECT 24.500 91.440 25.270 91.475 ;
        RECT 24.485 91.430 25.270 91.440 ;
        RECT 24.480 91.415 25.375 91.430 ;
        RECT 24.460 91.400 25.375 91.415 ;
        RECT 24.440 91.390 25.375 91.400 ;
        RECT 24.415 91.380 25.375 91.390 ;
        RECT 24.345 91.350 25.375 91.380 ;
        RECT 24.325 91.320 25.375 91.350 ;
        RECT 24.305 91.290 25.375 91.320 ;
        RECT 24.275 91.265 25.375 91.290 ;
        RECT 24.240 91.230 25.375 91.265 ;
        RECT 24.210 91.225 25.375 91.230 ;
        RECT 24.210 91.220 24.600 91.225 ;
        RECT 24.210 91.210 24.575 91.220 ;
        RECT 24.210 91.205 24.560 91.210 ;
        RECT 24.210 91.200 24.545 91.205 ;
        RECT 23.585 91.195 24.545 91.200 ;
        RECT 23.585 91.185 24.535 91.195 ;
        RECT 23.585 91.180 24.525 91.185 ;
        RECT 23.585 91.170 24.515 91.180 ;
        RECT 23.585 91.160 24.510 91.170 ;
        RECT 23.585 91.155 24.505 91.160 ;
        RECT 23.585 91.140 24.495 91.155 ;
        RECT 23.585 91.125 24.490 91.140 ;
        RECT 23.585 91.100 24.480 91.125 ;
        RECT 23.585 91.030 24.475 91.100 ;
        RECT 21.810 90.665 22.035 90.705 ;
        RECT 18.710 90.205 19.115 90.375 ;
        RECT 19.285 90.205 20.070 90.375 ;
        RECT 20.345 89.925 20.555 90.455 ;
        RECT 20.815 90.140 21.145 90.665 ;
        RECT 21.655 90.580 22.035 90.665 ;
        RECT 21.315 89.925 21.485 90.535 ;
        RECT 21.655 90.145 21.985 90.580 ;
        RECT 23.585 90.475 24.135 90.860 ;
        RECT 22.155 89.925 22.325 90.440 ;
        RECT 24.305 90.305 24.475 91.030 ;
        RECT 23.585 90.135 24.475 90.305 ;
        RECT 24.645 90.630 24.975 91.055 ;
        RECT 25.145 90.830 25.375 91.225 ;
        RECT 24.645 90.145 24.865 90.630 ;
        RECT 25.545 90.575 25.715 91.605 ;
        RECT 26.345 91.310 26.635 92.475 ;
        RECT 27.270 91.335 27.605 92.305 ;
        RECT 27.775 91.335 27.945 92.475 ;
        RECT 28.115 92.135 30.145 92.305 ;
        RECT 27.270 90.665 27.440 91.335 ;
        RECT 28.115 91.165 28.285 92.135 ;
        RECT 27.610 90.835 27.865 91.165 ;
        RECT 28.090 90.835 28.285 91.165 ;
        RECT 28.455 91.795 29.580 91.965 ;
        RECT 27.695 90.665 27.865 90.835 ;
        RECT 28.455 90.665 28.625 91.795 ;
        RECT 25.035 89.925 25.285 90.465 ;
        RECT 25.455 90.095 25.715 90.575 ;
        RECT 26.345 89.925 26.635 90.650 ;
        RECT 27.270 90.095 27.525 90.665 ;
        RECT 27.695 90.495 28.625 90.665 ;
        RECT 28.795 91.455 29.805 91.625 ;
        RECT 28.795 90.655 28.965 91.455 ;
        RECT 29.170 90.775 29.445 91.255 ;
        RECT 29.165 90.605 29.445 90.775 ;
        RECT 28.450 90.460 28.625 90.495 ;
        RECT 27.695 89.925 28.025 90.325 ;
        RECT 28.450 90.095 28.980 90.460 ;
        RECT 29.170 90.095 29.445 90.605 ;
        RECT 29.615 90.095 29.805 91.455 ;
        RECT 29.975 91.470 30.145 92.135 ;
        RECT 30.315 91.715 30.485 92.475 ;
        RECT 30.720 91.715 31.235 92.125 ;
        RECT 31.405 92.040 36.750 92.475 ;
        RECT 29.975 91.280 30.725 91.470 ;
        RECT 30.895 90.905 31.235 91.715 ;
        RECT 30.005 90.735 31.235 90.905 ;
        RECT 29.985 89.925 30.495 90.460 ;
        RECT 30.715 90.130 30.960 90.735 ;
        RECT 32.990 90.470 33.330 91.300 ;
        RECT 34.810 90.790 35.160 92.040 ;
        RECT 36.925 91.385 40.435 92.475 ;
        RECT 40.720 91.845 41.005 92.305 ;
        RECT 41.175 92.015 41.445 92.475 ;
        RECT 40.720 91.625 41.675 91.845 ;
        RECT 36.925 90.695 38.575 91.215 ;
        RECT 38.745 90.865 40.435 91.385 ;
        RECT 40.605 90.895 41.295 91.455 ;
        RECT 41.465 90.725 41.675 91.625 ;
        RECT 31.405 89.925 36.750 90.470 ;
        RECT 36.925 89.925 40.435 90.695 ;
        RECT 40.720 90.555 41.675 90.725 ;
        RECT 41.845 91.455 42.245 92.305 ;
        RECT 42.435 91.845 42.715 92.305 ;
        RECT 43.235 92.015 43.560 92.475 ;
        RECT 42.435 91.625 43.560 91.845 ;
        RECT 41.845 90.895 42.940 91.455 ;
        RECT 43.110 91.165 43.560 91.625 ;
        RECT 43.730 91.335 44.115 92.305 ;
        RECT 44.285 91.385 45.955 92.475 ;
        RECT 46.585 91.400 46.925 92.475 ;
        RECT 47.110 91.965 49.160 92.255 ;
        RECT 40.720 90.095 41.005 90.555 ;
        RECT 41.175 89.925 41.445 90.385 ;
        RECT 41.845 90.095 42.245 90.895 ;
        RECT 43.110 90.835 43.665 91.165 ;
        RECT 43.110 90.725 43.560 90.835 ;
        RECT 42.435 90.555 43.560 90.725 ;
        RECT 43.835 90.665 44.115 91.335 ;
        RECT 42.435 90.095 42.715 90.555 ;
        RECT 43.235 89.925 43.560 90.385 ;
        RECT 43.730 90.095 44.115 90.665 ;
        RECT 44.285 90.695 45.035 91.215 ;
        RECT 45.205 90.865 45.955 91.385 ;
        RECT 47.095 91.165 47.335 91.760 ;
        RECT 47.530 91.625 49.160 91.795 ;
        RECT 49.330 91.675 49.610 92.475 ;
        RECT 47.530 91.335 47.850 91.625 ;
        RECT 48.990 91.505 49.160 91.625 ;
        RECT 44.285 89.925 45.955 90.695 ;
        RECT 46.585 90.595 46.925 91.165 ;
        RECT 47.095 90.835 47.750 91.165 ;
        RECT 48.020 90.835 48.760 91.455 ;
        RECT 48.990 91.335 49.650 91.505 ;
        RECT 49.820 91.335 50.095 92.305 ;
        RECT 50.265 91.385 51.935 92.475 ;
        RECT 49.480 91.165 49.650 91.335 ;
        RECT 48.930 90.835 49.310 91.165 ;
        RECT 49.480 90.835 49.755 91.165 ;
        RECT 46.585 89.925 46.925 90.425 ;
        RECT 47.095 90.145 47.340 90.835 ;
        RECT 49.480 90.665 49.650 90.835 ;
        RECT 48.065 90.495 49.650 90.665 ;
        RECT 49.925 90.600 50.095 91.335 ;
        RECT 47.535 89.925 47.865 90.425 ;
        RECT 48.065 90.145 48.235 90.495 ;
        RECT 48.410 89.925 48.740 90.325 ;
        RECT 48.910 90.145 49.080 90.495 ;
        RECT 49.250 89.925 49.630 90.325 ;
        RECT 49.820 90.255 50.095 90.600 ;
        RECT 50.265 90.695 51.015 91.215 ;
        RECT 51.185 90.865 51.935 91.385 ;
        RECT 52.105 91.310 52.395 92.475 ;
        RECT 52.565 92.040 57.910 92.475 ;
        RECT 58.085 92.040 63.430 92.475 ;
        RECT 50.265 89.925 51.935 90.695 ;
        RECT 52.105 89.925 52.395 90.650 ;
        RECT 54.150 90.470 54.490 91.300 ;
        RECT 55.970 90.790 56.320 92.040 ;
        RECT 59.670 90.470 60.010 91.300 ;
        RECT 61.490 90.790 61.840 92.040 ;
        RECT 63.605 91.385 67.115 92.475 ;
        RECT 67.390 91.675 67.645 92.475 ;
        RECT 67.815 91.505 68.145 92.305 ;
        RECT 68.315 91.675 68.485 92.475 ;
        RECT 68.655 91.505 68.985 92.305 ;
        RECT 63.605 90.695 65.255 91.215 ;
        RECT 65.425 90.865 67.115 91.385 ;
        RECT 67.285 91.335 68.985 91.505 ;
        RECT 69.155 91.335 69.415 92.475 ;
        RECT 69.585 91.385 71.255 92.475 ;
        RECT 71.425 91.920 72.030 92.475 ;
        RECT 72.205 91.965 72.685 92.305 ;
        RECT 72.855 91.930 73.110 92.475 ;
        RECT 71.425 91.820 72.040 91.920 ;
        RECT 71.855 91.795 72.040 91.820 ;
        RECT 67.285 90.745 67.565 91.335 ;
        RECT 67.735 90.915 68.485 91.165 ;
        RECT 68.655 90.915 69.415 91.165 ;
        RECT 52.565 89.925 57.910 90.470 ;
        RECT 58.085 89.925 63.430 90.470 ;
        RECT 63.605 89.925 67.115 90.695 ;
        RECT 67.285 90.495 68.145 90.745 ;
        RECT 68.315 90.555 69.415 90.725 ;
        RECT 67.395 90.305 67.725 90.325 ;
        RECT 68.315 90.305 68.565 90.555 ;
        RECT 67.395 90.095 68.565 90.305 ;
        RECT 68.735 89.925 68.905 90.385 ;
        RECT 69.075 90.095 69.415 90.555 ;
        RECT 69.585 90.695 70.335 91.215 ;
        RECT 70.505 90.865 71.255 91.385 ;
        RECT 71.425 91.200 71.685 91.650 ;
        RECT 71.855 91.550 72.185 91.795 ;
        RECT 72.355 91.475 73.110 91.725 ;
        RECT 73.280 91.605 73.555 92.305 ;
        RECT 72.340 91.440 73.110 91.475 ;
        RECT 72.325 91.430 73.110 91.440 ;
        RECT 72.320 91.415 73.215 91.430 ;
        RECT 72.300 91.400 73.215 91.415 ;
        RECT 72.280 91.390 73.215 91.400 ;
        RECT 72.255 91.380 73.215 91.390 ;
        RECT 72.185 91.350 73.215 91.380 ;
        RECT 72.165 91.320 73.215 91.350 ;
        RECT 72.145 91.290 73.215 91.320 ;
        RECT 72.115 91.265 73.215 91.290 ;
        RECT 72.080 91.230 73.215 91.265 ;
        RECT 72.050 91.225 73.215 91.230 ;
        RECT 72.050 91.220 72.440 91.225 ;
        RECT 72.050 91.210 72.415 91.220 ;
        RECT 72.050 91.205 72.400 91.210 ;
        RECT 72.050 91.200 72.385 91.205 ;
        RECT 71.425 91.195 72.385 91.200 ;
        RECT 71.425 91.185 72.375 91.195 ;
        RECT 71.425 91.180 72.365 91.185 ;
        RECT 71.425 91.170 72.355 91.180 ;
        RECT 71.425 91.160 72.350 91.170 ;
        RECT 71.425 91.155 72.345 91.160 ;
        RECT 71.425 91.140 72.335 91.155 ;
        RECT 71.425 91.125 72.330 91.140 ;
        RECT 71.425 91.100 72.320 91.125 ;
        RECT 71.425 91.030 72.315 91.100 ;
        RECT 69.585 89.925 71.255 90.695 ;
        RECT 71.425 90.475 71.975 90.860 ;
        RECT 72.145 90.305 72.315 91.030 ;
        RECT 71.425 90.135 72.315 90.305 ;
        RECT 72.485 90.630 72.815 91.055 ;
        RECT 72.985 90.830 73.215 91.225 ;
        RECT 72.485 90.145 72.705 90.630 ;
        RECT 73.385 90.575 73.555 91.605 ;
        RECT 73.725 91.385 77.235 92.475 ;
        RECT 72.875 89.925 73.125 90.465 ;
        RECT 73.295 90.095 73.555 90.575 ;
        RECT 73.725 90.695 75.375 91.215 ;
        RECT 75.545 90.865 77.235 91.385 ;
        RECT 77.865 91.310 78.155 92.475 ;
        RECT 78.330 91.505 78.605 92.305 ;
        RECT 78.775 91.675 79.105 92.475 ;
        RECT 79.275 92.135 80.415 92.305 ;
        RECT 79.275 91.505 79.445 92.135 ;
        RECT 78.330 91.295 79.445 91.505 ;
        RECT 79.615 91.505 79.945 91.965 ;
        RECT 80.115 91.675 80.415 92.135 ;
        RECT 79.615 91.455 80.375 91.505 ;
        RECT 79.615 91.285 80.395 91.455 ;
        RECT 80.685 91.335 80.895 92.475 ;
        RECT 81.065 91.325 81.395 92.305 ;
        RECT 81.565 91.335 81.795 92.475 ;
        RECT 82.005 91.385 85.515 92.475 ;
        RECT 85.685 91.385 86.895 92.475 ;
        RECT 78.330 90.915 79.050 91.115 ;
        RECT 79.220 90.915 79.990 91.115 ;
        RECT 80.160 90.745 80.375 91.285 ;
        RECT 73.725 89.925 77.235 90.695 ;
        RECT 77.865 89.925 78.155 90.650 ;
        RECT 78.330 89.925 78.605 90.745 ;
        RECT 78.775 90.575 80.375 90.745 ;
        RECT 78.775 90.565 79.945 90.575 ;
        RECT 78.775 90.095 79.105 90.565 ;
        RECT 79.275 89.925 79.445 90.395 ;
        RECT 79.615 90.095 79.945 90.565 ;
        RECT 80.115 89.925 80.405 90.395 ;
        RECT 80.685 89.925 80.895 90.745 ;
        RECT 81.065 90.725 81.315 91.325 ;
        RECT 81.485 90.915 81.815 91.165 ;
        RECT 81.065 90.095 81.395 90.725 ;
        RECT 81.565 89.925 81.795 90.745 ;
        RECT 82.005 90.695 83.655 91.215 ;
        RECT 83.825 90.865 85.515 91.385 ;
        RECT 82.005 89.925 85.515 90.695 ;
        RECT 85.685 90.675 86.205 91.215 ;
        RECT 86.375 90.845 86.895 91.385 ;
        RECT 87.065 91.335 87.450 92.305 ;
        RECT 87.620 92.015 87.945 92.475 ;
        RECT 88.465 91.845 88.745 92.305 ;
        RECT 87.620 91.625 88.745 91.845 ;
        RECT 85.685 89.925 86.895 90.675 ;
        RECT 87.065 90.665 87.345 91.335 ;
        RECT 87.620 91.165 88.070 91.625 ;
        RECT 88.935 91.455 89.335 92.305 ;
        RECT 89.735 92.015 90.005 92.475 ;
        RECT 90.175 91.845 90.460 92.305 ;
        RECT 87.515 90.835 88.070 91.165 ;
        RECT 88.240 90.895 89.335 91.455 ;
        RECT 87.620 90.725 88.070 90.835 ;
        RECT 87.065 90.095 87.450 90.665 ;
        RECT 87.620 90.555 88.745 90.725 ;
        RECT 87.620 89.925 87.945 90.385 ;
        RECT 88.465 90.095 88.745 90.555 ;
        RECT 88.935 90.095 89.335 90.895 ;
        RECT 89.505 91.625 90.460 91.845 ;
        RECT 89.505 90.725 89.715 91.625 ;
        RECT 89.885 90.895 90.575 91.455 ;
        RECT 90.745 91.385 91.955 92.475 ;
        RECT 117.630 92.430 130.440 93.120 ;
        RECT 117.590 92.260 130.440 92.430 ;
        RECT 99.990 91.675 112.800 91.845 ;
        RECT 90.745 90.845 91.265 91.385 ;
        RECT 89.505 90.555 90.460 90.725 ;
        RECT 91.435 90.675 91.955 91.215 ;
        RECT 89.735 89.925 90.005 90.385 ;
        RECT 90.175 90.095 90.460 90.555 ;
        RECT 90.745 89.925 91.955 90.675 ;
        RECT 13.380 89.755 92.040 89.925 ;
        RECT 13.465 89.005 14.675 89.755 ;
        RECT 13.465 88.465 13.985 89.005 ;
        RECT 14.845 88.985 16.515 89.755 ;
        RECT 17.150 89.080 17.425 89.425 ;
        RECT 17.615 89.355 17.995 89.755 ;
        RECT 18.165 89.185 18.335 89.535 ;
        RECT 18.505 89.355 18.835 89.755 ;
        RECT 19.005 89.185 19.260 89.535 ;
        RECT 14.155 88.295 14.675 88.835 ;
        RECT 14.845 88.465 15.595 88.985 ;
        RECT 15.765 88.295 16.515 88.815 ;
        RECT 13.465 87.205 14.675 88.295 ;
        RECT 14.845 87.205 16.515 88.295 ;
        RECT 17.150 88.345 17.320 89.080 ;
        RECT 17.595 89.015 19.260 89.185 ;
        RECT 19.535 89.205 19.705 89.495 ;
        RECT 19.875 89.375 20.205 89.755 ;
        RECT 19.535 89.035 20.200 89.205 ;
        RECT 17.595 88.845 17.765 89.015 ;
        RECT 17.490 88.515 17.765 88.845 ;
        RECT 17.935 88.515 18.760 88.845 ;
        RECT 18.930 88.515 19.275 88.845 ;
        RECT 17.595 88.345 17.765 88.515 ;
        RECT 17.150 87.375 17.425 88.345 ;
        RECT 17.595 88.175 18.255 88.345 ;
        RECT 18.565 88.225 18.760 88.515 ;
        RECT 18.085 88.055 18.255 88.175 ;
        RECT 18.930 88.055 19.255 88.345 ;
        RECT 19.450 88.215 19.800 88.865 ;
        RECT 17.635 87.205 17.915 88.005 ;
        RECT 18.085 87.885 19.255 88.055 ;
        RECT 19.970 88.045 20.200 89.035 ;
        RECT 19.535 87.875 20.200 88.045 ;
        RECT 18.085 87.425 19.275 87.715 ;
        RECT 19.535 87.375 19.705 87.875 ;
        RECT 19.875 87.205 20.205 87.705 ;
        RECT 20.375 87.375 20.560 89.495 ;
        RECT 20.815 89.295 21.065 89.755 ;
        RECT 21.235 89.305 21.570 89.475 ;
        RECT 21.765 89.305 22.440 89.475 ;
        RECT 21.235 89.165 21.405 89.305 ;
        RECT 20.730 88.175 21.010 89.125 ;
        RECT 21.180 89.035 21.405 89.165 ;
        RECT 21.180 87.930 21.350 89.035 ;
        RECT 21.575 88.885 22.100 89.105 ;
        RECT 21.520 88.120 21.760 88.715 ;
        RECT 21.930 88.185 22.100 88.885 ;
        RECT 22.270 88.525 22.440 89.305 ;
        RECT 22.760 89.255 23.130 89.755 ;
        RECT 23.310 89.305 23.715 89.475 ;
        RECT 23.885 89.305 24.670 89.475 ;
        RECT 23.310 89.075 23.480 89.305 ;
        RECT 22.650 88.775 23.480 89.075 ;
        RECT 23.865 88.805 24.330 89.135 ;
        RECT 22.650 88.745 22.850 88.775 ;
        RECT 22.970 88.525 23.140 88.595 ;
        RECT 22.270 88.355 23.140 88.525 ;
        RECT 22.630 88.265 23.140 88.355 ;
        RECT 21.180 87.800 21.485 87.930 ;
        RECT 21.930 87.820 22.460 88.185 ;
        RECT 20.800 87.205 21.065 87.665 ;
        RECT 21.235 87.375 21.485 87.800 ;
        RECT 22.630 87.650 22.800 88.265 ;
        RECT 21.695 87.480 22.800 87.650 ;
        RECT 22.970 87.205 23.140 88.005 ;
        RECT 23.310 87.705 23.480 88.775 ;
        RECT 23.650 87.875 23.840 88.595 ;
        RECT 24.010 87.845 24.330 88.805 ;
        RECT 24.500 88.845 24.670 89.305 ;
        RECT 24.945 89.225 25.155 89.755 ;
        RECT 25.415 89.015 25.745 89.540 ;
        RECT 25.915 89.145 26.085 89.755 ;
        RECT 26.255 89.100 26.585 89.535 ;
        RECT 26.805 89.375 27.695 89.545 ;
        RECT 26.255 89.015 26.635 89.100 ;
        RECT 25.545 88.845 25.745 89.015 ;
        RECT 26.410 88.975 26.635 89.015 ;
        RECT 24.500 88.515 25.375 88.845 ;
        RECT 25.545 88.515 26.295 88.845 ;
        RECT 23.310 87.375 23.560 87.705 ;
        RECT 24.500 87.675 24.670 88.515 ;
        RECT 25.545 88.310 25.735 88.515 ;
        RECT 26.465 88.395 26.635 88.975 ;
        RECT 26.805 88.820 27.355 89.205 ;
        RECT 27.525 88.650 27.695 89.375 ;
        RECT 26.420 88.345 26.635 88.395 ;
        RECT 24.840 87.935 25.735 88.310 ;
        RECT 26.245 88.265 26.635 88.345 ;
        RECT 26.805 88.580 27.695 88.650 ;
        RECT 27.865 89.050 28.085 89.535 ;
        RECT 28.255 89.215 28.505 89.755 ;
        RECT 28.675 89.105 28.935 89.585 ;
        RECT 27.865 88.625 28.195 89.050 ;
        RECT 26.805 88.555 27.700 88.580 ;
        RECT 26.805 88.540 27.710 88.555 ;
        RECT 26.805 88.525 27.715 88.540 ;
        RECT 26.805 88.520 27.725 88.525 ;
        RECT 26.805 88.510 27.730 88.520 ;
        RECT 26.805 88.500 27.735 88.510 ;
        RECT 26.805 88.495 27.745 88.500 ;
        RECT 26.805 88.485 27.755 88.495 ;
        RECT 26.805 88.480 27.765 88.485 ;
        RECT 23.785 87.505 24.670 87.675 ;
        RECT 24.850 87.205 25.165 87.705 ;
        RECT 25.395 87.375 25.735 87.935 ;
        RECT 25.905 87.205 26.075 88.215 ;
        RECT 26.245 87.420 26.575 88.265 ;
        RECT 26.805 88.030 27.065 88.480 ;
        RECT 27.430 88.475 27.765 88.480 ;
        RECT 27.430 88.470 27.780 88.475 ;
        RECT 27.430 88.460 27.795 88.470 ;
        RECT 27.430 88.455 27.820 88.460 ;
        RECT 28.365 88.455 28.595 88.850 ;
        RECT 27.430 88.450 28.595 88.455 ;
        RECT 27.460 88.415 28.595 88.450 ;
        RECT 27.495 88.390 28.595 88.415 ;
        RECT 27.525 88.360 28.595 88.390 ;
        RECT 27.545 88.330 28.595 88.360 ;
        RECT 27.565 88.300 28.595 88.330 ;
        RECT 27.635 88.290 28.595 88.300 ;
        RECT 27.660 88.280 28.595 88.290 ;
        RECT 27.680 88.265 28.595 88.280 ;
        RECT 27.700 88.250 28.595 88.265 ;
        RECT 27.705 88.240 28.490 88.250 ;
        RECT 27.720 88.205 28.490 88.240 ;
        RECT 27.235 87.885 27.565 88.130 ;
        RECT 27.735 87.955 28.490 88.205 ;
        RECT 28.765 88.075 28.935 89.105 ;
        RECT 29.105 88.985 31.695 89.755 ;
        RECT 31.955 89.205 32.125 89.495 ;
        RECT 32.295 89.375 32.625 89.755 ;
        RECT 31.955 89.035 32.620 89.205 ;
        RECT 29.105 88.465 30.315 88.985 ;
        RECT 30.485 88.295 31.695 88.815 ;
        RECT 27.235 87.860 27.420 87.885 ;
        RECT 26.805 87.760 27.420 87.860 ;
        RECT 26.805 87.205 27.410 87.760 ;
        RECT 27.585 87.375 28.065 87.715 ;
        RECT 28.235 87.205 28.490 87.750 ;
        RECT 28.660 87.375 28.935 88.075 ;
        RECT 29.105 87.205 31.695 88.295 ;
        RECT 31.870 88.215 32.220 88.865 ;
        RECT 32.390 88.045 32.620 89.035 ;
        RECT 31.955 87.875 32.620 88.045 ;
        RECT 31.955 87.375 32.125 87.875 ;
        RECT 32.295 87.205 32.625 87.705 ;
        RECT 32.795 87.375 32.980 89.495 ;
        RECT 33.235 89.295 33.485 89.755 ;
        RECT 33.655 89.305 33.990 89.475 ;
        RECT 34.185 89.305 34.860 89.475 ;
        RECT 33.655 89.165 33.825 89.305 ;
        RECT 33.150 88.175 33.430 89.125 ;
        RECT 33.600 89.035 33.825 89.165 ;
        RECT 33.600 87.930 33.770 89.035 ;
        RECT 33.995 88.885 34.520 89.105 ;
        RECT 33.940 88.120 34.180 88.715 ;
        RECT 34.350 88.185 34.520 88.885 ;
        RECT 34.690 88.525 34.860 89.305 ;
        RECT 35.180 89.255 35.550 89.755 ;
        RECT 35.730 89.305 36.135 89.475 ;
        RECT 36.305 89.305 37.090 89.475 ;
        RECT 35.730 89.075 35.900 89.305 ;
        RECT 35.070 88.775 35.900 89.075 ;
        RECT 36.285 88.805 36.750 89.135 ;
        RECT 35.070 88.745 35.270 88.775 ;
        RECT 35.390 88.525 35.560 88.595 ;
        RECT 34.690 88.355 35.560 88.525 ;
        RECT 35.050 88.265 35.560 88.355 ;
        RECT 33.600 87.800 33.905 87.930 ;
        RECT 34.350 87.820 34.880 88.185 ;
        RECT 33.220 87.205 33.485 87.665 ;
        RECT 33.655 87.375 33.905 87.800 ;
        RECT 35.050 87.650 35.220 88.265 ;
        RECT 34.115 87.480 35.220 87.650 ;
        RECT 35.390 87.205 35.560 88.005 ;
        RECT 35.730 87.705 35.900 88.775 ;
        RECT 36.070 87.875 36.260 88.595 ;
        RECT 36.430 87.845 36.750 88.805 ;
        RECT 36.920 88.845 37.090 89.305 ;
        RECT 37.365 89.225 37.575 89.755 ;
        RECT 37.835 89.015 38.165 89.540 ;
        RECT 38.335 89.145 38.505 89.755 ;
        RECT 38.675 89.100 39.005 89.535 ;
        RECT 38.675 89.015 39.055 89.100 ;
        RECT 39.225 89.030 39.515 89.755 ;
        RECT 37.965 88.845 38.165 89.015 ;
        RECT 38.830 88.975 39.055 89.015 ;
        RECT 36.920 88.515 37.795 88.845 ;
        RECT 37.965 88.515 38.715 88.845 ;
        RECT 35.730 87.375 35.980 87.705 ;
        RECT 36.920 87.675 37.090 88.515 ;
        RECT 37.965 88.310 38.155 88.515 ;
        RECT 38.885 88.395 39.055 88.975 ;
        RECT 38.840 88.345 39.055 88.395 ;
        RECT 39.690 89.015 39.945 89.585 ;
        RECT 40.115 89.355 40.445 89.755 ;
        RECT 40.870 89.220 41.400 89.585 ;
        RECT 41.590 89.415 41.865 89.585 ;
        RECT 41.585 89.245 41.865 89.415 ;
        RECT 40.870 89.185 41.045 89.220 ;
        RECT 40.115 89.015 41.045 89.185 ;
        RECT 37.260 87.935 38.155 88.310 ;
        RECT 38.665 88.265 39.055 88.345 ;
        RECT 36.205 87.505 37.090 87.675 ;
        RECT 37.270 87.205 37.585 87.705 ;
        RECT 37.815 87.375 38.155 87.935 ;
        RECT 38.325 87.205 38.495 88.215 ;
        RECT 38.665 87.420 38.995 88.265 ;
        RECT 39.225 87.205 39.515 88.370 ;
        RECT 39.690 88.345 39.860 89.015 ;
        RECT 40.115 88.845 40.285 89.015 ;
        RECT 40.030 88.515 40.285 88.845 ;
        RECT 40.510 88.515 40.705 88.845 ;
        RECT 39.690 87.375 40.025 88.345 ;
        RECT 40.195 87.205 40.365 88.345 ;
        RECT 40.535 87.545 40.705 88.515 ;
        RECT 40.875 87.885 41.045 89.015 ;
        RECT 41.215 88.225 41.385 89.025 ;
        RECT 41.590 88.425 41.865 89.245 ;
        RECT 42.035 88.225 42.225 89.585 ;
        RECT 42.405 89.220 42.915 89.755 ;
        RECT 43.135 88.945 43.380 89.550 ;
        RECT 43.825 88.985 45.495 89.755 ;
        RECT 42.425 88.775 43.655 88.945 ;
        RECT 41.215 88.055 42.225 88.225 ;
        RECT 42.395 88.210 43.145 88.400 ;
        RECT 40.875 87.715 42.000 87.885 ;
        RECT 42.395 87.545 42.565 88.210 ;
        RECT 43.315 87.965 43.655 88.775 ;
        RECT 43.825 88.465 44.575 88.985 ;
        RECT 45.665 88.955 46.005 89.585 ;
        RECT 46.175 88.955 46.425 89.755 ;
        RECT 46.615 89.105 46.945 89.585 ;
        RECT 47.115 89.295 47.340 89.755 ;
        RECT 47.510 89.105 47.840 89.585 ;
        RECT 44.745 88.295 45.495 88.815 ;
        RECT 40.535 87.375 42.565 87.545 ;
        RECT 42.735 87.205 42.905 87.965 ;
        RECT 43.140 87.555 43.655 87.965 ;
        RECT 43.825 87.205 45.495 88.295 ;
        RECT 45.665 88.345 45.840 88.955 ;
        RECT 46.615 88.935 47.840 89.105 ;
        RECT 48.470 88.975 48.970 89.585 ;
        RECT 49.345 89.105 49.605 89.585 ;
        RECT 49.775 89.295 50.105 89.755 ;
        RECT 50.295 89.115 50.495 89.535 ;
        RECT 46.010 88.595 46.705 88.765 ;
        RECT 46.535 88.345 46.705 88.595 ;
        RECT 46.880 88.565 47.300 88.765 ;
        RECT 47.470 88.565 47.800 88.765 ;
        RECT 47.970 88.565 48.300 88.765 ;
        RECT 48.470 88.345 48.640 88.975 ;
        RECT 48.825 88.515 49.175 88.765 ;
        RECT 45.665 87.375 46.005 88.345 ;
        RECT 46.175 87.205 46.345 88.345 ;
        RECT 46.535 88.175 48.970 88.345 ;
        RECT 46.615 87.205 46.865 88.005 ;
        RECT 47.510 87.375 47.840 88.175 ;
        RECT 48.140 87.205 48.470 88.005 ;
        RECT 48.640 87.375 48.970 88.175 ;
        RECT 49.345 88.075 49.515 89.105 ;
        RECT 49.685 88.415 49.915 88.845 ;
        RECT 50.085 88.595 50.495 89.115 ;
        RECT 50.665 89.270 51.455 89.535 ;
        RECT 50.665 88.415 50.920 89.270 ;
        RECT 51.635 88.935 51.965 89.355 ;
        RECT 52.135 88.935 52.395 89.755 ;
        RECT 52.585 89.065 52.825 89.585 ;
        RECT 52.995 89.260 53.390 89.755 ;
        RECT 53.955 89.425 54.125 89.570 ;
        RECT 53.750 89.230 54.125 89.425 ;
        RECT 51.635 88.845 51.885 88.935 ;
        RECT 51.090 88.595 51.885 88.845 ;
        RECT 49.685 88.245 51.475 88.415 ;
        RECT 49.345 87.375 49.620 88.075 ;
        RECT 49.790 87.950 50.505 88.245 ;
        RECT 50.725 87.885 51.055 88.075 ;
        RECT 49.830 87.205 50.045 87.750 ;
        RECT 50.215 87.375 50.690 87.715 ;
        RECT 50.860 87.710 51.055 87.885 ;
        RECT 51.225 87.880 51.475 88.245 ;
        RECT 50.860 87.205 51.475 87.710 ;
        RECT 51.715 87.375 51.885 88.595 ;
        RECT 52.055 87.885 52.395 88.765 ;
        RECT 52.585 88.260 52.760 89.065 ;
        RECT 53.750 88.895 53.920 89.230 ;
        RECT 54.405 89.185 54.645 89.560 ;
        RECT 54.815 89.250 55.150 89.755 ;
        RECT 54.405 89.035 54.625 89.185 ;
        RECT 52.935 88.535 53.920 88.895 ;
        RECT 54.090 88.705 54.625 89.035 ;
        RECT 52.935 88.515 54.220 88.535 ;
        RECT 53.360 88.365 54.220 88.515 ;
        RECT 52.135 87.205 52.395 87.715 ;
        RECT 52.585 87.475 52.890 88.260 ;
        RECT 53.065 87.885 53.760 88.195 ;
        RECT 53.070 87.205 53.755 87.675 ;
        RECT 53.935 87.420 54.220 88.365 ;
        RECT 54.390 88.055 54.625 88.705 ;
        RECT 54.795 88.225 55.095 89.075 ;
        RECT 55.325 88.985 56.995 89.755 ;
        RECT 57.255 89.205 57.425 89.495 ;
        RECT 57.595 89.375 57.925 89.755 ;
        RECT 57.255 89.035 57.920 89.205 ;
        RECT 55.325 88.465 56.075 88.985 ;
        RECT 56.245 88.295 56.995 88.815 ;
        RECT 54.390 87.825 55.065 88.055 ;
        RECT 54.395 87.205 54.725 87.655 ;
        RECT 54.895 87.395 55.065 87.825 ;
        RECT 55.325 87.205 56.995 88.295 ;
        RECT 57.170 88.215 57.520 88.865 ;
        RECT 57.690 88.045 57.920 89.035 ;
        RECT 57.255 87.875 57.920 88.045 ;
        RECT 57.255 87.375 57.425 87.875 ;
        RECT 57.595 87.205 57.925 87.705 ;
        RECT 58.095 87.375 58.280 89.495 ;
        RECT 58.535 89.295 58.785 89.755 ;
        RECT 58.955 89.305 59.290 89.475 ;
        RECT 59.485 89.305 60.160 89.475 ;
        RECT 58.955 89.165 59.125 89.305 ;
        RECT 58.450 88.175 58.730 89.125 ;
        RECT 58.900 89.035 59.125 89.165 ;
        RECT 58.900 87.930 59.070 89.035 ;
        RECT 59.295 88.885 59.820 89.105 ;
        RECT 59.240 88.120 59.480 88.715 ;
        RECT 59.650 88.185 59.820 88.885 ;
        RECT 59.990 88.525 60.160 89.305 ;
        RECT 60.480 89.255 60.850 89.755 ;
        RECT 61.030 89.305 61.435 89.475 ;
        RECT 61.605 89.305 62.390 89.475 ;
        RECT 61.030 89.075 61.200 89.305 ;
        RECT 60.370 88.775 61.200 89.075 ;
        RECT 61.585 88.805 62.050 89.135 ;
        RECT 60.370 88.745 60.570 88.775 ;
        RECT 60.690 88.525 60.860 88.595 ;
        RECT 59.990 88.355 60.860 88.525 ;
        RECT 60.350 88.265 60.860 88.355 ;
        RECT 58.900 87.800 59.205 87.930 ;
        RECT 59.650 87.820 60.180 88.185 ;
        RECT 58.520 87.205 58.785 87.665 ;
        RECT 58.955 87.375 59.205 87.800 ;
        RECT 60.350 87.650 60.520 88.265 ;
        RECT 59.415 87.480 60.520 87.650 ;
        RECT 60.690 87.205 60.860 88.005 ;
        RECT 61.030 87.705 61.200 88.775 ;
        RECT 61.370 87.875 61.560 88.595 ;
        RECT 61.730 87.845 62.050 88.805 ;
        RECT 62.220 88.845 62.390 89.305 ;
        RECT 62.665 89.225 62.875 89.755 ;
        RECT 63.135 89.015 63.465 89.540 ;
        RECT 63.635 89.145 63.805 89.755 ;
        RECT 63.975 89.100 64.305 89.535 ;
        RECT 63.975 89.015 64.355 89.100 ;
        RECT 64.985 89.030 65.275 89.755 ;
        RECT 65.450 89.280 65.785 89.540 ;
        RECT 65.955 89.355 66.285 89.755 ;
        RECT 66.455 89.355 68.070 89.525 ;
        RECT 63.265 88.845 63.465 89.015 ;
        RECT 64.130 88.975 64.355 89.015 ;
        RECT 62.220 88.515 63.095 88.845 ;
        RECT 63.265 88.515 64.015 88.845 ;
        RECT 61.030 87.375 61.280 87.705 ;
        RECT 62.220 87.675 62.390 88.515 ;
        RECT 63.265 88.310 63.455 88.515 ;
        RECT 64.185 88.395 64.355 88.975 ;
        RECT 64.140 88.345 64.355 88.395 ;
        RECT 62.560 87.935 63.455 88.310 ;
        RECT 63.965 88.265 64.355 88.345 ;
        RECT 61.505 87.505 62.390 87.675 ;
        RECT 62.570 87.205 62.885 87.705 ;
        RECT 63.115 87.375 63.455 87.935 ;
        RECT 63.625 87.205 63.795 88.215 ;
        RECT 63.965 87.420 64.295 88.265 ;
        RECT 64.985 87.205 65.275 88.370 ;
        RECT 65.450 87.925 65.705 89.280 ;
        RECT 66.455 89.185 66.625 89.355 ;
        RECT 66.065 89.015 66.625 89.185 ;
        RECT 66.065 88.845 66.235 89.015 ;
        RECT 65.930 88.515 66.235 88.845 ;
        RECT 66.430 88.735 66.680 88.845 ;
        RECT 66.890 88.735 67.160 89.175 ;
        RECT 67.350 89.075 67.640 89.175 ;
        RECT 67.345 88.905 67.640 89.075 ;
        RECT 66.425 88.565 66.680 88.735 ;
        RECT 66.885 88.565 67.160 88.735 ;
        RECT 66.430 88.515 66.680 88.565 ;
        RECT 66.890 88.515 67.160 88.565 ;
        RECT 67.350 88.515 67.640 88.905 ;
        RECT 67.810 88.515 68.230 89.180 ;
        RECT 68.615 89.035 68.945 89.755 ;
        RECT 70.050 89.250 70.385 89.755 ;
        RECT 70.555 89.185 70.795 89.560 ;
        RECT 71.075 89.425 71.245 89.570 ;
        RECT 71.075 89.230 71.450 89.425 ;
        RECT 71.810 89.260 72.205 89.755 ;
        RECT 68.540 88.735 68.890 88.845 ;
        RECT 68.540 88.565 68.895 88.735 ;
        RECT 68.540 88.515 68.890 88.565 ;
        RECT 66.065 88.345 66.235 88.515 ;
        RECT 66.065 88.175 68.435 88.345 ;
        RECT 68.685 88.225 68.890 88.515 ;
        RECT 70.105 88.225 70.405 89.075 ;
        RECT 70.575 89.035 70.795 89.185 ;
        RECT 70.575 88.705 71.110 89.035 ;
        RECT 71.280 88.895 71.450 89.230 ;
        RECT 72.375 89.065 72.615 89.585 ;
        RECT 65.450 87.415 65.785 87.925 ;
        RECT 66.035 87.205 66.365 88.005 ;
        RECT 66.610 87.795 68.035 87.965 ;
        RECT 66.610 87.375 66.895 87.795 ;
        RECT 67.150 87.205 67.480 87.625 ;
        RECT 67.705 87.545 68.035 87.795 ;
        RECT 68.265 87.715 68.435 88.175 ;
        RECT 70.575 88.055 70.810 88.705 ;
        RECT 71.280 88.535 72.265 88.895 ;
        RECT 68.695 87.545 68.865 88.045 ;
        RECT 67.705 87.375 68.865 87.545 ;
        RECT 70.135 87.825 70.810 88.055 ;
        RECT 70.980 88.515 72.265 88.535 ;
        RECT 70.980 88.365 71.840 88.515 ;
        RECT 70.135 87.395 70.305 87.825 ;
        RECT 70.475 87.205 70.805 87.655 ;
        RECT 70.980 87.420 71.265 88.365 ;
        RECT 72.440 88.260 72.615 89.065 ;
        RECT 72.810 89.225 73.100 89.575 ;
        RECT 73.295 89.395 73.625 89.755 ;
        RECT 73.795 89.225 74.025 89.530 ;
        RECT 72.810 89.055 74.025 89.225 ;
        RECT 74.215 89.415 74.385 89.450 ;
        RECT 74.215 89.245 74.415 89.415 ;
        RECT 74.215 88.885 74.385 89.245 ;
        RECT 72.870 88.735 73.130 88.845 ;
        RECT 72.865 88.565 73.130 88.735 ;
        RECT 72.870 88.515 73.130 88.565 ;
        RECT 73.310 88.515 73.695 88.845 ;
        RECT 73.865 88.715 74.385 88.885 ;
        RECT 74.645 88.985 77.235 89.755 ;
        RECT 77.870 88.990 78.325 89.755 ;
        RECT 78.600 89.375 79.900 89.585 ;
        RECT 80.155 89.395 80.485 89.755 ;
        RECT 79.730 89.225 79.900 89.375 ;
        RECT 80.655 89.255 80.915 89.585 ;
        RECT 71.440 87.885 72.135 88.195 ;
        RECT 71.445 87.205 72.130 87.675 ;
        RECT 72.310 87.475 72.615 88.260 ;
        RECT 72.810 87.205 73.130 88.345 ;
        RECT 73.310 87.465 73.505 88.515 ;
        RECT 73.865 88.335 74.035 88.715 ;
        RECT 73.685 88.055 74.035 88.335 ;
        RECT 74.225 88.185 74.470 88.545 ;
        RECT 74.645 88.465 75.855 88.985 ;
        RECT 76.025 88.295 77.235 88.815 ;
        RECT 78.800 88.765 79.020 89.165 ;
        RECT 77.865 88.565 78.355 88.765 ;
        RECT 78.545 88.555 79.020 88.765 ;
        RECT 79.265 88.765 79.475 89.165 ;
        RECT 79.730 89.100 80.485 89.225 ;
        RECT 79.730 89.055 80.575 89.100 ;
        RECT 80.305 88.935 80.575 89.055 ;
        RECT 79.265 88.555 79.595 88.765 ;
        RECT 79.765 88.495 80.175 88.800 ;
        RECT 73.685 87.375 74.015 88.055 ;
        RECT 74.215 87.205 74.470 88.005 ;
        RECT 74.645 87.205 77.235 88.295 ;
        RECT 77.870 88.325 79.045 88.385 ;
        RECT 80.405 88.360 80.575 88.935 ;
        RECT 80.375 88.325 80.575 88.360 ;
        RECT 77.870 88.215 80.575 88.325 ;
        RECT 77.870 87.595 78.125 88.215 ;
        RECT 78.715 88.155 80.515 88.215 ;
        RECT 78.715 88.125 79.045 88.155 ;
        RECT 80.745 88.055 80.915 89.255 ;
        RECT 81.635 89.205 81.805 89.495 ;
        RECT 81.975 89.375 82.305 89.755 ;
        RECT 81.635 89.035 82.300 89.205 ;
        RECT 81.550 88.215 81.900 88.865 ;
        RECT 78.375 87.955 78.560 88.045 ;
        RECT 79.150 87.955 79.985 87.965 ;
        RECT 78.375 87.755 79.985 87.955 ;
        RECT 78.375 87.715 78.605 87.755 ;
        RECT 77.870 87.375 78.205 87.595 ;
        RECT 79.210 87.205 79.565 87.585 ;
        RECT 79.735 87.375 79.985 87.755 ;
        RECT 80.235 87.205 80.485 87.985 ;
        RECT 80.655 87.375 80.915 88.055 ;
        RECT 82.070 88.045 82.300 89.035 ;
        RECT 81.635 87.875 82.300 88.045 ;
        RECT 81.635 87.375 81.805 87.875 ;
        RECT 81.975 87.205 82.305 87.705 ;
        RECT 82.475 87.375 82.660 89.495 ;
        RECT 82.915 89.295 83.165 89.755 ;
        RECT 83.335 89.305 83.670 89.475 ;
        RECT 83.865 89.305 84.540 89.475 ;
        RECT 83.335 89.165 83.505 89.305 ;
        RECT 82.830 88.175 83.110 89.125 ;
        RECT 83.280 89.035 83.505 89.165 ;
        RECT 83.280 87.930 83.450 89.035 ;
        RECT 83.675 88.885 84.200 89.105 ;
        RECT 83.620 88.120 83.860 88.715 ;
        RECT 84.030 88.185 84.200 88.885 ;
        RECT 84.370 88.525 84.540 89.305 ;
        RECT 84.860 89.255 85.230 89.755 ;
        RECT 85.410 89.305 85.815 89.475 ;
        RECT 85.985 89.305 86.770 89.475 ;
        RECT 85.410 89.075 85.580 89.305 ;
        RECT 84.750 88.775 85.580 89.075 ;
        RECT 85.965 88.805 86.430 89.135 ;
        RECT 84.750 88.745 84.950 88.775 ;
        RECT 85.070 88.525 85.240 88.595 ;
        RECT 84.370 88.355 85.240 88.525 ;
        RECT 84.730 88.265 85.240 88.355 ;
        RECT 83.280 87.800 83.585 87.930 ;
        RECT 84.030 87.820 84.560 88.185 ;
        RECT 82.900 87.205 83.165 87.665 ;
        RECT 83.335 87.375 83.585 87.800 ;
        RECT 84.730 87.650 84.900 88.265 ;
        RECT 83.795 87.480 84.900 87.650 ;
        RECT 85.070 87.205 85.240 88.005 ;
        RECT 85.410 87.705 85.580 88.775 ;
        RECT 85.750 87.875 85.940 88.595 ;
        RECT 86.110 87.845 86.430 88.805 ;
        RECT 86.600 88.845 86.770 89.305 ;
        RECT 87.045 89.225 87.255 89.755 ;
        RECT 87.515 89.015 87.845 89.540 ;
        RECT 88.015 89.145 88.185 89.755 ;
        RECT 88.355 89.100 88.685 89.535 ;
        RECT 88.995 89.205 89.165 89.585 ;
        RECT 89.380 89.375 89.710 89.755 ;
        RECT 88.355 89.015 88.735 89.100 ;
        RECT 88.995 89.035 89.710 89.205 ;
        RECT 87.645 88.845 87.845 89.015 ;
        RECT 88.510 88.975 88.735 89.015 ;
        RECT 86.600 88.515 87.475 88.845 ;
        RECT 87.645 88.515 88.395 88.845 ;
        RECT 85.410 87.375 85.660 87.705 ;
        RECT 86.600 87.675 86.770 88.515 ;
        RECT 87.645 88.310 87.835 88.515 ;
        RECT 88.565 88.395 88.735 88.975 ;
        RECT 88.905 88.485 89.260 88.855 ;
        RECT 89.540 88.845 89.710 89.035 ;
        RECT 89.880 89.010 90.135 89.585 ;
        RECT 89.540 88.515 89.795 88.845 ;
        RECT 88.520 88.345 88.735 88.395 ;
        RECT 86.940 87.935 87.835 88.310 ;
        RECT 88.345 88.265 88.735 88.345 ;
        RECT 89.540 88.305 89.710 88.515 ;
        RECT 85.885 87.505 86.770 87.675 ;
        RECT 86.950 87.205 87.265 87.705 ;
        RECT 87.495 87.375 87.835 87.935 ;
        RECT 88.005 87.205 88.175 88.215 ;
        RECT 88.345 87.420 88.675 88.265 ;
        RECT 88.995 88.135 89.710 88.305 ;
        RECT 89.965 88.280 90.135 89.010 ;
        RECT 90.310 88.915 90.570 89.755 ;
        RECT 90.745 89.005 91.955 89.755 ;
        RECT 88.995 87.375 89.165 88.135 ;
        RECT 89.380 87.205 89.710 87.965 ;
        RECT 89.880 87.375 90.135 88.280 ;
        RECT 90.310 87.205 90.570 88.355 ;
        RECT 90.745 88.295 91.265 88.835 ;
        RECT 91.435 88.465 91.955 89.005 ;
        RECT 99.990 88.605 100.160 91.675 ;
        RECT 100.700 91.165 101.030 91.335 ;
        RECT 100.560 88.955 100.730 90.995 ;
        RECT 101.000 88.955 101.170 90.995 ;
        RECT 101.570 88.605 101.740 91.675 ;
        RECT 102.280 91.165 102.610 91.335 ;
        RECT 102.140 88.955 102.310 90.995 ;
        RECT 102.580 88.955 102.750 90.995 ;
        RECT 103.150 88.605 103.320 91.675 ;
        RECT 103.860 91.165 104.190 91.335 ;
        RECT 103.720 88.955 103.890 90.995 ;
        RECT 104.160 88.955 104.330 90.995 ;
        RECT 104.730 88.605 104.900 91.675 ;
        RECT 105.440 91.165 105.770 91.335 ;
        RECT 105.300 88.955 105.470 90.995 ;
        RECT 105.740 88.955 105.910 90.995 ;
        RECT 106.310 88.605 106.480 91.675 ;
        RECT 107.020 91.165 107.350 91.335 ;
        RECT 106.880 88.955 107.050 90.995 ;
        RECT 107.320 88.955 107.490 90.995 ;
        RECT 107.890 88.605 108.060 91.675 ;
        RECT 108.600 91.165 108.930 91.335 ;
        RECT 108.460 88.955 108.630 90.995 ;
        RECT 108.900 88.955 109.070 90.995 ;
        RECT 109.470 88.605 109.640 91.675 ;
        RECT 110.180 91.165 110.510 91.335 ;
        RECT 110.040 88.955 110.210 90.995 ;
        RECT 110.480 88.955 110.650 90.995 ;
        RECT 111.050 88.605 111.220 91.675 ;
        RECT 111.760 91.165 112.090 91.335 ;
        RECT 111.620 88.955 111.790 90.995 ;
        RECT 112.060 88.955 112.230 90.995 ;
        RECT 112.630 88.605 112.800 91.675 ;
        RECT 99.990 88.415 112.800 88.605 ;
        RECT 90.745 87.205 91.955 88.295 ;
        RECT 100.070 87.785 112.760 88.415 ;
        RECT 99.990 87.615 113.480 87.785 ;
        RECT 13.380 87.035 92.040 87.205 ;
        RECT 13.465 85.945 14.675 87.035 ;
        RECT 14.845 85.945 18.355 87.035 ;
        RECT 18.525 85.945 19.735 87.035 ;
        RECT 13.465 85.235 13.985 85.775 ;
        RECT 14.155 85.405 14.675 85.945 ;
        RECT 14.845 85.255 16.495 85.775 ;
        RECT 16.665 85.425 18.355 85.945 ;
        RECT 13.465 84.485 14.675 85.235 ;
        RECT 14.845 84.485 18.355 85.255 ;
        RECT 18.525 85.235 19.045 85.775 ;
        RECT 19.215 85.405 19.735 85.945 ;
        RECT 20.090 86.065 20.480 86.240 ;
        RECT 20.965 86.235 21.295 87.035 ;
        RECT 21.465 86.245 22.000 86.865 ;
        RECT 20.090 85.895 21.515 86.065 ;
        RECT 18.525 84.485 19.735 85.235 ;
        RECT 19.965 85.165 20.320 85.725 ;
        RECT 20.490 84.995 20.660 85.895 ;
        RECT 20.830 85.165 21.095 85.725 ;
        RECT 21.345 85.395 21.515 85.895 ;
        RECT 21.685 85.225 22.000 86.245 ;
        RECT 20.070 84.485 20.310 84.995 ;
        RECT 20.490 84.665 20.770 84.995 ;
        RECT 21.000 84.485 21.215 84.995 ;
        RECT 21.385 84.655 22.000 85.225 ;
        RECT 22.205 86.315 22.665 86.865 ;
        RECT 22.855 86.315 23.185 87.035 ;
        RECT 22.205 84.945 22.455 86.315 ;
        RECT 23.385 86.145 23.685 86.695 ;
        RECT 23.855 86.365 24.135 87.035 ;
        RECT 22.745 85.975 23.685 86.145 ;
        RECT 22.745 85.725 22.915 85.975 ;
        RECT 24.055 85.725 24.320 86.085 ;
        RECT 25.005 85.895 25.235 87.035 ;
        RECT 25.405 85.885 25.735 86.865 ;
        RECT 25.905 85.895 26.115 87.035 ;
        RECT 22.625 85.395 22.915 85.725 ;
        RECT 23.085 85.475 23.425 85.725 ;
        RECT 23.645 85.475 24.320 85.725 ;
        RECT 24.985 85.475 25.315 85.725 ;
        RECT 22.745 85.305 22.915 85.395 ;
        RECT 22.745 85.115 24.135 85.305 ;
        RECT 22.205 84.655 22.765 84.945 ;
        RECT 22.935 84.485 23.185 84.945 ;
        RECT 23.805 84.755 24.135 85.115 ;
        RECT 25.005 84.485 25.235 85.305 ;
        RECT 25.485 85.285 25.735 85.885 ;
        RECT 26.345 85.870 26.635 87.035 ;
        RECT 27.815 86.365 27.985 86.865 ;
        RECT 28.155 86.535 28.485 87.035 ;
        RECT 27.815 86.195 28.480 86.365 ;
        RECT 27.730 85.375 28.080 86.025 ;
        RECT 25.405 84.655 25.735 85.285 ;
        RECT 25.905 84.485 26.115 85.305 ;
        RECT 26.345 84.485 26.635 85.210 ;
        RECT 28.250 85.205 28.480 86.195 ;
        RECT 27.815 85.035 28.480 85.205 ;
        RECT 27.815 84.745 27.985 85.035 ;
        RECT 28.155 84.485 28.485 84.865 ;
        RECT 28.655 84.745 28.840 86.865 ;
        RECT 29.080 86.575 29.345 87.035 ;
        RECT 29.515 86.440 29.765 86.865 ;
        RECT 29.975 86.590 31.080 86.760 ;
        RECT 29.460 86.310 29.765 86.440 ;
        RECT 29.010 85.115 29.290 86.065 ;
        RECT 29.460 85.205 29.630 86.310 ;
        RECT 29.800 85.525 30.040 86.120 ;
        RECT 30.210 86.055 30.740 86.420 ;
        RECT 30.210 85.355 30.380 86.055 ;
        RECT 30.910 85.975 31.080 86.590 ;
        RECT 31.250 86.235 31.420 87.035 ;
        RECT 31.590 86.535 31.840 86.865 ;
        RECT 32.065 86.565 32.950 86.735 ;
        RECT 30.910 85.885 31.420 85.975 ;
        RECT 29.460 85.075 29.685 85.205 ;
        RECT 29.855 85.135 30.380 85.355 ;
        RECT 30.550 85.715 31.420 85.885 ;
        RECT 29.095 84.485 29.345 84.945 ;
        RECT 29.515 84.935 29.685 85.075 ;
        RECT 30.550 84.935 30.720 85.715 ;
        RECT 31.250 85.645 31.420 85.715 ;
        RECT 30.930 85.465 31.130 85.495 ;
        RECT 31.590 85.465 31.760 86.535 ;
        RECT 31.930 85.645 32.120 86.365 ;
        RECT 30.930 85.165 31.760 85.465 ;
        RECT 32.290 85.435 32.610 86.395 ;
        RECT 29.515 84.765 29.850 84.935 ;
        RECT 30.045 84.765 30.720 84.935 ;
        RECT 31.040 84.485 31.410 84.985 ;
        RECT 31.590 84.935 31.760 85.165 ;
        RECT 32.145 85.105 32.610 85.435 ;
        RECT 32.780 85.725 32.950 86.565 ;
        RECT 33.130 86.535 33.445 87.035 ;
        RECT 33.675 86.305 34.015 86.865 ;
        RECT 33.120 85.930 34.015 86.305 ;
        RECT 34.185 86.025 34.355 87.035 ;
        RECT 33.825 85.725 34.015 85.930 ;
        RECT 34.525 85.975 34.855 86.820 ;
        RECT 35.025 86.120 35.195 87.035 ;
        RECT 34.525 85.895 34.915 85.975 ;
        RECT 35.545 85.945 39.055 87.035 ;
        RECT 34.700 85.845 34.915 85.895 ;
        RECT 32.780 85.395 33.655 85.725 ;
        RECT 33.825 85.395 34.575 85.725 ;
        RECT 32.780 84.935 32.950 85.395 ;
        RECT 33.825 85.225 34.025 85.395 ;
        RECT 34.745 85.265 34.915 85.845 ;
        RECT 34.690 85.225 34.915 85.265 ;
        RECT 31.590 84.765 31.995 84.935 ;
        RECT 32.165 84.765 32.950 84.935 ;
        RECT 33.225 84.485 33.435 85.015 ;
        RECT 33.695 84.700 34.025 85.225 ;
        RECT 34.535 85.140 34.915 85.225 ;
        RECT 35.545 85.255 37.195 85.775 ;
        RECT 37.365 85.425 39.055 85.945 ;
        RECT 40.145 85.895 40.530 86.865 ;
        RECT 40.700 86.575 41.025 87.035 ;
        RECT 41.545 86.405 41.825 86.865 ;
        RECT 40.700 86.185 41.825 86.405 ;
        RECT 34.195 84.485 34.365 85.095 ;
        RECT 34.535 84.705 34.865 85.140 ;
        RECT 35.035 84.485 35.205 85.000 ;
        RECT 35.545 84.485 39.055 85.255 ;
        RECT 40.145 85.225 40.425 85.895 ;
        RECT 40.700 85.725 41.150 86.185 ;
        RECT 42.015 86.015 42.415 86.865 ;
        RECT 42.815 86.575 43.085 87.035 ;
        RECT 43.255 86.405 43.540 86.865 ;
        RECT 43.825 86.525 44.085 87.035 ;
        RECT 40.595 85.395 41.150 85.725 ;
        RECT 41.320 85.455 42.415 86.015 ;
        RECT 40.700 85.285 41.150 85.395 ;
        RECT 40.145 84.655 40.530 85.225 ;
        RECT 40.700 85.115 41.825 85.285 ;
        RECT 40.700 84.485 41.025 84.945 ;
        RECT 41.545 84.655 41.825 85.115 ;
        RECT 42.015 84.655 42.415 85.455 ;
        RECT 42.585 86.185 43.540 86.405 ;
        RECT 42.585 85.285 42.795 86.185 ;
        RECT 42.965 85.455 43.655 86.015 ;
        RECT 43.825 85.475 44.165 86.355 ;
        RECT 44.335 85.645 44.505 86.865 ;
        RECT 44.745 86.530 45.360 87.035 ;
        RECT 44.745 85.995 44.995 86.360 ;
        RECT 45.165 86.355 45.360 86.530 ;
        RECT 45.530 86.525 46.005 86.865 ;
        RECT 46.175 86.490 46.390 87.035 ;
        RECT 45.165 86.165 45.495 86.355 ;
        RECT 45.715 85.995 46.430 86.290 ;
        RECT 46.600 86.165 46.875 86.865 ;
        RECT 44.745 85.825 46.535 85.995 ;
        RECT 44.335 85.395 45.130 85.645 ;
        RECT 44.335 85.305 44.585 85.395 ;
        RECT 42.585 85.115 43.540 85.285 ;
        RECT 42.815 84.485 43.085 84.945 ;
        RECT 43.255 84.655 43.540 85.115 ;
        RECT 43.825 84.485 44.085 85.305 ;
        RECT 44.255 84.885 44.585 85.305 ;
        RECT 45.300 84.970 45.555 85.825 ;
        RECT 44.765 84.705 45.555 84.970 ;
        RECT 45.725 85.125 46.135 85.645 ;
        RECT 46.305 85.395 46.535 85.825 ;
        RECT 46.705 85.135 46.875 86.165 ;
        RECT 45.725 84.705 45.925 85.125 ;
        RECT 46.115 84.485 46.445 84.945 ;
        RECT 46.615 84.655 46.875 85.135 ;
        RECT 47.985 85.980 48.290 86.765 ;
        RECT 48.470 86.565 49.155 87.035 ;
        RECT 48.465 86.045 49.160 86.355 ;
        RECT 47.985 85.175 48.160 85.980 ;
        RECT 49.335 85.875 49.620 86.820 ;
        RECT 49.795 86.585 50.125 87.035 ;
        RECT 50.295 86.415 50.465 86.845 ;
        RECT 48.760 85.725 49.620 85.875 ;
        RECT 48.335 85.705 49.620 85.725 ;
        RECT 49.790 86.185 50.465 86.415 ;
        RECT 48.335 85.345 49.320 85.705 ;
        RECT 49.790 85.535 50.025 86.185 ;
        RECT 47.985 84.655 48.225 85.175 ;
        RECT 49.150 85.010 49.320 85.345 ;
        RECT 49.490 85.205 50.025 85.535 ;
        RECT 49.805 85.055 50.025 85.205 ;
        RECT 50.195 85.165 50.495 86.015 ;
        RECT 50.725 85.945 51.935 87.035 ;
        RECT 50.725 85.235 51.245 85.775 ;
        RECT 51.415 85.405 51.935 85.945 ;
        RECT 52.105 85.870 52.395 87.035 ;
        RECT 52.570 85.895 52.905 86.865 ;
        RECT 53.075 85.895 53.245 87.035 ;
        RECT 53.415 86.695 55.445 86.865 ;
        RECT 48.395 84.485 48.790 84.980 ;
        RECT 49.150 84.815 49.525 85.010 ;
        RECT 49.355 84.670 49.525 84.815 ;
        RECT 49.805 84.680 50.045 85.055 ;
        RECT 50.215 84.485 50.550 84.990 ;
        RECT 50.725 84.485 51.935 85.235 ;
        RECT 52.570 85.225 52.740 85.895 ;
        RECT 53.415 85.725 53.585 86.695 ;
        RECT 52.910 85.395 53.165 85.725 ;
        RECT 53.390 85.395 53.585 85.725 ;
        RECT 53.755 86.355 54.880 86.525 ;
        RECT 52.995 85.225 53.165 85.395 ;
        RECT 53.755 85.225 53.925 86.355 ;
        RECT 52.105 84.485 52.395 85.210 ;
        RECT 52.570 84.655 52.825 85.225 ;
        RECT 52.995 85.055 53.925 85.225 ;
        RECT 54.095 86.015 55.105 86.185 ;
        RECT 54.095 85.215 54.265 86.015 ;
        RECT 53.750 85.020 53.925 85.055 ;
        RECT 52.995 84.485 53.325 84.885 ;
        RECT 53.750 84.655 54.280 85.020 ;
        RECT 54.470 84.995 54.745 85.815 ;
        RECT 54.465 84.825 54.745 84.995 ;
        RECT 54.470 84.655 54.745 84.825 ;
        RECT 54.915 84.655 55.105 86.015 ;
        RECT 55.275 86.030 55.445 86.695 ;
        RECT 55.615 86.275 55.785 87.035 ;
        RECT 56.020 86.275 56.535 86.685 ;
        RECT 55.275 85.840 56.025 86.030 ;
        RECT 56.195 85.465 56.535 86.275 ;
        RECT 57.255 86.365 57.425 86.865 ;
        RECT 57.595 86.535 57.925 87.035 ;
        RECT 57.255 86.195 57.920 86.365 ;
        RECT 55.305 85.295 56.535 85.465 ;
        RECT 57.170 85.375 57.520 86.025 ;
        RECT 55.285 84.485 55.795 85.020 ;
        RECT 56.015 84.690 56.260 85.295 ;
        RECT 57.690 85.205 57.920 86.195 ;
        RECT 57.255 85.035 57.920 85.205 ;
        RECT 57.255 84.745 57.425 85.035 ;
        RECT 57.595 84.485 57.925 84.865 ;
        RECT 58.095 84.745 58.280 86.865 ;
        RECT 58.520 86.575 58.785 87.035 ;
        RECT 58.955 86.440 59.205 86.865 ;
        RECT 59.415 86.590 60.520 86.760 ;
        RECT 58.900 86.310 59.205 86.440 ;
        RECT 58.450 85.115 58.730 86.065 ;
        RECT 58.900 85.205 59.070 86.310 ;
        RECT 59.240 85.525 59.480 86.120 ;
        RECT 59.650 86.055 60.180 86.420 ;
        RECT 59.650 85.355 59.820 86.055 ;
        RECT 60.350 85.975 60.520 86.590 ;
        RECT 60.690 86.235 60.860 87.035 ;
        RECT 61.030 86.535 61.280 86.865 ;
        RECT 61.505 86.565 62.390 86.735 ;
        RECT 60.350 85.885 60.860 85.975 ;
        RECT 58.900 85.075 59.125 85.205 ;
        RECT 59.295 85.135 59.820 85.355 ;
        RECT 59.990 85.715 60.860 85.885 ;
        RECT 58.535 84.485 58.785 84.945 ;
        RECT 58.955 84.935 59.125 85.075 ;
        RECT 59.990 84.935 60.160 85.715 ;
        RECT 60.690 85.645 60.860 85.715 ;
        RECT 60.370 85.465 60.570 85.495 ;
        RECT 61.030 85.465 61.200 86.535 ;
        RECT 61.370 85.645 61.560 86.365 ;
        RECT 60.370 85.165 61.200 85.465 ;
        RECT 61.730 85.435 62.050 86.395 ;
        RECT 58.955 84.765 59.290 84.935 ;
        RECT 59.485 84.765 60.160 84.935 ;
        RECT 60.480 84.485 60.850 84.985 ;
        RECT 61.030 84.935 61.200 85.165 ;
        RECT 61.585 85.105 62.050 85.435 ;
        RECT 62.220 85.725 62.390 86.565 ;
        RECT 62.570 86.535 62.885 87.035 ;
        RECT 63.115 86.305 63.455 86.865 ;
        RECT 62.560 85.930 63.455 86.305 ;
        RECT 63.625 86.025 63.795 87.035 ;
        RECT 63.265 85.725 63.455 85.930 ;
        RECT 63.965 85.975 64.295 86.820 ;
        RECT 64.530 86.085 64.795 86.855 ;
        RECT 64.965 86.315 65.295 87.035 ;
        RECT 65.485 86.495 65.745 86.855 ;
        RECT 65.915 86.665 66.245 87.035 ;
        RECT 66.415 86.495 66.675 86.855 ;
        RECT 65.485 86.265 66.675 86.495 ;
        RECT 67.245 86.085 67.535 86.855 ;
        RECT 63.965 85.895 64.355 85.975 ;
        RECT 64.140 85.845 64.355 85.895 ;
        RECT 62.220 85.395 63.095 85.725 ;
        RECT 63.265 85.395 64.015 85.725 ;
        RECT 62.220 84.935 62.390 85.395 ;
        RECT 63.265 85.225 63.465 85.395 ;
        RECT 64.185 85.265 64.355 85.845 ;
        RECT 64.130 85.225 64.355 85.265 ;
        RECT 61.030 84.765 61.435 84.935 ;
        RECT 61.605 84.765 62.390 84.935 ;
        RECT 62.665 84.485 62.875 85.015 ;
        RECT 63.135 84.700 63.465 85.225 ;
        RECT 63.975 85.140 64.355 85.225 ;
        RECT 63.635 84.485 63.805 85.095 ;
        RECT 63.975 84.705 64.305 85.140 ;
        RECT 64.530 84.665 64.865 86.085 ;
        RECT 65.040 85.905 67.535 86.085 ;
        RECT 67.780 86.245 68.315 86.865 ;
        RECT 65.040 85.215 65.265 85.905 ;
        RECT 65.465 85.395 65.745 85.725 ;
        RECT 65.925 85.395 66.500 85.725 ;
        RECT 66.680 85.395 67.115 85.725 ;
        RECT 67.295 85.395 67.565 85.725 ;
        RECT 67.780 85.225 68.095 86.245 ;
        RECT 68.485 86.235 68.815 87.035 ;
        RECT 69.300 86.065 69.690 86.240 ;
        RECT 68.265 85.895 69.690 86.065 ;
        RECT 70.045 85.895 70.305 87.035 ;
        RECT 68.265 85.395 68.435 85.895 ;
        RECT 65.040 85.025 67.525 85.215 ;
        RECT 65.045 84.485 65.790 84.855 ;
        RECT 66.355 84.665 66.610 85.025 ;
        RECT 66.790 84.485 67.120 84.855 ;
        RECT 67.300 84.665 67.525 85.025 ;
        RECT 67.780 84.655 68.395 85.225 ;
        RECT 68.685 85.165 68.950 85.725 ;
        RECT 69.120 84.995 69.290 85.895 ;
        RECT 70.475 85.885 70.805 86.865 ;
        RECT 70.975 85.895 71.255 87.035 ;
        RECT 71.425 85.945 72.635 87.035 ;
        RECT 69.460 85.165 69.815 85.725 ;
        RECT 70.065 85.475 70.400 85.725 ;
        RECT 70.570 85.285 70.740 85.885 ;
        RECT 70.910 85.455 71.245 85.725 ;
        RECT 68.565 84.485 68.780 84.995 ;
        RECT 69.010 84.665 69.290 84.995 ;
        RECT 69.470 84.485 69.710 84.995 ;
        RECT 70.045 84.655 70.740 85.285 ;
        RECT 70.945 84.485 71.255 85.285 ;
        RECT 71.425 85.235 71.945 85.775 ;
        RECT 72.115 85.405 72.635 85.945 ;
        RECT 72.810 85.895 73.130 87.035 ;
        RECT 73.310 85.725 73.505 86.775 ;
        RECT 73.685 86.185 74.015 86.865 ;
        RECT 74.215 86.235 74.470 87.035 ;
        RECT 73.685 85.905 74.035 86.185 ;
        RECT 75.750 86.065 76.140 86.240 ;
        RECT 76.625 86.235 76.955 87.035 ;
        RECT 77.125 86.245 77.660 86.865 ;
        RECT 72.870 85.675 73.130 85.725 ;
        RECT 72.865 85.505 73.130 85.675 ;
        RECT 72.870 85.395 73.130 85.505 ;
        RECT 73.310 85.395 73.695 85.725 ;
        RECT 73.865 85.525 74.035 85.905 ;
        RECT 74.225 85.695 74.470 86.055 ;
        RECT 75.750 85.895 77.175 86.065 ;
        RECT 73.865 85.355 74.385 85.525 ;
        RECT 71.425 84.485 72.635 85.235 ;
        RECT 72.810 85.015 74.025 85.185 ;
        RECT 72.810 84.665 73.100 85.015 ;
        RECT 73.295 84.485 73.625 84.845 ;
        RECT 73.795 84.710 74.025 85.015 ;
        RECT 74.215 84.995 74.385 85.355 ;
        RECT 75.625 85.165 75.980 85.725 ;
        RECT 76.150 84.995 76.320 85.895 ;
        RECT 76.490 85.165 76.755 85.725 ;
        RECT 77.005 85.395 77.175 85.895 ;
        RECT 77.345 85.225 77.660 86.245 ;
        RECT 77.865 85.870 78.155 87.035 ;
        RECT 78.480 86.025 78.780 86.865 ;
        RECT 78.975 86.195 79.225 87.035 ;
        RECT 79.815 86.445 80.620 86.865 ;
        RECT 79.395 86.275 80.960 86.445 ;
        RECT 79.395 86.025 79.565 86.275 ;
        RECT 78.480 85.855 79.565 86.025 ;
        RECT 78.325 85.395 78.655 85.685 ;
        RECT 78.825 85.225 78.995 85.855 ;
        RECT 79.735 85.725 80.055 86.105 ;
        RECT 80.245 86.015 80.620 86.105 ;
        RECT 80.225 85.845 80.620 86.015 ;
        RECT 80.790 86.025 80.960 86.275 ;
        RECT 81.130 86.195 81.460 87.035 ;
        RECT 81.630 86.275 82.295 86.865 ;
        RECT 80.790 85.855 81.710 86.025 ;
        RECT 79.165 85.475 79.495 85.685 ;
        RECT 79.675 85.475 80.055 85.725 ;
        RECT 80.245 85.685 80.620 85.845 ;
        RECT 81.540 85.685 81.710 85.855 ;
        RECT 80.245 85.475 80.730 85.685 ;
        RECT 80.920 85.475 81.370 85.685 ;
        RECT 81.540 85.475 81.875 85.685 ;
        RECT 82.045 85.305 82.295 86.275 ;
        RECT 74.215 84.825 74.415 84.995 ;
        RECT 74.215 84.790 74.385 84.825 ;
        RECT 75.730 84.485 75.970 84.995 ;
        RECT 76.150 84.665 76.430 84.995 ;
        RECT 76.660 84.485 76.875 84.995 ;
        RECT 77.045 84.655 77.660 85.225 ;
        RECT 77.865 84.485 78.155 85.210 ;
        RECT 78.485 85.045 78.995 85.225 ;
        RECT 79.400 85.135 81.100 85.305 ;
        RECT 79.400 85.045 79.785 85.135 ;
        RECT 78.485 84.655 78.815 85.045 ;
        RECT 78.985 84.705 80.170 84.875 ;
        RECT 80.430 84.485 80.600 84.955 ;
        RECT 80.770 84.670 81.100 85.135 ;
        RECT 81.270 84.485 81.440 85.305 ;
        RECT 81.610 84.665 82.295 85.305 ;
        RECT 83.390 85.895 83.725 86.865 ;
        RECT 83.895 85.895 84.065 87.035 ;
        RECT 84.235 86.695 86.265 86.865 ;
        RECT 83.390 85.225 83.560 85.895 ;
        RECT 84.235 85.725 84.405 86.695 ;
        RECT 83.730 85.395 83.985 85.725 ;
        RECT 84.210 85.395 84.405 85.725 ;
        RECT 84.575 86.355 85.700 86.525 ;
        RECT 83.815 85.225 83.985 85.395 ;
        RECT 84.575 85.225 84.745 86.355 ;
        RECT 83.390 84.655 83.645 85.225 ;
        RECT 83.815 85.055 84.745 85.225 ;
        RECT 84.915 86.015 85.925 86.185 ;
        RECT 84.915 85.215 85.085 86.015 ;
        RECT 85.290 85.675 85.565 85.815 ;
        RECT 85.285 85.505 85.565 85.675 ;
        RECT 84.570 85.020 84.745 85.055 ;
        RECT 83.815 84.485 84.145 84.885 ;
        RECT 84.570 84.655 85.100 85.020 ;
        RECT 85.290 84.655 85.565 85.505 ;
        RECT 85.735 84.655 85.925 86.015 ;
        RECT 86.095 86.030 86.265 86.695 ;
        RECT 86.435 86.275 86.605 87.035 ;
        RECT 86.840 86.275 87.355 86.685 ;
        RECT 86.095 85.840 86.845 86.030 ;
        RECT 87.015 85.465 87.355 86.275 ;
        RECT 87.615 86.105 87.785 86.865 ;
        RECT 87.965 86.275 88.295 87.035 ;
        RECT 87.615 85.935 88.280 86.105 ;
        RECT 88.465 85.960 88.735 86.865 ;
        RECT 88.110 85.790 88.280 85.935 ;
        RECT 86.125 85.295 87.355 85.465 ;
        RECT 87.545 85.385 87.875 85.755 ;
        RECT 88.110 85.460 88.395 85.790 ;
        RECT 86.105 84.485 86.615 85.020 ;
        RECT 86.835 84.690 87.080 85.295 ;
        RECT 88.110 85.205 88.280 85.460 ;
        RECT 87.615 85.035 88.280 85.205 ;
        RECT 88.565 85.160 88.735 85.960 ;
        RECT 88.905 85.945 90.575 87.035 ;
        RECT 87.615 84.655 87.785 85.035 ;
        RECT 87.965 84.485 88.295 84.865 ;
        RECT 88.475 84.655 88.735 85.160 ;
        RECT 88.905 85.255 89.655 85.775 ;
        RECT 89.825 85.425 90.575 85.945 ;
        RECT 90.745 85.945 91.955 87.035 ;
        RECT 90.745 85.405 91.265 85.945 ;
        RECT 88.905 84.485 90.575 85.255 ;
        RECT 91.435 85.235 91.955 85.775 ;
        RECT 90.745 84.485 91.955 85.235 ;
        RECT 13.380 84.315 92.040 84.485 ;
        RECT 13.465 83.565 14.675 84.315 ;
        RECT 14.845 83.770 20.190 84.315 ;
        RECT 20.365 83.770 25.710 84.315 ;
        RECT 13.465 83.025 13.985 83.565 ;
        RECT 14.155 82.855 14.675 83.395 ;
        RECT 16.430 82.940 16.770 83.770 ;
        RECT 13.465 81.765 14.675 82.855 ;
        RECT 18.250 82.200 18.600 83.450 ;
        RECT 21.950 82.940 22.290 83.770 ;
        RECT 25.885 83.545 27.555 84.315 ;
        RECT 28.190 83.575 28.445 84.145 ;
        RECT 28.615 83.915 28.945 84.315 ;
        RECT 29.370 83.780 29.900 84.145 ;
        RECT 29.370 83.745 29.545 83.780 ;
        RECT 28.615 83.575 29.545 83.745 ;
        RECT 23.770 82.200 24.120 83.450 ;
        RECT 25.885 83.025 26.635 83.545 ;
        RECT 26.805 82.855 27.555 83.375 ;
        RECT 14.845 81.765 20.190 82.200 ;
        RECT 20.365 81.765 25.710 82.200 ;
        RECT 25.885 81.765 27.555 82.855 ;
        RECT 28.190 82.905 28.360 83.575 ;
        RECT 28.615 83.405 28.785 83.575 ;
        RECT 28.530 83.075 28.785 83.405 ;
        RECT 29.010 83.075 29.205 83.405 ;
        RECT 28.190 81.935 28.525 82.905 ;
        RECT 28.695 81.765 28.865 82.905 ;
        RECT 29.035 82.105 29.205 83.075 ;
        RECT 29.375 82.445 29.545 83.575 ;
        RECT 29.715 82.785 29.885 83.585 ;
        RECT 30.090 83.295 30.365 84.145 ;
        RECT 30.085 83.125 30.365 83.295 ;
        RECT 30.090 82.985 30.365 83.125 ;
        RECT 30.535 82.785 30.725 84.145 ;
        RECT 30.905 83.780 31.415 84.315 ;
        RECT 31.635 83.505 31.880 84.110 ;
        RECT 32.325 83.770 37.670 84.315 ;
        RECT 30.925 83.335 32.155 83.505 ;
        RECT 29.715 82.615 30.725 82.785 ;
        RECT 30.895 82.770 31.645 82.960 ;
        RECT 29.375 82.275 30.500 82.445 ;
        RECT 30.895 82.105 31.065 82.770 ;
        RECT 31.815 82.525 32.155 83.335 ;
        RECT 33.910 82.940 34.250 83.770 ;
        RECT 37.845 83.565 39.055 84.315 ;
        RECT 39.225 83.590 39.515 84.315 ;
        RECT 39.775 83.765 39.945 84.055 ;
        RECT 40.115 83.935 40.445 84.315 ;
        RECT 39.775 83.595 40.440 83.765 ;
        RECT 29.035 81.935 31.065 82.105 ;
        RECT 31.235 81.765 31.405 82.525 ;
        RECT 31.640 82.115 32.155 82.525 ;
        RECT 35.730 82.200 36.080 83.450 ;
        RECT 37.845 83.025 38.365 83.565 ;
        RECT 38.535 82.855 39.055 83.395 ;
        RECT 32.325 81.765 37.670 82.200 ;
        RECT 37.845 81.765 39.055 82.855 ;
        RECT 39.225 81.765 39.515 82.930 ;
        RECT 39.690 82.775 40.040 83.425 ;
        RECT 40.210 82.605 40.440 83.595 ;
        RECT 39.775 82.435 40.440 82.605 ;
        RECT 39.775 81.935 39.945 82.435 ;
        RECT 40.115 81.765 40.445 82.265 ;
        RECT 40.615 81.935 40.800 84.055 ;
        RECT 41.055 83.855 41.305 84.315 ;
        RECT 41.475 83.865 41.810 84.035 ;
        RECT 42.005 83.865 42.680 84.035 ;
        RECT 41.475 83.725 41.645 83.865 ;
        RECT 40.970 82.735 41.250 83.685 ;
        RECT 41.420 83.595 41.645 83.725 ;
        RECT 41.420 82.490 41.590 83.595 ;
        RECT 41.815 83.445 42.340 83.665 ;
        RECT 41.760 82.680 42.000 83.275 ;
        RECT 42.170 82.745 42.340 83.445 ;
        RECT 42.510 83.085 42.680 83.865 ;
        RECT 43.000 83.815 43.370 84.315 ;
        RECT 43.550 83.865 43.955 84.035 ;
        RECT 44.125 83.865 44.910 84.035 ;
        RECT 43.550 83.635 43.720 83.865 ;
        RECT 42.890 83.335 43.720 83.635 ;
        RECT 44.105 83.365 44.570 83.695 ;
        RECT 42.890 83.305 43.090 83.335 ;
        RECT 43.210 83.085 43.380 83.155 ;
        RECT 42.510 82.915 43.380 83.085 ;
        RECT 42.870 82.825 43.380 82.915 ;
        RECT 41.420 82.360 41.725 82.490 ;
        RECT 42.170 82.380 42.700 82.745 ;
        RECT 41.040 81.765 41.305 82.225 ;
        RECT 41.475 81.935 41.725 82.360 ;
        RECT 42.870 82.210 43.040 82.825 ;
        RECT 41.935 82.040 43.040 82.210 ;
        RECT 43.210 81.765 43.380 82.565 ;
        RECT 43.550 82.265 43.720 83.335 ;
        RECT 43.890 82.435 44.080 83.155 ;
        RECT 44.250 82.405 44.570 83.365 ;
        RECT 44.740 83.405 44.910 83.865 ;
        RECT 45.185 83.785 45.395 84.315 ;
        RECT 45.655 83.575 45.985 84.100 ;
        RECT 46.155 83.705 46.325 84.315 ;
        RECT 46.495 83.660 46.825 84.095 ;
        RECT 46.495 83.575 46.875 83.660 ;
        RECT 45.785 83.405 45.985 83.575 ;
        RECT 46.650 83.535 46.875 83.575 ;
        RECT 44.740 83.075 45.615 83.405 ;
        RECT 45.785 83.075 46.535 83.405 ;
        RECT 43.550 81.935 43.800 82.265 ;
        RECT 44.740 82.235 44.910 83.075 ;
        RECT 45.785 82.870 45.975 83.075 ;
        RECT 46.705 82.955 46.875 83.535 ;
        RECT 46.660 82.905 46.875 82.955 ;
        RECT 45.080 82.495 45.975 82.870 ;
        RECT 46.485 82.825 46.875 82.905 ;
        RECT 47.045 83.640 47.315 83.985 ;
        RECT 47.505 83.915 47.885 84.315 ;
        RECT 48.055 83.745 48.225 84.095 ;
        RECT 48.395 83.915 48.725 84.315 ;
        RECT 48.925 83.745 49.095 84.095 ;
        RECT 49.295 83.815 49.625 84.315 ;
        RECT 47.045 82.905 47.215 83.640 ;
        RECT 47.485 83.575 49.095 83.745 ;
        RECT 50.355 83.765 50.525 84.055 ;
        RECT 50.695 83.935 51.025 84.315 ;
        RECT 47.485 83.405 47.655 83.575 ;
        RECT 47.385 83.075 47.655 83.405 ;
        RECT 47.825 83.075 48.230 83.405 ;
        RECT 47.485 82.905 47.655 83.075 ;
        RECT 44.025 82.065 44.910 82.235 ;
        RECT 45.090 81.765 45.405 82.265 ;
        RECT 45.635 81.935 45.975 82.495 ;
        RECT 46.145 81.765 46.315 82.775 ;
        RECT 46.485 81.980 46.815 82.825 ;
        RECT 47.045 81.935 47.315 82.905 ;
        RECT 47.485 82.735 48.210 82.905 ;
        RECT 48.400 82.785 49.110 83.405 ;
        RECT 49.280 83.075 49.630 83.645 ;
        RECT 50.355 83.595 51.020 83.765 ;
        RECT 48.040 82.615 48.210 82.735 ;
        RECT 49.310 82.615 49.630 82.905 ;
        RECT 50.270 82.775 50.620 83.425 ;
        RECT 47.525 81.765 47.805 82.565 ;
        RECT 48.040 82.445 49.630 82.615 ;
        RECT 50.790 82.605 51.020 83.595 ;
        RECT 50.355 82.435 51.020 82.605 ;
        RECT 47.975 81.985 49.630 82.275 ;
        RECT 50.355 81.935 50.525 82.435 ;
        RECT 50.695 81.765 51.025 82.265 ;
        RECT 51.195 81.935 51.380 84.055 ;
        RECT 51.635 83.855 51.885 84.315 ;
        RECT 52.055 83.865 52.390 84.035 ;
        RECT 52.585 83.865 53.260 84.035 ;
        RECT 52.055 83.725 52.225 83.865 ;
        RECT 51.550 82.735 51.830 83.685 ;
        RECT 52.000 83.595 52.225 83.725 ;
        RECT 52.000 82.490 52.170 83.595 ;
        RECT 52.395 83.445 52.920 83.665 ;
        RECT 52.340 82.680 52.580 83.275 ;
        RECT 52.750 82.745 52.920 83.445 ;
        RECT 53.090 83.085 53.260 83.865 ;
        RECT 53.580 83.815 53.950 84.315 ;
        RECT 54.130 83.865 54.535 84.035 ;
        RECT 54.705 83.865 55.490 84.035 ;
        RECT 54.130 83.635 54.300 83.865 ;
        RECT 53.470 83.335 54.300 83.635 ;
        RECT 54.685 83.365 55.150 83.695 ;
        RECT 53.470 83.305 53.670 83.335 ;
        RECT 53.790 83.085 53.960 83.155 ;
        RECT 53.090 82.915 53.960 83.085 ;
        RECT 53.450 82.825 53.960 82.915 ;
        RECT 52.000 82.360 52.305 82.490 ;
        RECT 52.750 82.380 53.280 82.745 ;
        RECT 51.620 81.765 51.885 82.225 ;
        RECT 52.055 81.935 52.305 82.360 ;
        RECT 53.450 82.210 53.620 82.825 ;
        RECT 52.515 82.040 53.620 82.210 ;
        RECT 53.790 81.765 53.960 82.565 ;
        RECT 54.130 82.265 54.300 83.335 ;
        RECT 54.470 82.435 54.660 83.155 ;
        RECT 54.830 82.405 55.150 83.365 ;
        RECT 55.320 83.405 55.490 83.865 ;
        RECT 55.765 83.785 55.975 84.315 ;
        RECT 56.235 83.575 56.565 84.100 ;
        RECT 56.735 83.705 56.905 84.315 ;
        RECT 57.075 83.660 57.405 84.095 ;
        RECT 57.075 83.575 57.455 83.660 ;
        RECT 56.365 83.405 56.565 83.575 ;
        RECT 57.230 83.535 57.455 83.575 ;
        RECT 55.320 83.075 56.195 83.405 ;
        RECT 56.365 83.075 57.115 83.405 ;
        RECT 54.130 81.935 54.380 82.265 ;
        RECT 55.320 82.235 55.490 83.075 ;
        RECT 56.365 82.870 56.555 83.075 ;
        RECT 57.285 82.955 57.455 83.535 ;
        RECT 57.240 82.905 57.455 82.955 ;
        RECT 55.660 82.495 56.555 82.870 ;
        RECT 57.065 82.825 57.455 82.905 ;
        RECT 57.625 83.575 58.010 84.145 ;
        RECT 58.180 83.855 58.505 84.315 ;
        RECT 59.025 83.685 59.305 84.145 ;
        RECT 57.625 82.905 57.905 83.575 ;
        RECT 58.180 83.515 59.305 83.685 ;
        RECT 58.180 83.405 58.630 83.515 ;
        RECT 58.075 83.075 58.630 83.405 ;
        RECT 59.495 83.345 59.895 84.145 ;
        RECT 60.295 83.855 60.565 84.315 ;
        RECT 60.735 83.685 61.020 84.145 ;
        RECT 54.605 82.065 55.490 82.235 ;
        RECT 55.670 81.765 55.985 82.265 ;
        RECT 56.215 81.935 56.555 82.495 ;
        RECT 56.725 81.765 56.895 82.775 ;
        RECT 57.065 81.980 57.395 82.825 ;
        RECT 57.625 81.935 58.010 82.905 ;
        RECT 58.180 82.615 58.630 83.075 ;
        RECT 58.800 82.785 59.895 83.345 ;
        RECT 58.180 82.395 59.305 82.615 ;
        RECT 58.180 81.765 58.505 82.225 ;
        RECT 59.025 81.935 59.305 82.395 ;
        RECT 59.495 81.935 59.895 82.785 ;
        RECT 60.065 83.515 61.020 83.685 ;
        RECT 61.305 83.545 64.815 84.315 ;
        RECT 64.985 83.590 65.275 84.315 ;
        RECT 60.065 82.615 60.275 83.515 ;
        RECT 60.445 82.785 61.135 83.345 ;
        RECT 61.305 83.025 62.955 83.545 ;
        RECT 66.365 83.495 66.625 84.315 ;
        RECT 66.795 83.495 67.125 83.915 ;
        RECT 67.305 83.830 68.095 84.095 ;
        RECT 66.875 83.405 67.125 83.495 ;
        RECT 63.125 82.855 64.815 83.375 ;
        RECT 60.065 82.395 61.020 82.615 ;
        RECT 60.295 81.765 60.565 82.225 ;
        RECT 60.735 81.935 61.020 82.395 ;
        RECT 61.305 81.765 64.815 82.855 ;
        RECT 64.985 81.765 65.275 82.930 ;
        RECT 66.365 82.445 66.705 83.325 ;
        RECT 66.875 83.155 67.670 83.405 ;
        RECT 66.365 81.765 66.625 82.275 ;
        RECT 66.875 81.935 67.045 83.155 ;
        RECT 67.840 82.975 68.095 83.830 ;
        RECT 68.265 83.675 68.465 84.095 ;
        RECT 68.655 83.855 68.985 84.315 ;
        RECT 68.265 83.155 68.675 83.675 ;
        RECT 69.155 83.665 69.415 84.145 ;
        RECT 68.845 82.975 69.075 83.405 ;
        RECT 67.285 82.805 69.075 82.975 ;
        RECT 67.285 82.440 67.535 82.805 ;
        RECT 67.705 82.445 68.035 82.635 ;
        RECT 68.255 82.510 68.970 82.805 ;
        RECT 69.245 82.635 69.415 83.665 ;
        RECT 67.705 82.270 67.900 82.445 ;
        RECT 67.285 81.765 67.900 82.270 ;
        RECT 68.070 81.935 68.545 82.275 ;
        RECT 68.715 81.765 68.930 82.310 ;
        RECT 69.140 81.935 69.415 82.635 ;
        RECT 69.605 83.625 69.845 84.145 ;
        RECT 70.015 83.820 70.410 84.315 ;
        RECT 70.975 83.985 71.145 84.130 ;
        RECT 70.770 83.790 71.145 83.985 ;
        RECT 69.605 82.820 69.780 83.625 ;
        RECT 70.770 83.455 70.940 83.790 ;
        RECT 71.425 83.745 71.665 84.120 ;
        RECT 71.835 83.810 72.170 84.315 ;
        RECT 71.425 83.595 71.645 83.745 ;
        RECT 69.955 83.095 70.940 83.455 ;
        RECT 71.110 83.265 71.645 83.595 ;
        RECT 69.955 83.075 71.240 83.095 ;
        RECT 70.380 82.925 71.240 83.075 ;
        RECT 69.605 82.035 69.910 82.820 ;
        RECT 70.085 82.445 70.780 82.755 ;
        RECT 70.090 81.765 70.775 82.235 ;
        RECT 70.955 81.980 71.240 82.925 ;
        RECT 71.410 82.615 71.645 83.265 ;
        RECT 71.815 82.785 72.115 83.635 ;
        RECT 72.345 83.545 74.935 84.315 ;
        RECT 75.105 83.665 75.365 84.145 ;
        RECT 75.535 83.775 75.785 84.315 ;
        RECT 72.345 83.025 73.555 83.545 ;
        RECT 73.725 82.855 74.935 83.375 ;
        RECT 71.410 82.385 72.085 82.615 ;
        RECT 71.415 81.765 71.745 82.215 ;
        RECT 71.915 81.955 72.085 82.385 ;
        RECT 72.345 81.765 74.935 82.855 ;
        RECT 75.105 82.635 75.275 83.665 ;
        RECT 75.955 83.610 76.175 84.095 ;
        RECT 75.445 83.015 75.675 83.410 ;
        RECT 75.845 83.185 76.175 83.610 ;
        RECT 76.345 83.935 77.235 84.105 ;
        RECT 76.345 83.210 76.515 83.935 ;
        RECT 77.405 83.770 82.750 84.315 ;
        RECT 76.685 83.380 77.235 83.765 ;
        RECT 76.345 83.140 77.235 83.210 ;
        RECT 76.340 83.115 77.235 83.140 ;
        RECT 76.330 83.100 77.235 83.115 ;
        RECT 76.325 83.085 77.235 83.100 ;
        RECT 76.315 83.080 77.235 83.085 ;
        RECT 76.310 83.070 77.235 83.080 ;
        RECT 76.305 83.060 77.235 83.070 ;
        RECT 76.295 83.055 77.235 83.060 ;
        RECT 76.285 83.045 77.235 83.055 ;
        RECT 76.275 83.040 77.235 83.045 ;
        RECT 76.275 83.035 76.610 83.040 ;
        RECT 76.260 83.030 76.610 83.035 ;
        RECT 76.245 83.020 76.610 83.030 ;
        RECT 76.220 83.015 76.610 83.020 ;
        RECT 75.445 83.010 76.610 83.015 ;
        RECT 75.445 82.975 76.580 83.010 ;
        RECT 75.445 82.950 76.545 82.975 ;
        RECT 75.445 82.920 76.515 82.950 ;
        RECT 75.445 82.890 76.495 82.920 ;
        RECT 75.445 82.860 76.475 82.890 ;
        RECT 75.445 82.850 76.405 82.860 ;
        RECT 75.445 82.840 76.380 82.850 ;
        RECT 75.445 82.825 76.360 82.840 ;
        RECT 75.445 82.810 76.340 82.825 ;
        RECT 75.550 82.800 76.335 82.810 ;
        RECT 75.550 82.765 76.320 82.800 ;
        RECT 75.105 81.935 75.380 82.635 ;
        RECT 75.550 82.515 76.305 82.765 ;
        RECT 76.475 82.445 76.805 82.690 ;
        RECT 76.975 82.590 77.235 83.040 ;
        RECT 78.990 82.940 79.330 83.770 ;
        RECT 82.925 83.545 85.515 84.315 ;
        RECT 85.775 83.765 85.945 84.145 ;
        RECT 86.125 83.935 86.455 84.315 ;
        RECT 85.775 83.595 86.440 83.765 ;
        RECT 86.635 83.640 86.895 84.145 ;
        RECT 76.620 82.420 76.805 82.445 ;
        RECT 76.620 82.320 77.235 82.420 ;
        RECT 75.550 81.765 75.805 82.310 ;
        RECT 75.975 81.935 76.455 82.275 ;
        RECT 76.630 81.765 77.235 82.320 ;
        RECT 80.810 82.200 81.160 83.450 ;
        RECT 82.925 83.025 84.135 83.545 ;
        RECT 84.305 82.855 85.515 83.375 ;
        RECT 85.705 83.045 86.035 83.415 ;
        RECT 86.270 83.340 86.440 83.595 ;
        RECT 86.270 83.010 86.555 83.340 ;
        RECT 86.270 82.865 86.440 83.010 ;
        RECT 77.405 81.765 82.750 82.200 ;
        RECT 82.925 81.765 85.515 82.855 ;
        RECT 85.775 82.695 86.440 82.865 ;
        RECT 86.725 82.840 86.895 83.640 ;
        RECT 85.775 81.935 85.945 82.695 ;
        RECT 86.125 81.765 86.455 82.525 ;
        RECT 86.625 81.935 86.895 82.840 ;
        RECT 87.065 83.575 87.450 84.145 ;
        RECT 87.620 83.855 87.945 84.315 ;
        RECT 88.465 83.685 88.745 84.145 ;
        RECT 87.065 82.905 87.345 83.575 ;
        RECT 87.620 83.515 88.745 83.685 ;
        RECT 87.620 83.405 88.070 83.515 ;
        RECT 87.515 83.075 88.070 83.405 ;
        RECT 88.935 83.345 89.335 84.145 ;
        RECT 89.735 83.855 90.005 84.315 ;
        RECT 90.175 83.685 90.460 84.145 ;
        RECT 87.065 81.935 87.450 82.905 ;
        RECT 87.620 82.615 88.070 83.075 ;
        RECT 88.240 82.785 89.335 83.345 ;
        RECT 87.620 82.395 88.745 82.615 ;
        RECT 87.620 81.765 87.945 82.225 ;
        RECT 88.465 81.935 88.745 82.395 ;
        RECT 88.935 81.935 89.335 82.785 ;
        RECT 89.505 83.515 90.460 83.685 ;
        RECT 90.745 83.565 91.955 84.315 ;
        RECT 89.505 82.615 89.715 83.515 ;
        RECT 89.885 82.785 90.575 83.345 ;
        RECT 90.745 82.855 91.265 83.395 ;
        RECT 91.435 83.025 91.955 83.565 ;
        RECT 89.505 82.395 90.460 82.615 ;
        RECT 89.735 81.765 90.005 82.225 ;
        RECT 90.175 81.935 90.460 82.395 ;
        RECT 90.745 81.765 91.955 82.855 ;
        RECT 13.380 81.595 92.040 81.765 ;
        RECT 13.465 80.505 14.675 81.595 ;
        RECT 14.845 80.505 16.515 81.595 ;
        RECT 13.465 79.795 13.985 80.335 ;
        RECT 14.155 79.965 14.675 80.505 ;
        RECT 14.845 79.815 15.595 80.335 ;
        RECT 15.765 79.985 16.515 80.505 ;
        RECT 17.145 80.875 17.605 81.425 ;
        RECT 17.795 80.875 18.125 81.595 ;
        RECT 13.465 79.045 14.675 79.795 ;
        RECT 14.845 79.045 16.515 79.815 ;
        RECT 17.145 79.505 17.395 80.875 ;
        RECT 18.325 80.705 18.625 81.255 ;
        RECT 18.795 80.925 19.075 81.595 ;
        RECT 17.685 80.535 18.625 80.705 ;
        RECT 17.685 80.285 17.855 80.535 ;
        RECT 18.995 80.285 19.260 80.645 ;
        RECT 19.445 80.455 19.705 81.595 ;
        RECT 19.875 80.445 20.205 81.425 ;
        RECT 20.375 80.455 20.655 81.595 ;
        RECT 20.835 80.625 21.165 81.410 ;
        RECT 20.835 80.455 21.515 80.625 ;
        RECT 21.695 80.455 22.025 81.595 ;
        RECT 23.125 80.455 23.385 81.595 ;
        RECT 23.625 81.085 25.240 81.415 ;
        RECT 19.965 80.405 20.140 80.445 ;
        RECT 17.565 79.955 17.855 80.285 ;
        RECT 18.025 80.035 18.365 80.285 ;
        RECT 18.585 80.035 19.260 80.285 ;
        RECT 19.465 80.035 19.800 80.285 ;
        RECT 17.685 79.865 17.855 79.955 ;
        RECT 17.685 79.675 19.075 79.865 ;
        RECT 19.970 79.845 20.140 80.405 ;
        RECT 20.310 80.015 20.645 80.285 ;
        RECT 20.825 80.035 21.175 80.285 ;
        RECT 21.345 79.855 21.515 80.455 ;
        RECT 23.635 80.285 23.805 80.845 ;
        RECT 24.065 80.745 25.240 80.915 ;
        RECT 25.410 80.795 25.690 81.595 ;
        RECT 24.065 80.455 24.395 80.745 ;
        RECT 25.070 80.625 25.240 80.745 ;
        RECT 24.565 80.285 24.810 80.575 ;
        RECT 25.070 80.455 25.730 80.625 ;
        RECT 25.900 80.455 26.175 81.425 ;
        RECT 25.560 80.285 25.730 80.455 ;
        RECT 21.685 80.035 22.035 80.285 ;
        RECT 23.130 80.035 23.465 80.285 ;
        RECT 23.635 79.955 24.350 80.285 ;
        RECT 24.565 79.955 25.390 80.285 ;
        RECT 25.560 79.955 25.835 80.285 ;
        RECT 23.635 79.865 23.885 79.955 ;
        RECT 17.145 79.215 17.705 79.505 ;
        RECT 17.875 79.045 18.125 79.505 ;
        RECT 18.745 79.315 19.075 79.675 ;
        RECT 19.445 79.215 20.140 79.845 ;
        RECT 20.345 79.045 20.655 79.845 ;
        RECT 20.845 79.045 21.085 79.855 ;
        RECT 21.255 79.215 21.585 79.855 ;
        RECT 21.755 79.045 22.025 79.855 ;
        RECT 23.125 79.045 23.385 79.865 ;
        RECT 23.555 79.445 23.885 79.865 ;
        RECT 25.560 79.785 25.730 79.955 ;
        RECT 24.065 79.615 25.730 79.785 ;
        RECT 26.005 79.720 26.175 80.455 ;
        RECT 26.345 80.430 26.635 81.595 ;
        RECT 26.805 80.505 28.015 81.595 ;
        RECT 26.805 79.795 27.325 80.335 ;
        RECT 27.495 79.965 28.015 80.505 ;
        RECT 28.190 80.455 28.525 81.425 ;
        RECT 28.695 80.455 28.865 81.595 ;
        RECT 29.035 81.255 31.065 81.425 ;
        RECT 24.065 79.215 24.325 79.615 ;
        RECT 24.495 79.045 24.825 79.445 ;
        RECT 24.995 79.265 25.165 79.615 ;
        RECT 25.335 79.045 25.710 79.445 ;
        RECT 25.900 79.375 26.175 79.720 ;
        RECT 26.345 79.045 26.635 79.770 ;
        RECT 26.805 79.045 28.015 79.795 ;
        RECT 28.190 79.785 28.360 80.455 ;
        RECT 29.035 80.285 29.205 81.255 ;
        RECT 28.530 79.955 28.785 80.285 ;
        RECT 29.010 79.955 29.205 80.285 ;
        RECT 29.375 80.915 30.500 81.085 ;
        RECT 28.615 79.785 28.785 79.955 ;
        RECT 29.375 79.785 29.545 80.915 ;
        RECT 28.190 79.215 28.445 79.785 ;
        RECT 28.615 79.615 29.545 79.785 ;
        RECT 29.715 80.575 30.725 80.745 ;
        RECT 29.715 79.775 29.885 80.575 ;
        RECT 30.090 80.235 30.365 80.375 ;
        RECT 30.085 80.065 30.365 80.235 ;
        RECT 29.370 79.580 29.545 79.615 ;
        RECT 28.615 79.045 28.945 79.445 ;
        RECT 29.370 79.215 29.900 79.580 ;
        RECT 30.090 79.215 30.365 80.065 ;
        RECT 30.535 79.215 30.725 80.575 ;
        RECT 30.895 80.590 31.065 81.255 ;
        RECT 31.235 80.835 31.405 81.595 ;
        RECT 31.640 80.835 32.155 81.245 ;
        RECT 32.325 81.160 37.670 81.595 ;
        RECT 30.895 80.400 31.645 80.590 ;
        RECT 31.815 80.025 32.155 80.835 ;
        RECT 30.925 79.855 32.155 80.025 ;
        RECT 30.905 79.045 31.415 79.580 ;
        RECT 31.635 79.250 31.880 79.855 ;
        RECT 33.910 79.590 34.250 80.420 ;
        RECT 35.730 79.910 36.080 81.160 ;
        RECT 38.765 80.835 39.280 81.245 ;
        RECT 39.515 80.835 39.685 81.595 ;
        RECT 39.855 81.255 41.885 81.425 ;
        RECT 38.765 80.025 39.105 80.835 ;
        RECT 39.855 80.590 40.025 81.255 ;
        RECT 40.420 80.915 41.545 81.085 ;
        RECT 39.275 80.400 40.025 80.590 ;
        RECT 40.195 80.575 41.205 80.745 ;
        RECT 38.765 79.855 39.995 80.025 ;
        RECT 32.325 79.045 37.670 79.590 ;
        RECT 39.040 79.250 39.285 79.855 ;
        RECT 39.505 79.045 40.015 79.580 ;
        RECT 40.195 79.215 40.385 80.575 ;
        RECT 40.555 79.555 40.830 80.375 ;
        RECT 41.035 79.775 41.205 80.575 ;
        RECT 41.375 79.785 41.545 80.915 ;
        RECT 41.715 80.285 41.885 81.255 ;
        RECT 42.055 80.455 42.225 81.595 ;
        RECT 42.395 80.455 42.730 81.425 ;
        RECT 42.905 80.505 44.575 81.595 ;
        RECT 41.715 79.955 41.910 80.285 ;
        RECT 42.135 79.955 42.390 80.285 ;
        RECT 42.135 79.785 42.305 79.955 ;
        RECT 42.560 79.785 42.730 80.455 ;
        RECT 41.375 79.615 42.305 79.785 ;
        RECT 41.375 79.580 41.550 79.615 ;
        RECT 40.555 79.385 40.835 79.555 ;
        RECT 40.555 79.215 40.830 79.385 ;
        RECT 41.020 79.215 41.550 79.580 ;
        RECT 41.975 79.045 42.305 79.445 ;
        RECT 42.475 79.215 42.730 79.785 ;
        RECT 42.905 79.815 43.655 80.335 ;
        RECT 43.825 79.985 44.575 80.505 ;
        RECT 44.745 80.455 45.130 81.425 ;
        RECT 45.300 81.135 45.625 81.595 ;
        RECT 46.145 80.965 46.425 81.425 ;
        RECT 45.300 80.745 46.425 80.965 ;
        RECT 42.905 79.045 44.575 79.815 ;
        RECT 44.745 79.785 45.025 80.455 ;
        RECT 45.300 80.285 45.750 80.745 ;
        RECT 46.615 80.575 47.015 81.425 ;
        RECT 47.415 81.135 47.685 81.595 ;
        RECT 47.855 80.965 48.140 81.425 ;
        RECT 45.195 79.955 45.750 80.285 ;
        RECT 45.920 80.015 47.015 80.575 ;
        RECT 45.300 79.845 45.750 79.955 ;
        RECT 44.745 79.215 45.130 79.785 ;
        RECT 45.300 79.675 46.425 79.845 ;
        RECT 45.300 79.045 45.625 79.505 ;
        RECT 46.145 79.215 46.425 79.675 ;
        RECT 46.615 79.215 47.015 80.015 ;
        RECT 47.185 80.745 48.140 80.965 ;
        RECT 48.540 80.965 48.825 81.425 ;
        RECT 48.995 81.135 49.265 81.595 ;
        RECT 48.540 80.745 49.495 80.965 ;
        RECT 47.185 79.845 47.395 80.745 ;
        RECT 47.565 80.015 48.255 80.575 ;
        RECT 48.425 80.015 49.115 80.575 ;
        RECT 49.285 79.845 49.495 80.745 ;
        RECT 47.185 79.675 48.140 79.845 ;
        RECT 47.415 79.045 47.685 79.505 ;
        RECT 47.855 79.215 48.140 79.675 ;
        RECT 48.540 79.675 49.495 79.845 ;
        RECT 49.665 80.575 50.065 81.425 ;
        RECT 50.255 80.965 50.535 81.425 ;
        RECT 51.055 81.135 51.380 81.595 ;
        RECT 50.255 80.745 51.380 80.965 ;
        RECT 49.665 80.015 50.760 80.575 ;
        RECT 50.930 80.285 51.380 80.745 ;
        RECT 51.550 80.455 51.935 81.425 ;
        RECT 48.540 79.215 48.825 79.675 ;
        RECT 48.995 79.045 49.265 79.505 ;
        RECT 49.665 79.215 50.065 80.015 ;
        RECT 50.930 79.955 51.485 80.285 ;
        RECT 50.930 79.845 51.380 79.955 ;
        RECT 50.255 79.675 51.380 79.845 ;
        RECT 51.655 79.785 51.935 80.455 ;
        RECT 52.105 80.430 52.395 81.595 ;
        RECT 52.565 80.725 52.840 81.425 ;
        RECT 53.010 81.050 53.265 81.595 ;
        RECT 53.435 81.085 53.915 81.425 ;
        RECT 54.090 81.040 54.695 81.595 ;
        RECT 54.080 80.940 54.695 81.040 ;
        RECT 54.080 80.915 54.265 80.940 ;
        RECT 50.255 79.215 50.535 79.675 ;
        RECT 51.055 79.045 51.380 79.505 ;
        RECT 51.550 79.215 51.935 79.785 ;
        RECT 52.105 79.045 52.395 79.770 ;
        RECT 52.565 79.695 52.735 80.725 ;
        RECT 53.010 80.595 53.765 80.845 ;
        RECT 53.935 80.670 54.265 80.915 ;
        RECT 53.010 80.560 53.780 80.595 ;
        RECT 53.010 80.550 53.795 80.560 ;
        RECT 52.905 80.535 53.800 80.550 ;
        RECT 52.905 80.520 53.820 80.535 ;
        RECT 52.905 80.510 53.840 80.520 ;
        RECT 52.905 80.500 53.865 80.510 ;
        RECT 52.905 80.470 53.935 80.500 ;
        RECT 52.905 80.440 53.955 80.470 ;
        RECT 52.905 80.410 53.975 80.440 ;
        RECT 52.905 80.385 54.005 80.410 ;
        RECT 52.905 80.350 54.040 80.385 ;
        RECT 52.905 80.345 54.070 80.350 ;
        RECT 52.905 79.950 53.135 80.345 ;
        RECT 53.680 80.340 54.070 80.345 ;
        RECT 53.705 80.330 54.070 80.340 ;
        RECT 53.720 80.325 54.070 80.330 ;
        RECT 53.735 80.320 54.070 80.325 ;
        RECT 54.435 80.320 54.695 80.770 ;
        RECT 53.735 80.315 54.695 80.320 ;
        RECT 53.745 80.305 54.695 80.315 ;
        RECT 53.755 80.300 54.695 80.305 ;
        RECT 53.765 80.290 54.695 80.300 ;
        RECT 53.770 80.280 54.695 80.290 ;
        RECT 53.775 80.275 54.695 80.280 ;
        RECT 53.785 80.260 54.695 80.275 ;
        RECT 53.790 80.245 54.695 80.260 ;
        RECT 53.800 80.220 54.695 80.245 ;
        RECT 53.305 79.750 53.635 80.175 ;
        RECT 52.565 79.215 52.825 79.695 ;
        RECT 52.995 79.045 53.245 79.585 ;
        RECT 53.415 79.265 53.635 79.750 ;
        RECT 53.805 80.150 54.695 80.220 ;
        RECT 54.870 80.455 55.205 81.425 ;
        RECT 55.375 80.455 55.545 81.595 ;
        RECT 55.715 81.255 57.745 81.425 ;
        RECT 53.805 79.425 53.975 80.150 ;
        RECT 54.145 79.595 54.695 79.980 ;
        RECT 54.870 79.785 55.040 80.455 ;
        RECT 55.715 80.285 55.885 81.255 ;
        RECT 55.210 79.955 55.465 80.285 ;
        RECT 55.690 79.955 55.885 80.285 ;
        RECT 56.055 80.915 57.180 81.085 ;
        RECT 55.295 79.785 55.465 79.955 ;
        RECT 56.055 79.785 56.225 80.915 ;
        RECT 53.805 79.255 54.695 79.425 ;
        RECT 54.870 79.215 55.125 79.785 ;
        RECT 55.295 79.615 56.225 79.785 ;
        RECT 56.395 80.575 57.405 80.745 ;
        RECT 56.395 79.775 56.565 80.575 ;
        RECT 56.050 79.580 56.225 79.615 ;
        RECT 55.295 79.045 55.625 79.445 ;
        RECT 56.050 79.215 56.580 79.580 ;
        RECT 56.770 79.555 57.045 80.375 ;
        RECT 56.765 79.385 57.045 79.555 ;
        RECT 56.770 79.215 57.045 79.385 ;
        RECT 57.215 79.215 57.405 80.575 ;
        RECT 57.575 80.590 57.745 81.255 ;
        RECT 57.915 80.835 58.085 81.595 ;
        RECT 58.320 80.835 58.835 81.245 ;
        RECT 59.005 81.160 64.350 81.595 ;
        RECT 57.575 80.400 58.325 80.590 ;
        RECT 58.495 80.025 58.835 80.835 ;
        RECT 57.605 79.855 58.835 80.025 ;
        RECT 57.585 79.045 58.095 79.580 ;
        RECT 58.315 79.250 58.560 79.855 ;
        RECT 60.590 79.590 60.930 80.420 ;
        RECT 62.410 79.910 62.760 81.160 ;
        RECT 64.640 80.965 64.925 81.425 ;
        RECT 65.095 81.135 65.365 81.595 ;
        RECT 64.640 80.745 65.595 80.965 ;
        RECT 64.525 80.015 65.215 80.575 ;
        RECT 65.385 79.845 65.595 80.745 ;
        RECT 64.640 79.675 65.595 79.845 ;
        RECT 65.765 80.575 66.165 81.425 ;
        RECT 66.355 80.965 66.635 81.425 ;
        RECT 67.155 81.135 67.480 81.595 ;
        RECT 66.355 80.745 67.480 80.965 ;
        RECT 65.765 80.015 66.860 80.575 ;
        RECT 67.030 80.285 67.480 80.745 ;
        RECT 67.650 80.455 68.035 81.425 ;
        RECT 68.205 81.040 68.810 81.595 ;
        RECT 68.985 81.085 69.465 81.425 ;
        RECT 69.635 81.050 69.890 81.595 ;
        RECT 68.205 80.940 68.820 81.040 ;
        RECT 68.635 80.915 68.820 80.940 ;
        RECT 59.005 79.045 64.350 79.590 ;
        RECT 64.640 79.215 64.925 79.675 ;
        RECT 65.095 79.045 65.365 79.505 ;
        RECT 65.765 79.215 66.165 80.015 ;
        RECT 67.030 79.955 67.585 80.285 ;
        RECT 67.030 79.845 67.480 79.955 ;
        RECT 66.355 79.675 67.480 79.845 ;
        RECT 67.755 79.785 68.035 80.455 ;
        RECT 68.205 80.320 68.465 80.770 ;
        RECT 68.635 80.670 68.965 80.915 ;
        RECT 69.135 80.595 69.890 80.845 ;
        RECT 70.060 80.725 70.335 81.425 ;
        RECT 69.120 80.560 69.890 80.595 ;
        RECT 69.105 80.550 69.890 80.560 ;
        RECT 69.100 80.535 69.995 80.550 ;
        RECT 69.080 80.520 69.995 80.535 ;
        RECT 69.060 80.510 69.995 80.520 ;
        RECT 69.035 80.500 69.995 80.510 ;
        RECT 68.965 80.470 69.995 80.500 ;
        RECT 68.945 80.440 69.995 80.470 ;
        RECT 68.925 80.410 69.995 80.440 ;
        RECT 68.895 80.385 69.995 80.410 ;
        RECT 68.860 80.350 69.995 80.385 ;
        RECT 68.830 80.345 69.995 80.350 ;
        RECT 68.830 80.340 69.220 80.345 ;
        RECT 68.830 80.330 69.195 80.340 ;
        RECT 68.830 80.325 69.180 80.330 ;
        RECT 68.830 80.320 69.165 80.325 ;
        RECT 68.205 80.315 69.165 80.320 ;
        RECT 68.205 80.305 69.155 80.315 ;
        RECT 68.205 80.300 69.145 80.305 ;
        RECT 68.205 80.290 69.135 80.300 ;
        RECT 68.205 80.280 69.130 80.290 ;
        RECT 68.205 80.275 69.125 80.280 ;
        RECT 68.205 80.260 69.115 80.275 ;
        RECT 68.205 80.245 69.110 80.260 ;
        RECT 68.205 80.220 69.100 80.245 ;
        RECT 68.205 80.150 69.095 80.220 ;
        RECT 66.355 79.215 66.635 79.675 ;
        RECT 67.155 79.045 67.480 79.505 ;
        RECT 67.650 79.215 68.035 79.785 ;
        RECT 68.205 79.595 68.755 79.980 ;
        RECT 68.925 79.425 69.095 80.150 ;
        RECT 68.205 79.255 69.095 79.425 ;
        RECT 69.265 79.750 69.595 80.175 ;
        RECT 69.765 79.950 69.995 80.345 ;
        RECT 69.265 79.265 69.485 79.750 ;
        RECT 70.165 79.695 70.335 80.725 ;
        RECT 70.505 80.505 73.095 81.595 ;
        RECT 69.655 79.045 69.905 79.585 ;
        RECT 70.075 79.215 70.335 79.695 ;
        RECT 70.505 79.815 71.715 80.335 ;
        RECT 71.885 79.985 73.095 80.505 ;
        RECT 73.880 80.585 74.180 81.425 ;
        RECT 74.375 80.755 74.625 81.595 ;
        RECT 75.215 81.005 76.020 81.425 ;
        RECT 74.795 80.835 76.360 81.005 ;
        RECT 74.795 80.585 74.965 80.835 ;
        RECT 73.880 80.415 74.965 80.585 ;
        RECT 73.725 79.955 74.055 80.245 ;
        RECT 70.505 79.045 73.095 79.815 ;
        RECT 74.225 79.785 74.395 80.415 ;
        RECT 75.135 80.285 75.455 80.665 ;
        RECT 74.565 80.035 74.895 80.245 ;
        RECT 75.075 80.035 75.455 80.285 ;
        RECT 75.645 80.245 76.020 80.665 ;
        RECT 76.190 80.585 76.360 80.835 ;
        RECT 76.530 80.755 76.860 81.595 ;
        RECT 77.030 80.835 77.695 81.425 ;
        RECT 76.190 80.415 77.110 80.585 ;
        RECT 76.940 80.245 77.110 80.415 ;
        RECT 75.645 80.235 76.130 80.245 ;
        RECT 75.625 80.065 76.130 80.235 ;
        RECT 75.645 80.035 76.130 80.065 ;
        RECT 76.320 80.035 76.770 80.245 ;
        RECT 76.940 80.035 77.275 80.245 ;
        RECT 77.445 79.865 77.695 80.835 ;
        RECT 77.865 80.430 78.155 81.595 ;
        RECT 78.330 81.205 78.665 81.425 ;
        RECT 79.670 81.215 80.025 81.595 ;
        RECT 78.330 80.585 78.585 81.205 ;
        RECT 78.835 81.045 79.065 81.085 ;
        RECT 80.195 81.045 80.445 81.425 ;
        RECT 78.835 80.845 80.445 81.045 ;
        RECT 78.835 80.755 79.020 80.845 ;
        RECT 79.610 80.835 80.445 80.845 ;
        RECT 80.695 80.815 80.945 81.595 ;
        RECT 81.115 80.745 81.375 81.425 ;
        RECT 81.635 80.925 81.805 81.425 ;
        RECT 81.975 81.095 82.305 81.595 ;
        RECT 81.635 80.755 82.300 80.925 ;
        RECT 79.175 80.645 79.505 80.675 ;
        RECT 79.175 80.585 80.975 80.645 ;
        RECT 78.330 80.475 81.035 80.585 ;
        RECT 78.330 80.415 79.505 80.475 ;
        RECT 80.835 80.440 81.035 80.475 ;
        RECT 78.325 80.035 78.815 80.235 ;
        RECT 79.005 80.035 79.480 80.245 ;
        RECT 73.885 79.605 74.395 79.785 ;
        RECT 74.800 79.695 76.500 79.865 ;
        RECT 74.800 79.605 75.185 79.695 ;
        RECT 73.885 79.215 74.215 79.605 ;
        RECT 74.385 79.265 75.570 79.435 ;
        RECT 75.830 79.045 76.000 79.515 ;
        RECT 76.170 79.230 76.500 79.695 ;
        RECT 76.670 79.045 76.840 79.865 ;
        RECT 77.010 79.225 77.695 79.865 ;
        RECT 77.865 79.045 78.155 79.770 ;
        RECT 78.330 79.045 78.785 79.810 ;
        RECT 79.260 79.635 79.480 80.035 ;
        RECT 79.725 80.035 80.055 80.245 ;
        RECT 79.725 79.635 79.935 80.035 ;
        RECT 80.225 80.000 80.635 80.305 ;
        RECT 80.865 79.865 81.035 80.440 ;
        RECT 80.765 79.745 81.035 79.865 ;
        RECT 80.190 79.700 81.035 79.745 ;
        RECT 80.190 79.575 80.945 79.700 ;
        RECT 80.190 79.425 80.360 79.575 ;
        RECT 81.205 79.555 81.375 80.745 ;
        RECT 81.550 79.935 81.900 80.585 ;
        RECT 82.070 79.765 82.300 80.755 ;
        RECT 81.145 79.545 81.375 79.555 ;
        RECT 79.060 79.215 80.360 79.425 ;
        RECT 80.615 79.045 80.945 79.405 ;
        RECT 81.115 79.215 81.375 79.545 ;
        RECT 81.635 79.595 82.300 79.765 ;
        RECT 81.635 79.305 81.805 79.595 ;
        RECT 81.975 79.045 82.305 79.425 ;
        RECT 82.475 79.305 82.660 81.425 ;
        RECT 82.900 81.135 83.165 81.595 ;
        RECT 83.335 81.000 83.585 81.425 ;
        RECT 83.795 81.150 84.900 81.320 ;
        RECT 83.280 80.870 83.585 81.000 ;
        RECT 82.830 79.675 83.110 80.625 ;
        RECT 83.280 79.765 83.450 80.870 ;
        RECT 83.620 80.085 83.860 80.680 ;
        RECT 84.030 80.615 84.560 80.980 ;
        RECT 84.030 79.915 84.200 80.615 ;
        RECT 84.730 80.535 84.900 81.150 ;
        RECT 85.070 80.795 85.240 81.595 ;
        RECT 85.410 81.095 85.660 81.425 ;
        RECT 85.885 81.125 86.770 81.295 ;
        RECT 84.730 80.445 85.240 80.535 ;
        RECT 83.280 79.635 83.505 79.765 ;
        RECT 83.675 79.695 84.200 79.915 ;
        RECT 84.370 80.275 85.240 80.445 ;
        RECT 82.915 79.045 83.165 79.505 ;
        RECT 83.335 79.495 83.505 79.635 ;
        RECT 84.370 79.495 84.540 80.275 ;
        RECT 85.070 80.205 85.240 80.275 ;
        RECT 84.750 80.025 84.950 80.055 ;
        RECT 85.410 80.025 85.580 81.095 ;
        RECT 85.750 80.205 85.940 80.925 ;
        RECT 84.750 79.725 85.580 80.025 ;
        RECT 86.110 79.995 86.430 80.955 ;
        RECT 83.335 79.325 83.670 79.495 ;
        RECT 83.865 79.325 84.540 79.495 ;
        RECT 84.860 79.045 85.230 79.545 ;
        RECT 85.410 79.495 85.580 79.725 ;
        RECT 85.965 79.665 86.430 79.995 ;
        RECT 86.600 80.285 86.770 81.125 ;
        RECT 86.950 81.095 87.265 81.595 ;
        RECT 87.495 80.865 87.835 81.425 ;
        RECT 86.940 80.490 87.835 80.865 ;
        RECT 88.005 80.585 88.175 81.595 ;
        RECT 87.645 80.285 87.835 80.490 ;
        RECT 88.345 80.535 88.675 81.380 ;
        RECT 88.995 80.665 89.165 81.425 ;
        RECT 89.380 80.835 89.710 81.595 ;
        RECT 88.345 80.455 88.735 80.535 ;
        RECT 88.995 80.495 89.710 80.665 ;
        RECT 89.880 80.520 90.135 81.425 ;
        RECT 88.520 80.405 88.735 80.455 ;
        RECT 86.600 79.955 87.475 80.285 ;
        RECT 87.645 79.955 88.395 80.285 ;
        RECT 86.600 79.495 86.770 79.955 ;
        RECT 87.645 79.785 87.845 79.955 ;
        RECT 88.565 79.825 88.735 80.405 ;
        RECT 88.905 79.945 89.260 80.315 ;
        RECT 89.540 80.285 89.710 80.495 ;
        RECT 89.540 79.955 89.795 80.285 ;
        RECT 88.510 79.785 88.735 79.825 ;
        RECT 85.410 79.325 85.815 79.495 ;
        RECT 85.985 79.325 86.770 79.495 ;
        RECT 87.045 79.045 87.255 79.575 ;
        RECT 87.515 79.260 87.845 79.785 ;
        RECT 88.355 79.700 88.735 79.785 ;
        RECT 89.540 79.765 89.710 79.955 ;
        RECT 89.965 79.790 90.135 80.520 ;
        RECT 90.310 80.445 90.570 81.595 ;
        RECT 90.745 80.505 91.955 81.595 ;
        RECT 99.990 81.095 100.160 87.615 ;
        RECT 100.640 84.975 100.990 87.135 ;
        RECT 100.640 81.575 100.990 83.735 ;
        RECT 101.470 81.095 101.640 87.615 ;
        RECT 102.120 84.975 102.470 87.135 ;
        RECT 102.120 81.575 102.470 83.735 ;
        RECT 102.950 81.095 103.120 87.615 ;
        RECT 103.600 84.975 103.950 87.135 ;
        RECT 103.600 81.575 103.950 83.735 ;
        RECT 104.430 81.095 104.600 87.615 ;
        RECT 105.080 84.975 105.430 87.135 ;
        RECT 105.080 81.575 105.430 83.735 ;
        RECT 105.910 81.095 106.080 87.615 ;
        RECT 106.560 84.975 106.910 87.135 ;
        RECT 106.560 81.575 106.910 83.735 ;
        RECT 107.390 81.095 107.560 87.615 ;
        RECT 108.040 84.975 108.390 87.135 ;
        RECT 108.040 81.575 108.390 83.735 ;
        RECT 108.870 81.095 109.040 87.615 ;
        RECT 109.520 84.975 109.870 87.135 ;
        RECT 109.520 81.575 109.870 83.735 ;
        RECT 110.350 81.095 110.520 87.615 ;
        RECT 111.000 84.975 111.350 87.135 ;
        RECT 111.000 81.575 111.350 83.735 ;
        RECT 111.830 81.095 112.000 87.615 ;
        RECT 112.480 84.975 112.830 87.135 ;
        RECT 112.480 81.575 112.830 83.735 ;
        RECT 113.310 81.095 113.480 87.615 ;
        RECT 117.590 82.770 117.760 92.260 ;
        RECT 118.390 91.750 119.390 91.920 ;
        RECT 118.160 83.495 118.330 91.535 ;
        RECT 119.450 83.495 119.620 91.535 ;
        RECT 118.390 83.110 119.390 83.280 ;
        RECT 120.020 82.770 120.190 92.260 ;
        RECT 120.820 91.750 122.820 91.920 ;
        RECT 120.590 83.495 120.760 91.535 ;
        RECT 122.880 83.495 123.050 91.535 ;
        RECT 120.820 83.110 122.820 83.280 ;
        RECT 123.450 82.770 123.620 92.260 ;
        RECT 124.250 91.750 126.250 91.920 ;
        RECT 124.020 83.495 124.190 91.535 ;
        RECT 126.310 83.495 126.480 91.535 ;
        RECT 124.250 83.110 126.250 83.280 ;
        RECT 126.880 82.770 127.050 92.260 ;
        RECT 127.680 91.750 128.680 91.920 ;
        RECT 127.450 83.495 127.620 91.535 ;
        RECT 128.740 83.495 128.910 91.535 ;
        RECT 129.310 86.660 130.440 92.260 ;
        RECT 127.680 83.110 128.680 83.280 ;
        RECT 129.310 82.770 130.460 86.660 ;
        RECT 134.410 84.640 139.730 85.560 ;
        RECT 134.410 84.540 136.170 84.640 ;
        RECT 117.590 82.600 130.460 82.770 ;
        RECT 129.340 82.570 130.460 82.600 ;
        RECT 99.990 80.925 113.480 81.095 ;
        RECT 129.450 81.350 130.450 82.570 ;
        RECT 126.900 81.010 129.140 81.020 ;
        RECT 90.745 79.965 91.265 80.505 ;
        RECT 88.015 79.045 88.185 79.655 ;
        RECT 88.355 79.265 88.685 79.700 ;
        RECT 88.995 79.595 89.710 79.765 ;
        RECT 88.995 79.215 89.165 79.595 ;
        RECT 89.380 79.045 89.710 79.425 ;
        RECT 89.880 79.215 90.135 79.790 ;
        RECT 90.310 79.045 90.570 79.885 ;
        RECT 91.435 79.795 91.955 80.335 ;
        RECT 90.745 79.045 91.955 79.795 ;
        RECT 13.380 78.875 92.040 79.045 ;
        RECT 13.465 78.125 14.675 78.875 ;
        RECT 15.855 78.325 16.025 78.615 ;
        RECT 16.195 78.495 16.525 78.875 ;
        RECT 15.855 78.155 16.520 78.325 ;
        RECT 13.465 77.585 13.985 78.125 ;
        RECT 14.155 77.415 14.675 77.955 ;
        RECT 13.465 76.325 14.675 77.415 ;
        RECT 15.770 77.335 16.120 77.985 ;
        RECT 16.290 77.165 16.520 78.155 ;
        RECT 15.855 76.995 16.520 77.165 ;
        RECT 15.855 76.495 16.025 76.995 ;
        RECT 16.195 76.325 16.525 76.825 ;
        RECT 16.695 76.495 16.880 78.615 ;
        RECT 17.135 78.415 17.385 78.875 ;
        RECT 17.555 78.425 17.890 78.595 ;
        RECT 18.085 78.425 18.760 78.595 ;
        RECT 17.555 78.285 17.725 78.425 ;
        RECT 17.050 77.295 17.330 78.245 ;
        RECT 17.500 78.155 17.725 78.285 ;
        RECT 17.500 77.050 17.670 78.155 ;
        RECT 17.895 78.005 18.420 78.225 ;
        RECT 17.840 77.240 18.080 77.835 ;
        RECT 18.250 77.305 18.420 78.005 ;
        RECT 18.590 77.645 18.760 78.425 ;
        RECT 19.080 78.375 19.450 78.875 ;
        RECT 19.630 78.425 20.035 78.595 ;
        RECT 20.205 78.425 20.990 78.595 ;
        RECT 19.630 78.195 19.800 78.425 ;
        RECT 18.970 77.895 19.800 78.195 ;
        RECT 20.185 77.925 20.650 78.255 ;
        RECT 18.970 77.865 19.170 77.895 ;
        RECT 19.290 77.645 19.460 77.715 ;
        RECT 18.590 77.475 19.460 77.645 ;
        RECT 18.950 77.385 19.460 77.475 ;
        RECT 17.500 76.920 17.805 77.050 ;
        RECT 18.250 76.940 18.780 77.305 ;
        RECT 17.120 76.325 17.385 76.785 ;
        RECT 17.555 76.495 17.805 76.920 ;
        RECT 18.950 76.770 19.120 77.385 ;
        RECT 18.015 76.600 19.120 76.770 ;
        RECT 19.290 76.325 19.460 77.125 ;
        RECT 19.630 76.825 19.800 77.895 ;
        RECT 19.970 76.995 20.160 77.715 ;
        RECT 20.330 76.965 20.650 77.925 ;
        RECT 20.820 77.965 20.990 78.425 ;
        RECT 21.265 78.345 21.475 78.875 ;
        RECT 21.735 78.135 22.065 78.660 ;
        RECT 22.235 78.265 22.405 78.875 ;
        RECT 22.575 78.220 22.905 78.655 ;
        RECT 22.575 78.135 22.955 78.220 ;
        RECT 21.865 77.965 22.065 78.135 ;
        RECT 22.730 78.095 22.955 78.135 ;
        RECT 20.820 77.635 21.695 77.965 ;
        RECT 21.865 77.635 22.615 77.965 ;
        RECT 19.630 76.495 19.880 76.825 ;
        RECT 20.820 76.795 20.990 77.635 ;
        RECT 21.865 77.430 22.055 77.635 ;
        RECT 22.785 77.515 22.955 78.095 ;
        RECT 23.125 78.105 24.795 78.875 ;
        RECT 23.125 77.585 23.875 78.105 ;
        RECT 24.965 78.055 25.225 78.875 ;
        RECT 25.395 78.055 25.725 78.475 ;
        RECT 25.905 78.305 26.165 78.705 ;
        RECT 26.335 78.475 26.665 78.875 ;
        RECT 26.835 78.305 27.005 78.655 ;
        RECT 27.175 78.475 27.550 78.875 ;
        RECT 25.905 78.135 27.570 78.305 ;
        RECT 27.740 78.200 28.015 78.545 ;
        RECT 25.475 77.965 25.725 78.055 ;
        RECT 27.400 77.965 27.570 78.135 ;
        RECT 22.740 77.465 22.955 77.515 ;
        RECT 21.160 77.055 22.055 77.430 ;
        RECT 22.565 77.385 22.955 77.465 ;
        RECT 24.045 77.415 24.795 77.935 ;
        RECT 24.970 77.635 25.305 77.885 ;
        RECT 25.475 77.635 26.190 77.965 ;
        RECT 26.405 77.635 27.230 77.965 ;
        RECT 27.400 77.635 27.675 77.965 ;
        RECT 20.105 76.625 20.990 76.795 ;
        RECT 21.170 76.325 21.485 76.825 ;
        RECT 21.715 76.495 22.055 77.055 ;
        RECT 22.225 76.325 22.395 77.335 ;
        RECT 22.565 76.540 22.895 77.385 ;
        RECT 23.125 76.325 24.795 77.415 ;
        RECT 24.965 76.325 25.225 77.465 ;
        RECT 25.475 77.075 25.645 77.635 ;
        RECT 25.905 77.175 26.235 77.465 ;
        RECT 26.405 77.345 26.650 77.635 ;
        RECT 27.400 77.465 27.570 77.635 ;
        RECT 27.845 77.465 28.015 78.200 ;
        RECT 28.735 78.325 28.905 78.615 ;
        RECT 29.075 78.495 29.405 78.875 ;
        RECT 28.735 78.155 29.400 78.325 ;
        RECT 26.910 77.295 27.570 77.465 ;
        RECT 26.910 77.175 27.080 77.295 ;
        RECT 25.905 77.005 27.080 77.175 ;
        RECT 25.465 76.505 27.080 76.835 ;
        RECT 27.250 76.325 27.530 77.125 ;
        RECT 27.740 76.495 28.015 77.465 ;
        RECT 28.650 77.335 29.000 77.985 ;
        RECT 29.170 77.165 29.400 78.155 ;
        RECT 28.735 76.995 29.400 77.165 ;
        RECT 28.735 76.495 28.905 76.995 ;
        RECT 29.075 76.325 29.405 76.825 ;
        RECT 29.575 76.495 29.760 78.615 ;
        RECT 30.015 78.415 30.265 78.875 ;
        RECT 30.435 78.425 30.770 78.595 ;
        RECT 30.965 78.425 31.640 78.595 ;
        RECT 30.435 78.285 30.605 78.425 ;
        RECT 29.930 77.295 30.210 78.245 ;
        RECT 30.380 78.155 30.605 78.285 ;
        RECT 30.380 77.050 30.550 78.155 ;
        RECT 30.775 78.005 31.300 78.225 ;
        RECT 30.720 77.240 30.960 77.835 ;
        RECT 31.130 77.305 31.300 78.005 ;
        RECT 31.470 77.645 31.640 78.425 ;
        RECT 31.960 78.375 32.330 78.875 ;
        RECT 32.510 78.425 32.915 78.595 ;
        RECT 33.085 78.425 33.870 78.595 ;
        RECT 32.510 78.195 32.680 78.425 ;
        RECT 31.850 77.895 32.680 78.195 ;
        RECT 33.065 77.925 33.530 78.255 ;
        RECT 31.850 77.865 32.050 77.895 ;
        RECT 32.170 77.645 32.340 77.715 ;
        RECT 31.470 77.475 32.340 77.645 ;
        RECT 31.830 77.385 32.340 77.475 ;
        RECT 30.380 76.920 30.685 77.050 ;
        RECT 31.130 76.940 31.660 77.305 ;
        RECT 30.000 76.325 30.265 76.785 ;
        RECT 30.435 76.495 30.685 76.920 ;
        RECT 31.830 76.770 32.000 77.385 ;
        RECT 30.895 76.600 32.000 76.770 ;
        RECT 32.170 76.325 32.340 77.125 ;
        RECT 32.510 76.825 32.680 77.895 ;
        RECT 32.850 76.995 33.040 77.715 ;
        RECT 33.210 76.965 33.530 77.925 ;
        RECT 33.700 77.965 33.870 78.425 ;
        RECT 34.145 78.345 34.355 78.875 ;
        RECT 34.615 78.135 34.945 78.660 ;
        RECT 35.115 78.265 35.285 78.875 ;
        RECT 35.455 78.220 35.785 78.655 ;
        RECT 35.955 78.360 36.125 78.875 ;
        RECT 35.455 78.135 35.835 78.220 ;
        RECT 34.745 77.965 34.945 78.135 ;
        RECT 35.610 78.095 35.835 78.135 ;
        RECT 33.700 77.635 34.575 77.965 ;
        RECT 34.745 77.635 35.495 77.965 ;
        RECT 32.510 76.495 32.760 76.825 ;
        RECT 33.700 76.795 33.870 77.635 ;
        RECT 34.745 77.430 34.935 77.635 ;
        RECT 35.665 77.515 35.835 78.095 ;
        RECT 36.465 78.105 39.055 78.875 ;
        RECT 39.225 78.150 39.515 78.875 ;
        RECT 39.775 78.325 39.945 78.615 ;
        RECT 40.115 78.495 40.445 78.875 ;
        RECT 39.775 78.155 40.440 78.325 ;
        RECT 36.465 77.585 37.675 78.105 ;
        RECT 35.620 77.465 35.835 77.515 ;
        RECT 34.040 77.055 34.935 77.430 ;
        RECT 35.445 77.385 35.835 77.465 ;
        RECT 37.845 77.415 39.055 77.935 ;
        RECT 32.985 76.625 33.870 76.795 ;
        RECT 34.050 76.325 34.365 76.825 ;
        RECT 34.595 76.495 34.935 77.055 ;
        RECT 35.105 76.325 35.275 77.335 ;
        RECT 35.445 76.540 35.775 77.385 ;
        RECT 35.945 76.325 36.115 77.240 ;
        RECT 36.465 76.325 39.055 77.415 ;
        RECT 39.225 76.325 39.515 77.490 ;
        RECT 39.690 77.335 40.040 77.985 ;
        RECT 40.210 77.165 40.440 78.155 ;
        RECT 39.775 76.995 40.440 77.165 ;
        RECT 39.775 76.495 39.945 76.995 ;
        RECT 40.115 76.325 40.445 76.825 ;
        RECT 40.615 76.495 40.800 78.615 ;
        RECT 41.055 78.415 41.305 78.875 ;
        RECT 41.475 78.425 41.810 78.595 ;
        RECT 42.005 78.425 42.680 78.595 ;
        RECT 41.475 78.285 41.645 78.425 ;
        RECT 40.970 77.295 41.250 78.245 ;
        RECT 41.420 78.155 41.645 78.285 ;
        RECT 41.420 77.050 41.590 78.155 ;
        RECT 41.815 78.005 42.340 78.225 ;
        RECT 41.760 77.240 42.000 77.835 ;
        RECT 42.170 77.305 42.340 78.005 ;
        RECT 42.510 77.645 42.680 78.425 ;
        RECT 43.000 78.375 43.370 78.875 ;
        RECT 43.550 78.425 43.955 78.595 ;
        RECT 44.125 78.425 44.910 78.595 ;
        RECT 43.550 78.195 43.720 78.425 ;
        RECT 42.890 77.895 43.720 78.195 ;
        RECT 44.105 77.925 44.570 78.255 ;
        RECT 42.890 77.865 43.090 77.895 ;
        RECT 43.210 77.645 43.380 77.715 ;
        RECT 42.510 77.475 43.380 77.645 ;
        RECT 42.870 77.385 43.380 77.475 ;
        RECT 41.420 76.920 41.725 77.050 ;
        RECT 42.170 76.940 42.700 77.305 ;
        RECT 41.040 76.325 41.305 76.785 ;
        RECT 41.475 76.495 41.725 76.920 ;
        RECT 42.870 76.770 43.040 77.385 ;
        RECT 41.935 76.600 43.040 76.770 ;
        RECT 43.210 76.325 43.380 77.125 ;
        RECT 43.550 76.825 43.720 77.895 ;
        RECT 43.890 76.995 44.080 77.715 ;
        RECT 44.250 76.965 44.570 77.925 ;
        RECT 44.740 77.965 44.910 78.425 ;
        RECT 45.185 78.345 45.395 78.875 ;
        RECT 45.655 78.135 45.985 78.660 ;
        RECT 46.155 78.265 46.325 78.875 ;
        RECT 46.495 78.220 46.825 78.655 ;
        RECT 47.555 78.220 47.885 78.655 ;
        RECT 48.055 78.265 48.225 78.875 ;
        RECT 46.495 78.135 46.875 78.220 ;
        RECT 45.785 77.965 45.985 78.135 ;
        RECT 46.650 78.095 46.875 78.135 ;
        RECT 44.740 77.635 45.615 77.965 ;
        RECT 45.785 77.635 46.535 77.965 ;
        RECT 43.550 76.495 43.800 76.825 ;
        RECT 44.740 76.795 44.910 77.635 ;
        RECT 45.785 77.430 45.975 77.635 ;
        RECT 46.705 77.515 46.875 78.095 ;
        RECT 46.660 77.465 46.875 77.515 ;
        RECT 45.080 77.055 45.975 77.430 ;
        RECT 46.485 77.385 46.875 77.465 ;
        RECT 47.505 78.135 47.885 78.220 ;
        RECT 48.395 78.135 48.725 78.660 ;
        RECT 48.985 78.345 49.195 78.875 ;
        RECT 49.470 78.425 50.255 78.595 ;
        RECT 50.425 78.425 50.830 78.595 ;
        RECT 47.505 78.095 47.730 78.135 ;
        RECT 47.505 77.515 47.675 78.095 ;
        RECT 48.395 77.965 48.595 78.135 ;
        RECT 49.470 77.965 49.640 78.425 ;
        RECT 47.845 77.635 48.595 77.965 ;
        RECT 48.765 77.635 49.640 77.965 ;
        RECT 47.505 77.465 47.720 77.515 ;
        RECT 47.505 77.385 47.895 77.465 ;
        RECT 44.025 76.625 44.910 76.795 ;
        RECT 45.090 76.325 45.405 76.825 ;
        RECT 45.635 76.495 45.975 77.055 ;
        RECT 46.145 76.325 46.315 77.335 ;
        RECT 46.485 76.540 46.815 77.385 ;
        RECT 47.565 76.540 47.895 77.385 ;
        RECT 48.405 77.430 48.595 77.635 ;
        RECT 48.065 76.325 48.235 77.335 ;
        RECT 48.405 77.055 49.300 77.430 ;
        RECT 48.405 76.495 48.745 77.055 ;
        RECT 48.975 76.325 49.290 76.825 ;
        RECT 49.470 76.795 49.640 77.635 ;
        RECT 49.810 77.925 50.275 78.255 ;
        RECT 50.660 78.195 50.830 78.425 ;
        RECT 51.010 78.375 51.380 78.875 ;
        RECT 51.700 78.425 52.375 78.595 ;
        RECT 52.570 78.425 52.905 78.595 ;
        RECT 49.810 76.965 50.130 77.925 ;
        RECT 50.660 77.895 51.490 78.195 ;
        RECT 50.300 76.995 50.490 77.715 ;
        RECT 50.660 76.825 50.830 77.895 ;
        RECT 51.290 77.865 51.490 77.895 ;
        RECT 51.000 77.645 51.170 77.715 ;
        RECT 51.700 77.645 51.870 78.425 ;
        RECT 52.735 78.285 52.905 78.425 ;
        RECT 53.075 78.415 53.325 78.875 ;
        RECT 51.000 77.475 51.870 77.645 ;
        RECT 52.040 78.005 52.565 78.225 ;
        RECT 52.735 78.155 52.960 78.285 ;
        RECT 51.000 77.385 51.510 77.475 ;
        RECT 49.470 76.625 50.355 76.795 ;
        RECT 50.580 76.495 50.830 76.825 ;
        RECT 51.000 76.325 51.170 77.125 ;
        RECT 51.340 76.770 51.510 77.385 ;
        RECT 52.040 77.305 52.210 78.005 ;
        RECT 51.680 76.940 52.210 77.305 ;
        RECT 52.380 77.240 52.620 77.835 ;
        RECT 52.790 77.050 52.960 78.155 ;
        RECT 53.130 77.295 53.410 78.245 ;
        RECT 52.655 76.920 52.960 77.050 ;
        RECT 51.340 76.600 52.445 76.770 ;
        RECT 52.655 76.495 52.905 76.920 ;
        RECT 53.075 76.325 53.340 76.785 ;
        RECT 53.580 76.495 53.765 78.615 ;
        RECT 53.935 78.495 54.265 78.875 ;
        RECT 54.435 78.325 54.605 78.615 ;
        RECT 53.940 78.155 54.605 78.325 ;
        RECT 53.940 77.165 54.170 78.155 ;
        RECT 54.865 78.105 57.455 78.875 ;
        RECT 57.675 78.220 58.005 78.655 ;
        RECT 58.175 78.265 58.345 78.875 ;
        RECT 57.625 78.135 58.005 78.220 ;
        RECT 58.515 78.135 58.845 78.660 ;
        RECT 59.105 78.345 59.315 78.875 ;
        RECT 59.590 78.425 60.375 78.595 ;
        RECT 60.545 78.425 60.950 78.595 ;
        RECT 54.340 77.335 54.690 77.985 ;
        RECT 54.865 77.585 56.075 78.105 ;
        RECT 57.625 78.095 57.850 78.135 ;
        RECT 56.245 77.415 57.455 77.935 ;
        RECT 53.940 76.995 54.605 77.165 ;
        RECT 53.935 76.325 54.265 76.825 ;
        RECT 54.435 76.495 54.605 76.995 ;
        RECT 54.865 76.325 57.455 77.415 ;
        RECT 57.625 77.515 57.795 78.095 ;
        RECT 58.515 77.965 58.715 78.135 ;
        RECT 59.590 77.965 59.760 78.425 ;
        RECT 57.965 77.635 58.715 77.965 ;
        RECT 58.885 77.635 59.760 77.965 ;
        RECT 57.625 77.465 57.840 77.515 ;
        RECT 57.625 77.385 58.015 77.465 ;
        RECT 57.685 76.540 58.015 77.385 ;
        RECT 58.525 77.430 58.715 77.635 ;
        RECT 58.185 76.325 58.355 77.335 ;
        RECT 58.525 77.055 59.420 77.430 ;
        RECT 58.525 76.495 58.865 77.055 ;
        RECT 59.095 76.325 59.410 76.825 ;
        RECT 59.590 76.795 59.760 77.635 ;
        RECT 59.930 77.925 60.395 78.255 ;
        RECT 60.780 78.195 60.950 78.425 ;
        RECT 61.130 78.375 61.500 78.875 ;
        RECT 61.820 78.425 62.495 78.595 ;
        RECT 62.690 78.425 63.025 78.595 ;
        RECT 59.930 76.965 60.250 77.925 ;
        RECT 60.780 77.895 61.610 78.195 ;
        RECT 60.420 76.995 60.610 77.715 ;
        RECT 60.780 76.825 60.950 77.895 ;
        RECT 61.410 77.865 61.610 77.895 ;
        RECT 61.120 77.645 61.290 77.715 ;
        RECT 61.820 77.645 61.990 78.425 ;
        RECT 62.855 78.285 63.025 78.425 ;
        RECT 63.195 78.415 63.445 78.875 ;
        RECT 61.120 77.475 61.990 77.645 ;
        RECT 62.160 78.005 62.685 78.225 ;
        RECT 62.855 78.155 63.080 78.285 ;
        RECT 61.120 77.385 61.630 77.475 ;
        RECT 59.590 76.625 60.475 76.795 ;
        RECT 60.700 76.495 60.950 76.825 ;
        RECT 61.120 76.325 61.290 77.125 ;
        RECT 61.460 76.770 61.630 77.385 ;
        RECT 62.160 77.305 62.330 78.005 ;
        RECT 61.800 76.940 62.330 77.305 ;
        RECT 62.500 77.240 62.740 77.835 ;
        RECT 62.910 77.050 63.080 78.155 ;
        RECT 63.250 77.295 63.530 78.245 ;
        RECT 62.775 76.920 63.080 77.050 ;
        RECT 61.460 76.600 62.565 76.770 ;
        RECT 62.775 76.495 63.025 76.920 ;
        RECT 63.195 76.325 63.460 76.785 ;
        RECT 63.700 76.495 63.885 78.615 ;
        RECT 64.055 78.495 64.385 78.875 ;
        RECT 64.555 78.325 64.725 78.615 ;
        RECT 64.060 78.155 64.725 78.325 ;
        RECT 64.060 77.165 64.290 78.155 ;
        RECT 64.985 78.150 65.275 78.875 ;
        RECT 65.445 78.135 65.885 78.695 ;
        RECT 66.055 78.135 66.505 78.875 ;
        RECT 66.675 78.305 66.845 78.705 ;
        RECT 67.015 78.475 67.435 78.875 ;
        RECT 67.605 78.305 67.835 78.705 ;
        RECT 66.675 78.135 67.835 78.305 ;
        RECT 68.005 78.135 68.495 78.705 ;
        RECT 64.460 77.335 64.810 77.985 ;
        RECT 64.060 76.995 64.725 77.165 ;
        RECT 64.055 76.325 64.385 76.825 ;
        RECT 64.555 76.495 64.725 76.995 ;
        RECT 64.985 76.325 65.275 77.490 ;
        RECT 65.445 77.125 65.755 78.135 ;
        RECT 65.925 77.515 66.095 77.965 ;
        RECT 66.265 77.685 66.655 77.965 ;
        RECT 66.840 77.635 67.085 77.965 ;
        RECT 65.925 77.345 66.715 77.515 ;
        RECT 65.445 76.495 65.885 77.125 ;
        RECT 66.060 76.325 66.375 77.175 ;
        RECT 66.545 76.665 66.715 77.345 ;
        RECT 66.885 76.835 67.085 77.635 ;
        RECT 67.285 76.835 67.535 77.965 ;
        RECT 67.750 77.635 68.155 77.965 ;
        RECT 68.325 77.465 68.495 78.135 ;
        RECT 67.725 77.295 68.495 77.465 ;
        RECT 68.675 78.150 69.005 78.660 ;
        RECT 69.175 78.475 69.505 78.875 ;
        RECT 70.555 78.305 70.885 78.645 ;
        RECT 71.055 78.475 71.385 78.875 ;
        RECT 68.675 77.515 68.865 78.150 ;
        RECT 69.175 78.135 71.540 78.305 ;
        RECT 72.825 78.145 73.115 78.875 ;
        RECT 69.175 77.965 69.345 78.135 ;
        RECT 69.035 77.635 69.345 77.965 ;
        RECT 69.515 77.635 69.820 77.965 ;
        RECT 68.675 77.385 68.895 77.515 ;
        RECT 67.725 76.665 67.975 77.295 ;
        RECT 66.545 76.495 67.975 76.665 ;
        RECT 68.155 76.325 68.485 77.125 ;
        RECT 68.675 76.535 69.005 77.385 ;
        RECT 69.175 76.325 69.425 77.465 ;
        RECT 69.605 77.305 69.820 77.635 ;
        RECT 69.995 77.305 70.280 77.965 ;
        RECT 70.475 77.305 70.740 77.965 ;
        RECT 70.955 77.305 71.200 77.965 ;
        RECT 71.370 77.135 71.540 78.135 ;
        RECT 72.815 77.635 73.115 77.965 ;
        RECT 73.295 77.945 73.525 78.585 ;
        RECT 73.705 78.325 74.015 78.695 ;
        RECT 74.195 78.505 74.865 78.875 ;
        RECT 73.705 78.125 74.935 78.325 ;
        RECT 73.295 77.635 73.820 77.945 ;
        RECT 74.000 77.635 74.465 77.945 ;
        RECT 74.645 77.455 74.935 78.125 ;
        RECT 69.615 76.965 70.905 77.135 ;
        RECT 69.615 76.545 69.865 76.965 ;
        RECT 70.095 76.325 70.425 76.795 ;
        RECT 70.655 76.545 70.905 76.965 ;
        RECT 71.085 76.965 71.540 77.135 ;
        RECT 72.825 77.215 73.985 77.455 ;
        RECT 71.085 76.535 71.415 76.965 ;
        RECT 72.825 76.505 73.085 77.215 ;
        RECT 73.255 76.325 73.585 77.035 ;
        RECT 73.755 76.505 73.985 77.215 ;
        RECT 74.165 77.235 74.935 77.455 ;
        RECT 74.165 76.505 74.435 77.235 ;
        RECT 74.615 76.325 74.955 77.055 ;
        RECT 75.125 76.505 75.385 78.695 ;
        RECT 75.585 78.145 75.875 78.875 ;
        RECT 75.575 77.635 75.875 77.965 ;
        RECT 76.055 77.945 76.285 78.585 ;
        RECT 76.465 78.325 76.775 78.695 ;
        RECT 76.955 78.505 77.625 78.875 ;
        RECT 76.465 78.125 77.695 78.325 ;
        RECT 76.055 77.635 76.580 77.945 ;
        RECT 76.760 77.635 77.225 77.945 ;
        RECT 77.405 77.455 77.695 78.125 ;
        RECT 75.585 77.215 76.745 77.455 ;
        RECT 75.585 76.505 75.845 77.215 ;
        RECT 76.015 76.325 76.345 77.035 ;
        RECT 76.515 76.505 76.745 77.215 ;
        RECT 76.925 77.235 77.695 77.455 ;
        RECT 76.925 76.505 77.195 77.235 ;
        RECT 77.375 76.325 77.715 77.055 ;
        RECT 77.885 76.505 78.145 78.695 ;
        RECT 78.325 78.105 81.835 78.875 ;
        RECT 82.005 78.125 83.215 78.875 ;
        RECT 83.390 78.135 83.645 78.705 ;
        RECT 83.815 78.475 84.145 78.875 ;
        RECT 84.570 78.340 85.100 78.705 ;
        RECT 85.290 78.535 85.565 78.705 ;
        RECT 85.285 78.365 85.565 78.535 ;
        RECT 84.570 78.305 84.745 78.340 ;
        RECT 83.815 78.135 84.745 78.305 ;
        RECT 78.325 77.585 79.975 78.105 ;
        RECT 80.145 77.415 81.835 77.935 ;
        RECT 82.005 77.585 82.525 78.125 ;
        RECT 82.695 77.415 83.215 77.955 ;
        RECT 78.325 76.325 81.835 77.415 ;
        RECT 82.005 76.325 83.215 77.415 ;
        RECT 83.390 77.465 83.560 78.135 ;
        RECT 83.815 77.965 83.985 78.135 ;
        RECT 83.730 77.635 83.985 77.965 ;
        RECT 84.210 77.635 84.405 77.965 ;
        RECT 83.390 76.495 83.725 77.465 ;
        RECT 83.895 76.325 84.065 77.465 ;
        RECT 84.235 76.665 84.405 77.635 ;
        RECT 84.575 77.005 84.745 78.135 ;
        RECT 84.915 77.345 85.085 78.145 ;
        RECT 85.290 77.545 85.565 78.365 ;
        RECT 85.735 77.345 85.925 78.705 ;
        RECT 86.105 78.340 86.615 78.875 ;
        RECT 86.835 78.065 87.080 78.670 ;
        RECT 87.615 78.325 87.785 78.705 ;
        RECT 87.965 78.495 88.295 78.875 ;
        RECT 87.615 78.155 88.280 78.325 ;
        RECT 88.475 78.200 88.735 78.705 ;
        RECT 86.125 77.895 87.355 78.065 ;
        RECT 84.915 77.175 85.925 77.345 ;
        RECT 86.095 77.330 86.845 77.520 ;
        RECT 84.575 76.835 85.700 77.005 ;
        RECT 86.095 76.665 86.265 77.330 ;
        RECT 87.015 77.085 87.355 77.895 ;
        RECT 87.545 77.605 87.875 77.975 ;
        RECT 88.110 77.900 88.280 78.155 ;
        RECT 88.110 77.570 88.395 77.900 ;
        RECT 88.110 77.425 88.280 77.570 ;
        RECT 84.235 76.495 86.265 76.665 ;
        RECT 86.435 76.325 86.605 77.085 ;
        RECT 86.840 76.675 87.355 77.085 ;
        RECT 87.615 77.255 88.280 77.425 ;
        RECT 88.565 77.400 88.735 78.200 ;
        RECT 88.905 78.105 90.575 78.875 ;
        RECT 90.745 78.125 91.955 78.875 ;
        RECT 88.905 77.585 89.655 78.105 ;
        RECT 89.825 77.415 90.575 77.935 ;
        RECT 87.615 76.495 87.785 77.255 ;
        RECT 87.965 76.325 88.295 77.085 ;
        RECT 88.465 76.495 88.735 77.400 ;
        RECT 88.905 76.325 90.575 77.415 ;
        RECT 90.745 77.415 91.265 77.955 ;
        RECT 91.435 77.585 91.955 78.125 ;
        RECT 90.745 76.325 91.955 77.415 ;
        RECT 13.380 76.155 92.040 76.325 ;
        RECT 13.465 75.065 14.675 76.155 ;
        RECT 14.845 75.065 16.515 76.155 ;
        RECT 13.465 74.355 13.985 74.895 ;
        RECT 14.155 74.525 14.675 75.065 ;
        RECT 14.845 74.375 15.595 74.895 ;
        RECT 15.765 74.545 16.515 75.065 ;
        RECT 16.720 75.365 17.255 75.985 ;
        RECT 13.465 73.605 14.675 74.355 ;
        RECT 14.845 73.605 16.515 74.375 ;
        RECT 16.720 74.345 17.035 75.365 ;
        RECT 17.425 75.355 17.755 76.155 ;
        RECT 19.445 75.645 19.705 76.155 ;
        RECT 18.240 75.185 18.630 75.360 ;
        RECT 17.205 75.015 18.630 75.185 ;
        RECT 17.205 74.515 17.375 75.015 ;
        RECT 16.720 73.775 17.335 74.345 ;
        RECT 17.625 74.285 17.890 74.845 ;
        RECT 18.060 74.115 18.230 75.015 ;
        RECT 18.400 74.285 18.755 74.845 ;
        RECT 19.445 74.595 19.785 75.475 ;
        RECT 19.955 74.765 20.125 75.985 ;
        RECT 20.365 75.650 20.980 76.155 ;
        RECT 20.365 75.115 20.615 75.480 ;
        RECT 20.785 75.475 20.980 75.650 ;
        RECT 21.150 75.645 21.625 75.985 ;
        RECT 21.795 75.610 22.010 76.155 ;
        RECT 20.785 75.285 21.115 75.475 ;
        RECT 21.335 75.115 22.050 75.410 ;
        RECT 22.220 75.285 22.495 75.985 ;
        RECT 20.365 74.945 22.155 75.115 ;
        RECT 19.955 74.515 20.750 74.765 ;
        RECT 19.955 74.425 20.205 74.515 ;
        RECT 17.505 73.605 17.720 74.115 ;
        RECT 17.950 73.785 18.230 74.115 ;
        RECT 18.410 73.605 18.650 74.115 ;
        RECT 19.445 73.605 19.705 74.425 ;
        RECT 19.875 74.005 20.205 74.425 ;
        RECT 20.920 74.090 21.175 74.945 ;
        RECT 20.385 73.825 21.175 74.090 ;
        RECT 21.345 74.245 21.755 74.765 ;
        RECT 21.925 74.515 22.155 74.945 ;
        RECT 22.325 74.255 22.495 75.285 ;
        RECT 23.125 75.015 23.385 76.155 ;
        RECT 23.625 75.645 25.240 75.975 ;
        RECT 23.635 74.845 23.805 75.405 ;
        RECT 24.065 75.305 25.240 75.475 ;
        RECT 25.410 75.355 25.690 76.155 ;
        RECT 24.065 75.015 24.395 75.305 ;
        RECT 25.070 75.185 25.240 75.305 ;
        RECT 24.565 74.845 24.810 75.135 ;
        RECT 25.070 75.015 25.730 75.185 ;
        RECT 25.900 75.015 26.175 75.985 ;
        RECT 25.560 74.845 25.730 75.015 ;
        RECT 23.130 74.595 23.465 74.845 ;
        RECT 23.635 74.515 24.350 74.845 ;
        RECT 24.565 74.515 25.390 74.845 ;
        RECT 25.560 74.515 25.835 74.845 ;
        RECT 23.635 74.425 23.885 74.515 ;
        RECT 21.345 73.825 21.545 74.245 ;
        RECT 21.735 73.605 22.065 74.065 ;
        RECT 22.235 73.775 22.495 74.255 ;
        RECT 23.125 73.605 23.385 74.425 ;
        RECT 23.555 74.005 23.885 74.425 ;
        RECT 25.560 74.345 25.730 74.515 ;
        RECT 24.065 74.175 25.730 74.345 ;
        RECT 26.005 74.280 26.175 75.015 ;
        RECT 26.345 74.990 26.635 76.155 ;
        RECT 26.805 75.065 28.475 76.155 ;
        RECT 29.195 75.485 29.365 75.985 ;
        RECT 29.535 75.655 29.865 76.155 ;
        RECT 29.195 75.315 29.860 75.485 ;
        RECT 26.805 74.375 27.555 74.895 ;
        RECT 27.725 74.545 28.475 75.065 ;
        RECT 29.110 74.495 29.460 75.145 ;
        RECT 24.065 73.775 24.325 74.175 ;
        RECT 24.495 73.605 24.825 74.005 ;
        RECT 24.995 73.825 25.165 74.175 ;
        RECT 25.335 73.605 25.710 74.005 ;
        RECT 25.900 73.935 26.175 74.280 ;
        RECT 26.345 73.605 26.635 74.330 ;
        RECT 26.805 73.605 28.475 74.375 ;
        RECT 29.630 74.325 29.860 75.315 ;
        RECT 29.195 74.155 29.860 74.325 ;
        RECT 29.195 73.865 29.365 74.155 ;
        RECT 29.535 73.605 29.865 73.985 ;
        RECT 30.035 73.865 30.220 75.985 ;
        RECT 30.460 75.695 30.725 76.155 ;
        RECT 30.895 75.560 31.145 75.985 ;
        RECT 31.355 75.710 32.460 75.880 ;
        RECT 30.840 75.430 31.145 75.560 ;
        RECT 30.390 74.235 30.670 75.185 ;
        RECT 30.840 74.325 31.010 75.430 ;
        RECT 31.180 74.645 31.420 75.240 ;
        RECT 31.590 75.175 32.120 75.540 ;
        RECT 31.590 74.475 31.760 75.175 ;
        RECT 32.290 75.095 32.460 75.710 ;
        RECT 32.630 75.355 32.800 76.155 ;
        RECT 32.970 75.655 33.220 75.985 ;
        RECT 33.445 75.685 34.330 75.855 ;
        RECT 32.290 75.005 32.800 75.095 ;
        RECT 30.840 74.195 31.065 74.325 ;
        RECT 31.235 74.255 31.760 74.475 ;
        RECT 31.930 74.835 32.800 75.005 ;
        RECT 30.475 73.605 30.725 74.065 ;
        RECT 30.895 74.055 31.065 74.195 ;
        RECT 31.930 74.055 32.100 74.835 ;
        RECT 32.630 74.765 32.800 74.835 ;
        RECT 32.310 74.585 32.510 74.615 ;
        RECT 32.970 74.585 33.140 75.655 ;
        RECT 33.310 74.765 33.500 75.485 ;
        RECT 32.310 74.285 33.140 74.585 ;
        RECT 33.670 74.555 33.990 75.515 ;
        RECT 30.895 73.885 31.230 74.055 ;
        RECT 31.425 73.885 32.100 74.055 ;
        RECT 32.420 73.605 32.790 74.105 ;
        RECT 32.970 74.055 33.140 74.285 ;
        RECT 33.525 74.225 33.990 74.555 ;
        RECT 34.160 74.845 34.330 75.685 ;
        RECT 34.510 75.655 34.825 76.155 ;
        RECT 35.055 75.425 35.395 75.985 ;
        RECT 34.500 75.050 35.395 75.425 ;
        RECT 35.565 75.145 35.735 76.155 ;
        RECT 35.205 74.845 35.395 75.050 ;
        RECT 35.905 75.095 36.235 75.940 ;
        RECT 36.405 75.240 36.575 76.155 ;
        RECT 35.905 75.015 36.295 75.095 ;
        RECT 36.925 75.065 40.435 76.155 ;
        RECT 36.080 74.965 36.295 75.015 ;
        RECT 34.160 74.515 35.035 74.845 ;
        RECT 35.205 74.515 35.955 74.845 ;
        RECT 34.160 74.055 34.330 74.515 ;
        RECT 35.205 74.345 35.405 74.515 ;
        RECT 36.125 74.385 36.295 74.965 ;
        RECT 36.070 74.345 36.295 74.385 ;
        RECT 32.970 73.885 33.375 74.055 ;
        RECT 33.545 73.885 34.330 74.055 ;
        RECT 34.605 73.605 34.815 74.135 ;
        RECT 35.075 73.820 35.405 74.345 ;
        RECT 35.915 74.260 36.295 74.345 ;
        RECT 36.925 74.375 38.575 74.895 ;
        RECT 38.745 74.545 40.435 75.065 ;
        RECT 40.675 75.150 40.930 75.955 ;
        RECT 41.100 75.320 41.360 76.155 ;
        RECT 41.530 75.150 41.790 75.955 ;
        RECT 41.960 75.320 42.215 76.155 ;
        RECT 40.675 74.980 42.275 75.150 ;
        RECT 40.605 74.585 41.825 74.810 ;
        RECT 41.995 74.415 42.275 74.980 ;
        RECT 35.575 73.605 35.745 74.215 ;
        RECT 35.915 73.825 36.245 74.260 ;
        RECT 36.415 73.605 36.585 74.120 ;
        RECT 36.925 73.605 40.435 74.375 ;
        RECT 41.545 74.245 42.275 74.415 ;
        RECT 42.450 75.015 42.785 75.985 ;
        RECT 42.955 75.015 43.125 76.155 ;
        RECT 43.295 75.815 45.325 75.985 ;
        RECT 42.450 74.345 42.620 75.015 ;
        RECT 43.295 74.845 43.465 75.815 ;
        RECT 42.790 74.515 43.045 74.845 ;
        RECT 43.270 74.515 43.465 74.845 ;
        RECT 43.635 75.475 44.760 75.645 ;
        RECT 42.875 74.345 43.045 74.515 ;
        RECT 43.635 74.345 43.805 75.475 ;
        RECT 41.080 73.605 41.375 74.130 ;
        RECT 41.545 73.800 41.770 74.245 ;
        RECT 41.940 73.605 42.270 74.075 ;
        RECT 42.450 73.775 42.705 74.345 ;
        RECT 42.875 74.175 43.805 74.345 ;
        RECT 43.975 75.135 44.985 75.305 ;
        RECT 43.975 74.335 44.145 75.135 ;
        RECT 43.630 74.140 43.805 74.175 ;
        RECT 42.875 73.605 43.205 74.005 ;
        RECT 43.630 73.775 44.160 74.140 ;
        RECT 44.350 74.115 44.625 74.935 ;
        RECT 44.345 73.945 44.625 74.115 ;
        RECT 44.350 73.775 44.625 73.945 ;
        RECT 44.795 73.775 44.985 75.135 ;
        RECT 45.155 75.150 45.325 75.815 ;
        RECT 45.495 75.395 45.665 76.155 ;
        RECT 45.900 75.395 46.415 75.805 ;
        RECT 45.155 74.960 45.905 75.150 ;
        RECT 46.075 74.585 46.415 75.395 ;
        RECT 45.185 74.415 46.415 74.585 ;
        RECT 46.590 75.015 46.925 75.985 ;
        RECT 47.095 75.015 47.265 76.155 ;
        RECT 47.435 75.815 49.465 75.985 ;
        RECT 45.165 73.605 45.675 74.140 ;
        RECT 45.895 73.810 46.140 74.415 ;
        RECT 46.590 74.345 46.760 75.015 ;
        RECT 47.435 74.845 47.605 75.815 ;
        RECT 46.930 74.515 47.185 74.845 ;
        RECT 47.410 74.515 47.605 74.845 ;
        RECT 47.775 75.475 48.900 75.645 ;
        RECT 47.015 74.345 47.185 74.515 ;
        RECT 47.775 74.345 47.945 75.475 ;
        RECT 46.590 73.775 46.845 74.345 ;
        RECT 47.015 74.175 47.945 74.345 ;
        RECT 48.115 75.135 49.125 75.305 ;
        RECT 48.115 74.335 48.285 75.135 ;
        RECT 47.770 74.140 47.945 74.175 ;
        RECT 47.015 73.605 47.345 74.005 ;
        RECT 47.770 73.775 48.300 74.140 ;
        RECT 48.490 74.115 48.765 74.935 ;
        RECT 48.485 73.945 48.765 74.115 ;
        RECT 48.490 73.775 48.765 73.945 ;
        RECT 48.935 73.775 49.125 75.135 ;
        RECT 49.295 75.150 49.465 75.815 ;
        RECT 49.635 75.395 49.805 76.155 ;
        RECT 50.040 75.395 50.555 75.805 ;
        RECT 49.295 74.960 50.045 75.150 ;
        RECT 50.215 74.585 50.555 75.395 ;
        RECT 50.725 75.065 51.935 76.155 ;
        RECT 49.325 74.415 50.555 74.585 ;
        RECT 49.305 73.605 49.815 74.140 ;
        RECT 50.035 73.810 50.280 74.415 ;
        RECT 50.725 74.355 51.245 74.895 ;
        RECT 51.415 74.525 51.935 75.065 ;
        RECT 52.105 74.990 52.395 76.155 ;
        RECT 52.570 75.015 52.905 75.985 ;
        RECT 53.075 75.015 53.245 76.155 ;
        RECT 53.415 75.815 55.445 75.985 ;
        RECT 50.725 73.605 51.935 74.355 ;
        RECT 52.570 74.345 52.740 75.015 ;
        RECT 53.415 74.845 53.585 75.815 ;
        RECT 52.910 74.515 53.165 74.845 ;
        RECT 53.390 74.515 53.585 74.845 ;
        RECT 53.755 75.475 54.880 75.645 ;
        RECT 52.995 74.345 53.165 74.515 ;
        RECT 53.755 74.345 53.925 75.475 ;
        RECT 52.105 73.605 52.395 74.330 ;
        RECT 52.570 73.775 52.825 74.345 ;
        RECT 52.995 74.175 53.925 74.345 ;
        RECT 54.095 75.135 55.105 75.305 ;
        RECT 54.095 74.335 54.265 75.135 ;
        RECT 53.750 74.140 53.925 74.175 ;
        RECT 52.995 73.605 53.325 74.005 ;
        RECT 53.750 73.775 54.280 74.140 ;
        RECT 54.470 74.115 54.745 74.935 ;
        RECT 54.465 73.945 54.745 74.115 ;
        RECT 54.470 73.775 54.745 73.945 ;
        RECT 54.915 73.775 55.105 75.135 ;
        RECT 55.275 75.150 55.445 75.815 ;
        RECT 55.615 75.395 55.785 76.155 ;
        RECT 56.020 75.395 56.535 75.805 ;
        RECT 55.275 74.960 56.025 75.150 ;
        RECT 56.195 74.585 56.535 75.395 ;
        RECT 57.225 75.095 57.555 75.940 ;
        RECT 57.725 75.145 57.895 76.155 ;
        RECT 58.065 75.425 58.405 75.985 ;
        RECT 58.635 75.655 58.950 76.155 ;
        RECT 59.130 75.685 60.015 75.855 ;
        RECT 55.305 74.415 56.535 74.585 ;
        RECT 57.165 75.015 57.555 75.095 ;
        RECT 58.065 75.050 58.960 75.425 ;
        RECT 57.165 74.965 57.380 75.015 ;
        RECT 55.285 73.605 55.795 74.140 ;
        RECT 56.015 73.810 56.260 74.415 ;
        RECT 57.165 74.385 57.335 74.965 ;
        RECT 58.065 74.845 58.255 75.050 ;
        RECT 59.130 74.845 59.300 75.685 ;
        RECT 60.240 75.655 60.490 75.985 ;
        RECT 57.505 74.515 58.255 74.845 ;
        RECT 58.425 74.515 59.300 74.845 ;
        RECT 57.165 74.345 57.390 74.385 ;
        RECT 58.055 74.345 58.255 74.515 ;
        RECT 57.165 74.260 57.545 74.345 ;
        RECT 57.215 73.825 57.545 74.260 ;
        RECT 57.715 73.605 57.885 74.215 ;
        RECT 58.055 73.820 58.385 74.345 ;
        RECT 58.645 73.605 58.855 74.135 ;
        RECT 59.130 74.055 59.300 74.515 ;
        RECT 59.470 74.555 59.790 75.515 ;
        RECT 59.960 74.765 60.150 75.485 ;
        RECT 60.320 74.585 60.490 75.655 ;
        RECT 60.660 75.355 60.830 76.155 ;
        RECT 61.000 75.710 62.105 75.880 ;
        RECT 61.000 75.095 61.170 75.710 ;
        RECT 62.315 75.560 62.565 75.985 ;
        RECT 62.735 75.695 63.000 76.155 ;
        RECT 61.340 75.175 61.870 75.540 ;
        RECT 62.315 75.430 62.620 75.560 ;
        RECT 60.660 75.005 61.170 75.095 ;
        RECT 60.660 74.835 61.530 75.005 ;
        RECT 60.660 74.765 60.830 74.835 ;
        RECT 60.950 74.585 61.150 74.615 ;
        RECT 59.470 74.225 59.935 74.555 ;
        RECT 60.320 74.285 61.150 74.585 ;
        RECT 60.320 74.055 60.490 74.285 ;
        RECT 59.130 73.885 59.915 74.055 ;
        RECT 60.085 73.885 60.490 74.055 ;
        RECT 60.670 73.605 61.040 74.105 ;
        RECT 61.360 74.055 61.530 74.835 ;
        RECT 61.700 74.475 61.870 75.175 ;
        RECT 62.040 74.645 62.280 75.240 ;
        RECT 61.700 74.255 62.225 74.475 ;
        RECT 62.450 74.325 62.620 75.430 ;
        RECT 62.395 74.195 62.620 74.325 ;
        RECT 62.790 74.235 63.070 75.185 ;
        RECT 62.395 74.055 62.565 74.195 ;
        RECT 61.360 73.885 62.035 74.055 ;
        RECT 62.230 73.885 62.565 74.055 ;
        RECT 62.735 73.605 62.985 74.065 ;
        RECT 63.240 73.865 63.425 75.985 ;
        RECT 63.595 75.655 63.925 76.155 ;
        RECT 64.095 75.485 64.265 75.985 ;
        RECT 63.600 75.315 64.265 75.485 ;
        RECT 64.640 75.525 64.925 75.985 ;
        RECT 65.095 75.695 65.365 76.155 ;
        RECT 63.600 74.325 63.830 75.315 ;
        RECT 64.640 75.305 65.595 75.525 ;
        RECT 64.000 74.495 64.350 75.145 ;
        RECT 64.525 74.575 65.215 75.135 ;
        RECT 65.385 74.405 65.595 75.305 ;
        RECT 63.600 74.155 64.265 74.325 ;
        RECT 63.595 73.605 63.925 73.985 ;
        RECT 64.095 73.865 64.265 74.155 ;
        RECT 64.640 74.235 65.595 74.405 ;
        RECT 65.765 75.135 66.165 75.985 ;
        RECT 66.355 75.525 66.635 75.985 ;
        RECT 67.155 75.695 67.480 76.155 ;
        RECT 66.355 75.305 67.480 75.525 ;
        RECT 65.765 74.575 66.860 75.135 ;
        RECT 67.030 74.845 67.480 75.305 ;
        RECT 67.650 75.015 68.035 75.985 ;
        RECT 64.640 73.775 64.925 74.235 ;
        RECT 65.095 73.605 65.365 74.065 ;
        RECT 65.765 73.775 66.165 74.575 ;
        RECT 67.030 74.515 67.585 74.845 ;
        RECT 67.030 74.405 67.480 74.515 ;
        RECT 66.355 74.235 67.480 74.405 ;
        RECT 67.755 74.345 68.035 75.015 ;
        RECT 66.355 73.775 66.635 74.235 ;
        RECT 67.155 73.605 67.480 74.065 ;
        RECT 67.650 73.775 68.035 74.345 ;
        RECT 68.205 73.885 68.485 75.985 ;
        RECT 68.675 75.395 69.460 76.155 ;
        RECT 69.855 75.325 70.240 75.985 ;
        RECT 69.855 75.225 70.265 75.325 ;
        RECT 68.655 75.015 70.265 75.225 ;
        RECT 70.565 75.135 70.765 75.925 ;
        RECT 68.655 74.415 68.930 75.015 ;
        RECT 70.435 74.965 70.765 75.135 ;
        RECT 70.935 74.975 71.255 76.155 ;
        RECT 71.625 75.485 71.905 76.155 ;
        RECT 72.075 75.265 72.375 75.815 ;
        RECT 72.575 75.435 72.905 76.155 ;
        RECT 73.095 75.435 73.555 75.985 ;
        RECT 70.435 74.845 70.615 74.965 ;
        RECT 69.100 74.595 69.455 74.845 ;
        RECT 69.650 74.795 70.115 74.845 ;
        RECT 69.645 74.625 70.115 74.795 ;
        RECT 69.650 74.595 70.115 74.625 ;
        RECT 70.285 74.595 70.615 74.845 ;
        RECT 71.440 74.845 71.705 75.205 ;
        RECT 72.075 75.095 73.015 75.265 ;
        RECT 72.845 74.845 73.015 75.095 ;
        RECT 70.790 74.595 71.255 74.795 ;
        RECT 71.440 74.595 72.115 74.845 ;
        RECT 72.335 74.595 72.675 74.845 ;
        RECT 72.845 74.515 73.135 74.845 ;
        RECT 72.845 74.425 73.015 74.515 ;
        RECT 68.655 74.235 69.905 74.415 ;
        RECT 69.540 74.165 69.905 74.235 ;
        RECT 70.075 74.215 71.255 74.385 ;
        RECT 68.715 73.605 68.885 74.065 ;
        RECT 70.075 73.995 70.405 74.215 ;
        RECT 69.155 73.815 70.405 73.995 ;
        RECT 70.575 73.605 70.745 74.045 ;
        RECT 70.915 73.800 71.255 74.215 ;
        RECT 71.625 74.235 73.015 74.425 ;
        RECT 71.625 73.875 71.955 74.235 ;
        RECT 73.305 74.065 73.555 75.435 ;
        RECT 73.725 75.015 73.985 76.155 ;
        RECT 74.155 75.005 74.485 75.985 ;
        RECT 74.655 75.015 74.935 76.155 ;
        RECT 75.655 75.225 75.825 75.985 ;
        RECT 76.040 75.395 76.370 76.155 ;
        RECT 75.655 75.055 76.370 75.225 ;
        RECT 76.540 75.080 76.795 75.985 ;
        RECT 73.745 74.595 74.080 74.845 ;
        RECT 74.250 74.405 74.420 75.005 ;
        RECT 74.590 74.575 74.925 74.845 ;
        RECT 75.565 74.505 75.920 74.875 ;
        RECT 76.200 74.845 76.370 75.055 ;
        RECT 76.200 74.515 76.455 74.845 ;
        RECT 72.575 73.605 72.825 74.065 ;
        RECT 72.995 73.775 73.555 74.065 ;
        RECT 73.725 73.775 74.420 74.405 ;
        RECT 74.625 73.605 74.935 74.405 ;
        RECT 76.200 74.325 76.370 74.515 ;
        RECT 76.625 74.350 76.795 75.080 ;
        RECT 76.970 75.005 77.230 76.155 ;
        RECT 77.865 74.990 78.155 76.155 ;
        RECT 78.325 75.065 80.915 76.155 ;
        RECT 81.635 75.485 81.805 75.985 ;
        RECT 81.975 75.655 82.305 76.155 ;
        RECT 81.635 75.315 82.300 75.485 ;
        RECT 75.655 74.155 76.370 74.325 ;
        RECT 75.655 73.775 75.825 74.155 ;
        RECT 76.040 73.605 76.370 73.985 ;
        RECT 76.540 73.775 76.795 74.350 ;
        RECT 76.970 73.605 77.230 74.445 ;
        RECT 78.325 74.375 79.535 74.895 ;
        RECT 79.705 74.545 80.915 75.065 ;
        RECT 81.550 74.495 81.900 75.145 ;
        RECT 77.865 73.605 78.155 74.330 ;
        RECT 78.325 73.605 80.915 74.375 ;
        RECT 82.070 74.325 82.300 75.315 ;
        RECT 81.635 74.155 82.300 74.325 ;
        RECT 81.635 73.865 81.805 74.155 ;
        RECT 81.975 73.605 82.305 73.985 ;
        RECT 82.475 73.865 82.660 75.985 ;
        RECT 82.900 75.695 83.165 76.155 ;
        RECT 83.335 75.560 83.585 75.985 ;
        RECT 83.795 75.710 84.900 75.880 ;
        RECT 83.280 75.430 83.585 75.560 ;
        RECT 82.830 74.235 83.110 75.185 ;
        RECT 83.280 74.325 83.450 75.430 ;
        RECT 83.620 74.645 83.860 75.240 ;
        RECT 84.030 75.175 84.560 75.540 ;
        RECT 84.030 74.475 84.200 75.175 ;
        RECT 84.730 75.095 84.900 75.710 ;
        RECT 85.070 75.355 85.240 76.155 ;
        RECT 85.410 75.655 85.660 75.985 ;
        RECT 85.885 75.685 86.770 75.855 ;
        RECT 84.730 75.005 85.240 75.095 ;
        RECT 83.280 74.195 83.505 74.325 ;
        RECT 83.675 74.255 84.200 74.475 ;
        RECT 84.370 74.835 85.240 75.005 ;
        RECT 82.915 73.605 83.165 74.065 ;
        RECT 83.335 74.055 83.505 74.195 ;
        RECT 84.370 74.055 84.540 74.835 ;
        RECT 85.070 74.765 85.240 74.835 ;
        RECT 84.750 74.585 84.950 74.615 ;
        RECT 85.410 74.585 85.580 75.655 ;
        RECT 85.750 74.765 85.940 75.485 ;
        RECT 84.750 74.285 85.580 74.585 ;
        RECT 86.110 74.555 86.430 75.515 ;
        RECT 83.335 73.885 83.670 74.055 ;
        RECT 83.865 73.885 84.540 74.055 ;
        RECT 84.860 73.605 85.230 74.105 ;
        RECT 85.410 74.055 85.580 74.285 ;
        RECT 85.965 74.225 86.430 74.555 ;
        RECT 86.600 74.845 86.770 75.685 ;
        RECT 86.950 75.655 87.265 76.155 ;
        RECT 87.495 75.425 87.835 75.985 ;
        RECT 86.940 75.050 87.835 75.425 ;
        RECT 88.005 75.145 88.175 76.155 ;
        RECT 87.645 74.845 87.835 75.050 ;
        RECT 88.345 75.095 88.675 75.940 ;
        RECT 88.995 75.225 89.165 75.985 ;
        RECT 89.380 75.395 89.710 76.155 ;
        RECT 88.345 75.015 88.735 75.095 ;
        RECT 88.995 75.055 89.710 75.225 ;
        RECT 89.880 75.080 90.135 75.985 ;
        RECT 88.520 74.965 88.735 75.015 ;
        RECT 86.600 74.515 87.475 74.845 ;
        RECT 87.645 74.515 88.395 74.845 ;
        RECT 86.600 74.055 86.770 74.515 ;
        RECT 87.645 74.345 87.845 74.515 ;
        RECT 88.565 74.385 88.735 74.965 ;
        RECT 88.905 74.505 89.260 74.875 ;
        RECT 89.540 74.845 89.710 75.055 ;
        RECT 89.540 74.515 89.795 74.845 ;
        RECT 88.510 74.345 88.735 74.385 ;
        RECT 85.410 73.885 85.815 74.055 ;
        RECT 85.985 73.885 86.770 74.055 ;
        RECT 87.045 73.605 87.255 74.135 ;
        RECT 87.515 73.820 87.845 74.345 ;
        RECT 88.355 74.260 88.735 74.345 ;
        RECT 89.540 74.325 89.710 74.515 ;
        RECT 89.965 74.350 90.135 75.080 ;
        RECT 90.310 75.005 90.570 76.155 ;
        RECT 90.745 75.065 91.955 76.155 ;
        RECT 99.990 75.105 100.160 80.925 ;
        RECT 100.640 78.285 100.990 80.445 ;
        RECT 100.640 75.585 100.990 77.745 ;
        RECT 101.470 75.105 101.640 80.925 ;
        RECT 102.120 78.285 102.470 80.445 ;
        RECT 102.120 75.585 102.470 77.745 ;
        RECT 102.950 75.105 103.120 80.925 ;
        RECT 103.600 78.285 103.950 80.445 ;
        RECT 103.600 75.585 103.950 77.745 ;
        RECT 104.430 75.105 104.600 80.925 ;
        RECT 105.080 78.285 105.430 80.445 ;
        RECT 105.080 75.585 105.430 77.745 ;
        RECT 105.910 75.105 106.080 80.925 ;
        RECT 106.560 78.285 106.910 80.445 ;
        RECT 106.560 75.585 106.910 77.745 ;
        RECT 107.390 75.105 107.560 80.925 ;
        RECT 108.040 78.285 108.390 80.445 ;
        RECT 108.040 75.585 108.390 77.745 ;
        RECT 108.870 75.105 109.040 80.925 ;
        RECT 109.520 78.285 109.870 80.445 ;
        RECT 109.520 75.585 109.870 77.745 ;
        RECT 110.350 75.105 110.520 80.925 ;
        RECT 117.600 80.850 129.140 81.010 ;
        RECT 117.600 80.840 127.560 80.850 ;
        RECT 117.600 75.450 117.770 80.840 ;
        RECT 118.400 80.330 119.400 80.500 ;
        RECT 118.170 76.120 118.340 80.160 ;
        RECT 119.460 76.120 119.630 80.160 ;
        RECT 118.400 75.780 119.400 75.950 ;
        RECT 120.030 75.450 120.200 80.840 ;
        RECT 120.830 80.330 122.830 80.500 ;
        RECT 120.600 76.120 120.770 80.160 ;
        RECT 122.890 76.120 123.060 80.160 ;
        RECT 120.830 75.780 122.830 75.950 ;
        RECT 123.460 75.450 123.630 80.840 ;
        RECT 124.260 80.330 126.260 80.500 ;
        RECT 124.030 76.120 124.200 80.160 ;
        RECT 126.320 76.120 126.490 80.160 ;
        RECT 126.890 79.940 127.560 80.840 ;
        RECT 128.100 80.340 128.430 80.510 ;
        RECT 126.890 78.760 127.580 79.940 ;
        RECT 127.960 79.130 128.130 80.170 ;
        RECT 128.400 79.130 128.570 80.170 ;
        RECT 128.970 78.760 129.140 80.850 ;
        RECT 129.450 80.960 130.470 81.350 ;
        RECT 129.450 80.820 131.250 80.960 ;
        RECT 126.890 78.590 129.140 78.760 ;
        RECT 129.500 80.790 131.250 80.820 ;
        RECT 129.500 80.780 130.470 80.790 ;
        RECT 126.890 78.430 128.750 78.590 ;
        RECT 126.890 78.200 127.660 78.430 ;
        RECT 126.890 76.690 127.650 78.200 ;
        RECT 124.260 75.780 126.260 75.950 ;
        RECT 126.890 75.450 128.920 76.690 ;
        RECT 129.500 76.650 129.670 80.780 ;
        RECT 130.210 80.275 130.540 80.445 ;
        RECT 130.070 77.020 130.240 80.060 ;
        RECT 130.510 77.020 130.680 80.060 ;
        RECT 131.080 76.650 131.250 80.790 ;
        RECT 134.420 79.150 134.590 84.540 ;
        RECT 135.130 84.130 135.460 84.300 ;
        RECT 134.990 79.875 135.160 83.915 ;
        RECT 135.430 79.875 135.600 83.915 ;
        RECT 135.130 79.490 135.460 79.660 ;
        RECT 136.000 79.150 136.170 84.540 ;
        RECT 139.540 84.540 139.730 84.640 ;
        RECT 137.210 84.130 137.540 84.300 ;
        RECT 138.170 84.130 138.500 84.300 ;
        RECT 136.570 79.875 136.740 83.915 ;
        RECT 137.050 79.875 137.220 83.915 ;
        RECT 137.530 79.875 137.700 83.915 ;
        RECT 138.010 79.875 138.180 83.915 ;
        RECT 138.490 79.875 138.660 83.915 ;
        RECT 138.970 79.875 139.140 83.915 ;
        RECT 136.730 79.490 137.060 79.660 ;
        RECT 137.690 79.490 138.020 79.660 ;
        RECT 138.650 79.490 138.980 79.660 ;
        RECT 139.540 79.150 139.710 84.540 ;
        RECT 134.420 78.980 139.710 79.150 ;
        RECT 129.500 76.480 131.250 76.650 ;
        RECT 134.410 78.090 139.700 78.260 ;
        RECT 134.410 75.690 134.580 78.090 ;
        RECT 135.120 77.580 135.450 77.750 ;
        RECT 134.980 76.370 135.150 77.410 ;
        RECT 135.420 76.370 135.590 77.410 ;
        RECT 135.120 76.030 135.450 76.200 ;
        RECT 135.990 75.690 136.160 78.090 ;
        RECT 137.200 77.580 137.530 77.750 ;
        RECT 138.160 77.580 138.490 77.750 ;
        RECT 136.560 76.370 136.730 77.410 ;
        RECT 137.040 76.370 137.210 77.410 ;
        RECT 137.520 76.370 137.690 77.410 ;
        RECT 138.000 76.370 138.170 77.410 ;
        RECT 138.480 76.370 138.650 77.410 ;
        RECT 138.960 76.370 139.130 77.410 ;
        RECT 136.720 76.030 137.050 76.200 ;
        RECT 137.680 76.030 138.010 76.200 ;
        RECT 138.640 76.030 138.970 76.200 ;
        RECT 139.530 75.690 139.700 78.090 ;
        RECT 134.410 75.520 139.700 75.690 ;
        RECT 117.600 75.270 128.920 75.450 ;
        RECT 90.745 74.525 91.265 75.065 ;
        RECT 99.990 74.935 110.520 75.105 ;
        RECT 88.015 73.605 88.185 74.215 ;
        RECT 88.355 73.825 88.685 74.260 ;
        RECT 88.995 74.155 89.710 74.325 ;
        RECT 88.995 73.775 89.165 74.155 ;
        RECT 89.380 73.605 89.710 73.985 ;
        RECT 89.880 73.775 90.135 74.350 ;
        RECT 90.310 73.605 90.570 74.445 ;
        RECT 91.435 74.355 91.955 74.895 ;
        RECT 117.610 74.780 128.920 75.270 ;
        RECT 127.000 74.770 128.920 74.780 ;
        RECT 134.420 74.690 139.700 75.520 ;
        RECT 90.745 73.605 91.955 74.355 ;
        RECT 13.380 73.435 92.040 73.605 ;
        RECT 13.465 72.685 14.675 73.435 ;
        RECT 15.310 72.695 15.565 73.265 ;
        RECT 15.735 73.035 16.065 73.435 ;
        RECT 16.490 72.900 17.020 73.265 ;
        RECT 16.490 72.865 16.665 72.900 ;
        RECT 15.735 72.695 16.665 72.865 ;
        RECT 13.465 72.145 13.985 72.685 ;
        RECT 14.155 71.975 14.675 72.515 ;
        RECT 13.465 70.885 14.675 71.975 ;
        RECT 15.310 72.025 15.480 72.695 ;
        RECT 15.735 72.525 15.905 72.695 ;
        RECT 15.650 72.195 15.905 72.525 ;
        RECT 16.130 72.195 16.325 72.525 ;
        RECT 15.310 71.055 15.645 72.025 ;
        RECT 15.815 70.885 15.985 72.025 ;
        RECT 16.155 71.225 16.325 72.195 ;
        RECT 16.495 71.565 16.665 72.695 ;
        RECT 16.835 71.905 17.005 72.705 ;
        RECT 17.210 72.415 17.485 73.265 ;
        RECT 17.205 72.245 17.485 72.415 ;
        RECT 17.210 72.105 17.485 72.245 ;
        RECT 17.655 71.905 17.845 73.265 ;
        RECT 18.025 72.900 18.535 73.435 ;
        RECT 18.755 72.625 19.000 73.230 ;
        RECT 19.450 72.695 19.705 73.265 ;
        RECT 19.875 73.035 20.205 73.435 ;
        RECT 20.630 72.900 21.160 73.265 ;
        RECT 20.630 72.865 20.805 72.900 ;
        RECT 19.875 72.695 20.805 72.865 ;
        RECT 18.045 72.455 19.275 72.625 ;
        RECT 16.835 71.735 17.845 71.905 ;
        RECT 18.015 71.890 18.765 72.080 ;
        RECT 16.495 71.395 17.620 71.565 ;
        RECT 18.015 71.225 18.185 71.890 ;
        RECT 18.935 71.645 19.275 72.455 ;
        RECT 16.155 71.055 18.185 71.225 ;
        RECT 18.355 70.885 18.525 71.645 ;
        RECT 18.760 71.235 19.275 71.645 ;
        RECT 19.450 72.025 19.620 72.695 ;
        RECT 19.875 72.525 20.045 72.695 ;
        RECT 19.790 72.195 20.045 72.525 ;
        RECT 20.270 72.195 20.465 72.525 ;
        RECT 19.450 71.055 19.785 72.025 ;
        RECT 19.955 70.885 20.125 72.025 ;
        RECT 20.295 71.225 20.465 72.195 ;
        RECT 20.635 71.565 20.805 72.695 ;
        RECT 20.975 71.905 21.145 72.705 ;
        RECT 21.350 72.415 21.625 73.265 ;
        RECT 21.345 72.245 21.625 72.415 ;
        RECT 21.350 72.105 21.625 72.245 ;
        RECT 21.795 71.905 21.985 73.265 ;
        RECT 22.165 72.900 22.675 73.435 ;
        RECT 22.895 72.625 23.140 73.230 ;
        RECT 24.780 72.625 25.025 73.230 ;
        RECT 25.245 72.900 25.755 73.435 ;
        RECT 22.185 72.455 23.415 72.625 ;
        RECT 20.975 71.735 21.985 71.905 ;
        RECT 22.155 71.890 22.905 72.080 ;
        RECT 20.635 71.395 21.760 71.565 ;
        RECT 22.155 71.225 22.325 71.890 ;
        RECT 23.075 71.645 23.415 72.455 ;
        RECT 20.295 71.055 22.325 71.225 ;
        RECT 22.495 70.885 22.665 71.645 ;
        RECT 22.900 71.235 23.415 71.645 ;
        RECT 24.505 72.455 25.735 72.625 ;
        RECT 24.505 71.645 24.845 72.455 ;
        RECT 25.015 71.890 25.765 72.080 ;
        RECT 24.505 71.235 25.020 71.645 ;
        RECT 25.255 70.885 25.425 71.645 ;
        RECT 25.595 71.225 25.765 71.890 ;
        RECT 25.935 71.905 26.125 73.265 ;
        RECT 26.295 73.095 26.570 73.265 ;
        RECT 26.295 72.925 26.575 73.095 ;
        RECT 26.295 72.105 26.570 72.925 ;
        RECT 26.760 72.900 27.290 73.265 ;
        RECT 27.715 73.035 28.045 73.435 ;
        RECT 27.115 72.865 27.290 72.900 ;
        RECT 26.775 71.905 26.945 72.705 ;
        RECT 25.935 71.735 26.945 71.905 ;
        RECT 27.115 72.695 28.045 72.865 ;
        RECT 28.215 72.695 28.470 73.265 ;
        RECT 28.705 72.975 28.950 73.435 ;
        RECT 27.115 71.565 27.285 72.695 ;
        RECT 27.875 72.525 28.045 72.695 ;
        RECT 26.160 71.395 27.285 71.565 ;
        RECT 27.455 72.195 27.650 72.525 ;
        RECT 27.875 72.195 28.130 72.525 ;
        RECT 27.455 71.225 27.625 72.195 ;
        RECT 28.300 72.025 28.470 72.695 ;
        RECT 28.645 72.195 28.960 72.805 ;
        RECT 29.130 72.445 29.380 73.255 ;
        RECT 29.550 72.910 29.810 73.435 ;
        RECT 29.980 72.785 30.240 73.240 ;
        RECT 30.410 72.955 30.670 73.435 ;
        RECT 30.840 72.785 31.100 73.240 ;
        RECT 31.270 72.955 31.530 73.435 ;
        RECT 31.700 72.785 31.960 73.240 ;
        RECT 32.130 72.955 32.390 73.435 ;
        RECT 32.560 72.785 32.820 73.240 ;
        RECT 32.990 72.955 33.290 73.435 ;
        RECT 33.705 72.890 39.050 73.435 ;
        RECT 29.980 72.615 33.290 72.785 ;
        RECT 29.130 72.195 32.150 72.445 ;
        RECT 25.595 71.055 27.625 71.225 ;
        RECT 27.795 70.885 27.965 72.025 ;
        RECT 28.135 71.055 28.470 72.025 ;
        RECT 28.655 70.885 28.950 71.995 ;
        RECT 29.130 71.060 29.380 72.195 ;
        RECT 32.320 72.025 33.290 72.615 ;
        RECT 35.290 72.060 35.630 72.890 ;
        RECT 39.225 72.710 39.515 73.435 ;
        RECT 40.665 72.975 40.910 73.435 ;
        RECT 29.550 70.885 29.810 71.995 ;
        RECT 29.980 71.785 33.290 72.025 ;
        RECT 29.980 71.060 30.240 71.785 ;
        RECT 30.410 70.885 30.670 71.615 ;
        RECT 30.840 71.060 31.100 71.785 ;
        RECT 31.270 70.885 31.530 71.615 ;
        RECT 31.700 71.060 31.960 71.785 ;
        RECT 32.130 70.885 32.390 71.615 ;
        RECT 32.560 71.060 32.820 71.785 ;
        RECT 32.990 70.885 33.285 71.615 ;
        RECT 37.110 71.320 37.460 72.570 ;
        RECT 40.605 72.195 40.920 72.805 ;
        RECT 41.090 72.445 41.340 73.255 ;
        RECT 41.510 72.910 41.770 73.435 ;
        RECT 41.940 72.785 42.200 73.240 ;
        RECT 42.370 72.955 42.630 73.435 ;
        RECT 42.800 72.785 43.060 73.240 ;
        RECT 43.230 72.955 43.490 73.435 ;
        RECT 43.660 72.785 43.920 73.240 ;
        RECT 44.090 72.955 44.350 73.435 ;
        RECT 44.520 72.785 44.780 73.240 ;
        RECT 44.950 72.955 45.250 73.435 ;
        RECT 41.940 72.615 45.250 72.785 ;
        RECT 41.090 72.195 44.110 72.445 ;
        RECT 33.705 70.885 39.050 71.320 ;
        RECT 39.225 70.885 39.515 72.050 ;
        RECT 40.615 70.885 40.910 71.995 ;
        RECT 41.090 71.060 41.340 72.195 ;
        RECT 44.280 72.025 45.250 72.615 ;
        RECT 45.665 72.665 48.255 73.435 ;
        RECT 48.515 72.885 48.685 73.175 ;
        RECT 48.855 73.055 49.185 73.435 ;
        RECT 48.515 72.715 49.180 72.885 ;
        RECT 45.665 72.145 46.875 72.665 ;
        RECT 41.510 70.885 41.770 71.995 ;
        RECT 41.940 71.785 45.250 72.025 ;
        RECT 47.045 71.975 48.255 72.495 ;
        RECT 41.940 71.060 42.200 71.785 ;
        RECT 42.370 70.885 42.630 71.615 ;
        RECT 42.800 71.060 43.060 71.785 ;
        RECT 43.230 70.885 43.490 71.615 ;
        RECT 43.660 71.060 43.920 71.785 ;
        RECT 44.090 70.885 44.350 71.615 ;
        RECT 44.520 71.060 44.780 71.785 ;
        RECT 44.950 70.885 45.245 71.615 ;
        RECT 45.665 70.885 48.255 71.975 ;
        RECT 48.430 71.895 48.780 72.545 ;
        RECT 48.950 71.725 49.180 72.715 ;
        RECT 48.515 71.555 49.180 71.725 ;
        RECT 48.515 71.055 48.685 71.555 ;
        RECT 48.855 70.885 49.185 71.385 ;
        RECT 49.355 71.055 49.540 73.175 ;
        RECT 49.795 72.975 50.045 73.435 ;
        RECT 50.215 72.985 50.550 73.155 ;
        RECT 50.745 72.985 51.420 73.155 ;
        RECT 50.215 72.845 50.385 72.985 ;
        RECT 49.710 71.855 49.990 72.805 ;
        RECT 50.160 72.715 50.385 72.845 ;
        RECT 50.160 71.610 50.330 72.715 ;
        RECT 50.555 72.565 51.080 72.785 ;
        RECT 50.500 71.800 50.740 72.395 ;
        RECT 50.910 71.865 51.080 72.565 ;
        RECT 51.250 72.205 51.420 72.985 ;
        RECT 51.740 72.935 52.110 73.435 ;
        RECT 52.290 72.985 52.695 73.155 ;
        RECT 52.865 72.985 53.650 73.155 ;
        RECT 52.290 72.755 52.460 72.985 ;
        RECT 51.630 72.455 52.460 72.755 ;
        RECT 52.845 72.485 53.310 72.815 ;
        RECT 51.630 72.425 51.830 72.455 ;
        RECT 51.950 72.205 52.120 72.275 ;
        RECT 51.250 72.035 52.120 72.205 ;
        RECT 51.610 71.945 52.120 72.035 ;
        RECT 50.160 71.480 50.465 71.610 ;
        RECT 50.910 71.500 51.440 71.865 ;
        RECT 49.780 70.885 50.045 71.345 ;
        RECT 50.215 71.055 50.465 71.480 ;
        RECT 51.610 71.330 51.780 71.945 ;
        RECT 50.675 71.160 51.780 71.330 ;
        RECT 51.950 70.885 52.120 71.685 ;
        RECT 52.290 71.385 52.460 72.455 ;
        RECT 52.630 71.555 52.820 72.275 ;
        RECT 52.990 71.525 53.310 72.485 ;
        RECT 53.480 72.525 53.650 72.985 ;
        RECT 53.925 72.905 54.135 73.435 ;
        RECT 54.395 72.695 54.725 73.220 ;
        RECT 54.895 72.825 55.065 73.435 ;
        RECT 55.235 72.780 55.565 73.215 ;
        RECT 55.235 72.695 55.615 72.780 ;
        RECT 54.525 72.525 54.725 72.695 ;
        RECT 55.390 72.655 55.615 72.695 ;
        RECT 53.480 72.195 54.355 72.525 ;
        RECT 54.525 72.195 55.275 72.525 ;
        RECT 52.290 71.055 52.540 71.385 ;
        RECT 53.480 71.355 53.650 72.195 ;
        RECT 54.525 71.990 54.715 72.195 ;
        RECT 55.445 72.075 55.615 72.655 ;
        RECT 55.400 72.025 55.615 72.075 ;
        RECT 53.820 71.615 54.715 71.990 ;
        RECT 55.225 71.945 55.615 72.025 ;
        RECT 55.790 72.695 56.045 73.265 ;
        RECT 56.215 73.035 56.545 73.435 ;
        RECT 56.970 72.900 57.500 73.265 ;
        RECT 56.970 72.865 57.145 72.900 ;
        RECT 56.215 72.695 57.145 72.865 ;
        RECT 55.790 72.025 55.960 72.695 ;
        RECT 56.215 72.525 56.385 72.695 ;
        RECT 56.130 72.195 56.385 72.525 ;
        RECT 56.610 72.195 56.805 72.525 ;
        RECT 52.765 71.185 53.650 71.355 ;
        RECT 53.830 70.885 54.145 71.385 ;
        RECT 54.375 71.055 54.715 71.615 ;
        RECT 54.885 70.885 55.055 71.895 ;
        RECT 55.225 71.100 55.555 71.945 ;
        RECT 55.790 71.055 56.125 72.025 ;
        RECT 56.295 70.885 56.465 72.025 ;
        RECT 56.635 71.225 56.805 72.195 ;
        RECT 56.975 71.565 57.145 72.695 ;
        RECT 57.315 71.905 57.485 72.705 ;
        RECT 57.690 72.415 57.965 73.265 ;
        RECT 57.685 72.245 57.965 72.415 ;
        RECT 57.690 72.105 57.965 72.245 ;
        RECT 58.135 71.905 58.325 73.265 ;
        RECT 58.505 72.900 59.015 73.435 ;
        RECT 59.235 72.625 59.480 73.230 ;
        RECT 59.925 72.695 60.310 73.265 ;
        RECT 60.480 72.975 60.805 73.435 ;
        RECT 61.325 72.805 61.605 73.265 ;
        RECT 58.525 72.455 59.755 72.625 ;
        RECT 57.315 71.735 58.325 71.905 ;
        RECT 58.495 71.890 59.245 72.080 ;
        RECT 56.975 71.395 58.100 71.565 ;
        RECT 58.495 71.225 58.665 71.890 ;
        RECT 59.415 71.645 59.755 72.455 ;
        RECT 56.635 71.055 58.665 71.225 ;
        RECT 58.835 70.885 59.005 71.645 ;
        RECT 59.240 71.235 59.755 71.645 ;
        RECT 59.925 72.025 60.205 72.695 ;
        RECT 60.480 72.635 61.605 72.805 ;
        RECT 60.480 72.525 60.930 72.635 ;
        RECT 60.375 72.195 60.930 72.525 ;
        RECT 61.795 72.465 62.195 73.265 ;
        RECT 62.595 72.975 62.865 73.435 ;
        RECT 63.035 72.805 63.320 73.265 ;
        RECT 59.925 71.055 60.310 72.025 ;
        RECT 60.480 71.735 60.930 72.195 ;
        RECT 61.100 71.905 62.195 72.465 ;
        RECT 60.480 71.515 61.605 71.735 ;
        RECT 60.480 70.885 60.805 71.345 ;
        RECT 61.325 71.055 61.605 71.515 ;
        RECT 61.795 71.055 62.195 71.905 ;
        RECT 62.365 72.635 63.320 72.805 ;
        RECT 63.605 72.685 64.815 73.435 ;
        RECT 64.985 72.710 65.275 73.435 ;
        RECT 65.925 72.965 66.220 73.435 ;
        RECT 66.390 72.795 66.650 73.240 ;
        RECT 66.820 72.965 67.080 73.435 ;
        RECT 67.250 72.795 67.505 73.240 ;
        RECT 67.675 72.965 67.975 73.435 ;
        RECT 62.365 71.735 62.575 72.635 ;
        RECT 62.745 71.905 63.435 72.465 ;
        RECT 63.605 72.145 64.125 72.685 ;
        RECT 65.465 72.625 68.495 72.795 ;
        RECT 68.665 72.635 69.360 73.265 ;
        RECT 69.565 72.635 69.875 73.435 ;
        RECT 70.045 72.635 70.740 73.265 ;
        RECT 70.945 72.635 71.255 73.435 ;
        RECT 64.295 71.975 64.815 72.515 ;
        RECT 65.465 72.060 65.635 72.625 ;
        RECT 65.805 72.230 68.020 72.455 ;
        RECT 68.195 72.060 68.495 72.625 ;
        RECT 68.685 72.195 69.020 72.445 ;
        RECT 62.365 71.515 63.320 71.735 ;
        RECT 62.595 70.885 62.865 71.345 ;
        RECT 63.035 71.055 63.320 71.515 ;
        RECT 63.605 70.885 64.815 71.975 ;
        RECT 64.985 70.885 65.275 72.050 ;
        RECT 65.465 71.890 68.495 72.060 ;
        RECT 69.190 72.035 69.360 72.635 ;
        RECT 69.530 72.195 69.865 72.465 ;
        RECT 70.065 72.195 70.400 72.445 ;
        RECT 70.570 72.035 70.740 72.635 ;
        RECT 71.435 72.625 71.705 73.435 ;
        RECT 71.875 72.625 72.205 73.265 ;
        RECT 72.375 72.625 72.615 73.435 ;
        RECT 73.730 72.670 74.185 73.435 ;
        RECT 74.460 73.055 75.760 73.265 ;
        RECT 76.015 73.075 76.345 73.435 ;
        RECT 75.590 72.905 75.760 73.055 ;
        RECT 76.515 72.935 76.775 73.265 ;
        RECT 76.545 72.925 76.775 72.935 ;
        RECT 70.910 72.195 71.245 72.465 ;
        RECT 71.425 72.195 71.775 72.445 ;
        RECT 65.445 70.885 65.790 71.720 ;
        RECT 65.965 71.085 66.220 71.890 ;
        RECT 66.390 70.885 66.650 71.720 ;
        RECT 66.825 71.085 67.080 71.890 ;
        RECT 67.250 70.885 67.510 71.720 ;
        RECT 67.680 71.085 67.940 71.890 ;
        RECT 68.110 70.885 68.495 71.720 ;
        RECT 68.665 70.885 68.925 72.025 ;
        RECT 69.095 71.055 69.425 72.035 ;
        RECT 69.595 70.885 69.875 72.025 ;
        RECT 70.045 70.885 70.305 72.025 ;
        RECT 70.475 71.055 70.805 72.035 ;
        RECT 71.945 72.025 72.115 72.625 ;
        RECT 74.660 72.445 74.880 72.845 ;
        RECT 72.285 72.195 72.635 72.445 ;
        RECT 73.725 72.245 74.215 72.445 ;
        RECT 74.405 72.235 74.880 72.445 ;
        RECT 75.125 72.445 75.335 72.845 ;
        RECT 75.590 72.780 76.345 72.905 ;
        RECT 75.590 72.735 76.435 72.780 ;
        RECT 76.165 72.615 76.435 72.735 ;
        RECT 75.125 72.235 75.455 72.445 ;
        RECT 75.625 72.175 76.035 72.480 ;
        RECT 70.975 70.885 71.255 72.025 ;
        RECT 71.435 70.885 71.765 72.025 ;
        RECT 71.945 71.855 72.625 72.025 ;
        RECT 72.295 71.070 72.625 71.855 ;
        RECT 73.730 72.005 74.905 72.065 ;
        RECT 76.265 72.040 76.435 72.615 ;
        RECT 76.235 72.005 76.435 72.040 ;
        RECT 73.730 71.895 76.435 72.005 ;
        RECT 73.730 71.275 73.985 71.895 ;
        RECT 74.575 71.835 76.375 71.895 ;
        RECT 74.575 71.805 74.905 71.835 ;
        RECT 76.605 71.735 76.775 72.925 ;
        RECT 77.150 72.655 77.650 73.265 ;
        RECT 76.945 72.195 77.295 72.445 ;
        RECT 77.480 72.025 77.650 72.655 ;
        RECT 78.280 72.785 78.610 73.265 ;
        RECT 78.780 72.975 79.005 73.435 ;
        RECT 79.175 72.785 79.505 73.265 ;
        RECT 78.280 72.615 79.505 72.785 ;
        RECT 79.695 72.635 79.945 73.435 ;
        RECT 80.115 72.635 80.455 73.265 ;
        RECT 77.820 72.245 78.150 72.445 ;
        RECT 78.320 72.245 78.650 72.445 ;
        RECT 78.820 72.245 79.240 72.445 ;
        RECT 79.415 72.275 80.110 72.445 ;
        RECT 79.415 72.025 79.585 72.275 ;
        RECT 80.280 72.025 80.455 72.635 ;
        RECT 80.625 72.665 82.295 73.435 ;
        RECT 82.930 72.695 83.185 73.265 ;
        RECT 83.355 73.035 83.685 73.435 ;
        RECT 84.110 72.900 84.640 73.265 ;
        RECT 84.110 72.865 84.285 72.900 ;
        RECT 83.355 72.695 84.285 72.865 ;
        RECT 80.625 72.145 81.375 72.665 ;
        RECT 74.235 71.635 74.420 71.725 ;
        RECT 75.010 71.635 75.845 71.645 ;
        RECT 74.235 71.435 75.845 71.635 ;
        RECT 74.235 71.395 74.465 71.435 ;
        RECT 73.730 71.055 74.065 71.275 ;
        RECT 75.070 70.885 75.425 71.265 ;
        RECT 75.595 71.055 75.845 71.435 ;
        RECT 76.095 70.885 76.345 71.665 ;
        RECT 76.515 71.055 76.775 71.735 ;
        RECT 77.150 71.855 79.585 72.025 ;
        RECT 77.150 71.055 77.480 71.855 ;
        RECT 77.650 70.885 77.980 71.685 ;
        RECT 78.280 71.055 78.610 71.855 ;
        RECT 79.255 70.885 79.505 71.685 ;
        RECT 79.775 70.885 79.945 72.025 ;
        RECT 80.115 71.055 80.455 72.025 ;
        RECT 81.545 71.975 82.295 72.495 ;
        RECT 80.625 70.885 82.295 71.975 ;
        RECT 82.930 72.025 83.100 72.695 ;
        RECT 83.355 72.525 83.525 72.695 ;
        RECT 83.270 72.195 83.525 72.525 ;
        RECT 83.750 72.195 83.945 72.525 ;
        RECT 82.930 71.055 83.265 72.025 ;
        RECT 83.435 70.885 83.605 72.025 ;
        RECT 83.775 71.225 83.945 72.195 ;
        RECT 84.115 71.565 84.285 72.695 ;
        RECT 84.455 71.905 84.625 72.705 ;
        RECT 84.830 72.415 85.105 73.265 ;
        RECT 84.825 72.245 85.105 72.415 ;
        RECT 84.830 72.105 85.105 72.245 ;
        RECT 85.275 71.905 85.465 73.265 ;
        RECT 85.645 72.900 86.155 73.435 ;
        RECT 86.375 72.625 86.620 73.230 ;
        RECT 87.065 72.695 87.450 73.265 ;
        RECT 87.620 72.975 87.945 73.435 ;
        RECT 88.465 72.805 88.745 73.265 ;
        RECT 85.665 72.455 86.895 72.625 ;
        RECT 84.455 71.735 85.465 71.905 ;
        RECT 85.635 71.890 86.385 72.080 ;
        RECT 84.115 71.395 85.240 71.565 ;
        RECT 85.635 71.225 85.805 71.890 ;
        RECT 86.555 71.645 86.895 72.455 ;
        RECT 83.775 71.055 85.805 71.225 ;
        RECT 85.975 70.885 86.145 71.645 ;
        RECT 86.380 71.235 86.895 71.645 ;
        RECT 87.065 72.025 87.345 72.695 ;
        RECT 87.620 72.635 88.745 72.805 ;
        RECT 87.620 72.525 88.070 72.635 ;
        RECT 87.515 72.195 88.070 72.525 ;
        RECT 88.935 72.465 89.335 73.265 ;
        RECT 89.735 72.975 90.005 73.435 ;
        RECT 90.175 72.805 90.460 73.265 ;
        RECT 87.065 71.055 87.450 72.025 ;
        RECT 87.620 71.735 88.070 72.195 ;
        RECT 88.240 71.905 89.335 72.465 ;
        RECT 87.620 71.515 88.745 71.735 ;
        RECT 87.620 70.885 87.945 71.345 ;
        RECT 88.465 71.055 88.745 71.515 ;
        RECT 88.935 71.055 89.335 71.905 ;
        RECT 89.505 72.635 90.460 72.805 ;
        RECT 90.745 72.685 91.955 73.435 ;
        RECT 89.505 71.735 89.715 72.635 ;
        RECT 89.885 71.905 90.575 72.465 ;
        RECT 90.745 71.975 91.265 72.515 ;
        RECT 91.435 72.145 91.955 72.685 ;
        RECT 89.505 71.515 90.460 71.735 ;
        RECT 89.735 70.885 90.005 71.345 ;
        RECT 90.175 71.055 90.460 71.515 ;
        RECT 90.745 70.885 91.955 71.975 ;
        RECT 13.380 70.715 92.040 70.885 ;
        RECT 13.465 69.625 14.675 70.715 ;
        RECT 14.935 70.045 15.105 70.545 ;
        RECT 15.275 70.215 15.605 70.715 ;
        RECT 14.935 69.875 15.600 70.045 ;
        RECT 13.465 68.915 13.985 69.455 ;
        RECT 14.155 69.085 14.675 69.625 ;
        RECT 14.850 69.055 15.200 69.705 ;
        RECT 13.465 68.165 14.675 68.915 ;
        RECT 15.370 68.885 15.600 69.875 ;
        RECT 14.935 68.715 15.600 68.885 ;
        RECT 14.935 68.425 15.105 68.715 ;
        RECT 15.275 68.165 15.605 68.545 ;
        RECT 15.775 68.425 15.960 70.545 ;
        RECT 16.200 70.255 16.465 70.715 ;
        RECT 16.635 70.120 16.885 70.545 ;
        RECT 17.095 70.270 18.200 70.440 ;
        RECT 16.580 69.990 16.885 70.120 ;
        RECT 16.130 68.795 16.410 69.745 ;
        RECT 16.580 68.885 16.750 69.990 ;
        RECT 16.920 69.205 17.160 69.800 ;
        RECT 17.330 69.735 17.860 70.100 ;
        RECT 17.330 69.035 17.500 69.735 ;
        RECT 18.030 69.655 18.200 70.270 ;
        RECT 18.370 69.915 18.540 70.715 ;
        RECT 18.710 70.215 18.960 70.545 ;
        RECT 19.185 70.245 20.070 70.415 ;
        RECT 18.030 69.565 18.540 69.655 ;
        RECT 16.580 68.755 16.805 68.885 ;
        RECT 16.975 68.815 17.500 69.035 ;
        RECT 17.670 69.395 18.540 69.565 ;
        RECT 16.215 68.165 16.465 68.625 ;
        RECT 16.635 68.615 16.805 68.755 ;
        RECT 17.670 68.615 17.840 69.395 ;
        RECT 18.370 69.325 18.540 69.395 ;
        RECT 18.050 69.145 18.250 69.175 ;
        RECT 18.710 69.145 18.880 70.215 ;
        RECT 19.050 69.325 19.240 70.045 ;
        RECT 18.050 68.845 18.880 69.145 ;
        RECT 19.410 69.115 19.730 70.075 ;
        RECT 16.635 68.445 16.970 68.615 ;
        RECT 17.165 68.445 17.840 68.615 ;
        RECT 18.160 68.165 18.530 68.665 ;
        RECT 18.710 68.615 18.880 68.845 ;
        RECT 19.265 68.785 19.730 69.115 ;
        RECT 19.900 69.405 20.070 70.245 ;
        RECT 20.250 70.215 20.565 70.715 ;
        RECT 20.795 69.985 21.135 70.545 ;
        RECT 20.240 69.610 21.135 69.985 ;
        RECT 21.305 69.705 21.475 70.715 ;
        RECT 20.945 69.405 21.135 69.610 ;
        RECT 21.645 69.655 21.975 70.500 ;
        RECT 22.145 69.800 22.315 70.715 ;
        RECT 21.645 69.575 22.035 69.655 ;
        RECT 22.665 69.625 26.175 70.715 ;
        RECT 21.820 69.525 22.035 69.575 ;
        RECT 19.900 69.075 20.775 69.405 ;
        RECT 20.945 69.075 21.695 69.405 ;
        RECT 19.900 68.615 20.070 69.075 ;
        RECT 20.945 68.905 21.145 69.075 ;
        RECT 21.865 68.945 22.035 69.525 ;
        RECT 21.810 68.905 22.035 68.945 ;
        RECT 18.710 68.445 19.115 68.615 ;
        RECT 19.285 68.445 20.070 68.615 ;
        RECT 20.345 68.165 20.555 68.695 ;
        RECT 20.815 68.380 21.145 68.905 ;
        RECT 21.655 68.820 22.035 68.905 ;
        RECT 22.665 68.935 24.315 69.455 ;
        RECT 24.485 69.105 26.175 69.625 ;
        RECT 26.345 69.550 26.635 70.715 ;
        RECT 26.895 70.045 27.065 70.545 ;
        RECT 27.235 70.215 27.565 70.715 ;
        RECT 26.895 69.875 27.560 70.045 ;
        RECT 26.810 69.055 27.160 69.705 ;
        RECT 21.315 68.165 21.485 68.775 ;
        RECT 21.655 68.385 21.985 68.820 ;
        RECT 22.155 68.165 22.325 68.680 ;
        RECT 22.665 68.165 26.175 68.935 ;
        RECT 26.345 68.165 26.635 68.890 ;
        RECT 27.330 68.885 27.560 69.875 ;
        RECT 26.895 68.715 27.560 68.885 ;
        RECT 26.895 68.425 27.065 68.715 ;
        RECT 27.235 68.165 27.565 68.545 ;
        RECT 27.735 68.425 27.920 70.545 ;
        RECT 28.160 70.255 28.425 70.715 ;
        RECT 28.595 70.120 28.845 70.545 ;
        RECT 29.055 70.270 30.160 70.440 ;
        RECT 28.540 69.990 28.845 70.120 ;
        RECT 28.090 68.795 28.370 69.745 ;
        RECT 28.540 68.885 28.710 69.990 ;
        RECT 28.880 69.205 29.120 69.800 ;
        RECT 29.290 69.735 29.820 70.100 ;
        RECT 29.290 69.035 29.460 69.735 ;
        RECT 29.990 69.655 30.160 70.270 ;
        RECT 30.330 69.915 30.500 70.715 ;
        RECT 30.670 70.215 30.920 70.545 ;
        RECT 31.145 70.245 32.030 70.415 ;
        RECT 29.990 69.565 30.500 69.655 ;
        RECT 28.540 68.755 28.765 68.885 ;
        RECT 28.935 68.815 29.460 69.035 ;
        RECT 29.630 69.395 30.500 69.565 ;
        RECT 28.175 68.165 28.425 68.625 ;
        RECT 28.595 68.615 28.765 68.755 ;
        RECT 29.630 68.615 29.800 69.395 ;
        RECT 30.330 69.325 30.500 69.395 ;
        RECT 30.010 69.145 30.210 69.175 ;
        RECT 30.670 69.145 30.840 70.215 ;
        RECT 31.010 69.325 31.200 70.045 ;
        RECT 30.010 68.845 30.840 69.145 ;
        RECT 31.370 69.115 31.690 70.075 ;
        RECT 28.595 68.445 28.930 68.615 ;
        RECT 29.125 68.445 29.800 68.615 ;
        RECT 30.120 68.165 30.490 68.665 ;
        RECT 30.670 68.615 30.840 68.845 ;
        RECT 31.225 68.785 31.690 69.115 ;
        RECT 31.860 69.405 32.030 70.245 ;
        RECT 32.210 70.215 32.525 70.715 ;
        RECT 32.755 69.985 33.095 70.545 ;
        RECT 32.200 69.610 33.095 69.985 ;
        RECT 33.265 69.705 33.435 70.715 ;
        RECT 32.905 69.405 33.095 69.610 ;
        RECT 33.605 69.655 33.935 70.500 ;
        RECT 34.105 69.800 34.275 70.715 ;
        RECT 33.605 69.575 33.995 69.655 ;
        RECT 34.625 69.625 36.295 70.715 ;
        RECT 33.780 69.525 33.995 69.575 ;
        RECT 31.860 69.075 32.735 69.405 ;
        RECT 32.905 69.075 33.655 69.405 ;
        RECT 31.860 68.615 32.030 69.075 ;
        RECT 32.905 68.905 33.105 69.075 ;
        RECT 33.825 68.945 33.995 69.525 ;
        RECT 33.770 68.905 33.995 68.945 ;
        RECT 30.670 68.445 31.075 68.615 ;
        RECT 31.245 68.445 32.030 68.615 ;
        RECT 32.305 68.165 32.515 68.695 ;
        RECT 32.775 68.380 33.105 68.905 ;
        RECT 33.615 68.820 33.995 68.905 ;
        RECT 34.625 68.935 35.375 69.455 ;
        RECT 35.545 69.105 36.295 69.625 ;
        RECT 36.470 69.575 36.805 70.545 ;
        RECT 36.975 69.575 37.145 70.715 ;
        RECT 37.315 70.375 39.345 70.545 ;
        RECT 33.275 68.165 33.445 68.775 ;
        RECT 33.615 68.385 33.945 68.820 ;
        RECT 34.115 68.165 34.285 68.680 ;
        RECT 34.625 68.165 36.295 68.935 ;
        RECT 36.470 68.905 36.640 69.575 ;
        RECT 37.315 69.405 37.485 70.375 ;
        RECT 36.810 69.075 37.065 69.405 ;
        RECT 37.290 69.075 37.485 69.405 ;
        RECT 37.655 70.035 38.780 70.205 ;
        RECT 36.895 68.905 37.065 69.075 ;
        RECT 37.655 68.905 37.825 70.035 ;
        RECT 36.470 68.335 36.725 68.905 ;
        RECT 36.895 68.735 37.825 68.905 ;
        RECT 37.995 69.695 39.005 69.865 ;
        RECT 37.995 68.895 38.165 69.695 ;
        RECT 37.650 68.700 37.825 68.735 ;
        RECT 36.895 68.165 37.225 68.565 ;
        RECT 37.650 68.335 38.180 68.700 ;
        RECT 38.370 68.675 38.645 69.495 ;
        RECT 38.365 68.505 38.645 68.675 ;
        RECT 38.370 68.335 38.645 68.505 ;
        RECT 38.815 68.335 39.005 69.695 ;
        RECT 39.175 69.710 39.345 70.375 ;
        RECT 39.515 69.955 39.685 70.715 ;
        RECT 39.920 69.955 40.435 70.365 ;
        RECT 39.175 69.520 39.925 69.710 ;
        RECT 40.095 69.145 40.435 69.955 ;
        RECT 40.695 70.045 40.865 70.545 ;
        RECT 41.035 70.215 41.365 70.715 ;
        RECT 40.695 69.875 41.360 70.045 ;
        RECT 39.205 68.975 40.435 69.145 ;
        RECT 40.610 69.055 40.960 69.705 ;
        RECT 39.185 68.165 39.695 68.700 ;
        RECT 39.915 68.370 40.160 68.975 ;
        RECT 41.130 68.885 41.360 69.875 ;
        RECT 40.695 68.715 41.360 68.885 ;
        RECT 40.695 68.425 40.865 68.715 ;
        RECT 41.035 68.165 41.365 68.545 ;
        RECT 41.535 68.425 41.720 70.545 ;
        RECT 41.960 70.255 42.225 70.715 ;
        RECT 42.395 70.120 42.645 70.545 ;
        RECT 42.855 70.270 43.960 70.440 ;
        RECT 42.340 69.990 42.645 70.120 ;
        RECT 41.890 68.795 42.170 69.745 ;
        RECT 42.340 68.885 42.510 69.990 ;
        RECT 42.680 69.205 42.920 69.800 ;
        RECT 43.090 69.735 43.620 70.100 ;
        RECT 43.090 69.035 43.260 69.735 ;
        RECT 43.790 69.655 43.960 70.270 ;
        RECT 44.130 69.915 44.300 70.715 ;
        RECT 44.470 70.215 44.720 70.545 ;
        RECT 44.945 70.245 45.830 70.415 ;
        RECT 43.790 69.565 44.300 69.655 ;
        RECT 42.340 68.755 42.565 68.885 ;
        RECT 42.735 68.815 43.260 69.035 ;
        RECT 43.430 69.395 44.300 69.565 ;
        RECT 41.975 68.165 42.225 68.625 ;
        RECT 42.395 68.615 42.565 68.755 ;
        RECT 43.430 68.615 43.600 69.395 ;
        RECT 44.130 69.325 44.300 69.395 ;
        RECT 43.810 69.145 44.010 69.175 ;
        RECT 44.470 69.145 44.640 70.215 ;
        RECT 44.810 69.325 45.000 70.045 ;
        RECT 43.810 68.845 44.640 69.145 ;
        RECT 45.170 69.115 45.490 70.075 ;
        RECT 42.395 68.445 42.730 68.615 ;
        RECT 42.925 68.445 43.600 68.615 ;
        RECT 43.920 68.165 44.290 68.665 ;
        RECT 44.470 68.615 44.640 68.845 ;
        RECT 45.025 68.785 45.490 69.115 ;
        RECT 45.660 69.405 45.830 70.245 ;
        RECT 46.010 70.215 46.325 70.715 ;
        RECT 46.555 69.985 46.895 70.545 ;
        RECT 46.000 69.610 46.895 69.985 ;
        RECT 47.065 69.705 47.235 70.715 ;
        RECT 46.705 69.405 46.895 69.610 ;
        RECT 47.405 69.655 47.735 70.500 ;
        RECT 47.405 69.575 47.795 69.655 ;
        RECT 47.580 69.525 47.795 69.575 ;
        RECT 45.660 69.075 46.535 69.405 ;
        RECT 46.705 69.075 47.455 69.405 ;
        RECT 45.660 68.615 45.830 69.075 ;
        RECT 46.705 68.905 46.905 69.075 ;
        RECT 47.625 68.945 47.795 69.525 ;
        RECT 47.570 68.905 47.795 68.945 ;
        RECT 44.470 68.445 44.875 68.615 ;
        RECT 45.045 68.445 45.830 68.615 ;
        RECT 46.105 68.165 46.315 68.695 ;
        RECT 46.575 68.380 46.905 68.905 ;
        RECT 47.415 68.820 47.795 68.905 ;
        RECT 47.970 69.575 48.305 70.545 ;
        RECT 48.475 69.575 48.645 70.715 ;
        RECT 48.815 70.375 50.845 70.545 ;
        RECT 47.970 68.905 48.140 69.575 ;
        RECT 48.815 69.405 48.985 70.375 ;
        RECT 48.310 69.075 48.565 69.405 ;
        RECT 48.790 69.075 48.985 69.405 ;
        RECT 49.155 70.035 50.280 70.205 ;
        RECT 48.395 68.905 48.565 69.075 ;
        RECT 49.155 68.905 49.325 70.035 ;
        RECT 47.075 68.165 47.245 68.775 ;
        RECT 47.415 68.385 47.745 68.820 ;
        RECT 47.970 68.335 48.225 68.905 ;
        RECT 48.395 68.735 49.325 68.905 ;
        RECT 49.495 69.695 50.505 69.865 ;
        RECT 49.495 68.895 49.665 69.695 ;
        RECT 49.150 68.700 49.325 68.735 ;
        RECT 48.395 68.165 48.725 68.565 ;
        RECT 49.150 68.335 49.680 68.700 ;
        RECT 49.870 68.675 50.145 69.495 ;
        RECT 49.865 68.505 50.145 68.675 ;
        RECT 49.870 68.335 50.145 68.505 ;
        RECT 50.315 68.335 50.505 69.695 ;
        RECT 50.675 69.710 50.845 70.375 ;
        RECT 51.015 69.955 51.185 70.715 ;
        RECT 51.420 69.955 51.935 70.365 ;
        RECT 50.675 69.520 51.425 69.710 ;
        RECT 51.595 69.145 51.935 69.955 ;
        RECT 52.105 69.550 52.395 70.715 ;
        RECT 52.565 69.575 52.950 70.545 ;
        RECT 53.120 70.255 53.445 70.715 ;
        RECT 53.965 70.085 54.245 70.545 ;
        RECT 53.120 69.865 54.245 70.085 ;
        RECT 50.705 68.975 51.935 69.145 ;
        RECT 50.685 68.165 51.195 68.700 ;
        RECT 51.415 68.370 51.660 68.975 ;
        RECT 52.565 68.905 52.845 69.575 ;
        RECT 53.120 69.405 53.570 69.865 ;
        RECT 54.435 69.695 54.835 70.545 ;
        RECT 55.235 70.255 55.505 70.715 ;
        RECT 55.675 70.085 55.960 70.545 ;
        RECT 53.015 69.075 53.570 69.405 ;
        RECT 53.740 69.135 54.835 69.695 ;
        RECT 53.120 68.965 53.570 69.075 ;
        RECT 52.105 68.165 52.395 68.890 ;
        RECT 52.565 68.335 52.950 68.905 ;
        RECT 53.120 68.795 54.245 68.965 ;
        RECT 53.120 68.165 53.445 68.625 ;
        RECT 53.965 68.335 54.245 68.795 ;
        RECT 54.435 68.335 54.835 69.135 ;
        RECT 55.005 69.865 55.960 70.085 ;
        RECT 55.005 68.965 55.215 69.865 ;
        RECT 55.385 69.135 56.075 69.695 ;
        RECT 56.245 69.625 59.755 70.715 ;
        RECT 55.005 68.795 55.960 68.965 ;
        RECT 55.235 68.165 55.505 68.625 ;
        RECT 55.675 68.335 55.960 68.795 ;
        RECT 56.245 68.935 57.895 69.455 ;
        RECT 58.065 69.105 59.755 69.625 ;
        RECT 60.855 69.605 61.150 70.715 ;
        RECT 61.330 69.405 61.580 70.540 ;
        RECT 61.750 69.605 62.010 70.715 ;
        RECT 62.180 69.815 62.440 70.540 ;
        RECT 62.610 69.985 62.870 70.715 ;
        RECT 63.040 69.815 63.300 70.540 ;
        RECT 63.470 69.985 63.730 70.715 ;
        RECT 63.900 69.815 64.160 70.540 ;
        RECT 64.330 69.985 64.590 70.715 ;
        RECT 64.760 69.815 65.020 70.540 ;
        RECT 65.190 69.985 65.485 70.715 ;
        RECT 66.020 70.085 66.305 70.545 ;
        RECT 66.475 70.255 66.745 70.715 ;
        RECT 66.020 69.865 66.975 70.085 ;
        RECT 62.180 69.575 65.490 69.815 ;
        RECT 56.245 68.165 59.755 68.935 ;
        RECT 60.845 68.795 61.160 69.405 ;
        RECT 61.330 69.155 64.350 69.405 ;
        RECT 60.905 68.165 61.150 68.625 ;
        RECT 61.330 68.345 61.580 69.155 ;
        RECT 64.520 68.985 65.490 69.575 ;
        RECT 65.905 69.135 66.595 69.695 ;
        RECT 62.180 68.815 65.490 68.985 ;
        RECT 66.765 68.965 66.975 69.865 ;
        RECT 61.750 68.165 62.010 68.690 ;
        RECT 62.180 68.360 62.440 68.815 ;
        RECT 62.610 68.165 62.870 68.645 ;
        RECT 63.040 68.360 63.300 68.815 ;
        RECT 63.470 68.165 63.730 68.645 ;
        RECT 63.900 68.360 64.160 68.815 ;
        RECT 64.330 68.165 64.590 68.645 ;
        RECT 64.760 68.360 65.020 68.815 ;
        RECT 66.020 68.795 66.975 68.965 ;
        RECT 67.145 69.695 67.545 70.545 ;
        RECT 67.735 70.085 68.015 70.545 ;
        RECT 68.535 70.255 68.860 70.715 ;
        RECT 67.735 69.865 68.860 70.085 ;
        RECT 67.145 69.135 68.240 69.695 ;
        RECT 68.410 69.405 68.860 69.865 ;
        RECT 69.030 69.575 69.415 70.545 ;
        RECT 65.190 68.165 65.490 68.645 ;
        RECT 66.020 68.335 66.305 68.795 ;
        RECT 66.475 68.165 66.745 68.625 ;
        RECT 67.145 68.335 67.545 69.135 ;
        RECT 68.410 69.075 68.965 69.405 ;
        RECT 68.410 68.965 68.860 69.075 ;
        RECT 67.735 68.795 68.860 68.965 ;
        RECT 69.135 68.905 69.415 69.575 ;
        RECT 67.735 68.335 68.015 68.795 ;
        RECT 68.535 68.165 68.860 68.625 ;
        RECT 69.030 68.335 69.415 68.905 ;
        RECT 69.585 69.995 70.045 70.545 ;
        RECT 70.235 69.995 70.565 70.715 ;
        RECT 69.585 68.625 69.835 69.995 ;
        RECT 70.765 69.825 71.065 70.375 ;
        RECT 71.235 70.045 71.515 70.715 ;
        RECT 70.125 69.655 71.065 69.825 ;
        RECT 70.125 69.405 70.295 69.655 ;
        RECT 71.435 69.405 71.700 69.765 ;
        RECT 71.945 69.575 72.155 70.715 ;
        RECT 70.005 69.075 70.295 69.405 ;
        RECT 70.465 69.155 70.805 69.405 ;
        RECT 71.025 69.155 71.700 69.405 ;
        RECT 72.325 69.565 72.655 70.545 ;
        RECT 72.825 69.575 73.055 70.715 ;
        RECT 73.265 69.575 73.545 70.715 ;
        RECT 73.715 69.565 74.045 70.545 ;
        RECT 74.215 69.575 74.475 70.715 ;
        RECT 74.645 70.205 75.835 70.495 ;
        RECT 74.665 69.865 75.835 70.035 ;
        RECT 76.005 69.915 76.285 70.715 ;
        RECT 74.665 69.575 74.990 69.865 ;
        RECT 75.665 69.745 75.835 69.865 ;
        RECT 70.125 68.985 70.295 69.075 ;
        RECT 70.125 68.795 71.515 68.985 ;
        RECT 69.585 68.335 70.145 68.625 ;
        RECT 70.315 68.165 70.565 68.625 ;
        RECT 71.185 68.435 71.515 68.795 ;
        RECT 71.945 68.165 72.155 68.985 ;
        RECT 72.325 68.965 72.575 69.565 ;
        RECT 72.745 69.155 73.075 69.405 ;
        RECT 73.275 69.135 73.610 69.405 ;
        RECT 72.325 68.335 72.655 68.965 ;
        RECT 72.825 68.165 73.055 68.985 ;
        RECT 73.780 68.965 73.950 69.565 ;
        RECT 75.160 69.405 75.355 69.695 ;
        RECT 75.665 69.575 76.325 69.745 ;
        RECT 76.495 69.575 76.770 70.545 ;
        RECT 76.155 69.405 76.325 69.575 ;
        RECT 74.120 69.155 74.455 69.405 ;
        RECT 74.645 69.075 74.990 69.405 ;
        RECT 75.160 69.075 75.985 69.405 ;
        RECT 76.155 69.075 76.430 69.405 ;
        RECT 73.265 68.165 73.575 68.965 ;
        RECT 73.780 68.335 74.475 68.965 ;
        RECT 76.155 68.905 76.325 69.075 ;
        RECT 74.660 68.735 76.325 68.905 ;
        RECT 76.600 68.840 76.770 69.575 ;
        RECT 77.865 69.550 78.155 70.715 ;
        RECT 79.250 70.325 79.585 70.545 ;
        RECT 80.590 70.335 80.945 70.715 ;
        RECT 79.250 69.705 79.505 70.325 ;
        RECT 79.755 70.165 79.985 70.205 ;
        RECT 81.115 70.165 81.365 70.545 ;
        RECT 79.755 69.965 81.365 70.165 ;
        RECT 79.755 69.875 79.940 69.965 ;
        RECT 80.530 69.955 81.365 69.965 ;
        RECT 81.615 69.935 81.865 70.715 ;
        RECT 82.035 69.865 82.295 70.545 ;
        RECT 80.095 69.765 80.425 69.795 ;
        RECT 80.095 69.705 81.895 69.765 ;
        RECT 79.250 69.595 81.955 69.705 ;
        RECT 79.250 69.535 80.425 69.595 ;
        RECT 81.755 69.560 81.955 69.595 ;
        RECT 79.245 69.155 79.735 69.355 ;
        RECT 79.925 69.155 80.400 69.365 ;
        RECT 74.660 68.385 74.915 68.735 ;
        RECT 75.085 68.165 75.415 68.565 ;
        RECT 75.585 68.385 75.755 68.735 ;
        RECT 75.925 68.165 76.305 68.565 ;
        RECT 76.495 68.495 76.770 68.840 ;
        RECT 77.865 68.165 78.155 68.890 ;
        RECT 79.250 68.165 79.705 68.930 ;
        RECT 80.180 68.755 80.400 69.155 ;
        RECT 80.645 69.155 80.975 69.365 ;
        RECT 80.645 68.755 80.855 69.155 ;
        RECT 81.145 69.120 81.555 69.425 ;
        RECT 81.785 68.985 81.955 69.560 ;
        RECT 81.685 68.865 81.955 68.985 ;
        RECT 81.110 68.820 81.955 68.865 ;
        RECT 81.110 68.695 81.865 68.820 ;
        RECT 81.110 68.545 81.280 68.695 ;
        RECT 82.125 68.675 82.295 69.865 ;
        RECT 82.465 69.625 85.055 70.715 ;
        RECT 82.065 68.665 82.295 68.675 ;
        RECT 79.980 68.335 81.280 68.545 ;
        RECT 81.535 68.165 81.865 68.525 ;
        RECT 82.035 68.335 82.295 68.665 ;
        RECT 82.465 68.935 83.675 69.455 ;
        RECT 83.845 69.105 85.055 69.625 ;
        RECT 85.230 69.565 85.490 70.715 ;
        RECT 85.665 69.640 85.920 70.545 ;
        RECT 86.090 69.955 86.420 70.715 ;
        RECT 86.635 69.785 86.805 70.545 ;
        RECT 82.465 68.165 85.055 68.935 ;
        RECT 85.230 68.165 85.490 69.005 ;
        RECT 85.665 68.910 85.835 69.640 ;
        RECT 86.090 69.615 86.805 69.785 ;
        RECT 86.090 69.405 86.260 69.615 ;
        RECT 87.065 69.575 87.450 70.545 ;
        RECT 87.620 70.255 87.945 70.715 ;
        RECT 88.465 70.085 88.745 70.545 ;
        RECT 87.620 69.865 88.745 70.085 ;
        RECT 86.005 69.075 86.260 69.405 ;
        RECT 85.665 68.335 85.920 68.910 ;
        RECT 86.090 68.885 86.260 69.075 ;
        RECT 86.540 69.065 86.895 69.435 ;
        RECT 87.065 68.905 87.345 69.575 ;
        RECT 87.620 69.405 88.070 69.865 ;
        RECT 88.935 69.695 89.335 70.545 ;
        RECT 89.735 70.255 90.005 70.715 ;
        RECT 90.175 70.085 90.460 70.545 ;
        RECT 87.515 69.075 88.070 69.405 ;
        RECT 88.240 69.135 89.335 69.695 ;
        RECT 87.620 68.965 88.070 69.075 ;
        RECT 86.090 68.715 86.805 68.885 ;
        RECT 86.090 68.165 86.420 68.545 ;
        RECT 86.635 68.335 86.805 68.715 ;
        RECT 87.065 68.335 87.450 68.905 ;
        RECT 87.620 68.795 88.745 68.965 ;
        RECT 87.620 68.165 87.945 68.625 ;
        RECT 88.465 68.335 88.745 68.795 ;
        RECT 88.935 68.335 89.335 69.135 ;
        RECT 89.505 69.865 90.460 70.085 ;
        RECT 89.505 68.965 89.715 69.865 ;
        RECT 89.885 69.135 90.575 69.695 ;
        RECT 90.745 69.625 91.955 70.715 ;
        RECT 90.745 69.085 91.265 69.625 ;
        RECT 89.505 68.795 90.460 68.965 ;
        RECT 91.435 68.915 91.955 69.455 ;
        RECT 89.735 68.165 90.005 68.625 ;
        RECT 90.175 68.335 90.460 68.795 ;
        RECT 90.745 68.165 91.955 68.915 ;
        RECT 13.380 67.995 92.040 68.165 ;
        RECT 13.465 67.245 14.675 67.995 ;
        RECT 13.465 66.705 13.985 67.245 ;
        RECT 14.850 67.155 15.110 67.995 ;
        RECT 15.285 67.250 15.540 67.825 ;
        RECT 15.710 67.615 16.040 67.995 ;
        RECT 16.255 67.445 16.425 67.825 ;
        RECT 15.710 67.275 16.425 67.445 ;
        RECT 17.695 67.445 17.865 67.735 ;
        RECT 18.035 67.615 18.365 67.995 ;
        RECT 17.695 67.275 18.360 67.445 ;
        RECT 14.155 66.535 14.675 67.075 ;
        RECT 13.465 65.445 14.675 66.535 ;
        RECT 14.850 65.445 15.110 66.595 ;
        RECT 15.285 66.520 15.455 67.250 ;
        RECT 15.710 67.085 15.880 67.275 ;
        RECT 15.625 66.755 15.880 67.085 ;
        RECT 15.710 66.545 15.880 66.755 ;
        RECT 16.160 66.725 16.515 67.095 ;
        RECT 15.285 65.615 15.540 66.520 ;
        RECT 15.710 66.375 16.425 66.545 ;
        RECT 17.610 66.455 17.960 67.105 ;
        RECT 15.710 65.445 16.040 66.205 ;
        RECT 16.255 65.615 16.425 66.375 ;
        RECT 18.130 66.285 18.360 67.275 ;
        RECT 17.695 66.115 18.360 66.285 ;
        RECT 17.695 65.615 17.865 66.115 ;
        RECT 18.035 65.445 18.365 65.945 ;
        RECT 18.535 65.615 18.720 67.735 ;
        RECT 18.975 67.535 19.225 67.995 ;
        RECT 19.395 67.545 19.730 67.715 ;
        RECT 19.925 67.545 20.600 67.715 ;
        RECT 19.395 67.405 19.565 67.545 ;
        RECT 18.890 66.415 19.170 67.365 ;
        RECT 19.340 67.275 19.565 67.405 ;
        RECT 19.340 66.170 19.510 67.275 ;
        RECT 19.735 67.125 20.260 67.345 ;
        RECT 19.680 66.360 19.920 66.955 ;
        RECT 20.090 66.425 20.260 67.125 ;
        RECT 20.430 66.765 20.600 67.545 ;
        RECT 20.920 67.495 21.290 67.995 ;
        RECT 21.470 67.545 21.875 67.715 ;
        RECT 22.045 67.545 22.830 67.715 ;
        RECT 21.470 67.315 21.640 67.545 ;
        RECT 20.810 67.015 21.640 67.315 ;
        RECT 22.025 67.045 22.490 67.375 ;
        RECT 20.810 66.985 21.010 67.015 ;
        RECT 21.130 66.765 21.300 66.835 ;
        RECT 20.430 66.595 21.300 66.765 ;
        RECT 20.790 66.505 21.300 66.595 ;
        RECT 19.340 66.040 19.645 66.170 ;
        RECT 20.090 66.060 20.620 66.425 ;
        RECT 18.960 65.445 19.225 65.905 ;
        RECT 19.395 65.615 19.645 66.040 ;
        RECT 20.790 65.890 20.960 66.505 ;
        RECT 19.855 65.720 20.960 65.890 ;
        RECT 21.130 65.445 21.300 66.245 ;
        RECT 21.470 65.945 21.640 67.015 ;
        RECT 21.810 66.115 22.000 66.835 ;
        RECT 22.170 66.085 22.490 67.045 ;
        RECT 22.660 67.085 22.830 67.545 ;
        RECT 23.105 67.465 23.315 67.995 ;
        RECT 23.575 67.255 23.905 67.780 ;
        RECT 24.075 67.385 24.245 67.995 ;
        RECT 24.415 67.340 24.745 67.775 ;
        RECT 24.915 67.480 25.085 67.995 ;
        RECT 24.415 67.255 24.795 67.340 ;
        RECT 23.705 67.085 23.905 67.255 ;
        RECT 24.570 67.215 24.795 67.255 ;
        RECT 22.660 66.755 23.535 67.085 ;
        RECT 23.705 66.755 24.455 67.085 ;
        RECT 21.470 65.615 21.720 65.945 ;
        RECT 22.660 65.915 22.830 66.755 ;
        RECT 23.705 66.550 23.895 66.755 ;
        RECT 24.625 66.635 24.795 67.215 ;
        RECT 25.700 67.185 25.945 67.790 ;
        RECT 26.165 67.460 26.675 67.995 ;
        RECT 24.580 66.585 24.795 66.635 ;
        RECT 23.000 66.175 23.895 66.550 ;
        RECT 24.405 66.505 24.795 66.585 ;
        RECT 25.425 67.015 26.655 67.185 ;
        RECT 21.945 65.745 22.830 65.915 ;
        RECT 23.010 65.445 23.325 65.945 ;
        RECT 23.555 65.615 23.895 66.175 ;
        RECT 24.065 65.445 24.235 66.455 ;
        RECT 24.405 65.660 24.735 66.505 ;
        RECT 24.905 65.445 25.075 66.360 ;
        RECT 25.425 66.205 25.765 67.015 ;
        RECT 25.935 66.450 26.685 66.640 ;
        RECT 25.425 65.795 25.940 66.205 ;
        RECT 26.175 65.445 26.345 66.205 ;
        RECT 26.515 65.785 26.685 66.450 ;
        RECT 26.855 66.465 27.045 67.825 ;
        RECT 27.215 67.655 27.490 67.825 ;
        RECT 27.215 67.485 27.495 67.655 ;
        RECT 27.215 66.665 27.490 67.485 ;
        RECT 27.680 67.460 28.210 67.825 ;
        RECT 28.635 67.595 28.965 67.995 ;
        RECT 28.035 67.425 28.210 67.460 ;
        RECT 27.695 66.465 27.865 67.265 ;
        RECT 26.855 66.295 27.865 66.465 ;
        RECT 28.035 67.255 28.965 67.425 ;
        RECT 29.135 67.255 29.390 67.825 ;
        RECT 29.565 67.450 34.910 67.995 ;
        RECT 28.035 66.125 28.205 67.255 ;
        RECT 28.795 67.085 28.965 67.255 ;
        RECT 27.080 65.955 28.205 66.125 ;
        RECT 28.375 66.755 28.570 67.085 ;
        RECT 28.795 66.755 29.050 67.085 ;
        RECT 28.375 65.785 28.545 66.755 ;
        RECT 29.220 66.585 29.390 67.255 ;
        RECT 31.150 66.620 31.490 67.450 ;
        RECT 35.085 67.225 38.595 67.995 ;
        RECT 39.225 67.270 39.515 67.995 ;
        RECT 40.145 67.255 40.530 67.825 ;
        RECT 40.700 67.535 41.025 67.995 ;
        RECT 41.545 67.365 41.825 67.825 ;
        RECT 26.515 65.615 28.545 65.785 ;
        RECT 28.715 65.445 28.885 66.585 ;
        RECT 29.055 65.615 29.390 66.585 ;
        RECT 32.970 65.880 33.320 67.130 ;
        RECT 35.085 66.705 36.735 67.225 ;
        RECT 36.905 66.535 38.595 67.055 ;
        RECT 29.565 65.445 34.910 65.880 ;
        RECT 35.085 65.445 38.595 66.535 ;
        RECT 39.225 65.445 39.515 66.610 ;
        RECT 40.145 66.585 40.425 67.255 ;
        RECT 40.700 67.195 41.825 67.365 ;
        RECT 40.700 67.085 41.150 67.195 ;
        RECT 40.595 66.755 41.150 67.085 ;
        RECT 42.015 67.025 42.415 67.825 ;
        RECT 42.815 67.535 43.085 67.995 ;
        RECT 43.255 67.365 43.540 67.825 ;
        RECT 40.145 65.615 40.530 66.585 ;
        RECT 40.700 66.295 41.150 66.755 ;
        RECT 41.320 66.465 42.415 67.025 ;
        RECT 40.700 66.075 41.825 66.295 ;
        RECT 40.700 65.445 41.025 65.905 ;
        RECT 41.545 65.615 41.825 66.075 ;
        RECT 42.015 65.615 42.415 66.465 ;
        RECT 42.585 67.195 43.540 67.365 ;
        RECT 43.875 67.455 44.100 67.815 ;
        RECT 44.280 67.625 44.610 67.995 ;
        RECT 44.790 67.455 45.045 67.815 ;
        RECT 45.610 67.625 46.355 67.995 ;
        RECT 43.875 67.265 46.360 67.455 ;
        RECT 42.585 66.295 42.795 67.195 ;
        RECT 42.965 66.465 43.655 67.025 ;
        RECT 43.835 66.755 44.105 67.085 ;
        RECT 44.285 66.755 44.720 67.085 ;
        RECT 44.900 66.755 45.475 67.085 ;
        RECT 45.655 66.755 45.935 67.085 ;
        RECT 46.135 66.575 46.360 67.265 ;
        RECT 43.865 66.395 46.360 66.575 ;
        RECT 46.535 66.395 46.870 67.815 ;
        RECT 47.045 67.245 48.255 67.995 ;
        RECT 48.425 67.255 48.810 67.825 ;
        RECT 48.980 67.535 49.305 67.995 ;
        RECT 49.825 67.365 50.105 67.825 ;
        RECT 47.045 66.705 47.565 67.245 ;
        RECT 47.735 66.535 48.255 67.075 ;
        RECT 42.585 66.075 43.540 66.295 ;
        RECT 42.815 65.445 43.085 65.905 ;
        RECT 43.255 65.615 43.540 66.075 ;
        RECT 43.865 65.625 44.155 66.395 ;
        RECT 44.725 65.985 45.915 66.215 ;
        RECT 44.725 65.625 44.985 65.985 ;
        RECT 45.155 65.445 45.485 65.815 ;
        RECT 45.655 65.625 45.915 65.985 ;
        RECT 46.105 65.445 46.435 66.165 ;
        RECT 46.605 65.625 46.870 66.395 ;
        RECT 47.045 65.445 48.255 66.535 ;
        RECT 48.425 66.585 48.705 67.255 ;
        RECT 48.980 67.195 50.105 67.365 ;
        RECT 48.980 67.085 49.430 67.195 ;
        RECT 48.875 66.755 49.430 67.085 ;
        RECT 50.295 67.025 50.695 67.825 ;
        RECT 51.095 67.535 51.365 67.995 ;
        RECT 51.535 67.365 51.820 67.825 ;
        RECT 48.425 65.615 48.810 66.585 ;
        RECT 48.980 66.295 49.430 66.755 ;
        RECT 49.600 66.465 50.695 67.025 ;
        RECT 48.980 66.075 50.105 66.295 ;
        RECT 48.980 65.445 49.305 65.905 ;
        RECT 49.825 65.615 50.105 66.075 ;
        RECT 50.295 65.615 50.695 66.465 ;
        RECT 50.865 67.195 51.820 67.365 ;
        RECT 53.030 67.255 53.285 67.825 ;
        RECT 53.455 67.595 53.785 67.995 ;
        RECT 54.210 67.460 54.740 67.825 ;
        RECT 54.210 67.425 54.385 67.460 ;
        RECT 53.455 67.255 54.385 67.425 ;
        RECT 50.865 66.295 51.075 67.195 ;
        RECT 51.245 66.465 51.935 67.025 ;
        RECT 53.030 66.585 53.200 67.255 ;
        RECT 53.455 67.085 53.625 67.255 ;
        RECT 53.370 66.755 53.625 67.085 ;
        RECT 53.850 66.755 54.045 67.085 ;
        RECT 50.865 66.075 51.820 66.295 ;
        RECT 51.095 65.445 51.365 65.905 ;
        RECT 51.535 65.615 51.820 66.075 ;
        RECT 53.030 65.615 53.365 66.585 ;
        RECT 53.535 65.445 53.705 66.585 ;
        RECT 53.875 65.785 54.045 66.755 ;
        RECT 54.215 66.125 54.385 67.255 ;
        RECT 54.555 66.465 54.725 67.265 ;
        RECT 54.930 66.975 55.205 67.825 ;
        RECT 54.925 66.805 55.205 66.975 ;
        RECT 54.930 66.665 55.205 66.805 ;
        RECT 55.375 66.465 55.565 67.825 ;
        RECT 55.745 67.460 56.255 67.995 ;
        RECT 56.475 67.185 56.720 67.790 ;
        RECT 57.215 67.340 57.545 67.775 ;
        RECT 57.715 67.385 57.885 67.995 ;
        RECT 57.165 67.255 57.545 67.340 ;
        RECT 58.055 67.255 58.385 67.780 ;
        RECT 58.645 67.465 58.855 67.995 ;
        RECT 59.130 67.545 59.915 67.715 ;
        RECT 60.085 67.545 60.490 67.715 ;
        RECT 57.165 67.215 57.390 67.255 ;
        RECT 55.765 67.015 56.995 67.185 ;
        RECT 54.555 66.295 55.565 66.465 ;
        RECT 55.735 66.450 56.485 66.640 ;
        RECT 54.215 65.955 55.340 66.125 ;
        RECT 55.735 65.785 55.905 66.450 ;
        RECT 56.655 66.205 56.995 67.015 ;
        RECT 57.165 66.635 57.335 67.215 ;
        RECT 58.055 67.085 58.255 67.255 ;
        RECT 59.130 67.085 59.300 67.545 ;
        RECT 57.505 66.755 58.255 67.085 ;
        RECT 58.425 66.755 59.300 67.085 ;
        RECT 57.165 66.585 57.380 66.635 ;
        RECT 57.165 66.505 57.555 66.585 ;
        RECT 53.875 65.615 55.905 65.785 ;
        RECT 56.075 65.445 56.245 66.205 ;
        RECT 56.480 65.795 56.995 66.205 ;
        RECT 57.225 65.660 57.555 66.505 ;
        RECT 58.065 66.550 58.255 66.755 ;
        RECT 57.725 65.445 57.895 66.455 ;
        RECT 58.065 66.175 58.960 66.550 ;
        RECT 58.065 65.615 58.405 66.175 ;
        RECT 58.635 65.445 58.950 65.945 ;
        RECT 59.130 65.915 59.300 66.755 ;
        RECT 59.470 67.045 59.935 67.375 ;
        RECT 60.320 67.315 60.490 67.545 ;
        RECT 60.670 67.495 61.040 67.995 ;
        RECT 61.360 67.545 62.035 67.715 ;
        RECT 62.230 67.545 62.565 67.715 ;
        RECT 59.470 66.085 59.790 67.045 ;
        RECT 60.320 67.015 61.150 67.315 ;
        RECT 59.960 66.115 60.150 66.835 ;
        RECT 60.320 65.945 60.490 67.015 ;
        RECT 60.950 66.985 61.150 67.015 ;
        RECT 60.660 66.765 60.830 66.835 ;
        RECT 61.360 66.765 61.530 67.545 ;
        RECT 62.395 67.405 62.565 67.545 ;
        RECT 62.735 67.535 62.985 67.995 ;
        RECT 60.660 66.595 61.530 66.765 ;
        RECT 61.700 67.125 62.225 67.345 ;
        RECT 62.395 67.275 62.620 67.405 ;
        RECT 60.660 66.505 61.170 66.595 ;
        RECT 59.130 65.745 60.015 65.915 ;
        RECT 60.240 65.615 60.490 65.945 ;
        RECT 60.660 65.445 60.830 66.245 ;
        RECT 61.000 65.890 61.170 66.505 ;
        RECT 61.700 66.425 61.870 67.125 ;
        RECT 61.340 66.060 61.870 66.425 ;
        RECT 62.040 66.360 62.280 66.955 ;
        RECT 62.450 66.170 62.620 67.275 ;
        RECT 62.790 66.415 63.070 67.365 ;
        RECT 62.315 66.040 62.620 66.170 ;
        RECT 61.000 65.720 62.105 65.890 ;
        RECT 62.315 65.615 62.565 66.040 ;
        RECT 62.735 65.445 63.000 65.905 ;
        RECT 63.240 65.615 63.425 67.735 ;
        RECT 63.595 67.615 63.925 67.995 ;
        RECT 64.095 67.445 64.265 67.735 ;
        RECT 63.600 67.275 64.265 67.445 ;
        RECT 63.600 66.285 63.830 67.275 ;
        RECT 64.985 67.270 65.275 67.995 ;
        RECT 65.450 67.255 65.705 67.825 ;
        RECT 65.875 67.595 66.205 67.995 ;
        RECT 66.630 67.460 67.160 67.825 ;
        RECT 67.350 67.655 67.625 67.825 ;
        RECT 67.345 67.485 67.625 67.655 ;
        RECT 66.630 67.425 66.805 67.460 ;
        RECT 65.875 67.255 66.805 67.425 ;
        RECT 64.000 66.455 64.350 67.105 ;
        RECT 63.600 66.115 64.265 66.285 ;
        RECT 63.595 65.445 63.925 65.945 ;
        RECT 64.095 65.615 64.265 66.115 ;
        RECT 64.985 65.445 65.275 66.610 ;
        RECT 65.450 66.585 65.620 67.255 ;
        RECT 65.875 67.085 66.045 67.255 ;
        RECT 65.790 66.755 66.045 67.085 ;
        RECT 66.270 66.755 66.465 67.085 ;
        RECT 65.450 65.615 65.785 66.585 ;
        RECT 65.955 65.445 66.125 66.585 ;
        RECT 66.295 65.785 66.465 66.755 ;
        RECT 66.635 66.125 66.805 67.255 ;
        RECT 66.975 66.465 67.145 67.265 ;
        RECT 67.350 66.665 67.625 67.485 ;
        RECT 67.795 66.465 67.985 67.825 ;
        RECT 68.165 67.460 68.675 67.995 ;
        RECT 68.895 67.185 69.140 67.790 ;
        RECT 69.585 67.225 72.175 67.995 ;
        RECT 72.820 67.425 73.075 67.775 ;
        RECT 73.245 67.595 73.575 67.995 ;
        RECT 73.745 67.425 73.915 67.775 ;
        RECT 74.085 67.595 74.465 67.995 ;
        RECT 72.820 67.255 74.485 67.425 ;
        RECT 74.655 67.320 74.930 67.665 ;
        RECT 68.185 67.015 69.415 67.185 ;
        RECT 66.975 66.295 67.985 66.465 ;
        RECT 68.155 66.450 68.905 66.640 ;
        RECT 66.635 65.955 67.760 66.125 ;
        RECT 68.155 65.785 68.325 66.450 ;
        RECT 69.075 66.205 69.415 67.015 ;
        RECT 69.585 66.705 70.795 67.225 ;
        RECT 74.315 67.085 74.485 67.255 ;
        RECT 70.965 66.535 72.175 67.055 ;
        RECT 72.805 66.755 73.150 67.085 ;
        RECT 73.320 66.755 74.145 67.085 ;
        RECT 74.315 66.755 74.590 67.085 ;
        RECT 66.295 65.615 68.325 65.785 ;
        RECT 68.495 65.445 68.665 66.205 ;
        RECT 68.900 65.795 69.415 66.205 ;
        RECT 69.585 65.445 72.175 66.535 ;
        RECT 72.825 66.295 73.150 66.585 ;
        RECT 73.320 66.465 73.515 66.755 ;
        RECT 74.315 66.585 74.485 66.755 ;
        RECT 74.760 66.585 74.930 67.320 ;
        RECT 75.310 67.215 75.810 67.825 ;
        RECT 75.105 66.755 75.455 67.005 ;
        RECT 75.640 66.585 75.810 67.215 ;
        RECT 76.440 67.345 76.770 67.825 ;
        RECT 76.940 67.535 77.165 67.995 ;
        RECT 77.335 67.345 77.665 67.825 ;
        RECT 76.440 67.175 77.665 67.345 ;
        RECT 77.855 67.195 78.105 67.995 ;
        RECT 78.275 67.195 78.615 67.825 ;
        RECT 78.790 67.230 79.245 67.995 ;
        RECT 79.520 67.615 80.820 67.825 ;
        RECT 81.075 67.635 81.405 67.995 ;
        RECT 80.650 67.465 80.820 67.615 ;
        RECT 81.575 67.495 81.835 67.825 ;
        RECT 75.980 66.805 76.310 67.005 ;
        RECT 76.480 66.805 76.810 67.005 ;
        RECT 76.980 66.805 77.400 67.005 ;
        RECT 77.575 66.835 78.270 67.005 ;
        RECT 77.575 66.585 77.745 66.835 ;
        RECT 78.440 66.585 78.615 67.195 ;
        RECT 79.720 67.005 79.940 67.405 ;
        RECT 78.785 66.805 79.275 67.005 ;
        RECT 79.465 66.795 79.940 67.005 ;
        RECT 80.185 67.005 80.395 67.405 ;
        RECT 80.650 67.340 81.405 67.465 ;
        RECT 80.650 67.295 81.495 67.340 ;
        RECT 81.225 67.175 81.495 67.295 ;
        RECT 80.185 66.795 80.515 67.005 ;
        RECT 80.685 66.735 81.095 67.040 ;
        RECT 73.825 66.415 74.485 66.585 ;
        RECT 73.825 66.295 73.995 66.415 ;
        RECT 72.825 66.125 73.995 66.295 ;
        RECT 72.805 65.665 73.995 65.955 ;
        RECT 74.165 65.445 74.445 66.245 ;
        RECT 74.655 65.615 74.930 66.585 ;
        RECT 75.310 66.415 77.745 66.585 ;
        RECT 75.310 65.615 75.640 66.415 ;
        RECT 75.810 65.445 76.140 66.245 ;
        RECT 76.440 65.615 76.770 66.415 ;
        RECT 77.415 65.445 77.665 66.245 ;
        RECT 77.935 65.445 78.105 66.585 ;
        RECT 78.275 65.615 78.615 66.585 ;
        RECT 78.790 66.565 79.965 66.625 ;
        RECT 81.325 66.600 81.495 67.175 ;
        RECT 81.295 66.565 81.495 66.600 ;
        RECT 78.790 66.455 81.495 66.565 ;
        RECT 78.790 65.835 79.045 66.455 ;
        RECT 79.635 66.395 81.435 66.455 ;
        RECT 79.635 66.365 79.965 66.395 ;
        RECT 81.665 66.295 81.835 67.495 ;
        RECT 82.095 67.445 82.265 67.735 ;
        RECT 82.435 67.615 82.765 67.995 ;
        RECT 82.095 67.275 82.760 67.445 ;
        RECT 82.010 66.455 82.360 67.105 ;
        RECT 79.295 66.195 79.480 66.285 ;
        RECT 80.070 66.195 80.905 66.205 ;
        RECT 79.295 65.995 80.905 66.195 ;
        RECT 79.295 65.955 79.525 65.995 ;
        RECT 78.790 65.615 79.125 65.835 ;
        RECT 80.130 65.445 80.485 65.825 ;
        RECT 80.655 65.615 80.905 65.995 ;
        RECT 81.155 65.445 81.405 66.225 ;
        RECT 81.575 65.615 81.835 66.295 ;
        RECT 82.530 66.285 82.760 67.275 ;
        RECT 82.095 66.115 82.760 66.285 ;
        RECT 82.095 65.615 82.265 66.115 ;
        RECT 82.435 65.445 82.765 65.945 ;
        RECT 82.935 65.615 83.120 67.735 ;
        RECT 83.375 67.535 83.625 67.995 ;
        RECT 83.795 67.545 84.130 67.715 ;
        RECT 84.325 67.545 85.000 67.715 ;
        RECT 83.795 67.405 83.965 67.545 ;
        RECT 83.290 66.415 83.570 67.365 ;
        RECT 83.740 67.275 83.965 67.405 ;
        RECT 83.740 66.170 83.910 67.275 ;
        RECT 84.135 67.125 84.660 67.345 ;
        RECT 84.080 66.360 84.320 66.955 ;
        RECT 84.490 66.425 84.660 67.125 ;
        RECT 84.830 66.765 85.000 67.545 ;
        RECT 85.320 67.495 85.690 67.995 ;
        RECT 85.870 67.545 86.275 67.715 ;
        RECT 86.445 67.545 87.230 67.715 ;
        RECT 85.870 67.315 86.040 67.545 ;
        RECT 85.210 67.015 86.040 67.315 ;
        RECT 86.425 67.045 86.890 67.375 ;
        RECT 85.210 66.985 85.410 67.015 ;
        RECT 85.530 66.765 85.700 66.835 ;
        RECT 84.830 66.595 85.700 66.765 ;
        RECT 85.190 66.505 85.700 66.595 ;
        RECT 83.740 66.040 84.045 66.170 ;
        RECT 84.490 66.060 85.020 66.425 ;
        RECT 83.360 65.445 83.625 65.905 ;
        RECT 83.795 65.615 84.045 66.040 ;
        RECT 85.190 65.890 85.360 66.505 ;
        RECT 84.255 65.720 85.360 65.890 ;
        RECT 85.530 65.445 85.700 66.245 ;
        RECT 85.870 65.945 86.040 67.015 ;
        RECT 86.210 66.115 86.400 66.835 ;
        RECT 86.570 66.085 86.890 67.045 ;
        RECT 87.060 67.085 87.230 67.545 ;
        RECT 87.505 67.465 87.715 67.995 ;
        RECT 87.975 67.255 88.305 67.780 ;
        RECT 88.475 67.385 88.645 67.995 ;
        RECT 88.815 67.340 89.145 67.775 ;
        RECT 88.815 67.255 89.195 67.340 ;
        RECT 88.105 67.085 88.305 67.255 ;
        RECT 88.970 67.215 89.195 67.255 ;
        RECT 87.060 66.755 87.935 67.085 ;
        RECT 88.105 66.755 88.855 67.085 ;
        RECT 85.870 65.615 86.120 65.945 ;
        RECT 87.060 65.915 87.230 66.755 ;
        RECT 88.105 66.550 88.295 66.755 ;
        RECT 89.025 66.635 89.195 67.215 ;
        RECT 88.980 66.585 89.195 66.635 ;
        RECT 87.400 66.175 88.295 66.550 ;
        RECT 88.805 66.505 89.195 66.585 ;
        RECT 89.365 67.320 89.625 67.825 ;
        RECT 89.805 67.615 90.135 67.995 ;
        RECT 90.315 67.445 90.485 67.825 ;
        RECT 89.365 66.520 89.535 67.320 ;
        RECT 89.820 67.275 90.485 67.445 ;
        RECT 89.820 67.020 89.990 67.275 ;
        RECT 90.745 67.245 91.955 67.995 ;
        RECT 89.705 66.690 89.990 67.020 ;
        RECT 90.225 66.725 90.555 67.095 ;
        RECT 89.820 66.545 89.990 66.690 ;
        RECT 86.345 65.745 87.230 65.915 ;
        RECT 87.410 65.445 87.725 65.945 ;
        RECT 87.955 65.615 88.295 66.175 ;
        RECT 88.465 65.445 88.635 66.455 ;
        RECT 88.805 65.660 89.135 66.505 ;
        RECT 89.365 65.615 89.635 66.520 ;
        RECT 89.820 66.375 90.485 66.545 ;
        RECT 89.805 65.445 90.135 66.205 ;
        RECT 90.315 65.615 90.485 66.375 ;
        RECT 90.745 66.535 91.265 67.075 ;
        RECT 91.435 66.705 91.955 67.245 ;
        RECT 90.745 65.445 91.955 66.535 ;
        RECT 13.380 65.275 92.040 65.445 ;
        RECT 13.465 64.185 14.675 65.275 ;
        RECT 13.465 63.475 13.985 64.015 ;
        RECT 14.155 63.645 14.675 64.185 ;
        RECT 14.850 64.125 15.110 65.275 ;
        RECT 15.285 64.200 15.540 65.105 ;
        RECT 15.710 64.515 16.040 65.275 ;
        RECT 16.255 64.345 16.425 65.105 ;
        RECT 13.465 62.725 14.675 63.475 ;
        RECT 14.850 62.725 15.110 63.565 ;
        RECT 15.285 63.470 15.455 64.200 ;
        RECT 15.710 64.175 16.425 64.345 ;
        RECT 15.710 63.965 15.880 64.175 ;
        RECT 16.690 64.125 16.950 65.275 ;
        RECT 17.125 64.200 17.380 65.105 ;
        RECT 17.550 64.515 17.880 65.275 ;
        RECT 18.095 64.345 18.265 65.105 ;
        RECT 15.625 63.635 15.880 63.965 ;
        RECT 15.285 62.895 15.540 63.470 ;
        RECT 15.710 63.445 15.880 63.635 ;
        RECT 16.160 63.625 16.515 63.995 ;
        RECT 15.710 63.275 16.425 63.445 ;
        RECT 15.710 62.725 16.040 63.105 ;
        RECT 16.255 62.895 16.425 63.275 ;
        RECT 16.690 62.725 16.950 63.565 ;
        RECT 17.125 63.470 17.295 64.200 ;
        RECT 17.550 64.175 18.265 64.345 ;
        RECT 18.525 64.185 19.735 65.275 ;
        RECT 17.550 63.965 17.720 64.175 ;
        RECT 17.465 63.635 17.720 63.965 ;
        RECT 17.125 62.895 17.380 63.470 ;
        RECT 17.550 63.445 17.720 63.635 ;
        RECT 18.000 63.625 18.355 63.995 ;
        RECT 18.525 63.475 19.045 64.015 ;
        RECT 19.215 63.645 19.735 64.185 ;
        RECT 19.910 64.125 20.170 65.275 ;
        RECT 20.345 64.200 20.600 65.105 ;
        RECT 20.770 64.515 21.100 65.275 ;
        RECT 21.315 64.345 21.485 65.105 ;
        RECT 17.550 63.275 18.265 63.445 ;
        RECT 17.550 62.725 17.880 63.105 ;
        RECT 18.095 62.895 18.265 63.275 ;
        RECT 18.525 62.725 19.735 63.475 ;
        RECT 19.910 62.725 20.170 63.565 ;
        RECT 20.345 63.470 20.515 64.200 ;
        RECT 20.770 64.175 21.485 64.345 ;
        RECT 21.745 64.185 25.255 65.275 ;
        RECT 20.770 63.965 20.940 64.175 ;
        RECT 20.685 63.635 20.940 63.965 ;
        RECT 20.345 62.895 20.600 63.470 ;
        RECT 20.770 63.445 20.940 63.635 ;
        RECT 21.220 63.625 21.575 63.995 ;
        RECT 21.745 63.495 23.395 64.015 ;
        RECT 23.565 63.665 25.255 64.185 ;
        RECT 26.345 64.110 26.635 65.275 ;
        RECT 26.805 64.135 27.145 65.105 ;
        RECT 27.315 64.135 27.485 65.275 ;
        RECT 27.755 64.475 28.005 65.275 ;
        RECT 28.650 64.305 28.980 65.105 ;
        RECT 29.280 64.475 29.610 65.275 ;
        RECT 29.780 64.305 30.110 65.105 ;
        RECT 27.675 64.135 30.110 64.305 ;
        RECT 30.670 64.305 31.060 64.480 ;
        RECT 31.545 64.475 31.875 65.275 ;
        RECT 32.045 64.485 32.580 65.105 ;
        RECT 30.670 64.135 32.095 64.305 ;
        RECT 26.805 63.525 26.980 64.135 ;
        RECT 27.675 63.885 27.845 64.135 ;
        RECT 27.150 63.715 27.845 63.885 ;
        RECT 28.020 63.715 28.440 63.915 ;
        RECT 28.610 63.715 28.940 63.915 ;
        RECT 29.110 63.715 29.440 63.915 ;
        RECT 20.770 63.275 21.485 63.445 ;
        RECT 20.770 62.725 21.100 63.105 ;
        RECT 21.315 62.895 21.485 63.275 ;
        RECT 21.745 62.725 25.255 63.495 ;
        RECT 26.345 62.725 26.635 63.450 ;
        RECT 26.805 62.895 27.145 63.525 ;
        RECT 27.315 62.725 27.565 63.525 ;
        RECT 27.755 63.375 28.980 63.545 ;
        RECT 27.755 62.895 28.085 63.375 ;
        RECT 28.255 62.725 28.480 63.185 ;
        RECT 28.650 62.895 28.980 63.375 ;
        RECT 29.610 63.505 29.780 64.135 ;
        RECT 29.965 63.715 30.315 63.965 ;
        RECT 29.610 62.895 30.110 63.505 ;
        RECT 30.545 63.405 30.900 63.965 ;
        RECT 31.070 63.235 31.240 64.135 ;
        RECT 31.410 63.405 31.675 63.965 ;
        RECT 31.925 63.635 32.095 64.135 ;
        RECT 32.265 63.465 32.580 64.485 ;
        RECT 32.785 64.185 34.455 65.275 ;
        RECT 34.715 64.605 34.885 65.105 ;
        RECT 35.055 64.775 35.385 65.275 ;
        RECT 34.715 64.435 35.380 64.605 ;
        RECT 30.650 62.725 30.890 63.235 ;
        RECT 31.070 62.905 31.350 63.235 ;
        RECT 31.580 62.725 31.795 63.235 ;
        RECT 31.965 62.895 32.580 63.465 ;
        RECT 32.785 63.495 33.535 64.015 ;
        RECT 33.705 63.665 34.455 64.185 ;
        RECT 34.630 63.615 34.980 64.265 ;
        RECT 32.785 62.725 34.455 63.495 ;
        RECT 35.150 63.445 35.380 64.435 ;
        RECT 34.715 63.275 35.380 63.445 ;
        RECT 34.715 62.985 34.885 63.275 ;
        RECT 35.055 62.725 35.385 63.105 ;
        RECT 35.555 62.985 35.740 65.105 ;
        RECT 35.980 64.815 36.245 65.275 ;
        RECT 36.415 64.680 36.665 65.105 ;
        RECT 36.875 64.830 37.980 65.000 ;
        RECT 36.360 64.550 36.665 64.680 ;
        RECT 35.910 63.355 36.190 64.305 ;
        RECT 36.360 63.445 36.530 64.550 ;
        RECT 36.700 63.765 36.940 64.360 ;
        RECT 37.110 64.295 37.640 64.660 ;
        RECT 37.110 63.595 37.280 64.295 ;
        RECT 37.810 64.215 37.980 64.830 ;
        RECT 38.150 64.475 38.320 65.275 ;
        RECT 38.490 64.775 38.740 65.105 ;
        RECT 38.965 64.805 39.850 64.975 ;
        RECT 37.810 64.125 38.320 64.215 ;
        RECT 36.360 63.315 36.585 63.445 ;
        RECT 36.755 63.375 37.280 63.595 ;
        RECT 37.450 63.955 38.320 64.125 ;
        RECT 35.995 62.725 36.245 63.185 ;
        RECT 36.415 63.175 36.585 63.315 ;
        RECT 37.450 63.175 37.620 63.955 ;
        RECT 38.150 63.885 38.320 63.955 ;
        RECT 37.830 63.705 38.030 63.735 ;
        RECT 38.490 63.705 38.660 64.775 ;
        RECT 38.830 63.885 39.020 64.605 ;
        RECT 37.830 63.405 38.660 63.705 ;
        RECT 39.190 63.675 39.510 64.635 ;
        RECT 36.415 63.005 36.750 63.175 ;
        RECT 36.945 63.005 37.620 63.175 ;
        RECT 37.940 62.725 38.310 63.225 ;
        RECT 38.490 63.175 38.660 63.405 ;
        RECT 39.045 63.345 39.510 63.675 ;
        RECT 39.680 63.965 39.850 64.805 ;
        RECT 40.030 64.775 40.345 65.275 ;
        RECT 40.575 64.545 40.915 65.105 ;
        RECT 40.020 64.170 40.915 64.545 ;
        RECT 41.085 64.265 41.255 65.275 ;
        RECT 40.725 63.965 40.915 64.170 ;
        RECT 41.425 64.215 41.755 65.060 ;
        RECT 41.425 64.135 41.815 64.215 ;
        RECT 41.985 64.185 44.575 65.275 ;
        RECT 41.600 64.085 41.815 64.135 ;
        RECT 39.680 63.635 40.555 63.965 ;
        RECT 40.725 63.635 41.475 63.965 ;
        RECT 39.680 63.175 39.850 63.635 ;
        RECT 40.725 63.465 40.925 63.635 ;
        RECT 41.645 63.505 41.815 64.085 ;
        RECT 41.590 63.465 41.815 63.505 ;
        RECT 38.490 63.005 38.895 63.175 ;
        RECT 39.065 63.005 39.850 63.175 ;
        RECT 40.125 62.725 40.335 63.255 ;
        RECT 40.595 62.940 40.925 63.465 ;
        RECT 41.435 63.380 41.815 63.465 ;
        RECT 41.985 63.495 43.195 64.015 ;
        RECT 43.365 63.665 44.575 64.185 ;
        RECT 44.750 64.135 45.085 65.105 ;
        RECT 45.255 64.135 45.425 65.275 ;
        RECT 45.595 64.935 47.625 65.105 ;
        RECT 41.095 62.725 41.265 63.335 ;
        RECT 41.435 62.945 41.765 63.380 ;
        RECT 41.985 62.725 44.575 63.495 ;
        RECT 44.750 63.465 44.920 64.135 ;
        RECT 45.595 63.965 45.765 64.935 ;
        RECT 45.090 63.635 45.345 63.965 ;
        RECT 45.570 63.635 45.765 63.965 ;
        RECT 45.935 64.595 47.060 64.765 ;
        RECT 45.175 63.465 45.345 63.635 ;
        RECT 45.935 63.465 46.105 64.595 ;
        RECT 44.750 62.895 45.005 63.465 ;
        RECT 45.175 63.295 46.105 63.465 ;
        RECT 46.275 64.255 47.285 64.425 ;
        RECT 46.275 63.455 46.445 64.255 ;
        RECT 46.650 63.915 46.925 64.055 ;
        RECT 46.645 63.745 46.925 63.915 ;
        RECT 45.930 63.260 46.105 63.295 ;
        RECT 45.175 62.725 45.505 63.125 ;
        RECT 45.930 62.895 46.460 63.260 ;
        RECT 46.650 62.895 46.925 63.745 ;
        RECT 47.095 62.895 47.285 64.255 ;
        RECT 47.455 64.270 47.625 64.935 ;
        RECT 47.795 64.515 47.965 65.275 ;
        RECT 48.200 64.515 48.715 64.925 ;
        RECT 47.455 64.080 48.205 64.270 ;
        RECT 48.375 63.705 48.715 64.515 ;
        RECT 49.400 64.405 49.685 65.275 ;
        RECT 49.855 64.645 50.115 65.105 ;
        RECT 50.290 64.815 50.545 65.275 ;
        RECT 50.715 64.645 50.975 65.105 ;
        RECT 49.855 64.475 50.975 64.645 ;
        RECT 51.145 64.475 51.455 65.275 ;
        RECT 49.855 64.225 50.115 64.475 ;
        RECT 51.625 64.305 51.935 65.105 ;
        RECT 47.485 63.535 48.715 63.705 ;
        RECT 49.360 64.055 50.115 64.225 ;
        RECT 50.905 64.135 51.935 64.305 ;
        RECT 49.360 63.545 49.765 64.055 ;
        RECT 50.905 63.885 51.075 64.135 ;
        RECT 49.935 63.715 51.075 63.885 ;
        RECT 47.465 62.725 47.975 63.260 ;
        RECT 48.195 62.930 48.440 63.535 ;
        RECT 49.360 63.375 51.010 63.545 ;
        RECT 51.245 63.395 51.595 63.965 ;
        RECT 49.405 62.725 49.685 63.205 ;
        RECT 49.855 62.985 50.115 63.375 ;
        RECT 50.290 62.725 50.545 63.205 ;
        RECT 50.715 62.985 51.010 63.375 ;
        RECT 51.765 63.225 51.935 64.135 ;
        RECT 52.105 64.110 52.395 65.275 ;
        RECT 52.655 64.605 52.825 65.105 ;
        RECT 52.995 64.775 53.325 65.275 ;
        RECT 52.655 64.435 53.320 64.605 ;
        RECT 52.570 63.615 52.920 64.265 ;
        RECT 51.190 62.725 51.465 63.205 ;
        RECT 51.635 62.895 51.935 63.225 ;
        RECT 52.105 62.725 52.395 63.450 ;
        RECT 53.090 63.445 53.320 64.435 ;
        RECT 52.655 63.275 53.320 63.445 ;
        RECT 52.655 62.985 52.825 63.275 ;
        RECT 52.995 62.725 53.325 63.105 ;
        RECT 53.495 62.985 53.680 65.105 ;
        RECT 53.920 64.815 54.185 65.275 ;
        RECT 54.355 64.680 54.605 65.105 ;
        RECT 54.815 64.830 55.920 65.000 ;
        RECT 54.300 64.550 54.605 64.680 ;
        RECT 53.850 63.355 54.130 64.305 ;
        RECT 54.300 63.445 54.470 64.550 ;
        RECT 54.640 63.765 54.880 64.360 ;
        RECT 55.050 64.295 55.580 64.660 ;
        RECT 55.050 63.595 55.220 64.295 ;
        RECT 55.750 64.215 55.920 64.830 ;
        RECT 56.090 64.475 56.260 65.275 ;
        RECT 56.430 64.775 56.680 65.105 ;
        RECT 56.905 64.805 57.790 64.975 ;
        RECT 55.750 64.125 56.260 64.215 ;
        RECT 54.300 63.315 54.525 63.445 ;
        RECT 54.695 63.375 55.220 63.595 ;
        RECT 55.390 63.955 56.260 64.125 ;
        RECT 53.935 62.725 54.185 63.185 ;
        RECT 54.355 63.175 54.525 63.315 ;
        RECT 55.390 63.175 55.560 63.955 ;
        RECT 56.090 63.885 56.260 63.955 ;
        RECT 55.770 63.705 55.970 63.735 ;
        RECT 56.430 63.705 56.600 64.775 ;
        RECT 56.770 63.885 56.960 64.605 ;
        RECT 55.770 63.405 56.600 63.705 ;
        RECT 57.130 63.675 57.450 64.635 ;
        RECT 54.355 63.005 54.690 63.175 ;
        RECT 54.885 63.005 55.560 63.175 ;
        RECT 55.880 62.725 56.250 63.225 ;
        RECT 56.430 63.175 56.600 63.405 ;
        RECT 56.985 63.345 57.450 63.675 ;
        RECT 57.620 63.965 57.790 64.805 ;
        RECT 57.970 64.775 58.285 65.275 ;
        RECT 58.515 64.545 58.855 65.105 ;
        RECT 57.960 64.170 58.855 64.545 ;
        RECT 59.025 64.265 59.195 65.275 ;
        RECT 58.665 63.965 58.855 64.170 ;
        RECT 59.365 64.215 59.695 65.060 ;
        RECT 59.365 64.135 59.755 64.215 ;
        RECT 59.540 64.085 59.755 64.135 ;
        RECT 57.620 63.635 58.495 63.965 ;
        RECT 58.665 63.635 59.415 63.965 ;
        RECT 57.620 63.175 57.790 63.635 ;
        RECT 58.665 63.465 58.865 63.635 ;
        RECT 59.585 63.505 59.755 64.085 ;
        RECT 59.530 63.465 59.755 63.505 ;
        RECT 56.430 63.005 56.835 63.175 ;
        RECT 57.005 63.005 57.790 63.175 ;
        RECT 58.065 62.725 58.275 63.255 ;
        RECT 58.535 62.940 58.865 63.465 ;
        RECT 59.375 63.380 59.755 63.465 ;
        RECT 59.925 64.135 60.310 65.105 ;
        RECT 60.480 64.815 60.805 65.275 ;
        RECT 61.325 64.645 61.605 65.105 ;
        RECT 60.480 64.425 61.605 64.645 ;
        RECT 59.925 63.465 60.205 64.135 ;
        RECT 60.480 63.965 60.930 64.425 ;
        RECT 61.795 64.255 62.195 65.105 ;
        RECT 62.595 64.815 62.865 65.275 ;
        RECT 63.035 64.645 63.320 65.105 ;
        RECT 60.375 63.635 60.930 63.965 ;
        RECT 61.100 63.695 62.195 64.255 ;
        RECT 60.480 63.525 60.930 63.635 ;
        RECT 59.035 62.725 59.205 63.335 ;
        RECT 59.375 62.945 59.705 63.380 ;
        RECT 59.925 62.895 60.310 63.465 ;
        RECT 60.480 63.355 61.605 63.525 ;
        RECT 60.480 62.725 60.805 63.185 ;
        RECT 61.325 62.895 61.605 63.355 ;
        RECT 61.795 62.895 62.195 63.695 ;
        RECT 62.365 64.425 63.320 64.645 ;
        RECT 63.720 64.645 64.005 65.105 ;
        RECT 64.175 64.815 64.445 65.275 ;
        RECT 63.720 64.425 64.675 64.645 ;
        RECT 62.365 63.525 62.575 64.425 ;
        RECT 62.745 63.695 63.435 64.255 ;
        RECT 63.605 63.695 64.295 64.255 ;
        RECT 64.465 63.525 64.675 64.425 ;
        RECT 62.365 63.355 63.320 63.525 ;
        RECT 62.595 62.725 62.865 63.185 ;
        RECT 63.035 62.895 63.320 63.355 ;
        RECT 63.720 63.355 64.675 63.525 ;
        RECT 64.845 64.255 65.245 65.105 ;
        RECT 65.435 64.645 65.715 65.105 ;
        RECT 66.235 64.815 66.560 65.275 ;
        RECT 65.435 64.425 66.560 64.645 ;
        RECT 64.845 63.695 65.940 64.255 ;
        RECT 66.110 63.965 66.560 64.425 ;
        RECT 66.730 64.135 67.115 65.105 ;
        RECT 67.290 64.475 67.545 65.275 ;
        RECT 67.745 64.425 68.075 65.105 ;
        RECT 63.720 62.895 64.005 63.355 ;
        RECT 64.175 62.725 64.445 63.185 ;
        RECT 64.845 62.895 65.245 63.695 ;
        RECT 66.110 63.635 66.665 63.965 ;
        RECT 66.110 63.525 66.560 63.635 ;
        RECT 65.435 63.355 66.560 63.525 ;
        RECT 66.835 63.465 67.115 64.135 ;
        RECT 67.290 63.935 67.535 64.295 ;
        RECT 67.725 64.145 68.075 64.425 ;
        RECT 67.725 63.765 67.895 64.145 ;
        RECT 68.255 63.965 68.450 65.015 ;
        RECT 68.630 64.135 68.950 65.275 ;
        RECT 70.055 64.165 70.350 65.275 ;
        RECT 70.530 63.965 70.780 65.100 ;
        RECT 70.950 64.165 71.210 65.275 ;
        RECT 71.380 64.375 71.640 65.100 ;
        RECT 71.810 64.545 72.070 65.275 ;
        RECT 72.240 64.375 72.500 65.100 ;
        RECT 72.670 64.545 72.930 65.275 ;
        RECT 73.100 64.375 73.360 65.100 ;
        RECT 73.530 64.545 73.790 65.275 ;
        RECT 73.960 64.375 74.220 65.100 ;
        RECT 74.390 64.545 74.685 65.275 ;
        RECT 71.380 64.135 74.690 64.375 ;
        RECT 75.750 64.305 76.140 64.480 ;
        RECT 76.625 64.475 76.955 65.275 ;
        RECT 77.125 64.485 77.660 65.105 ;
        RECT 75.750 64.135 77.175 64.305 ;
        RECT 65.435 62.895 65.715 63.355 ;
        RECT 66.235 62.725 66.560 63.185 ;
        RECT 66.730 62.895 67.115 63.465 ;
        RECT 67.375 63.595 67.895 63.765 ;
        RECT 68.065 63.635 68.450 63.965 ;
        RECT 68.630 63.915 68.890 63.965 ;
        RECT 68.630 63.745 68.895 63.915 ;
        RECT 68.630 63.635 68.890 63.745 ;
        RECT 67.375 63.235 67.545 63.595 ;
        RECT 67.345 63.065 67.545 63.235 ;
        RECT 67.375 63.030 67.545 63.065 ;
        RECT 67.735 63.255 68.950 63.425 ;
        RECT 70.045 63.355 70.360 63.965 ;
        RECT 70.530 63.715 73.550 63.965 ;
        RECT 67.735 62.950 67.965 63.255 ;
        RECT 68.135 62.725 68.465 63.085 ;
        RECT 68.660 62.905 68.950 63.255 ;
        RECT 70.105 62.725 70.350 63.185 ;
        RECT 70.530 62.905 70.780 63.715 ;
        RECT 73.720 63.545 74.690 64.135 ;
        RECT 71.380 63.375 74.690 63.545 ;
        RECT 75.625 63.405 75.980 63.965 ;
        RECT 70.950 62.725 71.210 63.250 ;
        RECT 71.380 62.920 71.640 63.375 ;
        RECT 71.810 62.725 72.070 63.205 ;
        RECT 72.240 62.920 72.500 63.375 ;
        RECT 72.670 62.725 72.930 63.205 ;
        RECT 73.100 62.920 73.360 63.375 ;
        RECT 73.530 62.725 73.790 63.205 ;
        RECT 73.960 62.920 74.220 63.375 ;
        RECT 76.150 63.235 76.320 64.135 ;
        RECT 76.490 63.405 76.755 63.965 ;
        RECT 77.005 63.635 77.175 64.135 ;
        RECT 77.345 63.465 77.660 64.485 ;
        RECT 77.865 64.110 78.155 65.275 ;
        RECT 78.325 64.185 79.995 65.275 ;
        RECT 80.280 64.645 80.565 65.105 ;
        RECT 80.735 64.815 81.005 65.275 ;
        RECT 80.280 64.425 81.235 64.645 ;
        RECT 74.390 62.725 74.690 63.205 ;
        RECT 75.730 62.725 75.970 63.235 ;
        RECT 76.150 62.905 76.430 63.235 ;
        RECT 76.660 62.725 76.875 63.235 ;
        RECT 77.045 62.895 77.660 63.465 ;
        RECT 78.325 63.495 79.075 64.015 ;
        RECT 79.245 63.665 79.995 64.185 ;
        RECT 80.165 63.695 80.855 64.255 ;
        RECT 81.025 63.525 81.235 64.425 ;
        RECT 77.865 62.725 78.155 63.450 ;
        RECT 78.325 62.725 79.995 63.495 ;
        RECT 80.280 63.355 81.235 63.525 ;
        RECT 81.405 64.255 81.805 65.105 ;
        RECT 81.995 64.645 82.275 65.105 ;
        RECT 82.795 64.815 83.120 65.275 ;
        RECT 81.995 64.425 83.120 64.645 ;
        RECT 81.405 63.695 82.500 64.255 ;
        RECT 82.670 63.965 83.120 64.425 ;
        RECT 83.290 64.135 83.675 65.105 ;
        RECT 80.280 62.895 80.565 63.355 ;
        RECT 80.735 62.725 81.005 63.185 ;
        RECT 81.405 62.895 81.805 63.695 ;
        RECT 82.670 63.635 83.225 63.965 ;
        RECT 82.670 63.525 83.120 63.635 ;
        RECT 81.995 63.355 83.120 63.525 ;
        RECT 83.395 63.465 83.675 64.135 ;
        RECT 81.995 62.895 82.275 63.355 ;
        RECT 82.795 62.725 83.120 63.185 ;
        RECT 83.290 62.895 83.675 63.465 ;
        RECT 83.850 64.135 84.185 65.105 ;
        RECT 84.355 64.135 84.525 65.275 ;
        RECT 84.695 64.935 86.725 65.105 ;
        RECT 83.850 63.465 84.020 64.135 ;
        RECT 84.695 63.965 84.865 64.935 ;
        RECT 84.190 63.635 84.445 63.965 ;
        RECT 84.670 63.635 84.865 63.965 ;
        RECT 85.035 64.595 86.160 64.765 ;
        RECT 84.275 63.465 84.445 63.635 ;
        RECT 85.035 63.465 85.205 64.595 ;
        RECT 83.850 62.895 84.105 63.465 ;
        RECT 84.275 63.295 85.205 63.465 ;
        RECT 85.375 64.255 86.385 64.425 ;
        RECT 85.375 63.455 85.545 64.255 ;
        RECT 85.750 63.575 86.025 64.055 ;
        RECT 85.745 63.405 86.025 63.575 ;
        RECT 85.030 63.260 85.205 63.295 ;
        RECT 84.275 62.725 84.605 63.125 ;
        RECT 85.030 62.895 85.560 63.260 ;
        RECT 85.750 62.895 86.025 63.405 ;
        RECT 86.195 62.895 86.385 64.255 ;
        RECT 86.555 64.270 86.725 64.935 ;
        RECT 86.895 64.515 87.065 65.275 ;
        RECT 87.300 64.515 87.815 64.925 ;
        RECT 86.555 64.080 87.305 64.270 ;
        RECT 87.475 63.705 87.815 64.515 ;
        RECT 88.995 64.345 89.165 65.105 ;
        RECT 89.380 64.515 89.710 65.275 ;
        RECT 88.995 64.175 89.710 64.345 ;
        RECT 89.880 64.200 90.135 65.105 ;
        RECT 86.585 63.535 87.815 63.705 ;
        RECT 88.905 63.625 89.260 63.995 ;
        RECT 89.540 63.965 89.710 64.175 ;
        RECT 89.540 63.635 89.795 63.965 ;
        RECT 86.565 62.725 87.075 63.260 ;
        RECT 87.295 62.930 87.540 63.535 ;
        RECT 89.540 63.445 89.710 63.635 ;
        RECT 89.965 63.470 90.135 64.200 ;
        RECT 90.310 64.125 90.570 65.275 ;
        RECT 90.745 64.185 91.955 65.275 ;
        RECT 90.745 63.645 91.265 64.185 ;
        RECT 88.995 63.275 89.710 63.445 ;
        RECT 88.995 62.895 89.165 63.275 ;
        RECT 89.380 62.725 89.710 63.105 ;
        RECT 89.880 62.895 90.135 63.470 ;
        RECT 90.310 62.725 90.570 63.565 ;
        RECT 91.435 63.475 91.955 64.015 ;
        RECT 90.745 62.725 91.955 63.475 ;
        RECT 13.380 62.555 92.040 62.725 ;
        RECT 13.465 61.805 14.675 62.555 ;
        RECT 14.845 61.805 16.055 62.555 ;
        RECT 16.390 62.045 16.630 62.555 ;
        RECT 16.810 62.045 17.090 62.375 ;
        RECT 17.320 62.045 17.535 62.555 ;
        RECT 13.465 61.265 13.985 61.805 ;
        RECT 14.155 61.095 14.675 61.635 ;
        RECT 14.845 61.265 15.365 61.805 ;
        RECT 15.535 61.095 16.055 61.635 ;
        RECT 16.285 61.315 16.640 61.875 ;
        RECT 16.810 61.145 16.980 62.045 ;
        RECT 17.150 61.315 17.415 61.875 ;
        RECT 17.705 61.815 18.320 62.385 ;
        RECT 17.665 61.145 17.835 61.645 ;
        RECT 13.465 60.005 14.675 61.095 ;
        RECT 14.845 60.005 16.055 61.095 ;
        RECT 16.410 60.975 17.835 61.145 ;
        RECT 16.410 60.800 16.800 60.975 ;
        RECT 17.285 60.005 17.615 60.805 ;
        RECT 18.005 60.795 18.320 61.815 ;
        RECT 18.525 61.805 19.735 62.555 ;
        RECT 19.905 61.815 20.165 62.385 ;
        RECT 20.335 62.155 20.720 62.555 ;
        RECT 20.890 61.985 21.145 62.385 ;
        RECT 20.335 61.815 21.145 61.985 ;
        RECT 21.335 61.815 21.580 62.385 ;
        RECT 21.750 62.155 22.135 62.555 ;
        RECT 22.305 61.985 22.560 62.385 ;
        RECT 21.750 61.815 22.560 61.985 ;
        RECT 22.750 61.815 23.175 62.385 ;
        RECT 23.345 62.155 23.730 62.555 ;
        RECT 23.900 61.985 24.335 62.385 ;
        RECT 23.345 61.815 24.335 61.985 ;
        RECT 24.595 62.005 24.765 62.295 ;
        RECT 24.935 62.175 25.265 62.555 ;
        RECT 24.595 61.835 25.260 62.005 ;
        RECT 18.525 61.265 19.045 61.805 ;
        RECT 19.215 61.095 19.735 61.635 ;
        RECT 17.785 60.175 18.320 60.795 ;
        RECT 18.525 60.005 19.735 61.095 ;
        RECT 19.905 61.145 20.090 61.815 ;
        RECT 20.335 61.645 20.685 61.815 ;
        RECT 21.335 61.645 21.505 61.815 ;
        RECT 21.750 61.645 22.100 61.815 ;
        RECT 22.750 61.645 23.100 61.815 ;
        RECT 23.345 61.645 23.680 61.815 ;
        RECT 20.260 61.315 20.685 61.645 ;
        RECT 19.905 60.175 20.165 61.145 ;
        RECT 20.335 60.795 20.685 61.315 ;
        RECT 20.855 61.145 21.505 61.645 ;
        RECT 21.675 61.315 22.100 61.645 ;
        RECT 20.855 60.965 21.580 61.145 ;
        RECT 20.335 60.600 21.145 60.795 ;
        RECT 20.335 60.005 20.720 60.430 ;
        RECT 20.890 60.175 21.145 60.600 ;
        RECT 21.335 60.175 21.580 60.965 ;
        RECT 21.750 60.795 22.100 61.315 ;
        RECT 22.270 61.145 23.100 61.645 ;
        RECT 23.270 61.315 23.680 61.645 ;
        RECT 22.270 60.965 23.175 61.145 ;
        RECT 21.750 60.600 22.580 60.795 ;
        RECT 21.750 60.005 22.135 60.430 ;
        RECT 22.305 60.175 22.580 60.600 ;
        RECT 22.750 60.175 23.175 60.965 ;
        RECT 23.345 60.770 23.680 61.315 ;
        RECT 23.850 60.940 24.335 61.645 ;
        RECT 24.510 61.015 24.860 61.665 ;
        RECT 25.030 60.845 25.260 61.835 ;
        RECT 23.345 60.600 24.335 60.770 ;
        RECT 23.345 60.005 23.730 60.430 ;
        RECT 23.900 60.175 24.335 60.600 ;
        RECT 24.595 60.675 25.260 60.845 ;
        RECT 24.595 60.175 24.765 60.675 ;
        RECT 24.935 60.005 25.265 60.505 ;
        RECT 25.435 60.175 25.620 62.295 ;
        RECT 25.875 62.095 26.125 62.555 ;
        RECT 26.295 62.105 26.630 62.275 ;
        RECT 26.825 62.105 27.500 62.275 ;
        RECT 26.295 61.965 26.465 62.105 ;
        RECT 25.790 60.975 26.070 61.925 ;
        RECT 26.240 61.835 26.465 61.965 ;
        RECT 26.240 60.730 26.410 61.835 ;
        RECT 26.635 61.685 27.160 61.905 ;
        RECT 26.580 60.920 26.820 61.515 ;
        RECT 26.990 60.985 27.160 61.685 ;
        RECT 27.330 61.325 27.500 62.105 ;
        RECT 27.820 62.055 28.190 62.555 ;
        RECT 28.370 62.105 28.775 62.275 ;
        RECT 28.945 62.105 29.730 62.275 ;
        RECT 28.370 61.875 28.540 62.105 ;
        RECT 27.710 61.575 28.540 61.875 ;
        RECT 28.925 61.605 29.390 61.935 ;
        RECT 27.710 61.545 27.910 61.575 ;
        RECT 28.030 61.325 28.200 61.395 ;
        RECT 27.330 61.155 28.200 61.325 ;
        RECT 27.690 61.065 28.200 61.155 ;
        RECT 26.240 60.600 26.545 60.730 ;
        RECT 26.990 60.620 27.520 60.985 ;
        RECT 25.860 60.005 26.125 60.465 ;
        RECT 26.295 60.175 26.545 60.600 ;
        RECT 27.690 60.450 27.860 61.065 ;
        RECT 26.755 60.280 27.860 60.450 ;
        RECT 28.030 60.005 28.200 60.805 ;
        RECT 28.370 60.505 28.540 61.575 ;
        RECT 28.710 60.675 28.900 61.395 ;
        RECT 29.070 60.645 29.390 61.605 ;
        RECT 29.560 61.645 29.730 62.105 ;
        RECT 30.005 62.025 30.215 62.555 ;
        RECT 30.475 61.815 30.805 62.340 ;
        RECT 30.975 61.945 31.145 62.555 ;
        RECT 31.315 61.900 31.645 62.335 ;
        RECT 31.955 62.005 32.125 62.295 ;
        RECT 32.295 62.175 32.625 62.555 ;
        RECT 31.315 61.815 31.695 61.900 ;
        RECT 31.955 61.835 32.620 62.005 ;
        RECT 30.605 61.645 30.805 61.815 ;
        RECT 31.470 61.775 31.695 61.815 ;
        RECT 29.560 61.315 30.435 61.645 ;
        RECT 30.605 61.315 31.355 61.645 ;
        RECT 28.370 60.175 28.620 60.505 ;
        RECT 29.560 60.475 29.730 61.315 ;
        RECT 30.605 61.110 30.795 61.315 ;
        RECT 31.525 61.195 31.695 61.775 ;
        RECT 31.480 61.145 31.695 61.195 ;
        RECT 29.900 60.735 30.795 61.110 ;
        RECT 31.305 61.065 31.695 61.145 ;
        RECT 28.845 60.305 29.730 60.475 ;
        RECT 29.910 60.005 30.225 60.505 ;
        RECT 30.455 60.175 30.795 60.735 ;
        RECT 30.965 60.005 31.135 61.015 ;
        RECT 31.305 60.220 31.635 61.065 ;
        RECT 31.870 61.015 32.220 61.665 ;
        RECT 32.390 60.845 32.620 61.835 ;
        RECT 31.955 60.675 32.620 60.845 ;
        RECT 31.955 60.175 32.125 60.675 ;
        RECT 32.295 60.005 32.625 60.505 ;
        RECT 32.795 60.175 32.980 62.295 ;
        RECT 33.235 62.095 33.485 62.555 ;
        RECT 33.655 62.105 33.990 62.275 ;
        RECT 34.185 62.105 34.860 62.275 ;
        RECT 33.655 61.965 33.825 62.105 ;
        RECT 33.150 60.975 33.430 61.925 ;
        RECT 33.600 61.835 33.825 61.965 ;
        RECT 33.600 60.730 33.770 61.835 ;
        RECT 33.995 61.685 34.520 61.905 ;
        RECT 33.940 60.920 34.180 61.515 ;
        RECT 34.350 60.985 34.520 61.685 ;
        RECT 34.690 61.325 34.860 62.105 ;
        RECT 35.180 62.055 35.550 62.555 ;
        RECT 35.730 62.105 36.135 62.275 ;
        RECT 36.305 62.105 37.090 62.275 ;
        RECT 35.730 61.875 35.900 62.105 ;
        RECT 35.070 61.575 35.900 61.875 ;
        RECT 36.285 61.605 36.750 61.935 ;
        RECT 35.070 61.545 35.270 61.575 ;
        RECT 35.390 61.325 35.560 61.395 ;
        RECT 34.690 61.155 35.560 61.325 ;
        RECT 35.050 61.065 35.560 61.155 ;
        RECT 33.600 60.600 33.905 60.730 ;
        RECT 34.350 60.620 34.880 60.985 ;
        RECT 33.220 60.005 33.485 60.465 ;
        RECT 33.655 60.175 33.905 60.600 ;
        RECT 35.050 60.450 35.220 61.065 ;
        RECT 34.115 60.280 35.220 60.450 ;
        RECT 35.390 60.005 35.560 60.805 ;
        RECT 35.730 60.505 35.900 61.575 ;
        RECT 36.070 60.675 36.260 61.395 ;
        RECT 36.430 60.645 36.750 61.605 ;
        RECT 36.920 61.645 37.090 62.105 ;
        RECT 37.365 62.025 37.575 62.555 ;
        RECT 37.835 61.815 38.165 62.340 ;
        RECT 38.335 61.945 38.505 62.555 ;
        RECT 38.675 61.900 39.005 62.335 ;
        RECT 38.675 61.815 39.055 61.900 ;
        RECT 39.225 61.830 39.515 62.555 ;
        RECT 37.965 61.645 38.165 61.815 ;
        RECT 38.830 61.775 39.055 61.815 ;
        RECT 36.920 61.315 37.795 61.645 ;
        RECT 37.965 61.315 38.715 61.645 ;
        RECT 35.730 60.175 35.980 60.505 ;
        RECT 36.920 60.475 37.090 61.315 ;
        RECT 37.965 61.110 38.155 61.315 ;
        RECT 38.885 61.195 39.055 61.775 ;
        RECT 39.685 61.785 42.275 62.555 ;
        RECT 42.535 62.005 42.705 62.295 ;
        RECT 42.875 62.175 43.205 62.555 ;
        RECT 42.535 61.835 43.200 62.005 ;
        RECT 39.685 61.265 40.895 61.785 ;
        RECT 38.840 61.145 39.055 61.195 ;
        RECT 37.260 60.735 38.155 61.110 ;
        RECT 38.665 61.065 39.055 61.145 ;
        RECT 36.205 60.305 37.090 60.475 ;
        RECT 37.270 60.005 37.585 60.505 ;
        RECT 37.815 60.175 38.155 60.735 ;
        RECT 38.325 60.005 38.495 61.015 ;
        RECT 38.665 60.220 38.995 61.065 ;
        RECT 39.225 60.005 39.515 61.170 ;
        RECT 41.065 61.095 42.275 61.615 ;
        RECT 39.685 60.005 42.275 61.095 ;
        RECT 42.450 61.015 42.800 61.665 ;
        RECT 42.970 60.845 43.200 61.835 ;
        RECT 42.535 60.675 43.200 60.845 ;
        RECT 42.535 60.175 42.705 60.675 ;
        RECT 42.875 60.005 43.205 60.505 ;
        RECT 43.375 60.175 43.560 62.295 ;
        RECT 43.815 62.095 44.065 62.555 ;
        RECT 44.235 62.105 44.570 62.275 ;
        RECT 44.765 62.105 45.440 62.275 ;
        RECT 44.235 61.965 44.405 62.105 ;
        RECT 43.730 60.975 44.010 61.925 ;
        RECT 44.180 61.835 44.405 61.965 ;
        RECT 44.180 60.730 44.350 61.835 ;
        RECT 44.575 61.685 45.100 61.905 ;
        RECT 44.520 60.920 44.760 61.515 ;
        RECT 44.930 60.985 45.100 61.685 ;
        RECT 45.270 61.325 45.440 62.105 ;
        RECT 45.760 62.055 46.130 62.555 ;
        RECT 46.310 62.105 46.715 62.275 ;
        RECT 46.885 62.105 47.670 62.275 ;
        RECT 46.310 61.875 46.480 62.105 ;
        RECT 45.650 61.575 46.480 61.875 ;
        RECT 46.865 61.605 47.330 61.935 ;
        RECT 45.650 61.545 45.850 61.575 ;
        RECT 45.970 61.325 46.140 61.395 ;
        RECT 45.270 61.155 46.140 61.325 ;
        RECT 45.630 61.065 46.140 61.155 ;
        RECT 44.180 60.600 44.485 60.730 ;
        RECT 44.930 60.620 45.460 60.985 ;
        RECT 43.800 60.005 44.065 60.465 ;
        RECT 44.235 60.175 44.485 60.600 ;
        RECT 45.630 60.450 45.800 61.065 ;
        RECT 44.695 60.280 45.800 60.450 ;
        RECT 45.970 60.005 46.140 60.805 ;
        RECT 46.310 60.505 46.480 61.575 ;
        RECT 46.650 60.675 46.840 61.395 ;
        RECT 47.010 60.645 47.330 61.605 ;
        RECT 47.500 61.645 47.670 62.105 ;
        RECT 47.945 62.025 48.155 62.555 ;
        RECT 48.415 61.815 48.745 62.340 ;
        RECT 48.915 61.945 49.085 62.555 ;
        RECT 49.255 61.900 49.585 62.335 ;
        RECT 49.255 61.815 49.635 61.900 ;
        RECT 48.545 61.645 48.745 61.815 ;
        RECT 49.410 61.775 49.635 61.815 ;
        RECT 47.500 61.315 48.375 61.645 ;
        RECT 48.545 61.315 49.295 61.645 ;
        RECT 46.310 60.175 46.560 60.505 ;
        RECT 47.500 60.475 47.670 61.315 ;
        RECT 48.545 61.110 48.735 61.315 ;
        RECT 49.465 61.195 49.635 61.775 ;
        RECT 49.805 61.785 51.475 62.555 ;
        RECT 49.805 61.265 50.555 61.785 ;
        RECT 51.920 61.745 52.165 62.350 ;
        RECT 52.385 62.020 52.895 62.555 ;
        RECT 49.420 61.145 49.635 61.195 ;
        RECT 47.840 60.735 48.735 61.110 ;
        RECT 49.245 61.065 49.635 61.145 ;
        RECT 50.725 61.095 51.475 61.615 ;
        RECT 46.785 60.305 47.670 60.475 ;
        RECT 47.850 60.005 48.165 60.505 ;
        RECT 48.395 60.175 48.735 60.735 ;
        RECT 48.905 60.005 49.075 61.015 ;
        RECT 49.245 60.220 49.575 61.065 ;
        RECT 49.805 60.005 51.475 61.095 ;
        RECT 51.645 61.575 52.875 61.745 ;
        RECT 51.645 60.765 51.985 61.575 ;
        RECT 52.155 61.010 52.905 61.200 ;
        RECT 51.645 60.355 52.160 60.765 ;
        RECT 52.395 60.005 52.565 60.765 ;
        RECT 52.735 60.345 52.905 61.010 ;
        RECT 53.075 61.025 53.265 62.385 ;
        RECT 53.435 61.875 53.710 62.385 ;
        RECT 53.900 62.020 54.430 62.385 ;
        RECT 54.855 62.155 55.185 62.555 ;
        RECT 54.255 61.985 54.430 62.020 ;
        RECT 53.435 61.705 53.715 61.875 ;
        RECT 53.435 61.225 53.710 61.705 ;
        RECT 53.915 61.025 54.085 61.825 ;
        RECT 53.075 60.855 54.085 61.025 ;
        RECT 54.255 61.815 55.185 61.985 ;
        RECT 55.355 61.815 55.610 62.385 ;
        RECT 54.255 60.685 54.425 61.815 ;
        RECT 55.015 61.645 55.185 61.815 ;
        RECT 53.300 60.515 54.425 60.685 ;
        RECT 54.595 61.315 54.790 61.645 ;
        RECT 55.015 61.315 55.270 61.645 ;
        RECT 54.595 60.345 54.765 61.315 ;
        RECT 55.440 61.145 55.610 61.815 ;
        RECT 55.785 61.785 57.455 62.555 ;
        RECT 57.675 61.900 58.005 62.335 ;
        RECT 58.175 61.945 58.345 62.555 ;
        RECT 57.625 61.815 58.005 61.900 ;
        RECT 58.515 61.815 58.845 62.340 ;
        RECT 59.105 62.025 59.315 62.555 ;
        RECT 59.590 62.105 60.375 62.275 ;
        RECT 60.545 62.105 60.950 62.275 ;
        RECT 55.785 61.265 56.535 61.785 ;
        RECT 57.625 61.775 57.850 61.815 ;
        RECT 52.735 60.175 54.765 60.345 ;
        RECT 54.935 60.005 55.105 61.145 ;
        RECT 55.275 60.175 55.610 61.145 ;
        RECT 56.705 61.095 57.455 61.615 ;
        RECT 55.785 60.005 57.455 61.095 ;
        RECT 57.625 61.195 57.795 61.775 ;
        RECT 58.515 61.645 58.715 61.815 ;
        RECT 59.590 61.645 59.760 62.105 ;
        RECT 57.965 61.315 58.715 61.645 ;
        RECT 58.885 61.315 59.760 61.645 ;
        RECT 57.625 61.145 57.840 61.195 ;
        RECT 57.625 61.065 58.015 61.145 ;
        RECT 57.685 60.220 58.015 61.065 ;
        RECT 58.525 61.110 58.715 61.315 ;
        RECT 58.185 60.005 58.355 61.015 ;
        RECT 58.525 60.735 59.420 61.110 ;
        RECT 58.525 60.175 58.865 60.735 ;
        RECT 59.095 60.005 59.410 60.505 ;
        RECT 59.590 60.475 59.760 61.315 ;
        RECT 59.930 61.605 60.395 61.935 ;
        RECT 60.780 61.875 60.950 62.105 ;
        RECT 61.130 62.055 61.500 62.555 ;
        RECT 61.820 62.105 62.495 62.275 ;
        RECT 62.690 62.105 63.025 62.275 ;
        RECT 59.930 60.645 60.250 61.605 ;
        RECT 60.780 61.575 61.610 61.875 ;
        RECT 60.420 60.675 60.610 61.395 ;
        RECT 60.780 60.505 60.950 61.575 ;
        RECT 61.410 61.545 61.610 61.575 ;
        RECT 61.120 61.325 61.290 61.395 ;
        RECT 61.820 61.325 61.990 62.105 ;
        RECT 62.855 61.965 63.025 62.105 ;
        RECT 63.195 62.095 63.445 62.555 ;
        RECT 61.120 61.155 61.990 61.325 ;
        RECT 62.160 61.685 62.685 61.905 ;
        RECT 62.855 61.835 63.080 61.965 ;
        RECT 61.120 61.065 61.630 61.155 ;
        RECT 59.590 60.305 60.475 60.475 ;
        RECT 60.700 60.175 60.950 60.505 ;
        RECT 61.120 60.005 61.290 60.805 ;
        RECT 61.460 60.450 61.630 61.065 ;
        RECT 62.160 60.985 62.330 61.685 ;
        RECT 61.800 60.620 62.330 60.985 ;
        RECT 62.500 60.920 62.740 61.515 ;
        RECT 62.910 60.730 63.080 61.835 ;
        RECT 63.250 60.975 63.530 61.925 ;
        RECT 62.775 60.600 63.080 60.730 ;
        RECT 61.460 60.280 62.565 60.450 ;
        RECT 62.775 60.175 63.025 60.600 ;
        RECT 63.195 60.005 63.460 60.465 ;
        RECT 63.700 60.175 63.885 62.295 ;
        RECT 64.055 62.175 64.385 62.555 ;
        RECT 64.555 62.005 64.725 62.295 ;
        RECT 64.060 61.835 64.725 62.005 ;
        RECT 64.060 60.845 64.290 61.835 ;
        RECT 64.985 61.830 65.275 62.555 ;
        RECT 65.445 62.055 65.705 62.385 ;
        RECT 65.875 62.195 66.205 62.555 ;
        RECT 66.460 62.175 67.760 62.385 ;
        RECT 65.445 62.045 65.675 62.055 ;
        RECT 64.460 61.015 64.810 61.665 ;
        RECT 64.060 60.675 64.725 60.845 ;
        RECT 64.055 60.005 64.385 60.505 ;
        RECT 64.555 60.175 64.725 60.675 ;
        RECT 64.985 60.005 65.275 61.170 ;
        RECT 65.445 60.855 65.615 62.045 ;
        RECT 66.460 62.025 66.630 62.175 ;
        RECT 65.875 61.900 66.630 62.025 ;
        RECT 65.785 61.855 66.630 61.900 ;
        RECT 65.785 61.735 66.055 61.855 ;
        RECT 65.785 61.160 65.955 61.735 ;
        RECT 66.185 61.295 66.595 61.600 ;
        RECT 66.885 61.565 67.095 61.965 ;
        RECT 66.765 61.355 67.095 61.565 ;
        RECT 67.340 61.565 67.560 61.965 ;
        RECT 68.035 61.790 68.490 62.555 ;
        RECT 68.665 61.755 69.360 62.385 ;
        RECT 69.565 61.755 69.875 62.555 ;
        RECT 70.055 61.905 70.385 62.380 ;
        RECT 70.555 62.075 70.725 62.555 ;
        RECT 70.895 61.905 71.225 62.380 ;
        RECT 71.395 62.075 71.565 62.555 ;
        RECT 71.735 61.905 72.065 62.380 ;
        RECT 72.235 62.075 72.405 62.555 ;
        RECT 72.575 61.905 72.905 62.380 ;
        RECT 73.075 62.075 73.245 62.555 ;
        RECT 73.415 61.905 73.745 62.380 ;
        RECT 73.915 62.075 74.085 62.555 ;
        RECT 74.255 62.380 74.505 62.385 ;
        RECT 74.255 61.905 74.585 62.380 ;
        RECT 74.755 62.075 74.925 62.555 ;
        RECT 75.175 62.380 75.345 62.385 ;
        RECT 75.095 61.905 75.425 62.380 ;
        RECT 75.595 62.075 75.765 62.555 ;
        RECT 76.015 62.380 76.185 62.385 ;
        RECT 75.935 61.905 76.265 62.380 ;
        RECT 76.435 62.075 76.605 62.555 ;
        RECT 76.775 61.905 77.105 62.380 ;
        RECT 77.275 62.075 77.445 62.555 ;
        RECT 77.615 61.905 77.945 62.380 ;
        RECT 78.115 62.075 78.285 62.555 ;
        RECT 78.455 61.905 78.785 62.380 ;
        RECT 78.955 62.075 79.125 62.555 ;
        RECT 79.295 61.905 79.625 62.380 ;
        RECT 79.795 62.075 79.965 62.555 ;
        RECT 80.135 61.905 80.465 62.380 ;
        RECT 80.635 62.075 80.805 62.555 ;
        RECT 67.340 61.355 67.815 61.565 ;
        RECT 68.005 61.365 68.495 61.565 ;
        RECT 68.685 61.315 69.020 61.565 ;
        RECT 65.785 61.125 65.985 61.160 ;
        RECT 67.315 61.125 68.490 61.185 ;
        RECT 69.190 61.155 69.360 61.755 ;
        RECT 70.055 61.735 71.565 61.905 ;
        RECT 71.735 61.735 74.085 61.905 ;
        RECT 74.255 61.735 80.915 61.905 ;
        RECT 81.085 61.755 81.395 62.555 ;
        RECT 81.600 61.755 82.295 62.385 ;
        RECT 83.390 61.815 83.645 62.385 ;
        RECT 83.815 62.155 84.145 62.555 ;
        RECT 84.570 62.020 85.100 62.385 ;
        RECT 85.290 62.215 85.565 62.385 ;
        RECT 85.285 62.045 85.565 62.215 ;
        RECT 84.570 61.985 84.745 62.020 ;
        RECT 83.815 61.815 84.745 61.985 ;
        RECT 69.530 61.315 69.865 61.585 ;
        RECT 71.395 61.565 71.565 61.735 ;
        RECT 73.910 61.565 74.085 61.735 ;
        RECT 70.050 61.365 71.225 61.565 ;
        RECT 71.395 61.365 73.705 61.565 ;
        RECT 73.910 61.365 80.470 61.565 ;
        RECT 71.395 61.195 71.565 61.365 ;
        RECT 73.910 61.195 74.085 61.365 ;
        RECT 80.640 61.195 80.915 61.735 ;
        RECT 81.095 61.315 81.430 61.585 ;
        RECT 65.785 61.015 68.490 61.125 ;
        RECT 65.845 60.955 67.645 61.015 ;
        RECT 67.315 60.925 67.645 60.955 ;
        RECT 65.445 60.175 65.705 60.855 ;
        RECT 65.875 60.005 66.125 60.785 ;
        RECT 66.375 60.755 67.210 60.765 ;
        RECT 67.800 60.755 67.985 60.845 ;
        RECT 66.375 60.555 67.985 60.755 ;
        RECT 66.375 60.175 66.625 60.555 ;
        RECT 67.755 60.515 67.985 60.555 ;
        RECT 68.235 60.395 68.490 61.015 ;
        RECT 66.795 60.005 67.150 60.385 ;
        RECT 68.155 60.175 68.490 60.395 ;
        RECT 68.665 60.005 68.925 61.145 ;
        RECT 69.095 60.175 69.425 61.155 ;
        RECT 69.595 60.005 69.875 61.145 ;
        RECT 70.055 61.025 71.565 61.195 ;
        RECT 71.735 61.025 74.085 61.195 ;
        RECT 74.255 61.025 80.915 61.195 ;
        RECT 81.600 61.155 81.770 61.755 ;
        RECT 81.940 61.315 82.275 61.565 ;
        RECT 70.055 60.175 70.385 61.025 ;
        RECT 70.555 60.005 70.725 60.855 ;
        RECT 70.895 60.175 71.225 61.025 ;
        RECT 71.395 60.005 71.565 60.855 ;
        RECT 71.735 60.175 72.065 61.025 ;
        RECT 72.235 60.005 72.405 60.805 ;
        RECT 72.575 60.175 72.905 61.025 ;
        RECT 73.075 60.005 73.245 60.805 ;
        RECT 73.415 60.175 73.745 61.025 ;
        RECT 73.915 60.005 74.085 60.805 ;
        RECT 74.255 60.175 74.585 61.025 ;
        RECT 74.755 60.005 74.925 60.805 ;
        RECT 75.095 60.175 75.425 61.025 ;
        RECT 75.595 60.005 75.765 60.805 ;
        RECT 75.935 60.175 76.265 61.025 ;
        RECT 76.435 60.005 76.605 60.805 ;
        RECT 76.775 60.175 77.105 61.025 ;
        RECT 77.275 60.005 77.445 60.805 ;
        RECT 77.615 60.175 77.945 61.025 ;
        RECT 78.115 60.005 78.285 60.805 ;
        RECT 78.455 60.175 78.785 61.025 ;
        RECT 78.955 60.005 79.125 60.805 ;
        RECT 79.295 60.175 79.625 61.025 ;
        RECT 79.795 60.005 79.965 60.805 ;
        RECT 80.135 60.175 80.465 61.025 ;
        RECT 80.635 60.005 80.805 60.805 ;
        RECT 81.085 60.005 81.365 61.145 ;
        RECT 81.535 60.175 81.865 61.155 ;
        RECT 83.390 61.145 83.560 61.815 ;
        RECT 83.815 61.645 83.985 61.815 ;
        RECT 83.730 61.315 83.985 61.645 ;
        RECT 84.210 61.315 84.405 61.645 ;
        RECT 82.035 60.005 82.295 61.145 ;
        RECT 83.390 60.175 83.725 61.145 ;
        RECT 83.895 60.005 84.065 61.145 ;
        RECT 84.235 60.345 84.405 61.315 ;
        RECT 84.575 60.685 84.745 61.815 ;
        RECT 84.915 61.025 85.085 61.825 ;
        RECT 85.290 61.225 85.565 62.045 ;
        RECT 85.735 61.025 85.925 62.385 ;
        RECT 86.105 62.020 86.615 62.555 ;
        RECT 86.835 61.745 87.080 62.350 ;
        RECT 87.525 61.880 87.785 62.385 ;
        RECT 87.965 62.175 88.295 62.555 ;
        RECT 88.475 62.005 88.645 62.385 ;
        RECT 86.125 61.575 87.355 61.745 ;
        RECT 84.915 60.855 85.925 61.025 ;
        RECT 86.095 61.010 86.845 61.200 ;
        RECT 84.575 60.515 85.700 60.685 ;
        RECT 86.095 60.345 86.265 61.010 ;
        RECT 87.015 60.765 87.355 61.575 ;
        RECT 84.235 60.175 86.265 60.345 ;
        RECT 86.435 60.005 86.605 60.765 ;
        RECT 86.840 60.355 87.355 60.765 ;
        RECT 87.525 61.080 87.695 61.880 ;
        RECT 87.980 61.835 88.645 62.005 ;
        RECT 88.995 62.005 89.165 62.385 ;
        RECT 89.380 62.175 89.710 62.555 ;
        RECT 88.995 61.835 89.710 62.005 ;
        RECT 87.980 61.580 88.150 61.835 ;
        RECT 87.865 61.250 88.150 61.580 ;
        RECT 88.385 61.285 88.715 61.655 ;
        RECT 88.905 61.285 89.260 61.655 ;
        RECT 89.540 61.645 89.710 61.835 ;
        RECT 89.880 61.810 90.135 62.385 ;
        RECT 89.540 61.315 89.795 61.645 ;
        RECT 87.980 61.105 88.150 61.250 ;
        RECT 89.540 61.105 89.710 61.315 ;
        RECT 87.525 60.175 87.795 61.080 ;
        RECT 87.980 60.935 88.645 61.105 ;
        RECT 87.965 60.005 88.295 60.765 ;
        RECT 88.475 60.175 88.645 60.935 ;
        RECT 88.995 60.935 89.710 61.105 ;
        RECT 89.965 61.080 90.135 61.810 ;
        RECT 90.310 61.715 90.570 62.555 ;
        RECT 90.745 61.805 91.955 62.555 ;
        RECT 88.995 60.175 89.165 60.935 ;
        RECT 89.380 60.005 89.710 60.765 ;
        RECT 89.880 60.175 90.135 61.080 ;
        RECT 90.310 60.005 90.570 61.155 ;
        RECT 90.745 61.095 91.265 61.635 ;
        RECT 91.435 61.265 91.955 61.805 ;
        RECT 90.745 60.005 91.955 61.095 ;
        RECT 13.380 59.835 92.040 60.005 ;
        RECT 13.465 58.745 14.675 59.835 ;
        RECT 13.465 58.035 13.985 58.575 ;
        RECT 14.155 58.205 14.675 58.745 ;
        RECT 14.850 58.685 15.110 59.835 ;
        RECT 15.285 58.760 15.540 59.665 ;
        RECT 15.710 59.075 16.040 59.835 ;
        RECT 16.255 58.905 16.425 59.665 ;
        RECT 16.775 59.165 16.945 59.665 ;
        RECT 17.115 59.335 17.445 59.835 ;
        RECT 16.775 58.995 17.440 59.165 ;
        RECT 13.465 57.285 14.675 58.035 ;
        RECT 14.850 57.285 15.110 58.125 ;
        RECT 15.285 58.030 15.455 58.760 ;
        RECT 15.710 58.735 16.425 58.905 ;
        RECT 15.710 58.525 15.880 58.735 ;
        RECT 15.625 58.195 15.880 58.525 ;
        RECT 15.285 57.455 15.540 58.030 ;
        RECT 15.710 58.005 15.880 58.195 ;
        RECT 16.160 58.185 16.515 58.555 ;
        RECT 16.690 58.175 17.040 58.825 ;
        RECT 17.210 58.005 17.440 58.995 ;
        RECT 15.710 57.835 16.425 58.005 ;
        RECT 15.710 57.285 16.040 57.665 ;
        RECT 16.255 57.455 16.425 57.835 ;
        RECT 16.775 57.835 17.440 58.005 ;
        RECT 16.775 57.545 16.945 57.835 ;
        RECT 17.115 57.285 17.445 57.665 ;
        RECT 17.615 57.545 17.800 59.665 ;
        RECT 18.040 59.375 18.305 59.835 ;
        RECT 18.475 59.240 18.725 59.665 ;
        RECT 18.935 59.390 20.040 59.560 ;
        RECT 18.420 59.110 18.725 59.240 ;
        RECT 17.970 57.915 18.250 58.865 ;
        RECT 18.420 58.005 18.590 59.110 ;
        RECT 18.760 58.325 19.000 58.920 ;
        RECT 19.170 58.855 19.700 59.220 ;
        RECT 19.170 58.155 19.340 58.855 ;
        RECT 19.870 58.775 20.040 59.390 ;
        RECT 20.210 59.035 20.380 59.835 ;
        RECT 20.550 59.335 20.800 59.665 ;
        RECT 21.025 59.365 21.910 59.535 ;
        RECT 19.870 58.685 20.380 58.775 ;
        RECT 18.420 57.875 18.645 58.005 ;
        RECT 18.815 57.935 19.340 58.155 ;
        RECT 19.510 58.515 20.380 58.685 ;
        RECT 18.055 57.285 18.305 57.745 ;
        RECT 18.475 57.735 18.645 57.875 ;
        RECT 19.510 57.735 19.680 58.515 ;
        RECT 20.210 58.445 20.380 58.515 ;
        RECT 19.890 58.265 20.090 58.295 ;
        RECT 20.550 58.265 20.720 59.335 ;
        RECT 20.890 58.445 21.080 59.165 ;
        RECT 19.890 57.965 20.720 58.265 ;
        RECT 21.250 58.235 21.570 59.195 ;
        RECT 18.475 57.565 18.810 57.735 ;
        RECT 19.005 57.565 19.680 57.735 ;
        RECT 20.000 57.285 20.370 57.785 ;
        RECT 20.550 57.735 20.720 57.965 ;
        RECT 21.105 57.905 21.570 58.235 ;
        RECT 21.740 58.525 21.910 59.365 ;
        RECT 22.090 59.335 22.405 59.835 ;
        RECT 22.635 59.105 22.975 59.665 ;
        RECT 22.080 58.730 22.975 59.105 ;
        RECT 23.145 58.825 23.315 59.835 ;
        RECT 22.785 58.525 22.975 58.730 ;
        RECT 23.485 58.775 23.815 59.620 ;
        RECT 23.485 58.695 23.875 58.775 ;
        RECT 24.045 58.745 25.715 59.835 ;
        RECT 23.660 58.645 23.875 58.695 ;
        RECT 21.740 58.195 22.615 58.525 ;
        RECT 22.785 58.195 23.535 58.525 ;
        RECT 21.740 57.735 21.910 58.195 ;
        RECT 22.785 58.025 22.985 58.195 ;
        RECT 23.705 58.065 23.875 58.645 ;
        RECT 23.650 58.025 23.875 58.065 ;
        RECT 20.550 57.565 20.955 57.735 ;
        RECT 21.125 57.565 21.910 57.735 ;
        RECT 22.185 57.285 22.395 57.815 ;
        RECT 22.655 57.500 22.985 58.025 ;
        RECT 23.495 57.940 23.875 58.025 ;
        RECT 24.045 58.055 24.795 58.575 ;
        RECT 24.965 58.225 25.715 58.745 ;
        RECT 26.345 58.670 26.635 59.835 ;
        RECT 26.990 58.865 27.380 59.040 ;
        RECT 27.865 59.035 28.195 59.835 ;
        RECT 28.365 59.045 28.900 59.665 ;
        RECT 26.990 58.695 28.415 58.865 ;
        RECT 23.155 57.285 23.325 57.895 ;
        RECT 23.495 57.505 23.825 57.940 ;
        RECT 24.045 57.285 25.715 58.055 ;
        RECT 26.345 57.285 26.635 58.010 ;
        RECT 26.865 57.965 27.220 58.525 ;
        RECT 27.390 57.795 27.560 58.695 ;
        RECT 27.730 57.965 27.995 58.525 ;
        RECT 28.245 58.195 28.415 58.695 ;
        RECT 28.585 58.025 28.900 59.045 ;
        RECT 29.770 58.865 30.100 59.665 ;
        RECT 30.270 59.035 30.600 59.835 ;
        RECT 30.900 58.865 31.230 59.665 ;
        RECT 31.875 59.035 32.125 59.835 ;
        RECT 29.770 58.695 32.205 58.865 ;
        RECT 32.395 58.695 32.565 59.835 ;
        RECT 32.735 58.695 33.075 59.665 ;
        RECT 33.245 58.745 34.915 59.835 ;
        RECT 35.175 59.165 35.345 59.665 ;
        RECT 35.515 59.335 35.845 59.835 ;
        RECT 35.175 58.995 35.840 59.165 ;
        RECT 29.565 58.275 29.915 58.525 ;
        RECT 30.100 58.065 30.270 58.695 ;
        RECT 30.440 58.275 30.770 58.475 ;
        RECT 30.940 58.275 31.270 58.475 ;
        RECT 31.440 58.275 31.860 58.475 ;
        RECT 32.035 58.445 32.205 58.695 ;
        RECT 32.035 58.275 32.730 58.445 ;
        RECT 26.970 57.285 27.210 57.795 ;
        RECT 27.390 57.465 27.670 57.795 ;
        RECT 27.900 57.285 28.115 57.795 ;
        RECT 28.285 57.455 28.900 58.025 ;
        RECT 29.770 57.455 30.270 58.065 ;
        RECT 30.900 57.935 32.125 58.105 ;
        RECT 32.900 58.085 33.075 58.695 ;
        RECT 30.900 57.455 31.230 57.935 ;
        RECT 31.400 57.285 31.625 57.745 ;
        RECT 31.795 57.455 32.125 57.935 ;
        RECT 32.315 57.285 32.565 58.085 ;
        RECT 32.735 57.455 33.075 58.085 ;
        RECT 33.245 58.055 33.995 58.575 ;
        RECT 34.165 58.225 34.915 58.745 ;
        RECT 35.090 58.175 35.440 58.825 ;
        RECT 33.245 57.285 34.915 58.055 ;
        RECT 35.610 58.005 35.840 58.995 ;
        RECT 35.175 57.835 35.840 58.005 ;
        RECT 35.175 57.545 35.345 57.835 ;
        RECT 35.515 57.285 35.845 57.665 ;
        RECT 36.015 57.545 36.200 59.665 ;
        RECT 36.440 59.375 36.705 59.835 ;
        RECT 36.875 59.240 37.125 59.665 ;
        RECT 37.335 59.390 38.440 59.560 ;
        RECT 36.820 59.110 37.125 59.240 ;
        RECT 36.370 57.915 36.650 58.865 ;
        RECT 36.820 58.005 36.990 59.110 ;
        RECT 37.160 58.325 37.400 58.920 ;
        RECT 37.570 58.855 38.100 59.220 ;
        RECT 37.570 58.155 37.740 58.855 ;
        RECT 38.270 58.775 38.440 59.390 ;
        RECT 38.610 59.035 38.780 59.835 ;
        RECT 38.950 59.335 39.200 59.665 ;
        RECT 39.425 59.365 40.310 59.535 ;
        RECT 38.270 58.685 38.780 58.775 ;
        RECT 36.820 57.875 37.045 58.005 ;
        RECT 37.215 57.935 37.740 58.155 ;
        RECT 37.910 58.515 38.780 58.685 ;
        RECT 36.455 57.285 36.705 57.745 ;
        RECT 36.875 57.735 37.045 57.875 ;
        RECT 37.910 57.735 38.080 58.515 ;
        RECT 38.610 58.445 38.780 58.515 ;
        RECT 38.290 58.265 38.490 58.295 ;
        RECT 38.950 58.265 39.120 59.335 ;
        RECT 39.290 58.445 39.480 59.165 ;
        RECT 38.290 57.965 39.120 58.265 ;
        RECT 39.650 58.235 39.970 59.195 ;
        RECT 36.875 57.565 37.210 57.735 ;
        RECT 37.405 57.565 38.080 57.735 ;
        RECT 38.400 57.285 38.770 57.785 ;
        RECT 38.950 57.735 39.120 57.965 ;
        RECT 39.505 57.905 39.970 58.235 ;
        RECT 40.140 58.525 40.310 59.365 ;
        RECT 40.490 59.335 40.805 59.835 ;
        RECT 41.035 59.105 41.375 59.665 ;
        RECT 40.480 58.730 41.375 59.105 ;
        RECT 41.545 58.825 41.715 59.835 ;
        RECT 41.185 58.525 41.375 58.730 ;
        RECT 41.885 58.775 42.215 59.620 ;
        RECT 41.885 58.695 42.275 58.775 ;
        RECT 42.060 58.645 42.275 58.695 ;
        RECT 40.140 58.195 41.015 58.525 ;
        RECT 41.185 58.195 41.935 58.525 ;
        RECT 40.140 57.735 40.310 58.195 ;
        RECT 41.185 58.025 41.385 58.195 ;
        RECT 42.105 58.065 42.275 58.645 ;
        RECT 42.050 58.025 42.275 58.065 ;
        RECT 38.950 57.565 39.355 57.735 ;
        RECT 39.525 57.565 40.310 57.735 ;
        RECT 40.585 57.285 40.795 57.815 ;
        RECT 41.055 57.500 41.385 58.025 ;
        RECT 41.895 57.940 42.275 58.025 ;
        RECT 42.450 58.695 42.785 59.665 ;
        RECT 42.955 58.695 43.125 59.835 ;
        RECT 43.295 59.495 45.325 59.665 ;
        RECT 42.450 58.025 42.620 58.695 ;
        RECT 43.295 58.525 43.465 59.495 ;
        RECT 42.790 58.195 43.045 58.525 ;
        RECT 43.270 58.195 43.465 58.525 ;
        RECT 43.635 59.155 44.760 59.325 ;
        RECT 42.875 58.025 43.045 58.195 ;
        RECT 43.635 58.025 43.805 59.155 ;
        RECT 41.555 57.285 41.725 57.895 ;
        RECT 41.895 57.505 42.225 57.940 ;
        RECT 42.450 57.455 42.705 58.025 ;
        RECT 42.875 57.855 43.805 58.025 ;
        RECT 43.975 58.815 44.985 58.985 ;
        RECT 43.975 58.015 44.145 58.815 ;
        RECT 43.630 57.820 43.805 57.855 ;
        RECT 42.875 57.285 43.205 57.685 ;
        RECT 43.630 57.455 44.160 57.820 ;
        RECT 44.350 57.795 44.625 58.615 ;
        RECT 44.345 57.625 44.625 57.795 ;
        RECT 44.350 57.455 44.625 57.625 ;
        RECT 44.795 57.455 44.985 58.815 ;
        RECT 45.155 58.830 45.325 59.495 ;
        RECT 45.495 59.075 45.665 59.835 ;
        RECT 45.900 59.075 46.415 59.485 ;
        RECT 45.155 58.640 45.905 58.830 ;
        RECT 46.075 58.265 46.415 59.075 ;
        RECT 45.185 58.095 46.415 58.265 ;
        RECT 47.045 59.075 47.560 59.485 ;
        RECT 47.795 59.075 47.965 59.835 ;
        RECT 48.135 59.495 50.165 59.665 ;
        RECT 47.045 58.265 47.385 59.075 ;
        RECT 48.135 58.830 48.305 59.495 ;
        RECT 48.700 59.155 49.825 59.325 ;
        RECT 47.555 58.640 48.305 58.830 ;
        RECT 48.475 58.815 49.485 58.985 ;
        RECT 47.045 58.095 48.275 58.265 ;
        RECT 45.165 57.285 45.675 57.820 ;
        RECT 45.895 57.490 46.140 58.095 ;
        RECT 47.320 57.490 47.565 58.095 ;
        RECT 47.785 57.285 48.295 57.820 ;
        RECT 48.475 57.455 48.665 58.815 ;
        RECT 48.835 58.475 49.110 58.615 ;
        RECT 48.835 58.305 49.115 58.475 ;
        RECT 48.835 57.455 49.110 58.305 ;
        RECT 49.315 58.015 49.485 58.815 ;
        RECT 49.655 58.025 49.825 59.155 ;
        RECT 49.995 58.525 50.165 59.495 ;
        RECT 50.335 58.695 50.505 59.835 ;
        RECT 50.675 58.695 51.010 59.665 ;
        RECT 49.995 58.195 50.190 58.525 ;
        RECT 50.415 58.195 50.670 58.525 ;
        RECT 50.415 58.025 50.585 58.195 ;
        RECT 50.840 58.025 51.010 58.695 ;
        RECT 52.105 58.670 52.395 59.835 ;
        RECT 52.565 58.745 56.075 59.835 ;
        RECT 49.655 57.855 50.585 58.025 ;
        RECT 49.655 57.820 49.830 57.855 ;
        RECT 49.300 57.455 49.830 57.820 ;
        RECT 50.255 57.285 50.585 57.685 ;
        RECT 50.755 57.455 51.010 58.025 ;
        RECT 52.565 58.055 54.215 58.575 ;
        RECT 54.385 58.225 56.075 58.745 ;
        RECT 56.250 58.695 56.585 59.665 ;
        RECT 56.755 58.695 56.925 59.835 ;
        RECT 57.095 59.495 59.125 59.665 ;
        RECT 52.105 57.285 52.395 58.010 ;
        RECT 52.565 57.285 56.075 58.055 ;
        RECT 56.250 58.025 56.420 58.695 ;
        RECT 57.095 58.525 57.265 59.495 ;
        RECT 56.590 58.195 56.845 58.525 ;
        RECT 57.070 58.195 57.265 58.525 ;
        RECT 57.435 59.155 58.560 59.325 ;
        RECT 56.675 58.025 56.845 58.195 ;
        RECT 57.435 58.025 57.605 59.155 ;
        RECT 56.250 57.455 56.505 58.025 ;
        RECT 56.675 57.855 57.605 58.025 ;
        RECT 57.775 58.815 58.785 58.985 ;
        RECT 57.775 58.015 57.945 58.815 ;
        RECT 57.430 57.820 57.605 57.855 ;
        RECT 56.675 57.285 57.005 57.685 ;
        RECT 57.430 57.455 57.960 57.820 ;
        RECT 58.150 57.795 58.425 58.615 ;
        RECT 58.145 57.625 58.425 57.795 ;
        RECT 58.150 57.455 58.425 57.625 ;
        RECT 58.595 57.455 58.785 58.815 ;
        RECT 58.955 58.830 59.125 59.495 ;
        RECT 59.295 59.075 59.465 59.835 ;
        RECT 59.700 59.075 60.215 59.485 ;
        RECT 60.385 59.400 65.730 59.835 ;
        RECT 58.955 58.640 59.705 58.830 ;
        RECT 59.875 58.265 60.215 59.075 ;
        RECT 58.985 58.095 60.215 58.265 ;
        RECT 58.965 57.285 59.475 57.820 ;
        RECT 59.695 57.490 59.940 58.095 ;
        RECT 61.970 57.830 62.310 58.660 ;
        RECT 63.790 58.150 64.140 59.400 ;
        RECT 65.905 58.985 66.165 59.665 ;
        RECT 66.335 59.055 66.585 59.835 ;
        RECT 66.835 59.285 67.085 59.665 ;
        RECT 67.255 59.455 67.610 59.835 ;
        RECT 68.615 59.445 68.950 59.665 ;
        RECT 68.215 59.285 68.445 59.325 ;
        RECT 66.835 59.085 68.445 59.285 ;
        RECT 66.835 59.075 67.670 59.085 ;
        RECT 68.260 58.995 68.445 59.085 ;
        RECT 60.385 57.285 65.730 57.830 ;
        RECT 65.905 57.795 66.075 58.985 ;
        RECT 67.775 58.885 68.105 58.915 ;
        RECT 66.305 58.825 68.105 58.885 ;
        RECT 68.695 58.825 68.950 59.445 ;
        RECT 66.245 58.715 68.950 58.825 ;
        RECT 66.245 58.680 66.445 58.715 ;
        RECT 66.245 58.105 66.415 58.680 ;
        RECT 67.775 58.655 68.950 58.715 ;
        RECT 69.125 58.695 69.405 59.835 ;
        RECT 69.575 58.685 69.905 59.665 ;
        RECT 70.075 58.695 70.335 59.835 ;
        RECT 70.515 58.775 70.845 59.625 ;
        RECT 69.640 58.645 69.815 58.685 ;
        RECT 66.645 58.240 67.055 58.545 ;
        RECT 67.225 58.275 67.555 58.485 ;
        RECT 66.245 57.985 66.515 58.105 ;
        RECT 66.245 57.940 67.090 57.985 ;
        RECT 66.335 57.815 67.090 57.940 ;
        RECT 67.345 57.875 67.555 58.275 ;
        RECT 67.800 58.275 68.275 58.485 ;
        RECT 68.465 58.275 68.955 58.475 ;
        RECT 67.800 57.875 68.020 58.275 ;
        RECT 69.135 58.255 69.470 58.525 ;
        RECT 69.640 58.085 69.810 58.645 ;
        RECT 69.980 58.275 70.315 58.525 ;
        RECT 65.905 57.785 66.135 57.795 ;
        RECT 65.905 57.455 66.165 57.785 ;
        RECT 66.920 57.665 67.090 57.815 ;
        RECT 66.335 57.285 66.665 57.645 ;
        RECT 66.920 57.455 68.220 57.665 ;
        RECT 68.495 57.285 68.950 58.050 ;
        RECT 69.125 57.285 69.435 58.085 ;
        RECT 69.640 57.455 70.335 58.085 ;
        RECT 70.515 58.010 70.705 58.775 ;
        RECT 71.015 58.695 71.265 59.835 ;
        RECT 71.455 59.195 71.705 59.615 ;
        RECT 71.935 59.365 72.265 59.835 ;
        RECT 72.495 59.195 72.745 59.615 ;
        RECT 71.455 59.025 72.745 59.195 ;
        RECT 72.925 59.195 73.255 59.625 ;
        RECT 72.925 59.025 73.380 59.195 ;
        RECT 71.445 58.525 71.660 58.855 ;
        RECT 70.875 58.195 71.185 58.525 ;
        RECT 71.355 58.195 71.660 58.525 ;
        RECT 71.835 58.195 72.120 58.855 ;
        RECT 72.315 58.195 72.580 58.855 ;
        RECT 72.795 58.195 73.040 58.855 ;
        RECT 71.015 58.025 71.185 58.195 ;
        RECT 73.210 58.025 73.380 59.025 ;
        RECT 73.880 58.825 74.180 59.665 ;
        RECT 74.375 58.995 74.625 59.835 ;
        RECT 75.215 59.245 76.020 59.665 ;
        RECT 74.795 59.075 76.360 59.245 ;
        RECT 74.795 58.825 74.965 59.075 ;
        RECT 73.880 58.655 74.965 58.825 ;
        RECT 73.725 58.195 74.055 58.485 ;
        RECT 74.225 58.025 74.395 58.655 ;
        RECT 75.135 58.525 75.455 58.905 ;
        RECT 75.645 58.815 76.020 58.905 ;
        RECT 75.625 58.645 76.020 58.815 ;
        RECT 76.190 58.825 76.360 59.075 ;
        RECT 76.530 58.995 76.860 59.835 ;
        RECT 77.030 59.075 77.695 59.665 ;
        RECT 76.190 58.655 77.110 58.825 ;
        RECT 74.565 58.275 74.895 58.485 ;
        RECT 75.075 58.275 75.455 58.525 ;
        RECT 75.645 58.485 76.020 58.645 ;
        RECT 76.940 58.485 77.110 58.655 ;
        RECT 75.645 58.275 76.130 58.485 ;
        RECT 76.320 58.275 76.770 58.485 ;
        RECT 76.940 58.275 77.275 58.485 ;
        RECT 77.445 58.105 77.695 59.075 ;
        RECT 77.865 58.670 78.155 59.835 ;
        RECT 78.330 59.445 78.665 59.665 ;
        RECT 79.670 59.455 80.025 59.835 ;
        RECT 78.330 58.825 78.585 59.445 ;
        RECT 78.835 59.285 79.065 59.325 ;
        RECT 80.195 59.285 80.445 59.665 ;
        RECT 78.835 59.085 80.445 59.285 ;
        RECT 78.835 58.995 79.020 59.085 ;
        RECT 79.610 59.075 80.445 59.085 ;
        RECT 80.695 59.055 80.945 59.835 ;
        RECT 81.115 58.985 81.375 59.665 ;
        RECT 82.095 59.165 82.265 59.665 ;
        RECT 82.435 59.335 82.765 59.835 ;
        RECT 82.095 58.995 82.760 59.165 ;
        RECT 79.175 58.885 79.505 58.915 ;
        RECT 79.175 58.825 80.975 58.885 ;
        RECT 78.330 58.715 81.035 58.825 ;
        RECT 78.330 58.655 79.505 58.715 ;
        RECT 80.835 58.680 81.035 58.715 ;
        RECT 78.325 58.275 78.815 58.475 ;
        RECT 79.005 58.275 79.480 58.485 ;
        RECT 70.515 57.500 70.845 58.010 ;
        RECT 71.015 57.855 73.380 58.025 ;
        RECT 71.015 57.285 71.345 57.685 ;
        RECT 72.395 57.515 72.725 57.855 ;
        RECT 73.885 57.845 74.395 58.025 ;
        RECT 74.800 57.935 76.500 58.105 ;
        RECT 74.800 57.845 75.185 57.935 ;
        RECT 72.895 57.285 73.225 57.685 ;
        RECT 73.885 57.455 74.215 57.845 ;
        RECT 74.385 57.505 75.570 57.675 ;
        RECT 75.830 57.285 76.000 57.755 ;
        RECT 76.170 57.470 76.500 57.935 ;
        RECT 76.670 57.285 76.840 58.105 ;
        RECT 77.010 57.465 77.695 58.105 ;
        RECT 77.865 57.285 78.155 58.010 ;
        RECT 78.330 57.285 78.785 58.050 ;
        RECT 79.260 57.875 79.480 58.275 ;
        RECT 79.725 58.275 80.055 58.485 ;
        RECT 79.725 57.875 79.935 58.275 ;
        RECT 80.225 58.240 80.635 58.545 ;
        RECT 80.865 58.105 81.035 58.680 ;
        RECT 80.765 57.985 81.035 58.105 ;
        RECT 80.190 57.940 81.035 57.985 ;
        RECT 80.190 57.815 80.945 57.940 ;
        RECT 80.190 57.665 80.360 57.815 ;
        RECT 81.205 57.785 81.375 58.985 ;
        RECT 82.010 58.175 82.360 58.825 ;
        RECT 82.530 58.005 82.760 58.995 ;
        RECT 79.060 57.455 80.360 57.665 ;
        RECT 80.615 57.285 80.945 57.645 ;
        RECT 81.115 57.455 81.375 57.785 ;
        RECT 82.095 57.835 82.760 58.005 ;
        RECT 82.095 57.545 82.265 57.835 ;
        RECT 82.435 57.285 82.765 57.665 ;
        RECT 82.935 57.545 83.120 59.665 ;
        RECT 83.360 59.375 83.625 59.835 ;
        RECT 83.795 59.240 84.045 59.665 ;
        RECT 84.255 59.390 85.360 59.560 ;
        RECT 83.740 59.110 84.045 59.240 ;
        RECT 83.290 57.915 83.570 58.865 ;
        RECT 83.740 58.005 83.910 59.110 ;
        RECT 84.080 58.325 84.320 58.920 ;
        RECT 84.490 58.855 85.020 59.220 ;
        RECT 84.490 58.155 84.660 58.855 ;
        RECT 85.190 58.775 85.360 59.390 ;
        RECT 85.530 59.035 85.700 59.835 ;
        RECT 85.870 59.335 86.120 59.665 ;
        RECT 86.345 59.365 87.230 59.535 ;
        RECT 85.190 58.685 85.700 58.775 ;
        RECT 83.740 57.875 83.965 58.005 ;
        RECT 84.135 57.935 84.660 58.155 ;
        RECT 84.830 58.515 85.700 58.685 ;
        RECT 83.375 57.285 83.625 57.745 ;
        RECT 83.795 57.735 83.965 57.875 ;
        RECT 84.830 57.735 85.000 58.515 ;
        RECT 85.530 58.445 85.700 58.515 ;
        RECT 85.210 58.265 85.410 58.295 ;
        RECT 85.870 58.265 86.040 59.335 ;
        RECT 86.210 58.445 86.400 59.165 ;
        RECT 85.210 57.965 86.040 58.265 ;
        RECT 86.570 58.235 86.890 59.195 ;
        RECT 83.795 57.565 84.130 57.735 ;
        RECT 84.325 57.565 85.000 57.735 ;
        RECT 85.320 57.285 85.690 57.785 ;
        RECT 85.870 57.735 86.040 57.965 ;
        RECT 86.425 57.905 86.890 58.235 ;
        RECT 87.060 58.525 87.230 59.365 ;
        RECT 87.410 59.335 87.725 59.835 ;
        RECT 87.955 59.105 88.295 59.665 ;
        RECT 87.400 58.730 88.295 59.105 ;
        RECT 88.465 58.825 88.635 59.835 ;
        RECT 88.105 58.525 88.295 58.730 ;
        RECT 88.805 58.775 89.135 59.620 ;
        RECT 88.805 58.695 89.195 58.775 ;
        RECT 88.980 58.645 89.195 58.695 ;
        RECT 87.060 58.195 87.935 58.525 ;
        RECT 88.105 58.195 88.855 58.525 ;
        RECT 87.060 57.735 87.230 58.195 ;
        RECT 88.105 58.025 88.305 58.195 ;
        RECT 89.025 58.065 89.195 58.645 ;
        RECT 88.970 58.025 89.195 58.065 ;
        RECT 85.870 57.565 86.275 57.735 ;
        RECT 86.445 57.565 87.230 57.735 ;
        RECT 87.505 57.285 87.715 57.815 ;
        RECT 87.975 57.500 88.305 58.025 ;
        RECT 88.815 57.940 89.195 58.025 ;
        RECT 89.365 58.760 89.635 59.665 ;
        RECT 89.805 59.075 90.135 59.835 ;
        RECT 90.315 58.905 90.485 59.665 ;
        RECT 89.365 57.960 89.535 58.760 ;
        RECT 89.820 58.735 90.485 58.905 ;
        RECT 90.745 58.745 91.955 59.835 ;
        RECT 89.820 58.590 89.990 58.735 ;
        RECT 89.705 58.260 89.990 58.590 ;
        RECT 89.820 58.005 89.990 58.260 ;
        RECT 90.225 58.185 90.555 58.555 ;
        RECT 90.745 58.205 91.265 58.745 ;
        RECT 91.435 58.035 91.955 58.575 ;
        RECT 88.475 57.285 88.645 57.895 ;
        RECT 88.815 57.505 89.145 57.940 ;
        RECT 89.365 57.455 89.625 57.960 ;
        RECT 89.820 57.835 90.485 58.005 ;
        RECT 89.805 57.285 90.135 57.665 ;
        RECT 90.315 57.455 90.485 57.835 ;
        RECT 90.745 57.285 91.955 58.035 ;
        RECT 13.380 57.115 92.040 57.285 ;
        RECT 13.465 56.365 14.675 57.115 ;
        RECT 14.845 56.365 16.055 57.115 ;
        RECT 13.465 55.825 13.985 56.365 ;
        RECT 14.155 55.655 14.675 56.195 ;
        RECT 14.845 55.825 15.365 56.365 ;
        RECT 16.225 56.315 16.565 56.945 ;
        RECT 16.735 56.315 16.985 57.115 ;
        RECT 17.175 56.465 17.505 56.945 ;
        RECT 17.675 56.655 17.900 57.115 ;
        RECT 18.070 56.465 18.400 56.945 ;
        RECT 15.535 55.655 16.055 56.195 ;
        RECT 13.465 54.565 14.675 55.655 ;
        RECT 14.845 54.565 16.055 55.655 ;
        RECT 16.225 55.705 16.400 56.315 ;
        RECT 17.175 56.295 18.400 56.465 ;
        RECT 19.030 56.335 19.530 56.945 ;
        RECT 16.570 55.955 17.265 56.125 ;
        RECT 17.095 55.705 17.265 55.955 ;
        RECT 17.440 55.925 17.860 56.125 ;
        RECT 18.030 55.925 18.360 56.125 ;
        RECT 18.530 55.925 18.860 56.125 ;
        RECT 19.030 55.705 19.200 56.335 ;
        RECT 19.905 56.315 20.245 56.945 ;
        RECT 20.415 56.315 20.665 57.115 ;
        RECT 20.855 56.465 21.185 56.945 ;
        RECT 21.355 56.655 21.580 57.115 ;
        RECT 21.750 56.465 22.080 56.945 ;
        RECT 19.385 55.875 19.735 56.125 ;
        RECT 19.905 55.705 20.080 56.315 ;
        RECT 20.855 56.295 22.080 56.465 ;
        RECT 22.710 56.335 23.210 56.945 ;
        RECT 23.635 56.575 23.860 56.935 ;
        RECT 24.040 56.745 24.370 57.115 ;
        RECT 24.550 56.575 24.805 56.935 ;
        RECT 25.370 56.745 26.115 57.115 ;
        RECT 23.635 56.385 26.120 56.575 ;
        RECT 20.250 55.955 20.945 56.125 ;
        RECT 20.775 55.705 20.945 55.955 ;
        RECT 21.120 55.925 21.540 56.125 ;
        RECT 21.710 55.925 22.040 56.125 ;
        RECT 22.210 55.925 22.540 56.125 ;
        RECT 22.710 55.705 22.880 56.335 ;
        RECT 23.065 55.875 23.415 56.125 ;
        RECT 23.595 55.875 23.865 56.205 ;
        RECT 24.045 55.875 24.480 56.205 ;
        RECT 24.660 55.875 25.235 56.205 ;
        RECT 25.415 55.875 25.695 56.205 ;
        RECT 16.225 54.735 16.565 55.705 ;
        RECT 16.735 54.565 16.905 55.705 ;
        RECT 17.095 55.535 19.530 55.705 ;
        RECT 17.175 54.565 17.425 55.365 ;
        RECT 18.070 54.735 18.400 55.535 ;
        RECT 18.700 54.565 19.030 55.365 ;
        RECT 19.200 54.735 19.530 55.535 ;
        RECT 19.905 54.735 20.245 55.705 ;
        RECT 20.415 54.565 20.585 55.705 ;
        RECT 20.775 55.535 23.210 55.705 ;
        RECT 25.895 55.695 26.120 56.385 ;
        RECT 20.855 54.565 21.105 55.365 ;
        RECT 21.750 54.735 22.080 55.535 ;
        RECT 22.380 54.565 22.710 55.365 ;
        RECT 22.880 54.735 23.210 55.535 ;
        RECT 23.625 55.515 26.120 55.695 ;
        RECT 26.295 55.515 26.630 56.935 ;
        RECT 27.010 56.335 27.510 56.945 ;
        RECT 26.805 55.875 27.155 56.125 ;
        RECT 27.340 55.705 27.510 56.335 ;
        RECT 28.140 56.465 28.470 56.945 ;
        RECT 28.640 56.655 28.865 57.115 ;
        RECT 29.035 56.465 29.365 56.945 ;
        RECT 28.140 56.295 29.365 56.465 ;
        RECT 29.555 56.315 29.805 57.115 ;
        RECT 29.975 56.315 30.315 56.945 ;
        RECT 30.575 56.565 30.745 56.855 ;
        RECT 30.915 56.735 31.245 57.115 ;
        RECT 30.575 56.395 31.240 56.565 ;
        RECT 30.085 56.265 30.315 56.315 ;
        RECT 27.680 55.925 28.010 56.125 ;
        RECT 28.180 55.925 28.510 56.125 ;
        RECT 28.680 55.925 29.100 56.125 ;
        RECT 29.275 55.955 29.970 56.125 ;
        RECT 29.275 55.705 29.445 55.955 ;
        RECT 30.140 55.705 30.315 56.265 ;
        RECT 23.625 54.745 23.915 55.515 ;
        RECT 24.485 55.105 25.675 55.335 ;
        RECT 24.485 54.745 24.745 55.105 ;
        RECT 24.915 54.565 25.245 54.935 ;
        RECT 25.415 54.745 25.675 55.105 ;
        RECT 25.865 54.565 26.195 55.285 ;
        RECT 26.365 54.745 26.630 55.515 ;
        RECT 27.010 55.535 29.445 55.705 ;
        RECT 27.010 54.735 27.340 55.535 ;
        RECT 27.510 54.565 27.840 55.365 ;
        RECT 28.140 54.735 28.470 55.535 ;
        RECT 29.115 54.565 29.365 55.365 ;
        RECT 29.635 54.565 29.805 55.705 ;
        RECT 29.975 54.735 30.315 55.705 ;
        RECT 30.490 55.575 30.840 56.225 ;
        RECT 31.010 55.405 31.240 56.395 ;
        RECT 30.575 55.235 31.240 55.405 ;
        RECT 30.575 54.735 30.745 55.235 ;
        RECT 30.915 54.565 31.245 55.065 ;
        RECT 31.415 54.735 31.600 56.855 ;
        RECT 31.855 56.655 32.105 57.115 ;
        RECT 32.275 56.665 32.610 56.835 ;
        RECT 32.805 56.665 33.480 56.835 ;
        RECT 32.275 56.525 32.445 56.665 ;
        RECT 31.770 55.535 32.050 56.485 ;
        RECT 32.220 56.395 32.445 56.525 ;
        RECT 32.220 55.290 32.390 56.395 ;
        RECT 32.615 56.245 33.140 56.465 ;
        RECT 32.560 55.480 32.800 56.075 ;
        RECT 32.970 55.545 33.140 56.245 ;
        RECT 33.310 55.885 33.480 56.665 ;
        RECT 33.800 56.615 34.170 57.115 ;
        RECT 34.350 56.665 34.755 56.835 ;
        RECT 34.925 56.665 35.710 56.835 ;
        RECT 34.350 56.435 34.520 56.665 ;
        RECT 33.690 56.135 34.520 56.435 ;
        RECT 34.905 56.165 35.370 56.495 ;
        RECT 33.690 56.105 33.890 56.135 ;
        RECT 34.010 55.885 34.180 55.955 ;
        RECT 33.310 55.715 34.180 55.885 ;
        RECT 33.670 55.625 34.180 55.715 ;
        RECT 32.220 55.160 32.525 55.290 ;
        RECT 32.970 55.180 33.500 55.545 ;
        RECT 31.840 54.565 32.105 55.025 ;
        RECT 32.275 54.735 32.525 55.160 ;
        RECT 33.670 55.010 33.840 55.625 ;
        RECT 32.735 54.840 33.840 55.010 ;
        RECT 34.010 54.565 34.180 55.365 ;
        RECT 34.350 55.065 34.520 56.135 ;
        RECT 34.690 55.235 34.880 55.955 ;
        RECT 35.050 55.205 35.370 56.165 ;
        RECT 35.540 56.205 35.710 56.665 ;
        RECT 35.985 56.585 36.195 57.115 ;
        RECT 36.455 56.375 36.785 56.900 ;
        RECT 36.955 56.505 37.125 57.115 ;
        RECT 37.295 56.460 37.625 56.895 ;
        RECT 37.295 56.375 37.675 56.460 ;
        RECT 36.585 56.205 36.785 56.375 ;
        RECT 37.450 56.335 37.675 56.375 ;
        RECT 35.540 55.875 36.415 56.205 ;
        RECT 36.585 55.875 37.335 56.205 ;
        RECT 34.350 54.735 34.600 55.065 ;
        RECT 35.540 55.035 35.710 55.875 ;
        RECT 36.585 55.670 36.775 55.875 ;
        RECT 37.505 55.755 37.675 56.335 ;
        RECT 37.845 56.365 39.055 57.115 ;
        RECT 39.225 56.390 39.515 57.115 ;
        RECT 39.690 56.375 39.945 56.945 ;
        RECT 40.115 56.715 40.445 57.115 ;
        RECT 40.870 56.580 41.400 56.945 ;
        RECT 40.870 56.545 41.045 56.580 ;
        RECT 40.115 56.375 41.045 56.545 ;
        RECT 37.845 55.825 38.365 56.365 ;
        RECT 37.460 55.705 37.675 55.755 ;
        RECT 35.880 55.295 36.775 55.670 ;
        RECT 37.285 55.625 37.675 55.705 ;
        RECT 38.535 55.655 39.055 56.195 ;
        RECT 34.825 54.865 35.710 55.035 ;
        RECT 35.890 54.565 36.205 55.065 ;
        RECT 36.435 54.735 36.775 55.295 ;
        RECT 36.945 54.565 37.115 55.575 ;
        RECT 37.285 54.780 37.615 55.625 ;
        RECT 37.845 54.565 39.055 55.655 ;
        RECT 39.225 54.565 39.515 55.730 ;
        RECT 39.690 55.705 39.860 56.375 ;
        RECT 40.115 56.205 40.285 56.375 ;
        RECT 40.030 55.875 40.285 56.205 ;
        RECT 40.510 55.875 40.705 56.205 ;
        RECT 39.690 54.735 40.025 55.705 ;
        RECT 40.195 54.565 40.365 55.705 ;
        RECT 40.535 54.905 40.705 55.875 ;
        RECT 40.875 55.245 41.045 56.375 ;
        RECT 41.215 55.585 41.385 56.385 ;
        RECT 41.590 56.095 41.865 56.945 ;
        RECT 41.585 55.925 41.865 56.095 ;
        RECT 41.590 55.785 41.865 55.925 ;
        RECT 42.035 55.585 42.225 56.945 ;
        RECT 42.405 56.580 42.915 57.115 ;
        RECT 43.135 56.305 43.380 56.910 ;
        RECT 43.825 56.375 44.210 56.945 ;
        RECT 44.380 56.655 44.705 57.115 ;
        RECT 45.225 56.485 45.505 56.945 ;
        RECT 42.425 56.135 43.655 56.305 ;
        RECT 41.215 55.415 42.225 55.585 ;
        RECT 42.395 55.570 43.145 55.760 ;
        RECT 40.875 55.075 42.000 55.245 ;
        RECT 42.395 54.905 42.565 55.570 ;
        RECT 43.315 55.325 43.655 56.135 ;
        RECT 40.535 54.735 42.565 54.905 ;
        RECT 42.735 54.565 42.905 55.325 ;
        RECT 43.140 54.915 43.655 55.325 ;
        RECT 43.825 55.705 44.105 56.375 ;
        RECT 44.380 56.315 45.505 56.485 ;
        RECT 44.380 56.205 44.830 56.315 ;
        RECT 44.275 55.875 44.830 56.205 ;
        RECT 45.695 56.145 46.095 56.945 ;
        RECT 46.495 56.655 46.765 57.115 ;
        RECT 46.935 56.485 47.220 56.945 ;
        RECT 43.825 54.735 44.210 55.705 ;
        RECT 44.380 55.415 44.830 55.875 ;
        RECT 45.000 55.585 46.095 56.145 ;
        RECT 44.380 55.195 45.505 55.415 ;
        RECT 44.380 54.565 44.705 55.025 ;
        RECT 45.225 54.735 45.505 55.195 ;
        RECT 45.695 54.735 46.095 55.585 ;
        RECT 46.265 56.315 47.220 56.485 ;
        RECT 46.265 55.415 46.475 56.315 ;
        RECT 46.645 55.585 47.335 56.145 ;
        RECT 47.510 55.515 47.845 56.935 ;
        RECT 48.025 56.745 48.770 57.115 ;
        RECT 49.335 56.575 49.590 56.935 ;
        RECT 49.770 56.745 50.100 57.115 ;
        RECT 50.280 56.575 50.505 56.935 ;
        RECT 48.020 56.385 50.505 56.575 ;
        RECT 48.020 55.695 48.245 56.385 ;
        RECT 50.725 56.345 52.395 57.115 ;
        RECT 52.570 56.375 52.825 56.945 ;
        RECT 52.995 56.715 53.325 57.115 ;
        RECT 53.750 56.580 54.280 56.945 ;
        RECT 53.750 56.545 53.925 56.580 ;
        RECT 52.995 56.375 53.925 56.545 ;
        RECT 48.445 55.875 48.725 56.205 ;
        RECT 48.905 55.875 49.480 56.205 ;
        RECT 49.660 55.875 50.095 56.205 ;
        RECT 50.275 55.875 50.545 56.205 ;
        RECT 50.725 55.825 51.475 56.345 ;
        RECT 48.020 55.515 50.515 55.695 ;
        RECT 51.645 55.655 52.395 56.175 ;
        RECT 46.265 55.195 47.220 55.415 ;
        RECT 46.495 54.565 46.765 55.025 ;
        RECT 46.935 54.735 47.220 55.195 ;
        RECT 47.510 54.745 47.775 55.515 ;
        RECT 47.945 54.565 48.275 55.285 ;
        RECT 48.465 55.105 49.655 55.335 ;
        RECT 48.465 54.745 48.725 55.105 ;
        RECT 48.895 54.565 49.225 54.935 ;
        RECT 49.395 54.745 49.655 55.105 ;
        RECT 50.225 54.745 50.515 55.515 ;
        RECT 50.725 54.565 52.395 55.655 ;
        RECT 52.570 55.705 52.740 56.375 ;
        RECT 52.995 56.205 53.165 56.375 ;
        RECT 52.910 55.875 53.165 56.205 ;
        RECT 53.390 55.875 53.585 56.205 ;
        RECT 52.570 54.735 52.905 55.705 ;
        RECT 53.075 54.565 53.245 55.705 ;
        RECT 53.415 54.905 53.585 55.875 ;
        RECT 53.755 55.245 53.925 56.375 ;
        RECT 54.095 55.585 54.265 56.385 ;
        RECT 54.470 56.095 54.745 56.945 ;
        RECT 54.465 55.925 54.745 56.095 ;
        RECT 54.470 55.785 54.745 55.925 ;
        RECT 54.915 55.585 55.105 56.945 ;
        RECT 55.285 56.580 55.795 57.115 ;
        RECT 56.015 56.305 56.260 56.910 ;
        RECT 56.705 56.375 57.090 56.945 ;
        RECT 57.260 56.655 57.585 57.115 ;
        RECT 58.105 56.485 58.385 56.945 ;
        RECT 55.305 56.135 56.535 56.305 ;
        RECT 54.095 55.415 55.105 55.585 ;
        RECT 55.275 55.570 56.025 55.760 ;
        RECT 53.755 55.075 54.880 55.245 ;
        RECT 55.275 54.905 55.445 55.570 ;
        RECT 56.195 55.325 56.535 56.135 ;
        RECT 53.415 54.735 55.445 54.905 ;
        RECT 55.615 54.565 55.785 55.325 ;
        RECT 56.020 54.915 56.535 55.325 ;
        RECT 56.705 55.705 56.985 56.375 ;
        RECT 57.260 56.315 58.385 56.485 ;
        RECT 57.260 56.205 57.710 56.315 ;
        RECT 57.155 55.875 57.710 56.205 ;
        RECT 58.575 56.145 58.975 56.945 ;
        RECT 59.375 56.655 59.645 57.115 ;
        RECT 59.815 56.485 60.100 56.945 ;
        RECT 56.705 54.735 57.090 55.705 ;
        RECT 57.260 55.415 57.710 55.875 ;
        RECT 57.880 55.585 58.975 56.145 ;
        RECT 57.260 55.195 58.385 55.415 ;
        RECT 57.260 54.565 57.585 55.025 ;
        RECT 58.105 54.735 58.385 55.195 ;
        RECT 58.575 54.735 58.975 55.585 ;
        RECT 59.145 56.315 60.100 56.485 ;
        RECT 60.845 56.375 61.230 56.945 ;
        RECT 61.400 56.655 61.725 57.115 ;
        RECT 62.245 56.485 62.525 56.945 ;
        RECT 59.145 55.415 59.355 56.315 ;
        RECT 59.525 55.585 60.215 56.145 ;
        RECT 60.845 55.705 61.125 56.375 ;
        RECT 61.400 56.315 62.525 56.485 ;
        RECT 61.400 56.205 61.850 56.315 ;
        RECT 61.295 55.875 61.850 56.205 ;
        RECT 62.715 56.145 63.115 56.945 ;
        RECT 63.515 56.655 63.785 57.115 ;
        RECT 63.955 56.485 64.240 56.945 ;
        RECT 59.145 55.195 60.100 55.415 ;
        RECT 59.375 54.565 59.645 55.025 ;
        RECT 59.815 54.735 60.100 55.195 ;
        RECT 60.845 54.735 61.230 55.705 ;
        RECT 61.400 55.415 61.850 55.875 ;
        RECT 62.020 55.585 63.115 56.145 ;
        RECT 61.400 55.195 62.525 55.415 ;
        RECT 61.400 54.565 61.725 55.025 ;
        RECT 62.245 54.735 62.525 55.195 ;
        RECT 62.715 54.735 63.115 55.585 ;
        RECT 63.285 56.315 64.240 56.485 ;
        RECT 64.985 56.390 65.275 57.115 ;
        RECT 65.560 56.485 65.845 56.945 ;
        RECT 66.015 56.655 66.285 57.115 ;
        RECT 65.560 56.315 66.515 56.485 ;
        RECT 63.285 55.415 63.495 56.315 ;
        RECT 63.665 55.585 64.355 56.145 ;
        RECT 63.285 55.195 64.240 55.415 ;
        RECT 63.515 54.565 63.785 55.025 ;
        RECT 63.955 54.735 64.240 55.195 ;
        RECT 64.985 54.565 65.275 55.730 ;
        RECT 65.445 55.585 66.135 56.145 ;
        RECT 66.305 55.415 66.515 56.315 ;
        RECT 65.560 55.195 66.515 55.415 ;
        RECT 66.685 56.145 67.085 56.945 ;
        RECT 67.275 56.485 67.555 56.945 ;
        RECT 68.075 56.655 68.400 57.115 ;
        RECT 67.275 56.315 68.400 56.485 ;
        RECT 68.570 56.375 68.955 56.945 ;
        RECT 69.135 56.605 70.365 56.945 ;
        RECT 70.535 56.625 70.790 57.115 ;
        RECT 69.135 56.375 69.465 56.605 ;
        RECT 67.950 56.205 68.400 56.315 ;
        RECT 66.685 55.585 67.780 56.145 ;
        RECT 67.950 55.875 68.505 56.205 ;
        RECT 65.560 54.735 65.845 55.195 ;
        RECT 66.015 54.565 66.285 55.025 ;
        RECT 66.685 54.735 67.085 55.585 ;
        RECT 67.950 55.415 68.400 55.875 ;
        RECT 68.675 55.705 68.955 56.375 ;
        RECT 69.125 55.875 69.435 56.205 ;
        RECT 69.640 55.875 70.015 56.435 ;
        RECT 70.185 55.705 70.365 56.605 ;
        RECT 70.550 55.875 70.770 56.455 ;
        RECT 71.055 56.435 71.225 56.810 ;
        RECT 71.025 56.265 71.225 56.435 ;
        RECT 71.415 56.585 71.645 56.890 ;
        RECT 71.815 56.755 72.145 57.115 ;
        RECT 72.340 56.585 72.630 56.935 ;
        RECT 73.765 56.605 74.165 57.115 ;
        RECT 71.415 56.415 72.630 56.585 ;
        RECT 74.740 56.500 74.910 56.945 ;
        RECT 75.080 56.715 75.800 57.115 ;
        RECT 75.970 56.545 76.140 56.945 ;
        RECT 76.375 56.670 76.805 57.115 ;
        RECT 71.055 56.245 71.225 56.265 ;
        RECT 71.055 56.075 71.575 56.245 ;
        RECT 67.275 55.195 68.400 55.415 ;
        RECT 67.275 54.735 67.555 55.195 ;
        RECT 68.075 54.565 68.400 55.025 ;
        RECT 68.570 54.735 68.955 55.705 ;
        RECT 69.135 55.535 70.365 55.705 ;
        RECT 69.135 54.735 69.465 55.535 ;
        RECT 69.635 54.565 69.865 55.365 ;
        RECT 70.035 54.735 70.365 55.535 ;
        RECT 70.535 54.565 70.790 55.705 ;
        RECT 70.970 55.545 71.215 55.905 ;
        RECT 71.405 55.695 71.575 56.075 ;
        RECT 71.745 55.875 72.130 56.205 ;
        RECT 72.310 56.095 72.570 56.205 ;
        RECT 72.310 55.925 72.575 56.095 ;
        RECT 72.310 55.875 72.570 55.925 ;
        RECT 71.405 55.415 71.755 55.695 ;
        RECT 70.970 54.565 71.225 55.365 ;
        RECT 71.425 54.735 71.755 55.415 ;
        RECT 71.935 54.825 72.130 55.875 ;
        RECT 72.310 54.565 72.630 55.705 ;
        RECT 73.780 55.545 74.040 56.435 ;
        RECT 74.240 55.845 74.500 56.435 ;
        RECT 74.740 56.330 75.090 56.500 ;
        RECT 74.240 55.545 74.720 55.845 ;
        RECT 73.805 55.195 74.745 55.365 ;
        RECT 73.805 54.735 73.985 55.195 ;
        RECT 74.155 54.565 74.405 55.025 ;
        RECT 74.575 54.945 74.745 55.195 ;
        RECT 74.920 55.305 75.090 56.330 ;
        RECT 75.260 56.375 76.140 56.545 ;
        RECT 76.975 56.390 77.235 56.945 ;
        RECT 75.260 55.655 75.430 56.375 ;
        RECT 75.620 55.825 75.910 56.205 ;
        RECT 75.260 55.485 75.780 55.655 ;
        RECT 76.080 55.585 76.410 56.205 ;
        RECT 76.635 55.875 76.890 56.205 ;
        RECT 74.920 55.135 75.330 55.305 ;
        RECT 75.610 55.295 75.780 55.485 ;
        RECT 76.635 55.395 76.805 55.875 ;
        RECT 77.060 55.675 77.235 56.390 ;
        RECT 77.425 56.385 77.755 57.115 ;
        RECT 77.925 56.205 78.135 56.825 ;
        RECT 78.315 56.405 78.745 56.935 ;
        RECT 77.440 55.855 77.730 56.205 ;
        RECT 77.925 55.855 78.320 56.205 ;
        RECT 78.500 56.155 78.745 56.405 ;
        RECT 78.925 56.335 79.155 57.115 ;
        RECT 79.335 56.485 79.715 56.935 ;
        RECT 80.715 56.565 80.885 56.855 ;
        RECT 81.055 56.735 81.385 57.115 ;
        RECT 78.500 55.855 79.035 56.155 ;
        RECT 79.335 56.035 79.565 56.485 ;
        RECT 80.715 56.395 81.380 56.565 ;
        RECT 75.075 55.000 75.330 55.135 ;
        RECT 76.045 55.225 76.805 55.395 ;
        RECT 76.045 55.000 76.215 55.225 ;
        RECT 74.575 54.775 74.905 54.945 ;
        RECT 75.075 54.830 76.215 55.000 ;
        RECT 75.075 54.735 75.330 54.830 ;
        RECT 76.475 54.565 76.805 54.965 ;
        RECT 76.975 54.735 77.235 55.675 ;
        RECT 77.495 55.475 78.535 55.675 ;
        RECT 77.495 54.745 77.665 55.475 ;
        RECT 77.845 54.565 78.175 55.295 ;
        RECT 78.345 54.745 78.535 55.475 ;
        RECT 78.705 54.745 79.035 55.855 ;
        RECT 79.225 55.355 79.565 56.035 ;
        RECT 79.745 55.535 79.975 56.225 ;
        RECT 80.630 55.575 80.980 56.225 ;
        RECT 81.150 55.405 81.380 56.395 ;
        RECT 79.225 55.155 79.985 55.355 ;
        RECT 79.225 54.565 79.555 54.975 ;
        RECT 79.725 54.765 79.985 55.155 ;
        RECT 80.715 55.235 81.380 55.405 ;
        RECT 80.715 54.735 80.885 55.235 ;
        RECT 81.055 54.565 81.385 55.065 ;
        RECT 81.555 54.735 81.740 56.855 ;
        RECT 81.995 56.655 82.245 57.115 ;
        RECT 82.415 56.665 82.750 56.835 ;
        RECT 82.945 56.665 83.620 56.835 ;
        RECT 82.415 56.525 82.585 56.665 ;
        RECT 81.910 55.535 82.190 56.485 ;
        RECT 82.360 56.395 82.585 56.525 ;
        RECT 82.360 55.290 82.530 56.395 ;
        RECT 82.755 56.245 83.280 56.465 ;
        RECT 82.700 55.480 82.940 56.075 ;
        RECT 83.110 55.545 83.280 56.245 ;
        RECT 83.450 55.885 83.620 56.665 ;
        RECT 83.940 56.615 84.310 57.115 ;
        RECT 84.490 56.665 84.895 56.835 ;
        RECT 85.065 56.665 85.850 56.835 ;
        RECT 84.490 56.435 84.660 56.665 ;
        RECT 83.830 56.135 84.660 56.435 ;
        RECT 85.045 56.165 85.510 56.495 ;
        RECT 83.830 56.105 84.030 56.135 ;
        RECT 84.150 55.885 84.320 55.955 ;
        RECT 83.450 55.715 84.320 55.885 ;
        RECT 83.810 55.625 84.320 55.715 ;
        RECT 82.360 55.160 82.665 55.290 ;
        RECT 83.110 55.180 83.640 55.545 ;
        RECT 81.980 54.565 82.245 55.025 ;
        RECT 82.415 54.735 82.665 55.160 ;
        RECT 83.810 55.010 83.980 55.625 ;
        RECT 82.875 54.840 83.980 55.010 ;
        RECT 84.150 54.565 84.320 55.365 ;
        RECT 84.490 55.065 84.660 56.135 ;
        RECT 84.830 55.235 85.020 55.955 ;
        RECT 85.190 55.205 85.510 56.165 ;
        RECT 85.680 56.205 85.850 56.665 ;
        RECT 86.125 56.585 86.335 57.115 ;
        RECT 86.595 56.375 86.925 56.900 ;
        RECT 87.095 56.505 87.265 57.115 ;
        RECT 87.435 56.460 87.765 56.895 ;
        RECT 88.995 56.565 89.165 56.945 ;
        RECT 89.380 56.735 89.710 57.115 ;
        RECT 87.435 56.375 87.815 56.460 ;
        RECT 88.995 56.395 89.710 56.565 ;
        RECT 86.725 56.205 86.925 56.375 ;
        RECT 87.590 56.335 87.815 56.375 ;
        RECT 85.680 55.875 86.555 56.205 ;
        RECT 86.725 55.875 87.475 56.205 ;
        RECT 84.490 54.735 84.740 55.065 ;
        RECT 85.680 55.035 85.850 55.875 ;
        RECT 86.725 55.670 86.915 55.875 ;
        RECT 87.645 55.755 87.815 56.335 ;
        RECT 88.905 55.845 89.260 56.215 ;
        RECT 89.540 56.205 89.710 56.395 ;
        RECT 89.880 56.370 90.135 56.945 ;
        RECT 89.540 55.875 89.795 56.205 ;
        RECT 87.600 55.705 87.815 55.755 ;
        RECT 86.020 55.295 86.915 55.670 ;
        RECT 87.425 55.625 87.815 55.705 ;
        RECT 89.540 55.665 89.710 55.875 ;
        RECT 84.965 54.865 85.850 55.035 ;
        RECT 86.030 54.565 86.345 55.065 ;
        RECT 86.575 54.735 86.915 55.295 ;
        RECT 87.085 54.565 87.255 55.575 ;
        RECT 87.425 54.780 87.755 55.625 ;
        RECT 88.995 55.495 89.710 55.665 ;
        RECT 89.965 55.640 90.135 56.370 ;
        RECT 90.310 56.275 90.570 57.115 ;
        RECT 90.745 56.365 91.955 57.115 ;
        RECT 88.995 54.735 89.165 55.495 ;
        RECT 89.380 54.565 89.710 55.325 ;
        RECT 89.880 54.735 90.135 55.640 ;
        RECT 90.310 54.565 90.570 55.715 ;
        RECT 90.745 55.655 91.265 56.195 ;
        RECT 91.435 55.825 91.955 56.365 ;
        RECT 90.745 54.565 91.955 55.655 ;
        RECT 13.380 54.395 92.040 54.565 ;
        RECT 13.465 53.305 14.675 54.395 ;
        RECT 13.465 52.595 13.985 53.135 ;
        RECT 14.155 52.765 14.675 53.305 ;
        RECT 15.030 53.425 15.420 53.600 ;
        RECT 15.905 53.595 16.235 54.395 ;
        RECT 16.405 53.605 16.940 54.225 ;
        RECT 15.030 53.255 16.455 53.425 ;
        RECT 13.465 51.845 14.675 52.595 ;
        RECT 14.905 52.525 15.260 53.085 ;
        RECT 15.430 52.355 15.600 53.255 ;
        RECT 15.770 52.525 16.035 53.085 ;
        RECT 16.285 52.755 16.455 53.255 ;
        RECT 16.625 52.585 16.940 53.605 ;
        RECT 17.235 53.725 17.405 54.225 ;
        RECT 17.575 53.895 17.905 54.395 ;
        RECT 17.235 53.555 17.900 53.725 ;
        RECT 17.150 52.735 17.500 53.385 ;
        RECT 15.010 51.845 15.250 52.355 ;
        RECT 15.430 52.025 15.710 52.355 ;
        RECT 15.940 51.845 16.155 52.355 ;
        RECT 16.325 52.015 16.940 52.585 ;
        RECT 17.670 52.565 17.900 53.555 ;
        RECT 17.235 52.395 17.900 52.565 ;
        RECT 17.235 52.105 17.405 52.395 ;
        RECT 17.575 51.845 17.905 52.225 ;
        RECT 18.075 52.105 18.260 54.225 ;
        RECT 18.500 53.935 18.765 54.395 ;
        RECT 18.935 53.800 19.185 54.225 ;
        RECT 19.395 53.950 20.500 54.120 ;
        RECT 18.880 53.670 19.185 53.800 ;
        RECT 18.430 52.475 18.710 53.425 ;
        RECT 18.880 52.565 19.050 53.670 ;
        RECT 19.220 52.885 19.460 53.480 ;
        RECT 19.630 53.415 20.160 53.780 ;
        RECT 19.630 52.715 19.800 53.415 ;
        RECT 20.330 53.335 20.500 53.950 ;
        RECT 20.670 53.595 20.840 54.395 ;
        RECT 21.010 53.895 21.260 54.225 ;
        RECT 21.485 53.925 22.370 54.095 ;
        RECT 20.330 53.245 20.840 53.335 ;
        RECT 18.880 52.435 19.105 52.565 ;
        RECT 19.275 52.495 19.800 52.715 ;
        RECT 19.970 53.075 20.840 53.245 ;
        RECT 18.515 51.845 18.765 52.305 ;
        RECT 18.935 52.295 19.105 52.435 ;
        RECT 19.970 52.295 20.140 53.075 ;
        RECT 20.670 53.005 20.840 53.075 ;
        RECT 20.350 52.825 20.550 52.855 ;
        RECT 21.010 52.825 21.180 53.895 ;
        RECT 21.350 53.005 21.540 53.725 ;
        RECT 20.350 52.525 21.180 52.825 ;
        RECT 21.710 52.795 22.030 53.755 ;
        RECT 18.935 52.125 19.270 52.295 ;
        RECT 19.465 52.125 20.140 52.295 ;
        RECT 20.460 51.845 20.830 52.345 ;
        RECT 21.010 52.295 21.180 52.525 ;
        RECT 21.565 52.465 22.030 52.795 ;
        RECT 22.200 53.085 22.370 53.925 ;
        RECT 22.550 53.895 22.865 54.395 ;
        RECT 23.095 53.665 23.435 54.225 ;
        RECT 22.540 53.290 23.435 53.665 ;
        RECT 23.605 53.385 23.775 54.395 ;
        RECT 23.245 53.085 23.435 53.290 ;
        RECT 23.945 53.335 24.275 54.180 ;
        RECT 23.945 53.255 24.335 53.335 ;
        RECT 24.505 53.305 26.175 54.395 ;
        RECT 24.120 53.205 24.335 53.255 ;
        RECT 22.200 52.755 23.075 53.085 ;
        RECT 23.245 52.755 23.995 53.085 ;
        RECT 22.200 52.295 22.370 52.755 ;
        RECT 23.245 52.585 23.445 52.755 ;
        RECT 24.165 52.625 24.335 53.205 ;
        RECT 24.110 52.585 24.335 52.625 ;
        RECT 21.010 52.125 21.415 52.295 ;
        RECT 21.585 52.125 22.370 52.295 ;
        RECT 22.645 51.845 22.855 52.375 ;
        RECT 23.115 52.060 23.445 52.585 ;
        RECT 23.955 52.500 24.335 52.585 ;
        RECT 24.505 52.615 25.255 53.135 ;
        RECT 25.425 52.785 26.175 53.305 ;
        RECT 26.345 53.230 26.635 54.395 ;
        RECT 26.815 53.285 27.110 54.395 ;
        RECT 27.290 53.085 27.540 54.220 ;
        RECT 27.710 53.285 27.970 54.395 ;
        RECT 28.140 53.495 28.400 54.220 ;
        RECT 28.570 53.665 28.830 54.395 ;
        RECT 29.000 53.495 29.260 54.220 ;
        RECT 29.430 53.665 29.690 54.395 ;
        RECT 29.860 53.495 30.120 54.220 ;
        RECT 30.290 53.665 30.550 54.395 ;
        RECT 30.720 53.495 30.980 54.220 ;
        RECT 31.150 53.665 31.445 54.395 ;
        RECT 28.140 53.255 31.450 53.495 ;
        RECT 31.905 53.445 32.195 54.215 ;
        RECT 32.765 53.855 33.025 54.215 ;
        RECT 33.195 54.025 33.525 54.395 ;
        RECT 33.695 53.855 33.955 54.215 ;
        RECT 32.765 53.625 33.955 53.855 ;
        RECT 34.145 53.675 34.475 54.395 ;
        RECT 34.645 53.445 34.910 54.215 ;
        RECT 35.085 53.960 40.430 54.395 ;
        RECT 40.605 53.960 45.950 54.395 ;
        RECT 31.905 53.265 34.400 53.445 ;
        RECT 23.615 51.845 23.785 52.455 ;
        RECT 23.955 52.065 24.285 52.500 ;
        RECT 24.505 51.845 26.175 52.615 ;
        RECT 26.345 51.845 26.635 52.570 ;
        RECT 26.805 52.475 27.120 53.085 ;
        RECT 27.290 52.835 30.310 53.085 ;
        RECT 26.865 51.845 27.110 52.305 ;
        RECT 27.290 52.025 27.540 52.835 ;
        RECT 30.480 52.665 31.450 53.255 ;
        RECT 31.875 52.755 32.145 53.085 ;
        RECT 32.325 52.755 32.760 53.085 ;
        RECT 32.940 52.755 33.515 53.085 ;
        RECT 33.695 52.755 33.975 53.085 ;
        RECT 28.140 52.495 31.450 52.665 ;
        RECT 34.175 52.575 34.400 53.265 ;
        RECT 27.710 51.845 27.970 52.370 ;
        RECT 28.140 52.040 28.400 52.495 ;
        RECT 28.570 51.845 28.830 52.325 ;
        RECT 29.000 52.040 29.260 52.495 ;
        RECT 29.430 51.845 29.690 52.325 ;
        RECT 29.860 52.040 30.120 52.495 ;
        RECT 30.290 51.845 30.550 52.325 ;
        RECT 30.720 52.040 30.980 52.495 ;
        RECT 31.915 52.385 34.400 52.575 ;
        RECT 31.150 51.845 31.450 52.325 ;
        RECT 31.915 52.025 32.140 52.385 ;
        RECT 32.320 51.845 32.650 52.215 ;
        RECT 32.830 52.025 33.085 52.385 ;
        RECT 33.650 51.845 34.395 52.215 ;
        RECT 34.575 52.025 34.910 53.445 ;
        RECT 36.670 52.390 37.010 53.220 ;
        RECT 38.490 52.710 38.840 53.960 ;
        RECT 42.190 52.390 42.530 53.220 ;
        RECT 44.010 52.710 44.360 53.960 ;
        RECT 46.125 53.305 48.715 54.395 ;
        RECT 46.125 52.615 47.335 53.135 ;
        RECT 47.505 52.785 48.715 53.305 ;
        RECT 48.890 53.445 49.155 54.215 ;
        RECT 49.325 53.675 49.655 54.395 ;
        RECT 49.845 53.855 50.105 54.215 ;
        RECT 50.275 54.025 50.605 54.395 ;
        RECT 50.775 53.855 51.035 54.215 ;
        RECT 49.845 53.625 51.035 53.855 ;
        RECT 51.605 53.445 51.895 54.215 ;
        RECT 35.085 51.845 40.430 52.390 ;
        RECT 40.605 51.845 45.950 52.390 ;
        RECT 46.125 51.845 48.715 52.615 ;
        RECT 48.890 52.025 49.225 53.445 ;
        RECT 49.400 53.265 51.895 53.445 ;
        RECT 49.400 52.575 49.625 53.265 ;
        RECT 52.105 53.230 52.395 54.395 ;
        RECT 53.575 53.725 53.745 54.225 ;
        RECT 53.915 53.895 54.245 54.395 ;
        RECT 53.575 53.555 54.240 53.725 ;
        RECT 49.825 52.755 50.105 53.085 ;
        RECT 50.285 52.755 50.860 53.085 ;
        RECT 51.040 52.755 51.475 53.085 ;
        RECT 51.655 52.755 51.925 53.085 ;
        RECT 53.490 52.735 53.840 53.385 ;
        RECT 49.400 52.385 51.885 52.575 ;
        RECT 49.405 51.845 50.150 52.215 ;
        RECT 50.715 52.025 50.970 52.385 ;
        RECT 51.150 51.845 51.480 52.215 ;
        RECT 51.660 52.025 51.885 52.385 ;
        RECT 52.105 51.845 52.395 52.570 ;
        RECT 54.010 52.565 54.240 53.555 ;
        RECT 53.575 52.395 54.240 52.565 ;
        RECT 53.575 52.105 53.745 52.395 ;
        RECT 53.915 51.845 54.245 52.225 ;
        RECT 54.415 52.105 54.600 54.225 ;
        RECT 54.840 53.935 55.105 54.395 ;
        RECT 55.275 53.800 55.525 54.225 ;
        RECT 55.735 53.950 56.840 54.120 ;
        RECT 55.220 53.670 55.525 53.800 ;
        RECT 54.770 52.475 55.050 53.425 ;
        RECT 55.220 52.565 55.390 53.670 ;
        RECT 55.560 52.885 55.800 53.480 ;
        RECT 55.970 53.415 56.500 53.780 ;
        RECT 55.970 52.715 56.140 53.415 ;
        RECT 56.670 53.335 56.840 53.950 ;
        RECT 57.010 53.595 57.180 54.395 ;
        RECT 57.350 53.895 57.600 54.225 ;
        RECT 57.825 53.925 58.710 54.095 ;
        RECT 56.670 53.245 57.180 53.335 ;
        RECT 55.220 52.435 55.445 52.565 ;
        RECT 55.615 52.495 56.140 52.715 ;
        RECT 56.310 53.075 57.180 53.245 ;
        RECT 54.855 51.845 55.105 52.305 ;
        RECT 55.275 52.295 55.445 52.435 ;
        RECT 56.310 52.295 56.480 53.075 ;
        RECT 57.010 53.005 57.180 53.075 ;
        RECT 56.690 52.825 56.890 52.855 ;
        RECT 57.350 52.825 57.520 53.895 ;
        RECT 57.690 53.005 57.880 53.725 ;
        RECT 56.690 52.525 57.520 52.825 ;
        RECT 58.050 52.795 58.370 53.755 ;
        RECT 55.275 52.125 55.610 52.295 ;
        RECT 55.805 52.125 56.480 52.295 ;
        RECT 56.800 51.845 57.170 52.345 ;
        RECT 57.350 52.295 57.520 52.525 ;
        RECT 57.905 52.465 58.370 52.795 ;
        RECT 58.540 53.085 58.710 53.925 ;
        RECT 58.890 53.895 59.205 54.395 ;
        RECT 59.435 53.665 59.775 54.225 ;
        RECT 58.880 53.290 59.775 53.665 ;
        RECT 59.945 53.385 60.115 54.395 ;
        RECT 59.585 53.085 59.775 53.290 ;
        RECT 60.285 53.335 60.615 54.180 ;
        RECT 60.905 53.335 61.235 54.180 ;
        RECT 61.405 53.385 61.575 54.395 ;
        RECT 61.745 53.665 62.085 54.225 ;
        RECT 62.315 53.895 62.630 54.395 ;
        RECT 62.810 53.925 63.695 54.095 ;
        RECT 60.285 53.255 60.675 53.335 ;
        RECT 60.460 53.205 60.675 53.255 ;
        RECT 58.540 52.755 59.415 53.085 ;
        RECT 59.585 52.755 60.335 53.085 ;
        RECT 58.540 52.295 58.710 52.755 ;
        RECT 59.585 52.585 59.785 52.755 ;
        RECT 60.505 52.625 60.675 53.205 ;
        RECT 60.450 52.585 60.675 52.625 ;
        RECT 57.350 52.125 57.755 52.295 ;
        RECT 57.925 52.125 58.710 52.295 ;
        RECT 58.985 51.845 59.195 52.375 ;
        RECT 59.455 52.060 59.785 52.585 ;
        RECT 60.295 52.500 60.675 52.585 ;
        RECT 60.845 53.255 61.235 53.335 ;
        RECT 61.745 53.290 62.640 53.665 ;
        RECT 60.845 53.205 61.060 53.255 ;
        RECT 60.845 52.625 61.015 53.205 ;
        RECT 61.745 53.085 61.935 53.290 ;
        RECT 62.810 53.085 62.980 53.925 ;
        RECT 63.920 53.895 64.170 54.225 ;
        RECT 61.185 52.755 61.935 53.085 ;
        RECT 62.105 52.755 62.980 53.085 ;
        RECT 60.845 52.585 61.070 52.625 ;
        RECT 61.735 52.585 61.935 52.755 ;
        RECT 60.845 52.500 61.225 52.585 ;
        RECT 59.955 51.845 60.125 52.455 ;
        RECT 60.295 52.065 60.625 52.500 ;
        RECT 60.895 52.065 61.225 52.500 ;
        RECT 61.395 51.845 61.565 52.455 ;
        RECT 61.735 52.060 62.065 52.585 ;
        RECT 62.325 51.845 62.535 52.375 ;
        RECT 62.810 52.295 62.980 52.755 ;
        RECT 63.150 52.795 63.470 53.755 ;
        RECT 63.640 53.005 63.830 53.725 ;
        RECT 64.000 52.825 64.170 53.895 ;
        RECT 64.340 53.595 64.510 54.395 ;
        RECT 64.680 53.950 65.785 54.120 ;
        RECT 64.680 53.335 64.850 53.950 ;
        RECT 65.995 53.800 66.245 54.225 ;
        RECT 66.415 53.935 66.680 54.395 ;
        RECT 65.020 53.415 65.550 53.780 ;
        RECT 65.995 53.670 66.300 53.800 ;
        RECT 64.340 53.245 64.850 53.335 ;
        RECT 64.340 53.075 65.210 53.245 ;
        RECT 64.340 53.005 64.510 53.075 ;
        RECT 64.630 52.825 64.830 52.855 ;
        RECT 63.150 52.465 63.615 52.795 ;
        RECT 64.000 52.525 64.830 52.825 ;
        RECT 64.000 52.295 64.170 52.525 ;
        RECT 62.810 52.125 63.595 52.295 ;
        RECT 63.765 52.125 64.170 52.295 ;
        RECT 64.350 51.845 64.720 52.345 ;
        RECT 65.040 52.295 65.210 53.075 ;
        RECT 65.380 52.715 65.550 53.415 ;
        RECT 65.720 52.885 65.960 53.480 ;
        RECT 65.380 52.495 65.905 52.715 ;
        RECT 66.130 52.565 66.300 53.670 ;
        RECT 66.075 52.435 66.300 52.565 ;
        RECT 66.470 52.475 66.750 53.425 ;
        RECT 66.075 52.295 66.245 52.435 ;
        RECT 65.040 52.125 65.715 52.295 ;
        RECT 65.910 52.125 66.245 52.295 ;
        RECT 66.415 51.845 66.665 52.305 ;
        RECT 66.920 52.105 67.105 54.225 ;
        RECT 67.275 53.895 67.605 54.395 ;
        RECT 67.775 53.725 67.945 54.225 ;
        RECT 67.280 53.555 67.945 53.725 ;
        RECT 67.280 52.565 67.510 53.555 ;
        RECT 67.680 52.735 68.030 53.385 ;
        RECT 68.265 53.335 68.595 54.180 ;
        RECT 68.765 53.385 68.935 54.395 ;
        RECT 69.105 53.665 69.445 54.225 ;
        RECT 69.675 53.895 69.990 54.395 ;
        RECT 70.170 53.925 71.055 54.095 ;
        RECT 68.205 53.255 68.595 53.335 ;
        RECT 69.105 53.290 70.000 53.665 ;
        RECT 68.205 53.205 68.420 53.255 ;
        RECT 68.205 52.625 68.375 53.205 ;
        RECT 69.105 53.085 69.295 53.290 ;
        RECT 70.170 53.085 70.340 53.925 ;
        RECT 71.280 53.895 71.530 54.225 ;
        RECT 68.545 52.755 69.295 53.085 ;
        RECT 69.465 52.755 70.340 53.085 ;
        RECT 68.205 52.585 68.430 52.625 ;
        RECT 69.095 52.585 69.295 52.755 ;
        RECT 67.280 52.395 67.945 52.565 ;
        RECT 68.205 52.500 68.585 52.585 ;
        RECT 67.275 51.845 67.605 52.225 ;
        RECT 67.775 52.105 67.945 52.395 ;
        RECT 68.255 52.065 68.585 52.500 ;
        RECT 68.755 51.845 68.925 52.455 ;
        RECT 69.095 52.060 69.425 52.585 ;
        RECT 69.685 51.845 69.895 52.375 ;
        RECT 70.170 52.295 70.340 52.755 ;
        RECT 70.510 52.795 70.830 53.755 ;
        RECT 71.000 53.005 71.190 53.725 ;
        RECT 71.360 52.825 71.530 53.895 ;
        RECT 71.700 53.595 71.870 54.395 ;
        RECT 72.040 53.950 73.145 54.120 ;
        RECT 72.040 53.335 72.210 53.950 ;
        RECT 73.355 53.800 73.605 54.225 ;
        RECT 73.775 53.935 74.040 54.395 ;
        RECT 72.380 53.415 72.910 53.780 ;
        RECT 73.355 53.670 73.660 53.800 ;
        RECT 71.700 53.245 72.210 53.335 ;
        RECT 71.700 53.075 72.570 53.245 ;
        RECT 71.700 53.005 71.870 53.075 ;
        RECT 71.990 52.825 72.190 52.855 ;
        RECT 70.510 52.465 70.975 52.795 ;
        RECT 71.360 52.525 72.190 52.825 ;
        RECT 71.360 52.295 71.530 52.525 ;
        RECT 70.170 52.125 70.955 52.295 ;
        RECT 71.125 52.125 71.530 52.295 ;
        RECT 71.710 51.845 72.080 52.345 ;
        RECT 72.400 52.295 72.570 53.075 ;
        RECT 72.740 52.715 72.910 53.415 ;
        RECT 73.080 52.885 73.320 53.480 ;
        RECT 72.740 52.495 73.265 52.715 ;
        RECT 73.490 52.565 73.660 53.670 ;
        RECT 73.435 52.435 73.660 52.565 ;
        RECT 73.830 52.475 74.110 53.425 ;
        RECT 73.435 52.295 73.605 52.435 ;
        RECT 72.400 52.125 73.075 52.295 ;
        RECT 73.270 52.125 73.605 52.295 ;
        RECT 73.775 51.845 74.025 52.305 ;
        RECT 74.280 52.105 74.465 54.225 ;
        RECT 74.635 53.895 74.965 54.395 ;
        RECT 75.135 53.725 75.305 54.225 ;
        RECT 74.640 53.555 75.305 53.725 ;
        RECT 74.640 52.565 74.870 53.555 ;
        RECT 75.040 52.735 75.390 53.385 ;
        RECT 75.565 53.255 75.845 54.395 ;
        RECT 76.015 53.245 76.345 54.225 ;
        RECT 76.515 53.255 76.775 54.395 ;
        RECT 75.575 52.815 75.910 53.085 ;
        RECT 76.080 52.645 76.250 53.245 ;
        RECT 77.865 53.230 78.155 54.395 ;
        RECT 78.325 53.255 78.710 54.225 ;
        RECT 78.880 53.935 79.205 54.395 ;
        RECT 79.725 53.765 80.005 54.225 ;
        RECT 78.880 53.545 80.005 53.765 ;
        RECT 76.420 52.835 76.755 53.085 ;
        RECT 74.640 52.395 75.305 52.565 ;
        RECT 74.635 51.845 74.965 52.225 ;
        RECT 75.135 52.105 75.305 52.395 ;
        RECT 75.565 51.845 75.875 52.645 ;
        RECT 76.080 52.015 76.775 52.645 ;
        RECT 78.325 52.585 78.605 53.255 ;
        RECT 78.880 53.085 79.330 53.545 ;
        RECT 80.195 53.375 80.595 54.225 ;
        RECT 80.995 53.935 81.265 54.395 ;
        RECT 81.435 53.765 81.720 54.225 ;
        RECT 78.775 52.755 79.330 53.085 ;
        RECT 79.500 52.815 80.595 53.375 ;
        RECT 78.880 52.645 79.330 52.755 ;
        RECT 77.865 51.845 78.155 52.570 ;
        RECT 78.325 52.015 78.710 52.585 ;
        RECT 78.880 52.475 80.005 52.645 ;
        RECT 78.880 51.845 79.205 52.305 ;
        RECT 79.725 52.015 80.005 52.475 ;
        RECT 80.195 52.015 80.595 52.815 ;
        RECT 80.765 53.545 81.720 53.765 ;
        RECT 80.765 52.645 80.975 53.545 ;
        RECT 81.145 52.815 81.835 53.375 ;
        RECT 82.470 53.255 82.805 54.225 ;
        RECT 82.975 53.255 83.145 54.395 ;
        RECT 83.315 54.055 85.345 54.225 ;
        RECT 80.765 52.475 81.720 52.645 ;
        RECT 80.995 51.845 81.265 52.305 ;
        RECT 81.435 52.015 81.720 52.475 ;
        RECT 82.470 52.585 82.640 53.255 ;
        RECT 83.315 53.085 83.485 54.055 ;
        RECT 82.810 52.755 83.065 53.085 ;
        RECT 83.290 52.755 83.485 53.085 ;
        RECT 83.655 53.715 84.780 53.885 ;
        RECT 82.895 52.585 83.065 52.755 ;
        RECT 83.655 52.585 83.825 53.715 ;
        RECT 82.470 52.015 82.725 52.585 ;
        RECT 82.895 52.415 83.825 52.585 ;
        RECT 83.995 53.375 85.005 53.545 ;
        RECT 83.995 52.575 84.165 53.375 ;
        RECT 83.650 52.380 83.825 52.415 ;
        RECT 82.895 51.845 83.225 52.245 ;
        RECT 83.650 52.015 84.180 52.380 ;
        RECT 84.370 52.355 84.645 53.175 ;
        RECT 84.365 52.185 84.645 52.355 ;
        RECT 84.370 52.015 84.645 52.185 ;
        RECT 84.815 52.015 85.005 53.375 ;
        RECT 85.175 53.390 85.345 54.055 ;
        RECT 85.515 53.635 85.685 54.395 ;
        RECT 85.920 53.635 86.435 54.045 ;
        RECT 85.175 53.200 85.925 53.390 ;
        RECT 86.095 52.825 86.435 53.635 ;
        RECT 85.205 52.655 86.435 52.825 ;
        RECT 86.605 53.255 86.990 54.225 ;
        RECT 87.160 53.935 87.485 54.395 ;
        RECT 88.005 53.765 88.285 54.225 ;
        RECT 87.160 53.545 88.285 53.765 ;
        RECT 85.185 51.845 85.695 52.380 ;
        RECT 85.915 52.050 86.160 52.655 ;
        RECT 86.605 52.585 86.885 53.255 ;
        RECT 87.160 53.085 87.610 53.545 ;
        RECT 88.475 53.375 88.875 54.225 ;
        RECT 89.275 53.935 89.545 54.395 ;
        RECT 89.715 53.765 90.000 54.225 ;
        RECT 87.055 52.755 87.610 53.085 ;
        RECT 87.780 52.815 88.875 53.375 ;
        RECT 87.160 52.645 87.610 52.755 ;
        RECT 86.605 52.015 86.990 52.585 ;
        RECT 87.160 52.475 88.285 52.645 ;
        RECT 87.160 51.845 87.485 52.305 ;
        RECT 88.005 52.015 88.285 52.475 ;
        RECT 88.475 52.015 88.875 52.815 ;
        RECT 89.045 53.545 90.000 53.765 ;
        RECT 89.045 52.645 89.255 53.545 ;
        RECT 89.425 52.815 90.115 53.375 ;
        RECT 90.745 53.305 91.955 54.395 ;
        RECT 90.745 52.765 91.265 53.305 ;
        RECT 89.045 52.475 90.000 52.645 ;
        RECT 91.435 52.595 91.955 53.135 ;
        RECT 89.275 51.845 89.545 52.305 ;
        RECT 89.715 52.015 90.000 52.475 ;
        RECT 90.745 51.845 91.955 52.595 ;
        RECT 13.380 51.675 92.040 51.845 ;
        RECT 13.465 50.925 14.675 51.675 ;
        RECT 13.465 50.385 13.985 50.925 ;
        RECT 14.850 50.835 15.110 51.675 ;
        RECT 15.285 50.930 15.540 51.505 ;
        RECT 15.710 51.295 16.040 51.675 ;
        RECT 16.255 51.125 16.425 51.505 ;
        RECT 15.710 50.955 16.425 51.125 ;
        RECT 14.155 50.215 14.675 50.755 ;
        RECT 13.465 49.125 14.675 50.215 ;
        RECT 14.850 49.125 15.110 50.275 ;
        RECT 15.285 50.200 15.455 50.930 ;
        RECT 15.710 50.765 15.880 50.955 ;
        RECT 16.690 50.835 16.950 51.675 ;
        RECT 17.125 50.930 17.380 51.505 ;
        RECT 17.550 51.295 17.880 51.675 ;
        RECT 18.095 51.125 18.265 51.505 ;
        RECT 18.525 51.130 23.870 51.675 ;
        RECT 24.670 51.165 24.910 51.675 ;
        RECT 25.090 51.165 25.370 51.495 ;
        RECT 25.600 51.165 25.815 51.675 ;
        RECT 17.550 50.955 18.265 51.125 ;
        RECT 15.625 50.435 15.880 50.765 ;
        RECT 15.710 50.225 15.880 50.435 ;
        RECT 16.160 50.405 16.515 50.775 ;
        RECT 15.285 49.295 15.540 50.200 ;
        RECT 15.710 50.055 16.425 50.225 ;
        RECT 15.710 49.125 16.040 49.885 ;
        RECT 16.255 49.295 16.425 50.055 ;
        RECT 16.690 49.125 16.950 50.275 ;
        RECT 17.125 50.200 17.295 50.930 ;
        RECT 17.550 50.765 17.720 50.955 ;
        RECT 17.465 50.435 17.720 50.765 ;
        RECT 17.550 50.225 17.720 50.435 ;
        RECT 18.000 50.405 18.355 50.775 ;
        RECT 20.110 50.300 20.450 51.130 ;
        RECT 17.125 49.295 17.380 50.200 ;
        RECT 17.550 50.055 18.265 50.225 ;
        RECT 17.550 49.125 17.880 49.885 ;
        RECT 18.095 49.295 18.265 50.055 ;
        RECT 21.930 49.560 22.280 50.810 ;
        RECT 24.565 50.435 24.920 50.995 ;
        RECT 25.090 50.265 25.260 51.165 ;
        RECT 25.430 50.435 25.695 50.995 ;
        RECT 25.985 50.935 26.600 51.505 ;
        RECT 27.050 51.195 27.350 51.675 ;
        RECT 27.520 51.025 27.780 51.480 ;
        RECT 27.950 51.195 28.210 51.675 ;
        RECT 28.380 51.025 28.640 51.480 ;
        RECT 28.810 51.195 29.070 51.675 ;
        RECT 29.240 51.025 29.500 51.480 ;
        RECT 29.670 51.195 29.930 51.675 ;
        RECT 30.100 51.025 30.360 51.480 ;
        RECT 30.530 51.150 30.790 51.675 ;
        RECT 25.945 50.265 26.115 50.765 ;
        RECT 24.690 50.095 26.115 50.265 ;
        RECT 24.690 49.920 25.080 50.095 ;
        RECT 18.525 49.125 23.870 49.560 ;
        RECT 25.565 49.125 25.895 49.925 ;
        RECT 26.285 49.915 26.600 50.935 ;
        RECT 27.050 50.855 30.360 51.025 ;
        RECT 27.050 50.265 28.020 50.855 ;
        RECT 30.960 50.685 31.210 51.495 ;
        RECT 31.390 51.215 31.635 51.675 ;
        RECT 32.030 51.165 32.270 51.675 ;
        RECT 32.450 51.165 32.730 51.495 ;
        RECT 32.960 51.165 33.175 51.675 ;
        RECT 28.190 50.435 31.210 50.685 ;
        RECT 31.380 50.435 31.695 51.045 ;
        RECT 31.925 50.435 32.280 50.995 ;
        RECT 27.050 50.025 30.360 50.265 ;
        RECT 26.065 49.295 26.600 49.915 ;
        RECT 27.055 49.125 27.350 49.855 ;
        RECT 27.520 49.300 27.780 50.025 ;
        RECT 27.950 49.125 28.210 49.855 ;
        RECT 28.380 49.300 28.640 50.025 ;
        RECT 28.810 49.125 29.070 49.855 ;
        RECT 29.240 49.300 29.500 50.025 ;
        RECT 29.670 49.125 29.930 49.855 ;
        RECT 30.100 49.300 30.360 50.025 ;
        RECT 30.530 49.125 30.790 50.235 ;
        RECT 30.960 49.300 31.210 50.435 ;
        RECT 32.450 50.265 32.620 51.165 ;
        RECT 32.790 50.435 33.055 50.995 ;
        RECT 33.345 50.935 33.960 51.505 ;
        RECT 33.305 50.265 33.475 50.765 ;
        RECT 31.390 49.125 31.685 50.235 ;
        RECT 32.050 50.095 33.475 50.265 ;
        RECT 32.050 49.920 32.440 50.095 ;
        RECT 32.925 49.125 33.255 49.925 ;
        RECT 33.645 49.915 33.960 50.935 ;
        RECT 34.165 50.905 35.835 51.675 ;
        RECT 36.525 51.205 36.825 51.675 ;
        RECT 36.995 51.035 37.250 51.480 ;
        RECT 37.420 51.205 37.680 51.675 ;
        RECT 37.850 51.035 38.110 51.480 ;
        RECT 38.280 51.205 38.575 51.675 ;
        RECT 34.165 50.385 34.915 50.905 ;
        RECT 36.005 50.865 39.035 51.035 ;
        RECT 39.225 50.950 39.515 51.675 ;
        RECT 35.085 50.215 35.835 50.735 ;
        RECT 33.425 49.295 33.960 49.915 ;
        RECT 34.165 49.125 35.835 50.215 ;
        RECT 36.005 50.300 36.305 50.865 ;
        RECT 36.480 50.470 38.695 50.695 ;
        RECT 38.865 50.300 39.035 50.865 ;
        RECT 36.005 50.130 39.035 50.300 ;
        RECT 36.005 49.125 36.390 49.960 ;
        RECT 36.560 49.325 36.820 50.130 ;
        RECT 36.990 49.125 37.250 49.960 ;
        RECT 37.420 49.325 37.675 50.130 ;
        RECT 37.850 49.125 38.110 49.960 ;
        RECT 38.280 49.325 38.535 50.130 ;
        RECT 38.710 49.125 39.055 49.960 ;
        RECT 39.225 49.125 39.515 50.290 ;
        RECT 40.150 50.075 40.485 51.495 ;
        RECT 40.665 51.305 41.410 51.675 ;
        RECT 41.975 51.135 42.230 51.495 ;
        RECT 42.410 51.305 42.740 51.675 ;
        RECT 42.920 51.135 43.145 51.495 ;
        RECT 40.660 50.945 43.145 51.135 ;
        RECT 43.915 51.125 44.085 51.415 ;
        RECT 44.255 51.295 44.585 51.675 ;
        RECT 43.915 50.955 44.580 51.125 ;
        RECT 40.660 50.255 40.885 50.945 ;
        RECT 41.085 50.435 41.365 50.765 ;
        RECT 41.545 50.435 42.120 50.765 ;
        RECT 42.300 50.435 42.735 50.765 ;
        RECT 42.915 50.435 43.185 50.765 ;
        RECT 40.660 50.075 43.155 50.255 ;
        RECT 43.830 50.135 44.180 50.785 ;
        RECT 40.150 49.305 40.415 50.075 ;
        RECT 40.585 49.125 40.915 49.845 ;
        RECT 41.105 49.665 42.295 49.895 ;
        RECT 41.105 49.305 41.365 49.665 ;
        RECT 41.535 49.125 41.865 49.495 ;
        RECT 42.035 49.305 42.295 49.665 ;
        RECT 42.865 49.305 43.155 50.075 ;
        RECT 44.350 49.965 44.580 50.955 ;
        RECT 43.915 49.795 44.580 49.965 ;
        RECT 43.915 49.295 44.085 49.795 ;
        RECT 44.255 49.125 44.585 49.625 ;
        RECT 44.755 49.295 44.940 51.415 ;
        RECT 45.195 51.215 45.445 51.675 ;
        RECT 45.615 51.225 45.950 51.395 ;
        RECT 46.145 51.225 46.820 51.395 ;
        RECT 45.615 51.085 45.785 51.225 ;
        RECT 45.110 50.095 45.390 51.045 ;
        RECT 45.560 50.955 45.785 51.085 ;
        RECT 45.560 49.850 45.730 50.955 ;
        RECT 45.955 50.805 46.480 51.025 ;
        RECT 45.900 50.040 46.140 50.635 ;
        RECT 46.310 50.105 46.480 50.805 ;
        RECT 46.650 50.445 46.820 51.225 ;
        RECT 47.140 51.175 47.510 51.675 ;
        RECT 47.690 51.225 48.095 51.395 ;
        RECT 48.265 51.225 49.050 51.395 ;
        RECT 47.690 50.995 47.860 51.225 ;
        RECT 47.030 50.695 47.860 50.995 ;
        RECT 48.245 50.725 48.710 51.055 ;
        RECT 47.030 50.665 47.230 50.695 ;
        RECT 47.350 50.445 47.520 50.515 ;
        RECT 46.650 50.275 47.520 50.445 ;
        RECT 47.010 50.185 47.520 50.275 ;
        RECT 45.560 49.720 45.865 49.850 ;
        RECT 46.310 49.740 46.840 50.105 ;
        RECT 45.180 49.125 45.445 49.585 ;
        RECT 45.615 49.295 45.865 49.720 ;
        RECT 47.010 49.570 47.180 50.185 ;
        RECT 46.075 49.400 47.180 49.570 ;
        RECT 47.350 49.125 47.520 49.925 ;
        RECT 47.690 49.625 47.860 50.695 ;
        RECT 48.030 49.795 48.220 50.515 ;
        RECT 48.390 49.765 48.710 50.725 ;
        RECT 48.880 50.765 49.050 51.225 ;
        RECT 49.325 51.145 49.535 51.675 ;
        RECT 49.795 50.935 50.125 51.460 ;
        RECT 50.295 51.065 50.465 51.675 ;
        RECT 50.635 51.020 50.965 51.455 ;
        RECT 51.275 51.125 51.445 51.415 ;
        RECT 51.615 51.295 51.945 51.675 ;
        RECT 50.635 50.935 51.015 51.020 ;
        RECT 51.275 50.955 51.940 51.125 ;
        RECT 49.925 50.765 50.125 50.935 ;
        RECT 50.790 50.895 51.015 50.935 ;
        RECT 48.880 50.435 49.755 50.765 ;
        RECT 49.925 50.435 50.675 50.765 ;
        RECT 47.690 49.295 47.940 49.625 ;
        RECT 48.880 49.595 49.050 50.435 ;
        RECT 49.925 50.230 50.115 50.435 ;
        RECT 50.845 50.315 51.015 50.895 ;
        RECT 50.800 50.265 51.015 50.315 ;
        RECT 49.220 49.855 50.115 50.230 ;
        RECT 50.625 50.185 51.015 50.265 ;
        RECT 48.165 49.425 49.050 49.595 ;
        RECT 49.230 49.125 49.545 49.625 ;
        RECT 49.775 49.295 50.115 49.855 ;
        RECT 50.285 49.125 50.455 50.135 ;
        RECT 50.625 49.340 50.955 50.185 ;
        RECT 51.190 50.135 51.540 50.785 ;
        RECT 51.710 49.965 51.940 50.955 ;
        RECT 51.275 49.795 51.940 49.965 ;
        RECT 51.275 49.295 51.445 49.795 ;
        RECT 51.615 49.125 51.945 49.625 ;
        RECT 52.115 49.295 52.300 51.415 ;
        RECT 52.555 51.215 52.805 51.675 ;
        RECT 52.975 51.225 53.310 51.395 ;
        RECT 53.505 51.225 54.180 51.395 ;
        RECT 52.975 51.085 53.145 51.225 ;
        RECT 52.470 50.095 52.750 51.045 ;
        RECT 52.920 50.955 53.145 51.085 ;
        RECT 52.920 49.850 53.090 50.955 ;
        RECT 53.315 50.805 53.840 51.025 ;
        RECT 53.260 50.040 53.500 50.635 ;
        RECT 53.670 50.105 53.840 50.805 ;
        RECT 54.010 50.445 54.180 51.225 ;
        RECT 54.500 51.175 54.870 51.675 ;
        RECT 55.050 51.225 55.455 51.395 ;
        RECT 55.625 51.225 56.410 51.395 ;
        RECT 55.050 50.995 55.220 51.225 ;
        RECT 54.390 50.695 55.220 50.995 ;
        RECT 55.605 50.725 56.070 51.055 ;
        RECT 54.390 50.665 54.590 50.695 ;
        RECT 54.710 50.445 54.880 50.515 ;
        RECT 54.010 50.275 54.880 50.445 ;
        RECT 54.370 50.185 54.880 50.275 ;
        RECT 52.920 49.720 53.225 49.850 ;
        RECT 53.670 49.740 54.200 50.105 ;
        RECT 52.540 49.125 52.805 49.585 ;
        RECT 52.975 49.295 53.225 49.720 ;
        RECT 54.370 49.570 54.540 50.185 ;
        RECT 53.435 49.400 54.540 49.570 ;
        RECT 54.710 49.125 54.880 49.925 ;
        RECT 55.050 49.625 55.220 50.695 ;
        RECT 55.390 49.795 55.580 50.515 ;
        RECT 55.750 49.765 56.070 50.725 ;
        RECT 56.240 50.765 56.410 51.225 ;
        RECT 56.685 51.145 56.895 51.675 ;
        RECT 57.155 50.935 57.485 51.460 ;
        RECT 57.655 51.065 57.825 51.675 ;
        RECT 57.995 51.020 58.325 51.455 ;
        RECT 57.995 50.935 58.375 51.020 ;
        RECT 57.285 50.765 57.485 50.935 ;
        RECT 58.150 50.895 58.375 50.935 ;
        RECT 56.240 50.435 57.115 50.765 ;
        RECT 57.285 50.435 58.035 50.765 ;
        RECT 55.050 49.295 55.300 49.625 ;
        RECT 56.240 49.595 56.410 50.435 ;
        RECT 57.285 50.230 57.475 50.435 ;
        RECT 58.205 50.315 58.375 50.895 ;
        RECT 58.160 50.265 58.375 50.315 ;
        RECT 56.580 49.855 57.475 50.230 ;
        RECT 57.985 50.185 58.375 50.265 ;
        RECT 58.550 50.935 58.805 51.505 ;
        RECT 58.975 51.275 59.305 51.675 ;
        RECT 59.730 51.140 60.260 51.505 ;
        RECT 60.450 51.335 60.725 51.505 ;
        RECT 60.445 51.165 60.725 51.335 ;
        RECT 59.730 51.105 59.905 51.140 ;
        RECT 58.975 50.935 59.905 51.105 ;
        RECT 58.550 50.265 58.720 50.935 ;
        RECT 58.975 50.765 59.145 50.935 ;
        RECT 58.890 50.435 59.145 50.765 ;
        RECT 59.370 50.435 59.565 50.765 ;
        RECT 55.525 49.425 56.410 49.595 ;
        RECT 56.590 49.125 56.905 49.625 ;
        RECT 57.135 49.295 57.475 49.855 ;
        RECT 57.645 49.125 57.815 50.135 ;
        RECT 57.985 49.340 58.315 50.185 ;
        RECT 58.550 49.295 58.885 50.265 ;
        RECT 59.055 49.125 59.225 50.265 ;
        RECT 59.395 49.465 59.565 50.435 ;
        RECT 59.735 49.805 59.905 50.935 ;
        RECT 60.075 50.145 60.245 50.945 ;
        RECT 60.450 50.345 60.725 51.165 ;
        RECT 60.895 50.145 61.085 51.505 ;
        RECT 61.265 51.140 61.775 51.675 ;
        RECT 61.995 50.865 62.240 51.470 ;
        RECT 62.685 50.905 64.355 51.675 ;
        RECT 64.985 50.950 65.275 51.675 ;
        RECT 65.445 51.130 70.790 51.675 ;
        RECT 70.965 51.130 76.310 51.675 ;
        RECT 61.285 50.695 62.515 50.865 ;
        RECT 60.075 49.975 61.085 50.145 ;
        RECT 61.255 50.130 62.005 50.320 ;
        RECT 59.735 49.635 60.860 49.805 ;
        RECT 61.255 49.465 61.425 50.130 ;
        RECT 62.175 49.885 62.515 50.695 ;
        RECT 62.685 50.385 63.435 50.905 ;
        RECT 63.605 50.215 64.355 50.735 ;
        RECT 67.030 50.300 67.370 51.130 ;
        RECT 59.395 49.295 61.425 49.465 ;
        RECT 61.595 49.125 61.765 49.885 ;
        RECT 62.000 49.475 62.515 49.885 ;
        RECT 62.685 49.125 64.355 50.215 ;
        RECT 64.985 49.125 65.275 50.290 ;
        RECT 68.850 49.560 69.200 50.810 ;
        RECT 72.550 50.300 72.890 51.130 ;
        RECT 76.485 50.905 78.155 51.675 ;
        RECT 74.370 49.560 74.720 50.810 ;
        RECT 76.485 50.385 77.235 50.905 ;
        RECT 78.365 50.855 78.595 51.675 ;
        RECT 78.765 50.875 79.095 51.505 ;
        RECT 77.405 50.215 78.155 50.735 ;
        RECT 78.345 50.435 78.675 50.685 ;
        RECT 78.845 50.275 79.095 50.875 ;
        RECT 79.265 50.855 79.475 51.675 ;
        RECT 79.705 51.130 85.050 51.675 ;
        RECT 81.290 50.300 81.630 51.130 ;
        RECT 85.225 50.905 88.735 51.675 ;
        RECT 89.365 51.000 89.625 51.505 ;
        RECT 89.805 51.295 90.135 51.675 ;
        RECT 90.315 51.125 90.485 51.505 ;
        RECT 65.445 49.125 70.790 49.560 ;
        RECT 70.965 49.125 76.310 49.560 ;
        RECT 76.485 49.125 78.155 50.215 ;
        RECT 78.365 49.125 78.595 50.265 ;
        RECT 78.765 49.295 79.095 50.275 ;
        RECT 79.265 49.125 79.475 50.265 ;
        RECT 83.110 49.560 83.460 50.810 ;
        RECT 85.225 50.385 86.875 50.905 ;
        RECT 87.045 50.215 88.735 50.735 ;
        RECT 79.705 49.125 85.050 49.560 ;
        RECT 85.225 49.125 88.735 50.215 ;
        RECT 89.365 50.200 89.535 51.000 ;
        RECT 89.820 50.955 90.485 51.125 ;
        RECT 89.820 50.700 89.990 50.955 ;
        RECT 90.745 50.925 91.955 51.675 ;
        RECT 89.705 50.370 89.990 50.700 ;
        RECT 90.225 50.405 90.555 50.775 ;
        RECT 89.820 50.225 89.990 50.370 ;
        RECT 89.365 49.295 89.635 50.200 ;
        RECT 89.820 50.055 90.485 50.225 ;
        RECT 89.805 49.125 90.135 49.885 ;
        RECT 90.315 49.295 90.485 50.055 ;
        RECT 90.745 50.215 91.265 50.755 ;
        RECT 91.435 50.385 91.955 50.925 ;
        RECT 90.745 49.125 91.955 50.215 ;
        RECT 13.380 48.955 92.040 49.125 ;
        RECT 13.465 47.865 14.675 48.955 ;
        RECT 13.465 47.155 13.985 47.695 ;
        RECT 14.155 47.325 14.675 47.865 ;
        RECT 14.850 47.805 15.110 48.955 ;
        RECT 15.285 47.880 15.540 48.785 ;
        RECT 15.710 48.195 16.040 48.955 ;
        RECT 16.255 48.025 16.425 48.785 ;
        RECT 13.465 46.405 14.675 47.155 ;
        RECT 14.850 46.405 15.110 47.245 ;
        RECT 15.285 47.150 15.455 47.880 ;
        RECT 15.710 47.855 16.425 48.025 ;
        RECT 17.810 47.985 18.140 48.785 ;
        RECT 18.310 48.155 18.640 48.955 ;
        RECT 18.940 47.985 19.270 48.785 ;
        RECT 19.915 48.155 20.165 48.955 ;
        RECT 15.710 47.645 15.880 47.855 ;
        RECT 17.810 47.815 20.245 47.985 ;
        RECT 20.435 47.815 20.605 48.955 ;
        RECT 20.775 47.815 21.115 48.785 ;
        RECT 15.625 47.315 15.880 47.645 ;
        RECT 15.285 46.575 15.540 47.150 ;
        RECT 15.710 47.125 15.880 47.315 ;
        RECT 16.160 47.305 16.515 47.675 ;
        RECT 17.605 47.395 17.955 47.645 ;
        RECT 18.140 47.185 18.310 47.815 ;
        RECT 18.480 47.395 18.810 47.595 ;
        RECT 18.980 47.395 19.310 47.595 ;
        RECT 19.480 47.395 19.900 47.595 ;
        RECT 20.075 47.565 20.245 47.815 ;
        RECT 20.075 47.395 20.770 47.565 ;
        RECT 15.710 46.955 16.425 47.125 ;
        RECT 15.710 46.405 16.040 46.785 ;
        RECT 16.255 46.575 16.425 46.955 ;
        RECT 17.810 46.575 18.310 47.185 ;
        RECT 18.940 47.055 20.165 47.225 ;
        RECT 20.940 47.205 21.115 47.815 ;
        RECT 21.290 47.805 21.550 48.955 ;
        RECT 21.725 47.880 21.980 48.785 ;
        RECT 22.150 48.195 22.480 48.955 ;
        RECT 22.695 48.025 22.865 48.785 ;
        RECT 18.940 46.575 19.270 47.055 ;
        RECT 19.440 46.405 19.665 46.865 ;
        RECT 19.835 46.575 20.165 47.055 ;
        RECT 20.355 46.405 20.605 47.205 ;
        RECT 20.775 46.575 21.115 47.205 ;
        RECT 21.290 46.405 21.550 47.245 ;
        RECT 21.725 47.150 21.895 47.880 ;
        RECT 22.150 47.855 22.865 48.025 ;
        RECT 23.125 47.865 25.715 48.955 ;
        RECT 22.150 47.645 22.320 47.855 ;
        RECT 22.065 47.315 22.320 47.645 ;
        RECT 21.725 46.575 21.980 47.150 ;
        RECT 22.150 47.125 22.320 47.315 ;
        RECT 22.600 47.305 22.955 47.675 ;
        RECT 23.125 47.175 24.335 47.695 ;
        RECT 24.505 47.345 25.715 47.865 ;
        RECT 26.345 47.790 26.635 48.955 ;
        RECT 27.470 47.985 27.800 48.785 ;
        RECT 27.970 48.155 28.300 48.955 ;
        RECT 28.600 47.985 28.930 48.785 ;
        RECT 29.575 48.155 29.825 48.955 ;
        RECT 27.470 47.815 29.905 47.985 ;
        RECT 30.095 47.815 30.265 48.955 ;
        RECT 30.435 47.815 30.775 48.785 ;
        RECT 31.035 48.285 31.205 48.785 ;
        RECT 31.375 48.455 31.705 48.955 ;
        RECT 31.035 48.115 31.700 48.285 ;
        RECT 27.265 47.395 27.615 47.645 ;
        RECT 27.800 47.185 27.970 47.815 ;
        RECT 28.140 47.395 28.470 47.595 ;
        RECT 28.640 47.395 28.970 47.595 ;
        RECT 29.140 47.395 29.560 47.595 ;
        RECT 29.735 47.565 29.905 47.815 ;
        RECT 29.735 47.395 30.430 47.565 ;
        RECT 30.600 47.255 30.775 47.815 ;
        RECT 30.950 47.295 31.300 47.945 ;
        RECT 22.150 46.955 22.865 47.125 ;
        RECT 22.150 46.405 22.480 46.785 ;
        RECT 22.695 46.575 22.865 46.955 ;
        RECT 23.125 46.405 25.715 47.175 ;
        RECT 26.345 46.405 26.635 47.130 ;
        RECT 27.470 46.575 27.970 47.185 ;
        RECT 28.600 47.055 29.825 47.225 ;
        RECT 30.545 47.205 30.775 47.255 ;
        RECT 28.600 46.575 28.930 47.055 ;
        RECT 29.100 46.405 29.325 46.865 ;
        RECT 29.495 46.575 29.825 47.055 ;
        RECT 30.015 46.405 30.265 47.205 ;
        RECT 30.435 46.575 30.775 47.205 ;
        RECT 31.470 47.125 31.700 48.115 ;
        RECT 31.035 46.955 31.700 47.125 ;
        RECT 31.035 46.665 31.205 46.955 ;
        RECT 31.375 46.405 31.705 46.785 ;
        RECT 31.875 46.665 32.060 48.785 ;
        RECT 32.300 48.495 32.565 48.955 ;
        RECT 32.735 48.360 32.985 48.785 ;
        RECT 33.195 48.510 34.300 48.680 ;
        RECT 32.680 48.230 32.985 48.360 ;
        RECT 32.230 47.035 32.510 47.985 ;
        RECT 32.680 47.125 32.850 48.230 ;
        RECT 33.020 47.445 33.260 48.040 ;
        RECT 33.430 47.975 33.960 48.340 ;
        RECT 33.430 47.275 33.600 47.975 ;
        RECT 34.130 47.895 34.300 48.510 ;
        RECT 34.470 48.155 34.640 48.955 ;
        RECT 34.810 48.455 35.060 48.785 ;
        RECT 35.285 48.485 36.170 48.655 ;
        RECT 34.130 47.805 34.640 47.895 ;
        RECT 32.680 46.995 32.905 47.125 ;
        RECT 33.075 47.055 33.600 47.275 ;
        RECT 33.770 47.635 34.640 47.805 ;
        RECT 32.315 46.405 32.565 46.865 ;
        RECT 32.735 46.855 32.905 46.995 ;
        RECT 33.770 46.855 33.940 47.635 ;
        RECT 34.470 47.565 34.640 47.635 ;
        RECT 34.150 47.385 34.350 47.415 ;
        RECT 34.810 47.385 34.980 48.455 ;
        RECT 35.150 47.565 35.340 48.285 ;
        RECT 34.150 47.085 34.980 47.385 ;
        RECT 35.510 47.355 35.830 48.315 ;
        RECT 32.735 46.685 33.070 46.855 ;
        RECT 33.265 46.685 33.940 46.855 ;
        RECT 34.260 46.405 34.630 46.905 ;
        RECT 34.810 46.855 34.980 47.085 ;
        RECT 35.365 47.025 35.830 47.355 ;
        RECT 36.000 47.645 36.170 48.485 ;
        RECT 36.350 48.455 36.665 48.955 ;
        RECT 36.895 48.225 37.235 48.785 ;
        RECT 36.340 47.850 37.235 48.225 ;
        RECT 37.405 47.945 37.575 48.955 ;
        RECT 37.045 47.645 37.235 47.850 ;
        RECT 37.745 47.895 38.075 48.740 ;
        RECT 38.395 48.285 38.565 48.785 ;
        RECT 38.735 48.455 39.065 48.955 ;
        RECT 38.395 48.115 39.060 48.285 ;
        RECT 37.745 47.815 38.135 47.895 ;
        RECT 37.920 47.765 38.135 47.815 ;
        RECT 36.000 47.315 36.875 47.645 ;
        RECT 37.045 47.315 37.795 47.645 ;
        RECT 36.000 46.855 36.170 47.315 ;
        RECT 37.045 47.145 37.245 47.315 ;
        RECT 37.965 47.185 38.135 47.765 ;
        RECT 38.310 47.295 38.660 47.945 ;
        RECT 37.910 47.145 38.135 47.185 ;
        RECT 34.810 46.685 35.215 46.855 ;
        RECT 35.385 46.685 36.170 46.855 ;
        RECT 36.445 46.405 36.655 46.935 ;
        RECT 36.915 46.620 37.245 47.145 ;
        RECT 37.755 47.060 38.135 47.145 ;
        RECT 38.830 47.125 39.060 48.115 ;
        RECT 37.415 46.405 37.585 47.015 ;
        RECT 37.755 46.625 38.085 47.060 ;
        RECT 38.395 46.955 39.060 47.125 ;
        RECT 38.395 46.665 38.565 46.955 ;
        RECT 38.735 46.405 39.065 46.785 ;
        RECT 39.235 46.665 39.420 48.785 ;
        RECT 39.660 48.495 39.925 48.955 ;
        RECT 40.095 48.360 40.345 48.785 ;
        RECT 40.555 48.510 41.660 48.680 ;
        RECT 40.040 48.230 40.345 48.360 ;
        RECT 39.590 47.035 39.870 47.985 ;
        RECT 40.040 47.125 40.210 48.230 ;
        RECT 40.380 47.445 40.620 48.040 ;
        RECT 40.790 47.975 41.320 48.340 ;
        RECT 40.790 47.275 40.960 47.975 ;
        RECT 41.490 47.895 41.660 48.510 ;
        RECT 41.830 48.155 42.000 48.955 ;
        RECT 42.170 48.455 42.420 48.785 ;
        RECT 42.645 48.485 43.530 48.655 ;
        RECT 41.490 47.805 42.000 47.895 ;
        RECT 40.040 46.995 40.265 47.125 ;
        RECT 40.435 47.055 40.960 47.275 ;
        RECT 41.130 47.635 42.000 47.805 ;
        RECT 39.675 46.405 39.925 46.865 ;
        RECT 40.095 46.855 40.265 46.995 ;
        RECT 41.130 46.855 41.300 47.635 ;
        RECT 41.830 47.565 42.000 47.635 ;
        RECT 41.510 47.385 41.710 47.415 ;
        RECT 42.170 47.385 42.340 48.455 ;
        RECT 42.510 47.565 42.700 48.285 ;
        RECT 41.510 47.085 42.340 47.385 ;
        RECT 42.870 47.355 43.190 48.315 ;
        RECT 40.095 46.685 40.430 46.855 ;
        RECT 40.625 46.685 41.300 46.855 ;
        RECT 41.620 46.405 41.990 46.905 ;
        RECT 42.170 46.855 42.340 47.085 ;
        RECT 42.725 47.025 43.190 47.355 ;
        RECT 43.360 47.645 43.530 48.485 ;
        RECT 43.710 48.455 44.025 48.955 ;
        RECT 44.255 48.225 44.595 48.785 ;
        RECT 43.700 47.850 44.595 48.225 ;
        RECT 44.765 47.945 44.935 48.955 ;
        RECT 44.405 47.645 44.595 47.850 ;
        RECT 45.105 47.895 45.435 48.740 ;
        RECT 45.105 47.815 45.495 47.895 ;
        RECT 45.280 47.765 45.495 47.815 ;
        RECT 43.360 47.315 44.235 47.645 ;
        RECT 44.405 47.315 45.155 47.645 ;
        RECT 43.360 46.855 43.530 47.315 ;
        RECT 44.405 47.145 44.605 47.315 ;
        RECT 45.325 47.185 45.495 47.765 ;
        RECT 45.270 47.145 45.495 47.185 ;
        RECT 42.170 46.685 42.575 46.855 ;
        RECT 42.745 46.685 43.530 46.855 ;
        RECT 43.805 46.405 44.015 46.935 ;
        RECT 44.275 46.620 44.605 47.145 ;
        RECT 45.115 47.060 45.495 47.145 ;
        RECT 45.670 47.815 46.005 48.785 ;
        RECT 46.175 47.815 46.345 48.955 ;
        RECT 46.515 48.615 48.545 48.785 ;
        RECT 45.670 47.145 45.840 47.815 ;
        RECT 46.515 47.645 46.685 48.615 ;
        RECT 46.010 47.315 46.265 47.645 ;
        RECT 46.490 47.315 46.685 47.645 ;
        RECT 46.855 48.275 47.980 48.445 ;
        RECT 46.095 47.145 46.265 47.315 ;
        RECT 46.855 47.145 47.025 48.275 ;
        RECT 44.775 46.405 44.945 47.015 ;
        RECT 45.115 46.625 45.445 47.060 ;
        RECT 45.670 46.575 45.925 47.145 ;
        RECT 46.095 46.975 47.025 47.145 ;
        RECT 47.195 47.935 48.205 48.105 ;
        RECT 47.195 47.135 47.365 47.935 ;
        RECT 47.570 47.255 47.845 47.735 ;
        RECT 47.565 47.085 47.845 47.255 ;
        RECT 46.850 46.940 47.025 46.975 ;
        RECT 46.095 46.405 46.425 46.805 ;
        RECT 46.850 46.575 47.380 46.940 ;
        RECT 47.570 46.575 47.845 47.085 ;
        RECT 48.015 46.575 48.205 47.935 ;
        RECT 48.375 47.950 48.545 48.615 ;
        RECT 48.715 48.195 48.885 48.955 ;
        RECT 49.120 48.195 49.635 48.605 ;
        RECT 48.375 47.760 49.125 47.950 ;
        RECT 49.295 47.385 49.635 48.195 ;
        RECT 49.805 47.865 51.475 48.955 ;
        RECT 48.405 47.215 49.635 47.385 ;
        RECT 48.385 46.405 48.895 46.940 ;
        RECT 49.115 46.610 49.360 47.215 ;
        RECT 49.805 47.175 50.555 47.695 ;
        RECT 50.725 47.345 51.475 47.865 ;
        RECT 52.105 47.790 52.395 48.955 ;
        RECT 52.565 47.815 52.950 48.785 ;
        RECT 53.120 48.495 53.445 48.955 ;
        RECT 53.965 48.325 54.245 48.785 ;
        RECT 53.120 48.105 54.245 48.325 ;
        RECT 49.805 46.405 51.475 47.175 ;
        RECT 52.565 47.145 52.845 47.815 ;
        RECT 53.120 47.645 53.570 48.105 ;
        RECT 54.435 47.935 54.835 48.785 ;
        RECT 55.235 48.495 55.505 48.955 ;
        RECT 55.675 48.325 55.960 48.785 ;
        RECT 56.245 48.450 56.875 48.955 ;
        RECT 53.015 47.315 53.570 47.645 ;
        RECT 53.740 47.375 54.835 47.935 ;
        RECT 53.120 47.205 53.570 47.315 ;
        RECT 52.105 46.405 52.395 47.130 ;
        RECT 52.565 46.575 52.950 47.145 ;
        RECT 53.120 47.035 54.245 47.205 ;
        RECT 53.120 46.405 53.445 46.865 ;
        RECT 53.965 46.575 54.245 47.035 ;
        RECT 54.435 46.575 54.835 47.375 ;
        RECT 55.005 48.105 55.960 48.325 ;
        RECT 55.005 47.205 55.215 48.105 ;
        RECT 55.385 47.375 56.075 47.935 ;
        RECT 56.260 47.915 56.515 48.280 ;
        RECT 56.685 48.275 56.875 48.450 ;
        RECT 57.055 48.445 57.530 48.785 ;
        RECT 56.685 48.085 57.015 48.275 ;
        RECT 57.240 47.915 57.490 48.210 ;
        RECT 57.715 48.110 57.930 48.955 ;
        RECT 58.130 48.115 58.405 48.785 ;
        RECT 56.260 47.745 58.050 47.915 ;
        RECT 58.235 47.765 58.405 48.115 ;
        RECT 58.575 47.945 58.835 48.955 ;
        RECT 59.005 47.985 59.275 48.755 ;
        RECT 59.445 48.175 59.775 48.955 ;
        RECT 59.980 48.350 60.165 48.755 ;
        RECT 60.335 48.530 60.670 48.955 ;
        RECT 59.980 48.175 60.645 48.350 ;
        RECT 59.005 47.815 60.135 47.985 ;
        RECT 55.005 47.035 55.960 47.205 ;
        RECT 56.245 47.085 56.630 47.565 ;
        RECT 55.235 46.405 55.505 46.865 ;
        RECT 55.675 46.575 55.960 47.035 ;
        RECT 56.800 46.890 57.055 47.745 ;
        RECT 56.265 46.625 57.055 46.890 ;
        RECT 57.225 47.070 57.635 47.565 ;
        RECT 57.820 47.315 58.050 47.745 ;
        RECT 58.220 47.245 58.835 47.765 ;
        RECT 57.225 46.625 57.455 47.070 ;
        RECT 58.220 47.035 58.390 47.245 ;
        RECT 57.635 46.405 57.965 46.900 ;
        RECT 58.140 46.575 58.390 47.035 ;
        RECT 58.560 46.405 58.835 47.065 ;
        RECT 59.005 46.905 59.175 47.815 ;
        RECT 59.345 47.065 59.705 47.645 ;
        RECT 59.885 47.315 60.135 47.815 ;
        RECT 60.305 47.145 60.645 48.175 ;
        RECT 60.845 47.865 62.055 48.955 ;
        RECT 59.960 46.975 60.645 47.145 ;
        RECT 60.845 47.155 61.365 47.695 ;
        RECT 61.535 47.325 62.055 47.865 ;
        RECT 62.225 48.105 62.485 48.785 ;
        RECT 62.655 48.175 62.905 48.955 ;
        RECT 63.155 48.405 63.405 48.785 ;
        RECT 63.575 48.575 63.930 48.955 ;
        RECT 64.935 48.565 65.270 48.785 ;
        RECT 64.535 48.405 64.765 48.445 ;
        RECT 63.155 48.205 64.765 48.405 ;
        RECT 63.155 48.195 63.990 48.205 ;
        RECT 64.580 48.115 64.765 48.205 ;
        RECT 59.005 46.575 59.265 46.905 ;
        RECT 59.475 46.405 59.750 46.885 ;
        RECT 59.960 46.575 60.165 46.975 ;
        RECT 60.335 46.405 60.670 46.805 ;
        RECT 60.845 46.405 62.055 47.155 ;
        RECT 62.225 46.905 62.395 48.105 ;
        RECT 64.095 48.005 64.425 48.035 ;
        RECT 62.625 47.945 64.425 48.005 ;
        RECT 65.015 47.945 65.270 48.565 ;
        RECT 65.445 48.360 65.880 48.785 ;
        RECT 66.050 48.530 66.435 48.955 ;
        RECT 65.445 48.190 66.435 48.360 ;
        RECT 62.565 47.835 65.270 47.945 ;
        RECT 62.565 47.800 62.765 47.835 ;
        RECT 62.565 47.225 62.735 47.800 ;
        RECT 64.095 47.775 65.270 47.835 ;
        RECT 62.965 47.360 63.375 47.665 ;
        RECT 63.545 47.395 63.875 47.605 ;
        RECT 62.565 47.105 62.835 47.225 ;
        RECT 62.565 47.060 63.410 47.105 ;
        RECT 62.655 46.935 63.410 47.060 ;
        RECT 63.665 46.995 63.875 47.395 ;
        RECT 64.120 47.395 64.595 47.605 ;
        RECT 64.785 47.395 65.275 47.595 ;
        RECT 64.120 46.995 64.340 47.395 ;
        RECT 65.445 47.315 65.930 48.020 ;
        RECT 66.100 47.645 66.435 48.190 ;
        RECT 66.605 47.995 67.030 48.785 ;
        RECT 67.200 48.360 67.475 48.785 ;
        RECT 67.645 48.530 68.030 48.955 ;
        RECT 67.200 48.165 68.030 48.360 ;
        RECT 66.605 47.815 67.510 47.995 ;
        RECT 66.100 47.315 66.510 47.645 ;
        RECT 66.680 47.315 67.510 47.815 ;
        RECT 67.680 47.645 68.030 48.165 ;
        RECT 68.200 47.995 68.445 48.785 ;
        RECT 68.635 48.360 68.890 48.785 ;
        RECT 69.060 48.530 69.445 48.955 ;
        RECT 68.635 48.165 69.445 48.360 ;
        RECT 68.200 47.815 68.925 47.995 ;
        RECT 67.680 47.315 68.105 47.645 ;
        RECT 68.275 47.315 68.925 47.815 ;
        RECT 69.095 47.645 69.445 48.165 ;
        RECT 69.615 47.815 69.875 48.785 ;
        RECT 69.095 47.315 69.520 47.645 ;
        RECT 62.225 46.575 62.485 46.905 ;
        RECT 63.240 46.785 63.410 46.935 ;
        RECT 62.655 46.405 62.985 46.765 ;
        RECT 63.240 46.575 64.540 46.785 ;
        RECT 64.815 46.405 65.270 47.170 ;
        RECT 66.100 47.145 66.435 47.315 ;
        RECT 66.680 47.145 67.030 47.315 ;
        RECT 67.680 47.145 68.030 47.315 ;
        RECT 68.275 47.145 68.445 47.315 ;
        RECT 69.095 47.145 69.445 47.315 ;
        RECT 69.690 47.145 69.875 47.815 ;
        RECT 70.050 48.565 70.385 48.785 ;
        RECT 71.390 48.575 71.745 48.955 ;
        RECT 70.050 47.945 70.305 48.565 ;
        RECT 70.555 48.405 70.785 48.445 ;
        RECT 71.915 48.405 72.165 48.785 ;
        RECT 70.555 48.205 72.165 48.405 ;
        RECT 70.555 48.115 70.740 48.205 ;
        RECT 71.330 48.195 72.165 48.205 ;
        RECT 72.415 48.175 72.665 48.955 ;
        RECT 72.835 48.105 73.095 48.785 ;
        RECT 70.895 48.005 71.225 48.035 ;
        RECT 70.895 47.945 72.695 48.005 ;
        RECT 70.050 47.835 72.755 47.945 ;
        RECT 70.050 47.775 71.225 47.835 ;
        RECT 72.555 47.800 72.755 47.835 ;
        RECT 70.045 47.395 70.535 47.595 ;
        RECT 70.725 47.395 71.200 47.605 ;
        RECT 65.445 46.975 66.435 47.145 ;
        RECT 65.445 46.575 65.880 46.975 ;
        RECT 66.050 46.405 66.435 46.805 ;
        RECT 66.605 46.575 67.030 47.145 ;
        RECT 67.220 46.975 68.030 47.145 ;
        RECT 67.220 46.575 67.475 46.975 ;
        RECT 67.645 46.405 68.030 46.805 ;
        RECT 68.200 46.575 68.445 47.145 ;
        RECT 68.635 46.975 69.445 47.145 ;
        RECT 68.635 46.575 68.890 46.975 ;
        RECT 69.060 46.405 69.445 46.805 ;
        RECT 69.615 46.575 69.875 47.145 ;
        RECT 70.050 46.405 70.505 47.170 ;
        RECT 70.980 46.995 71.200 47.395 ;
        RECT 71.445 47.395 71.775 47.605 ;
        RECT 71.445 46.995 71.655 47.395 ;
        RECT 71.945 47.360 72.355 47.665 ;
        RECT 72.585 47.225 72.755 47.800 ;
        RECT 72.485 47.105 72.755 47.225 ;
        RECT 71.910 47.060 72.755 47.105 ;
        RECT 71.910 46.935 72.665 47.060 ;
        RECT 71.910 46.785 72.080 46.935 ;
        RECT 72.925 46.905 73.095 48.105 ;
        RECT 70.780 46.575 72.080 46.785 ;
        RECT 72.335 46.405 72.665 46.765 ;
        RECT 72.835 46.575 73.095 46.905 ;
        RECT 73.300 48.165 73.835 48.785 ;
        RECT 73.300 47.145 73.615 48.165 ;
        RECT 74.005 48.155 74.335 48.955 ;
        RECT 74.820 47.985 75.210 48.160 ;
        RECT 73.785 47.815 75.210 47.985 ;
        RECT 75.565 47.865 77.235 48.955 ;
        RECT 73.785 47.315 73.955 47.815 ;
        RECT 73.300 46.575 73.915 47.145 ;
        RECT 74.205 47.085 74.470 47.645 ;
        RECT 74.640 46.915 74.810 47.815 ;
        RECT 74.980 47.085 75.335 47.645 ;
        RECT 75.565 47.175 76.315 47.695 ;
        RECT 76.485 47.345 77.235 47.865 ;
        RECT 77.865 47.790 78.155 48.955 ;
        RECT 78.530 47.985 78.860 48.785 ;
        RECT 79.030 48.155 79.360 48.955 ;
        RECT 79.660 47.985 79.990 48.785 ;
        RECT 80.635 48.155 80.885 48.955 ;
        RECT 78.530 47.815 80.965 47.985 ;
        RECT 81.155 47.815 81.325 48.955 ;
        RECT 81.495 47.815 81.835 48.785 ;
        RECT 82.005 48.520 87.350 48.955 ;
        RECT 78.325 47.395 78.675 47.645 ;
        RECT 78.860 47.185 79.030 47.815 ;
        RECT 79.200 47.395 79.530 47.595 ;
        RECT 79.700 47.395 80.030 47.595 ;
        RECT 80.200 47.395 80.620 47.595 ;
        RECT 80.795 47.565 80.965 47.815 ;
        RECT 80.795 47.395 81.490 47.565 ;
        RECT 74.085 46.405 74.300 46.915 ;
        RECT 74.530 46.585 74.810 46.915 ;
        RECT 74.990 46.405 75.230 46.915 ;
        RECT 75.565 46.405 77.235 47.175 ;
        RECT 77.865 46.405 78.155 47.130 ;
        RECT 78.530 46.575 79.030 47.185 ;
        RECT 79.660 47.055 80.885 47.225 ;
        RECT 81.660 47.205 81.835 47.815 ;
        RECT 79.660 46.575 79.990 47.055 ;
        RECT 80.160 46.405 80.385 46.865 ;
        RECT 80.555 46.575 80.885 47.055 ;
        RECT 81.075 46.405 81.325 47.205 ;
        RECT 81.495 46.575 81.835 47.205 ;
        RECT 83.590 46.950 83.930 47.780 ;
        RECT 85.410 47.270 85.760 48.520 ;
        RECT 87.525 47.865 90.115 48.955 ;
        RECT 87.525 47.175 88.735 47.695 ;
        RECT 88.905 47.345 90.115 47.865 ;
        RECT 90.745 47.865 91.955 48.955 ;
        RECT 90.745 47.325 91.265 47.865 ;
        RECT 82.005 46.405 87.350 46.950 ;
        RECT 87.525 46.405 90.115 47.175 ;
        RECT 91.435 47.155 91.955 47.695 ;
        RECT 90.745 46.405 91.955 47.155 ;
        RECT 13.380 46.235 92.040 46.405 ;
        RECT 13.465 45.485 14.675 46.235 ;
        RECT 14.845 45.485 16.055 46.235 ;
        RECT 16.390 45.725 16.630 46.235 ;
        RECT 16.810 45.725 17.090 46.055 ;
        RECT 17.320 45.725 17.535 46.235 ;
        RECT 13.465 44.945 13.985 45.485 ;
        RECT 14.155 44.775 14.675 45.315 ;
        RECT 14.845 44.945 15.365 45.485 ;
        RECT 15.535 44.775 16.055 45.315 ;
        RECT 16.285 44.995 16.640 45.555 ;
        RECT 16.810 44.825 16.980 45.725 ;
        RECT 17.150 44.995 17.415 45.555 ;
        RECT 17.705 45.495 18.320 46.065 ;
        RECT 18.615 45.685 18.785 45.975 ;
        RECT 18.955 45.855 19.285 46.235 ;
        RECT 18.615 45.515 19.280 45.685 ;
        RECT 17.665 44.825 17.835 45.325 ;
        RECT 13.465 43.685 14.675 44.775 ;
        RECT 14.845 43.685 16.055 44.775 ;
        RECT 16.410 44.655 17.835 44.825 ;
        RECT 16.410 44.480 16.800 44.655 ;
        RECT 17.285 43.685 17.615 44.485 ;
        RECT 18.005 44.475 18.320 45.495 ;
        RECT 18.530 44.695 18.880 45.345 ;
        RECT 19.050 44.525 19.280 45.515 ;
        RECT 17.785 43.855 18.320 44.475 ;
        RECT 18.615 44.355 19.280 44.525 ;
        RECT 18.615 43.855 18.785 44.355 ;
        RECT 18.955 43.685 19.285 44.185 ;
        RECT 19.455 43.855 19.640 45.975 ;
        RECT 19.895 45.775 20.145 46.235 ;
        RECT 20.315 45.785 20.650 45.955 ;
        RECT 20.845 45.785 21.520 45.955 ;
        RECT 20.315 45.645 20.485 45.785 ;
        RECT 19.810 44.655 20.090 45.605 ;
        RECT 20.260 45.515 20.485 45.645 ;
        RECT 20.260 44.410 20.430 45.515 ;
        RECT 20.655 45.365 21.180 45.585 ;
        RECT 20.600 44.600 20.840 45.195 ;
        RECT 21.010 44.665 21.180 45.365 ;
        RECT 21.350 45.005 21.520 45.785 ;
        RECT 21.840 45.735 22.210 46.235 ;
        RECT 22.390 45.785 22.795 45.955 ;
        RECT 22.965 45.785 23.750 45.955 ;
        RECT 22.390 45.555 22.560 45.785 ;
        RECT 21.730 45.255 22.560 45.555 ;
        RECT 22.945 45.285 23.410 45.615 ;
        RECT 21.730 45.225 21.930 45.255 ;
        RECT 22.050 45.005 22.220 45.075 ;
        RECT 21.350 44.835 22.220 45.005 ;
        RECT 21.710 44.745 22.220 44.835 ;
        RECT 20.260 44.280 20.565 44.410 ;
        RECT 21.010 44.300 21.540 44.665 ;
        RECT 19.880 43.685 20.145 44.145 ;
        RECT 20.315 43.855 20.565 44.280 ;
        RECT 21.710 44.130 21.880 44.745 ;
        RECT 20.775 43.960 21.880 44.130 ;
        RECT 22.050 43.685 22.220 44.485 ;
        RECT 22.390 44.185 22.560 45.255 ;
        RECT 22.730 44.355 22.920 45.075 ;
        RECT 23.090 44.325 23.410 45.285 ;
        RECT 23.580 45.325 23.750 45.785 ;
        RECT 24.025 45.705 24.235 46.235 ;
        RECT 24.495 45.495 24.825 46.020 ;
        RECT 24.995 45.625 25.165 46.235 ;
        RECT 25.335 45.580 25.665 46.015 ;
        RECT 26.050 45.725 26.290 46.235 ;
        RECT 26.470 45.725 26.750 46.055 ;
        RECT 26.980 45.725 27.195 46.235 ;
        RECT 25.335 45.495 25.715 45.580 ;
        RECT 24.625 45.325 24.825 45.495 ;
        RECT 25.490 45.455 25.715 45.495 ;
        RECT 23.580 44.995 24.455 45.325 ;
        RECT 24.625 44.995 25.375 45.325 ;
        RECT 22.390 43.855 22.640 44.185 ;
        RECT 23.580 44.155 23.750 44.995 ;
        RECT 24.625 44.790 24.815 44.995 ;
        RECT 25.545 44.875 25.715 45.455 ;
        RECT 25.945 44.995 26.300 45.555 ;
        RECT 25.500 44.825 25.715 44.875 ;
        RECT 26.470 44.825 26.640 45.725 ;
        RECT 26.810 44.995 27.075 45.555 ;
        RECT 27.365 45.495 27.980 46.065 ;
        RECT 27.325 44.825 27.495 45.325 ;
        RECT 23.920 44.415 24.815 44.790 ;
        RECT 25.325 44.745 25.715 44.825 ;
        RECT 22.865 43.985 23.750 44.155 ;
        RECT 23.930 43.685 24.245 44.185 ;
        RECT 24.475 43.855 24.815 44.415 ;
        RECT 24.985 43.685 25.155 44.695 ;
        RECT 25.325 43.900 25.655 44.745 ;
        RECT 26.070 44.655 27.495 44.825 ;
        RECT 26.070 44.480 26.460 44.655 ;
        RECT 26.945 43.685 27.275 44.485 ;
        RECT 27.665 44.475 27.980 45.495 ;
        RECT 28.390 45.455 28.890 46.065 ;
        RECT 28.185 44.995 28.535 45.245 ;
        RECT 28.720 44.825 28.890 45.455 ;
        RECT 29.520 45.585 29.850 46.065 ;
        RECT 30.020 45.775 30.245 46.235 ;
        RECT 30.415 45.585 30.745 46.065 ;
        RECT 29.520 45.415 30.745 45.585 ;
        RECT 30.935 45.435 31.185 46.235 ;
        RECT 31.355 45.435 31.695 46.065 ;
        RECT 31.955 45.685 32.125 45.975 ;
        RECT 32.295 45.855 32.625 46.235 ;
        RECT 31.955 45.515 32.620 45.685 ;
        RECT 29.060 45.045 29.390 45.245 ;
        RECT 29.560 45.045 29.890 45.245 ;
        RECT 30.060 45.045 30.480 45.245 ;
        RECT 30.655 45.075 31.350 45.245 ;
        RECT 30.655 44.825 30.825 45.075 ;
        RECT 31.520 44.875 31.695 45.435 ;
        RECT 31.465 44.825 31.695 44.875 ;
        RECT 27.445 43.855 27.980 44.475 ;
        RECT 28.390 44.655 30.825 44.825 ;
        RECT 28.390 43.855 28.720 44.655 ;
        RECT 28.890 43.685 29.220 44.485 ;
        RECT 29.520 43.855 29.850 44.655 ;
        RECT 30.495 43.685 30.745 44.485 ;
        RECT 31.015 43.685 31.185 44.825 ;
        RECT 31.355 43.855 31.695 44.825 ;
        RECT 31.870 44.695 32.220 45.345 ;
        RECT 32.390 44.525 32.620 45.515 ;
        RECT 31.955 44.355 32.620 44.525 ;
        RECT 31.955 43.855 32.125 44.355 ;
        RECT 32.295 43.685 32.625 44.185 ;
        RECT 32.795 43.855 32.980 45.975 ;
        RECT 33.235 45.775 33.485 46.235 ;
        RECT 33.655 45.785 33.990 45.955 ;
        RECT 34.185 45.785 34.860 45.955 ;
        RECT 33.655 45.645 33.825 45.785 ;
        RECT 33.150 44.655 33.430 45.605 ;
        RECT 33.600 45.515 33.825 45.645 ;
        RECT 33.600 44.410 33.770 45.515 ;
        RECT 33.995 45.365 34.520 45.585 ;
        RECT 33.940 44.600 34.180 45.195 ;
        RECT 34.350 44.665 34.520 45.365 ;
        RECT 34.690 45.005 34.860 45.785 ;
        RECT 35.180 45.735 35.550 46.235 ;
        RECT 35.730 45.785 36.135 45.955 ;
        RECT 36.305 45.785 37.090 45.955 ;
        RECT 35.730 45.555 35.900 45.785 ;
        RECT 35.070 45.255 35.900 45.555 ;
        RECT 36.285 45.285 36.750 45.615 ;
        RECT 35.070 45.225 35.270 45.255 ;
        RECT 35.390 45.005 35.560 45.075 ;
        RECT 34.690 44.835 35.560 45.005 ;
        RECT 35.050 44.745 35.560 44.835 ;
        RECT 33.600 44.280 33.905 44.410 ;
        RECT 34.350 44.300 34.880 44.665 ;
        RECT 33.220 43.685 33.485 44.145 ;
        RECT 33.655 43.855 33.905 44.280 ;
        RECT 35.050 44.130 35.220 44.745 ;
        RECT 34.115 43.960 35.220 44.130 ;
        RECT 35.390 43.685 35.560 44.485 ;
        RECT 35.730 44.185 35.900 45.255 ;
        RECT 36.070 44.355 36.260 45.075 ;
        RECT 36.430 44.325 36.750 45.285 ;
        RECT 36.920 45.325 37.090 45.785 ;
        RECT 37.365 45.705 37.575 46.235 ;
        RECT 37.835 45.495 38.165 46.020 ;
        RECT 38.335 45.625 38.505 46.235 ;
        RECT 38.675 45.580 39.005 46.015 ;
        RECT 38.675 45.495 39.055 45.580 ;
        RECT 39.225 45.510 39.515 46.235 ;
        RECT 39.745 45.775 39.990 46.235 ;
        RECT 37.965 45.325 38.165 45.495 ;
        RECT 38.830 45.455 39.055 45.495 ;
        RECT 36.920 44.995 37.795 45.325 ;
        RECT 37.965 44.995 38.715 45.325 ;
        RECT 35.730 43.855 35.980 44.185 ;
        RECT 36.920 44.155 37.090 44.995 ;
        RECT 37.965 44.790 38.155 44.995 ;
        RECT 38.885 44.875 39.055 45.455 ;
        RECT 39.685 44.995 40.000 45.605 ;
        RECT 40.170 45.245 40.420 46.055 ;
        RECT 40.590 45.710 40.850 46.235 ;
        RECT 41.020 45.585 41.280 46.040 ;
        RECT 41.450 45.755 41.710 46.235 ;
        RECT 41.880 45.585 42.140 46.040 ;
        RECT 42.310 45.755 42.570 46.235 ;
        RECT 42.740 45.585 43.000 46.040 ;
        RECT 43.170 45.755 43.430 46.235 ;
        RECT 43.600 45.585 43.860 46.040 ;
        RECT 44.030 45.755 44.330 46.235 ;
        RECT 41.020 45.415 44.330 45.585 ;
        RECT 40.170 44.995 43.190 45.245 ;
        RECT 38.840 44.825 39.055 44.875 ;
        RECT 37.260 44.415 38.155 44.790 ;
        RECT 38.665 44.745 39.055 44.825 ;
        RECT 36.205 43.985 37.090 44.155 ;
        RECT 37.270 43.685 37.585 44.185 ;
        RECT 37.815 43.855 38.155 44.415 ;
        RECT 38.325 43.685 38.495 44.695 ;
        RECT 38.665 43.900 38.995 44.745 ;
        RECT 39.225 43.685 39.515 44.850 ;
        RECT 39.695 43.685 39.990 44.795 ;
        RECT 40.170 43.860 40.420 44.995 ;
        RECT 43.360 44.825 44.330 45.415 ;
        RECT 40.590 43.685 40.850 44.795 ;
        RECT 41.020 44.585 44.330 44.825 ;
        RECT 44.745 45.495 45.130 46.065 ;
        RECT 45.300 45.775 45.625 46.235 ;
        RECT 46.145 45.605 46.425 46.065 ;
        RECT 44.745 44.825 45.025 45.495 ;
        RECT 45.300 45.435 46.425 45.605 ;
        RECT 45.300 45.325 45.750 45.435 ;
        RECT 45.195 44.995 45.750 45.325 ;
        RECT 46.615 45.265 47.015 46.065 ;
        RECT 47.415 45.775 47.685 46.235 ;
        RECT 47.855 45.605 48.140 46.065 ;
        RECT 41.020 43.860 41.280 44.585 ;
        RECT 41.450 43.685 41.710 44.415 ;
        RECT 41.880 43.860 42.140 44.585 ;
        RECT 42.310 43.685 42.570 44.415 ;
        RECT 42.740 43.860 43.000 44.585 ;
        RECT 43.170 43.685 43.430 44.415 ;
        RECT 43.600 43.860 43.860 44.585 ;
        RECT 44.030 43.685 44.325 44.415 ;
        RECT 44.745 43.855 45.130 44.825 ;
        RECT 45.300 44.535 45.750 44.995 ;
        RECT 45.920 44.705 47.015 45.265 ;
        RECT 45.300 44.315 46.425 44.535 ;
        RECT 45.300 43.685 45.625 44.145 ;
        RECT 46.145 43.855 46.425 44.315 ;
        RECT 46.615 43.855 47.015 44.705 ;
        RECT 47.185 45.435 48.140 45.605 ;
        RECT 48.425 45.735 48.725 46.065 ;
        RECT 48.895 45.755 49.170 46.235 ;
        RECT 47.185 44.535 47.395 45.435 ;
        RECT 47.565 44.705 48.255 45.265 ;
        RECT 48.425 44.825 48.595 45.735 ;
        RECT 49.350 45.585 49.645 45.975 ;
        RECT 49.815 45.755 50.070 46.235 ;
        RECT 50.245 45.585 50.505 45.975 ;
        RECT 50.675 45.755 50.955 46.235 ;
        RECT 48.765 44.995 49.115 45.565 ;
        RECT 49.350 45.415 51.000 45.585 ;
        RECT 51.190 45.415 51.465 46.235 ;
        RECT 51.635 45.595 51.965 46.065 ;
        RECT 52.135 45.765 52.305 46.235 ;
        RECT 52.475 45.595 52.805 46.065 ;
        RECT 52.975 45.765 53.685 46.235 ;
        RECT 53.855 45.595 54.185 46.065 ;
        RECT 54.355 45.765 54.645 46.235 ;
        RECT 51.635 45.415 54.695 45.595 ;
        RECT 49.285 45.075 50.425 45.245 ;
        RECT 49.285 44.825 49.455 45.075 ;
        RECT 50.595 44.905 51.000 45.415 ;
        RECT 51.235 45.035 52.065 45.245 ;
        RECT 52.235 45.035 53.285 45.245 ;
        RECT 53.475 45.035 54.065 45.245 ;
        RECT 48.425 44.655 49.455 44.825 ;
        RECT 50.245 44.735 51.000 44.905 ;
        RECT 47.185 44.315 48.140 44.535 ;
        RECT 47.415 43.685 47.685 44.145 ;
        RECT 47.855 43.855 48.140 44.315 ;
        RECT 48.425 43.855 48.735 44.655 ;
        RECT 50.245 44.485 50.505 44.735 ;
        RECT 51.250 44.695 53.185 44.865 ;
        RECT 53.475 44.695 53.740 45.035 ;
        RECT 54.235 44.865 54.695 45.415 ;
        RECT 54.865 45.465 56.535 46.235 ;
        RECT 56.715 45.745 57.045 46.235 ;
        RECT 57.215 45.640 57.835 46.065 ;
        RECT 54.865 44.945 55.615 45.465 ;
        RECT 53.935 44.695 54.695 44.865 ;
        RECT 55.785 44.775 56.535 45.295 ;
        RECT 56.705 44.995 57.045 45.575 ;
        RECT 57.215 45.305 57.575 45.640 ;
        RECT 58.295 45.545 58.625 46.235 ;
        RECT 60.495 45.855 61.665 46.065 ;
        RECT 60.495 45.835 60.825 45.855 ;
        RECT 60.385 45.415 61.245 45.665 ;
        RECT 61.415 45.605 61.665 45.855 ;
        RECT 61.835 45.775 62.005 46.235 ;
        RECT 62.175 45.605 62.515 46.065 ;
        RECT 61.415 45.435 62.515 45.605 ;
        RECT 62.685 45.465 64.355 46.235 ;
        RECT 64.985 45.510 65.275 46.235 ;
        RECT 65.445 45.465 67.115 46.235 ;
        RECT 67.290 45.765 67.620 46.235 ;
        RECT 67.790 45.595 68.015 46.040 ;
        RECT 68.185 45.710 68.480 46.235 ;
        RECT 69.185 45.775 69.430 46.235 ;
        RECT 57.215 45.025 58.635 45.305 ;
        RECT 48.905 43.685 49.215 44.485 ;
        RECT 49.385 44.315 50.505 44.485 ;
        RECT 49.385 43.855 49.645 44.315 ;
        RECT 49.815 43.685 50.070 44.145 ;
        RECT 50.245 43.855 50.505 44.315 ;
        RECT 50.675 43.685 50.960 44.555 ;
        RECT 51.250 43.855 51.505 44.695 ;
        RECT 51.675 43.685 51.925 44.525 ;
        RECT 52.095 43.855 52.345 44.695 ;
        RECT 52.515 44.025 52.765 44.525 ;
        RECT 52.935 44.195 53.185 44.695 ;
        RECT 53.515 44.025 53.725 44.525 ;
        RECT 53.935 44.195 54.145 44.695 ;
        RECT 54.315 44.025 54.565 44.525 ;
        RECT 52.515 43.855 54.565 44.025 ;
        RECT 54.865 43.685 56.535 44.775 ;
        RECT 56.715 43.685 57.045 44.825 ;
        RECT 57.215 43.855 57.575 45.025 ;
        RECT 57.775 43.685 58.105 44.855 ;
        RECT 58.305 43.855 58.635 45.025 ;
        RECT 58.835 43.685 59.165 44.855 ;
        RECT 60.385 44.825 60.665 45.415 ;
        RECT 60.835 44.995 61.585 45.245 ;
        RECT 61.755 44.995 62.515 45.245 ;
        RECT 62.685 44.945 63.435 45.465 ;
        RECT 60.385 44.655 62.085 44.825 ;
        RECT 60.490 43.685 60.745 44.485 ;
        RECT 60.915 43.855 61.245 44.655 ;
        RECT 61.415 43.685 61.585 44.485 ;
        RECT 61.755 43.855 62.085 44.655 ;
        RECT 62.255 43.685 62.515 44.825 ;
        RECT 63.605 44.775 64.355 45.295 ;
        RECT 65.445 44.945 66.195 45.465 ;
        RECT 67.285 45.425 68.015 45.595 ;
        RECT 62.685 43.685 64.355 44.775 ;
        RECT 64.985 43.685 65.275 44.850 ;
        RECT 66.365 44.775 67.115 45.295 ;
        RECT 65.445 43.685 67.115 44.775 ;
        RECT 67.285 44.860 67.565 45.425 ;
        RECT 67.735 45.030 68.955 45.255 ;
        RECT 69.125 44.995 69.440 45.605 ;
        RECT 69.610 45.245 69.860 46.055 ;
        RECT 70.030 45.710 70.290 46.235 ;
        RECT 70.460 45.585 70.720 46.040 ;
        RECT 70.890 45.755 71.150 46.235 ;
        RECT 71.320 45.585 71.580 46.040 ;
        RECT 71.750 45.755 72.010 46.235 ;
        RECT 72.180 45.585 72.440 46.040 ;
        RECT 72.610 45.755 72.870 46.235 ;
        RECT 73.040 45.585 73.300 46.040 ;
        RECT 73.470 45.755 73.770 46.235 ;
        RECT 74.275 45.685 74.445 45.975 ;
        RECT 74.615 45.855 74.945 46.235 ;
        RECT 70.460 45.415 73.770 45.585 ;
        RECT 74.275 45.515 74.940 45.685 ;
        RECT 69.610 44.995 72.630 45.245 ;
        RECT 67.285 44.690 68.885 44.860 ;
        RECT 67.345 43.685 67.600 44.520 ;
        RECT 67.770 43.885 68.030 44.690 ;
        RECT 68.200 43.685 68.460 44.520 ;
        RECT 68.630 43.885 68.885 44.690 ;
        RECT 69.135 43.685 69.430 44.795 ;
        RECT 69.610 43.860 69.860 44.995 ;
        RECT 72.800 44.825 73.770 45.415 ;
        RECT 70.030 43.685 70.290 44.795 ;
        RECT 70.460 44.585 73.770 44.825 ;
        RECT 74.190 44.695 74.540 45.345 ;
        RECT 70.460 43.860 70.720 44.585 ;
        RECT 70.890 43.685 71.150 44.415 ;
        RECT 71.320 43.860 71.580 44.585 ;
        RECT 71.750 43.685 72.010 44.415 ;
        RECT 72.180 43.860 72.440 44.585 ;
        RECT 72.610 43.685 72.870 44.415 ;
        RECT 73.040 43.860 73.300 44.585 ;
        RECT 74.710 44.525 74.940 45.515 ;
        RECT 73.470 43.685 73.765 44.415 ;
        RECT 74.275 44.355 74.940 44.525 ;
        RECT 74.275 43.855 74.445 44.355 ;
        RECT 74.615 43.685 74.945 44.185 ;
        RECT 75.115 43.855 75.300 45.975 ;
        RECT 75.555 45.775 75.805 46.235 ;
        RECT 75.975 45.785 76.310 45.955 ;
        RECT 76.505 45.785 77.180 45.955 ;
        RECT 75.975 45.645 76.145 45.785 ;
        RECT 75.470 44.655 75.750 45.605 ;
        RECT 75.920 45.515 76.145 45.645 ;
        RECT 75.920 44.410 76.090 45.515 ;
        RECT 76.315 45.365 76.840 45.585 ;
        RECT 76.260 44.600 76.500 45.195 ;
        RECT 76.670 44.665 76.840 45.365 ;
        RECT 77.010 45.005 77.180 45.785 ;
        RECT 77.500 45.735 77.870 46.235 ;
        RECT 78.050 45.785 78.455 45.955 ;
        RECT 78.625 45.785 79.410 45.955 ;
        RECT 78.050 45.555 78.220 45.785 ;
        RECT 77.390 45.255 78.220 45.555 ;
        RECT 78.605 45.285 79.070 45.615 ;
        RECT 77.390 45.225 77.590 45.255 ;
        RECT 77.710 45.005 77.880 45.075 ;
        RECT 77.010 44.835 77.880 45.005 ;
        RECT 77.370 44.745 77.880 44.835 ;
        RECT 75.920 44.280 76.225 44.410 ;
        RECT 76.670 44.300 77.200 44.665 ;
        RECT 75.540 43.685 75.805 44.145 ;
        RECT 75.975 43.855 76.225 44.280 ;
        RECT 77.370 44.130 77.540 44.745 ;
        RECT 76.435 43.960 77.540 44.130 ;
        RECT 77.710 43.685 77.880 44.485 ;
        RECT 78.050 44.185 78.220 45.255 ;
        RECT 78.390 44.355 78.580 45.075 ;
        RECT 78.750 44.325 79.070 45.285 ;
        RECT 79.240 45.325 79.410 45.785 ;
        RECT 79.685 45.705 79.895 46.235 ;
        RECT 80.155 45.495 80.485 46.020 ;
        RECT 80.655 45.625 80.825 46.235 ;
        RECT 80.995 45.580 81.325 46.015 ;
        RECT 81.545 45.690 86.890 46.235 ;
        RECT 80.995 45.495 81.375 45.580 ;
        RECT 80.285 45.325 80.485 45.495 ;
        RECT 81.150 45.455 81.375 45.495 ;
        RECT 79.240 44.995 80.115 45.325 ;
        RECT 80.285 44.995 81.035 45.325 ;
        RECT 78.050 43.855 78.300 44.185 ;
        RECT 79.240 44.155 79.410 44.995 ;
        RECT 80.285 44.790 80.475 44.995 ;
        RECT 81.205 44.875 81.375 45.455 ;
        RECT 81.160 44.825 81.375 44.875 ;
        RECT 83.130 44.860 83.470 45.690 ;
        RECT 87.065 45.465 88.735 46.235 ;
        RECT 88.995 45.685 89.165 46.065 ;
        RECT 89.380 45.855 89.710 46.235 ;
        RECT 88.995 45.515 89.710 45.685 ;
        RECT 79.580 44.415 80.475 44.790 ;
        RECT 80.985 44.745 81.375 44.825 ;
        RECT 78.525 43.985 79.410 44.155 ;
        RECT 79.590 43.685 79.905 44.185 ;
        RECT 80.135 43.855 80.475 44.415 ;
        RECT 80.645 43.685 80.815 44.695 ;
        RECT 80.985 43.900 81.315 44.745 ;
        RECT 84.950 44.120 85.300 45.370 ;
        RECT 87.065 44.945 87.815 45.465 ;
        RECT 87.985 44.775 88.735 45.295 ;
        RECT 88.905 44.965 89.260 45.335 ;
        RECT 89.540 45.325 89.710 45.515 ;
        RECT 89.880 45.490 90.135 46.065 ;
        RECT 89.540 44.995 89.795 45.325 ;
        RECT 89.540 44.785 89.710 44.995 ;
        RECT 81.545 43.685 86.890 44.120 ;
        RECT 87.065 43.685 88.735 44.775 ;
        RECT 88.995 44.615 89.710 44.785 ;
        RECT 89.965 44.760 90.135 45.490 ;
        RECT 90.310 45.395 90.570 46.235 ;
        RECT 90.745 45.485 91.955 46.235 ;
        RECT 88.995 43.855 89.165 44.615 ;
        RECT 89.380 43.685 89.710 44.445 ;
        RECT 89.880 43.855 90.135 44.760 ;
        RECT 90.310 43.685 90.570 44.835 ;
        RECT 90.745 44.775 91.265 45.315 ;
        RECT 91.435 44.945 91.955 45.485 ;
        RECT 90.745 43.685 91.955 44.775 ;
        RECT 13.380 43.515 92.040 43.685 ;
        RECT 13.465 42.425 14.675 43.515 ;
        RECT 14.935 42.845 15.105 43.345 ;
        RECT 15.275 43.015 15.605 43.515 ;
        RECT 14.935 42.675 15.600 42.845 ;
        RECT 13.465 41.715 13.985 42.255 ;
        RECT 14.155 41.885 14.675 42.425 ;
        RECT 14.850 41.855 15.200 42.505 ;
        RECT 13.465 40.965 14.675 41.715 ;
        RECT 15.370 41.685 15.600 42.675 ;
        RECT 14.935 41.515 15.600 41.685 ;
        RECT 14.935 41.225 15.105 41.515 ;
        RECT 15.275 40.965 15.605 41.345 ;
        RECT 15.775 41.225 15.960 43.345 ;
        RECT 16.200 43.055 16.465 43.515 ;
        RECT 16.635 42.920 16.885 43.345 ;
        RECT 17.095 43.070 18.200 43.240 ;
        RECT 16.580 42.790 16.885 42.920 ;
        RECT 16.130 41.595 16.410 42.545 ;
        RECT 16.580 41.685 16.750 42.790 ;
        RECT 16.920 42.005 17.160 42.600 ;
        RECT 17.330 42.535 17.860 42.900 ;
        RECT 17.330 41.835 17.500 42.535 ;
        RECT 18.030 42.455 18.200 43.070 ;
        RECT 18.370 42.715 18.540 43.515 ;
        RECT 18.710 43.015 18.960 43.345 ;
        RECT 19.185 43.045 20.070 43.215 ;
        RECT 18.030 42.365 18.540 42.455 ;
        RECT 16.580 41.555 16.805 41.685 ;
        RECT 16.975 41.615 17.500 41.835 ;
        RECT 17.670 42.195 18.540 42.365 ;
        RECT 16.215 40.965 16.465 41.425 ;
        RECT 16.635 41.415 16.805 41.555 ;
        RECT 17.670 41.415 17.840 42.195 ;
        RECT 18.370 42.125 18.540 42.195 ;
        RECT 18.050 41.945 18.250 41.975 ;
        RECT 18.710 41.945 18.880 43.015 ;
        RECT 19.050 42.125 19.240 42.845 ;
        RECT 18.050 41.645 18.880 41.945 ;
        RECT 19.410 41.915 19.730 42.875 ;
        RECT 16.635 41.245 16.970 41.415 ;
        RECT 17.165 41.245 17.840 41.415 ;
        RECT 18.160 40.965 18.530 41.465 ;
        RECT 18.710 41.415 18.880 41.645 ;
        RECT 19.265 41.585 19.730 41.915 ;
        RECT 19.900 42.205 20.070 43.045 ;
        RECT 20.250 43.015 20.565 43.515 ;
        RECT 20.795 42.785 21.135 43.345 ;
        RECT 20.240 42.410 21.135 42.785 ;
        RECT 21.305 42.505 21.475 43.515 ;
        RECT 20.945 42.205 21.135 42.410 ;
        RECT 21.645 42.455 21.975 43.300 ;
        RECT 21.645 42.375 22.035 42.455 ;
        RECT 21.820 42.325 22.035 42.375 ;
        RECT 22.210 42.365 22.470 43.515 ;
        RECT 22.645 42.440 22.900 43.345 ;
        RECT 23.070 42.755 23.400 43.515 ;
        RECT 23.615 42.585 23.785 43.345 ;
        RECT 19.900 41.875 20.775 42.205 ;
        RECT 20.945 41.875 21.695 42.205 ;
        RECT 19.900 41.415 20.070 41.875 ;
        RECT 20.945 41.705 21.145 41.875 ;
        RECT 21.865 41.745 22.035 42.325 ;
        RECT 21.810 41.705 22.035 41.745 ;
        RECT 18.710 41.245 19.115 41.415 ;
        RECT 19.285 41.245 20.070 41.415 ;
        RECT 20.345 40.965 20.555 41.495 ;
        RECT 20.815 41.180 21.145 41.705 ;
        RECT 21.655 41.620 22.035 41.705 ;
        RECT 21.315 40.965 21.485 41.575 ;
        RECT 21.655 41.185 21.985 41.620 ;
        RECT 22.210 40.965 22.470 41.805 ;
        RECT 22.645 41.710 22.815 42.440 ;
        RECT 23.070 42.415 23.785 42.585 ;
        RECT 24.045 42.425 25.715 43.515 ;
        RECT 23.070 42.205 23.240 42.415 ;
        RECT 22.985 41.875 23.240 42.205 ;
        RECT 22.645 41.135 22.900 41.710 ;
        RECT 23.070 41.685 23.240 41.875 ;
        RECT 23.520 41.865 23.875 42.235 ;
        RECT 24.045 41.735 24.795 42.255 ;
        RECT 24.965 41.905 25.715 42.425 ;
        RECT 26.345 42.350 26.635 43.515 ;
        RECT 26.845 42.565 27.135 43.335 ;
        RECT 27.705 42.975 27.965 43.335 ;
        RECT 28.135 43.145 28.465 43.515 ;
        RECT 28.635 42.975 28.895 43.335 ;
        RECT 27.705 42.745 28.895 42.975 ;
        RECT 29.085 42.795 29.415 43.515 ;
        RECT 29.585 42.565 29.850 43.335 ;
        RECT 30.130 43.055 30.300 43.515 ;
        RECT 30.470 42.885 30.800 43.345 ;
        RECT 26.845 42.385 29.340 42.565 ;
        RECT 26.815 41.875 27.085 42.205 ;
        RECT 27.265 41.875 27.700 42.205 ;
        RECT 27.880 41.875 28.455 42.205 ;
        RECT 28.635 41.875 28.915 42.205 ;
        RECT 23.070 41.515 23.785 41.685 ;
        RECT 23.070 40.965 23.400 41.345 ;
        RECT 23.615 41.135 23.785 41.515 ;
        RECT 24.045 40.965 25.715 41.735 ;
        RECT 29.115 41.695 29.340 42.385 ;
        RECT 26.345 40.965 26.635 41.690 ;
        RECT 26.855 41.505 29.340 41.695 ;
        RECT 26.855 41.145 27.080 41.505 ;
        RECT 27.260 40.965 27.590 41.335 ;
        RECT 27.770 41.145 28.025 41.505 ;
        RECT 28.590 40.965 29.335 41.335 ;
        RECT 29.515 41.145 29.850 42.565 ;
        RECT 30.025 42.715 30.800 42.885 ;
        RECT 30.970 42.715 31.140 43.515 ;
        RECT 30.025 41.705 30.455 42.715 ;
        RECT 31.725 42.545 32.085 42.720 ;
        RECT 30.625 42.375 32.085 42.545 ;
        RECT 32.365 42.375 32.595 43.515 ;
        RECT 30.625 41.875 30.795 42.375 ;
        RECT 30.025 41.535 30.720 41.705 ;
        RECT 30.965 41.645 31.375 42.205 ;
        RECT 30.050 40.965 30.380 41.365 ;
        RECT 30.550 41.265 30.720 41.535 ;
        RECT 31.545 41.475 31.725 42.375 ;
        RECT 32.765 42.365 33.095 43.345 ;
        RECT 33.265 42.375 33.475 43.515 ;
        RECT 33.705 43.080 39.050 43.515 ;
        RECT 31.895 42.155 32.090 42.205 ;
        RECT 31.895 41.985 32.095 42.155 ;
        RECT 31.895 41.645 32.090 41.985 ;
        RECT 32.345 41.955 32.675 42.205 ;
        RECT 30.890 40.965 31.205 41.475 ;
        RECT 31.435 41.135 31.725 41.475 ;
        RECT 31.895 40.965 32.135 41.475 ;
        RECT 32.365 40.965 32.595 41.785 ;
        RECT 32.845 41.765 33.095 42.365 ;
        RECT 32.765 41.135 33.095 41.765 ;
        RECT 33.265 40.965 33.475 41.785 ;
        RECT 35.290 41.510 35.630 42.340 ;
        RECT 37.110 41.830 37.460 43.080 ;
        RECT 39.690 42.375 40.025 43.345 ;
        RECT 40.195 42.375 40.365 43.515 ;
        RECT 40.535 43.175 42.565 43.345 ;
        RECT 39.690 41.705 39.860 42.375 ;
        RECT 40.535 42.205 40.705 43.175 ;
        RECT 40.030 41.875 40.285 42.205 ;
        RECT 40.510 41.875 40.705 42.205 ;
        RECT 40.875 42.835 42.000 43.005 ;
        RECT 40.115 41.705 40.285 41.875 ;
        RECT 40.875 41.705 41.045 42.835 ;
        RECT 33.705 40.965 39.050 41.510 ;
        RECT 39.690 41.135 39.945 41.705 ;
        RECT 40.115 41.535 41.045 41.705 ;
        RECT 41.215 42.495 42.225 42.665 ;
        RECT 41.215 41.695 41.385 42.495 ;
        RECT 41.590 42.155 41.865 42.295 ;
        RECT 41.585 41.985 41.865 42.155 ;
        RECT 40.870 41.500 41.045 41.535 ;
        RECT 40.115 40.965 40.445 41.365 ;
        RECT 40.870 41.135 41.400 41.500 ;
        RECT 41.590 41.135 41.865 41.985 ;
        RECT 42.035 41.135 42.225 42.495 ;
        RECT 42.395 42.510 42.565 43.175 ;
        RECT 42.735 42.755 42.905 43.515 ;
        RECT 43.140 42.755 43.655 43.165 ;
        RECT 42.395 42.320 43.145 42.510 ;
        RECT 43.315 41.945 43.655 42.755 ;
        RECT 44.835 42.845 45.005 43.345 ;
        RECT 45.175 43.015 45.505 43.515 ;
        RECT 44.835 42.675 45.500 42.845 ;
        RECT 42.425 41.775 43.655 41.945 ;
        RECT 44.750 41.855 45.100 42.505 ;
        RECT 42.405 40.965 42.915 41.500 ;
        RECT 43.135 41.170 43.380 41.775 ;
        RECT 45.270 41.685 45.500 42.675 ;
        RECT 44.835 41.515 45.500 41.685 ;
        RECT 44.835 41.225 45.005 41.515 ;
        RECT 45.175 40.965 45.505 41.345 ;
        RECT 45.675 41.225 45.860 43.345 ;
        RECT 46.100 43.055 46.365 43.515 ;
        RECT 46.535 42.920 46.785 43.345 ;
        RECT 46.995 43.070 48.100 43.240 ;
        RECT 46.480 42.790 46.785 42.920 ;
        RECT 46.030 41.595 46.310 42.545 ;
        RECT 46.480 41.685 46.650 42.790 ;
        RECT 46.820 42.005 47.060 42.600 ;
        RECT 47.230 42.535 47.760 42.900 ;
        RECT 47.230 41.835 47.400 42.535 ;
        RECT 47.930 42.455 48.100 43.070 ;
        RECT 48.270 42.715 48.440 43.515 ;
        RECT 48.610 43.015 48.860 43.345 ;
        RECT 49.085 43.045 49.970 43.215 ;
        RECT 47.930 42.365 48.440 42.455 ;
        RECT 46.480 41.555 46.705 41.685 ;
        RECT 46.875 41.615 47.400 41.835 ;
        RECT 47.570 42.195 48.440 42.365 ;
        RECT 46.115 40.965 46.365 41.425 ;
        RECT 46.535 41.415 46.705 41.555 ;
        RECT 47.570 41.415 47.740 42.195 ;
        RECT 48.270 42.125 48.440 42.195 ;
        RECT 47.950 41.945 48.150 41.975 ;
        RECT 48.610 41.945 48.780 43.015 ;
        RECT 48.950 42.125 49.140 42.845 ;
        RECT 47.950 41.645 48.780 41.945 ;
        RECT 49.310 41.915 49.630 42.875 ;
        RECT 46.535 41.245 46.870 41.415 ;
        RECT 47.065 41.245 47.740 41.415 ;
        RECT 48.060 40.965 48.430 41.465 ;
        RECT 48.610 41.415 48.780 41.645 ;
        RECT 49.165 41.585 49.630 41.915 ;
        RECT 49.800 42.205 49.970 43.045 ;
        RECT 50.150 43.015 50.465 43.515 ;
        RECT 50.695 42.785 51.035 43.345 ;
        RECT 50.140 42.410 51.035 42.785 ;
        RECT 51.205 42.505 51.375 43.515 ;
        RECT 50.845 42.205 51.035 42.410 ;
        RECT 51.545 42.455 51.875 43.300 ;
        RECT 51.545 42.375 51.935 42.455 ;
        RECT 51.720 42.325 51.935 42.375 ;
        RECT 52.105 42.350 52.395 43.515 ;
        RECT 52.605 42.375 52.835 43.515 ;
        RECT 53.005 42.365 53.335 43.345 ;
        RECT 53.505 42.375 53.715 43.515 ;
        RECT 54.035 42.845 54.205 43.345 ;
        RECT 54.375 43.015 54.705 43.515 ;
        RECT 54.035 42.675 54.700 42.845 ;
        RECT 49.800 41.875 50.675 42.205 ;
        RECT 50.845 41.875 51.595 42.205 ;
        RECT 49.800 41.415 49.970 41.875 ;
        RECT 50.845 41.705 51.045 41.875 ;
        RECT 51.765 41.745 51.935 42.325 ;
        RECT 52.585 41.955 52.915 42.205 ;
        RECT 51.710 41.705 51.935 41.745 ;
        RECT 48.610 41.245 49.015 41.415 ;
        RECT 49.185 41.245 49.970 41.415 ;
        RECT 50.245 40.965 50.455 41.495 ;
        RECT 50.715 41.180 51.045 41.705 ;
        RECT 51.555 41.620 51.935 41.705 ;
        RECT 51.215 40.965 51.385 41.575 ;
        RECT 51.555 41.185 51.885 41.620 ;
        RECT 52.105 40.965 52.395 41.690 ;
        RECT 52.605 40.965 52.835 41.785 ;
        RECT 53.085 41.765 53.335 42.365 ;
        RECT 53.950 41.855 54.300 42.505 ;
        RECT 53.005 41.135 53.335 41.765 ;
        RECT 53.505 40.965 53.715 41.785 ;
        RECT 54.470 41.685 54.700 42.675 ;
        RECT 54.035 41.515 54.700 41.685 ;
        RECT 54.035 41.225 54.205 41.515 ;
        RECT 54.375 40.965 54.705 41.345 ;
        RECT 54.875 41.225 55.060 43.345 ;
        RECT 55.300 43.055 55.565 43.515 ;
        RECT 55.735 42.920 55.985 43.345 ;
        RECT 56.195 43.070 57.300 43.240 ;
        RECT 55.680 42.790 55.985 42.920 ;
        RECT 55.230 41.595 55.510 42.545 ;
        RECT 55.680 41.685 55.850 42.790 ;
        RECT 56.020 42.005 56.260 42.600 ;
        RECT 56.430 42.535 56.960 42.900 ;
        RECT 56.430 41.835 56.600 42.535 ;
        RECT 57.130 42.455 57.300 43.070 ;
        RECT 57.470 42.715 57.640 43.515 ;
        RECT 57.810 43.015 58.060 43.345 ;
        RECT 58.285 43.045 59.170 43.215 ;
        RECT 57.130 42.365 57.640 42.455 ;
        RECT 55.680 41.555 55.905 41.685 ;
        RECT 56.075 41.615 56.600 41.835 ;
        RECT 56.770 42.195 57.640 42.365 ;
        RECT 55.315 40.965 55.565 41.425 ;
        RECT 55.735 41.415 55.905 41.555 ;
        RECT 56.770 41.415 56.940 42.195 ;
        RECT 57.470 42.125 57.640 42.195 ;
        RECT 57.150 41.945 57.350 41.975 ;
        RECT 57.810 41.945 57.980 43.015 ;
        RECT 58.150 42.125 58.340 42.845 ;
        RECT 57.150 41.645 57.980 41.945 ;
        RECT 58.510 41.915 58.830 42.875 ;
        RECT 55.735 41.245 56.070 41.415 ;
        RECT 56.265 41.245 56.940 41.415 ;
        RECT 57.260 40.965 57.630 41.465 ;
        RECT 57.810 41.415 57.980 41.645 ;
        RECT 58.365 41.585 58.830 41.915 ;
        RECT 59.000 42.205 59.170 43.045 ;
        RECT 59.350 43.015 59.665 43.515 ;
        RECT 59.895 42.785 60.235 43.345 ;
        RECT 59.340 42.410 60.235 42.785 ;
        RECT 60.405 42.505 60.575 43.515 ;
        RECT 60.045 42.205 60.235 42.410 ;
        RECT 60.745 42.455 61.075 43.300 ;
        RECT 62.315 42.845 62.485 43.345 ;
        RECT 62.655 43.015 62.985 43.515 ;
        RECT 62.315 42.675 62.980 42.845 ;
        RECT 60.745 42.375 61.135 42.455 ;
        RECT 60.920 42.325 61.135 42.375 ;
        RECT 59.000 41.875 59.875 42.205 ;
        RECT 60.045 41.875 60.795 42.205 ;
        RECT 59.000 41.415 59.170 41.875 ;
        RECT 60.045 41.705 60.245 41.875 ;
        RECT 60.965 41.745 61.135 42.325 ;
        RECT 62.230 41.855 62.580 42.505 ;
        RECT 60.910 41.705 61.135 41.745 ;
        RECT 57.810 41.245 58.215 41.415 ;
        RECT 58.385 41.245 59.170 41.415 ;
        RECT 59.445 40.965 59.655 41.495 ;
        RECT 59.915 41.180 60.245 41.705 ;
        RECT 60.755 41.620 61.135 41.705 ;
        RECT 62.750 41.685 62.980 42.675 ;
        RECT 60.415 40.965 60.585 41.575 ;
        RECT 60.755 41.185 61.085 41.620 ;
        RECT 62.315 41.515 62.980 41.685 ;
        RECT 62.315 41.225 62.485 41.515 ;
        RECT 62.655 40.965 62.985 41.345 ;
        RECT 63.155 41.225 63.340 43.345 ;
        RECT 63.580 43.055 63.845 43.515 ;
        RECT 64.015 42.920 64.265 43.345 ;
        RECT 64.475 43.070 65.580 43.240 ;
        RECT 63.960 42.790 64.265 42.920 ;
        RECT 63.510 41.595 63.790 42.545 ;
        RECT 63.960 41.685 64.130 42.790 ;
        RECT 64.300 42.005 64.540 42.600 ;
        RECT 64.710 42.535 65.240 42.900 ;
        RECT 64.710 41.835 64.880 42.535 ;
        RECT 65.410 42.455 65.580 43.070 ;
        RECT 65.750 42.715 65.920 43.515 ;
        RECT 66.090 43.015 66.340 43.345 ;
        RECT 66.565 43.045 67.450 43.215 ;
        RECT 65.410 42.365 65.920 42.455 ;
        RECT 63.960 41.555 64.185 41.685 ;
        RECT 64.355 41.615 64.880 41.835 ;
        RECT 65.050 42.195 65.920 42.365 ;
        RECT 63.595 40.965 63.845 41.425 ;
        RECT 64.015 41.415 64.185 41.555 ;
        RECT 65.050 41.415 65.220 42.195 ;
        RECT 65.750 42.125 65.920 42.195 ;
        RECT 65.430 41.945 65.630 41.975 ;
        RECT 66.090 41.945 66.260 43.015 ;
        RECT 66.430 42.125 66.620 42.845 ;
        RECT 65.430 41.645 66.260 41.945 ;
        RECT 66.790 41.915 67.110 42.875 ;
        RECT 64.015 41.245 64.350 41.415 ;
        RECT 64.545 41.245 65.220 41.415 ;
        RECT 65.540 40.965 65.910 41.465 ;
        RECT 66.090 41.415 66.260 41.645 ;
        RECT 66.645 41.585 67.110 41.915 ;
        RECT 67.280 42.205 67.450 43.045 ;
        RECT 67.630 43.015 67.945 43.515 ;
        RECT 68.175 42.785 68.515 43.345 ;
        RECT 67.620 42.410 68.515 42.785 ;
        RECT 68.685 42.505 68.855 43.515 ;
        RECT 68.325 42.205 68.515 42.410 ;
        RECT 69.025 42.455 69.355 43.300 ;
        RECT 70.710 42.545 71.040 43.345 ;
        RECT 71.210 42.715 71.540 43.515 ;
        RECT 71.840 42.545 72.170 43.345 ;
        RECT 72.815 42.715 73.065 43.515 ;
        RECT 69.025 42.375 69.415 42.455 ;
        RECT 70.710 42.375 73.145 42.545 ;
        RECT 73.335 42.375 73.505 43.515 ;
        RECT 73.675 42.375 74.015 43.345 ;
        RECT 74.370 42.545 74.760 42.720 ;
        RECT 75.245 42.715 75.575 43.515 ;
        RECT 75.745 42.725 76.280 43.345 ;
        RECT 74.370 42.375 75.795 42.545 ;
        RECT 69.200 42.325 69.415 42.375 ;
        RECT 67.280 41.875 68.155 42.205 ;
        RECT 68.325 41.875 69.075 42.205 ;
        RECT 67.280 41.415 67.450 41.875 ;
        RECT 68.325 41.705 68.525 41.875 ;
        RECT 69.245 41.745 69.415 42.325 ;
        RECT 70.505 41.955 70.855 42.205 ;
        RECT 71.040 41.745 71.210 42.375 ;
        RECT 71.380 41.955 71.710 42.155 ;
        RECT 71.880 41.955 72.210 42.155 ;
        RECT 72.380 41.955 72.800 42.155 ;
        RECT 72.975 42.125 73.145 42.375 ;
        RECT 72.975 41.955 73.670 42.125 ;
        RECT 69.190 41.705 69.415 41.745 ;
        RECT 66.090 41.245 66.495 41.415 ;
        RECT 66.665 41.245 67.450 41.415 ;
        RECT 67.725 40.965 67.935 41.495 ;
        RECT 68.195 41.180 68.525 41.705 ;
        RECT 69.035 41.620 69.415 41.705 ;
        RECT 68.695 40.965 68.865 41.575 ;
        RECT 69.035 41.185 69.365 41.620 ;
        RECT 70.710 41.135 71.210 41.745 ;
        RECT 71.840 41.615 73.065 41.785 ;
        RECT 73.840 41.765 74.015 42.375 ;
        RECT 71.840 41.135 72.170 41.615 ;
        RECT 72.340 40.965 72.565 41.425 ;
        RECT 72.735 41.135 73.065 41.615 ;
        RECT 73.255 40.965 73.505 41.765 ;
        RECT 73.675 41.135 74.015 41.765 ;
        RECT 74.245 41.645 74.600 42.205 ;
        RECT 74.770 41.475 74.940 42.375 ;
        RECT 75.110 41.645 75.375 42.205 ;
        RECT 75.625 41.875 75.795 42.375 ;
        RECT 75.965 41.705 76.280 42.725 ;
        RECT 76.485 42.425 77.695 43.515 ;
        RECT 74.350 40.965 74.590 41.475 ;
        RECT 74.770 41.145 75.050 41.475 ;
        RECT 75.280 40.965 75.495 41.475 ;
        RECT 75.665 41.135 76.280 41.705 ;
        RECT 76.485 41.715 77.005 42.255 ;
        RECT 77.175 41.885 77.695 42.425 ;
        RECT 77.865 42.350 78.155 43.515 ;
        RECT 78.415 42.845 78.585 43.345 ;
        RECT 78.755 43.015 79.085 43.515 ;
        RECT 78.415 42.675 79.080 42.845 ;
        RECT 78.330 41.855 78.680 42.505 ;
        RECT 76.485 40.965 77.695 41.715 ;
        RECT 77.865 40.965 78.155 41.690 ;
        RECT 78.850 41.685 79.080 42.675 ;
        RECT 78.415 41.515 79.080 41.685 ;
        RECT 78.415 41.225 78.585 41.515 ;
        RECT 78.755 40.965 79.085 41.345 ;
        RECT 79.255 41.225 79.440 43.345 ;
        RECT 79.680 43.055 79.945 43.515 ;
        RECT 80.115 42.920 80.365 43.345 ;
        RECT 80.575 43.070 81.680 43.240 ;
        RECT 80.060 42.790 80.365 42.920 ;
        RECT 79.610 41.595 79.890 42.545 ;
        RECT 80.060 41.685 80.230 42.790 ;
        RECT 80.400 42.005 80.640 42.600 ;
        RECT 80.810 42.535 81.340 42.900 ;
        RECT 80.810 41.835 80.980 42.535 ;
        RECT 81.510 42.455 81.680 43.070 ;
        RECT 81.850 42.715 82.020 43.515 ;
        RECT 82.190 43.015 82.440 43.345 ;
        RECT 82.665 43.045 83.550 43.215 ;
        RECT 81.510 42.365 82.020 42.455 ;
        RECT 80.060 41.555 80.285 41.685 ;
        RECT 80.455 41.615 80.980 41.835 ;
        RECT 81.150 42.195 82.020 42.365 ;
        RECT 79.695 40.965 79.945 41.425 ;
        RECT 80.115 41.415 80.285 41.555 ;
        RECT 81.150 41.415 81.320 42.195 ;
        RECT 81.850 42.125 82.020 42.195 ;
        RECT 81.530 41.945 81.730 41.975 ;
        RECT 82.190 41.945 82.360 43.015 ;
        RECT 82.530 42.125 82.720 42.845 ;
        RECT 81.530 41.645 82.360 41.945 ;
        RECT 82.890 41.915 83.210 42.875 ;
        RECT 80.115 41.245 80.450 41.415 ;
        RECT 80.645 41.245 81.320 41.415 ;
        RECT 81.640 40.965 82.010 41.465 ;
        RECT 82.190 41.415 82.360 41.645 ;
        RECT 82.745 41.585 83.210 41.915 ;
        RECT 83.380 42.205 83.550 43.045 ;
        RECT 83.730 43.015 84.045 43.515 ;
        RECT 84.275 42.785 84.615 43.345 ;
        RECT 83.720 42.410 84.615 42.785 ;
        RECT 84.785 42.505 84.955 43.515 ;
        RECT 84.425 42.205 84.615 42.410 ;
        RECT 85.125 42.455 85.455 43.300 ;
        RECT 85.125 42.375 85.515 42.455 ;
        RECT 85.685 42.425 89.195 43.515 ;
        RECT 89.365 42.425 90.575 43.515 ;
        RECT 85.300 42.325 85.515 42.375 ;
        RECT 83.380 41.875 84.255 42.205 ;
        RECT 84.425 41.875 85.175 42.205 ;
        RECT 83.380 41.415 83.550 41.875 ;
        RECT 84.425 41.705 84.625 41.875 ;
        RECT 85.345 41.745 85.515 42.325 ;
        RECT 85.290 41.705 85.515 41.745 ;
        RECT 82.190 41.245 82.595 41.415 ;
        RECT 82.765 41.245 83.550 41.415 ;
        RECT 83.825 40.965 84.035 41.495 ;
        RECT 84.295 41.180 84.625 41.705 ;
        RECT 85.135 41.620 85.515 41.705 ;
        RECT 85.685 41.735 87.335 42.255 ;
        RECT 87.505 41.905 89.195 42.425 ;
        RECT 84.795 40.965 84.965 41.575 ;
        RECT 85.135 41.185 85.465 41.620 ;
        RECT 85.685 40.965 89.195 41.735 ;
        RECT 89.365 41.715 89.885 42.255 ;
        RECT 90.055 41.885 90.575 42.425 ;
        RECT 90.745 42.425 91.955 43.515 ;
        RECT 90.745 41.885 91.265 42.425 ;
        RECT 91.435 41.715 91.955 42.255 ;
        RECT 89.365 40.965 90.575 41.715 ;
        RECT 90.745 40.965 91.955 41.715 ;
        RECT 13.380 40.795 92.040 40.965 ;
        RECT 13.465 40.045 14.675 40.795 ;
        RECT 13.465 39.505 13.985 40.045 ;
        RECT 15.765 39.995 16.105 40.625 ;
        RECT 16.275 39.995 16.525 40.795 ;
        RECT 16.715 40.145 17.045 40.625 ;
        RECT 17.215 40.335 17.440 40.795 ;
        RECT 17.610 40.145 17.940 40.625 ;
        RECT 14.155 39.335 14.675 39.875 ;
        RECT 13.465 38.245 14.675 39.335 ;
        RECT 15.765 39.385 15.940 39.995 ;
        RECT 16.715 39.975 17.940 40.145 ;
        RECT 18.570 40.015 19.070 40.625 ;
        RECT 19.480 40.055 20.095 40.625 ;
        RECT 20.265 40.285 20.480 40.795 ;
        RECT 20.710 40.285 20.990 40.615 ;
        RECT 21.170 40.285 21.410 40.795 ;
        RECT 16.110 39.635 16.805 39.805 ;
        RECT 16.635 39.385 16.805 39.635 ;
        RECT 16.980 39.605 17.400 39.805 ;
        RECT 17.570 39.605 17.900 39.805 ;
        RECT 18.070 39.605 18.400 39.805 ;
        RECT 18.570 39.385 18.740 40.015 ;
        RECT 18.925 39.555 19.275 39.805 ;
        RECT 15.765 38.415 16.105 39.385 ;
        RECT 16.275 38.245 16.445 39.385 ;
        RECT 16.635 39.215 19.070 39.385 ;
        RECT 16.715 38.245 16.965 39.045 ;
        RECT 17.610 38.415 17.940 39.215 ;
        RECT 18.240 38.245 18.570 39.045 ;
        RECT 18.740 38.415 19.070 39.215 ;
        RECT 19.480 39.035 19.795 40.055 ;
        RECT 19.965 39.385 20.135 39.885 ;
        RECT 20.385 39.555 20.650 40.115 ;
        RECT 20.820 39.385 20.990 40.285 ;
        RECT 21.160 39.555 21.515 40.115 ;
        RECT 21.750 40.030 22.205 40.795 ;
        RECT 22.480 40.415 23.780 40.625 ;
        RECT 24.035 40.435 24.365 40.795 ;
        RECT 23.610 40.265 23.780 40.415 ;
        RECT 24.535 40.295 24.795 40.625 ;
        RECT 24.565 40.285 24.795 40.295 ;
        RECT 22.680 39.805 22.900 40.205 ;
        RECT 21.745 39.605 22.235 39.805 ;
        RECT 22.425 39.595 22.900 39.805 ;
        RECT 23.145 39.805 23.355 40.205 ;
        RECT 23.610 40.140 24.365 40.265 ;
        RECT 23.610 40.095 24.455 40.140 ;
        RECT 24.185 39.975 24.455 40.095 ;
        RECT 23.145 39.595 23.475 39.805 ;
        RECT 23.645 39.535 24.055 39.840 ;
        RECT 19.965 39.215 21.390 39.385 ;
        RECT 19.480 38.415 20.015 39.035 ;
        RECT 20.185 38.245 20.515 39.045 ;
        RECT 21.000 39.040 21.390 39.215 ;
        RECT 21.750 39.365 22.925 39.425 ;
        RECT 24.285 39.400 24.455 39.975 ;
        RECT 24.255 39.365 24.455 39.400 ;
        RECT 21.750 39.255 24.455 39.365 ;
        RECT 21.750 38.635 22.005 39.255 ;
        RECT 22.595 39.195 24.395 39.255 ;
        RECT 22.595 39.165 22.925 39.195 ;
        RECT 24.625 39.095 24.795 40.285 ;
        RECT 24.965 40.025 28.475 40.795 ;
        RECT 24.965 39.505 26.615 40.025 ;
        RECT 29.125 39.985 29.365 40.795 ;
        RECT 29.535 39.985 29.865 40.625 ;
        RECT 30.035 39.985 30.305 40.795 ;
        RECT 30.485 40.045 31.695 40.795 ;
        RECT 31.865 40.335 32.425 40.625 ;
        RECT 32.595 40.335 32.845 40.795 ;
        RECT 26.785 39.335 28.475 39.855 ;
        RECT 29.105 39.555 29.455 39.805 ;
        RECT 29.625 39.385 29.795 39.985 ;
        RECT 29.965 39.555 30.315 39.805 ;
        RECT 30.485 39.505 31.005 40.045 ;
        RECT 22.255 38.995 22.440 39.085 ;
        RECT 23.030 38.995 23.865 39.005 ;
        RECT 22.255 38.795 23.865 38.995 ;
        RECT 22.255 38.755 22.485 38.795 ;
        RECT 21.750 38.415 22.085 38.635 ;
        RECT 23.090 38.245 23.445 38.625 ;
        RECT 23.615 38.415 23.865 38.795 ;
        RECT 24.115 38.245 24.365 39.025 ;
        RECT 24.535 38.415 24.795 39.095 ;
        RECT 24.965 38.245 28.475 39.335 ;
        RECT 29.115 39.215 29.795 39.385 ;
        RECT 29.115 38.430 29.445 39.215 ;
        RECT 29.975 38.245 30.305 39.385 ;
        RECT 31.175 39.335 31.695 39.875 ;
        RECT 30.485 38.245 31.695 39.335 ;
        RECT 31.865 38.965 32.115 40.335 ;
        RECT 33.465 40.165 33.795 40.525 ;
        RECT 32.405 39.975 33.795 40.165 ;
        RECT 34.165 40.025 37.675 40.795 ;
        RECT 37.845 40.045 39.055 40.795 ;
        RECT 39.225 40.070 39.515 40.795 ;
        RECT 32.405 39.885 32.575 39.975 ;
        RECT 32.285 39.555 32.575 39.885 ;
        RECT 32.745 39.555 33.085 39.805 ;
        RECT 33.305 39.555 33.980 39.805 ;
        RECT 32.405 39.305 32.575 39.555 ;
        RECT 32.405 39.135 33.345 39.305 ;
        RECT 33.715 39.195 33.980 39.555 ;
        RECT 34.165 39.505 35.815 40.025 ;
        RECT 35.985 39.335 37.675 39.855 ;
        RECT 37.845 39.505 38.365 40.045 ;
        RECT 39.685 40.025 41.355 40.795 ;
        RECT 38.535 39.335 39.055 39.875 ;
        RECT 39.685 39.505 40.435 40.025 ;
        RECT 31.865 38.415 32.325 38.965 ;
        RECT 32.515 38.245 32.845 38.965 ;
        RECT 33.045 38.585 33.345 39.135 ;
        RECT 33.515 38.245 33.795 38.915 ;
        RECT 34.165 38.245 37.675 39.335 ;
        RECT 37.845 38.245 39.055 39.335 ;
        RECT 39.225 38.245 39.515 39.410 ;
        RECT 40.605 39.335 41.355 39.855 ;
        RECT 39.685 38.245 41.355 39.335 ;
        RECT 41.530 39.195 41.865 40.615 ;
        RECT 42.045 40.425 42.790 40.795 ;
        RECT 43.355 40.255 43.610 40.615 ;
        RECT 43.790 40.425 44.120 40.795 ;
        RECT 44.300 40.255 44.525 40.615 ;
        RECT 42.040 40.065 44.525 40.255 ;
        RECT 42.040 39.375 42.265 40.065 ;
        RECT 44.745 40.025 47.335 40.795 ;
        RECT 47.970 40.055 48.225 40.625 ;
        RECT 48.395 40.395 48.725 40.795 ;
        RECT 49.150 40.260 49.680 40.625 ;
        RECT 49.870 40.455 50.145 40.625 ;
        RECT 49.865 40.285 50.145 40.455 ;
        RECT 49.150 40.225 49.325 40.260 ;
        RECT 48.395 40.055 49.325 40.225 ;
        RECT 42.465 39.555 42.745 39.885 ;
        RECT 42.925 39.555 43.500 39.885 ;
        RECT 43.680 39.555 44.115 39.885 ;
        RECT 44.295 39.555 44.565 39.885 ;
        RECT 44.745 39.505 45.955 40.025 ;
        RECT 42.040 39.195 44.535 39.375 ;
        RECT 46.125 39.335 47.335 39.855 ;
        RECT 41.530 38.425 41.795 39.195 ;
        RECT 41.965 38.245 42.295 38.965 ;
        RECT 42.485 38.785 43.675 39.015 ;
        RECT 42.485 38.425 42.745 38.785 ;
        RECT 42.915 38.245 43.245 38.615 ;
        RECT 43.415 38.425 43.675 38.785 ;
        RECT 44.245 38.425 44.535 39.195 ;
        RECT 44.745 38.245 47.335 39.335 ;
        RECT 47.970 39.385 48.140 40.055 ;
        RECT 48.395 39.885 48.565 40.055 ;
        RECT 48.310 39.555 48.565 39.885 ;
        RECT 48.790 39.555 48.985 39.885 ;
        RECT 47.970 38.415 48.305 39.385 ;
        RECT 48.475 38.245 48.645 39.385 ;
        RECT 48.815 38.585 48.985 39.555 ;
        RECT 49.155 38.925 49.325 40.055 ;
        RECT 49.495 39.265 49.665 40.065 ;
        RECT 49.870 39.465 50.145 40.285 ;
        RECT 50.315 39.265 50.505 40.625 ;
        RECT 50.685 40.260 51.195 40.795 ;
        RECT 51.415 39.985 51.660 40.590 ;
        RECT 52.105 40.135 52.380 40.795 ;
        RECT 52.550 40.165 52.800 40.625 ;
        RECT 52.975 40.300 53.305 40.795 ;
        RECT 50.705 39.815 51.935 39.985 ;
        RECT 52.550 39.955 52.720 40.165 ;
        RECT 53.485 40.130 53.715 40.575 ;
        RECT 49.495 39.095 50.505 39.265 ;
        RECT 50.675 39.250 51.425 39.440 ;
        RECT 49.155 38.755 50.280 38.925 ;
        RECT 50.675 38.585 50.845 39.250 ;
        RECT 51.595 39.005 51.935 39.815 ;
        RECT 52.105 39.435 52.720 39.955 ;
        RECT 52.890 39.455 53.120 39.885 ;
        RECT 53.305 39.635 53.715 40.130 ;
        RECT 53.885 40.310 54.675 40.575 ;
        RECT 53.885 39.455 54.140 40.310 ;
        RECT 54.310 39.635 54.695 40.115 ;
        RECT 55.385 39.975 55.595 40.795 ;
        RECT 55.765 39.995 56.095 40.625 ;
        RECT 48.815 38.415 50.845 38.585 ;
        RECT 51.015 38.245 51.185 39.005 ;
        RECT 51.420 38.595 51.935 39.005 ;
        RECT 52.105 38.245 52.365 39.255 ;
        RECT 52.535 39.085 52.705 39.435 ;
        RECT 52.890 39.285 54.680 39.455 ;
        RECT 55.765 39.395 56.015 39.995 ;
        RECT 56.265 39.975 56.495 40.795 ;
        RECT 56.950 40.315 57.250 40.795 ;
        RECT 57.420 40.145 57.680 40.600 ;
        RECT 57.850 40.315 58.110 40.795 ;
        RECT 58.280 40.145 58.540 40.600 ;
        RECT 58.710 40.315 58.970 40.795 ;
        RECT 59.140 40.145 59.400 40.600 ;
        RECT 59.570 40.315 59.830 40.795 ;
        RECT 60.000 40.145 60.260 40.600 ;
        RECT 60.430 40.270 60.690 40.795 ;
        RECT 56.950 39.975 60.260 40.145 ;
        RECT 56.185 39.555 56.515 39.805 ;
        RECT 52.535 38.415 52.810 39.085 ;
        RECT 53.010 38.245 53.225 39.090 ;
        RECT 53.450 38.990 53.700 39.285 ;
        RECT 53.925 38.925 54.255 39.115 ;
        RECT 53.410 38.415 53.885 38.755 ;
        RECT 54.065 38.750 54.255 38.925 ;
        RECT 54.425 38.920 54.680 39.285 ;
        RECT 54.065 38.245 54.695 38.750 ;
        RECT 55.385 38.245 55.595 39.385 ;
        RECT 55.765 38.415 56.095 39.395 ;
        RECT 56.950 39.385 57.920 39.975 ;
        RECT 60.860 39.805 61.110 40.615 ;
        RECT 61.290 40.335 61.535 40.795 ;
        RECT 61.965 40.165 62.295 40.525 ;
        RECT 62.925 40.335 63.175 40.795 ;
        RECT 63.345 40.335 63.895 40.625 ;
        RECT 58.090 39.555 61.110 39.805 ;
        RECT 61.280 39.555 61.595 40.165 ;
        RECT 61.965 39.975 63.355 40.165 ;
        RECT 63.185 39.885 63.355 39.975 ;
        RECT 61.765 39.555 62.455 39.805 ;
        RECT 62.685 39.555 63.015 39.805 ;
        RECT 63.185 39.555 63.475 39.885 ;
        RECT 56.265 38.245 56.495 39.385 ;
        RECT 56.950 39.145 60.260 39.385 ;
        RECT 56.955 38.245 57.250 38.975 ;
        RECT 57.420 38.420 57.680 39.145 ;
        RECT 57.850 38.245 58.110 38.975 ;
        RECT 58.280 38.420 58.540 39.145 ;
        RECT 58.710 38.245 58.970 38.975 ;
        RECT 59.140 38.420 59.400 39.145 ;
        RECT 59.570 38.245 59.830 38.975 ;
        RECT 60.000 38.420 60.260 39.145 ;
        RECT 60.430 38.245 60.690 39.355 ;
        RECT 60.860 38.420 61.110 39.555 ;
        RECT 61.290 38.245 61.585 39.355 ;
        RECT 61.765 39.115 62.080 39.555 ;
        RECT 63.185 39.305 63.355 39.555 ;
        RECT 62.415 39.135 63.355 39.305 ;
        RECT 61.965 38.245 62.245 38.915 ;
        RECT 62.415 38.585 62.715 39.135 ;
        RECT 63.645 38.965 63.895 40.335 ;
        RECT 64.065 39.995 64.355 40.795 ;
        RECT 64.985 40.070 65.275 40.795 ;
        RECT 65.445 39.995 65.785 40.625 ;
        RECT 65.955 39.995 66.205 40.795 ;
        RECT 66.395 40.145 66.725 40.625 ;
        RECT 66.895 40.335 67.120 40.795 ;
        RECT 67.290 40.145 67.620 40.625 ;
        RECT 62.925 38.245 63.255 38.965 ;
        RECT 63.445 38.415 63.895 38.965 ;
        RECT 64.065 38.245 64.355 39.385 ;
        RECT 64.985 38.245 65.275 39.410 ;
        RECT 65.445 39.385 65.620 39.995 ;
        RECT 66.395 39.975 67.620 40.145 ;
        RECT 68.250 40.015 68.750 40.625 ;
        RECT 69.750 40.285 69.990 40.795 ;
        RECT 70.170 40.285 70.450 40.615 ;
        RECT 70.680 40.285 70.895 40.795 ;
        RECT 65.790 39.635 66.485 39.805 ;
        RECT 66.315 39.385 66.485 39.635 ;
        RECT 66.660 39.605 67.080 39.805 ;
        RECT 67.250 39.605 67.580 39.805 ;
        RECT 67.750 39.605 68.080 39.805 ;
        RECT 68.250 39.385 68.420 40.015 ;
        RECT 68.605 39.555 68.955 39.805 ;
        RECT 69.645 39.555 70.000 40.115 ;
        RECT 70.170 39.385 70.340 40.285 ;
        RECT 70.510 39.555 70.775 40.115 ;
        RECT 71.065 40.055 71.680 40.625 ;
        RECT 71.025 39.385 71.195 39.885 ;
        RECT 65.445 38.415 65.785 39.385 ;
        RECT 65.955 38.245 66.125 39.385 ;
        RECT 66.315 39.215 68.750 39.385 ;
        RECT 66.395 38.245 66.645 39.045 ;
        RECT 67.290 38.415 67.620 39.215 ;
        RECT 67.920 38.245 68.250 39.045 ;
        RECT 68.420 38.415 68.750 39.215 ;
        RECT 69.770 39.215 71.195 39.385 ;
        RECT 69.770 39.040 70.160 39.215 ;
        RECT 70.645 38.245 70.975 39.045 ;
        RECT 71.365 39.035 71.680 40.055 ;
        RECT 71.885 40.165 72.225 40.625 ;
        RECT 72.395 40.335 72.565 40.795 ;
        RECT 72.735 40.415 73.905 40.625 ;
        RECT 72.735 40.165 72.985 40.415 ;
        RECT 73.575 40.395 73.905 40.415 ;
        RECT 71.885 39.995 72.985 40.165 ;
        RECT 73.155 39.975 74.015 40.225 ;
        RECT 74.385 40.165 74.715 40.525 ;
        RECT 75.335 40.335 75.585 40.795 ;
        RECT 75.755 40.335 76.315 40.625 ;
        RECT 74.385 39.975 75.775 40.165 ;
        RECT 71.885 39.555 72.645 39.805 ;
        RECT 72.815 39.555 73.565 39.805 ;
        RECT 73.735 39.385 74.015 39.975 ;
        RECT 75.605 39.885 75.775 39.975 ;
        RECT 71.145 38.415 71.680 39.035 ;
        RECT 71.885 38.245 72.145 39.385 ;
        RECT 72.315 39.215 74.015 39.385 ;
        RECT 74.200 39.555 74.875 39.805 ;
        RECT 75.095 39.555 75.435 39.805 ;
        RECT 75.605 39.555 75.895 39.885 ;
        RECT 72.315 38.415 72.645 39.215 ;
        RECT 72.815 38.245 72.985 39.045 ;
        RECT 73.155 38.415 73.485 39.215 ;
        RECT 74.200 39.195 74.465 39.555 ;
        RECT 75.605 39.305 75.775 39.555 ;
        RECT 74.835 39.135 75.775 39.305 ;
        RECT 73.655 38.245 73.910 39.045 ;
        RECT 74.385 38.245 74.665 38.915 ;
        RECT 74.835 38.585 75.135 39.135 ;
        RECT 76.065 38.965 76.315 40.335 ;
        RECT 76.485 40.025 79.995 40.795 ;
        RECT 76.485 39.505 78.135 40.025 ;
        RECT 80.370 40.015 80.870 40.625 ;
        RECT 78.305 39.335 79.995 39.855 ;
        RECT 80.165 39.555 80.515 39.805 ;
        RECT 80.700 39.385 80.870 40.015 ;
        RECT 81.500 40.145 81.830 40.625 ;
        RECT 82.000 40.335 82.225 40.795 ;
        RECT 82.395 40.145 82.725 40.625 ;
        RECT 81.500 39.975 82.725 40.145 ;
        RECT 82.915 39.995 83.165 40.795 ;
        RECT 83.335 39.995 83.675 40.625 ;
        RECT 81.040 39.605 81.370 39.805 ;
        RECT 81.540 39.605 81.870 39.805 ;
        RECT 82.040 39.605 82.460 39.805 ;
        RECT 82.635 39.635 83.330 39.805 ;
        RECT 82.635 39.385 82.805 39.635 ;
        RECT 83.500 39.385 83.675 39.995 ;
        RECT 75.335 38.245 75.665 38.965 ;
        RECT 75.855 38.415 76.315 38.965 ;
        RECT 76.485 38.245 79.995 39.335 ;
        RECT 80.370 39.215 82.805 39.385 ;
        RECT 80.370 38.415 80.700 39.215 ;
        RECT 80.870 38.245 81.200 39.045 ;
        RECT 81.500 38.415 81.830 39.215 ;
        RECT 82.475 38.245 82.725 39.045 ;
        RECT 82.995 38.245 83.165 39.385 ;
        RECT 83.335 38.415 83.675 39.385 ;
        RECT 83.845 40.120 84.105 40.625 ;
        RECT 84.285 40.415 84.615 40.795 ;
        RECT 84.795 40.245 84.965 40.625 ;
        RECT 85.225 40.250 90.570 40.795 ;
        RECT 83.845 39.320 84.025 40.120 ;
        RECT 84.300 40.075 84.965 40.245 ;
        RECT 84.300 39.820 84.470 40.075 ;
        RECT 84.195 39.490 84.470 39.820 ;
        RECT 84.695 39.525 85.035 39.895 ;
        RECT 84.300 39.345 84.470 39.490 ;
        RECT 86.810 39.420 87.150 40.250 ;
        RECT 90.745 40.045 91.955 40.795 ;
        RECT 83.845 38.415 84.115 39.320 ;
        RECT 84.300 39.175 84.975 39.345 ;
        RECT 84.285 38.245 84.615 39.005 ;
        RECT 84.795 38.415 84.975 39.175 ;
        RECT 88.630 38.680 88.980 39.930 ;
        RECT 90.745 39.335 91.265 39.875 ;
        RECT 91.435 39.505 91.955 40.045 ;
        RECT 85.225 38.245 90.570 38.680 ;
        RECT 90.745 38.245 91.955 39.335 ;
        RECT 13.380 38.075 92.040 38.245 ;
        RECT 13.465 36.985 14.675 38.075 ;
        RECT 14.845 36.985 17.435 38.075 ;
        RECT 18.155 37.405 18.325 37.905 ;
        RECT 18.495 37.575 18.825 38.075 ;
        RECT 18.155 37.235 18.820 37.405 ;
        RECT 13.465 36.275 13.985 36.815 ;
        RECT 14.155 36.445 14.675 36.985 ;
        RECT 14.845 36.295 16.055 36.815 ;
        RECT 16.225 36.465 17.435 36.985 ;
        RECT 18.070 36.415 18.420 37.065 ;
        RECT 13.465 35.525 14.675 36.275 ;
        RECT 14.845 35.525 17.435 36.295 ;
        RECT 18.590 36.245 18.820 37.235 ;
        RECT 18.155 36.075 18.820 36.245 ;
        RECT 18.155 35.785 18.325 36.075 ;
        RECT 18.495 35.525 18.825 35.905 ;
        RECT 18.995 35.785 19.180 37.905 ;
        RECT 19.420 37.615 19.685 38.075 ;
        RECT 19.855 37.480 20.105 37.905 ;
        RECT 20.315 37.630 21.420 37.800 ;
        RECT 19.800 37.350 20.105 37.480 ;
        RECT 19.350 36.155 19.630 37.105 ;
        RECT 19.800 36.245 19.970 37.350 ;
        RECT 20.140 36.565 20.380 37.160 ;
        RECT 20.550 37.095 21.080 37.460 ;
        RECT 20.550 36.395 20.720 37.095 ;
        RECT 21.250 37.015 21.420 37.630 ;
        RECT 21.590 37.275 21.760 38.075 ;
        RECT 21.930 37.575 22.180 37.905 ;
        RECT 22.405 37.605 23.290 37.775 ;
        RECT 21.250 36.925 21.760 37.015 ;
        RECT 19.800 36.115 20.025 36.245 ;
        RECT 20.195 36.175 20.720 36.395 ;
        RECT 20.890 36.755 21.760 36.925 ;
        RECT 19.435 35.525 19.685 35.985 ;
        RECT 19.855 35.975 20.025 36.115 ;
        RECT 20.890 35.975 21.060 36.755 ;
        RECT 21.590 36.685 21.760 36.755 ;
        RECT 21.270 36.505 21.470 36.535 ;
        RECT 21.930 36.505 22.100 37.575 ;
        RECT 22.270 36.685 22.460 37.405 ;
        RECT 21.270 36.205 22.100 36.505 ;
        RECT 22.630 36.475 22.950 37.435 ;
        RECT 19.855 35.805 20.190 35.975 ;
        RECT 20.385 35.805 21.060 35.975 ;
        RECT 21.380 35.525 21.750 36.025 ;
        RECT 21.930 35.975 22.100 36.205 ;
        RECT 22.485 36.145 22.950 36.475 ;
        RECT 23.120 36.765 23.290 37.605 ;
        RECT 23.470 37.575 23.785 38.075 ;
        RECT 24.015 37.345 24.355 37.905 ;
        RECT 23.460 36.970 24.355 37.345 ;
        RECT 24.525 37.065 24.695 38.075 ;
        RECT 24.165 36.765 24.355 36.970 ;
        RECT 24.865 37.015 25.195 37.860 ;
        RECT 24.865 36.935 25.255 37.015 ;
        RECT 25.040 36.885 25.255 36.935 ;
        RECT 26.345 36.910 26.635 38.075 ;
        RECT 26.840 37.285 27.375 37.905 ;
        RECT 23.120 36.435 23.995 36.765 ;
        RECT 24.165 36.435 24.915 36.765 ;
        RECT 23.120 35.975 23.290 36.435 ;
        RECT 24.165 36.265 24.365 36.435 ;
        RECT 25.085 36.305 25.255 36.885 ;
        RECT 25.030 36.265 25.255 36.305 ;
        RECT 21.930 35.805 22.335 35.975 ;
        RECT 22.505 35.805 23.290 35.975 ;
        RECT 23.565 35.525 23.775 36.055 ;
        RECT 24.035 35.740 24.365 36.265 ;
        RECT 24.875 36.180 25.255 36.265 ;
        RECT 26.840 36.265 27.155 37.285 ;
        RECT 27.545 37.275 27.875 38.075 ;
        RECT 28.360 37.105 28.750 37.280 ;
        RECT 27.325 36.935 28.750 37.105 ;
        RECT 30.230 37.105 30.560 37.905 ;
        RECT 30.730 37.275 31.060 38.075 ;
        RECT 31.360 37.105 31.690 37.905 ;
        RECT 32.335 37.275 32.585 38.075 ;
        RECT 30.230 36.935 32.665 37.105 ;
        RECT 32.855 36.935 33.025 38.075 ;
        RECT 33.195 36.935 33.535 37.905 ;
        RECT 33.810 37.275 34.065 38.075 ;
        RECT 34.235 37.105 34.565 37.905 ;
        RECT 34.735 37.275 34.905 38.075 ;
        RECT 35.075 37.105 35.405 37.905 ;
        RECT 27.325 36.435 27.495 36.935 ;
        RECT 24.535 35.525 24.705 36.135 ;
        RECT 24.875 35.745 25.205 36.180 ;
        RECT 26.345 35.525 26.635 36.250 ;
        RECT 26.840 35.695 27.455 36.265 ;
        RECT 27.745 36.205 28.010 36.765 ;
        RECT 28.180 36.035 28.350 36.935 ;
        RECT 28.520 36.205 28.875 36.765 ;
        RECT 30.025 36.515 30.375 36.765 ;
        RECT 30.560 36.305 30.730 36.935 ;
        RECT 30.900 36.515 31.230 36.715 ;
        RECT 31.400 36.515 31.730 36.715 ;
        RECT 31.900 36.515 32.320 36.715 ;
        RECT 32.495 36.685 32.665 36.935 ;
        RECT 32.495 36.515 33.190 36.685 ;
        RECT 27.625 35.525 27.840 36.035 ;
        RECT 28.070 35.705 28.350 36.035 ;
        RECT 28.530 35.525 28.770 36.035 ;
        RECT 30.230 35.695 30.730 36.305 ;
        RECT 31.360 36.175 32.585 36.345 ;
        RECT 33.360 36.325 33.535 36.935 ;
        RECT 31.360 35.695 31.690 36.175 ;
        RECT 31.860 35.525 32.085 35.985 ;
        RECT 32.255 35.695 32.585 36.175 ;
        RECT 32.775 35.525 33.025 36.325 ;
        RECT 33.195 35.695 33.535 36.325 ;
        RECT 33.705 36.935 35.405 37.105 ;
        RECT 35.575 36.935 35.835 38.075 ;
        RECT 36.005 36.985 37.675 38.075 ;
        RECT 37.905 37.015 38.235 37.860 ;
        RECT 38.405 37.065 38.575 38.075 ;
        RECT 38.745 37.345 39.085 37.905 ;
        RECT 39.315 37.575 39.630 38.075 ;
        RECT 39.810 37.605 40.695 37.775 ;
        RECT 33.705 36.345 33.985 36.935 ;
        RECT 34.155 36.515 34.905 36.765 ;
        RECT 35.075 36.515 35.835 36.765 ;
        RECT 33.705 36.095 34.565 36.345 ;
        RECT 34.735 36.155 35.835 36.325 ;
        RECT 33.815 35.905 34.145 35.925 ;
        RECT 34.735 35.905 34.985 36.155 ;
        RECT 33.815 35.695 34.985 35.905 ;
        RECT 35.155 35.525 35.325 35.985 ;
        RECT 35.495 35.695 35.835 36.155 ;
        RECT 36.005 36.295 36.755 36.815 ;
        RECT 36.925 36.465 37.675 36.985 ;
        RECT 37.845 36.935 38.235 37.015 ;
        RECT 38.745 36.970 39.640 37.345 ;
        RECT 37.845 36.885 38.060 36.935 ;
        RECT 37.845 36.305 38.015 36.885 ;
        RECT 38.745 36.765 38.935 36.970 ;
        RECT 39.810 36.765 39.980 37.605 ;
        RECT 40.920 37.575 41.170 37.905 ;
        RECT 38.185 36.435 38.935 36.765 ;
        RECT 39.105 36.435 39.980 36.765 ;
        RECT 36.005 35.525 37.675 36.295 ;
        RECT 37.845 36.265 38.070 36.305 ;
        RECT 38.735 36.265 38.935 36.435 ;
        RECT 37.845 36.180 38.225 36.265 ;
        RECT 37.895 35.745 38.225 36.180 ;
        RECT 38.395 35.525 38.565 36.135 ;
        RECT 38.735 35.740 39.065 36.265 ;
        RECT 39.325 35.525 39.535 36.055 ;
        RECT 39.810 35.975 39.980 36.435 ;
        RECT 40.150 36.475 40.470 37.435 ;
        RECT 40.640 36.685 40.830 37.405 ;
        RECT 41.000 36.505 41.170 37.575 ;
        RECT 41.340 37.275 41.510 38.075 ;
        RECT 41.680 37.630 42.785 37.800 ;
        RECT 41.680 37.015 41.850 37.630 ;
        RECT 42.995 37.480 43.245 37.905 ;
        RECT 43.415 37.615 43.680 38.075 ;
        RECT 42.020 37.095 42.550 37.460 ;
        RECT 42.995 37.350 43.300 37.480 ;
        RECT 41.340 36.925 41.850 37.015 ;
        RECT 41.340 36.755 42.210 36.925 ;
        RECT 41.340 36.685 41.510 36.755 ;
        RECT 41.630 36.505 41.830 36.535 ;
        RECT 40.150 36.145 40.615 36.475 ;
        RECT 41.000 36.205 41.830 36.505 ;
        RECT 41.000 35.975 41.170 36.205 ;
        RECT 39.810 35.805 40.595 35.975 ;
        RECT 40.765 35.805 41.170 35.975 ;
        RECT 41.350 35.525 41.720 36.025 ;
        RECT 42.040 35.975 42.210 36.755 ;
        RECT 42.380 36.395 42.550 37.095 ;
        RECT 42.720 36.565 42.960 37.160 ;
        RECT 42.380 36.175 42.905 36.395 ;
        RECT 43.130 36.245 43.300 37.350 ;
        RECT 43.075 36.115 43.300 36.245 ;
        RECT 43.470 36.155 43.750 37.105 ;
        RECT 43.075 35.975 43.245 36.115 ;
        RECT 42.040 35.805 42.715 35.975 ;
        RECT 42.910 35.805 43.245 35.975 ;
        RECT 43.415 35.525 43.665 35.985 ;
        RECT 43.920 35.785 44.105 37.905 ;
        RECT 44.275 37.575 44.605 38.075 ;
        RECT 44.775 37.405 44.945 37.905 ;
        RECT 44.280 37.235 44.945 37.405 ;
        RECT 44.280 36.245 44.510 37.235 ;
        RECT 44.680 36.415 45.030 37.065 ;
        RECT 45.205 36.935 45.545 37.905 ;
        RECT 45.715 36.935 45.885 38.075 ;
        RECT 46.155 37.275 46.405 38.075 ;
        RECT 47.050 37.105 47.380 37.905 ;
        RECT 47.680 37.275 48.010 38.075 ;
        RECT 48.180 37.105 48.510 37.905 ;
        RECT 46.075 36.935 48.510 37.105 ;
        RECT 48.885 36.985 51.475 38.075 ;
        RECT 45.205 36.375 45.380 36.935 ;
        RECT 46.075 36.685 46.245 36.935 ;
        RECT 45.550 36.515 46.245 36.685 ;
        RECT 46.420 36.515 46.840 36.715 ;
        RECT 47.010 36.515 47.340 36.715 ;
        RECT 47.510 36.515 47.840 36.715 ;
        RECT 45.205 36.325 45.435 36.375 ;
        RECT 44.280 36.075 44.945 36.245 ;
        RECT 44.275 35.525 44.605 35.905 ;
        RECT 44.775 35.785 44.945 36.075 ;
        RECT 45.205 35.695 45.545 36.325 ;
        RECT 45.715 35.525 45.965 36.325 ;
        RECT 46.155 36.175 47.380 36.345 ;
        RECT 46.155 35.695 46.485 36.175 ;
        RECT 46.655 35.525 46.880 35.985 ;
        RECT 47.050 35.695 47.380 36.175 ;
        RECT 48.010 36.305 48.180 36.935 ;
        RECT 48.365 36.515 48.715 36.765 ;
        RECT 48.010 35.695 48.510 36.305 ;
        RECT 48.885 36.295 50.095 36.815 ;
        RECT 50.265 36.465 51.475 36.985 ;
        RECT 52.105 36.910 52.395 38.075 ;
        RECT 52.565 36.985 55.155 38.075 ;
        RECT 52.565 36.295 53.775 36.815 ;
        RECT 53.945 36.465 55.155 36.985 ;
        RECT 55.330 36.935 55.665 37.905 ;
        RECT 55.835 36.935 56.005 38.075 ;
        RECT 56.175 37.735 58.205 37.905 ;
        RECT 48.885 35.525 51.475 36.295 ;
        RECT 52.105 35.525 52.395 36.250 ;
        RECT 52.565 35.525 55.155 36.295 ;
        RECT 55.330 36.265 55.500 36.935 ;
        RECT 56.175 36.765 56.345 37.735 ;
        RECT 55.670 36.435 55.925 36.765 ;
        RECT 56.150 36.435 56.345 36.765 ;
        RECT 56.515 37.395 57.640 37.565 ;
        RECT 55.755 36.265 55.925 36.435 ;
        RECT 56.515 36.265 56.685 37.395 ;
        RECT 55.330 35.695 55.585 36.265 ;
        RECT 55.755 36.095 56.685 36.265 ;
        RECT 56.855 37.055 57.865 37.225 ;
        RECT 56.855 36.255 57.025 37.055 ;
        RECT 57.230 36.375 57.505 36.855 ;
        RECT 57.225 36.205 57.505 36.375 ;
        RECT 56.510 36.060 56.685 36.095 ;
        RECT 55.755 35.525 56.085 35.925 ;
        RECT 56.510 35.695 57.040 36.060 ;
        RECT 57.230 35.695 57.505 36.205 ;
        RECT 57.675 35.695 57.865 37.055 ;
        RECT 58.035 37.070 58.205 37.735 ;
        RECT 58.375 37.315 58.545 38.075 ;
        RECT 58.780 37.315 59.295 37.725 ;
        RECT 58.035 36.880 58.785 37.070 ;
        RECT 58.955 36.505 59.295 37.315 ;
        RECT 58.065 36.335 59.295 36.505 ;
        RECT 59.465 36.935 59.850 37.905 ;
        RECT 60.020 37.615 60.345 38.075 ;
        RECT 60.865 37.445 61.145 37.905 ;
        RECT 60.020 37.225 61.145 37.445 ;
        RECT 58.045 35.525 58.555 36.060 ;
        RECT 58.775 35.730 59.020 36.335 ;
        RECT 59.465 36.265 59.745 36.935 ;
        RECT 60.020 36.765 60.470 37.225 ;
        RECT 61.335 37.055 61.735 37.905 ;
        RECT 62.135 37.615 62.405 38.075 ;
        RECT 62.575 37.445 62.860 37.905 ;
        RECT 59.915 36.435 60.470 36.765 ;
        RECT 60.640 36.495 61.735 37.055 ;
        RECT 60.020 36.325 60.470 36.435 ;
        RECT 59.465 35.695 59.850 36.265 ;
        RECT 60.020 36.155 61.145 36.325 ;
        RECT 60.020 35.525 60.345 35.985 ;
        RECT 60.865 35.695 61.145 36.155 ;
        RECT 61.335 35.695 61.735 36.495 ;
        RECT 61.905 37.225 62.860 37.445 ;
        RECT 61.905 36.325 62.115 37.225 ;
        RECT 63.145 37.105 63.415 37.875 ;
        RECT 63.585 37.295 63.915 38.075 ;
        RECT 64.120 37.470 64.305 37.875 ;
        RECT 64.475 37.650 64.810 38.075 ;
        RECT 64.985 37.640 70.330 38.075 ;
        RECT 64.120 37.295 64.785 37.470 ;
        RECT 62.285 36.495 62.975 37.055 ;
        RECT 63.145 36.935 64.275 37.105 ;
        RECT 61.905 36.155 62.860 36.325 ;
        RECT 62.135 35.525 62.405 35.985 ;
        RECT 62.575 35.695 62.860 36.155 ;
        RECT 63.145 36.025 63.315 36.935 ;
        RECT 63.485 36.185 63.845 36.765 ;
        RECT 64.025 36.435 64.275 36.935 ;
        RECT 64.445 36.265 64.785 37.295 ;
        RECT 64.100 36.095 64.785 36.265 ;
        RECT 63.145 35.695 63.405 36.025 ;
        RECT 63.615 35.525 63.890 36.005 ;
        RECT 64.100 35.695 64.305 36.095 ;
        RECT 66.570 36.070 66.910 36.900 ;
        RECT 68.390 36.390 68.740 37.640 ;
        RECT 70.505 36.985 74.015 38.075 ;
        RECT 74.185 36.985 75.395 38.075 ;
        RECT 70.505 36.295 72.155 36.815 ;
        RECT 72.325 36.465 74.015 36.985 ;
        RECT 64.475 35.525 64.810 35.925 ;
        RECT 64.985 35.525 70.330 36.070 ;
        RECT 70.505 35.525 74.015 36.295 ;
        RECT 74.185 36.275 74.705 36.815 ;
        RECT 74.875 36.445 75.395 36.985 ;
        RECT 75.750 37.105 76.140 37.280 ;
        RECT 76.625 37.275 76.955 38.075 ;
        RECT 77.125 37.285 77.660 37.905 ;
        RECT 75.750 36.935 77.175 37.105 ;
        RECT 74.185 35.525 75.395 36.275 ;
        RECT 75.625 36.205 75.980 36.765 ;
        RECT 76.150 36.035 76.320 36.935 ;
        RECT 76.490 36.205 76.755 36.765 ;
        RECT 77.005 36.435 77.175 36.935 ;
        RECT 77.345 36.265 77.660 37.285 ;
        RECT 77.865 36.910 78.155 38.075 ;
        RECT 79.450 37.105 79.780 37.905 ;
        RECT 79.950 37.275 80.280 38.075 ;
        RECT 80.580 37.105 80.910 37.905 ;
        RECT 81.555 37.275 81.805 38.075 ;
        RECT 79.450 36.935 81.885 37.105 ;
        RECT 82.075 36.935 82.245 38.075 ;
        RECT 82.415 36.935 82.755 37.905 ;
        RECT 83.015 37.405 83.185 37.905 ;
        RECT 83.355 37.575 83.685 38.075 ;
        RECT 83.015 37.235 83.680 37.405 ;
        RECT 79.245 36.515 79.595 36.765 ;
        RECT 79.780 36.305 79.950 36.935 ;
        RECT 80.120 36.515 80.450 36.715 ;
        RECT 80.620 36.515 80.950 36.715 ;
        RECT 81.120 36.515 81.540 36.715 ;
        RECT 81.715 36.685 81.885 36.935 ;
        RECT 81.715 36.515 82.410 36.685 ;
        RECT 82.580 36.375 82.755 36.935 ;
        RECT 82.930 36.415 83.280 37.065 ;
        RECT 75.730 35.525 75.970 36.035 ;
        RECT 76.150 35.705 76.430 36.035 ;
        RECT 76.660 35.525 76.875 36.035 ;
        RECT 77.045 35.695 77.660 36.265 ;
        RECT 77.865 35.525 78.155 36.250 ;
        RECT 79.450 35.695 79.950 36.305 ;
        RECT 80.580 36.175 81.805 36.345 ;
        RECT 82.525 36.325 82.755 36.375 ;
        RECT 80.580 35.695 80.910 36.175 ;
        RECT 81.080 35.525 81.305 35.985 ;
        RECT 81.475 35.695 81.805 36.175 ;
        RECT 81.995 35.525 82.245 36.325 ;
        RECT 82.415 35.695 82.755 36.325 ;
        RECT 83.450 36.245 83.680 37.235 ;
        RECT 83.015 36.075 83.680 36.245 ;
        RECT 83.015 35.785 83.185 36.075 ;
        RECT 83.355 35.525 83.685 35.905 ;
        RECT 83.855 35.785 84.040 37.905 ;
        RECT 84.280 37.615 84.545 38.075 ;
        RECT 84.715 37.480 84.965 37.905 ;
        RECT 85.175 37.630 86.280 37.800 ;
        RECT 84.660 37.350 84.965 37.480 ;
        RECT 84.210 36.155 84.490 37.105 ;
        RECT 84.660 36.245 84.830 37.350 ;
        RECT 85.000 36.565 85.240 37.160 ;
        RECT 85.410 37.095 85.940 37.460 ;
        RECT 85.410 36.395 85.580 37.095 ;
        RECT 86.110 37.015 86.280 37.630 ;
        RECT 86.450 37.275 86.620 38.075 ;
        RECT 86.790 37.575 87.040 37.905 ;
        RECT 87.265 37.605 88.150 37.775 ;
        RECT 86.110 36.925 86.620 37.015 ;
        RECT 84.660 36.115 84.885 36.245 ;
        RECT 85.055 36.175 85.580 36.395 ;
        RECT 85.750 36.755 86.620 36.925 ;
        RECT 84.295 35.525 84.545 35.985 ;
        RECT 84.715 35.975 84.885 36.115 ;
        RECT 85.750 35.975 85.920 36.755 ;
        RECT 86.450 36.685 86.620 36.755 ;
        RECT 86.130 36.505 86.330 36.535 ;
        RECT 86.790 36.505 86.960 37.575 ;
        RECT 87.130 36.685 87.320 37.405 ;
        RECT 86.130 36.205 86.960 36.505 ;
        RECT 87.490 36.475 87.810 37.435 ;
        RECT 84.715 35.805 85.050 35.975 ;
        RECT 85.245 35.805 85.920 35.975 ;
        RECT 86.240 35.525 86.610 36.025 ;
        RECT 86.790 35.975 86.960 36.205 ;
        RECT 87.345 36.145 87.810 36.475 ;
        RECT 87.980 36.765 88.150 37.605 ;
        RECT 88.330 37.575 88.645 38.075 ;
        RECT 88.875 37.345 89.215 37.905 ;
        RECT 88.320 36.970 89.215 37.345 ;
        RECT 89.385 37.065 89.555 38.075 ;
        RECT 89.025 36.765 89.215 36.970 ;
        RECT 89.725 37.015 90.055 37.860 ;
        RECT 89.725 36.935 90.115 37.015 ;
        RECT 89.900 36.885 90.115 36.935 ;
        RECT 87.980 36.435 88.855 36.765 ;
        RECT 89.025 36.435 89.775 36.765 ;
        RECT 87.980 35.975 88.150 36.435 ;
        RECT 89.025 36.265 89.225 36.435 ;
        RECT 89.945 36.305 90.115 36.885 ;
        RECT 90.745 36.985 91.955 38.075 ;
        RECT 90.745 36.445 91.265 36.985 ;
        RECT 89.890 36.265 90.115 36.305 ;
        RECT 91.435 36.275 91.955 36.815 ;
        RECT 86.790 35.805 87.195 35.975 ;
        RECT 87.365 35.805 88.150 35.975 ;
        RECT 88.425 35.525 88.635 36.055 ;
        RECT 88.895 35.740 89.225 36.265 ;
        RECT 89.735 36.180 90.115 36.265 ;
        RECT 89.395 35.525 89.565 36.135 ;
        RECT 89.735 35.745 90.065 36.180 ;
        RECT 90.745 35.525 91.955 36.275 ;
        RECT 13.380 35.355 92.040 35.525 ;
        RECT 13.465 34.605 14.675 35.355 ;
        RECT 14.845 34.810 20.190 35.355 ;
        RECT 13.465 34.065 13.985 34.605 ;
        RECT 14.155 33.895 14.675 34.435 ;
        RECT 16.430 33.980 16.770 34.810 ;
        RECT 21.285 34.555 21.625 35.185 ;
        RECT 21.795 34.555 22.045 35.355 ;
        RECT 22.235 34.705 22.565 35.185 ;
        RECT 22.735 34.895 22.960 35.355 ;
        RECT 23.130 34.705 23.460 35.185 ;
        RECT 13.465 32.805 14.675 33.895 ;
        RECT 18.250 33.240 18.600 34.490 ;
        RECT 21.285 33.945 21.460 34.555 ;
        RECT 22.235 34.535 23.460 34.705 ;
        RECT 24.090 34.575 24.590 35.185 ;
        RECT 25.055 34.805 25.225 35.185 ;
        RECT 25.440 34.975 25.770 35.355 ;
        RECT 25.055 34.635 25.770 34.805 ;
        RECT 21.630 34.195 22.325 34.365 ;
        RECT 22.155 33.945 22.325 34.195 ;
        RECT 22.500 34.165 22.920 34.365 ;
        RECT 23.090 34.165 23.420 34.365 ;
        RECT 23.590 34.165 23.920 34.365 ;
        RECT 24.090 33.945 24.260 34.575 ;
        RECT 24.445 34.115 24.795 34.365 ;
        RECT 24.965 34.085 25.320 34.455 ;
        RECT 25.600 34.445 25.770 34.635 ;
        RECT 25.940 34.610 26.195 35.185 ;
        RECT 25.600 34.115 25.855 34.445 ;
        RECT 14.845 32.805 20.190 33.240 ;
        RECT 21.285 32.975 21.625 33.945 ;
        RECT 21.795 32.805 21.965 33.945 ;
        RECT 22.155 33.775 24.590 33.945 ;
        RECT 25.600 33.905 25.770 34.115 ;
        RECT 22.235 32.805 22.485 33.605 ;
        RECT 23.130 32.975 23.460 33.775 ;
        RECT 23.760 32.805 24.090 33.605 ;
        RECT 24.260 32.975 24.590 33.775 ;
        RECT 25.055 33.735 25.770 33.905 ;
        RECT 26.025 33.880 26.195 34.610 ;
        RECT 26.370 34.515 26.630 35.355 ;
        RECT 26.805 34.585 28.475 35.355 ;
        RECT 28.810 34.845 29.050 35.355 ;
        RECT 29.230 34.845 29.510 35.175 ;
        RECT 29.740 34.845 29.955 35.355 ;
        RECT 26.805 34.065 27.555 34.585 ;
        RECT 25.055 32.975 25.225 33.735 ;
        RECT 25.440 32.805 25.770 33.565 ;
        RECT 25.940 32.975 26.195 33.880 ;
        RECT 26.370 32.805 26.630 33.955 ;
        RECT 27.725 33.895 28.475 34.415 ;
        RECT 28.705 34.115 29.060 34.675 ;
        RECT 29.230 33.945 29.400 34.845 ;
        RECT 29.570 34.115 29.835 34.675 ;
        RECT 30.125 34.615 30.740 35.185 ;
        RECT 31.035 34.805 31.205 35.095 ;
        RECT 31.375 34.975 31.705 35.355 ;
        RECT 31.035 34.635 31.700 34.805 ;
        RECT 30.085 33.945 30.255 34.445 ;
        RECT 26.805 32.805 28.475 33.895 ;
        RECT 28.830 33.775 30.255 33.945 ;
        RECT 28.830 33.600 29.220 33.775 ;
        RECT 29.705 32.805 30.035 33.605 ;
        RECT 30.425 33.595 30.740 34.615 ;
        RECT 30.950 33.815 31.300 34.465 ;
        RECT 31.470 33.645 31.700 34.635 ;
        RECT 30.205 32.975 30.740 33.595 ;
        RECT 31.035 33.475 31.700 33.645 ;
        RECT 31.035 32.975 31.205 33.475 ;
        RECT 31.375 32.805 31.705 33.305 ;
        RECT 31.875 32.975 32.060 35.095 ;
        RECT 32.315 34.895 32.565 35.355 ;
        RECT 32.735 34.905 33.070 35.075 ;
        RECT 33.265 34.905 33.940 35.075 ;
        RECT 32.735 34.765 32.905 34.905 ;
        RECT 32.230 33.775 32.510 34.725 ;
        RECT 32.680 34.635 32.905 34.765 ;
        RECT 32.680 33.530 32.850 34.635 ;
        RECT 33.075 34.485 33.600 34.705 ;
        RECT 33.020 33.720 33.260 34.315 ;
        RECT 33.430 33.785 33.600 34.485 ;
        RECT 33.770 34.125 33.940 34.905 ;
        RECT 34.260 34.855 34.630 35.355 ;
        RECT 34.810 34.905 35.215 35.075 ;
        RECT 35.385 34.905 36.170 35.075 ;
        RECT 34.810 34.675 34.980 34.905 ;
        RECT 34.150 34.375 34.980 34.675 ;
        RECT 35.365 34.405 35.830 34.735 ;
        RECT 34.150 34.345 34.350 34.375 ;
        RECT 34.470 34.125 34.640 34.195 ;
        RECT 33.770 33.955 34.640 34.125 ;
        RECT 34.130 33.865 34.640 33.955 ;
        RECT 32.680 33.400 32.985 33.530 ;
        RECT 33.430 33.420 33.960 33.785 ;
        RECT 32.300 32.805 32.565 33.265 ;
        RECT 32.735 32.975 32.985 33.400 ;
        RECT 34.130 33.250 34.300 33.865 ;
        RECT 33.195 33.080 34.300 33.250 ;
        RECT 34.470 32.805 34.640 33.605 ;
        RECT 34.810 33.305 34.980 34.375 ;
        RECT 35.150 33.475 35.340 34.195 ;
        RECT 35.510 33.445 35.830 34.405 ;
        RECT 36.000 34.445 36.170 34.905 ;
        RECT 36.445 34.825 36.655 35.355 ;
        RECT 36.915 34.615 37.245 35.140 ;
        RECT 37.415 34.745 37.585 35.355 ;
        RECT 37.755 34.700 38.085 35.135 ;
        RECT 37.755 34.615 38.135 34.700 ;
        RECT 39.225 34.630 39.515 35.355 ;
        RECT 37.045 34.445 37.245 34.615 ;
        RECT 37.910 34.575 38.135 34.615 ;
        RECT 39.690 34.590 40.145 35.355 ;
        RECT 40.420 34.975 41.720 35.185 ;
        RECT 41.975 34.995 42.305 35.355 ;
        RECT 41.550 34.825 41.720 34.975 ;
        RECT 42.475 34.855 42.735 35.185 ;
        RECT 42.505 34.845 42.735 34.855 ;
        RECT 43.070 34.845 43.310 35.355 ;
        RECT 43.490 34.845 43.770 35.175 ;
        RECT 44.000 34.845 44.215 35.355 ;
        RECT 36.000 34.115 36.875 34.445 ;
        RECT 37.045 34.115 37.795 34.445 ;
        RECT 34.810 32.975 35.060 33.305 ;
        RECT 36.000 33.275 36.170 34.115 ;
        RECT 37.045 33.910 37.235 34.115 ;
        RECT 37.965 33.995 38.135 34.575 ;
        RECT 40.620 34.365 40.840 34.765 ;
        RECT 39.685 34.165 40.175 34.365 ;
        RECT 40.365 34.155 40.840 34.365 ;
        RECT 41.085 34.365 41.295 34.765 ;
        RECT 41.550 34.700 42.305 34.825 ;
        RECT 41.550 34.655 42.395 34.700 ;
        RECT 42.125 34.535 42.395 34.655 ;
        RECT 41.085 34.155 41.415 34.365 ;
        RECT 41.585 34.095 41.995 34.400 ;
        RECT 37.920 33.945 38.135 33.995 ;
        RECT 36.340 33.535 37.235 33.910 ;
        RECT 37.745 33.865 38.135 33.945 ;
        RECT 35.285 33.105 36.170 33.275 ;
        RECT 36.350 32.805 36.665 33.305 ;
        RECT 36.895 32.975 37.235 33.535 ;
        RECT 37.405 32.805 37.575 33.815 ;
        RECT 37.745 33.020 38.075 33.865 ;
        RECT 39.225 32.805 39.515 33.970 ;
        RECT 39.690 33.925 40.865 33.985 ;
        RECT 42.225 33.960 42.395 34.535 ;
        RECT 42.195 33.925 42.395 33.960 ;
        RECT 39.690 33.815 42.395 33.925 ;
        RECT 39.690 33.195 39.945 33.815 ;
        RECT 40.535 33.755 42.335 33.815 ;
        RECT 40.535 33.725 40.865 33.755 ;
        RECT 42.565 33.655 42.735 34.845 ;
        RECT 42.965 34.115 43.320 34.675 ;
        RECT 43.490 33.945 43.660 34.845 ;
        RECT 43.830 34.115 44.095 34.675 ;
        RECT 44.385 34.615 45.000 35.185 ;
        RECT 45.205 34.810 50.550 35.355 ;
        RECT 44.345 33.945 44.515 34.445 ;
        RECT 40.195 33.555 40.380 33.645 ;
        RECT 40.970 33.555 41.805 33.565 ;
        RECT 40.195 33.355 41.805 33.555 ;
        RECT 40.195 33.315 40.425 33.355 ;
        RECT 39.690 32.975 40.025 33.195 ;
        RECT 41.030 32.805 41.385 33.185 ;
        RECT 41.555 32.975 41.805 33.355 ;
        RECT 42.055 32.805 42.305 33.585 ;
        RECT 42.475 32.975 42.735 33.655 ;
        RECT 43.090 33.775 44.515 33.945 ;
        RECT 43.090 33.600 43.480 33.775 ;
        RECT 43.965 32.805 44.295 33.605 ;
        RECT 44.685 33.595 45.000 34.615 ;
        RECT 46.790 33.980 47.130 34.810 ;
        RECT 50.725 34.585 52.395 35.355 ;
        RECT 44.465 32.975 45.000 33.595 ;
        RECT 48.610 33.240 48.960 34.490 ;
        RECT 50.725 34.065 51.475 34.585 ;
        RECT 52.570 34.535 52.845 35.355 ;
        RECT 53.015 34.715 53.345 35.185 ;
        RECT 53.515 34.885 53.685 35.355 ;
        RECT 53.855 34.715 54.185 35.185 ;
        RECT 54.355 34.885 55.065 35.355 ;
        RECT 55.235 34.715 55.565 35.185 ;
        RECT 55.735 34.885 56.025 35.355 ;
        RECT 53.015 34.535 56.075 34.715 ;
        RECT 51.645 33.895 52.395 34.415 ;
        RECT 52.615 34.155 53.445 34.365 ;
        RECT 53.615 34.155 54.665 34.365 ;
        RECT 54.855 34.155 55.445 34.365 ;
        RECT 45.205 32.805 50.550 33.240 ;
        RECT 50.725 32.805 52.395 33.895 ;
        RECT 52.630 33.815 54.565 33.985 ;
        RECT 54.855 33.815 55.120 34.155 ;
        RECT 55.615 33.985 56.075 34.535 ;
        RECT 56.245 34.605 57.455 35.355 ;
        RECT 57.715 34.805 57.885 35.095 ;
        RECT 58.055 34.975 58.385 35.355 ;
        RECT 57.715 34.635 58.380 34.805 ;
        RECT 56.245 34.065 56.765 34.605 ;
        RECT 55.315 33.815 56.075 33.985 ;
        RECT 56.935 33.895 57.455 34.435 ;
        RECT 52.630 32.975 52.885 33.815 ;
        RECT 53.055 32.805 53.305 33.645 ;
        RECT 53.475 32.975 53.725 33.815 ;
        RECT 53.895 33.145 54.145 33.645 ;
        RECT 54.315 33.315 54.565 33.815 ;
        RECT 54.895 33.145 55.105 33.645 ;
        RECT 55.315 33.315 55.525 33.815 ;
        RECT 55.695 33.145 55.945 33.645 ;
        RECT 53.895 32.975 55.945 33.145 ;
        RECT 56.245 32.805 57.455 33.895 ;
        RECT 57.630 33.815 57.980 34.465 ;
        RECT 58.150 33.645 58.380 34.635 ;
        RECT 57.715 33.475 58.380 33.645 ;
        RECT 57.715 32.975 57.885 33.475 ;
        RECT 58.055 32.805 58.385 33.305 ;
        RECT 58.555 32.975 58.740 35.095 ;
        RECT 58.995 34.895 59.245 35.355 ;
        RECT 59.415 34.905 59.750 35.075 ;
        RECT 59.945 34.905 60.620 35.075 ;
        RECT 59.415 34.765 59.585 34.905 ;
        RECT 58.910 33.775 59.190 34.725 ;
        RECT 59.360 34.635 59.585 34.765 ;
        RECT 59.360 33.530 59.530 34.635 ;
        RECT 59.755 34.485 60.280 34.705 ;
        RECT 59.700 33.720 59.940 34.315 ;
        RECT 60.110 33.785 60.280 34.485 ;
        RECT 60.450 34.125 60.620 34.905 ;
        RECT 60.940 34.855 61.310 35.355 ;
        RECT 61.490 34.905 61.895 35.075 ;
        RECT 62.065 34.905 62.850 35.075 ;
        RECT 61.490 34.675 61.660 34.905 ;
        RECT 60.830 34.375 61.660 34.675 ;
        RECT 62.045 34.405 62.510 34.735 ;
        RECT 60.830 34.345 61.030 34.375 ;
        RECT 61.150 34.125 61.320 34.195 ;
        RECT 60.450 33.955 61.320 34.125 ;
        RECT 60.810 33.865 61.320 33.955 ;
        RECT 59.360 33.400 59.665 33.530 ;
        RECT 60.110 33.420 60.640 33.785 ;
        RECT 58.980 32.805 59.245 33.265 ;
        RECT 59.415 32.975 59.665 33.400 ;
        RECT 60.810 33.250 60.980 33.865 ;
        RECT 59.875 33.080 60.980 33.250 ;
        RECT 61.150 32.805 61.320 33.605 ;
        RECT 61.490 33.305 61.660 34.375 ;
        RECT 61.830 33.475 62.020 34.195 ;
        RECT 62.190 33.445 62.510 34.405 ;
        RECT 62.680 34.445 62.850 34.905 ;
        RECT 63.125 34.825 63.335 35.355 ;
        RECT 63.595 34.615 63.925 35.140 ;
        RECT 64.095 34.745 64.265 35.355 ;
        RECT 64.435 34.700 64.765 35.135 ;
        RECT 64.435 34.615 64.815 34.700 ;
        RECT 64.985 34.630 65.275 35.355 ;
        RECT 63.725 34.445 63.925 34.615 ;
        RECT 64.590 34.575 64.815 34.615 ;
        RECT 62.680 34.115 63.555 34.445 ;
        RECT 63.725 34.115 64.475 34.445 ;
        RECT 61.490 32.975 61.740 33.305 ;
        RECT 62.680 33.275 62.850 34.115 ;
        RECT 63.725 33.910 63.915 34.115 ;
        RECT 64.645 33.995 64.815 34.575 ;
        RECT 65.445 34.585 68.955 35.355 ;
        RECT 65.445 34.065 67.095 34.585 ;
        RECT 69.585 34.555 69.875 35.355 ;
        RECT 70.045 34.895 70.595 35.185 ;
        RECT 70.765 34.895 71.015 35.355 ;
        RECT 64.600 33.945 64.815 33.995 ;
        RECT 63.020 33.535 63.915 33.910 ;
        RECT 64.425 33.865 64.815 33.945 ;
        RECT 61.965 33.105 62.850 33.275 ;
        RECT 63.030 32.805 63.345 33.305 ;
        RECT 63.575 32.975 63.915 33.535 ;
        RECT 64.085 32.805 64.255 33.815 ;
        RECT 64.425 33.020 64.755 33.865 ;
        RECT 64.985 32.805 65.275 33.970 ;
        RECT 67.265 33.895 68.955 34.415 ;
        RECT 65.445 32.805 68.955 33.895 ;
        RECT 69.585 32.805 69.875 33.945 ;
        RECT 70.045 33.525 70.295 34.895 ;
        RECT 71.645 34.725 71.975 35.085 ;
        RECT 70.585 34.535 71.975 34.725 ;
        RECT 72.345 34.725 72.685 35.185 ;
        RECT 72.855 34.895 73.025 35.355 ;
        RECT 73.195 34.975 74.365 35.185 ;
        RECT 73.195 34.725 73.445 34.975 ;
        RECT 74.035 34.955 74.365 34.975 ;
        RECT 72.345 34.555 73.445 34.725 ;
        RECT 73.615 34.535 74.475 34.785 ;
        RECT 70.585 34.445 70.755 34.535 ;
        RECT 70.465 34.115 70.755 34.445 ;
        RECT 70.925 34.115 71.255 34.365 ;
        RECT 71.485 34.115 72.175 34.365 ;
        RECT 72.345 34.115 73.105 34.365 ;
        RECT 73.275 34.115 74.025 34.365 ;
        RECT 70.585 33.865 70.755 34.115 ;
        RECT 70.585 33.695 71.525 33.865 ;
        RECT 70.045 32.975 70.495 33.525 ;
        RECT 70.685 32.805 71.015 33.525 ;
        RECT 71.225 33.145 71.525 33.695 ;
        RECT 71.860 33.675 72.175 34.115 ;
        RECT 74.195 33.945 74.475 34.535 ;
        RECT 74.645 34.585 76.315 35.355 ;
        RECT 77.110 34.845 77.350 35.355 ;
        RECT 77.530 34.845 77.810 35.175 ;
        RECT 78.040 34.845 78.255 35.355 ;
        RECT 74.645 34.065 75.395 34.585 ;
        RECT 71.695 32.805 71.975 33.475 ;
        RECT 72.345 32.805 72.605 33.945 ;
        RECT 72.775 33.775 74.475 33.945 ;
        RECT 75.565 33.895 76.315 34.415 ;
        RECT 77.005 34.115 77.360 34.675 ;
        RECT 77.530 33.945 77.700 34.845 ;
        RECT 77.870 34.115 78.135 34.675 ;
        RECT 78.425 34.615 79.040 35.185 ;
        RECT 78.385 33.945 78.555 34.445 ;
        RECT 72.775 32.975 73.105 33.775 ;
        RECT 73.275 32.805 73.445 33.605 ;
        RECT 73.615 32.975 73.945 33.775 ;
        RECT 74.115 32.805 74.370 33.605 ;
        RECT 74.645 32.805 76.315 33.895 ;
        RECT 77.130 33.775 78.555 33.945 ;
        RECT 77.130 33.600 77.520 33.775 ;
        RECT 78.005 32.805 78.335 33.605 ;
        RECT 78.725 33.595 79.040 34.615 ;
        RECT 78.505 32.975 79.040 33.595 ;
        RECT 79.245 34.855 79.505 35.185 ;
        RECT 79.675 34.995 80.005 35.355 ;
        RECT 80.260 34.975 81.560 35.185 ;
        RECT 79.245 33.655 79.415 34.855 ;
        RECT 80.260 34.825 80.430 34.975 ;
        RECT 79.675 34.700 80.430 34.825 ;
        RECT 79.585 34.655 80.430 34.700 ;
        RECT 79.585 34.535 79.855 34.655 ;
        RECT 79.585 33.960 79.755 34.535 ;
        RECT 79.985 34.095 80.395 34.400 ;
        RECT 80.685 34.365 80.895 34.765 ;
        RECT 80.565 34.155 80.895 34.365 ;
        RECT 81.140 34.365 81.360 34.765 ;
        RECT 81.835 34.590 82.290 35.355 ;
        RECT 83.475 34.805 83.645 35.095 ;
        RECT 83.815 34.975 84.145 35.355 ;
        RECT 83.475 34.635 84.140 34.805 ;
        RECT 81.140 34.155 81.615 34.365 ;
        RECT 81.805 34.165 82.295 34.365 ;
        RECT 79.585 33.925 79.785 33.960 ;
        RECT 81.115 33.925 82.290 33.985 ;
        RECT 79.585 33.815 82.290 33.925 ;
        RECT 83.390 33.815 83.740 34.465 ;
        RECT 79.645 33.755 81.445 33.815 ;
        RECT 81.115 33.725 81.445 33.755 ;
        RECT 79.245 32.975 79.505 33.655 ;
        RECT 79.675 32.805 79.925 33.585 ;
        RECT 80.175 33.555 81.010 33.565 ;
        RECT 81.600 33.555 81.785 33.645 ;
        RECT 80.175 33.355 81.785 33.555 ;
        RECT 80.175 32.975 80.425 33.355 ;
        RECT 81.555 33.315 81.785 33.355 ;
        RECT 82.035 33.195 82.290 33.815 ;
        RECT 83.910 33.645 84.140 34.635 ;
        RECT 80.595 32.805 80.950 33.185 ;
        RECT 81.955 32.975 82.290 33.195 ;
        RECT 83.475 33.475 84.140 33.645 ;
        RECT 83.475 32.975 83.645 33.475 ;
        RECT 83.815 32.805 84.145 33.305 ;
        RECT 84.315 32.975 84.500 35.095 ;
        RECT 84.755 34.895 85.005 35.355 ;
        RECT 85.175 34.905 85.510 35.075 ;
        RECT 85.705 34.905 86.380 35.075 ;
        RECT 85.175 34.765 85.345 34.905 ;
        RECT 84.670 33.775 84.950 34.725 ;
        RECT 85.120 34.635 85.345 34.765 ;
        RECT 85.120 33.530 85.290 34.635 ;
        RECT 85.515 34.485 86.040 34.705 ;
        RECT 85.460 33.720 85.700 34.315 ;
        RECT 85.870 33.785 86.040 34.485 ;
        RECT 86.210 34.125 86.380 34.905 ;
        RECT 86.700 34.855 87.070 35.355 ;
        RECT 87.250 34.905 87.655 35.075 ;
        RECT 87.825 34.905 88.610 35.075 ;
        RECT 87.250 34.675 87.420 34.905 ;
        RECT 86.590 34.375 87.420 34.675 ;
        RECT 87.805 34.405 88.270 34.735 ;
        RECT 86.590 34.345 86.790 34.375 ;
        RECT 86.910 34.125 87.080 34.195 ;
        RECT 86.210 33.955 87.080 34.125 ;
        RECT 86.570 33.865 87.080 33.955 ;
        RECT 85.120 33.400 85.425 33.530 ;
        RECT 85.870 33.420 86.400 33.785 ;
        RECT 84.740 32.805 85.005 33.265 ;
        RECT 85.175 32.975 85.425 33.400 ;
        RECT 86.570 33.250 86.740 33.865 ;
        RECT 85.635 33.080 86.740 33.250 ;
        RECT 86.910 32.805 87.080 33.605 ;
        RECT 87.250 33.305 87.420 34.375 ;
        RECT 87.590 33.475 87.780 34.195 ;
        RECT 87.950 33.445 88.270 34.405 ;
        RECT 88.440 34.445 88.610 34.905 ;
        RECT 88.885 34.825 89.095 35.355 ;
        RECT 89.355 34.615 89.685 35.140 ;
        RECT 89.855 34.745 90.025 35.355 ;
        RECT 90.195 34.700 90.525 35.135 ;
        RECT 90.195 34.615 90.575 34.700 ;
        RECT 89.485 34.445 89.685 34.615 ;
        RECT 90.350 34.575 90.575 34.615 ;
        RECT 90.745 34.605 91.955 35.355 ;
        RECT 88.440 34.115 89.315 34.445 ;
        RECT 89.485 34.115 90.235 34.445 ;
        RECT 87.250 32.975 87.500 33.305 ;
        RECT 88.440 33.275 88.610 34.115 ;
        RECT 89.485 33.910 89.675 34.115 ;
        RECT 90.405 33.995 90.575 34.575 ;
        RECT 90.360 33.945 90.575 33.995 ;
        RECT 88.780 33.535 89.675 33.910 ;
        RECT 90.185 33.865 90.575 33.945 ;
        RECT 90.745 33.895 91.265 34.435 ;
        RECT 91.435 34.065 91.955 34.605 ;
        RECT 87.725 33.105 88.610 33.275 ;
        RECT 88.790 32.805 89.105 33.305 ;
        RECT 89.335 32.975 89.675 33.535 ;
        RECT 89.845 32.805 90.015 33.815 ;
        RECT 90.185 33.020 90.515 33.865 ;
        RECT 90.745 32.805 91.955 33.895 ;
        RECT 13.380 32.635 92.040 32.805 ;
        RECT 13.465 31.545 14.675 32.635 ;
        RECT 13.465 30.835 13.985 31.375 ;
        RECT 14.155 31.005 14.675 31.545 ;
        RECT 14.850 31.485 15.110 32.635 ;
        RECT 15.285 31.560 15.540 32.465 ;
        RECT 15.710 31.875 16.040 32.635 ;
        RECT 16.255 31.705 16.425 32.465 ;
        RECT 13.465 30.085 14.675 30.835 ;
        RECT 14.850 30.085 15.110 30.925 ;
        RECT 15.285 30.830 15.455 31.560 ;
        RECT 15.710 31.535 16.425 31.705 ;
        RECT 17.180 31.845 17.715 32.465 ;
        RECT 15.710 31.325 15.880 31.535 ;
        RECT 15.625 30.995 15.880 31.325 ;
        RECT 15.285 30.255 15.540 30.830 ;
        RECT 15.710 30.805 15.880 30.995 ;
        RECT 16.160 30.985 16.515 31.355 ;
        RECT 17.180 30.825 17.495 31.845 ;
        RECT 17.885 31.835 18.215 32.635 ;
        RECT 18.700 31.665 19.090 31.840 ;
        RECT 17.665 31.495 19.090 31.665 ;
        RECT 19.445 31.545 21.115 32.635 ;
        RECT 17.665 30.995 17.835 31.495 ;
        RECT 15.710 30.635 16.425 30.805 ;
        RECT 15.710 30.085 16.040 30.465 ;
        RECT 16.255 30.255 16.425 30.635 ;
        RECT 17.180 30.255 17.795 30.825 ;
        RECT 18.085 30.765 18.350 31.325 ;
        RECT 18.520 30.595 18.690 31.495 ;
        RECT 18.860 30.765 19.215 31.325 ;
        RECT 19.445 30.855 20.195 31.375 ;
        RECT 20.365 31.025 21.115 31.545 ;
        RECT 21.745 31.495 22.085 32.465 ;
        RECT 22.255 31.495 22.425 32.635 ;
        RECT 22.695 31.835 22.945 32.635 ;
        RECT 23.590 31.665 23.920 32.465 ;
        RECT 24.220 31.835 24.550 32.635 ;
        RECT 24.720 31.665 25.050 32.465 ;
        RECT 22.615 31.495 25.050 31.665 ;
        RECT 21.745 30.885 21.920 31.495 ;
        RECT 22.615 31.245 22.785 31.495 ;
        RECT 22.090 31.075 22.785 31.245 ;
        RECT 22.960 31.075 23.380 31.275 ;
        RECT 23.550 31.075 23.880 31.275 ;
        RECT 24.050 31.075 24.380 31.275 ;
        RECT 17.965 30.085 18.180 30.595 ;
        RECT 18.410 30.265 18.690 30.595 ;
        RECT 18.870 30.085 19.110 30.595 ;
        RECT 19.445 30.085 21.115 30.855 ;
        RECT 21.745 30.255 22.085 30.885 ;
        RECT 22.255 30.085 22.505 30.885 ;
        RECT 22.695 30.735 23.920 30.905 ;
        RECT 22.695 30.255 23.025 30.735 ;
        RECT 23.195 30.085 23.420 30.545 ;
        RECT 23.590 30.255 23.920 30.735 ;
        RECT 24.550 30.865 24.720 31.495 ;
        RECT 26.345 31.470 26.635 32.635 ;
        RECT 26.805 32.200 32.150 32.635 ;
        RECT 32.325 32.200 37.670 32.635 ;
        RECT 37.845 32.200 43.190 32.635 ;
        RECT 24.905 31.075 25.255 31.325 ;
        RECT 24.550 30.255 25.050 30.865 ;
        RECT 26.345 30.085 26.635 30.810 ;
        RECT 28.390 30.630 28.730 31.460 ;
        RECT 30.210 30.950 30.560 32.200 ;
        RECT 33.910 30.630 34.250 31.460 ;
        RECT 35.730 30.950 36.080 32.200 ;
        RECT 39.430 30.630 39.770 31.460 ;
        RECT 41.250 30.950 41.600 32.200 ;
        RECT 44.470 31.665 44.860 31.840 ;
        RECT 45.345 31.835 45.675 32.635 ;
        RECT 45.845 31.845 46.380 32.465 ;
        RECT 44.470 31.495 45.895 31.665 ;
        RECT 44.345 30.765 44.700 31.325 ;
        RECT 26.805 30.085 32.150 30.630 ;
        RECT 32.325 30.085 37.670 30.630 ;
        RECT 37.845 30.085 43.190 30.630 ;
        RECT 44.870 30.595 45.040 31.495 ;
        RECT 45.210 30.765 45.475 31.325 ;
        RECT 45.725 30.995 45.895 31.495 ;
        RECT 46.065 30.825 46.380 31.845 ;
        RECT 46.585 31.545 48.255 32.635 ;
        RECT 44.450 30.085 44.690 30.595 ;
        RECT 44.870 30.265 45.150 30.595 ;
        RECT 45.380 30.085 45.595 30.595 ;
        RECT 45.765 30.255 46.380 30.825 ;
        RECT 46.585 30.855 47.335 31.375 ;
        RECT 47.505 31.025 48.255 31.545 ;
        RECT 48.890 32.245 49.225 32.465 ;
        RECT 50.230 32.255 50.585 32.635 ;
        RECT 48.890 31.625 49.145 32.245 ;
        RECT 49.395 32.085 49.625 32.125 ;
        RECT 50.755 32.085 51.005 32.465 ;
        RECT 49.395 31.885 51.005 32.085 ;
        RECT 49.395 31.795 49.580 31.885 ;
        RECT 50.170 31.875 51.005 31.885 ;
        RECT 51.255 31.855 51.505 32.635 ;
        RECT 51.675 31.785 51.935 32.465 ;
        RECT 49.735 31.685 50.065 31.715 ;
        RECT 49.735 31.625 51.535 31.685 ;
        RECT 48.890 31.515 51.595 31.625 ;
        RECT 48.890 31.455 50.065 31.515 ;
        RECT 51.395 31.480 51.595 31.515 ;
        RECT 48.885 31.075 49.375 31.275 ;
        RECT 49.565 31.075 50.040 31.285 ;
        RECT 46.585 30.085 48.255 30.855 ;
        RECT 48.890 30.085 49.345 30.850 ;
        RECT 49.820 30.675 50.040 31.075 ;
        RECT 50.285 31.075 50.615 31.285 ;
        RECT 50.285 30.675 50.495 31.075 ;
        RECT 50.785 31.040 51.195 31.345 ;
        RECT 51.425 30.905 51.595 31.480 ;
        RECT 51.325 30.785 51.595 30.905 ;
        RECT 50.750 30.740 51.595 30.785 ;
        RECT 50.750 30.615 51.505 30.740 ;
        RECT 50.750 30.465 50.920 30.615 ;
        RECT 51.765 30.585 51.935 31.785 ;
        RECT 52.105 31.470 52.395 32.635 ;
        RECT 52.565 31.545 53.775 32.635 ;
        RECT 52.565 30.835 53.085 31.375 ;
        RECT 53.255 31.005 53.775 31.545 ;
        RECT 54.150 31.665 54.480 32.465 ;
        RECT 54.650 31.835 54.980 32.635 ;
        RECT 55.280 31.665 55.610 32.465 ;
        RECT 56.255 31.835 56.505 32.635 ;
        RECT 54.150 31.495 56.585 31.665 ;
        RECT 56.775 31.495 56.945 32.635 ;
        RECT 57.115 31.495 57.455 32.465 ;
        RECT 53.945 31.075 54.295 31.325 ;
        RECT 54.480 30.865 54.650 31.495 ;
        RECT 54.820 31.075 55.150 31.275 ;
        RECT 55.320 31.075 55.650 31.275 ;
        RECT 55.820 31.075 56.240 31.275 ;
        RECT 56.415 31.245 56.585 31.495 ;
        RECT 56.415 31.075 57.110 31.245 ;
        RECT 49.620 30.255 50.920 30.465 ;
        RECT 51.175 30.085 51.505 30.445 ;
        RECT 51.675 30.255 51.935 30.585 ;
        RECT 52.105 30.085 52.395 30.810 ;
        RECT 52.565 30.085 53.775 30.835 ;
        RECT 54.150 30.255 54.650 30.865 ;
        RECT 55.280 30.735 56.505 30.905 ;
        RECT 57.280 30.885 57.455 31.495 ;
        RECT 55.280 30.255 55.610 30.735 ;
        RECT 55.780 30.085 56.005 30.545 ;
        RECT 56.175 30.255 56.505 30.735 ;
        RECT 56.695 30.085 56.945 30.885 ;
        RECT 57.115 30.255 57.455 30.885 ;
        RECT 57.660 31.845 58.195 32.465 ;
        RECT 57.660 30.825 57.975 31.845 ;
        RECT 58.365 31.835 58.695 32.635 ;
        RECT 60.015 31.965 60.185 32.465 ;
        RECT 60.355 32.135 60.685 32.635 ;
        RECT 59.180 31.665 59.570 31.840 ;
        RECT 60.015 31.795 60.680 31.965 ;
        RECT 58.145 31.495 59.570 31.665 ;
        RECT 58.145 30.995 58.315 31.495 ;
        RECT 57.660 30.255 58.275 30.825 ;
        RECT 58.565 30.765 58.830 31.325 ;
        RECT 59.000 30.595 59.170 31.495 ;
        RECT 59.340 30.765 59.695 31.325 ;
        RECT 59.930 30.975 60.280 31.625 ;
        RECT 60.450 30.805 60.680 31.795 ;
        RECT 60.015 30.635 60.680 30.805 ;
        RECT 58.445 30.085 58.660 30.595 ;
        RECT 58.890 30.265 59.170 30.595 ;
        RECT 59.350 30.085 59.590 30.595 ;
        RECT 60.015 30.345 60.185 30.635 ;
        RECT 60.355 30.085 60.685 30.465 ;
        RECT 60.855 30.345 61.040 32.465 ;
        RECT 61.280 32.175 61.545 32.635 ;
        RECT 61.715 32.040 61.965 32.465 ;
        RECT 62.175 32.190 63.280 32.360 ;
        RECT 61.660 31.910 61.965 32.040 ;
        RECT 61.210 30.715 61.490 31.665 ;
        RECT 61.660 30.805 61.830 31.910 ;
        RECT 62.000 31.125 62.240 31.720 ;
        RECT 62.410 31.655 62.940 32.020 ;
        RECT 62.410 30.955 62.580 31.655 ;
        RECT 63.110 31.575 63.280 32.190 ;
        RECT 63.450 31.835 63.620 32.635 ;
        RECT 63.790 32.135 64.040 32.465 ;
        RECT 64.265 32.165 65.150 32.335 ;
        RECT 63.110 31.485 63.620 31.575 ;
        RECT 61.660 30.675 61.885 30.805 ;
        RECT 62.055 30.735 62.580 30.955 ;
        RECT 62.750 31.315 63.620 31.485 ;
        RECT 61.295 30.085 61.545 30.545 ;
        RECT 61.715 30.535 61.885 30.675 ;
        RECT 62.750 30.535 62.920 31.315 ;
        RECT 63.450 31.245 63.620 31.315 ;
        RECT 63.130 31.065 63.330 31.095 ;
        RECT 63.790 31.065 63.960 32.135 ;
        RECT 64.130 31.245 64.320 31.965 ;
        RECT 63.130 30.765 63.960 31.065 ;
        RECT 64.490 31.035 64.810 31.995 ;
        RECT 61.715 30.365 62.050 30.535 ;
        RECT 62.245 30.365 62.920 30.535 ;
        RECT 63.240 30.085 63.610 30.585 ;
        RECT 63.790 30.535 63.960 30.765 ;
        RECT 64.345 30.705 64.810 31.035 ;
        RECT 64.980 31.325 65.150 32.165 ;
        RECT 65.330 32.135 65.645 32.635 ;
        RECT 65.875 31.905 66.215 32.465 ;
        RECT 65.320 31.530 66.215 31.905 ;
        RECT 66.385 31.625 66.555 32.635 ;
        RECT 66.025 31.325 66.215 31.530 ;
        RECT 66.725 31.575 67.055 32.420 ;
        RECT 67.320 31.845 67.855 32.465 ;
        RECT 66.725 31.495 67.115 31.575 ;
        RECT 66.900 31.445 67.115 31.495 ;
        RECT 64.980 30.995 65.855 31.325 ;
        RECT 66.025 30.995 66.775 31.325 ;
        RECT 64.980 30.535 65.150 30.995 ;
        RECT 66.025 30.825 66.225 30.995 ;
        RECT 66.945 30.865 67.115 31.445 ;
        RECT 66.890 30.825 67.115 30.865 ;
        RECT 63.790 30.365 64.195 30.535 ;
        RECT 64.365 30.365 65.150 30.535 ;
        RECT 65.425 30.085 65.635 30.615 ;
        RECT 65.895 30.300 66.225 30.825 ;
        RECT 66.735 30.740 67.115 30.825 ;
        RECT 67.320 30.825 67.635 31.845 ;
        RECT 68.025 31.835 68.355 32.635 ;
        RECT 69.675 31.965 69.845 32.465 ;
        RECT 70.015 32.135 70.345 32.635 ;
        RECT 68.840 31.665 69.230 31.840 ;
        RECT 69.675 31.795 70.340 31.965 ;
        RECT 67.805 31.495 69.230 31.665 ;
        RECT 67.805 30.995 67.975 31.495 ;
        RECT 66.395 30.085 66.565 30.695 ;
        RECT 66.735 30.305 67.065 30.740 ;
        RECT 67.320 30.255 67.935 30.825 ;
        RECT 68.225 30.765 68.490 31.325 ;
        RECT 68.660 30.595 68.830 31.495 ;
        RECT 69.000 30.765 69.355 31.325 ;
        RECT 69.590 30.975 69.940 31.625 ;
        RECT 70.110 30.805 70.340 31.795 ;
        RECT 69.675 30.635 70.340 30.805 ;
        RECT 68.105 30.085 68.320 30.595 ;
        RECT 68.550 30.265 68.830 30.595 ;
        RECT 69.010 30.085 69.250 30.595 ;
        RECT 69.675 30.345 69.845 30.635 ;
        RECT 70.015 30.085 70.345 30.465 ;
        RECT 70.515 30.345 70.700 32.465 ;
        RECT 70.940 32.175 71.205 32.635 ;
        RECT 71.375 32.040 71.625 32.465 ;
        RECT 71.835 32.190 72.940 32.360 ;
        RECT 71.320 31.910 71.625 32.040 ;
        RECT 70.870 30.715 71.150 31.665 ;
        RECT 71.320 30.805 71.490 31.910 ;
        RECT 71.660 31.125 71.900 31.720 ;
        RECT 72.070 31.655 72.600 32.020 ;
        RECT 72.070 30.955 72.240 31.655 ;
        RECT 72.770 31.575 72.940 32.190 ;
        RECT 73.110 31.835 73.280 32.635 ;
        RECT 73.450 32.135 73.700 32.465 ;
        RECT 73.925 32.165 74.810 32.335 ;
        RECT 72.770 31.485 73.280 31.575 ;
        RECT 71.320 30.675 71.545 30.805 ;
        RECT 71.715 30.735 72.240 30.955 ;
        RECT 72.410 31.315 73.280 31.485 ;
        RECT 70.955 30.085 71.205 30.545 ;
        RECT 71.375 30.535 71.545 30.675 ;
        RECT 72.410 30.535 72.580 31.315 ;
        RECT 73.110 31.245 73.280 31.315 ;
        RECT 72.790 31.065 72.990 31.095 ;
        RECT 73.450 31.065 73.620 32.135 ;
        RECT 73.790 31.245 73.980 31.965 ;
        RECT 72.790 30.765 73.620 31.065 ;
        RECT 74.150 31.035 74.470 31.995 ;
        RECT 71.375 30.365 71.710 30.535 ;
        RECT 71.905 30.365 72.580 30.535 ;
        RECT 72.900 30.085 73.270 30.585 ;
        RECT 73.450 30.535 73.620 30.765 ;
        RECT 74.005 30.705 74.470 31.035 ;
        RECT 74.640 31.325 74.810 32.165 ;
        RECT 74.990 32.135 75.305 32.635 ;
        RECT 75.535 31.905 75.875 32.465 ;
        RECT 74.980 31.530 75.875 31.905 ;
        RECT 76.045 31.625 76.215 32.635 ;
        RECT 75.685 31.325 75.875 31.530 ;
        RECT 76.385 31.575 76.715 32.420 ;
        RECT 76.385 31.495 76.775 31.575 ;
        RECT 76.560 31.445 76.775 31.495 ;
        RECT 77.865 31.470 78.155 32.635 ;
        RECT 78.970 31.665 79.360 31.840 ;
        RECT 79.845 31.835 80.175 32.635 ;
        RECT 80.345 31.845 80.880 32.465 ;
        RECT 81.085 32.200 86.430 32.635 ;
        RECT 78.970 31.495 80.395 31.665 ;
        RECT 74.640 30.995 75.515 31.325 ;
        RECT 75.685 30.995 76.435 31.325 ;
        RECT 74.640 30.535 74.810 30.995 ;
        RECT 75.685 30.825 75.885 30.995 ;
        RECT 76.605 30.865 76.775 31.445 ;
        RECT 76.550 30.825 76.775 30.865 ;
        RECT 73.450 30.365 73.855 30.535 ;
        RECT 74.025 30.365 74.810 30.535 ;
        RECT 75.085 30.085 75.295 30.615 ;
        RECT 75.555 30.300 75.885 30.825 ;
        RECT 76.395 30.740 76.775 30.825 ;
        RECT 76.055 30.085 76.225 30.695 ;
        RECT 76.395 30.305 76.725 30.740 ;
        RECT 77.865 30.085 78.155 30.810 ;
        RECT 78.845 30.765 79.200 31.325 ;
        RECT 79.370 30.595 79.540 31.495 ;
        RECT 79.710 30.765 79.975 31.325 ;
        RECT 80.225 30.995 80.395 31.495 ;
        RECT 80.565 30.825 80.880 31.845 ;
        RECT 78.950 30.085 79.190 30.595 ;
        RECT 79.370 30.265 79.650 30.595 ;
        RECT 79.880 30.085 80.095 30.595 ;
        RECT 80.265 30.255 80.880 30.825 ;
        RECT 82.670 30.630 83.010 31.460 ;
        RECT 84.490 30.950 84.840 32.200 ;
        RECT 86.605 31.545 88.275 32.635 ;
        RECT 86.605 30.855 87.355 31.375 ;
        RECT 87.525 31.025 88.275 31.545 ;
        RECT 88.995 31.705 89.165 32.465 ;
        RECT 89.380 31.875 89.710 32.635 ;
        RECT 88.995 31.535 89.710 31.705 ;
        RECT 89.880 31.560 90.135 32.465 ;
        RECT 88.905 30.985 89.260 31.355 ;
        RECT 89.540 31.325 89.710 31.535 ;
        RECT 89.540 30.995 89.795 31.325 ;
        RECT 81.085 30.085 86.430 30.630 ;
        RECT 86.605 30.085 88.275 30.855 ;
        RECT 89.540 30.805 89.710 30.995 ;
        RECT 89.965 30.830 90.135 31.560 ;
        RECT 90.310 31.485 90.570 32.635 ;
        RECT 90.745 31.545 91.955 32.635 ;
        RECT 90.745 31.005 91.265 31.545 ;
        RECT 88.995 30.635 89.710 30.805 ;
        RECT 88.995 30.255 89.165 30.635 ;
        RECT 89.380 30.085 89.710 30.465 ;
        RECT 89.880 30.255 90.135 30.830 ;
        RECT 90.310 30.085 90.570 30.925 ;
        RECT 91.435 30.835 91.955 31.375 ;
        RECT 90.745 30.085 91.955 30.835 ;
        RECT 13.380 29.915 92.040 30.085 ;
        RECT 13.465 29.165 14.675 29.915 ;
        RECT 13.465 28.625 13.985 29.165 ;
        RECT 15.305 29.115 15.645 29.745 ;
        RECT 15.815 29.115 16.065 29.915 ;
        RECT 16.255 29.265 16.585 29.745 ;
        RECT 16.755 29.455 16.980 29.915 ;
        RECT 17.150 29.265 17.480 29.745 ;
        RECT 14.155 28.455 14.675 28.995 ;
        RECT 13.465 27.365 14.675 28.455 ;
        RECT 15.305 28.505 15.480 29.115 ;
        RECT 16.255 29.095 17.480 29.265 ;
        RECT 18.110 29.135 18.610 29.745 ;
        RECT 19.075 29.365 19.245 29.655 ;
        RECT 19.415 29.535 19.745 29.915 ;
        RECT 19.075 29.195 19.740 29.365 ;
        RECT 15.650 28.755 16.345 28.925 ;
        RECT 16.175 28.505 16.345 28.755 ;
        RECT 16.520 28.725 16.940 28.925 ;
        RECT 17.110 28.725 17.440 28.925 ;
        RECT 17.610 28.725 17.940 28.925 ;
        RECT 18.110 28.505 18.280 29.135 ;
        RECT 18.465 28.675 18.815 28.925 ;
        RECT 15.305 27.535 15.645 28.505 ;
        RECT 15.815 27.365 15.985 28.505 ;
        RECT 16.175 28.335 18.610 28.505 ;
        RECT 18.990 28.375 19.340 29.025 ;
        RECT 16.255 27.365 16.505 28.165 ;
        RECT 17.150 27.535 17.480 28.335 ;
        RECT 17.780 27.365 18.110 28.165 ;
        RECT 18.280 27.535 18.610 28.335 ;
        RECT 19.510 28.205 19.740 29.195 ;
        RECT 19.075 28.035 19.740 28.205 ;
        RECT 19.075 27.535 19.245 28.035 ;
        RECT 19.415 27.365 19.745 27.865 ;
        RECT 19.915 27.535 20.100 29.655 ;
        RECT 20.355 29.455 20.605 29.915 ;
        RECT 20.775 29.465 21.110 29.635 ;
        RECT 21.305 29.465 21.980 29.635 ;
        RECT 20.775 29.325 20.945 29.465 ;
        RECT 20.270 28.335 20.550 29.285 ;
        RECT 20.720 29.195 20.945 29.325 ;
        RECT 20.720 28.090 20.890 29.195 ;
        RECT 21.115 29.045 21.640 29.265 ;
        RECT 21.060 28.280 21.300 28.875 ;
        RECT 21.470 28.345 21.640 29.045 ;
        RECT 21.810 28.685 21.980 29.465 ;
        RECT 22.300 29.415 22.670 29.915 ;
        RECT 22.850 29.465 23.255 29.635 ;
        RECT 23.425 29.465 24.210 29.635 ;
        RECT 22.850 29.235 23.020 29.465 ;
        RECT 22.190 28.935 23.020 29.235 ;
        RECT 23.405 28.965 23.870 29.295 ;
        RECT 22.190 28.905 22.390 28.935 ;
        RECT 22.510 28.685 22.680 28.755 ;
        RECT 21.810 28.515 22.680 28.685 ;
        RECT 22.170 28.425 22.680 28.515 ;
        RECT 20.720 27.960 21.025 28.090 ;
        RECT 21.470 27.980 22.000 28.345 ;
        RECT 20.340 27.365 20.605 27.825 ;
        RECT 20.775 27.535 21.025 27.960 ;
        RECT 22.170 27.810 22.340 28.425 ;
        RECT 21.235 27.640 22.340 27.810 ;
        RECT 22.510 27.365 22.680 28.165 ;
        RECT 22.850 27.865 23.020 28.935 ;
        RECT 23.190 28.035 23.380 28.755 ;
        RECT 23.550 28.005 23.870 28.965 ;
        RECT 24.040 29.005 24.210 29.465 ;
        RECT 24.485 29.385 24.695 29.915 ;
        RECT 24.955 29.175 25.285 29.700 ;
        RECT 25.455 29.305 25.625 29.915 ;
        RECT 25.795 29.260 26.125 29.695 ;
        RECT 25.795 29.175 26.175 29.260 ;
        RECT 25.085 29.005 25.285 29.175 ;
        RECT 25.950 29.135 26.175 29.175 ;
        RECT 24.040 28.675 24.915 29.005 ;
        RECT 25.085 28.675 25.835 29.005 ;
        RECT 22.850 27.535 23.100 27.865 ;
        RECT 24.040 27.835 24.210 28.675 ;
        RECT 25.085 28.470 25.275 28.675 ;
        RECT 26.005 28.555 26.175 29.135 ;
        RECT 25.960 28.505 26.175 28.555 ;
        RECT 24.380 28.095 25.275 28.470 ;
        RECT 25.785 28.425 26.175 28.505 ;
        RECT 26.380 29.175 26.995 29.745 ;
        RECT 27.165 29.405 27.380 29.915 ;
        RECT 27.610 29.405 27.890 29.735 ;
        RECT 28.070 29.405 28.310 29.915 ;
        RECT 23.325 27.665 24.210 27.835 ;
        RECT 24.390 27.365 24.705 27.865 ;
        RECT 24.935 27.535 25.275 28.095 ;
        RECT 25.445 27.365 25.615 28.375 ;
        RECT 25.785 27.580 26.115 28.425 ;
        RECT 26.380 28.155 26.695 29.175 ;
        RECT 26.865 28.505 27.035 29.005 ;
        RECT 27.285 28.675 27.550 29.235 ;
        RECT 27.720 28.505 27.890 29.405 ;
        RECT 28.060 28.675 28.415 29.235 ;
        RECT 29.105 29.115 29.445 29.745 ;
        RECT 29.615 29.115 29.865 29.915 ;
        RECT 30.055 29.265 30.385 29.745 ;
        RECT 30.555 29.455 30.780 29.915 ;
        RECT 30.950 29.265 31.280 29.745 ;
        RECT 29.105 28.505 29.280 29.115 ;
        RECT 30.055 29.095 31.280 29.265 ;
        RECT 31.910 29.135 32.410 29.745 ;
        RECT 33.450 29.135 33.950 29.745 ;
        RECT 29.450 28.755 30.145 28.925 ;
        RECT 29.975 28.505 30.145 28.755 ;
        RECT 30.320 28.725 30.740 28.925 ;
        RECT 30.910 28.725 31.240 28.925 ;
        RECT 31.410 28.725 31.740 28.925 ;
        RECT 31.910 28.505 32.080 29.135 ;
        RECT 32.265 28.675 32.615 28.925 ;
        RECT 33.245 28.675 33.595 28.925 ;
        RECT 33.780 28.505 33.950 29.135 ;
        RECT 34.580 29.265 34.910 29.745 ;
        RECT 35.080 29.455 35.305 29.915 ;
        RECT 35.475 29.265 35.805 29.745 ;
        RECT 34.580 29.095 35.805 29.265 ;
        RECT 35.995 29.115 36.245 29.915 ;
        RECT 36.415 29.115 36.755 29.745 ;
        RECT 37.090 29.405 37.330 29.915 ;
        RECT 37.510 29.405 37.790 29.735 ;
        RECT 38.020 29.405 38.235 29.915 ;
        RECT 34.120 28.725 34.450 28.925 ;
        RECT 34.620 28.725 34.950 28.925 ;
        RECT 35.120 28.725 35.540 28.925 ;
        RECT 35.715 28.755 36.410 28.925 ;
        RECT 35.715 28.505 35.885 28.755 ;
        RECT 36.580 28.505 36.755 29.115 ;
        RECT 36.985 28.675 37.340 29.235 ;
        RECT 37.510 28.505 37.680 29.405 ;
        RECT 37.850 28.675 38.115 29.235 ;
        RECT 38.405 29.175 39.020 29.745 ;
        RECT 39.225 29.190 39.515 29.915 ;
        RECT 38.365 28.505 38.535 29.005 ;
        RECT 26.865 28.335 28.290 28.505 ;
        RECT 26.380 27.535 26.915 28.155 ;
        RECT 27.085 27.365 27.415 28.165 ;
        RECT 27.900 28.160 28.290 28.335 ;
        RECT 29.105 27.535 29.445 28.505 ;
        RECT 29.615 27.365 29.785 28.505 ;
        RECT 29.975 28.335 32.410 28.505 ;
        RECT 30.055 27.365 30.305 28.165 ;
        RECT 30.950 27.535 31.280 28.335 ;
        RECT 31.580 27.365 31.910 28.165 ;
        RECT 32.080 27.535 32.410 28.335 ;
        RECT 33.450 28.335 35.885 28.505 ;
        RECT 33.450 27.535 33.780 28.335 ;
        RECT 33.950 27.365 34.280 28.165 ;
        RECT 34.580 27.535 34.910 28.335 ;
        RECT 35.555 27.365 35.805 28.165 ;
        RECT 36.075 27.365 36.245 28.505 ;
        RECT 36.415 27.535 36.755 28.505 ;
        RECT 37.110 28.335 38.535 28.505 ;
        RECT 37.110 28.160 37.500 28.335 ;
        RECT 37.985 27.365 38.315 28.165 ;
        RECT 38.705 28.155 39.020 29.175 ;
        RECT 39.685 29.145 42.275 29.915 ;
        RECT 42.535 29.365 42.705 29.655 ;
        RECT 42.875 29.535 43.205 29.915 ;
        RECT 42.535 29.195 43.200 29.365 ;
        RECT 39.685 28.625 40.895 29.145 ;
        RECT 38.485 27.535 39.020 28.155 ;
        RECT 39.225 27.365 39.515 28.530 ;
        RECT 41.065 28.455 42.275 28.975 ;
        RECT 39.685 27.365 42.275 28.455 ;
        RECT 42.450 28.375 42.800 29.025 ;
        RECT 42.970 28.205 43.200 29.195 ;
        RECT 42.535 28.035 43.200 28.205 ;
        RECT 42.535 27.535 42.705 28.035 ;
        RECT 42.875 27.365 43.205 27.865 ;
        RECT 43.375 27.535 43.560 29.655 ;
        RECT 43.815 29.455 44.065 29.915 ;
        RECT 44.235 29.465 44.570 29.635 ;
        RECT 44.765 29.465 45.440 29.635 ;
        RECT 44.235 29.325 44.405 29.465 ;
        RECT 43.730 28.335 44.010 29.285 ;
        RECT 44.180 29.195 44.405 29.325 ;
        RECT 44.180 28.090 44.350 29.195 ;
        RECT 44.575 29.045 45.100 29.265 ;
        RECT 44.520 28.280 44.760 28.875 ;
        RECT 44.930 28.345 45.100 29.045 ;
        RECT 45.270 28.685 45.440 29.465 ;
        RECT 45.760 29.415 46.130 29.915 ;
        RECT 46.310 29.465 46.715 29.635 ;
        RECT 46.885 29.465 47.670 29.635 ;
        RECT 46.310 29.235 46.480 29.465 ;
        RECT 45.650 28.935 46.480 29.235 ;
        RECT 46.865 28.965 47.330 29.295 ;
        RECT 45.650 28.905 45.850 28.935 ;
        RECT 45.970 28.685 46.140 28.755 ;
        RECT 45.270 28.515 46.140 28.685 ;
        RECT 45.630 28.425 46.140 28.515 ;
        RECT 44.180 27.960 44.485 28.090 ;
        RECT 44.930 27.980 45.460 28.345 ;
        RECT 43.800 27.365 44.065 27.825 ;
        RECT 44.235 27.535 44.485 27.960 ;
        RECT 45.630 27.810 45.800 28.425 ;
        RECT 44.695 27.640 45.800 27.810 ;
        RECT 45.970 27.365 46.140 28.165 ;
        RECT 46.310 27.865 46.480 28.935 ;
        RECT 46.650 28.035 46.840 28.755 ;
        RECT 47.010 28.005 47.330 28.965 ;
        RECT 47.500 29.005 47.670 29.465 ;
        RECT 47.945 29.385 48.155 29.915 ;
        RECT 48.415 29.175 48.745 29.700 ;
        RECT 48.915 29.305 49.085 29.915 ;
        RECT 49.255 29.260 49.585 29.695 ;
        RECT 49.255 29.175 49.635 29.260 ;
        RECT 48.545 29.005 48.745 29.175 ;
        RECT 49.410 29.135 49.635 29.175 ;
        RECT 47.500 28.675 48.375 29.005 ;
        RECT 48.545 28.675 49.295 29.005 ;
        RECT 46.310 27.535 46.560 27.865 ;
        RECT 47.500 27.835 47.670 28.675 ;
        RECT 48.545 28.470 48.735 28.675 ;
        RECT 49.465 28.555 49.635 29.135 ;
        RECT 49.805 29.165 51.015 29.915 ;
        RECT 51.275 29.365 51.445 29.655 ;
        RECT 51.615 29.535 51.945 29.915 ;
        RECT 51.275 29.195 51.940 29.365 ;
        RECT 49.805 28.625 50.325 29.165 ;
        RECT 49.420 28.505 49.635 28.555 ;
        RECT 47.840 28.095 48.735 28.470 ;
        RECT 49.245 28.425 49.635 28.505 ;
        RECT 50.495 28.455 51.015 28.995 ;
        RECT 46.785 27.665 47.670 27.835 ;
        RECT 47.850 27.365 48.165 27.865 ;
        RECT 48.395 27.535 48.735 28.095 ;
        RECT 48.905 27.365 49.075 28.375 ;
        RECT 49.245 27.580 49.575 28.425 ;
        RECT 49.805 27.365 51.015 28.455 ;
        RECT 51.190 28.375 51.540 29.025 ;
        RECT 51.710 28.205 51.940 29.195 ;
        RECT 51.275 28.035 51.940 28.205 ;
        RECT 51.275 27.535 51.445 28.035 ;
        RECT 51.615 27.365 51.945 27.865 ;
        RECT 52.115 27.535 52.300 29.655 ;
        RECT 52.555 29.455 52.805 29.915 ;
        RECT 52.975 29.465 53.310 29.635 ;
        RECT 53.505 29.465 54.180 29.635 ;
        RECT 52.975 29.325 53.145 29.465 ;
        RECT 52.470 28.335 52.750 29.285 ;
        RECT 52.920 29.195 53.145 29.325 ;
        RECT 52.920 28.090 53.090 29.195 ;
        RECT 53.315 29.045 53.840 29.265 ;
        RECT 53.260 28.280 53.500 28.875 ;
        RECT 53.670 28.345 53.840 29.045 ;
        RECT 54.010 28.685 54.180 29.465 ;
        RECT 54.500 29.415 54.870 29.915 ;
        RECT 55.050 29.465 55.455 29.635 ;
        RECT 55.625 29.465 56.410 29.635 ;
        RECT 55.050 29.235 55.220 29.465 ;
        RECT 54.390 28.935 55.220 29.235 ;
        RECT 55.605 28.965 56.070 29.295 ;
        RECT 54.390 28.905 54.590 28.935 ;
        RECT 54.710 28.685 54.880 28.755 ;
        RECT 54.010 28.515 54.880 28.685 ;
        RECT 54.370 28.425 54.880 28.515 ;
        RECT 52.920 27.960 53.225 28.090 ;
        RECT 53.670 27.980 54.200 28.345 ;
        RECT 52.540 27.365 52.805 27.825 ;
        RECT 52.975 27.535 53.225 27.960 ;
        RECT 54.370 27.810 54.540 28.425 ;
        RECT 53.435 27.640 54.540 27.810 ;
        RECT 54.710 27.365 54.880 28.165 ;
        RECT 55.050 27.865 55.220 28.935 ;
        RECT 55.390 28.035 55.580 28.755 ;
        RECT 55.750 28.005 56.070 28.965 ;
        RECT 56.240 29.005 56.410 29.465 ;
        RECT 56.685 29.385 56.895 29.915 ;
        RECT 57.155 29.175 57.485 29.700 ;
        RECT 57.655 29.305 57.825 29.915 ;
        RECT 57.995 29.260 58.325 29.695 ;
        RECT 57.995 29.175 58.375 29.260 ;
        RECT 57.285 29.005 57.485 29.175 ;
        RECT 58.150 29.135 58.375 29.175 ;
        RECT 56.240 28.675 57.115 29.005 ;
        RECT 57.285 28.675 58.035 29.005 ;
        RECT 55.050 27.535 55.300 27.865 ;
        RECT 56.240 27.835 56.410 28.675 ;
        RECT 57.285 28.470 57.475 28.675 ;
        RECT 58.205 28.555 58.375 29.135 ;
        RECT 58.160 28.505 58.375 28.555 ;
        RECT 56.580 28.095 57.475 28.470 ;
        RECT 57.985 28.425 58.375 28.505 ;
        RECT 59.005 29.115 59.345 29.745 ;
        RECT 59.515 29.115 59.765 29.915 ;
        RECT 59.955 29.265 60.285 29.745 ;
        RECT 60.455 29.455 60.680 29.915 ;
        RECT 60.850 29.265 61.180 29.745 ;
        RECT 59.005 28.505 59.180 29.115 ;
        RECT 59.955 29.095 61.180 29.265 ;
        RECT 61.810 29.135 62.310 29.745 ;
        RECT 62.720 29.175 63.335 29.745 ;
        RECT 63.505 29.405 63.720 29.915 ;
        RECT 63.950 29.405 64.230 29.735 ;
        RECT 64.410 29.405 64.650 29.915 ;
        RECT 59.350 28.755 60.045 28.925 ;
        RECT 59.875 28.505 60.045 28.755 ;
        RECT 60.220 28.725 60.640 28.925 ;
        RECT 60.810 28.725 61.140 28.925 ;
        RECT 61.310 28.725 61.640 28.925 ;
        RECT 61.810 28.505 61.980 29.135 ;
        RECT 62.165 28.675 62.515 28.925 ;
        RECT 55.525 27.665 56.410 27.835 ;
        RECT 56.590 27.365 56.905 27.865 ;
        RECT 57.135 27.535 57.475 28.095 ;
        RECT 57.645 27.365 57.815 28.375 ;
        RECT 57.985 27.580 58.315 28.425 ;
        RECT 59.005 27.535 59.345 28.505 ;
        RECT 59.515 27.365 59.685 28.505 ;
        RECT 59.875 28.335 62.310 28.505 ;
        RECT 59.955 27.365 60.205 28.165 ;
        RECT 60.850 27.535 61.180 28.335 ;
        RECT 61.480 27.365 61.810 28.165 ;
        RECT 61.980 27.535 62.310 28.335 ;
        RECT 62.720 28.155 63.035 29.175 ;
        RECT 63.205 28.505 63.375 29.005 ;
        RECT 63.625 28.675 63.890 29.235 ;
        RECT 64.060 28.505 64.230 29.405 ;
        RECT 64.400 28.675 64.755 29.235 ;
        RECT 64.985 29.190 65.275 29.915 ;
        RECT 66.365 29.415 66.625 29.745 ;
        RECT 66.795 29.555 67.125 29.915 ;
        RECT 67.380 29.535 68.680 29.745 ;
        RECT 66.365 29.405 66.595 29.415 ;
        RECT 63.205 28.335 64.630 28.505 ;
        RECT 62.720 27.535 63.255 28.155 ;
        RECT 63.425 27.365 63.755 28.165 ;
        RECT 64.240 28.160 64.630 28.335 ;
        RECT 64.985 27.365 65.275 28.530 ;
        RECT 66.365 28.215 66.535 29.405 ;
        RECT 67.380 29.385 67.550 29.535 ;
        RECT 66.795 29.260 67.550 29.385 ;
        RECT 66.705 29.215 67.550 29.260 ;
        RECT 66.705 29.095 66.975 29.215 ;
        RECT 66.705 28.520 66.875 29.095 ;
        RECT 67.105 28.655 67.515 28.960 ;
        RECT 67.805 28.925 68.015 29.325 ;
        RECT 67.685 28.715 68.015 28.925 ;
        RECT 68.260 28.925 68.480 29.325 ;
        RECT 68.955 29.150 69.410 29.915 ;
        RECT 69.790 29.135 70.290 29.745 ;
        RECT 68.260 28.715 68.735 28.925 ;
        RECT 68.925 28.725 69.415 28.925 ;
        RECT 69.585 28.675 69.935 28.925 ;
        RECT 66.705 28.485 66.905 28.520 ;
        RECT 68.235 28.485 69.410 28.545 ;
        RECT 70.120 28.505 70.290 29.135 ;
        RECT 70.920 29.265 71.250 29.745 ;
        RECT 71.420 29.455 71.645 29.915 ;
        RECT 71.815 29.265 72.145 29.745 ;
        RECT 70.920 29.095 72.145 29.265 ;
        RECT 72.335 29.115 72.585 29.915 ;
        RECT 72.755 29.115 73.095 29.745 ;
        RECT 70.460 28.725 70.790 28.925 ;
        RECT 70.960 28.725 71.290 28.925 ;
        RECT 71.460 28.725 71.880 28.925 ;
        RECT 72.055 28.755 72.750 28.925 ;
        RECT 72.055 28.505 72.225 28.755 ;
        RECT 72.920 28.505 73.095 29.115 ;
        RECT 73.265 29.145 74.935 29.915 ;
        RECT 75.655 29.365 75.825 29.655 ;
        RECT 75.995 29.535 76.325 29.915 ;
        RECT 75.655 29.195 76.320 29.365 ;
        RECT 73.265 28.625 74.015 29.145 ;
        RECT 66.705 28.375 69.410 28.485 ;
        RECT 66.765 28.315 68.565 28.375 ;
        RECT 68.235 28.285 68.565 28.315 ;
        RECT 66.365 27.535 66.625 28.215 ;
        RECT 66.795 27.365 67.045 28.145 ;
        RECT 67.295 28.115 68.130 28.125 ;
        RECT 68.720 28.115 68.905 28.205 ;
        RECT 67.295 27.915 68.905 28.115 ;
        RECT 67.295 27.535 67.545 27.915 ;
        RECT 68.675 27.875 68.905 27.915 ;
        RECT 69.155 27.755 69.410 28.375 ;
        RECT 67.715 27.365 68.070 27.745 ;
        RECT 69.075 27.535 69.410 27.755 ;
        RECT 69.790 28.335 72.225 28.505 ;
        RECT 69.790 27.535 70.120 28.335 ;
        RECT 70.290 27.365 70.620 28.165 ;
        RECT 70.920 27.535 71.250 28.335 ;
        RECT 71.895 27.365 72.145 28.165 ;
        RECT 72.415 27.365 72.585 28.505 ;
        RECT 72.755 27.535 73.095 28.505 ;
        RECT 74.185 28.455 74.935 28.975 ;
        RECT 73.265 27.365 74.935 28.455 ;
        RECT 75.570 28.375 75.920 29.025 ;
        RECT 76.090 28.205 76.320 29.195 ;
        RECT 75.655 28.035 76.320 28.205 ;
        RECT 75.655 27.535 75.825 28.035 ;
        RECT 75.995 27.365 76.325 27.865 ;
        RECT 76.495 27.535 76.680 29.655 ;
        RECT 76.935 29.455 77.185 29.915 ;
        RECT 77.355 29.465 77.690 29.635 ;
        RECT 77.885 29.465 78.560 29.635 ;
        RECT 77.355 29.325 77.525 29.465 ;
        RECT 76.850 28.335 77.130 29.285 ;
        RECT 77.300 29.195 77.525 29.325 ;
        RECT 77.300 28.090 77.470 29.195 ;
        RECT 77.695 29.045 78.220 29.265 ;
        RECT 77.640 28.280 77.880 28.875 ;
        RECT 78.050 28.345 78.220 29.045 ;
        RECT 78.390 28.685 78.560 29.465 ;
        RECT 78.880 29.415 79.250 29.915 ;
        RECT 79.430 29.465 79.835 29.635 ;
        RECT 80.005 29.465 80.790 29.635 ;
        RECT 79.430 29.235 79.600 29.465 ;
        RECT 78.770 28.935 79.600 29.235 ;
        RECT 79.985 28.965 80.450 29.295 ;
        RECT 78.770 28.905 78.970 28.935 ;
        RECT 79.090 28.685 79.260 28.755 ;
        RECT 78.390 28.515 79.260 28.685 ;
        RECT 78.750 28.425 79.260 28.515 ;
        RECT 77.300 27.960 77.605 28.090 ;
        RECT 78.050 27.980 78.580 28.345 ;
        RECT 76.920 27.365 77.185 27.825 ;
        RECT 77.355 27.535 77.605 27.960 ;
        RECT 78.750 27.810 78.920 28.425 ;
        RECT 77.815 27.640 78.920 27.810 ;
        RECT 79.090 27.365 79.260 28.165 ;
        RECT 79.430 27.865 79.600 28.935 ;
        RECT 79.770 28.035 79.960 28.755 ;
        RECT 80.130 28.005 80.450 28.965 ;
        RECT 80.620 29.005 80.790 29.465 ;
        RECT 81.065 29.385 81.275 29.915 ;
        RECT 81.535 29.175 81.865 29.700 ;
        RECT 82.035 29.305 82.205 29.915 ;
        RECT 82.375 29.260 82.705 29.695 ;
        RECT 82.925 29.415 83.185 29.745 ;
        RECT 83.355 29.555 83.685 29.915 ;
        RECT 83.940 29.535 85.240 29.745 ;
        RECT 82.375 29.175 82.755 29.260 ;
        RECT 81.665 29.005 81.865 29.175 ;
        RECT 82.530 29.135 82.755 29.175 ;
        RECT 80.620 28.675 81.495 29.005 ;
        RECT 81.665 28.675 82.415 29.005 ;
        RECT 79.430 27.535 79.680 27.865 ;
        RECT 80.620 27.835 80.790 28.675 ;
        RECT 81.665 28.470 81.855 28.675 ;
        RECT 82.585 28.555 82.755 29.135 ;
        RECT 82.540 28.505 82.755 28.555 ;
        RECT 80.960 28.095 81.855 28.470 ;
        RECT 82.365 28.425 82.755 28.505 ;
        RECT 79.905 27.665 80.790 27.835 ;
        RECT 80.970 27.365 81.285 27.865 ;
        RECT 81.515 27.535 81.855 28.095 ;
        RECT 82.025 27.365 82.195 28.375 ;
        RECT 82.365 27.580 82.695 28.425 ;
        RECT 82.925 28.215 83.095 29.415 ;
        RECT 83.940 29.385 84.110 29.535 ;
        RECT 83.355 29.260 84.110 29.385 ;
        RECT 83.265 29.215 84.110 29.260 ;
        RECT 83.265 29.095 83.535 29.215 ;
        RECT 83.265 28.520 83.435 29.095 ;
        RECT 83.665 28.655 84.075 28.960 ;
        RECT 84.365 28.925 84.575 29.325 ;
        RECT 84.245 28.715 84.575 28.925 ;
        RECT 84.820 28.925 85.040 29.325 ;
        RECT 85.515 29.150 85.970 29.915 ;
        RECT 86.145 29.145 89.655 29.915 ;
        RECT 90.745 29.165 91.955 29.915 ;
        RECT 84.820 28.715 85.295 28.925 ;
        RECT 85.485 28.725 85.975 28.925 ;
        RECT 86.145 28.625 87.795 29.145 ;
        RECT 83.265 28.485 83.465 28.520 ;
        RECT 84.795 28.485 85.970 28.545 ;
        RECT 83.265 28.375 85.970 28.485 ;
        RECT 87.965 28.455 89.655 28.975 ;
        RECT 83.325 28.315 85.125 28.375 ;
        RECT 84.795 28.285 85.125 28.315 ;
        RECT 82.925 27.535 83.185 28.215 ;
        RECT 83.355 27.365 83.605 28.145 ;
        RECT 83.855 28.115 84.690 28.125 ;
        RECT 85.280 28.115 85.465 28.205 ;
        RECT 83.855 27.915 85.465 28.115 ;
        RECT 83.855 27.535 84.105 27.915 ;
        RECT 85.235 27.875 85.465 27.915 ;
        RECT 85.715 27.755 85.970 28.375 ;
        RECT 84.275 27.365 84.630 27.745 ;
        RECT 85.635 27.535 85.970 27.755 ;
        RECT 86.145 27.365 89.655 28.455 ;
        RECT 90.745 28.455 91.265 28.995 ;
        RECT 91.435 28.625 91.955 29.165 ;
        RECT 90.745 27.365 91.955 28.455 ;
        RECT 13.380 27.195 92.040 27.365 ;
        RECT 13.465 26.105 14.675 27.195 ;
        RECT 14.935 26.525 15.105 27.025 ;
        RECT 15.275 26.695 15.605 27.195 ;
        RECT 14.935 26.355 15.600 26.525 ;
        RECT 13.465 25.395 13.985 25.935 ;
        RECT 14.155 25.565 14.675 26.105 ;
        RECT 14.850 25.535 15.200 26.185 ;
        RECT 13.465 24.645 14.675 25.395 ;
        RECT 15.370 25.365 15.600 26.355 ;
        RECT 14.935 25.195 15.600 25.365 ;
        RECT 14.935 24.905 15.105 25.195 ;
        RECT 15.275 24.645 15.605 25.025 ;
        RECT 15.775 24.905 15.960 27.025 ;
        RECT 16.200 26.735 16.465 27.195 ;
        RECT 16.635 26.600 16.885 27.025 ;
        RECT 17.095 26.750 18.200 26.920 ;
        RECT 16.580 26.470 16.885 26.600 ;
        RECT 16.130 25.275 16.410 26.225 ;
        RECT 16.580 25.365 16.750 26.470 ;
        RECT 16.920 25.685 17.160 26.280 ;
        RECT 17.330 26.215 17.860 26.580 ;
        RECT 17.330 25.515 17.500 26.215 ;
        RECT 18.030 26.135 18.200 26.750 ;
        RECT 18.370 26.395 18.540 27.195 ;
        RECT 18.710 26.695 18.960 27.025 ;
        RECT 19.185 26.725 20.070 26.895 ;
        RECT 18.030 26.045 18.540 26.135 ;
        RECT 16.580 25.235 16.805 25.365 ;
        RECT 16.975 25.295 17.500 25.515 ;
        RECT 17.670 25.875 18.540 26.045 ;
        RECT 16.215 24.645 16.465 25.105 ;
        RECT 16.635 25.095 16.805 25.235 ;
        RECT 17.670 25.095 17.840 25.875 ;
        RECT 18.370 25.805 18.540 25.875 ;
        RECT 18.050 25.625 18.250 25.655 ;
        RECT 18.710 25.625 18.880 26.695 ;
        RECT 19.050 25.805 19.240 26.525 ;
        RECT 18.050 25.325 18.880 25.625 ;
        RECT 19.410 25.595 19.730 26.555 ;
        RECT 16.635 24.925 16.970 25.095 ;
        RECT 17.165 24.925 17.840 25.095 ;
        RECT 18.160 24.645 18.530 25.145 ;
        RECT 18.710 25.095 18.880 25.325 ;
        RECT 19.265 25.265 19.730 25.595 ;
        RECT 19.900 25.885 20.070 26.725 ;
        RECT 20.250 26.695 20.565 27.195 ;
        RECT 20.795 26.465 21.135 27.025 ;
        RECT 20.240 26.090 21.135 26.465 ;
        RECT 21.305 26.185 21.475 27.195 ;
        RECT 20.945 25.885 21.135 26.090 ;
        RECT 21.645 26.135 21.975 26.980 ;
        RECT 22.210 26.805 22.545 27.025 ;
        RECT 23.550 26.815 23.905 27.195 ;
        RECT 22.210 26.185 22.465 26.805 ;
        RECT 22.715 26.645 22.945 26.685 ;
        RECT 24.075 26.645 24.325 27.025 ;
        RECT 22.715 26.445 24.325 26.645 ;
        RECT 22.715 26.355 22.900 26.445 ;
        RECT 23.490 26.435 24.325 26.445 ;
        RECT 24.575 26.415 24.825 27.195 ;
        RECT 24.995 26.345 25.255 27.025 ;
        RECT 23.055 26.245 23.385 26.275 ;
        RECT 23.055 26.185 24.855 26.245 ;
        RECT 21.645 26.055 22.035 26.135 ;
        RECT 21.820 26.005 22.035 26.055 ;
        RECT 22.210 26.075 24.915 26.185 ;
        RECT 22.210 26.015 23.385 26.075 ;
        RECT 24.715 26.040 24.915 26.075 ;
        RECT 19.900 25.555 20.775 25.885 ;
        RECT 20.945 25.555 21.695 25.885 ;
        RECT 19.900 25.095 20.070 25.555 ;
        RECT 20.945 25.385 21.145 25.555 ;
        RECT 21.865 25.425 22.035 26.005 ;
        RECT 22.205 25.635 22.695 25.835 ;
        RECT 22.885 25.635 23.360 25.845 ;
        RECT 21.810 25.385 22.035 25.425 ;
        RECT 18.710 24.925 19.115 25.095 ;
        RECT 19.285 24.925 20.070 25.095 ;
        RECT 20.345 24.645 20.555 25.175 ;
        RECT 20.815 24.860 21.145 25.385 ;
        RECT 21.655 25.300 22.035 25.385 ;
        RECT 21.315 24.645 21.485 25.255 ;
        RECT 21.655 24.865 21.985 25.300 ;
        RECT 22.210 24.645 22.665 25.410 ;
        RECT 23.140 25.235 23.360 25.635 ;
        RECT 23.605 25.635 23.935 25.845 ;
        RECT 23.605 25.235 23.815 25.635 ;
        RECT 24.105 25.600 24.515 25.905 ;
        RECT 24.745 25.465 24.915 26.040 ;
        RECT 24.645 25.345 24.915 25.465 ;
        RECT 24.070 25.300 24.915 25.345 ;
        RECT 24.070 25.175 24.825 25.300 ;
        RECT 24.070 25.025 24.240 25.175 ;
        RECT 25.085 25.145 25.255 26.345 ;
        RECT 26.345 26.030 26.635 27.195 ;
        RECT 26.805 26.105 28.015 27.195 ;
        RECT 28.275 26.525 28.445 27.025 ;
        RECT 28.615 26.695 28.945 27.195 ;
        RECT 28.275 26.355 28.940 26.525 ;
        RECT 26.805 25.395 27.325 25.935 ;
        RECT 27.495 25.565 28.015 26.105 ;
        RECT 28.190 25.535 28.540 26.185 ;
        RECT 22.940 24.815 24.240 25.025 ;
        RECT 24.495 24.645 24.825 25.005 ;
        RECT 24.995 24.815 25.255 25.145 ;
        RECT 26.345 24.645 26.635 25.370 ;
        RECT 26.805 24.645 28.015 25.395 ;
        RECT 28.710 25.365 28.940 26.355 ;
        RECT 28.275 25.195 28.940 25.365 ;
        RECT 28.275 24.905 28.445 25.195 ;
        RECT 28.615 24.645 28.945 25.025 ;
        RECT 29.115 24.905 29.300 27.025 ;
        RECT 29.540 26.735 29.805 27.195 ;
        RECT 29.975 26.600 30.225 27.025 ;
        RECT 30.435 26.750 31.540 26.920 ;
        RECT 29.920 26.470 30.225 26.600 ;
        RECT 29.470 25.275 29.750 26.225 ;
        RECT 29.920 25.365 30.090 26.470 ;
        RECT 30.260 25.685 30.500 26.280 ;
        RECT 30.670 26.215 31.200 26.580 ;
        RECT 30.670 25.515 30.840 26.215 ;
        RECT 31.370 26.135 31.540 26.750 ;
        RECT 31.710 26.395 31.880 27.195 ;
        RECT 32.050 26.695 32.300 27.025 ;
        RECT 32.525 26.725 33.410 26.895 ;
        RECT 31.370 26.045 31.880 26.135 ;
        RECT 29.920 25.235 30.145 25.365 ;
        RECT 30.315 25.295 30.840 25.515 ;
        RECT 31.010 25.875 31.880 26.045 ;
        RECT 29.555 24.645 29.805 25.105 ;
        RECT 29.975 25.095 30.145 25.235 ;
        RECT 31.010 25.095 31.180 25.875 ;
        RECT 31.710 25.805 31.880 25.875 ;
        RECT 31.390 25.625 31.590 25.655 ;
        RECT 32.050 25.625 32.220 26.695 ;
        RECT 32.390 25.805 32.580 26.525 ;
        RECT 31.390 25.325 32.220 25.625 ;
        RECT 32.750 25.595 33.070 26.555 ;
        RECT 29.975 24.925 30.310 25.095 ;
        RECT 30.505 24.925 31.180 25.095 ;
        RECT 31.500 24.645 31.870 25.145 ;
        RECT 32.050 25.095 32.220 25.325 ;
        RECT 32.605 25.265 33.070 25.595 ;
        RECT 33.240 25.885 33.410 26.725 ;
        RECT 33.590 26.695 33.905 27.195 ;
        RECT 34.135 26.465 34.475 27.025 ;
        RECT 33.580 26.090 34.475 26.465 ;
        RECT 34.645 26.185 34.815 27.195 ;
        RECT 34.285 25.885 34.475 26.090 ;
        RECT 34.985 26.135 35.315 26.980 ;
        RECT 35.635 26.525 35.805 27.025 ;
        RECT 35.975 26.695 36.305 27.195 ;
        RECT 35.635 26.355 36.300 26.525 ;
        RECT 34.985 26.055 35.375 26.135 ;
        RECT 35.160 26.005 35.375 26.055 ;
        RECT 33.240 25.555 34.115 25.885 ;
        RECT 34.285 25.555 35.035 25.885 ;
        RECT 33.240 25.095 33.410 25.555 ;
        RECT 34.285 25.385 34.485 25.555 ;
        RECT 35.205 25.425 35.375 26.005 ;
        RECT 35.550 25.535 35.900 26.185 ;
        RECT 35.150 25.385 35.375 25.425 ;
        RECT 32.050 24.925 32.455 25.095 ;
        RECT 32.625 24.925 33.410 25.095 ;
        RECT 33.685 24.645 33.895 25.175 ;
        RECT 34.155 24.860 34.485 25.385 ;
        RECT 34.995 25.300 35.375 25.385 ;
        RECT 36.070 25.365 36.300 26.355 ;
        RECT 34.655 24.645 34.825 25.255 ;
        RECT 34.995 24.865 35.325 25.300 ;
        RECT 35.635 25.195 36.300 25.365 ;
        RECT 35.635 24.905 35.805 25.195 ;
        RECT 35.975 24.645 36.305 25.025 ;
        RECT 36.475 24.905 36.660 27.025 ;
        RECT 36.900 26.735 37.165 27.195 ;
        RECT 37.335 26.600 37.585 27.025 ;
        RECT 37.795 26.750 38.900 26.920 ;
        RECT 37.280 26.470 37.585 26.600 ;
        RECT 36.830 25.275 37.110 26.225 ;
        RECT 37.280 25.365 37.450 26.470 ;
        RECT 37.620 25.685 37.860 26.280 ;
        RECT 38.030 26.215 38.560 26.580 ;
        RECT 38.030 25.515 38.200 26.215 ;
        RECT 38.730 26.135 38.900 26.750 ;
        RECT 39.070 26.395 39.240 27.195 ;
        RECT 39.410 26.695 39.660 27.025 ;
        RECT 39.885 26.725 40.770 26.895 ;
        RECT 38.730 26.045 39.240 26.135 ;
        RECT 37.280 25.235 37.505 25.365 ;
        RECT 37.675 25.295 38.200 25.515 ;
        RECT 38.370 25.875 39.240 26.045 ;
        RECT 36.915 24.645 37.165 25.105 ;
        RECT 37.335 25.095 37.505 25.235 ;
        RECT 38.370 25.095 38.540 25.875 ;
        RECT 39.070 25.805 39.240 25.875 ;
        RECT 38.750 25.625 38.950 25.655 ;
        RECT 39.410 25.625 39.580 26.695 ;
        RECT 39.750 25.805 39.940 26.525 ;
        RECT 38.750 25.325 39.580 25.625 ;
        RECT 40.110 25.595 40.430 26.555 ;
        RECT 37.335 24.925 37.670 25.095 ;
        RECT 37.865 24.925 38.540 25.095 ;
        RECT 38.860 24.645 39.230 25.145 ;
        RECT 39.410 25.095 39.580 25.325 ;
        RECT 39.965 25.265 40.430 25.595 ;
        RECT 40.600 25.885 40.770 26.725 ;
        RECT 40.950 26.695 41.265 27.195 ;
        RECT 41.495 26.465 41.835 27.025 ;
        RECT 40.940 26.090 41.835 26.465 ;
        RECT 42.005 26.185 42.175 27.195 ;
        RECT 41.645 25.885 41.835 26.090 ;
        RECT 42.345 26.135 42.675 26.980 ;
        RECT 42.345 26.055 42.735 26.135 ;
        RECT 42.520 26.005 42.735 26.055 ;
        RECT 40.600 25.555 41.475 25.885 ;
        RECT 41.645 25.555 42.395 25.885 ;
        RECT 40.600 25.095 40.770 25.555 ;
        RECT 41.645 25.385 41.845 25.555 ;
        RECT 42.565 25.425 42.735 26.005 ;
        RECT 42.510 25.385 42.735 25.425 ;
        RECT 39.410 24.925 39.815 25.095 ;
        RECT 39.985 24.925 40.770 25.095 ;
        RECT 41.045 24.645 41.255 25.175 ;
        RECT 41.515 24.860 41.845 25.385 ;
        RECT 42.355 25.300 42.735 25.385 ;
        RECT 43.825 26.055 44.165 27.025 ;
        RECT 44.335 26.055 44.505 27.195 ;
        RECT 44.775 26.395 45.025 27.195 ;
        RECT 45.670 26.225 46.000 27.025 ;
        RECT 46.300 26.395 46.630 27.195 ;
        RECT 46.800 26.225 47.130 27.025 ;
        RECT 44.695 26.055 47.130 26.225 ;
        RECT 47.505 26.105 49.175 27.195 ;
        RECT 43.825 25.445 44.000 26.055 ;
        RECT 44.695 25.805 44.865 26.055 ;
        RECT 44.170 25.635 44.865 25.805 ;
        RECT 45.040 25.635 45.460 25.835 ;
        RECT 45.630 25.635 45.960 25.835 ;
        RECT 46.130 25.635 46.460 25.835 ;
        RECT 42.015 24.645 42.185 25.255 ;
        RECT 42.355 24.865 42.685 25.300 ;
        RECT 43.825 24.815 44.165 25.445 ;
        RECT 44.335 24.645 44.585 25.445 ;
        RECT 44.775 25.295 46.000 25.465 ;
        RECT 44.775 24.815 45.105 25.295 ;
        RECT 45.275 24.645 45.500 25.105 ;
        RECT 45.670 24.815 46.000 25.295 ;
        RECT 46.630 25.425 46.800 26.055 ;
        RECT 46.985 25.635 47.335 25.885 ;
        RECT 46.630 24.815 47.130 25.425 ;
        RECT 47.505 25.415 48.255 25.935 ;
        RECT 48.425 25.585 49.175 26.105 ;
        RECT 49.990 26.225 50.380 26.400 ;
        RECT 50.865 26.395 51.195 27.195 ;
        RECT 51.365 26.405 51.900 27.025 ;
        RECT 49.990 26.055 51.415 26.225 ;
        RECT 47.505 24.645 49.175 25.415 ;
        RECT 49.865 25.325 50.220 25.885 ;
        RECT 50.390 25.155 50.560 26.055 ;
        RECT 50.730 25.325 50.995 25.885 ;
        RECT 51.245 25.555 51.415 26.055 ;
        RECT 51.585 25.385 51.900 26.405 ;
        RECT 52.105 26.030 52.395 27.195 ;
        RECT 52.565 26.055 52.905 27.025 ;
        RECT 53.075 26.055 53.245 27.195 ;
        RECT 53.515 26.395 53.765 27.195 ;
        RECT 54.410 26.225 54.740 27.025 ;
        RECT 55.040 26.395 55.370 27.195 ;
        RECT 55.540 26.225 55.870 27.025 ;
        RECT 53.435 26.055 55.870 26.225 ;
        RECT 56.245 26.105 57.915 27.195 ;
        RECT 49.970 24.645 50.210 25.155 ;
        RECT 50.390 24.825 50.670 25.155 ;
        RECT 50.900 24.645 51.115 25.155 ;
        RECT 51.285 24.815 51.900 25.385 ;
        RECT 52.565 25.445 52.740 26.055 ;
        RECT 53.435 25.805 53.605 26.055 ;
        RECT 52.910 25.635 53.605 25.805 ;
        RECT 53.780 25.635 54.200 25.835 ;
        RECT 54.370 25.635 54.700 25.835 ;
        RECT 54.870 25.635 55.200 25.835 ;
        RECT 52.105 24.645 52.395 25.370 ;
        RECT 52.565 24.815 52.905 25.445 ;
        RECT 53.075 24.645 53.325 25.445 ;
        RECT 53.515 25.295 54.740 25.465 ;
        RECT 53.515 24.815 53.845 25.295 ;
        RECT 54.015 24.645 54.240 25.105 ;
        RECT 54.410 24.815 54.740 25.295 ;
        RECT 55.370 25.425 55.540 26.055 ;
        RECT 55.725 25.635 56.075 25.885 ;
        RECT 55.370 24.815 55.870 25.425 ;
        RECT 56.245 25.415 56.995 25.935 ;
        RECT 57.165 25.585 57.915 26.105 ;
        RECT 58.090 26.045 58.350 27.195 ;
        RECT 58.525 26.120 58.780 27.025 ;
        RECT 58.950 26.435 59.280 27.195 ;
        RECT 59.495 26.265 59.665 27.025 ;
        RECT 59.925 26.760 65.270 27.195 ;
        RECT 65.445 26.760 70.790 27.195 ;
        RECT 56.245 24.645 57.915 25.415 ;
        RECT 58.090 24.645 58.350 25.485 ;
        RECT 58.525 25.390 58.695 26.120 ;
        RECT 58.950 26.095 59.665 26.265 ;
        RECT 58.950 25.885 59.120 26.095 ;
        RECT 58.865 25.555 59.120 25.885 ;
        RECT 58.525 24.815 58.780 25.390 ;
        RECT 58.950 25.365 59.120 25.555 ;
        RECT 59.400 25.545 59.755 25.915 ;
        RECT 58.950 25.195 59.665 25.365 ;
        RECT 58.950 24.645 59.280 25.025 ;
        RECT 59.495 24.815 59.665 25.195 ;
        RECT 61.510 25.190 61.850 26.020 ;
        RECT 63.330 25.510 63.680 26.760 ;
        RECT 67.030 25.190 67.370 26.020 ;
        RECT 68.850 25.510 69.200 26.760 ;
        RECT 70.965 26.105 74.475 27.195 ;
        RECT 70.965 25.415 72.615 25.935 ;
        RECT 72.785 25.585 74.475 26.105 ;
        RECT 75.750 26.225 76.140 26.400 ;
        RECT 76.625 26.395 76.955 27.195 ;
        RECT 77.125 26.405 77.660 27.025 ;
        RECT 75.750 26.055 77.175 26.225 ;
        RECT 59.925 24.645 65.270 25.190 ;
        RECT 65.445 24.645 70.790 25.190 ;
        RECT 70.965 24.645 74.475 25.415 ;
        RECT 75.625 25.325 75.980 25.885 ;
        RECT 76.150 25.155 76.320 26.055 ;
        RECT 76.490 25.325 76.755 25.885 ;
        RECT 77.005 25.555 77.175 26.055 ;
        RECT 77.345 25.385 77.660 26.405 ;
        RECT 77.865 26.030 78.155 27.195 ;
        RECT 78.325 26.055 78.665 27.025 ;
        RECT 78.835 26.055 79.005 27.195 ;
        RECT 79.275 26.395 79.525 27.195 ;
        RECT 80.170 26.225 80.500 27.025 ;
        RECT 80.800 26.395 81.130 27.195 ;
        RECT 81.300 26.225 81.630 27.025 ;
        RECT 79.195 26.055 81.630 26.225 ;
        RECT 82.005 26.105 83.215 27.195 ;
        RECT 83.475 26.525 83.645 27.025 ;
        RECT 83.815 26.695 84.145 27.195 ;
        RECT 83.475 26.355 84.140 26.525 ;
        RECT 75.730 24.645 75.970 25.155 ;
        RECT 76.150 24.825 76.430 25.155 ;
        RECT 76.660 24.645 76.875 25.155 ;
        RECT 77.045 24.815 77.660 25.385 ;
        RECT 78.325 25.445 78.500 26.055 ;
        RECT 79.195 25.805 79.365 26.055 ;
        RECT 78.670 25.635 79.365 25.805 ;
        RECT 79.540 25.635 79.960 25.835 ;
        RECT 80.130 25.635 80.460 25.835 ;
        RECT 80.630 25.635 80.960 25.835 ;
        RECT 77.865 24.645 78.155 25.370 ;
        RECT 78.325 24.815 78.665 25.445 ;
        RECT 78.835 24.645 79.085 25.445 ;
        RECT 79.275 25.295 80.500 25.465 ;
        RECT 79.275 24.815 79.605 25.295 ;
        RECT 79.775 24.645 80.000 25.105 ;
        RECT 80.170 24.815 80.500 25.295 ;
        RECT 81.130 25.425 81.300 26.055 ;
        RECT 81.485 25.635 81.835 25.885 ;
        RECT 81.130 24.815 81.630 25.425 ;
        RECT 82.005 25.395 82.525 25.935 ;
        RECT 82.695 25.565 83.215 26.105 ;
        RECT 83.390 25.535 83.740 26.185 ;
        RECT 82.005 24.645 83.215 25.395 ;
        RECT 83.910 25.365 84.140 26.355 ;
        RECT 83.475 25.195 84.140 25.365 ;
        RECT 83.475 24.905 83.645 25.195 ;
        RECT 83.815 24.645 84.145 25.025 ;
        RECT 84.315 24.905 84.500 27.025 ;
        RECT 84.740 26.735 85.005 27.195 ;
        RECT 85.175 26.600 85.425 27.025 ;
        RECT 85.635 26.750 86.740 26.920 ;
        RECT 85.120 26.470 85.425 26.600 ;
        RECT 84.670 25.275 84.950 26.225 ;
        RECT 85.120 25.365 85.290 26.470 ;
        RECT 85.460 25.685 85.700 26.280 ;
        RECT 85.870 26.215 86.400 26.580 ;
        RECT 85.870 25.515 86.040 26.215 ;
        RECT 86.570 26.135 86.740 26.750 ;
        RECT 86.910 26.395 87.080 27.195 ;
        RECT 87.250 26.695 87.500 27.025 ;
        RECT 87.725 26.725 88.610 26.895 ;
        RECT 86.570 26.045 87.080 26.135 ;
        RECT 85.120 25.235 85.345 25.365 ;
        RECT 85.515 25.295 86.040 25.515 ;
        RECT 86.210 25.875 87.080 26.045 ;
        RECT 84.755 24.645 85.005 25.105 ;
        RECT 85.175 25.095 85.345 25.235 ;
        RECT 86.210 25.095 86.380 25.875 ;
        RECT 86.910 25.805 87.080 25.875 ;
        RECT 86.590 25.625 86.790 25.655 ;
        RECT 87.250 25.625 87.420 26.695 ;
        RECT 87.590 25.805 87.780 26.525 ;
        RECT 86.590 25.325 87.420 25.625 ;
        RECT 87.950 25.595 88.270 26.555 ;
        RECT 85.175 24.925 85.510 25.095 ;
        RECT 85.705 24.925 86.380 25.095 ;
        RECT 86.700 24.645 87.070 25.145 ;
        RECT 87.250 25.095 87.420 25.325 ;
        RECT 87.805 25.265 88.270 25.595 ;
        RECT 88.440 25.885 88.610 26.725 ;
        RECT 88.790 26.695 89.105 27.195 ;
        RECT 89.335 26.465 89.675 27.025 ;
        RECT 88.780 26.090 89.675 26.465 ;
        RECT 89.845 26.185 90.015 27.195 ;
        RECT 89.485 25.885 89.675 26.090 ;
        RECT 90.185 26.135 90.515 26.980 ;
        RECT 90.185 26.055 90.575 26.135 ;
        RECT 90.360 26.005 90.575 26.055 ;
        RECT 88.440 25.555 89.315 25.885 ;
        RECT 89.485 25.555 90.235 25.885 ;
        RECT 88.440 25.095 88.610 25.555 ;
        RECT 89.485 25.385 89.685 25.555 ;
        RECT 90.405 25.425 90.575 26.005 ;
        RECT 90.745 26.105 91.955 27.195 ;
        RECT 90.745 25.565 91.265 26.105 ;
        RECT 90.350 25.385 90.575 25.425 ;
        RECT 91.435 25.395 91.955 25.935 ;
        RECT 87.250 24.925 87.655 25.095 ;
        RECT 87.825 24.925 88.610 25.095 ;
        RECT 88.885 24.645 89.095 25.175 ;
        RECT 89.355 24.860 89.685 25.385 ;
        RECT 90.195 25.300 90.575 25.385 ;
        RECT 89.855 24.645 90.025 25.255 ;
        RECT 90.195 24.865 90.525 25.300 ;
        RECT 90.745 24.645 91.955 25.395 ;
        RECT 13.380 24.475 92.040 24.645 ;
        RECT 13.465 23.725 14.675 24.475 ;
        RECT 13.465 23.185 13.985 23.725 ;
        RECT 14.850 23.635 15.110 24.475 ;
        RECT 15.285 23.730 15.540 24.305 ;
        RECT 15.710 24.095 16.040 24.475 ;
        RECT 16.255 23.925 16.425 24.305 ;
        RECT 15.710 23.755 16.425 23.925 ;
        RECT 14.155 23.015 14.675 23.555 ;
        RECT 13.465 21.925 14.675 23.015 ;
        RECT 14.850 21.925 15.110 23.075 ;
        RECT 15.285 23.000 15.455 23.730 ;
        RECT 15.710 23.565 15.880 23.755 ;
        RECT 16.685 23.725 17.895 24.475 ;
        RECT 15.625 23.235 15.880 23.565 ;
        RECT 15.710 23.025 15.880 23.235 ;
        RECT 16.160 23.205 16.515 23.575 ;
        RECT 16.685 23.185 17.205 23.725 ;
        RECT 18.070 23.635 18.330 24.475 ;
        RECT 18.505 23.730 18.760 24.305 ;
        RECT 18.930 24.095 19.260 24.475 ;
        RECT 19.475 23.925 19.645 24.305 ;
        RECT 18.930 23.755 19.645 23.925 ;
        RECT 15.285 22.095 15.540 23.000 ;
        RECT 15.710 22.855 16.425 23.025 ;
        RECT 17.375 23.015 17.895 23.555 ;
        RECT 15.710 21.925 16.040 22.685 ;
        RECT 16.255 22.095 16.425 22.855 ;
        RECT 16.685 21.925 17.895 23.015 ;
        RECT 18.070 21.925 18.330 23.075 ;
        RECT 18.505 23.000 18.675 23.730 ;
        RECT 18.930 23.565 19.100 23.755 ;
        RECT 19.910 23.635 20.170 24.475 ;
        RECT 20.345 23.730 20.600 24.305 ;
        RECT 20.770 24.095 21.100 24.475 ;
        RECT 21.315 23.925 21.485 24.305 ;
        RECT 20.770 23.755 21.485 23.925 ;
        RECT 18.845 23.235 19.100 23.565 ;
        RECT 18.930 23.025 19.100 23.235 ;
        RECT 19.380 23.205 19.735 23.575 ;
        RECT 18.505 22.095 18.760 23.000 ;
        RECT 18.930 22.855 19.645 23.025 ;
        RECT 18.930 21.925 19.260 22.685 ;
        RECT 19.475 22.095 19.645 22.855 ;
        RECT 19.910 21.925 20.170 23.075 ;
        RECT 20.345 23.000 20.515 23.730 ;
        RECT 20.770 23.565 20.940 23.755 ;
        RECT 22.670 23.710 23.125 24.475 ;
        RECT 23.400 24.095 24.700 24.305 ;
        RECT 24.955 24.115 25.285 24.475 ;
        RECT 24.530 23.945 24.700 24.095 ;
        RECT 25.455 23.975 25.715 24.305 ;
        RECT 20.685 23.235 20.940 23.565 ;
        RECT 20.770 23.025 20.940 23.235 ;
        RECT 21.220 23.205 21.575 23.575 ;
        RECT 23.600 23.485 23.820 23.885 ;
        RECT 22.665 23.285 23.155 23.485 ;
        RECT 23.345 23.275 23.820 23.485 ;
        RECT 24.065 23.485 24.275 23.885 ;
        RECT 24.530 23.820 25.285 23.945 ;
        RECT 24.530 23.775 25.375 23.820 ;
        RECT 25.105 23.655 25.375 23.775 ;
        RECT 24.065 23.275 24.395 23.485 ;
        RECT 24.565 23.215 24.975 23.520 ;
        RECT 22.670 23.045 23.845 23.105 ;
        RECT 25.205 23.080 25.375 23.655 ;
        RECT 25.175 23.045 25.375 23.080 ;
        RECT 20.345 22.095 20.600 23.000 ;
        RECT 20.770 22.855 21.485 23.025 ;
        RECT 20.770 21.925 21.100 22.685 ;
        RECT 21.315 22.095 21.485 22.855 ;
        RECT 22.670 22.935 25.375 23.045 ;
        RECT 22.670 22.315 22.925 22.935 ;
        RECT 23.515 22.875 25.315 22.935 ;
        RECT 23.515 22.845 23.845 22.875 ;
        RECT 25.545 22.775 25.715 23.975 ;
        RECT 25.975 23.925 26.145 24.305 ;
        RECT 26.360 24.095 26.690 24.475 ;
        RECT 25.975 23.755 26.690 23.925 ;
        RECT 25.885 23.205 26.240 23.575 ;
        RECT 26.520 23.565 26.690 23.755 ;
        RECT 26.860 23.730 27.115 24.305 ;
        RECT 26.520 23.235 26.775 23.565 ;
        RECT 26.520 23.025 26.690 23.235 ;
        RECT 23.175 22.675 23.360 22.765 ;
        RECT 23.950 22.675 24.785 22.685 ;
        RECT 23.175 22.475 24.785 22.675 ;
        RECT 23.175 22.435 23.405 22.475 ;
        RECT 22.670 22.095 23.005 22.315 ;
        RECT 24.010 21.925 24.365 22.305 ;
        RECT 24.535 22.095 24.785 22.475 ;
        RECT 25.035 21.925 25.285 22.705 ;
        RECT 25.455 22.095 25.715 22.775 ;
        RECT 25.975 22.855 26.690 23.025 ;
        RECT 26.945 23.000 27.115 23.730 ;
        RECT 27.290 23.635 27.550 24.475 ;
        RECT 28.810 23.965 29.050 24.475 ;
        RECT 29.230 23.965 29.510 24.295 ;
        RECT 29.740 23.965 29.955 24.475 ;
        RECT 28.705 23.235 29.060 23.795 ;
        RECT 25.975 22.095 26.145 22.855 ;
        RECT 26.360 21.925 26.690 22.685 ;
        RECT 26.860 22.095 27.115 23.000 ;
        RECT 27.290 21.925 27.550 23.075 ;
        RECT 29.230 23.065 29.400 23.965 ;
        RECT 29.570 23.235 29.835 23.795 ;
        RECT 30.125 23.735 30.740 24.305 ;
        RECT 30.945 23.930 36.290 24.475 ;
        RECT 30.085 23.065 30.255 23.565 ;
        RECT 28.830 22.895 30.255 23.065 ;
        RECT 28.830 22.720 29.220 22.895 ;
        RECT 29.705 21.925 30.035 22.725 ;
        RECT 30.425 22.715 30.740 23.735 ;
        RECT 32.530 23.100 32.870 23.930 ;
        RECT 36.465 23.705 39.055 24.475 ;
        RECT 39.225 23.750 39.515 24.475 ;
        RECT 39.685 23.705 41.355 24.475 ;
        RECT 41.530 23.710 41.985 24.475 ;
        RECT 42.260 24.095 43.560 24.305 ;
        RECT 43.815 24.115 44.145 24.475 ;
        RECT 43.390 23.945 43.560 24.095 ;
        RECT 44.315 23.975 44.575 24.305 ;
        RECT 30.205 22.095 30.740 22.715 ;
        RECT 34.350 22.360 34.700 23.610 ;
        RECT 36.465 23.185 37.675 23.705 ;
        RECT 37.845 23.015 39.055 23.535 ;
        RECT 39.685 23.185 40.435 23.705 ;
        RECT 30.945 21.925 36.290 22.360 ;
        RECT 36.465 21.925 39.055 23.015 ;
        RECT 39.225 21.925 39.515 23.090 ;
        RECT 40.605 23.015 41.355 23.535 ;
        RECT 42.460 23.485 42.680 23.885 ;
        RECT 41.525 23.285 42.015 23.485 ;
        RECT 42.205 23.275 42.680 23.485 ;
        RECT 42.925 23.485 43.135 23.885 ;
        RECT 43.390 23.820 44.145 23.945 ;
        RECT 43.390 23.775 44.235 23.820 ;
        RECT 43.965 23.655 44.235 23.775 ;
        RECT 42.925 23.275 43.255 23.485 ;
        RECT 43.425 23.215 43.835 23.520 ;
        RECT 39.685 21.925 41.355 23.015 ;
        RECT 41.530 23.045 42.705 23.105 ;
        RECT 44.065 23.080 44.235 23.655 ;
        RECT 44.035 23.045 44.235 23.080 ;
        RECT 41.530 22.935 44.235 23.045 ;
        RECT 41.530 22.315 41.785 22.935 ;
        RECT 42.375 22.875 44.175 22.935 ;
        RECT 42.375 22.845 42.705 22.875 ;
        RECT 44.405 22.775 44.575 23.975 ;
        RECT 44.745 23.725 45.955 24.475 ;
        RECT 44.745 23.185 45.265 23.725 ;
        RECT 46.130 23.710 46.585 24.475 ;
        RECT 46.860 24.095 48.160 24.305 ;
        RECT 48.415 24.115 48.745 24.475 ;
        RECT 47.990 23.945 48.160 24.095 ;
        RECT 48.915 23.975 49.175 24.305 ;
        RECT 45.435 23.015 45.955 23.555 ;
        RECT 47.060 23.485 47.280 23.885 ;
        RECT 46.125 23.285 46.615 23.485 ;
        RECT 46.805 23.275 47.280 23.485 ;
        RECT 47.525 23.485 47.735 23.885 ;
        RECT 47.990 23.820 48.745 23.945 ;
        RECT 47.990 23.775 48.835 23.820 ;
        RECT 48.565 23.655 48.835 23.775 ;
        RECT 47.525 23.275 47.855 23.485 ;
        RECT 48.025 23.215 48.435 23.520 ;
        RECT 42.035 22.675 42.220 22.765 ;
        RECT 42.810 22.675 43.645 22.685 ;
        RECT 42.035 22.475 43.645 22.675 ;
        RECT 42.035 22.435 42.265 22.475 ;
        RECT 41.530 22.095 41.865 22.315 ;
        RECT 42.870 21.925 43.225 22.305 ;
        RECT 43.395 22.095 43.645 22.475 ;
        RECT 43.895 21.925 44.145 22.705 ;
        RECT 44.315 22.095 44.575 22.775 ;
        RECT 44.745 21.925 45.955 23.015 ;
        RECT 46.130 23.045 47.305 23.105 ;
        RECT 48.665 23.080 48.835 23.655 ;
        RECT 48.635 23.045 48.835 23.080 ;
        RECT 46.130 22.935 48.835 23.045 ;
        RECT 46.130 22.315 46.385 22.935 ;
        RECT 46.975 22.875 48.775 22.935 ;
        RECT 46.975 22.845 47.305 22.875 ;
        RECT 49.005 22.775 49.175 23.975 ;
        RECT 49.345 23.930 54.690 24.475 ;
        RECT 50.930 23.100 51.270 23.930 ;
        RECT 54.865 23.705 58.375 24.475 ;
        RECT 46.635 22.675 46.820 22.765 ;
        RECT 47.410 22.675 48.245 22.685 ;
        RECT 46.635 22.475 48.245 22.675 ;
        RECT 46.635 22.435 46.865 22.475 ;
        RECT 46.130 22.095 46.465 22.315 ;
        RECT 47.470 21.925 47.825 22.305 ;
        RECT 47.995 22.095 48.245 22.475 ;
        RECT 48.495 21.925 48.745 22.705 ;
        RECT 48.915 22.095 49.175 22.775 ;
        RECT 52.750 22.360 53.100 23.610 ;
        RECT 54.865 23.185 56.515 23.705 ;
        RECT 59.005 23.675 59.345 24.305 ;
        RECT 59.515 23.675 59.765 24.475 ;
        RECT 59.955 23.825 60.285 24.305 ;
        RECT 60.455 24.015 60.680 24.475 ;
        RECT 60.850 23.825 61.180 24.305 ;
        RECT 56.685 23.015 58.375 23.535 ;
        RECT 49.345 21.925 54.690 22.360 ;
        RECT 54.865 21.925 58.375 23.015 ;
        RECT 59.005 23.065 59.180 23.675 ;
        RECT 59.955 23.655 61.180 23.825 ;
        RECT 61.810 23.695 62.310 24.305 ;
        RECT 62.720 23.735 63.335 24.305 ;
        RECT 63.505 23.965 63.720 24.475 ;
        RECT 63.950 23.965 64.230 24.295 ;
        RECT 64.410 23.965 64.650 24.475 ;
        RECT 59.350 23.315 60.045 23.485 ;
        RECT 59.875 23.065 60.045 23.315 ;
        RECT 60.220 23.285 60.640 23.485 ;
        RECT 60.810 23.285 61.140 23.485 ;
        RECT 61.310 23.285 61.640 23.485 ;
        RECT 61.810 23.065 61.980 23.695 ;
        RECT 62.165 23.235 62.515 23.485 ;
        RECT 59.005 22.095 59.345 23.065 ;
        RECT 59.515 21.925 59.685 23.065 ;
        RECT 59.875 22.895 62.310 23.065 ;
        RECT 59.955 21.925 60.205 22.725 ;
        RECT 60.850 22.095 61.180 22.895 ;
        RECT 61.480 21.925 61.810 22.725 ;
        RECT 61.980 22.095 62.310 22.895 ;
        RECT 62.720 22.715 63.035 23.735 ;
        RECT 63.205 23.065 63.375 23.565 ;
        RECT 63.625 23.235 63.890 23.795 ;
        RECT 64.060 23.065 64.230 23.965 ;
        RECT 64.400 23.235 64.755 23.795 ;
        RECT 64.985 23.750 65.275 24.475 ;
        RECT 65.445 23.975 65.705 24.305 ;
        RECT 65.875 24.115 66.205 24.475 ;
        RECT 66.460 24.095 67.760 24.305 ;
        RECT 63.205 22.895 64.630 23.065 ;
        RECT 62.720 22.095 63.255 22.715 ;
        RECT 63.425 21.925 63.755 22.725 ;
        RECT 64.240 22.720 64.630 22.895 ;
        RECT 64.985 21.925 65.275 23.090 ;
        RECT 65.445 22.775 65.615 23.975 ;
        RECT 66.460 23.945 66.630 24.095 ;
        RECT 65.875 23.820 66.630 23.945 ;
        RECT 65.785 23.775 66.630 23.820 ;
        RECT 65.785 23.655 66.055 23.775 ;
        RECT 65.785 23.080 65.955 23.655 ;
        RECT 66.185 23.215 66.595 23.520 ;
        RECT 66.885 23.485 67.095 23.885 ;
        RECT 66.765 23.275 67.095 23.485 ;
        RECT 67.340 23.485 67.560 23.885 ;
        RECT 68.035 23.710 68.490 24.475 ;
        RECT 68.665 23.675 69.005 24.305 ;
        RECT 69.175 23.675 69.425 24.475 ;
        RECT 69.615 23.825 69.945 24.305 ;
        RECT 70.115 24.015 70.340 24.475 ;
        RECT 70.510 23.825 70.840 24.305 ;
        RECT 67.340 23.275 67.815 23.485 ;
        RECT 68.005 23.285 68.495 23.485 ;
        RECT 65.785 23.045 65.985 23.080 ;
        RECT 67.315 23.045 68.490 23.105 ;
        RECT 65.785 22.935 68.490 23.045 ;
        RECT 65.845 22.875 67.645 22.935 ;
        RECT 67.315 22.845 67.645 22.875 ;
        RECT 65.445 22.095 65.705 22.775 ;
        RECT 65.875 21.925 66.125 22.705 ;
        RECT 66.375 22.675 67.210 22.685 ;
        RECT 67.800 22.675 67.985 22.765 ;
        RECT 66.375 22.475 67.985 22.675 ;
        RECT 66.375 22.095 66.625 22.475 ;
        RECT 67.755 22.435 67.985 22.475 ;
        RECT 68.235 22.315 68.490 22.935 ;
        RECT 66.795 21.925 67.150 22.305 ;
        RECT 68.155 22.095 68.490 22.315 ;
        RECT 68.665 23.065 68.840 23.675 ;
        RECT 69.615 23.655 70.840 23.825 ;
        RECT 71.470 23.695 71.970 24.305 ;
        RECT 72.380 23.735 72.995 24.305 ;
        RECT 73.165 23.965 73.380 24.475 ;
        RECT 73.610 23.965 73.890 24.295 ;
        RECT 74.070 23.965 74.310 24.475 ;
        RECT 69.010 23.315 69.705 23.485 ;
        RECT 69.535 23.065 69.705 23.315 ;
        RECT 69.880 23.285 70.300 23.485 ;
        RECT 70.470 23.285 70.800 23.485 ;
        RECT 70.970 23.285 71.300 23.485 ;
        RECT 71.470 23.065 71.640 23.695 ;
        RECT 71.825 23.235 72.175 23.485 ;
        RECT 68.665 22.095 69.005 23.065 ;
        RECT 69.175 21.925 69.345 23.065 ;
        RECT 69.535 22.895 71.970 23.065 ;
        RECT 69.615 21.925 69.865 22.725 ;
        RECT 70.510 22.095 70.840 22.895 ;
        RECT 71.140 21.925 71.470 22.725 ;
        RECT 71.640 22.095 71.970 22.895 ;
        RECT 72.380 22.715 72.695 23.735 ;
        RECT 72.865 23.065 73.035 23.565 ;
        RECT 73.285 23.235 73.550 23.795 ;
        RECT 73.720 23.065 73.890 23.965 ;
        RECT 74.060 23.235 74.415 23.795 ;
        RECT 74.645 23.705 76.315 24.475 ;
        RECT 76.945 23.975 77.205 24.305 ;
        RECT 77.375 24.115 77.705 24.475 ;
        RECT 77.960 24.095 79.260 24.305 ;
        RECT 74.645 23.185 75.395 23.705 ;
        RECT 72.865 22.895 74.290 23.065 ;
        RECT 75.565 23.015 76.315 23.535 ;
        RECT 72.380 22.095 72.915 22.715 ;
        RECT 73.085 21.925 73.415 22.725 ;
        RECT 73.900 22.720 74.290 22.895 ;
        RECT 74.645 21.925 76.315 23.015 ;
        RECT 76.945 22.775 77.115 23.975 ;
        RECT 77.960 23.945 78.130 24.095 ;
        RECT 77.375 23.820 78.130 23.945 ;
        RECT 77.285 23.775 78.130 23.820 ;
        RECT 77.285 23.655 77.555 23.775 ;
        RECT 77.285 23.080 77.455 23.655 ;
        RECT 77.685 23.215 78.095 23.520 ;
        RECT 78.385 23.485 78.595 23.885 ;
        RECT 78.265 23.275 78.595 23.485 ;
        RECT 78.840 23.485 79.060 23.885 ;
        RECT 79.535 23.710 79.990 24.475 ;
        RECT 80.370 23.695 80.870 24.305 ;
        RECT 78.840 23.275 79.315 23.485 ;
        RECT 79.505 23.285 79.995 23.485 ;
        RECT 80.165 23.235 80.515 23.485 ;
        RECT 77.285 23.045 77.485 23.080 ;
        RECT 78.815 23.045 79.990 23.105 ;
        RECT 80.700 23.065 80.870 23.695 ;
        RECT 81.500 23.825 81.830 24.305 ;
        RECT 82.000 24.015 82.225 24.475 ;
        RECT 82.395 23.825 82.725 24.305 ;
        RECT 81.500 23.655 82.725 23.825 ;
        RECT 82.915 23.675 83.165 24.475 ;
        RECT 83.335 23.675 83.675 24.305 ;
        RECT 81.040 23.285 81.370 23.485 ;
        RECT 81.540 23.285 81.870 23.485 ;
        RECT 82.040 23.285 82.460 23.485 ;
        RECT 82.635 23.315 83.330 23.485 ;
        RECT 82.635 23.065 82.805 23.315 ;
        RECT 83.500 23.115 83.675 23.675 ;
        RECT 83.845 23.725 85.055 24.475 ;
        RECT 85.315 23.925 85.485 24.305 ;
        RECT 85.700 24.095 86.030 24.475 ;
        RECT 85.315 23.755 86.030 23.925 ;
        RECT 83.845 23.185 84.365 23.725 ;
        RECT 83.445 23.065 83.675 23.115 ;
        RECT 77.285 22.935 79.990 23.045 ;
        RECT 77.345 22.875 79.145 22.935 ;
        RECT 78.815 22.845 79.145 22.875 ;
        RECT 76.945 22.095 77.205 22.775 ;
        RECT 77.375 21.925 77.625 22.705 ;
        RECT 77.875 22.675 78.710 22.685 ;
        RECT 79.300 22.675 79.485 22.765 ;
        RECT 77.875 22.475 79.485 22.675 ;
        RECT 77.875 22.095 78.125 22.475 ;
        RECT 79.255 22.435 79.485 22.475 ;
        RECT 79.735 22.315 79.990 22.935 ;
        RECT 78.295 21.925 78.650 22.305 ;
        RECT 79.655 22.095 79.990 22.315 ;
        RECT 80.370 22.895 82.805 23.065 ;
        RECT 80.370 22.095 80.700 22.895 ;
        RECT 80.870 21.925 81.200 22.725 ;
        RECT 81.500 22.095 81.830 22.895 ;
        RECT 82.475 21.925 82.725 22.725 ;
        RECT 82.995 21.925 83.165 23.065 ;
        RECT 83.335 22.095 83.675 23.065 ;
        RECT 84.535 23.015 85.055 23.555 ;
        RECT 85.225 23.205 85.580 23.575 ;
        RECT 85.860 23.565 86.030 23.755 ;
        RECT 86.200 23.730 86.455 24.305 ;
        RECT 85.860 23.235 86.115 23.565 ;
        RECT 85.860 23.025 86.030 23.235 ;
        RECT 83.845 21.925 85.055 23.015 ;
        RECT 85.315 22.855 86.030 23.025 ;
        RECT 86.285 23.000 86.455 23.730 ;
        RECT 86.630 23.635 86.890 24.475 ;
        RECT 87.155 23.925 87.325 24.305 ;
        RECT 87.540 24.095 87.870 24.475 ;
        RECT 87.155 23.755 87.870 23.925 ;
        RECT 87.065 23.205 87.420 23.575 ;
        RECT 87.700 23.565 87.870 23.755 ;
        RECT 88.040 23.730 88.295 24.305 ;
        RECT 87.700 23.235 87.955 23.565 ;
        RECT 85.315 22.095 85.485 22.855 ;
        RECT 85.700 21.925 86.030 22.685 ;
        RECT 86.200 22.095 86.455 23.000 ;
        RECT 86.630 21.925 86.890 23.075 ;
        RECT 87.700 23.025 87.870 23.235 ;
        RECT 87.155 22.855 87.870 23.025 ;
        RECT 88.125 23.000 88.295 23.730 ;
        RECT 88.470 23.635 88.730 24.475 ;
        RECT 88.910 23.635 89.170 24.475 ;
        RECT 89.345 23.730 89.600 24.305 ;
        RECT 89.770 24.095 90.100 24.475 ;
        RECT 90.315 23.925 90.485 24.305 ;
        RECT 89.770 23.755 90.485 23.925 ;
        RECT 87.155 22.095 87.325 22.855 ;
        RECT 87.540 21.925 87.870 22.685 ;
        RECT 88.040 22.095 88.295 23.000 ;
        RECT 88.470 21.925 88.730 23.075 ;
        RECT 88.910 21.925 89.170 23.075 ;
        RECT 89.345 23.000 89.515 23.730 ;
        RECT 89.770 23.565 89.940 23.755 ;
        RECT 90.745 23.725 91.955 24.475 ;
        RECT 89.685 23.235 89.940 23.565 ;
        RECT 89.770 23.025 89.940 23.235 ;
        RECT 90.220 23.205 90.575 23.575 ;
        RECT 89.345 22.095 89.600 23.000 ;
        RECT 89.770 22.855 90.485 23.025 ;
        RECT 89.770 21.925 90.100 22.685 ;
        RECT 90.315 22.095 90.485 22.855 ;
        RECT 90.745 23.015 91.265 23.555 ;
        RECT 91.435 23.185 91.955 23.725 ;
        RECT 90.745 21.925 91.955 23.015 ;
        RECT 13.380 21.755 92.040 21.925 ;
        RECT 13.465 20.665 14.675 21.755 ;
        RECT 13.465 19.955 13.985 20.495 ;
        RECT 14.155 20.125 14.675 20.665 ;
        RECT 15.305 20.615 15.645 21.585 ;
        RECT 15.815 20.615 15.985 21.755 ;
        RECT 16.255 20.955 16.505 21.755 ;
        RECT 17.150 20.785 17.480 21.585 ;
        RECT 17.780 20.955 18.110 21.755 ;
        RECT 18.280 20.785 18.610 21.585 ;
        RECT 16.175 20.615 18.610 20.785 ;
        RECT 15.305 20.005 15.480 20.615 ;
        RECT 16.175 20.365 16.345 20.615 ;
        RECT 15.650 20.195 16.345 20.365 ;
        RECT 16.520 20.195 16.940 20.395 ;
        RECT 17.110 20.195 17.440 20.395 ;
        RECT 17.610 20.195 17.940 20.395 ;
        RECT 13.465 19.205 14.675 19.955 ;
        RECT 15.305 19.375 15.645 20.005 ;
        RECT 15.815 19.205 16.065 20.005 ;
        RECT 16.255 19.855 17.480 20.025 ;
        RECT 16.255 19.375 16.585 19.855 ;
        RECT 16.755 19.205 16.980 19.665 ;
        RECT 17.150 19.375 17.480 19.855 ;
        RECT 18.110 19.985 18.280 20.615 ;
        RECT 19.910 20.605 20.170 21.755 ;
        RECT 20.345 20.680 20.600 21.585 ;
        RECT 20.770 20.995 21.100 21.755 ;
        RECT 21.315 20.825 21.485 21.585 ;
        RECT 18.465 20.195 18.815 20.445 ;
        RECT 18.110 19.375 18.610 19.985 ;
        RECT 19.910 19.205 20.170 20.045 ;
        RECT 20.345 19.950 20.515 20.680 ;
        RECT 20.770 20.655 21.485 20.825 ;
        RECT 20.770 20.445 20.940 20.655 ;
        RECT 21.745 20.615 22.085 21.585 ;
        RECT 22.255 20.615 22.425 21.755 ;
        RECT 22.695 20.955 22.945 21.755 ;
        RECT 23.590 20.785 23.920 21.585 ;
        RECT 24.220 20.955 24.550 21.755 ;
        RECT 24.720 20.785 25.050 21.585 ;
        RECT 22.615 20.615 25.050 20.785 ;
        RECT 20.685 20.115 20.940 20.445 ;
        RECT 20.345 19.375 20.600 19.950 ;
        RECT 20.770 19.925 20.940 20.115 ;
        RECT 21.220 20.105 21.575 20.475 ;
        RECT 21.745 20.005 21.920 20.615 ;
        RECT 22.615 20.365 22.785 20.615 ;
        RECT 22.090 20.195 22.785 20.365 ;
        RECT 22.960 20.195 23.380 20.395 ;
        RECT 23.550 20.195 23.880 20.395 ;
        RECT 24.050 20.195 24.380 20.395 ;
        RECT 20.770 19.755 21.485 19.925 ;
        RECT 20.770 19.205 21.100 19.585 ;
        RECT 21.315 19.375 21.485 19.755 ;
        RECT 21.745 19.375 22.085 20.005 ;
        RECT 22.255 19.205 22.505 20.005 ;
        RECT 22.695 19.855 23.920 20.025 ;
        RECT 22.695 19.375 23.025 19.855 ;
        RECT 23.195 19.205 23.420 19.665 ;
        RECT 23.590 19.375 23.920 19.855 ;
        RECT 24.550 19.985 24.720 20.615 ;
        RECT 26.345 20.590 26.635 21.755 ;
        RECT 27.470 20.785 27.800 21.585 ;
        RECT 27.970 20.955 28.300 21.755 ;
        RECT 28.600 20.785 28.930 21.585 ;
        RECT 29.575 20.955 29.825 21.755 ;
        RECT 27.470 20.615 29.905 20.785 ;
        RECT 30.095 20.615 30.265 21.755 ;
        RECT 30.435 20.615 30.775 21.585 ;
        RECT 31.150 20.785 31.480 21.585 ;
        RECT 31.650 20.955 31.980 21.755 ;
        RECT 32.280 20.785 32.610 21.585 ;
        RECT 33.255 20.955 33.505 21.755 ;
        RECT 31.150 20.615 33.585 20.785 ;
        RECT 33.775 20.615 33.945 21.755 ;
        RECT 34.115 20.615 34.455 21.585 ;
        RECT 34.715 21.085 34.885 21.585 ;
        RECT 35.055 21.255 35.385 21.755 ;
        RECT 34.715 20.915 35.380 21.085 ;
        RECT 24.905 20.195 25.255 20.445 ;
        RECT 27.265 20.195 27.615 20.445 ;
        RECT 27.800 19.985 27.970 20.615 ;
        RECT 28.140 20.195 28.470 20.395 ;
        RECT 28.640 20.195 28.970 20.395 ;
        RECT 29.140 20.195 29.560 20.395 ;
        RECT 29.735 20.365 29.905 20.615 ;
        RECT 29.735 20.195 30.430 20.365 ;
        RECT 24.550 19.375 25.050 19.985 ;
        RECT 26.345 19.205 26.635 19.930 ;
        RECT 27.470 19.375 27.970 19.985 ;
        RECT 28.600 19.855 29.825 20.025 ;
        RECT 30.600 20.005 30.775 20.615 ;
        RECT 30.945 20.195 31.295 20.445 ;
        RECT 28.600 19.375 28.930 19.855 ;
        RECT 29.100 19.205 29.325 19.665 ;
        RECT 29.495 19.375 29.825 19.855 ;
        RECT 30.015 19.205 30.265 20.005 ;
        RECT 30.435 19.375 30.775 20.005 ;
        RECT 31.480 19.985 31.650 20.615 ;
        RECT 31.820 20.195 32.150 20.395 ;
        RECT 32.320 20.195 32.650 20.395 ;
        RECT 32.820 20.195 33.240 20.395 ;
        RECT 33.415 20.365 33.585 20.615 ;
        RECT 33.415 20.195 34.110 20.365 ;
        RECT 34.280 20.055 34.455 20.615 ;
        RECT 34.630 20.095 34.980 20.745 ;
        RECT 31.150 19.375 31.650 19.985 ;
        RECT 32.280 19.855 33.505 20.025 ;
        RECT 34.225 20.005 34.455 20.055 ;
        RECT 32.280 19.375 32.610 19.855 ;
        RECT 32.780 19.205 33.005 19.665 ;
        RECT 33.175 19.375 33.505 19.855 ;
        RECT 33.695 19.205 33.945 20.005 ;
        RECT 34.115 19.375 34.455 20.005 ;
        RECT 35.150 19.925 35.380 20.915 ;
        RECT 34.715 19.755 35.380 19.925 ;
        RECT 34.715 19.465 34.885 19.755 ;
        RECT 35.055 19.205 35.385 19.585 ;
        RECT 35.555 19.465 35.740 21.585 ;
        RECT 35.980 21.295 36.245 21.755 ;
        RECT 36.415 21.160 36.665 21.585 ;
        RECT 36.875 21.310 37.980 21.480 ;
        RECT 36.360 21.030 36.665 21.160 ;
        RECT 35.910 19.835 36.190 20.785 ;
        RECT 36.360 19.925 36.530 21.030 ;
        RECT 36.700 20.245 36.940 20.840 ;
        RECT 37.110 20.775 37.640 21.140 ;
        RECT 37.110 20.075 37.280 20.775 ;
        RECT 37.810 20.695 37.980 21.310 ;
        RECT 38.150 20.955 38.320 21.755 ;
        RECT 38.490 21.255 38.740 21.585 ;
        RECT 38.965 21.285 39.850 21.455 ;
        RECT 37.810 20.605 38.320 20.695 ;
        RECT 36.360 19.795 36.585 19.925 ;
        RECT 36.755 19.855 37.280 20.075 ;
        RECT 37.450 20.435 38.320 20.605 ;
        RECT 35.995 19.205 36.245 19.665 ;
        RECT 36.415 19.655 36.585 19.795 ;
        RECT 37.450 19.655 37.620 20.435 ;
        RECT 38.150 20.365 38.320 20.435 ;
        RECT 37.830 20.185 38.030 20.215 ;
        RECT 38.490 20.185 38.660 21.255 ;
        RECT 38.830 20.365 39.020 21.085 ;
        RECT 37.830 19.885 38.660 20.185 ;
        RECT 39.190 20.155 39.510 21.115 ;
        RECT 36.415 19.485 36.750 19.655 ;
        RECT 36.945 19.485 37.620 19.655 ;
        RECT 37.940 19.205 38.310 19.705 ;
        RECT 38.490 19.655 38.660 19.885 ;
        RECT 39.045 19.825 39.510 20.155 ;
        RECT 39.680 20.445 39.850 21.285 ;
        RECT 40.030 21.255 40.345 21.755 ;
        RECT 40.575 21.025 40.915 21.585 ;
        RECT 40.020 20.650 40.915 21.025 ;
        RECT 41.085 20.745 41.255 21.755 ;
        RECT 40.725 20.445 40.915 20.650 ;
        RECT 41.425 20.695 41.755 21.540 ;
        RECT 41.425 20.615 41.815 20.695 ;
        RECT 41.600 20.565 41.815 20.615 ;
        RECT 39.680 20.115 40.555 20.445 ;
        RECT 40.725 20.115 41.475 20.445 ;
        RECT 39.680 19.655 39.850 20.115 ;
        RECT 40.725 19.945 40.925 20.115 ;
        RECT 41.645 19.985 41.815 20.565 ;
        RECT 41.590 19.945 41.815 19.985 ;
        RECT 38.490 19.485 38.895 19.655 ;
        RECT 39.065 19.485 39.850 19.655 ;
        RECT 40.125 19.205 40.335 19.735 ;
        RECT 40.595 19.420 40.925 19.945 ;
        RECT 41.435 19.860 41.815 19.945 ;
        RECT 42.905 20.615 43.245 21.585 ;
        RECT 43.415 20.615 43.585 21.755 ;
        RECT 43.855 20.955 44.105 21.755 ;
        RECT 44.750 20.785 45.080 21.585 ;
        RECT 45.380 20.955 45.710 21.755 ;
        RECT 45.880 20.785 46.210 21.585 ;
        RECT 43.775 20.615 46.210 20.785 ;
        RECT 46.585 20.665 48.255 21.755 ;
        RECT 42.905 20.005 43.080 20.615 ;
        RECT 43.775 20.365 43.945 20.615 ;
        RECT 43.250 20.195 43.945 20.365 ;
        RECT 44.120 20.195 44.540 20.395 ;
        RECT 44.710 20.195 45.040 20.395 ;
        RECT 45.210 20.195 45.540 20.395 ;
        RECT 41.095 19.205 41.265 19.815 ;
        RECT 41.435 19.425 41.765 19.860 ;
        RECT 42.905 19.375 43.245 20.005 ;
        RECT 43.415 19.205 43.665 20.005 ;
        RECT 43.855 19.855 45.080 20.025 ;
        RECT 43.855 19.375 44.185 19.855 ;
        RECT 44.355 19.205 44.580 19.665 ;
        RECT 44.750 19.375 45.080 19.855 ;
        RECT 45.710 19.985 45.880 20.615 ;
        RECT 46.065 20.195 46.415 20.445 ;
        RECT 45.710 19.375 46.210 19.985 ;
        RECT 46.585 19.975 47.335 20.495 ;
        RECT 47.505 20.145 48.255 20.665 ;
        RECT 48.425 20.615 48.765 21.585 ;
        RECT 48.935 20.615 49.105 21.755 ;
        RECT 49.375 20.955 49.625 21.755 ;
        RECT 50.270 20.785 50.600 21.585 ;
        RECT 50.900 20.955 51.230 21.755 ;
        RECT 51.400 20.785 51.730 21.585 ;
        RECT 49.295 20.615 51.730 20.785 ;
        RECT 48.425 20.005 48.600 20.615 ;
        RECT 49.295 20.365 49.465 20.615 ;
        RECT 48.770 20.195 49.465 20.365 ;
        RECT 49.640 20.195 50.060 20.395 ;
        RECT 50.230 20.195 50.560 20.395 ;
        RECT 50.730 20.195 51.060 20.395 ;
        RECT 46.585 19.205 48.255 19.975 ;
        RECT 48.425 19.375 48.765 20.005 ;
        RECT 48.935 19.205 49.185 20.005 ;
        RECT 49.375 19.855 50.600 20.025 ;
        RECT 49.375 19.375 49.705 19.855 ;
        RECT 49.875 19.205 50.100 19.665 ;
        RECT 50.270 19.375 50.600 19.855 ;
        RECT 51.230 19.985 51.400 20.615 ;
        RECT 52.105 20.590 52.395 21.755 ;
        RECT 52.565 20.665 54.235 21.755 ;
        RECT 51.585 20.195 51.935 20.445 ;
        RECT 51.230 19.375 51.730 19.985 ;
        RECT 52.565 19.975 53.315 20.495 ;
        RECT 53.485 20.145 54.235 20.665 ;
        RECT 54.865 20.615 55.205 21.585 ;
        RECT 55.375 20.615 55.545 21.755 ;
        RECT 55.815 20.955 56.065 21.755 ;
        RECT 56.710 20.785 57.040 21.585 ;
        RECT 57.340 20.955 57.670 21.755 ;
        RECT 57.840 20.785 58.170 21.585 ;
        RECT 58.635 21.085 58.805 21.585 ;
        RECT 58.975 21.255 59.305 21.755 ;
        RECT 58.635 20.915 59.300 21.085 ;
        RECT 55.735 20.615 58.170 20.785 ;
        RECT 54.865 20.005 55.040 20.615 ;
        RECT 55.735 20.365 55.905 20.615 ;
        RECT 55.210 20.195 55.905 20.365 ;
        RECT 56.080 20.195 56.500 20.395 ;
        RECT 56.670 20.195 57.000 20.395 ;
        RECT 57.170 20.195 57.500 20.395 ;
        RECT 52.105 19.205 52.395 19.930 ;
        RECT 52.565 19.205 54.235 19.975 ;
        RECT 54.865 19.375 55.205 20.005 ;
        RECT 55.375 19.205 55.625 20.005 ;
        RECT 55.815 19.855 57.040 20.025 ;
        RECT 55.815 19.375 56.145 19.855 ;
        RECT 56.315 19.205 56.540 19.665 ;
        RECT 56.710 19.375 57.040 19.855 ;
        RECT 57.670 19.985 57.840 20.615 ;
        RECT 58.025 20.195 58.375 20.445 ;
        RECT 58.550 20.095 58.900 20.745 ;
        RECT 57.670 19.375 58.170 19.985 ;
        RECT 59.070 19.925 59.300 20.915 ;
        RECT 58.635 19.755 59.300 19.925 ;
        RECT 58.635 19.465 58.805 19.755 ;
        RECT 58.975 19.205 59.305 19.585 ;
        RECT 59.475 19.465 59.660 21.585 ;
        RECT 59.900 21.295 60.165 21.755 ;
        RECT 60.335 21.160 60.585 21.585 ;
        RECT 60.795 21.310 61.900 21.480 ;
        RECT 60.280 21.030 60.585 21.160 ;
        RECT 59.830 19.835 60.110 20.785 ;
        RECT 60.280 19.925 60.450 21.030 ;
        RECT 60.620 20.245 60.860 20.840 ;
        RECT 61.030 20.775 61.560 21.140 ;
        RECT 61.030 20.075 61.200 20.775 ;
        RECT 61.730 20.695 61.900 21.310 ;
        RECT 62.070 20.955 62.240 21.755 ;
        RECT 62.410 21.255 62.660 21.585 ;
        RECT 62.885 21.285 63.770 21.455 ;
        RECT 61.730 20.605 62.240 20.695 ;
        RECT 60.280 19.795 60.505 19.925 ;
        RECT 60.675 19.855 61.200 20.075 ;
        RECT 61.370 20.435 62.240 20.605 ;
        RECT 59.915 19.205 60.165 19.665 ;
        RECT 60.335 19.655 60.505 19.795 ;
        RECT 61.370 19.655 61.540 20.435 ;
        RECT 62.070 20.365 62.240 20.435 ;
        RECT 61.750 20.185 61.950 20.215 ;
        RECT 62.410 20.185 62.580 21.255 ;
        RECT 62.750 20.365 62.940 21.085 ;
        RECT 61.750 19.885 62.580 20.185 ;
        RECT 63.110 20.155 63.430 21.115 ;
        RECT 60.335 19.485 60.670 19.655 ;
        RECT 60.865 19.485 61.540 19.655 ;
        RECT 61.860 19.205 62.230 19.705 ;
        RECT 62.410 19.655 62.580 19.885 ;
        RECT 62.965 19.825 63.430 20.155 ;
        RECT 63.600 20.445 63.770 21.285 ;
        RECT 63.950 21.255 64.265 21.755 ;
        RECT 64.495 21.025 64.835 21.585 ;
        RECT 63.940 20.650 64.835 21.025 ;
        RECT 65.005 20.745 65.175 21.755 ;
        RECT 64.645 20.445 64.835 20.650 ;
        RECT 65.345 20.695 65.675 21.540 ;
        RECT 65.995 21.085 66.165 21.585 ;
        RECT 66.335 21.255 66.665 21.755 ;
        RECT 65.995 20.915 66.660 21.085 ;
        RECT 65.345 20.615 65.735 20.695 ;
        RECT 65.520 20.565 65.735 20.615 ;
        RECT 63.600 20.115 64.475 20.445 ;
        RECT 64.645 20.115 65.395 20.445 ;
        RECT 63.600 19.655 63.770 20.115 ;
        RECT 64.645 19.945 64.845 20.115 ;
        RECT 65.565 19.985 65.735 20.565 ;
        RECT 65.910 20.095 66.260 20.745 ;
        RECT 65.510 19.945 65.735 19.985 ;
        RECT 62.410 19.485 62.815 19.655 ;
        RECT 62.985 19.485 63.770 19.655 ;
        RECT 64.045 19.205 64.255 19.735 ;
        RECT 64.515 19.420 64.845 19.945 ;
        RECT 65.355 19.860 65.735 19.945 ;
        RECT 66.430 19.925 66.660 20.915 ;
        RECT 65.015 19.205 65.185 19.815 ;
        RECT 65.355 19.425 65.685 19.860 ;
        RECT 65.995 19.755 66.660 19.925 ;
        RECT 65.995 19.465 66.165 19.755 ;
        RECT 66.335 19.205 66.665 19.585 ;
        RECT 66.835 19.465 67.020 21.585 ;
        RECT 67.260 21.295 67.525 21.755 ;
        RECT 67.695 21.160 67.945 21.585 ;
        RECT 68.155 21.310 69.260 21.480 ;
        RECT 67.640 21.030 67.945 21.160 ;
        RECT 67.190 19.835 67.470 20.785 ;
        RECT 67.640 19.925 67.810 21.030 ;
        RECT 67.980 20.245 68.220 20.840 ;
        RECT 68.390 20.775 68.920 21.140 ;
        RECT 68.390 20.075 68.560 20.775 ;
        RECT 69.090 20.695 69.260 21.310 ;
        RECT 69.430 20.955 69.600 21.755 ;
        RECT 69.770 21.255 70.020 21.585 ;
        RECT 70.245 21.285 71.130 21.455 ;
        RECT 69.090 20.605 69.600 20.695 ;
        RECT 67.640 19.795 67.865 19.925 ;
        RECT 68.035 19.855 68.560 20.075 ;
        RECT 68.730 20.435 69.600 20.605 ;
        RECT 67.275 19.205 67.525 19.665 ;
        RECT 67.695 19.655 67.865 19.795 ;
        RECT 68.730 19.655 68.900 20.435 ;
        RECT 69.430 20.365 69.600 20.435 ;
        RECT 69.110 20.185 69.310 20.215 ;
        RECT 69.770 20.185 69.940 21.255 ;
        RECT 70.110 20.365 70.300 21.085 ;
        RECT 69.110 19.885 69.940 20.185 ;
        RECT 70.470 20.155 70.790 21.115 ;
        RECT 67.695 19.485 68.030 19.655 ;
        RECT 68.225 19.485 68.900 19.655 ;
        RECT 69.220 19.205 69.590 19.705 ;
        RECT 69.770 19.655 69.940 19.885 ;
        RECT 70.325 19.825 70.790 20.155 ;
        RECT 70.960 20.445 71.130 21.285 ;
        RECT 71.310 21.255 71.625 21.755 ;
        RECT 71.855 21.025 72.195 21.585 ;
        RECT 71.300 20.650 72.195 21.025 ;
        RECT 72.365 20.745 72.535 21.755 ;
        RECT 72.005 20.445 72.195 20.650 ;
        RECT 72.705 20.695 73.035 21.540 ;
        RECT 72.705 20.615 73.095 20.695 ;
        RECT 72.880 20.565 73.095 20.615 ;
        RECT 70.960 20.115 71.835 20.445 ;
        RECT 72.005 20.115 72.755 20.445 ;
        RECT 70.960 19.655 71.130 20.115 ;
        RECT 72.005 19.945 72.205 20.115 ;
        RECT 72.925 19.985 73.095 20.565 ;
        RECT 72.870 19.945 73.095 19.985 ;
        RECT 69.770 19.485 70.175 19.655 ;
        RECT 70.345 19.485 71.130 19.655 ;
        RECT 71.405 19.205 71.615 19.735 ;
        RECT 71.875 19.420 72.205 19.945 ;
        RECT 72.715 19.860 73.095 19.945 ;
        RECT 73.265 20.615 73.605 21.585 ;
        RECT 73.775 20.615 73.945 21.755 ;
        RECT 74.215 20.955 74.465 21.755 ;
        RECT 75.110 20.785 75.440 21.585 ;
        RECT 75.740 20.955 76.070 21.755 ;
        RECT 76.240 20.785 76.570 21.585 ;
        RECT 74.135 20.615 76.570 20.785 ;
        RECT 73.265 20.005 73.440 20.615 ;
        RECT 74.135 20.365 74.305 20.615 ;
        RECT 73.610 20.195 74.305 20.365 ;
        RECT 74.480 20.195 74.900 20.395 ;
        RECT 75.070 20.195 75.400 20.395 ;
        RECT 75.570 20.195 75.900 20.395 ;
        RECT 72.375 19.205 72.545 19.815 ;
        RECT 72.715 19.425 73.045 19.860 ;
        RECT 73.265 19.375 73.605 20.005 ;
        RECT 73.775 19.205 74.025 20.005 ;
        RECT 74.215 19.855 75.440 20.025 ;
        RECT 74.215 19.375 74.545 19.855 ;
        RECT 74.715 19.205 74.940 19.665 ;
        RECT 75.110 19.375 75.440 19.855 ;
        RECT 76.070 19.985 76.240 20.615 ;
        RECT 77.865 20.590 78.155 21.755 ;
        RECT 78.990 20.785 79.320 21.585 ;
        RECT 79.490 20.955 79.820 21.755 ;
        RECT 80.120 20.785 80.450 21.585 ;
        RECT 81.095 20.955 81.345 21.755 ;
        RECT 78.990 20.615 81.425 20.785 ;
        RECT 81.615 20.615 81.785 21.755 ;
        RECT 81.955 20.615 82.295 21.585 ;
        RECT 82.670 20.785 83.000 21.585 ;
        RECT 83.170 20.955 83.500 21.755 ;
        RECT 83.800 20.785 84.130 21.585 ;
        RECT 84.775 20.955 85.025 21.755 ;
        RECT 82.670 20.615 85.105 20.785 ;
        RECT 85.295 20.615 85.465 21.755 ;
        RECT 85.635 20.615 85.975 21.585 ;
        RECT 86.235 20.825 86.405 21.585 ;
        RECT 86.620 20.995 86.950 21.755 ;
        RECT 86.235 20.655 86.950 20.825 ;
        RECT 87.120 20.680 87.375 21.585 ;
        RECT 76.425 20.195 76.775 20.445 ;
        RECT 78.785 20.195 79.135 20.445 ;
        RECT 79.320 19.985 79.490 20.615 ;
        RECT 79.660 20.195 79.990 20.395 ;
        RECT 80.160 20.195 80.490 20.395 ;
        RECT 80.660 20.195 81.080 20.395 ;
        RECT 81.255 20.365 81.425 20.615 ;
        RECT 81.255 20.195 81.950 20.365 ;
        RECT 76.070 19.375 76.570 19.985 ;
        RECT 77.865 19.205 78.155 19.930 ;
        RECT 78.990 19.375 79.490 19.985 ;
        RECT 80.120 19.855 81.345 20.025 ;
        RECT 82.120 20.005 82.295 20.615 ;
        RECT 82.465 20.195 82.815 20.445 ;
        RECT 80.120 19.375 80.450 19.855 ;
        RECT 80.620 19.205 80.845 19.665 ;
        RECT 81.015 19.375 81.345 19.855 ;
        RECT 81.535 19.205 81.785 20.005 ;
        RECT 81.955 19.375 82.295 20.005 ;
        RECT 83.000 19.985 83.170 20.615 ;
        RECT 83.340 20.195 83.670 20.395 ;
        RECT 83.840 20.195 84.170 20.395 ;
        RECT 84.340 20.195 84.760 20.395 ;
        RECT 84.935 20.365 85.105 20.615 ;
        RECT 84.935 20.195 85.630 20.365 ;
        RECT 82.670 19.375 83.170 19.985 ;
        RECT 83.800 19.855 85.025 20.025 ;
        RECT 85.800 20.005 85.975 20.615 ;
        RECT 86.145 20.105 86.500 20.475 ;
        RECT 86.780 20.445 86.950 20.655 ;
        RECT 86.780 20.115 87.035 20.445 ;
        RECT 83.800 19.375 84.130 19.855 ;
        RECT 84.300 19.205 84.525 19.665 ;
        RECT 84.695 19.375 85.025 19.855 ;
        RECT 85.215 19.205 85.465 20.005 ;
        RECT 85.635 19.375 85.975 20.005 ;
        RECT 86.780 19.925 86.950 20.115 ;
        RECT 87.205 19.950 87.375 20.680 ;
        RECT 87.550 20.605 87.810 21.755 ;
        RECT 88.075 20.825 88.245 21.585 ;
        RECT 88.460 20.995 88.790 21.755 ;
        RECT 88.075 20.655 88.790 20.825 ;
        RECT 88.960 20.680 89.215 21.585 ;
        RECT 87.985 20.105 88.340 20.475 ;
        RECT 88.620 20.445 88.790 20.655 ;
        RECT 88.620 20.115 88.875 20.445 ;
        RECT 86.235 19.755 86.950 19.925 ;
        RECT 86.235 19.375 86.405 19.755 ;
        RECT 86.620 19.205 86.950 19.585 ;
        RECT 87.120 19.375 87.375 19.950 ;
        RECT 87.550 19.205 87.810 20.045 ;
        RECT 88.620 19.925 88.790 20.115 ;
        RECT 89.045 19.950 89.215 20.680 ;
        RECT 89.390 20.605 89.650 21.755 ;
        RECT 90.745 20.665 91.955 21.755 ;
        RECT 90.745 20.125 91.265 20.665 ;
        RECT 88.075 19.755 88.790 19.925 ;
        RECT 88.075 19.375 88.245 19.755 ;
        RECT 88.460 19.205 88.790 19.585 ;
        RECT 88.960 19.375 89.215 19.950 ;
        RECT 89.390 19.205 89.650 20.045 ;
        RECT 91.435 19.955 91.955 20.495 ;
        RECT 90.745 19.205 91.955 19.955 ;
        RECT 13.380 19.035 92.040 19.205 ;
        RECT 13.465 18.285 14.675 19.035 ;
        RECT 15.930 18.525 16.170 19.035 ;
        RECT 16.350 18.525 16.630 18.855 ;
        RECT 16.860 18.525 17.075 19.035 ;
        RECT 13.465 17.745 13.985 18.285 ;
        RECT 14.155 17.575 14.675 18.115 ;
        RECT 15.825 17.795 16.180 18.355 ;
        RECT 16.350 17.625 16.520 18.525 ;
        RECT 16.690 17.795 16.955 18.355 ;
        RECT 17.245 18.295 17.860 18.865 ;
        RECT 17.205 17.625 17.375 18.125 ;
        RECT 13.465 16.485 14.675 17.575 ;
        RECT 15.950 17.455 17.375 17.625 ;
        RECT 15.950 17.280 16.340 17.455 ;
        RECT 16.825 16.485 17.155 17.285 ;
        RECT 17.545 17.275 17.860 18.295 ;
        RECT 18.065 18.285 19.275 19.035 ;
        RECT 19.535 18.485 19.705 18.775 ;
        RECT 19.875 18.655 20.205 19.035 ;
        RECT 19.535 18.315 20.200 18.485 ;
        RECT 18.065 17.745 18.585 18.285 ;
        RECT 18.755 17.575 19.275 18.115 ;
        RECT 17.325 16.655 17.860 17.275 ;
        RECT 18.065 16.485 19.275 17.575 ;
        RECT 19.450 17.495 19.800 18.145 ;
        RECT 19.970 17.325 20.200 18.315 ;
        RECT 19.535 17.155 20.200 17.325 ;
        RECT 19.535 16.655 19.705 17.155 ;
        RECT 19.875 16.485 20.205 16.985 ;
        RECT 20.375 16.655 20.560 18.775 ;
        RECT 20.815 18.575 21.065 19.035 ;
        RECT 21.235 18.585 21.570 18.755 ;
        RECT 21.765 18.585 22.440 18.755 ;
        RECT 21.235 18.445 21.405 18.585 ;
        RECT 20.730 17.455 21.010 18.405 ;
        RECT 21.180 18.315 21.405 18.445 ;
        RECT 21.180 17.210 21.350 18.315 ;
        RECT 21.575 18.165 22.100 18.385 ;
        RECT 21.520 17.400 21.760 17.995 ;
        RECT 21.930 17.465 22.100 18.165 ;
        RECT 22.270 17.805 22.440 18.585 ;
        RECT 22.760 18.535 23.130 19.035 ;
        RECT 23.310 18.585 23.715 18.755 ;
        RECT 23.885 18.585 24.670 18.755 ;
        RECT 23.310 18.355 23.480 18.585 ;
        RECT 22.650 18.055 23.480 18.355 ;
        RECT 23.865 18.085 24.330 18.415 ;
        RECT 22.650 18.025 22.850 18.055 ;
        RECT 22.970 17.805 23.140 17.875 ;
        RECT 22.270 17.635 23.140 17.805 ;
        RECT 22.630 17.545 23.140 17.635 ;
        RECT 21.180 17.080 21.485 17.210 ;
        RECT 21.930 17.100 22.460 17.465 ;
        RECT 20.800 16.485 21.065 16.945 ;
        RECT 21.235 16.655 21.485 17.080 ;
        RECT 22.630 16.930 22.800 17.545 ;
        RECT 21.695 16.760 22.800 16.930 ;
        RECT 22.970 16.485 23.140 17.285 ;
        RECT 23.310 16.985 23.480 18.055 ;
        RECT 23.650 17.155 23.840 17.875 ;
        RECT 24.010 17.125 24.330 18.085 ;
        RECT 24.500 18.125 24.670 18.585 ;
        RECT 24.945 18.505 25.155 19.035 ;
        RECT 25.415 18.295 25.745 18.820 ;
        RECT 25.915 18.425 26.085 19.035 ;
        RECT 26.255 18.380 26.585 18.815 ;
        RECT 26.970 18.525 27.210 19.035 ;
        RECT 27.390 18.525 27.670 18.855 ;
        RECT 27.900 18.525 28.115 19.035 ;
        RECT 26.255 18.295 26.635 18.380 ;
        RECT 25.545 18.125 25.745 18.295 ;
        RECT 26.410 18.255 26.635 18.295 ;
        RECT 24.500 17.795 25.375 18.125 ;
        RECT 25.545 17.795 26.295 18.125 ;
        RECT 23.310 16.655 23.560 16.985 ;
        RECT 24.500 16.955 24.670 17.795 ;
        RECT 25.545 17.590 25.735 17.795 ;
        RECT 26.465 17.675 26.635 18.255 ;
        RECT 26.865 17.795 27.220 18.355 ;
        RECT 26.420 17.625 26.635 17.675 ;
        RECT 27.390 17.625 27.560 18.525 ;
        RECT 27.730 17.795 27.995 18.355 ;
        RECT 28.285 18.295 28.900 18.865 ;
        RECT 29.195 18.485 29.365 18.775 ;
        RECT 29.535 18.655 29.865 19.035 ;
        RECT 29.195 18.315 29.860 18.485 ;
        RECT 28.245 17.625 28.415 18.125 ;
        RECT 24.840 17.215 25.735 17.590 ;
        RECT 26.245 17.545 26.635 17.625 ;
        RECT 23.785 16.785 24.670 16.955 ;
        RECT 24.850 16.485 25.165 16.985 ;
        RECT 25.395 16.655 25.735 17.215 ;
        RECT 25.905 16.485 26.075 17.495 ;
        RECT 26.245 16.700 26.575 17.545 ;
        RECT 26.990 17.455 28.415 17.625 ;
        RECT 26.990 17.280 27.380 17.455 ;
        RECT 27.865 16.485 28.195 17.285 ;
        RECT 28.585 17.275 28.900 18.295 ;
        RECT 29.110 17.495 29.460 18.145 ;
        RECT 29.630 17.325 29.860 18.315 ;
        RECT 28.365 16.655 28.900 17.275 ;
        RECT 29.195 17.155 29.860 17.325 ;
        RECT 29.195 16.655 29.365 17.155 ;
        RECT 29.535 16.485 29.865 16.985 ;
        RECT 30.035 16.655 30.220 18.775 ;
        RECT 30.475 18.575 30.725 19.035 ;
        RECT 30.895 18.585 31.230 18.755 ;
        RECT 31.425 18.585 32.100 18.755 ;
        RECT 30.895 18.445 31.065 18.585 ;
        RECT 30.390 17.455 30.670 18.405 ;
        RECT 30.840 18.315 31.065 18.445 ;
        RECT 30.840 17.210 31.010 18.315 ;
        RECT 31.235 18.165 31.760 18.385 ;
        RECT 31.180 17.400 31.420 17.995 ;
        RECT 31.590 17.465 31.760 18.165 ;
        RECT 31.930 17.805 32.100 18.585 ;
        RECT 32.420 18.535 32.790 19.035 ;
        RECT 32.970 18.585 33.375 18.755 ;
        RECT 33.545 18.585 34.330 18.755 ;
        RECT 32.970 18.355 33.140 18.585 ;
        RECT 32.310 18.055 33.140 18.355 ;
        RECT 33.525 18.085 33.990 18.415 ;
        RECT 32.310 18.025 32.510 18.055 ;
        RECT 32.630 17.805 32.800 17.875 ;
        RECT 31.930 17.635 32.800 17.805 ;
        RECT 32.290 17.545 32.800 17.635 ;
        RECT 30.840 17.080 31.145 17.210 ;
        RECT 31.590 17.100 32.120 17.465 ;
        RECT 30.460 16.485 30.725 16.945 ;
        RECT 30.895 16.655 31.145 17.080 ;
        RECT 32.290 16.930 32.460 17.545 ;
        RECT 31.355 16.760 32.460 16.930 ;
        RECT 32.630 16.485 32.800 17.285 ;
        RECT 32.970 16.985 33.140 18.055 ;
        RECT 33.310 17.155 33.500 17.875 ;
        RECT 33.670 17.125 33.990 18.085 ;
        RECT 34.160 18.125 34.330 18.585 ;
        RECT 34.605 18.505 34.815 19.035 ;
        RECT 35.075 18.295 35.405 18.820 ;
        RECT 35.575 18.425 35.745 19.035 ;
        RECT 35.915 18.380 36.245 18.815 ;
        RECT 35.915 18.295 36.295 18.380 ;
        RECT 35.205 18.125 35.405 18.295 ;
        RECT 36.070 18.255 36.295 18.295 ;
        RECT 34.160 17.795 35.035 18.125 ;
        RECT 35.205 17.795 35.955 18.125 ;
        RECT 32.970 16.655 33.220 16.985 ;
        RECT 34.160 16.955 34.330 17.795 ;
        RECT 35.205 17.590 35.395 17.795 ;
        RECT 36.125 17.675 36.295 18.255 ;
        RECT 36.080 17.625 36.295 17.675 ;
        RECT 34.500 17.215 35.395 17.590 ;
        RECT 35.905 17.545 36.295 17.625 ;
        RECT 36.500 18.295 37.115 18.865 ;
        RECT 37.285 18.525 37.500 19.035 ;
        RECT 37.730 18.525 38.010 18.855 ;
        RECT 38.190 18.525 38.430 19.035 ;
        RECT 33.445 16.785 34.330 16.955 ;
        RECT 34.510 16.485 34.825 16.985 ;
        RECT 35.055 16.655 35.395 17.215 ;
        RECT 35.565 16.485 35.735 17.495 ;
        RECT 35.905 16.700 36.235 17.545 ;
        RECT 36.500 17.275 36.815 18.295 ;
        RECT 36.985 17.625 37.155 18.125 ;
        RECT 37.405 17.795 37.670 18.355 ;
        RECT 37.840 17.625 38.010 18.525 ;
        RECT 38.180 17.795 38.535 18.355 ;
        RECT 39.225 18.310 39.515 19.035 ;
        RECT 40.195 18.380 40.525 18.815 ;
        RECT 40.695 18.425 40.865 19.035 ;
        RECT 40.145 18.295 40.525 18.380 ;
        RECT 41.035 18.295 41.365 18.820 ;
        RECT 41.625 18.505 41.835 19.035 ;
        RECT 42.110 18.585 42.895 18.755 ;
        RECT 43.065 18.585 43.470 18.755 ;
        RECT 40.145 18.255 40.370 18.295 ;
        RECT 40.145 17.675 40.315 18.255 ;
        RECT 41.035 18.125 41.235 18.295 ;
        RECT 42.110 18.125 42.280 18.585 ;
        RECT 40.485 17.795 41.235 18.125 ;
        RECT 41.405 17.795 42.280 18.125 ;
        RECT 36.985 17.455 38.410 17.625 ;
        RECT 36.500 16.655 37.035 17.275 ;
        RECT 37.205 16.485 37.535 17.285 ;
        RECT 38.020 17.280 38.410 17.455 ;
        RECT 39.225 16.485 39.515 17.650 ;
        RECT 40.145 17.625 40.360 17.675 ;
        RECT 40.145 17.545 40.535 17.625 ;
        RECT 40.205 16.700 40.535 17.545 ;
        RECT 41.045 17.590 41.235 17.795 ;
        RECT 40.705 16.485 40.875 17.495 ;
        RECT 41.045 17.215 41.940 17.590 ;
        RECT 41.045 16.655 41.385 17.215 ;
        RECT 41.615 16.485 41.930 16.985 ;
        RECT 42.110 16.955 42.280 17.795 ;
        RECT 42.450 18.085 42.915 18.415 ;
        RECT 43.300 18.355 43.470 18.585 ;
        RECT 43.650 18.535 44.020 19.035 ;
        RECT 44.340 18.585 45.015 18.755 ;
        RECT 45.210 18.585 45.545 18.755 ;
        RECT 42.450 17.125 42.770 18.085 ;
        RECT 43.300 18.055 44.130 18.355 ;
        RECT 42.940 17.155 43.130 17.875 ;
        RECT 43.300 16.985 43.470 18.055 ;
        RECT 43.930 18.025 44.130 18.055 ;
        RECT 43.640 17.805 43.810 17.875 ;
        RECT 44.340 17.805 44.510 18.585 ;
        RECT 45.375 18.445 45.545 18.585 ;
        RECT 45.715 18.575 45.965 19.035 ;
        RECT 43.640 17.635 44.510 17.805 ;
        RECT 44.680 18.165 45.205 18.385 ;
        RECT 45.375 18.315 45.600 18.445 ;
        RECT 43.640 17.545 44.150 17.635 ;
        RECT 42.110 16.785 42.995 16.955 ;
        RECT 43.220 16.655 43.470 16.985 ;
        RECT 43.640 16.485 43.810 17.285 ;
        RECT 43.980 16.930 44.150 17.545 ;
        RECT 44.680 17.465 44.850 18.165 ;
        RECT 44.320 17.100 44.850 17.465 ;
        RECT 45.020 17.400 45.260 17.995 ;
        RECT 45.430 17.210 45.600 18.315 ;
        RECT 45.770 17.455 46.050 18.405 ;
        RECT 45.295 17.080 45.600 17.210 ;
        RECT 43.980 16.760 45.085 16.930 ;
        RECT 45.295 16.655 45.545 17.080 ;
        RECT 45.715 16.485 45.980 16.945 ;
        RECT 46.220 16.655 46.405 18.775 ;
        RECT 46.575 18.655 46.905 19.035 ;
        RECT 47.075 18.485 47.245 18.775 ;
        RECT 46.580 18.315 47.245 18.485 ;
        RECT 48.055 18.485 48.225 18.775 ;
        RECT 48.395 18.655 48.725 19.035 ;
        RECT 48.055 18.315 48.720 18.485 ;
        RECT 46.580 17.325 46.810 18.315 ;
        RECT 46.980 17.495 47.330 18.145 ;
        RECT 47.970 17.495 48.320 18.145 ;
        RECT 48.490 17.325 48.720 18.315 ;
        RECT 46.580 17.155 47.245 17.325 ;
        RECT 46.575 16.485 46.905 16.985 ;
        RECT 47.075 16.655 47.245 17.155 ;
        RECT 48.055 17.155 48.720 17.325 ;
        RECT 48.055 16.655 48.225 17.155 ;
        RECT 48.395 16.485 48.725 16.985 ;
        RECT 48.895 16.655 49.080 18.775 ;
        RECT 49.335 18.575 49.585 19.035 ;
        RECT 49.755 18.585 50.090 18.755 ;
        RECT 50.285 18.585 50.960 18.755 ;
        RECT 49.755 18.445 49.925 18.585 ;
        RECT 49.250 17.455 49.530 18.405 ;
        RECT 49.700 18.315 49.925 18.445 ;
        RECT 49.700 17.210 49.870 18.315 ;
        RECT 50.095 18.165 50.620 18.385 ;
        RECT 50.040 17.400 50.280 17.995 ;
        RECT 50.450 17.465 50.620 18.165 ;
        RECT 50.790 17.805 50.960 18.585 ;
        RECT 51.280 18.535 51.650 19.035 ;
        RECT 51.830 18.585 52.235 18.755 ;
        RECT 52.405 18.585 53.190 18.755 ;
        RECT 51.830 18.355 52.000 18.585 ;
        RECT 51.170 18.055 52.000 18.355 ;
        RECT 52.385 18.085 52.850 18.415 ;
        RECT 51.170 18.025 51.370 18.055 ;
        RECT 51.490 17.805 51.660 17.875 ;
        RECT 50.790 17.635 51.660 17.805 ;
        RECT 51.150 17.545 51.660 17.635 ;
        RECT 49.700 17.080 50.005 17.210 ;
        RECT 50.450 17.100 50.980 17.465 ;
        RECT 49.320 16.485 49.585 16.945 ;
        RECT 49.755 16.655 50.005 17.080 ;
        RECT 51.150 16.930 51.320 17.545 ;
        RECT 50.215 16.760 51.320 16.930 ;
        RECT 51.490 16.485 51.660 17.285 ;
        RECT 51.830 16.985 52.000 18.055 ;
        RECT 52.170 17.155 52.360 17.875 ;
        RECT 52.530 17.125 52.850 18.085 ;
        RECT 53.020 18.125 53.190 18.585 ;
        RECT 53.465 18.505 53.675 19.035 ;
        RECT 53.935 18.295 54.265 18.820 ;
        RECT 54.435 18.425 54.605 19.035 ;
        RECT 54.775 18.380 55.105 18.815 ;
        RECT 55.415 18.485 55.585 18.775 ;
        RECT 55.755 18.655 56.085 19.035 ;
        RECT 54.775 18.295 55.155 18.380 ;
        RECT 55.415 18.315 56.080 18.485 ;
        RECT 54.065 18.125 54.265 18.295 ;
        RECT 54.930 18.255 55.155 18.295 ;
        RECT 53.020 17.795 53.895 18.125 ;
        RECT 54.065 17.795 54.815 18.125 ;
        RECT 51.830 16.655 52.080 16.985 ;
        RECT 53.020 16.955 53.190 17.795 ;
        RECT 54.065 17.590 54.255 17.795 ;
        RECT 54.985 17.675 55.155 18.255 ;
        RECT 54.940 17.625 55.155 17.675 ;
        RECT 53.360 17.215 54.255 17.590 ;
        RECT 54.765 17.545 55.155 17.625 ;
        RECT 52.305 16.785 53.190 16.955 ;
        RECT 53.370 16.485 53.685 16.985 ;
        RECT 53.915 16.655 54.255 17.215 ;
        RECT 54.425 16.485 54.595 17.495 ;
        RECT 54.765 16.700 55.095 17.545 ;
        RECT 55.330 17.495 55.680 18.145 ;
        RECT 55.850 17.325 56.080 18.315 ;
        RECT 55.415 17.155 56.080 17.325 ;
        RECT 55.415 16.655 55.585 17.155 ;
        RECT 55.755 16.485 56.085 16.985 ;
        RECT 56.255 16.655 56.440 18.775 ;
        RECT 56.695 18.575 56.945 19.035 ;
        RECT 57.115 18.585 57.450 18.755 ;
        RECT 57.645 18.585 58.320 18.755 ;
        RECT 57.115 18.445 57.285 18.585 ;
        RECT 56.610 17.455 56.890 18.405 ;
        RECT 57.060 18.315 57.285 18.445 ;
        RECT 57.060 17.210 57.230 18.315 ;
        RECT 57.455 18.165 57.980 18.385 ;
        RECT 57.400 17.400 57.640 17.995 ;
        RECT 57.810 17.465 57.980 18.165 ;
        RECT 58.150 17.805 58.320 18.585 ;
        RECT 58.640 18.535 59.010 19.035 ;
        RECT 59.190 18.585 59.595 18.755 ;
        RECT 59.765 18.585 60.550 18.755 ;
        RECT 59.190 18.355 59.360 18.585 ;
        RECT 58.530 18.055 59.360 18.355 ;
        RECT 59.745 18.085 60.210 18.415 ;
        RECT 58.530 18.025 58.730 18.055 ;
        RECT 58.850 17.805 59.020 17.875 ;
        RECT 58.150 17.635 59.020 17.805 ;
        RECT 58.510 17.545 59.020 17.635 ;
        RECT 57.060 17.080 57.365 17.210 ;
        RECT 57.810 17.100 58.340 17.465 ;
        RECT 56.680 16.485 56.945 16.945 ;
        RECT 57.115 16.655 57.365 17.080 ;
        RECT 58.510 16.930 58.680 17.545 ;
        RECT 57.575 16.760 58.680 16.930 ;
        RECT 58.850 16.485 59.020 17.285 ;
        RECT 59.190 16.985 59.360 18.055 ;
        RECT 59.530 17.155 59.720 17.875 ;
        RECT 59.890 17.125 60.210 18.085 ;
        RECT 60.380 18.125 60.550 18.585 ;
        RECT 60.825 18.505 61.035 19.035 ;
        RECT 61.295 18.295 61.625 18.820 ;
        RECT 61.795 18.425 61.965 19.035 ;
        RECT 62.135 18.380 62.465 18.815 ;
        RECT 62.135 18.295 62.515 18.380 ;
        RECT 61.425 18.125 61.625 18.295 ;
        RECT 62.290 18.255 62.515 18.295 ;
        RECT 60.380 17.795 61.255 18.125 ;
        RECT 61.425 17.795 62.175 18.125 ;
        RECT 59.190 16.655 59.440 16.985 ;
        RECT 60.380 16.955 60.550 17.795 ;
        RECT 61.425 17.590 61.615 17.795 ;
        RECT 62.345 17.675 62.515 18.255 ;
        RECT 62.300 17.625 62.515 17.675 ;
        RECT 60.720 17.215 61.615 17.590 ;
        RECT 62.125 17.545 62.515 17.625 ;
        RECT 62.720 18.295 63.335 18.865 ;
        RECT 63.505 18.525 63.720 19.035 ;
        RECT 63.950 18.525 64.230 18.855 ;
        RECT 64.410 18.525 64.650 19.035 ;
        RECT 59.665 16.785 60.550 16.955 ;
        RECT 60.730 16.485 61.045 16.985 ;
        RECT 61.275 16.655 61.615 17.215 ;
        RECT 61.785 16.485 61.955 17.495 ;
        RECT 62.125 16.700 62.455 17.545 ;
        RECT 62.720 17.275 63.035 18.295 ;
        RECT 63.205 17.625 63.375 18.125 ;
        RECT 63.625 17.795 63.890 18.355 ;
        RECT 64.060 17.625 64.230 18.525 ;
        RECT 64.400 17.795 64.755 18.355 ;
        RECT 64.985 18.310 65.275 19.035 ;
        RECT 65.445 18.535 65.705 18.865 ;
        RECT 65.875 18.675 66.205 19.035 ;
        RECT 66.460 18.655 67.760 18.865 ;
        RECT 63.205 17.455 64.630 17.625 ;
        RECT 62.720 16.655 63.255 17.275 ;
        RECT 63.425 16.485 63.755 17.285 ;
        RECT 64.240 17.280 64.630 17.455 ;
        RECT 64.985 16.485 65.275 17.650 ;
        RECT 65.445 17.335 65.615 18.535 ;
        RECT 66.460 18.505 66.630 18.655 ;
        RECT 65.875 18.380 66.630 18.505 ;
        RECT 65.785 18.335 66.630 18.380 ;
        RECT 65.785 18.215 66.055 18.335 ;
        RECT 65.785 17.640 65.955 18.215 ;
        RECT 66.185 17.775 66.595 18.080 ;
        RECT 66.885 18.045 67.095 18.445 ;
        RECT 66.765 17.835 67.095 18.045 ;
        RECT 67.340 18.045 67.560 18.445 ;
        RECT 68.035 18.270 68.490 19.035 ;
        RECT 68.665 18.285 69.875 19.035 ;
        RECT 70.135 18.485 70.305 18.775 ;
        RECT 70.475 18.655 70.805 19.035 ;
        RECT 70.135 18.315 70.800 18.485 ;
        RECT 67.340 17.835 67.815 18.045 ;
        RECT 68.005 17.845 68.495 18.045 ;
        RECT 68.665 17.745 69.185 18.285 ;
        RECT 65.785 17.605 65.985 17.640 ;
        RECT 67.315 17.605 68.490 17.665 ;
        RECT 65.785 17.495 68.490 17.605 ;
        RECT 69.355 17.575 69.875 18.115 ;
        RECT 65.845 17.435 67.645 17.495 ;
        RECT 67.315 17.405 67.645 17.435 ;
        RECT 65.445 16.655 65.705 17.335 ;
        RECT 65.875 16.485 66.125 17.265 ;
        RECT 66.375 17.235 67.210 17.245 ;
        RECT 67.800 17.235 67.985 17.325 ;
        RECT 66.375 17.035 67.985 17.235 ;
        RECT 66.375 16.655 66.625 17.035 ;
        RECT 67.755 16.995 67.985 17.035 ;
        RECT 68.235 16.875 68.490 17.495 ;
        RECT 66.795 16.485 67.150 16.865 ;
        RECT 68.155 16.655 68.490 16.875 ;
        RECT 68.665 16.485 69.875 17.575 ;
        RECT 70.050 17.495 70.400 18.145 ;
        RECT 70.570 17.325 70.800 18.315 ;
        RECT 70.135 17.155 70.800 17.325 ;
        RECT 70.135 16.655 70.305 17.155 ;
        RECT 70.475 16.485 70.805 16.985 ;
        RECT 70.975 16.655 71.160 18.775 ;
        RECT 71.415 18.575 71.665 19.035 ;
        RECT 71.835 18.585 72.170 18.755 ;
        RECT 72.365 18.585 73.040 18.755 ;
        RECT 71.835 18.445 72.005 18.585 ;
        RECT 71.330 17.455 71.610 18.405 ;
        RECT 71.780 18.315 72.005 18.445 ;
        RECT 71.780 17.210 71.950 18.315 ;
        RECT 72.175 18.165 72.700 18.385 ;
        RECT 72.120 17.400 72.360 17.995 ;
        RECT 72.530 17.465 72.700 18.165 ;
        RECT 72.870 17.805 73.040 18.585 ;
        RECT 73.360 18.535 73.730 19.035 ;
        RECT 73.910 18.585 74.315 18.755 ;
        RECT 74.485 18.585 75.270 18.755 ;
        RECT 73.910 18.355 74.080 18.585 ;
        RECT 73.250 18.055 74.080 18.355 ;
        RECT 74.465 18.085 74.930 18.415 ;
        RECT 73.250 18.025 73.450 18.055 ;
        RECT 73.570 17.805 73.740 17.875 ;
        RECT 72.870 17.635 73.740 17.805 ;
        RECT 73.230 17.545 73.740 17.635 ;
        RECT 71.780 17.080 72.085 17.210 ;
        RECT 72.530 17.100 73.060 17.465 ;
        RECT 71.400 16.485 71.665 16.945 ;
        RECT 71.835 16.655 72.085 17.080 ;
        RECT 73.230 16.930 73.400 17.545 ;
        RECT 72.295 16.760 73.400 16.930 ;
        RECT 73.570 16.485 73.740 17.285 ;
        RECT 73.910 16.985 74.080 18.055 ;
        RECT 74.250 17.155 74.440 17.875 ;
        RECT 74.610 17.125 74.930 18.085 ;
        RECT 75.100 18.125 75.270 18.585 ;
        RECT 75.545 18.505 75.755 19.035 ;
        RECT 76.015 18.295 76.345 18.820 ;
        RECT 76.515 18.425 76.685 19.035 ;
        RECT 76.855 18.380 77.185 18.815 ;
        RECT 77.570 18.525 77.810 19.035 ;
        RECT 77.990 18.525 78.270 18.855 ;
        RECT 78.500 18.525 78.715 19.035 ;
        RECT 76.855 18.295 77.235 18.380 ;
        RECT 76.145 18.125 76.345 18.295 ;
        RECT 77.010 18.255 77.235 18.295 ;
        RECT 75.100 17.795 75.975 18.125 ;
        RECT 76.145 17.795 76.895 18.125 ;
        RECT 73.910 16.655 74.160 16.985 ;
        RECT 75.100 16.955 75.270 17.795 ;
        RECT 76.145 17.590 76.335 17.795 ;
        RECT 77.065 17.675 77.235 18.255 ;
        RECT 77.465 17.795 77.820 18.355 ;
        RECT 77.020 17.625 77.235 17.675 ;
        RECT 77.990 17.625 78.160 18.525 ;
        RECT 78.330 17.795 78.595 18.355 ;
        RECT 78.885 18.295 79.500 18.865 ;
        RECT 78.845 17.625 79.015 18.125 ;
        RECT 75.440 17.215 76.335 17.590 ;
        RECT 76.845 17.545 77.235 17.625 ;
        RECT 74.385 16.785 75.270 16.955 ;
        RECT 75.450 16.485 75.765 16.985 ;
        RECT 75.995 16.655 76.335 17.215 ;
        RECT 76.505 16.485 76.675 17.495 ;
        RECT 76.845 16.700 77.175 17.545 ;
        RECT 77.590 17.455 79.015 17.625 ;
        RECT 77.590 17.280 77.980 17.455 ;
        RECT 78.465 16.485 78.795 17.285 ;
        RECT 79.185 17.275 79.500 18.295 ;
        RECT 79.705 18.285 80.915 19.035 ;
        RECT 81.175 18.485 81.345 18.775 ;
        RECT 81.515 18.655 81.845 19.035 ;
        RECT 81.175 18.315 81.840 18.485 ;
        RECT 79.705 17.745 80.225 18.285 ;
        RECT 80.395 17.575 80.915 18.115 ;
        RECT 78.965 16.655 79.500 17.275 ;
        RECT 79.705 16.485 80.915 17.575 ;
        RECT 81.090 17.495 81.440 18.145 ;
        RECT 81.610 17.325 81.840 18.315 ;
        RECT 81.175 17.155 81.840 17.325 ;
        RECT 81.175 16.655 81.345 17.155 ;
        RECT 81.515 16.485 81.845 16.985 ;
        RECT 82.015 16.655 82.200 18.775 ;
        RECT 82.455 18.575 82.705 19.035 ;
        RECT 82.875 18.585 83.210 18.755 ;
        RECT 83.405 18.585 84.080 18.755 ;
        RECT 82.875 18.445 83.045 18.585 ;
        RECT 82.370 17.455 82.650 18.405 ;
        RECT 82.820 18.315 83.045 18.445 ;
        RECT 82.820 17.210 82.990 18.315 ;
        RECT 83.215 18.165 83.740 18.385 ;
        RECT 83.160 17.400 83.400 17.995 ;
        RECT 83.570 17.465 83.740 18.165 ;
        RECT 83.910 17.805 84.080 18.585 ;
        RECT 84.400 18.535 84.770 19.035 ;
        RECT 84.950 18.585 85.355 18.755 ;
        RECT 85.525 18.585 86.310 18.755 ;
        RECT 84.950 18.355 85.120 18.585 ;
        RECT 84.290 18.055 85.120 18.355 ;
        RECT 85.505 18.085 85.970 18.415 ;
        RECT 84.290 18.025 84.490 18.055 ;
        RECT 84.610 17.805 84.780 17.875 ;
        RECT 83.910 17.635 84.780 17.805 ;
        RECT 84.270 17.545 84.780 17.635 ;
        RECT 82.820 17.080 83.125 17.210 ;
        RECT 83.570 17.100 84.100 17.465 ;
        RECT 82.440 16.485 82.705 16.945 ;
        RECT 82.875 16.655 83.125 17.080 ;
        RECT 84.270 16.930 84.440 17.545 ;
        RECT 83.335 16.760 84.440 16.930 ;
        RECT 84.610 16.485 84.780 17.285 ;
        RECT 84.950 16.985 85.120 18.055 ;
        RECT 85.290 17.155 85.480 17.875 ;
        RECT 85.650 17.125 85.970 18.085 ;
        RECT 86.140 18.125 86.310 18.585 ;
        RECT 86.585 18.505 86.795 19.035 ;
        RECT 87.055 18.295 87.385 18.820 ;
        RECT 87.555 18.425 87.725 19.035 ;
        RECT 87.895 18.380 88.225 18.815 ;
        RECT 88.535 18.485 88.705 18.865 ;
        RECT 88.920 18.655 89.250 19.035 ;
        RECT 87.895 18.295 88.275 18.380 ;
        RECT 88.535 18.315 89.250 18.485 ;
        RECT 87.185 18.125 87.385 18.295 ;
        RECT 88.050 18.255 88.275 18.295 ;
        RECT 86.140 17.795 87.015 18.125 ;
        RECT 87.185 17.795 87.935 18.125 ;
        RECT 84.950 16.655 85.200 16.985 ;
        RECT 86.140 16.955 86.310 17.795 ;
        RECT 87.185 17.590 87.375 17.795 ;
        RECT 88.105 17.675 88.275 18.255 ;
        RECT 88.445 17.765 88.800 18.135 ;
        RECT 89.080 18.125 89.250 18.315 ;
        RECT 89.420 18.290 89.675 18.865 ;
        RECT 89.080 17.795 89.335 18.125 ;
        RECT 88.060 17.625 88.275 17.675 ;
        RECT 86.480 17.215 87.375 17.590 ;
        RECT 87.885 17.545 88.275 17.625 ;
        RECT 89.080 17.585 89.250 17.795 ;
        RECT 85.425 16.785 86.310 16.955 ;
        RECT 86.490 16.485 86.805 16.985 ;
        RECT 87.035 16.655 87.375 17.215 ;
        RECT 87.545 16.485 87.715 17.495 ;
        RECT 87.885 16.700 88.215 17.545 ;
        RECT 88.535 17.415 89.250 17.585 ;
        RECT 89.505 17.560 89.675 18.290 ;
        RECT 89.850 18.195 90.110 19.035 ;
        RECT 90.745 18.285 91.955 19.035 ;
        RECT 88.535 16.655 88.705 17.415 ;
        RECT 88.920 16.485 89.250 17.245 ;
        RECT 89.420 16.655 89.675 17.560 ;
        RECT 89.850 16.485 90.110 17.635 ;
        RECT 90.745 17.575 91.265 18.115 ;
        RECT 91.435 17.745 91.955 18.285 ;
        RECT 90.745 16.485 91.955 17.575 ;
        RECT 13.380 16.315 92.040 16.485 ;
        RECT 13.465 15.225 14.675 16.315 ;
        RECT 14.935 15.645 15.105 16.145 ;
        RECT 15.275 15.815 15.605 16.315 ;
        RECT 14.935 15.475 15.600 15.645 ;
        RECT 13.465 14.515 13.985 15.055 ;
        RECT 14.155 14.685 14.675 15.225 ;
        RECT 14.850 14.655 15.200 15.305 ;
        RECT 13.465 13.765 14.675 14.515 ;
        RECT 15.370 14.485 15.600 15.475 ;
        RECT 14.935 14.315 15.600 14.485 ;
        RECT 14.935 14.025 15.105 14.315 ;
        RECT 15.275 13.765 15.605 14.145 ;
        RECT 15.775 14.025 15.960 16.145 ;
        RECT 16.200 15.855 16.465 16.315 ;
        RECT 16.635 15.720 16.885 16.145 ;
        RECT 17.095 15.870 18.200 16.040 ;
        RECT 16.580 15.590 16.885 15.720 ;
        RECT 16.130 14.395 16.410 15.345 ;
        RECT 16.580 14.485 16.750 15.590 ;
        RECT 16.920 14.805 17.160 15.400 ;
        RECT 17.330 15.335 17.860 15.700 ;
        RECT 17.330 14.635 17.500 15.335 ;
        RECT 18.030 15.255 18.200 15.870 ;
        RECT 18.370 15.515 18.540 16.315 ;
        RECT 18.710 15.815 18.960 16.145 ;
        RECT 19.185 15.845 20.070 16.015 ;
        RECT 18.030 15.165 18.540 15.255 ;
        RECT 16.580 14.355 16.805 14.485 ;
        RECT 16.975 14.415 17.500 14.635 ;
        RECT 17.670 14.995 18.540 15.165 ;
        RECT 16.215 13.765 16.465 14.225 ;
        RECT 16.635 14.215 16.805 14.355 ;
        RECT 17.670 14.215 17.840 14.995 ;
        RECT 18.370 14.925 18.540 14.995 ;
        RECT 18.050 14.745 18.250 14.775 ;
        RECT 18.710 14.745 18.880 15.815 ;
        RECT 19.050 14.925 19.240 15.645 ;
        RECT 18.050 14.445 18.880 14.745 ;
        RECT 19.410 14.715 19.730 15.675 ;
        RECT 16.635 14.045 16.970 14.215 ;
        RECT 17.165 14.045 17.840 14.215 ;
        RECT 18.160 13.765 18.530 14.265 ;
        RECT 18.710 14.215 18.880 14.445 ;
        RECT 19.265 14.385 19.730 14.715 ;
        RECT 19.900 15.005 20.070 15.845 ;
        RECT 20.250 15.815 20.565 16.315 ;
        RECT 20.795 15.585 21.135 16.145 ;
        RECT 20.240 15.210 21.135 15.585 ;
        RECT 21.305 15.305 21.475 16.315 ;
        RECT 20.945 15.005 21.135 15.210 ;
        RECT 21.645 15.255 21.975 16.100 ;
        RECT 23.160 15.525 23.695 16.145 ;
        RECT 21.645 15.175 22.035 15.255 ;
        RECT 21.820 15.125 22.035 15.175 ;
        RECT 19.900 14.675 20.775 15.005 ;
        RECT 20.945 14.675 21.695 15.005 ;
        RECT 19.900 14.215 20.070 14.675 ;
        RECT 20.945 14.505 21.145 14.675 ;
        RECT 21.865 14.545 22.035 15.125 ;
        RECT 21.810 14.505 22.035 14.545 ;
        RECT 18.710 14.045 19.115 14.215 ;
        RECT 19.285 14.045 20.070 14.215 ;
        RECT 20.345 13.765 20.555 14.295 ;
        RECT 20.815 13.980 21.145 14.505 ;
        RECT 21.655 14.420 22.035 14.505 ;
        RECT 23.160 14.505 23.475 15.525 ;
        RECT 23.865 15.515 24.195 16.315 ;
        RECT 24.680 15.345 25.070 15.520 ;
        RECT 23.645 15.175 25.070 15.345 ;
        RECT 23.645 14.675 23.815 15.175 ;
        RECT 21.315 13.765 21.485 14.375 ;
        RECT 21.655 13.985 21.985 14.420 ;
        RECT 23.160 13.935 23.775 14.505 ;
        RECT 24.065 14.445 24.330 15.005 ;
        RECT 24.500 14.275 24.670 15.175 ;
        RECT 26.345 15.150 26.635 16.315 ;
        RECT 27.730 15.165 27.990 16.315 ;
        RECT 28.165 15.240 28.420 16.145 ;
        RECT 28.590 15.555 28.920 16.315 ;
        RECT 29.135 15.385 29.305 16.145 ;
        RECT 24.840 14.445 25.195 15.005 ;
        RECT 23.945 13.765 24.160 14.275 ;
        RECT 24.390 13.945 24.670 14.275 ;
        RECT 24.850 13.765 25.090 14.275 ;
        RECT 26.345 13.765 26.635 14.490 ;
        RECT 27.730 13.765 27.990 14.605 ;
        RECT 28.165 14.510 28.335 15.240 ;
        RECT 28.590 15.215 29.305 15.385 ;
        RECT 28.590 15.005 28.760 15.215 ;
        RECT 30.030 15.165 30.290 16.315 ;
        RECT 30.465 15.240 30.720 16.145 ;
        RECT 30.890 15.555 31.220 16.315 ;
        RECT 31.435 15.385 31.605 16.145 ;
        RECT 28.505 14.675 28.760 15.005 ;
        RECT 28.165 13.935 28.420 14.510 ;
        RECT 28.590 14.485 28.760 14.675 ;
        RECT 29.040 14.665 29.395 15.035 ;
        RECT 28.590 14.315 29.305 14.485 ;
        RECT 28.590 13.765 28.920 14.145 ;
        RECT 29.135 13.935 29.305 14.315 ;
        RECT 30.030 13.765 30.290 14.605 ;
        RECT 30.465 14.510 30.635 15.240 ;
        RECT 30.890 15.215 31.605 15.385 ;
        RECT 30.890 15.005 31.060 15.215 ;
        RECT 31.870 15.165 32.130 16.315 ;
        RECT 32.305 15.240 32.560 16.145 ;
        RECT 32.730 15.555 33.060 16.315 ;
        RECT 33.275 15.385 33.445 16.145 ;
        RECT 30.805 14.675 31.060 15.005 ;
        RECT 30.465 13.935 30.720 14.510 ;
        RECT 30.890 14.485 31.060 14.675 ;
        RECT 31.340 14.665 31.695 15.035 ;
        RECT 30.890 14.315 31.605 14.485 ;
        RECT 30.890 13.765 31.220 14.145 ;
        RECT 31.435 13.935 31.605 14.315 ;
        RECT 31.870 13.765 32.130 14.605 ;
        RECT 32.305 14.510 32.475 15.240 ;
        RECT 32.730 15.215 33.445 15.385 ;
        RECT 32.730 15.005 32.900 15.215 ;
        RECT 33.710 15.165 33.970 16.315 ;
        RECT 34.145 15.240 34.400 16.145 ;
        RECT 34.570 15.555 34.900 16.315 ;
        RECT 35.115 15.385 35.285 16.145 ;
        RECT 32.645 14.675 32.900 15.005 ;
        RECT 32.305 13.935 32.560 14.510 ;
        RECT 32.730 14.485 32.900 14.675 ;
        RECT 33.180 14.665 33.535 15.035 ;
        RECT 32.730 14.315 33.445 14.485 ;
        RECT 32.730 13.765 33.060 14.145 ;
        RECT 33.275 13.935 33.445 14.315 ;
        RECT 33.710 13.765 33.970 14.605 ;
        RECT 34.145 14.510 34.315 15.240 ;
        RECT 34.570 15.215 35.285 15.385 ;
        RECT 34.570 15.005 34.740 15.215 ;
        RECT 35.550 15.165 35.810 16.315 ;
        RECT 35.985 15.240 36.240 16.145 ;
        RECT 36.410 15.555 36.740 16.315 ;
        RECT 36.955 15.385 37.125 16.145 ;
        RECT 34.485 14.675 34.740 15.005 ;
        RECT 34.145 13.935 34.400 14.510 ;
        RECT 34.570 14.485 34.740 14.675 ;
        RECT 35.020 14.665 35.375 15.035 ;
        RECT 34.570 14.315 35.285 14.485 ;
        RECT 34.570 13.765 34.900 14.145 ;
        RECT 35.115 13.935 35.285 14.315 ;
        RECT 35.550 13.765 35.810 14.605 ;
        RECT 35.985 14.510 36.155 15.240 ;
        RECT 36.410 15.215 37.125 15.385 ;
        RECT 36.410 15.005 36.580 15.215 ;
        RECT 37.390 15.165 37.650 16.315 ;
        RECT 37.825 15.240 38.080 16.145 ;
        RECT 38.250 15.555 38.580 16.315 ;
        RECT 38.795 15.385 38.965 16.145 ;
        RECT 36.325 14.675 36.580 15.005 ;
        RECT 35.985 13.935 36.240 14.510 ;
        RECT 36.410 14.485 36.580 14.675 ;
        RECT 36.860 14.665 37.215 15.035 ;
        RECT 36.410 14.315 37.125 14.485 ;
        RECT 36.410 13.765 36.740 14.145 ;
        RECT 36.955 13.935 37.125 14.315 ;
        RECT 37.390 13.765 37.650 14.605 ;
        RECT 37.825 14.510 37.995 15.240 ;
        RECT 38.250 15.215 38.965 15.385 ;
        RECT 38.250 15.005 38.420 15.215 ;
        RECT 39.225 15.150 39.515 16.315 ;
        RECT 40.610 15.925 40.945 16.145 ;
        RECT 41.950 15.935 42.305 16.315 ;
        RECT 40.610 15.305 40.865 15.925 ;
        RECT 41.115 15.765 41.345 15.805 ;
        RECT 42.475 15.765 42.725 16.145 ;
        RECT 41.115 15.565 42.725 15.765 ;
        RECT 41.115 15.475 41.300 15.565 ;
        RECT 41.890 15.555 42.725 15.565 ;
        RECT 42.975 15.535 43.225 16.315 ;
        RECT 43.395 15.465 43.655 16.145 ;
        RECT 41.455 15.365 41.785 15.395 ;
        RECT 41.455 15.305 43.255 15.365 ;
        RECT 40.610 15.195 43.315 15.305 ;
        RECT 40.610 15.135 41.785 15.195 ;
        RECT 43.115 15.160 43.315 15.195 ;
        RECT 38.165 14.675 38.420 15.005 ;
        RECT 37.825 13.935 38.080 14.510 ;
        RECT 38.250 14.485 38.420 14.675 ;
        RECT 38.700 14.665 39.055 15.035 ;
        RECT 40.605 14.755 41.095 14.955 ;
        RECT 41.285 14.755 41.760 14.965 ;
        RECT 38.250 14.315 38.965 14.485 ;
        RECT 38.250 13.765 38.580 14.145 ;
        RECT 38.795 13.935 38.965 14.315 ;
        RECT 39.225 13.765 39.515 14.490 ;
        RECT 40.610 13.765 41.065 14.530 ;
        RECT 41.540 14.355 41.760 14.755 ;
        RECT 42.005 14.755 42.335 14.965 ;
        RECT 42.005 14.355 42.215 14.755 ;
        RECT 42.505 14.720 42.915 15.025 ;
        RECT 43.145 14.585 43.315 15.160 ;
        RECT 43.045 14.465 43.315 14.585 ;
        RECT 42.470 14.420 43.315 14.465 ;
        RECT 42.470 14.295 43.225 14.420 ;
        RECT 42.470 14.145 42.640 14.295 ;
        RECT 43.485 14.265 43.655 15.465 ;
        RECT 44.010 15.345 44.400 15.520 ;
        RECT 44.885 15.515 45.215 16.315 ;
        RECT 45.385 15.525 45.920 16.145 ;
        RECT 44.010 15.175 45.435 15.345 ;
        RECT 43.885 14.445 44.240 15.005 ;
        RECT 44.410 14.275 44.580 15.175 ;
        RECT 44.750 14.445 45.015 15.005 ;
        RECT 45.265 14.675 45.435 15.175 ;
        RECT 45.605 14.505 45.920 15.525 ;
        RECT 46.130 15.165 46.390 16.315 ;
        RECT 46.565 15.240 46.820 16.145 ;
        RECT 46.990 15.555 47.320 16.315 ;
        RECT 47.535 15.385 47.705 16.145 ;
        RECT 41.340 13.935 42.640 14.145 ;
        RECT 42.895 13.765 43.225 14.125 ;
        RECT 43.395 13.935 43.655 14.265 ;
        RECT 43.990 13.765 44.230 14.275 ;
        RECT 44.410 13.945 44.690 14.275 ;
        RECT 44.920 13.765 45.135 14.275 ;
        RECT 45.305 13.935 45.920 14.505 ;
        RECT 46.130 13.765 46.390 14.605 ;
        RECT 46.565 14.510 46.735 15.240 ;
        RECT 46.990 15.215 47.705 15.385 ;
        RECT 48.055 15.385 48.225 16.145 ;
        RECT 48.440 15.555 48.770 16.315 ;
        RECT 48.055 15.215 48.770 15.385 ;
        RECT 48.940 15.240 49.195 16.145 ;
        RECT 46.990 15.005 47.160 15.215 ;
        RECT 46.905 14.675 47.160 15.005 ;
        RECT 46.565 13.935 46.820 14.510 ;
        RECT 46.990 14.485 47.160 14.675 ;
        RECT 47.440 14.665 47.795 15.035 ;
        RECT 47.965 14.665 48.320 15.035 ;
        RECT 48.600 15.005 48.770 15.215 ;
        RECT 48.600 14.675 48.855 15.005 ;
        RECT 48.600 14.485 48.770 14.675 ;
        RECT 49.025 14.510 49.195 15.240 ;
        RECT 49.370 15.165 49.630 16.315 ;
        RECT 49.990 15.345 50.380 15.520 ;
        RECT 50.865 15.515 51.195 16.315 ;
        RECT 51.365 15.525 51.900 16.145 ;
        RECT 49.990 15.175 51.415 15.345 ;
        RECT 46.990 14.315 47.705 14.485 ;
        RECT 46.990 13.765 47.320 14.145 ;
        RECT 47.535 13.935 47.705 14.315 ;
        RECT 48.055 14.315 48.770 14.485 ;
        RECT 48.055 13.935 48.225 14.315 ;
        RECT 48.440 13.765 48.770 14.145 ;
        RECT 48.940 13.935 49.195 14.510 ;
        RECT 49.370 13.765 49.630 14.605 ;
        RECT 49.865 14.445 50.220 15.005 ;
        RECT 50.390 14.275 50.560 15.175 ;
        RECT 50.730 14.445 50.995 15.005 ;
        RECT 51.245 14.675 51.415 15.175 ;
        RECT 51.585 14.505 51.900 15.525 ;
        RECT 52.105 15.150 52.395 16.315 ;
        RECT 53.490 15.165 53.750 16.315 ;
        RECT 53.925 15.240 54.180 16.145 ;
        RECT 54.350 15.555 54.680 16.315 ;
        RECT 54.895 15.385 55.065 16.145 ;
        RECT 49.970 13.765 50.210 14.275 ;
        RECT 50.390 13.945 50.670 14.275 ;
        RECT 50.900 13.765 51.115 14.275 ;
        RECT 51.285 13.935 51.900 14.505 ;
        RECT 52.105 13.765 52.395 14.490 ;
        RECT 53.490 13.765 53.750 14.605 ;
        RECT 53.925 14.510 54.095 15.240 ;
        RECT 54.350 15.215 55.065 15.385 ;
        RECT 55.325 15.225 56.535 16.315 ;
        RECT 54.350 15.005 54.520 15.215 ;
        RECT 54.265 14.675 54.520 15.005 ;
        RECT 53.925 13.935 54.180 14.510 ;
        RECT 54.350 14.485 54.520 14.675 ;
        RECT 54.800 14.665 55.155 15.035 ;
        RECT 55.325 14.515 55.845 15.055 ;
        RECT 56.015 14.685 56.535 15.225 ;
        RECT 56.710 15.165 56.970 16.315 ;
        RECT 57.145 15.240 57.400 16.145 ;
        RECT 57.570 15.555 57.900 16.315 ;
        RECT 58.115 15.385 58.285 16.145 ;
        RECT 54.350 14.315 55.065 14.485 ;
        RECT 54.350 13.765 54.680 14.145 ;
        RECT 54.895 13.935 55.065 14.315 ;
        RECT 55.325 13.765 56.535 14.515 ;
        RECT 56.710 13.765 56.970 14.605 ;
        RECT 57.145 14.510 57.315 15.240 ;
        RECT 57.570 15.215 58.285 15.385 ;
        RECT 58.545 15.225 59.755 16.315 ;
        RECT 57.570 15.005 57.740 15.215 ;
        RECT 57.485 14.675 57.740 15.005 ;
        RECT 57.145 13.935 57.400 14.510 ;
        RECT 57.570 14.485 57.740 14.675 ;
        RECT 58.020 14.665 58.375 15.035 ;
        RECT 58.545 14.515 59.065 15.055 ;
        RECT 59.235 14.685 59.755 15.225 ;
        RECT 60.015 15.385 60.185 16.145 ;
        RECT 60.400 15.555 60.730 16.315 ;
        RECT 60.015 15.215 60.730 15.385 ;
        RECT 60.900 15.240 61.155 16.145 ;
        RECT 59.925 14.665 60.280 15.035 ;
        RECT 60.560 15.005 60.730 15.215 ;
        RECT 60.560 14.675 60.815 15.005 ;
        RECT 57.570 14.315 58.285 14.485 ;
        RECT 57.570 13.765 57.900 14.145 ;
        RECT 58.115 13.935 58.285 14.315 ;
        RECT 58.545 13.765 59.755 14.515 ;
        RECT 60.560 14.485 60.730 14.675 ;
        RECT 60.985 14.510 61.155 15.240 ;
        RECT 61.330 15.165 61.590 16.315 ;
        RECT 61.765 15.225 62.975 16.315 ;
        RECT 60.015 14.315 60.730 14.485 ;
        RECT 60.015 13.935 60.185 14.315 ;
        RECT 60.400 13.765 60.730 14.145 ;
        RECT 60.900 13.935 61.155 14.510 ;
        RECT 61.330 13.765 61.590 14.605 ;
        RECT 61.765 14.515 62.285 15.055 ;
        RECT 62.455 14.685 62.975 15.225 ;
        RECT 63.150 15.165 63.410 16.315 ;
        RECT 63.585 15.240 63.840 16.145 ;
        RECT 64.010 15.555 64.340 16.315 ;
        RECT 64.555 15.385 64.725 16.145 ;
        RECT 61.765 13.765 62.975 14.515 ;
        RECT 63.150 13.765 63.410 14.605 ;
        RECT 63.585 14.510 63.755 15.240 ;
        RECT 64.010 15.215 64.725 15.385 ;
        RECT 64.010 15.005 64.180 15.215 ;
        RECT 64.985 15.150 65.275 16.315 ;
        RECT 66.370 15.165 66.630 16.315 ;
        RECT 66.805 15.240 67.060 16.145 ;
        RECT 67.230 15.555 67.560 16.315 ;
        RECT 67.775 15.385 67.945 16.145 ;
        RECT 63.925 14.675 64.180 15.005 ;
        RECT 63.585 13.935 63.840 14.510 ;
        RECT 64.010 14.485 64.180 14.675 ;
        RECT 64.460 14.665 64.815 15.035 ;
        RECT 64.010 14.315 64.725 14.485 ;
        RECT 64.010 13.765 64.340 14.145 ;
        RECT 64.555 13.935 64.725 14.315 ;
        RECT 64.985 13.765 65.275 14.490 ;
        RECT 66.370 13.765 66.630 14.605 ;
        RECT 66.805 14.510 66.975 15.240 ;
        RECT 67.230 15.215 67.945 15.385 ;
        RECT 68.205 15.225 69.415 16.315 ;
        RECT 67.230 15.005 67.400 15.215 ;
        RECT 67.145 14.675 67.400 15.005 ;
        RECT 66.805 13.935 67.060 14.510 ;
        RECT 67.230 14.485 67.400 14.675 ;
        RECT 67.680 14.665 68.035 15.035 ;
        RECT 68.205 14.515 68.725 15.055 ;
        RECT 68.895 14.685 69.415 15.225 ;
        RECT 69.590 15.165 69.850 16.315 ;
        RECT 70.025 15.240 70.280 16.145 ;
        RECT 70.450 15.555 70.780 16.315 ;
        RECT 70.995 15.385 71.165 16.145 ;
        RECT 67.230 14.315 67.945 14.485 ;
        RECT 67.230 13.765 67.560 14.145 ;
        RECT 67.775 13.935 67.945 14.315 ;
        RECT 68.205 13.765 69.415 14.515 ;
        RECT 69.590 13.765 69.850 14.605 ;
        RECT 70.025 14.510 70.195 15.240 ;
        RECT 70.450 15.215 71.165 15.385 ;
        RECT 71.425 15.225 72.635 16.315 ;
        RECT 70.450 15.005 70.620 15.215 ;
        RECT 70.365 14.675 70.620 15.005 ;
        RECT 70.025 13.935 70.280 14.510 ;
        RECT 70.450 14.485 70.620 14.675 ;
        RECT 70.900 14.665 71.255 15.035 ;
        RECT 71.425 14.515 71.945 15.055 ;
        RECT 72.115 14.685 72.635 15.225 ;
        RECT 72.895 15.385 73.065 16.145 ;
        RECT 73.280 15.555 73.610 16.315 ;
        RECT 72.895 15.215 73.610 15.385 ;
        RECT 73.780 15.240 74.035 16.145 ;
        RECT 72.805 14.665 73.160 15.035 ;
        RECT 73.440 15.005 73.610 15.215 ;
        RECT 73.440 14.675 73.695 15.005 ;
        RECT 70.450 14.315 71.165 14.485 ;
        RECT 70.450 13.765 70.780 14.145 ;
        RECT 70.995 13.935 71.165 14.315 ;
        RECT 71.425 13.765 72.635 14.515 ;
        RECT 73.440 14.485 73.610 14.675 ;
        RECT 73.865 14.510 74.035 15.240 ;
        RECT 74.210 15.165 74.470 16.315 ;
        RECT 74.645 15.225 75.855 16.315 ;
        RECT 72.895 14.315 73.610 14.485 ;
        RECT 72.895 13.935 73.065 14.315 ;
        RECT 73.280 13.765 73.610 14.145 ;
        RECT 73.780 13.935 74.035 14.510 ;
        RECT 74.210 13.765 74.470 14.605 ;
        RECT 74.645 14.515 75.165 15.055 ;
        RECT 75.335 14.685 75.855 15.225 ;
        RECT 76.030 15.165 76.290 16.315 ;
        RECT 76.465 15.240 76.720 16.145 ;
        RECT 76.890 15.555 77.220 16.315 ;
        RECT 77.435 15.385 77.605 16.145 ;
        RECT 74.645 13.765 75.855 14.515 ;
        RECT 76.030 13.765 76.290 14.605 ;
        RECT 76.465 14.510 76.635 15.240 ;
        RECT 76.890 15.215 77.605 15.385 ;
        RECT 76.890 15.005 77.060 15.215 ;
        RECT 77.865 15.150 78.155 16.315 ;
        RECT 78.510 15.345 78.900 15.520 ;
        RECT 79.385 15.515 79.715 16.315 ;
        RECT 79.885 15.525 80.420 16.145 ;
        RECT 78.510 15.175 79.935 15.345 ;
        RECT 76.805 14.675 77.060 15.005 ;
        RECT 76.465 13.935 76.720 14.510 ;
        RECT 76.890 14.485 77.060 14.675 ;
        RECT 77.340 14.665 77.695 15.035 ;
        RECT 76.890 14.315 77.605 14.485 ;
        RECT 76.890 13.765 77.220 14.145 ;
        RECT 77.435 13.935 77.605 14.315 ;
        RECT 77.865 13.765 78.155 14.490 ;
        RECT 78.385 14.445 78.740 15.005 ;
        RECT 78.910 14.275 79.080 15.175 ;
        RECT 79.250 14.445 79.515 15.005 ;
        RECT 79.765 14.675 79.935 15.175 ;
        RECT 80.105 14.505 80.420 15.525 ;
        RECT 80.810 15.345 81.200 15.520 ;
        RECT 81.685 15.515 82.015 16.315 ;
        RECT 82.185 15.525 82.720 16.145 ;
        RECT 80.810 15.175 82.235 15.345 ;
        RECT 78.490 13.765 78.730 14.275 ;
        RECT 78.910 13.945 79.190 14.275 ;
        RECT 79.420 13.765 79.635 14.275 ;
        RECT 79.805 13.935 80.420 14.505 ;
        RECT 80.685 14.445 81.040 15.005 ;
        RECT 81.210 14.275 81.380 15.175 ;
        RECT 81.550 14.445 81.815 15.005 ;
        RECT 82.065 14.675 82.235 15.175 ;
        RECT 82.405 14.505 82.720 15.525 ;
        RECT 83.475 15.645 83.645 16.145 ;
        RECT 83.815 15.815 84.145 16.315 ;
        RECT 83.475 15.475 84.140 15.645 ;
        RECT 83.390 14.655 83.740 15.305 ;
        RECT 80.790 13.765 81.030 14.275 ;
        RECT 81.210 13.945 81.490 14.275 ;
        RECT 81.720 13.765 81.935 14.275 ;
        RECT 82.105 13.935 82.720 14.505 ;
        RECT 83.910 14.485 84.140 15.475 ;
        RECT 83.475 14.315 84.140 14.485 ;
        RECT 83.475 14.025 83.645 14.315 ;
        RECT 83.815 13.765 84.145 14.145 ;
        RECT 84.315 14.025 84.500 16.145 ;
        RECT 84.740 15.855 85.005 16.315 ;
        RECT 85.175 15.720 85.425 16.145 ;
        RECT 85.635 15.870 86.740 16.040 ;
        RECT 85.120 15.590 85.425 15.720 ;
        RECT 84.670 14.395 84.950 15.345 ;
        RECT 85.120 14.485 85.290 15.590 ;
        RECT 85.460 14.805 85.700 15.400 ;
        RECT 85.870 15.335 86.400 15.700 ;
        RECT 85.870 14.635 86.040 15.335 ;
        RECT 86.570 15.255 86.740 15.870 ;
        RECT 86.910 15.515 87.080 16.315 ;
        RECT 87.250 15.815 87.500 16.145 ;
        RECT 87.725 15.845 88.610 16.015 ;
        RECT 86.570 15.165 87.080 15.255 ;
        RECT 85.120 14.355 85.345 14.485 ;
        RECT 85.515 14.415 86.040 14.635 ;
        RECT 86.210 14.995 87.080 15.165 ;
        RECT 84.755 13.765 85.005 14.225 ;
        RECT 85.175 14.215 85.345 14.355 ;
        RECT 86.210 14.215 86.380 14.995 ;
        RECT 86.910 14.925 87.080 14.995 ;
        RECT 86.590 14.745 86.790 14.775 ;
        RECT 87.250 14.745 87.420 15.815 ;
        RECT 87.590 14.925 87.780 15.645 ;
        RECT 86.590 14.445 87.420 14.745 ;
        RECT 87.950 14.715 88.270 15.675 ;
        RECT 85.175 14.045 85.510 14.215 ;
        RECT 85.705 14.045 86.380 14.215 ;
        RECT 86.700 13.765 87.070 14.265 ;
        RECT 87.250 14.215 87.420 14.445 ;
        RECT 87.805 14.385 88.270 14.715 ;
        RECT 88.440 15.005 88.610 15.845 ;
        RECT 88.790 15.815 89.105 16.315 ;
        RECT 89.335 15.585 89.675 16.145 ;
        RECT 88.780 15.210 89.675 15.585 ;
        RECT 89.845 15.305 90.015 16.315 ;
        RECT 89.485 15.005 89.675 15.210 ;
        RECT 90.185 15.255 90.515 16.100 ;
        RECT 90.185 15.175 90.575 15.255 ;
        RECT 90.360 15.125 90.575 15.175 ;
        RECT 88.440 14.675 89.315 15.005 ;
        RECT 89.485 14.675 90.235 15.005 ;
        RECT 88.440 14.215 88.610 14.675 ;
        RECT 89.485 14.505 89.685 14.675 ;
        RECT 90.405 14.545 90.575 15.125 ;
        RECT 90.745 15.225 91.955 16.315 ;
        RECT 90.745 14.685 91.265 15.225 ;
        RECT 90.350 14.505 90.575 14.545 ;
        RECT 91.435 14.515 91.955 15.055 ;
        RECT 87.250 14.045 87.655 14.215 ;
        RECT 87.825 14.045 88.610 14.215 ;
        RECT 88.885 13.765 89.095 14.295 ;
        RECT 89.355 13.980 89.685 14.505 ;
        RECT 90.195 14.420 90.575 14.505 ;
        RECT 89.855 13.765 90.025 14.375 ;
        RECT 90.195 13.985 90.525 14.420 ;
        RECT 90.745 13.765 91.955 14.515 ;
        RECT 13.380 13.595 92.040 13.765 ;
      LAYER met1 ;
        RECT 149.710 221.830 149.970 222.150 ;
        RECT 149.150 220.770 149.410 221.090 ;
        RECT 115.800 220.285 116.060 220.605 ;
        RECT 110.950 206.310 111.210 206.630 ;
        RECT 109.950 205.860 110.210 206.180 ;
        RECT 13.380 201.120 92.040 201.600 ;
        RECT 51.170 200.920 51.490 200.980 ;
        RECT 59.005 200.920 59.295 200.965 ;
        RECT 51.170 200.780 59.295 200.920 ;
        RECT 51.170 200.720 51.490 200.780 ;
        RECT 59.005 200.735 59.295 200.780 ;
        RECT 62.670 199.900 62.990 199.960 ;
        RECT 63.145 199.900 63.435 199.945 ;
        RECT 62.670 199.760 63.435 199.900 ;
        RECT 62.670 199.700 62.990 199.760 ;
        RECT 63.145 199.715 63.435 199.760 ;
        RECT 72.330 199.900 72.650 199.960 ;
        RECT 73.725 199.900 74.015 199.945 ;
        RECT 72.330 199.760 74.015 199.900 ;
        RECT 72.330 199.700 72.650 199.760 ;
        RECT 73.725 199.715 74.015 199.760 ;
        RECT 48.870 199.560 49.190 199.620 ;
        RECT 59.925 199.560 60.215 199.605 ;
        RECT 48.870 199.420 60.215 199.560 ;
        RECT 48.870 199.360 49.190 199.420 ;
        RECT 59.925 199.375 60.215 199.420 ;
        RECT 58.070 199.020 58.390 199.280 ;
        RECT 58.925 199.220 59.215 199.265 ;
        RECT 61.750 199.220 62.070 199.280 ;
        RECT 58.925 199.080 62.070 199.220 ;
        RECT 58.925 199.035 59.215 199.080 ;
        RECT 61.750 199.020 62.070 199.080 ;
        RECT 64.065 199.220 64.355 199.265 ;
        RECT 64.510 199.220 64.830 199.280 ;
        RECT 64.065 199.080 64.830 199.220 ;
        RECT 64.065 199.035 64.355 199.080 ;
        RECT 64.510 199.020 64.830 199.080 ;
        RECT 70.950 199.220 71.270 199.280 ;
        RECT 72.805 199.220 73.095 199.265 ;
        RECT 70.950 199.080 73.095 199.220 ;
        RECT 70.950 199.020 71.270 199.080 ;
        RECT 72.805 199.035 73.095 199.080 ;
        RECT 13.380 198.400 92.040 198.880 ;
        RECT 45.665 198.015 45.955 198.245 ;
        RECT 58.070 198.200 58.390 198.260 ;
        RECT 58.070 198.060 58.760 198.200 ;
        RECT 42.890 197.860 43.210 197.920 ;
        RECT 44.730 197.905 45.050 197.920 ;
        RECT 43.825 197.860 44.115 197.905 ;
        RECT 42.890 197.720 44.115 197.860 ;
        RECT 42.890 197.660 43.210 197.720 ;
        RECT 43.825 197.675 44.115 197.720 ;
        RECT 44.730 197.675 45.115 197.905 ;
        RECT 45.740 197.860 45.880 198.015 ;
        RECT 58.070 198.000 58.390 198.060 ;
        RECT 58.620 197.905 58.760 198.060 ;
        RECT 47.350 197.860 47.640 197.905 ;
        RECT 45.740 197.720 47.640 197.860 ;
        RECT 47.350 197.675 47.640 197.720 ;
        RECT 58.500 197.675 58.790 197.905 ;
        RECT 42.430 197.320 42.750 197.580 ;
        RECT 43.350 197.320 43.670 197.580 ;
        RECT 43.900 197.520 44.040 197.675 ;
        RECT 44.730 197.660 45.050 197.675 ;
        RECT 48.870 197.520 49.190 197.580 ;
        RECT 43.900 197.380 49.190 197.520 ;
        RECT 48.870 197.320 49.190 197.380 ;
        RECT 71.410 197.520 71.730 197.580 ;
        RECT 73.310 197.520 73.600 197.565 ;
        RECT 71.410 197.380 73.600 197.520 ;
        RECT 71.410 197.320 71.730 197.380 ;
        RECT 73.310 197.335 73.600 197.380 ;
        RECT 38.290 197.180 38.610 197.240 ;
        RECT 46.125 197.180 46.415 197.225 ;
        RECT 38.290 197.040 46.415 197.180 ;
        RECT 38.290 196.980 38.610 197.040 ;
        RECT 46.125 196.995 46.415 197.040 ;
        RECT 47.005 197.180 47.295 197.225 ;
        RECT 48.195 197.180 48.485 197.225 ;
        RECT 50.715 197.180 51.005 197.225 ;
        RECT 47.005 197.040 51.005 197.180 ;
        RECT 47.005 196.995 47.295 197.040 ;
        RECT 48.195 196.995 48.485 197.040 ;
        RECT 50.715 196.995 51.005 197.040 ;
        RECT 56.690 197.180 57.010 197.240 ;
        RECT 57.165 197.180 57.455 197.225 ;
        RECT 56.690 197.040 57.455 197.180 ;
        RECT 56.690 196.980 57.010 197.040 ;
        RECT 57.165 196.995 57.455 197.040 ;
        RECT 58.045 197.180 58.335 197.225 ;
        RECT 59.235 197.180 59.525 197.225 ;
        RECT 61.755 197.180 62.045 197.225 ;
        RECT 58.045 197.040 62.045 197.180 ;
        RECT 58.045 196.995 58.335 197.040 ;
        RECT 59.235 196.995 59.525 197.040 ;
        RECT 61.755 196.995 62.045 197.040 ;
        RECT 70.055 197.180 70.345 197.225 ;
        RECT 72.575 197.180 72.865 197.225 ;
        RECT 73.765 197.180 74.055 197.225 ;
        RECT 70.055 197.040 74.055 197.180 ;
        RECT 70.055 196.995 70.345 197.040 ;
        RECT 72.575 196.995 72.865 197.040 ;
        RECT 73.765 196.995 74.055 197.040 ;
        RECT 74.645 197.180 74.935 197.225 ;
        RECT 77.390 197.180 77.710 197.240 ;
        RECT 74.645 197.040 77.710 197.180 ;
        RECT 74.645 196.995 74.935 197.040 ;
        RECT 77.390 196.980 77.710 197.040 ;
        RECT 46.610 196.840 46.900 196.885 ;
        RECT 48.710 196.840 49.000 196.885 ;
        RECT 50.280 196.840 50.570 196.885 ;
        RECT 46.610 196.700 50.570 196.840 ;
        RECT 46.610 196.655 46.900 196.700 ;
        RECT 48.710 196.655 49.000 196.700 ;
        RECT 50.280 196.655 50.570 196.700 ;
        RECT 57.650 196.840 57.940 196.885 ;
        RECT 59.750 196.840 60.040 196.885 ;
        RECT 61.320 196.840 61.610 196.885 ;
        RECT 57.650 196.700 61.610 196.840 ;
        RECT 57.650 196.655 57.940 196.700 ;
        RECT 59.750 196.655 60.040 196.700 ;
        RECT 61.320 196.655 61.610 196.700 ;
        RECT 70.490 196.840 70.780 196.885 ;
        RECT 72.060 196.840 72.350 196.885 ;
        RECT 74.160 196.840 74.450 196.885 ;
        RECT 70.490 196.700 74.450 196.840 ;
        RECT 70.490 196.655 70.780 196.700 ;
        RECT 72.060 196.655 72.350 196.700 ;
        RECT 74.160 196.655 74.450 196.700 ;
        RECT 43.350 196.300 43.670 196.560 ;
        RECT 44.745 196.500 45.035 196.545 ;
        RECT 47.490 196.500 47.810 196.560 ;
        RECT 44.745 196.360 47.810 196.500 ;
        RECT 44.745 196.315 45.035 196.360 ;
        RECT 47.490 196.300 47.810 196.360 ;
        RECT 49.330 196.500 49.650 196.560 ;
        RECT 53.025 196.500 53.315 196.545 ;
        RECT 49.330 196.360 53.315 196.500 ;
        RECT 49.330 196.300 49.650 196.360 ;
        RECT 53.025 196.315 53.315 196.360 ;
        RECT 63.130 196.500 63.450 196.560 ;
        RECT 64.065 196.500 64.355 196.545 ;
        RECT 63.130 196.360 64.355 196.500 ;
        RECT 63.130 196.300 63.450 196.360 ;
        RECT 64.065 196.315 64.355 196.360 ;
        RECT 67.745 196.500 68.035 196.545 ;
        RECT 68.190 196.500 68.510 196.560 ;
        RECT 67.745 196.360 68.510 196.500 ;
        RECT 67.745 196.315 68.035 196.360 ;
        RECT 68.190 196.300 68.510 196.360 ;
        RECT 13.380 195.680 92.040 196.160 ;
        RECT 46.570 195.480 46.890 195.540 ;
        RECT 47.045 195.480 47.335 195.525 ;
        RECT 46.570 195.340 47.335 195.480 ;
        RECT 46.570 195.280 46.890 195.340 ;
        RECT 47.045 195.295 47.335 195.340 ;
        RECT 47.490 195.480 47.810 195.540 ;
        RECT 50.725 195.480 51.015 195.525 ;
        RECT 51.170 195.480 51.490 195.540 ;
        RECT 47.490 195.340 51.490 195.480 ;
        RECT 47.490 195.280 47.810 195.340 ;
        RECT 50.725 195.295 51.015 195.340 ;
        RECT 51.170 195.280 51.490 195.340 ;
        RECT 61.750 195.280 62.070 195.540 ;
        RECT 68.205 195.480 68.495 195.525 ;
        RECT 68.650 195.480 68.970 195.540 ;
        RECT 68.205 195.340 68.970 195.480 ;
        RECT 68.205 195.295 68.495 195.340 ;
        RECT 68.650 195.280 68.970 195.340 ;
        RECT 69.125 195.480 69.415 195.525 ;
        RECT 71.410 195.480 71.730 195.540 ;
        RECT 69.125 195.340 71.730 195.480 ;
        RECT 69.125 195.295 69.415 195.340 ;
        RECT 71.410 195.280 71.730 195.340 ;
        RECT 38.790 195.140 39.080 195.185 ;
        RECT 40.890 195.140 41.180 195.185 ;
        RECT 42.460 195.140 42.750 195.185 ;
        RECT 38.790 195.000 42.750 195.140 ;
        RECT 38.790 194.955 39.080 195.000 ;
        RECT 40.890 194.955 41.180 195.000 ;
        RECT 42.460 194.955 42.750 195.000 ;
        RECT 44.730 195.140 45.050 195.200 ;
        RECT 48.425 195.140 48.715 195.185 ;
        RECT 44.730 195.000 48.715 195.140 ;
        RECT 44.730 194.940 45.050 195.000 ;
        RECT 48.425 194.955 48.715 195.000 ;
        RECT 53.050 195.140 53.340 195.185 ;
        RECT 55.150 195.140 55.440 195.185 ;
        RECT 56.720 195.140 57.010 195.185 ;
        RECT 53.050 195.000 57.010 195.140 ;
        RECT 53.050 194.955 53.340 195.000 ;
        RECT 55.150 194.955 55.440 195.000 ;
        RECT 56.720 194.955 57.010 195.000 ;
        RECT 73.250 195.140 73.540 195.185 ;
        RECT 74.820 195.140 75.110 195.185 ;
        RECT 76.920 195.140 77.210 195.185 ;
        RECT 73.250 195.000 77.210 195.140 ;
        RECT 73.250 194.955 73.540 195.000 ;
        RECT 74.820 194.955 75.110 195.000 ;
        RECT 76.920 194.955 77.210 195.000 ;
        RECT 38.290 194.600 38.610 194.860 ;
        RECT 39.185 194.800 39.475 194.845 ;
        RECT 40.375 194.800 40.665 194.845 ;
        RECT 42.895 194.800 43.185 194.845 ;
        RECT 53.445 194.800 53.735 194.845 ;
        RECT 54.635 194.800 54.925 194.845 ;
        RECT 57.155 194.800 57.445 194.845 ;
        RECT 63.605 194.800 63.895 194.845 ;
        RECT 39.185 194.660 43.185 194.800 ;
        RECT 39.185 194.615 39.475 194.660 ;
        RECT 40.375 194.615 40.665 194.660 ;
        RECT 42.895 194.615 43.185 194.660 ;
        RECT 46.200 194.660 49.560 194.800 ;
        RECT 39.640 194.120 39.930 194.165 ;
        RECT 41.050 194.120 41.370 194.180 ;
        RECT 39.640 193.980 41.370 194.120 ;
        RECT 39.640 193.935 39.930 193.980 ;
        RECT 41.050 193.920 41.370 193.980 ;
        RECT 46.200 193.840 46.340 194.660 ;
        RECT 48.410 194.260 48.730 194.520 ;
        RECT 49.420 194.505 49.560 194.660 ;
        RECT 53.445 194.660 57.445 194.800 ;
        RECT 53.445 194.615 53.735 194.660 ;
        RECT 54.635 194.615 54.925 194.660 ;
        RECT 57.155 194.615 57.445 194.660 ;
        RECT 61.840 194.660 63.895 194.800 ;
        RECT 49.345 194.275 49.635 194.505 ;
        RECT 50.250 194.460 50.570 194.520 ;
        RECT 52.565 194.460 52.855 194.505 ;
        RECT 56.690 194.460 57.010 194.520 ;
        RECT 50.250 194.320 57.010 194.460 ;
        RECT 50.250 194.260 50.570 194.320 ;
        RECT 52.565 194.275 52.855 194.320 ;
        RECT 56.690 194.260 57.010 194.320 ;
        RECT 60.830 194.260 61.150 194.520 ;
        RECT 61.840 194.505 61.980 194.660 ;
        RECT 63.605 194.615 63.895 194.660 ;
        RECT 72.815 194.800 73.105 194.845 ;
        RECT 75.335 194.800 75.625 194.845 ;
        RECT 76.525 194.800 76.815 194.845 ;
        RECT 72.815 194.660 76.815 194.800 ;
        RECT 72.815 194.615 73.105 194.660 ;
        RECT 75.335 194.615 75.625 194.660 ;
        RECT 76.525 194.615 76.815 194.660 ;
        RECT 77.390 194.600 77.710 194.860 ;
        RECT 61.765 194.275 62.055 194.505 ;
        RECT 63.130 194.260 63.450 194.520 ;
        RECT 64.065 194.460 64.355 194.505 ;
        RECT 65.430 194.460 65.750 194.520 ;
        RECT 65.905 194.460 66.195 194.505 ;
        RECT 64.065 194.320 66.195 194.460 ;
        RECT 64.065 194.275 64.355 194.320 ;
        RECT 65.430 194.260 65.750 194.320 ;
        RECT 65.905 194.275 66.195 194.320 ;
        RECT 66.825 194.460 67.115 194.505 ;
        RECT 68.650 194.460 68.970 194.520 ;
        RECT 66.825 194.320 68.970 194.460 ;
        RECT 66.825 194.275 67.115 194.320 ;
        RECT 68.650 194.260 68.970 194.320 ;
        RECT 47.965 193.935 48.255 194.165 ;
        RECT 48.870 194.120 49.190 194.180 ;
        RECT 49.805 194.120 50.095 194.165 ;
        RECT 53.790 194.120 54.080 194.165 ;
        RECT 48.870 193.980 50.095 194.120 ;
        RECT 45.205 193.780 45.495 193.825 ;
        RECT 45.650 193.780 45.970 193.840 ;
        RECT 45.205 193.640 45.970 193.780 ;
        RECT 45.205 193.595 45.495 193.640 ;
        RECT 45.650 193.580 45.970 193.640 ;
        RECT 46.110 193.580 46.430 193.840 ;
        RECT 47.030 193.825 47.350 193.840 ;
        RECT 46.965 193.595 47.350 193.825 ;
        RECT 48.040 193.780 48.180 193.935 ;
        RECT 48.870 193.920 49.190 193.980 ;
        RECT 49.805 193.935 50.095 193.980 ;
        RECT 51.720 193.980 54.080 194.120 ;
        RECT 49.330 193.780 49.650 193.840 ;
        RECT 48.040 193.640 49.650 193.780 ;
        RECT 47.030 193.580 47.350 193.595 ;
        RECT 49.330 193.580 49.650 193.640 ;
        RECT 50.710 193.825 51.030 193.840 ;
        RECT 51.720 193.825 51.860 193.980 ;
        RECT 53.790 193.935 54.080 193.980 ;
        RECT 67.270 193.920 67.590 194.180 ;
        RECT 73.250 194.120 73.570 194.180 ;
        RECT 76.070 194.120 76.360 194.165 ;
        RECT 73.250 193.980 76.360 194.120 ;
        RECT 73.250 193.920 73.570 193.980 ;
        RECT 76.070 193.935 76.360 193.980 ;
        RECT 50.710 193.595 51.095 193.825 ;
        RECT 51.645 193.595 51.935 193.825 ;
        RECT 50.710 193.580 51.030 193.595 ;
        RECT 59.450 193.580 59.770 193.840 ;
        RECT 66.365 193.780 66.655 193.825 ;
        RECT 68.285 193.780 68.575 193.825 ;
        RECT 66.365 193.640 68.575 193.780 ;
        RECT 66.365 193.595 66.655 193.640 ;
        RECT 68.285 193.595 68.575 193.640 ;
        RECT 69.570 193.780 69.890 193.840 ;
        RECT 70.505 193.780 70.795 193.825 ;
        RECT 69.570 193.640 70.795 193.780 ;
        RECT 69.570 193.580 69.890 193.640 ;
        RECT 70.505 193.595 70.795 193.640 ;
        RECT 13.380 192.960 92.040 193.440 ;
        RECT 41.050 192.560 41.370 192.820 ;
        RECT 41.905 192.760 42.195 192.805 ;
        RECT 43.350 192.760 43.670 192.820 ;
        RECT 41.905 192.620 43.670 192.760 ;
        RECT 41.905 192.575 42.195 192.620 ;
        RECT 43.350 192.560 43.670 192.620 ;
        RECT 43.810 192.560 44.130 192.820 ;
        RECT 46.110 192.560 46.430 192.820 ;
        RECT 48.410 192.805 48.730 192.820 ;
        RECT 48.410 192.760 48.745 192.805 ;
        RECT 48.245 192.620 48.745 192.760 ;
        RECT 48.410 192.575 48.745 192.620 ;
        RECT 48.885 192.760 49.175 192.805 ;
        RECT 51.630 192.760 51.950 192.820 ;
        RECT 57.610 192.760 57.930 192.820 ;
        RECT 59.450 192.760 59.770 192.820 ;
        RECT 48.885 192.620 59.770 192.760 ;
        RECT 48.885 192.575 49.175 192.620 ;
        RECT 48.410 192.560 48.730 192.575 ;
        RECT 51.630 192.560 51.950 192.620 ;
        RECT 57.610 192.560 57.930 192.620 ;
        RECT 59.450 192.560 59.770 192.620 ;
        RECT 60.830 192.760 61.150 192.820 ;
        RECT 68.205 192.760 68.495 192.805 ;
        RECT 60.830 192.620 68.495 192.760 ;
        RECT 60.830 192.560 61.150 192.620 ;
        RECT 68.205 192.575 68.495 192.620 ;
        RECT 69.110 192.760 69.430 192.820 ;
        RECT 71.425 192.760 71.715 192.805 ;
        RECT 69.110 192.620 71.715 192.760 ;
        RECT 69.110 192.560 69.430 192.620 ;
        RECT 71.425 192.575 71.715 192.620 ;
        RECT 73.250 192.560 73.570 192.820 ;
        RECT 42.890 192.220 43.210 192.480 ;
        RECT 46.200 192.420 46.340 192.560 ;
        RECT 43.440 192.280 46.340 192.420 ;
        RECT 46.585 192.420 46.875 192.465 ;
        RECT 47.030 192.420 47.350 192.480 ;
        RECT 46.585 192.280 49.560 192.420 ;
        RECT 43.440 192.125 43.580 192.280 ;
        RECT 46.585 192.235 46.875 192.280 ;
        RECT 47.030 192.220 47.350 192.280 ;
        RECT 43.365 191.895 43.655 192.125 ;
        RECT 44.285 192.080 44.575 192.125 ;
        RECT 45.650 192.080 45.970 192.140 ;
        RECT 44.285 191.940 45.970 192.080 ;
        RECT 44.285 191.895 44.575 191.940 ;
        RECT 45.650 191.880 45.970 191.940 ;
        RECT 46.110 191.880 46.430 192.140 ;
        RECT 49.420 192.125 49.560 192.280 ;
        RECT 51.630 192.125 51.950 192.140 ;
        RECT 47.965 192.080 48.255 192.125 ;
        RECT 49.345 192.080 49.635 192.125 ;
        RECT 51.630 192.080 51.970 192.125 ;
        RECT 47.965 191.940 48.640 192.080 ;
        RECT 47.965 191.895 48.255 191.940 ;
        RECT 44.745 191.400 45.035 191.445 ;
        RECT 48.500 191.400 48.640 191.940 ;
        RECT 49.345 191.940 51.355 192.080 ;
        RECT 49.345 191.895 49.635 191.940 ;
        RECT 49.805 191.740 50.095 191.785 ;
        RECT 50.710 191.740 51.030 191.800 ;
        RECT 49.805 191.600 51.030 191.740 ;
        RECT 51.215 191.740 51.355 191.940 ;
        RECT 51.630 191.940 52.145 192.080 ;
        RECT 51.630 191.895 51.970 191.940 ;
        RECT 51.630 191.880 51.950 191.895 ;
        RECT 52.105 191.740 52.395 191.785 ;
        RECT 60.920 191.740 61.060 192.560 ;
        RECT 110.010 192.545 110.150 205.860 ;
        RECT 111.010 201.530 111.150 206.310 ;
        RECT 111.360 205.830 111.620 206.150 ;
        RECT 111.420 202.635 111.560 205.830 ;
        RECT 111.330 202.375 111.650 202.635 ;
        RECT 111.010 201.390 111.640 201.530 ;
        RECT 111.500 198.530 111.640 201.390 ;
        RECT 111.410 198.200 111.740 198.530 ;
        RECT 64.065 192.420 64.355 192.465 ;
        RECT 70.950 192.420 71.270 192.480 ;
        RECT 64.065 192.280 71.270 192.420 ;
        RECT 64.065 192.235 64.355 192.280 ;
        RECT 70.950 192.220 71.270 192.280 ;
        RECT 72.345 192.420 72.635 192.465 ;
        RECT 75.565 192.420 75.855 192.465 ;
        RECT 72.345 192.280 75.855 192.420 ;
        RECT 72.345 192.235 72.635 192.280 ;
        RECT 75.565 192.235 75.855 192.280 ;
        RECT 109.950 192.225 110.210 192.545 ;
        RECT 63.130 192.080 63.450 192.140 ;
        RECT 65.445 192.080 65.735 192.125 ;
        RECT 66.365 192.080 66.655 192.125 ;
        RECT 63.130 191.940 65.735 192.080 ;
        RECT 63.130 191.880 63.450 191.940 ;
        RECT 65.445 191.895 65.735 191.940 ;
        RECT 65.980 191.940 66.655 192.080 ;
        RECT 51.215 191.600 61.060 191.740 ;
        RECT 64.050 191.740 64.370 191.800 ;
        RECT 65.980 191.740 66.120 191.940 ;
        RECT 66.365 191.895 66.655 191.940 ;
        RECT 66.825 191.895 67.115 192.125 ;
        RECT 67.285 191.895 67.575 192.125 ;
        RECT 68.190 192.080 68.510 192.140 ;
        RECT 68.665 192.080 68.955 192.125 ;
        RECT 68.190 191.940 68.955 192.080 ;
        RECT 66.900 191.740 67.040 191.895 ;
        RECT 64.050 191.600 66.120 191.740 ;
        RECT 66.440 191.600 67.040 191.740 ;
        RECT 67.360 191.740 67.500 191.895 ;
        RECT 68.190 191.880 68.510 191.940 ;
        RECT 68.665 191.895 68.955 191.940 ;
        RECT 69.570 191.880 69.890 192.140 ;
        RECT 70.045 192.080 70.335 192.125 ;
        RECT 70.045 191.940 70.720 192.080 ;
        RECT 70.045 191.895 70.335 191.940 ;
        RECT 70.580 191.740 70.720 191.940 ;
        RECT 71.870 191.880 72.190 192.140 ;
        RECT 73.725 191.895 74.015 192.125 ;
        RECT 70.950 191.740 71.270 191.800 ;
        RECT 73.800 191.740 73.940 191.895 ;
        RECT 74.630 191.880 74.950 192.140 ;
        RECT 67.360 191.600 73.940 191.740 ;
        RECT 49.805 191.555 50.095 191.600 ;
        RECT 50.710 191.540 51.030 191.600 ;
        RECT 52.105 191.555 52.395 191.600 ;
        RECT 64.050 191.540 64.370 191.600 ;
        RECT 66.440 191.460 66.580 191.600 ;
        RECT 70.950 191.540 71.270 191.600 ;
        RECT 49.330 191.400 49.650 191.460 ;
        RECT 44.745 191.260 49.650 191.400 ;
        RECT 44.745 191.215 45.035 191.260 ;
        RECT 49.330 191.200 49.650 191.260 ;
        RECT 66.350 191.200 66.670 191.460 ;
        RECT 68.650 191.200 68.970 191.460 ;
        RECT 70.505 191.400 70.795 191.445 ;
        RECT 69.890 191.260 70.795 191.400 ;
        RECT 41.970 190.860 42.290 191.120 ;
        RECT 42.430 191.060 42.750 191.120 ;
        RECT 47.505 191.060 47.795 191.105 ;
        RECT 42.430 190.920 47.795 191.060 ;
        RECT 42.430 190.860 42.750 190.920 ;
        RECT 47.505 190.875 47.795 190.920 ;
        RECT 62.210 191.060 62.530 191.120 ;
        RECT 62.685 191.060 62.975 191.105 ;
        RECT 62.210 190.920 62.975 191.060 ;
        RECT 62.210 190.860 62.530 190.920 ;
        RECT 62.685 190.875 62.975 190.920 ;
        RECT 63.590 191.060 63.910 191.120 ;
        RECT 67.270 191.060 67.590 191.120 ;
        RECT 69.890 191.060 70.030 191.260 ;
        RECT 70.505 191.215 70.795 191.260 ;
        RECT 63.590 190.920 70.030 191.060 ;
        RECT 63.590 190.860 63.910 190.920 ;
        RECT 67.270 190.860 67.590 190.920 ;
        RECT 13.380 190.240 92.040 190.720 ;
        RECT 41.970 190.040 42.290 190.100 ;
        RECT 42.445 190.040 42.735 190.085 ;
        RECT 51.170 190.040 51.490 190.100 ;
        RECT 41.970 189.900 51.490 190.040 ;
        RECT 41.970 189.840 42.290 189.900 ;
        RECT 42.445 189.855 42.735 189.900 ;
        RECT 51.170 189.840 51.490 189.900 ;
        RECT 65.430 189.840 65.750 190.100 ;
        RECT 66.350 189.840 66.670 190.100 ;
        RECT 71.425 190.040 71.715 190.085 ;
        RECT 71.870 190.040 72.190 190.100 ;
        RECT 71.425 189.900 72.190 190.040 ;
        RECT 71.425 189.855 71.715 189.900 ;
        RECT 71.870 189.840 72.190 189.900 ;
        RECT 58.545 189.700 58.835 189.745 ;
        RECT 60.830 189.700 61.150 189.760 ;
        RECT 58.545 189.560 61.150 189.700 ;
        RECT 58.545 189.515 58.835 189.560 ;
        RECT 60.830 189.500 61.150 189.560 ;
        RECT 62.210 189.700 62.530 189.760 ;
        RECT 62.210 189.560 64.740 189.700 ;
        RECT 62.210 189.500 62.530 189.560 ;
        RECT 64.600 189.405 64.740 189.560 ;
        RECT 61.305 189.360 61.595 189.405 ;
        RECT 57.700 189.220 60.600 189.360 ;
        RECT 57.700 189.080 57.840 189.220 ;
        RECT 42.890 188.820 43.210 189.080 ;
        RECT 57.150 188.820 57.470 189.080 ;
        RECT 57.610 188.820 57.930 189.080 ;
        RECT 60.460 189.065 60.600 189.220 ;
        RECT 61.305 189.220 63.360 189.360 ;
        RECT 61.305 189.175 61.595 189.220 ;
        RECT 63.220 189.080 63.360 189.220 ;
        RECT 64.525 189.175 64.815 189.405 ;
        RECT 66.350 189.360 66.670 189.420 ;
        RECT 69.570 189.360 69.890 189.420 ;
        RECT 66.350 189.220 72.100 189.360 ;
        RECT 66.350 189.160 66.670 189.220 ;
        RECT 69.570 189.160 69.890 189.220 ;
        RECT 59.925 189.020 60.215 189.065 ;
        RECT 58.160 188.880 60.215 189.020 ;
        RECT 42.980 188.680 43.120 188.820 ;
        RECT 43.365 188.680 43.655 188.725 ;
        RECT 42.980 188.540 43.655 188.680 ;
        RECT 57.240 188.680 57.380 188.820 ;
        RECT 58.160 188.680 58.300 188.880 ;
        RECT 59.925 188.835 60.215 188.880 ;
        RECT 60.385 188.835 60.675 189.065 ;
        RECT 61.750 188.820 62.070 189.080 ;
        RECT 63.130 188.820 63.450 189.080 ;
        RECT 64.050 188.820 64.370 189.080 ;
        RECT 70.950 189.020 71.270 189.080 ;
        RECT 71.960 189.065 72.100 189.220 ;
        RECT 66.900 188.880 71.270 189.020 ;
        RECT 57.240 188.540 58.300 188.680 ;
        RECT 58.545 188.680 58.835 188.725 ;
        RECT 62.225 188.680 62.515 188.725 ;
        RECT 58.545 188.540 62.515 188.680 ;
        RECT 43.365 188.495 43.655 188.540 ;
        RECT 58.545 188.495 58.835 188.540 ;
        RECT 62.225 188.495 62.515 188.540 ;
        RECT 66.285 188.680 66.575 188.725 ;
        RECT 66.900 188.680 67.040 188.880 ;
        RECT 70.950 188.820 71.270 188.880 ;
        RECT 71.885 189.020 72.175 189.065 ;
        RECT 74.630 189.020 74.950 189.080 ;
        RECT 71.885 188.880 74.950 189.020 ;
        RECT 71.885 188.835 72.175 188.880 ;
        RECT 74.630 188.820 74.950 188.880 ;
        RECT 66.285 188.540 67.040 188.680 ;
        RECT 67.285 188.680 67.575 188.725 ;
        RECT 68.190 188.680 68.510 188.740 ;
        RECT 67.285 188.540 68.510 188.680 ;
        RECT 71.040 188.680 71.180 188.820 ;
        RECT 72.790 188.680 73.110 188.740 ;
        RECT 71.040 188.540 73.110 188.680 ;
        RECT 66.285 188.495 66.575 188.540 ;
        RECT 67.285 188.495 67.575 188.540 ;
        RECT 41.510 188.140 41.830 188.400 ;
        RECT 42.365 188.340 42.655 188.385 ;
        RECT 42.890 188.340 43.210 188.400 ;
        RECT 42.365 188.200 43.210 188.340 ;
        RECT 42.365 188.155 42.655 188.200 ;
        RECT 42.890 188.140 43.210 188.200 ;
        RECT 58.070 188.340 58.390 188.400 ;
        RECT 59.005 188.340 59.295 188.385 ;
        RECT 58.070 188.200 59.295 188.340 ;
        RECT 58.070 188.140 58.390 188.200 ;
        RECT 59.005 188.155 59.295 188.200 ;
        RECT 64.050 188.340 64.370 188.400 ;
        RECT 67.360 188.340 67.500 188.495 ;
        RECT 68.190 188.480 68.510 188.540 ;
        RECT 72.790 188.480 73.110 188.540 ;
        RECT 64.050 188.200 67.500 188.340 ;
        RECT 64.050 188.140 64.370 188.200 ;
        RECT 13.380 187.520 92.040 188.000 ;
        RECT 57.165 187.320 57.455 187.365 ;
        RECT 57.610 187.320 57.930 187.380 ;
        RECT 57.165 187.180 57.930 187.320 ;
        RECT 57.165 187.135 57.455 187.180 ;
        RECT 57.610 187.120 57.930 187.180 ;
        RECT 22.650 187.025 22.970 187.040 ;
        RECT 22.585 186.795 22.970 187.025 ;
        RECT 23.585 186.795 23.875 187.025 ;
        RECT 41.020 186.980 41.310 187.025 ;
        RECT 41.510 186.980 41.830 187.040 ;
        RECT 41.020 186.840 41.830 186.980 ;
        RECT 41.020 186.795 41.310 186.840 ;
        RECT 22.650 186.780 22.970 186.795 ;
        RECT 18.050 186.300 18.370 186.360 ;
        RECT 23.660 186.300 23.800 186.795 ;
        RECT 41.510 186.780 41.830 186.840 ;
        RECT 53.010 186.980 53.330 187.040 ;
        RECT 63.590 186.980 63.910 187.040 ;
        RECT 53.010 186.840 63.910 186.980 ;
        RECT 53.010 186.780 53.330 186.840 ;
        RECT 63.590 186.780 63.910 186.840 ;
        RECT 28.170 186.640 28.490 186.700 ;
        RECT 29.005 186.640 29.295 186.685 ;
        RECT 28.170 186.500 29.295 186.640 ;
        RECT 28.170 186.440 28.490 186.500 ;
        RECT 29.005 186.455 29.295 186.500 ;
        RECT 38.290 186.640 38.610 186.700 ;
        RECT 39.685 186.640 39.975 186.685 ;
        RECT 38.290 186.500 39.975 186.640 ;
        RECT 38.290 186.440 38.610 186.500 ;
        RECT 39.685 186.455 39.975 186.500 ;
        RECT 56.705 186.455 56.995 186.685 ;
        RECT 18.050 186.160 23.800 186.300 ;
        RECT 25.870 186.300 26.190 186.360 ;
        RECT 27.725 186.300 28.015 186.345 ;
        RECT 25.870 186.160 28.015 186.300 ;
        RECT 18.050 186.100 18.370 186.160 ;
        RECT 25.870 186.100 26.190 186.160 ;
        RECT 27.725 186.115 28.015 186.160 ;
        RECT 28.605 186.300 28.895 186.345 ;
        RECT 29.795 186.300 30.085 186.345 ;
        RECT 32.315 186.300 32.605 186.345 ;
        RECT 28.605 186.160 32.605 186.300 ;
        RECT 28.605 186.115 28.895 186.160 ;
        RECT 29.795 186.115 30.085 186.160 ;
        RECT 32.315 186.115 32.605 186.160 ;
        RECT 40.565 186.300 40.855 186.345 ;
        RECT 41.755 186.300 42.045 186.345 ;
        RECT 44.275 186.300 44.565 186.345 ;
        RECT 40.565 186.160 44.565 186.300 ;
        RECT 56.780 186.300 56.920 186.455 ;
        RECT 58.070 186.440 58.390 186.700 ;
        RECT 59.910 186.640 60.230 186.700 ;
        RECT 60.845 186.640 61.135 186.685 ;
        RECT 59.910 186.500 61.135 186.640 ;
        RECT 59.910 186.440 60.230 186.500 ;
        RECT 60.845 186.455 61.135 186.500 ;
        RECT 61.305 186.640 61.595 186.685 ;
        RECT 64.050 186.640 64.370 186.700 ;
        RECT 61.305 186.500 64.370 186.640 ;
        RECT 61.305 186.455 61.595 186.500 ;
        RECT 64.050 186.440 64.370 186.500 ;
        RECT 57.150 186.300 57.470 186.360 ;
        RECT 58.990 186.300 59.310 186.360 ;
        RECT 56.780 186.160 59.310 186.300 ;
        RECT 40.565 186.115 40.855 186.160 ;
        RECT 41.755 186.115 42.045 186.160 ;
        RECT 44.275 186.115 44.565 186.160 ;
        RECT 57.150 186.100 57.470 186.160 ;
        RECT 58.990 186.100 59.310 186.160 ;
        RECT 62.225 186.300 62.515 186.345 ;
        RECT 66.350 186.300 66.670 186.360 ;
        RECT 62.225 186.160 66.670 186.300 ;
        RECT 62.225 186.115 62.515 186.160 ;
        RECT 66.350 186.100 66.670 186.160 ;
        RECT 28.210 185.960 28.500 186.005 ;
        RECT 30.310 185.960 30.600 186.005 ;
        RECT 31.880 185.960 32.170 186.005 ;
        RECT 28.210 185.820 32.170 185.960 ;
        RECT 28.210 185.775 28.500 185.820 ;
        RECT 30.310 185.775 30.600 185.820 ;
        RECT 31.880 185.775 32.170 185.820 ;
        RECT 40.170 185.960 40.460 186.005 ;
        RECT 42.270 185.960 42.560 186.005 ;
        RECT 43.840 185.960 44.130 186.005 ;
        RECT 40.170 185.820 44.130 185.960 ;
        RECT 40.170 185.775 40.460 185.820 ;
        RECT 42.270 185.775 42.560 185.820 ;
        RECT 43.840 185.775 44.130 185.820 ;
        RECT 47.490 185.960 47.810 186.020 ;
        RECT 48.870 185.960 49.190 186.020 ;
        RECT 68.650 185.960 68.970 186.020 ;
        RECT 47.490 185.820 68.970 185.960 ;
        RECT 47.490 185.760 47.810 185.820 ;
        RECT 48.870 185.760 49.190 185.820 ;
        RECT 68.650 185.760 68.970 185.820 ;
        RECT 21.730 185.420 22.050 185.680 ;
        RECT 22.665 185.620 22.955 185.665 ;
        RECT 27.710 185.620 28.030 185.680 ;
        RECT 22.665 185.480 28.030 185.620 ;
        RECT 22.665 185.435 22.955 185.480 ;
        RECT 27.710 185.420 28.030 185.480 ;
        RECT 34.610 185.420 34.930 185.680 ;
        RECT 44.270 185.620 44.590 185.680 ;
        RECT 46.585 185.620 46.875 185.665 ;
        RECT 44.270 185.480 46.875 185.620 ;
        RECT 44.270 185.420 44.590 185.480 ;
        RECT 46.585 185.435 46.875 185.480 ;
        RECT 58.085 185.620 58.375 185.665 ;
        RECT 60.370 185.620 60.690 185.680 ;
        RECT 58.085 185.480 60.690 185.620 ;
        RECT 58.085 185.435 58.375 185.480 ;
        RECT 60.370 185.420 60.690 185.480 ;
        RECT 61.750 185.420 62.070 185.680 ;
        RECT 13.380 184.800 92.040 185.280 ;
        RECT 18.050 184.400 18.370 184.660 ;
        RECT 27.725 184.600 28.015 184.645 ;
        RECT 28.170 184.600 28.490 184.660 ;
        RECT 27.725 184.460 28.490 184.600 ;
        RECT 27.725 184.415 28.015 184.460 ;
        RECT 28.170 184.400 28.490 184.460 ;
        RECT 28.630 184.400 28.950 184.660 ;
        RECT 38.305 184.600 38.595 184.645 ;
        RECT 29.180 184.460 38.595 184.600 ;
        RECT 21.730 184.260 22.020 184.305 ;
        RECT 23.300 184.260 23.590 184.305 ;
        RECT 25.400 184.260 25.690 184.305 ;
        RECT 21.730 184.120 25.690 184.260 ;
        RECT 21.730 184.075 22.020 184.120 ;
        RECT 23.300 184.075 23.590 184.120 ;
        RECT 25.400 184.075 25.690 184.120 ;
        RECT 21.295 183.920 21.585 183.965 ;
        RECT 23.815 183.920 24.105 183.965 ;
        RECT 25.005 183.920 25.295 183.965 ;
        RECT 21.295 183.780 25.295 183.920 ;
        RECT 21.295 183.735 21.585 183.780 ;
        RECT 23.815 183.735 24.105 183.780 ;
        RECT 25.005 183.735 25.295 183.780 ;
        RECT 17.605 183.395 17.895 183.625 ;
        RECT 17.680 183.240 17.820 183.395 ;
        RECT 18.510 183.380 18.830 183.640 ;
        RECT 21.730 183.580 22.050 183.640 ;
        RECT 24.550 183.580 24.840 183.625 ;
        RECT 21.730 183.440 24.840 183.580 ;
        RECT 21.730 183.380 22.050 183.440 ;
        RECT 24.550 183.395 24.840 183.440 ;
        RECT 25.870 183.380 26.190 183.640 ;
        RECT 28.565 183.240 28.855 183.285 ;
        RECT 29.180 183.240 29.320 184.460 ;
        RECT 38.305 184.415 38.595 184.460 ;
        RECT 42.890 184.400 43.210 184.660 ;
        RECT 58.070 184.600 58.390 184.660 ;
        RECT 64.970 184.600 65.290 184.660 ;
        RECT 58.070 184.460 65.290 184.600 ;
        RECT 58.070 184.400 58.390 184.460 ;
        RECT 31.020 184.120 36.680 184.260 ;
        RECT 30.470 183.580 30.790 183.640 ;
        RECT 31.020 183.625 31.160 184.120 ;
        RECT 31.390 183.920 31.710 183.980 ;
        RECT 31.390 183.780 34.380 183.920 ;
        RECT 31.390 183.720 31.710 183.780 ;
        RECT 30.945 183.580 31.235 183.625 ;
        RECT 30.470 183.440 31.235 183.580 ;
        RECT 30.470 183.380 30.790 183.440 ;
        RECT 30.945 183.395 31.235 183.440 ;
        RECT 31.850 183.380 32.170 183.640 ;
        RECT 32.310 183.380 32.630 183.640 ;
        RECT 34.240 183.625 34.380 183.780 ;
        RECT 34.165 183.580 34.455 183.625 ;
        RECT 34.610 183.580 34.930 183.640 ;
        RECT 34.165 183.440 34.930 183.580 ;
        RECT 35.160 183.590 35.300 184.120 ;
        RECT 36.540 183.920 36.680 184.120 ;
        RECT 41.525 183.920 41.815 183.965 ;
        RECT 42.430 183.920 42.750 183.980 ;
        RECT 36.540 183.780 39.900 183.920 ;
        RECT 35.545 183.590 35.835 183.625 ;
        RECT 35.160 183.450 35.835 183.590 ;
        RECT 34.165 183.395 34.455 183.440 ;
        RECT 34.610 183.380 34.930 183.440 ;
        RECT 35.545 183.395 35.835 183.450 ;
        RECT 35.990 183.380 36.310 183.640 ;
        RECT 36.540 183.580 36.680 183.780 ;
        RECT 36.925 183.580 37.215 183.625 ;
        RECT 36.540 183.440 37.215 183.580 ;
        RECT 36.925 183.395 37.215 183.440 ;
        RECT 37.370 183.380 37.690 183.640 ;
        RECT 39.760 183.625 39.900 183.780 ;
        RECT 41.525 183.780 42.750 183.920 ;
        RECT 41.525 183.735 41.815 183.780 ;
        RECT 42.430 183.720 42.750 183.780 ;
        RECT 38.305 183.580 38.595 183.625 ;
        RECT 38.305 183.440 39.440 183.580 ;
        RECT 38.305 183.395 38.595 183.440 ;
        RECT 17.680 183.100 19.200 183.240 ;
        RECT 19.060 182.945 19.200 183.100 ;
        RECT 28.565 183.100 29.320 183.240 ;
        RECT 29.565 183.240 29.855 183.285 ;
        RECT 33.245 183.240 33.535 183.285 ;
        RECT 33.690 183.240 34.010 183.300 ;
        RECT 29.565 183.100 34.010 183.240 ;
        RECT 34.700 183.240 34.840 183.380 ;
        RECT 38.765 183.240 39.055 183.285 ;
        RECT 34.700 183.100 39.055 183.240 ;
        RECT 28.565 183.055 28.855 183.100 ;
        RECT 29.565 183.055 29.855 183.100 ;
        RECT 33.245 183.055 33.535 183.100 ;
        RECT 33.690 183.040 34.010 183.100 ;
        RECT 38.765 183.055 39.055 183.100 ;
        RECT 18.985 182.900 19.275 182.945 ;
        RECT 24.030 182.900 24.350 182.960 ;
        RECT 18.985 182.760 24.350 182.900 ;
        RECT 18.985 182.715 19.275 182.760 ;
        RECT 24.030 182.700 24.350 182.760 ;
        RECT 30.025 182.900 30.315 182.945 ;
        RECT 30.930 182.900 31.250 182.960 ;
        RECT 30.025 182.760 31.250 182.900 ;
        RECT 30.025 182.715 30.315 182.760 ;
        RECT 30.930 182.700 31.250 182.760 ;
        RECT 32.770 182.900 33.090 182.960 ;
        RECT 34.610 182.900 34.930 182.960 ;
        RECT 35.085 182.900 35.375 182.945 ;
        RECT 39.300 182.900 39.440 183.440 ;
        RECT 39.685 183.395 39.975 183.625 ;
        RECT 41.065 183.580 41.355 183.625 ;
        RECT 43.810 183.580 44.130 183.640 ;
        RECT 41.065 183.440 44.130 183.580 ;
        RECT 41.065 183.395 41.355 183.440 ;
        RECT 43.810 183.380 44.130 183.440 ;
        RECT 53.470 183.380 53.790 183.640 ;
        RECT 54.865 183.580 55.155 183.625 ;
        RECT 57.610 183.580 57.930 183.640 ;
        RECT 59.540 183.625 59.680 184.460 ;
        RECT 64.970 184.400 65.290 184.460 ;
        RECT 68.650 184.600 68.970 184.660 ;
        RECT 69.125 184.600 69.415 184.645 ;
        RECT 68.650 184.460 69.415 184.600 ;
        RECT 68.650 184.400 68.970 184.460 ;
        RECT 69.125 184.415 69.415 184.460 ;
        RECT 60.845 184.260 61.135 184.305 ;
        RECT 61.750 184.260 62.070 184.320 ;
        RECT 60.845 184.120 62.070 184.260 ;
        RECT 60.845 184.075 61.135 184.120 ;
        RECT 61.750 184.060 62.070 184.120 ;
        RECT 68.190 184.260 68.510 184.320 ;
        RECT 70.505 184.260 70.795 184.305 ;
        RECT 68.190 184.120 70.795 184.260 ;
        RECT 68.190 184.060 68.510 184.120 ;
        RECT 70.505 184.075 70.795 184.120 ;
        RECT 73.250 184.260 73.540 184.305 ;
        RECT 74.820 184.260 75.110 184.305 ;
        RECT 76.920 184.260 77.210 184.305 ;
        RECT 73.250 184.120 77.210 184.260 ;
        RECT 73.250 184.075 73.540 184.120 ;
        RECT 74.820 184.075 75.110 184.120 ;
        RECT 76.920 184.075 77.210 184.120 ;
        RECT 62.760 183.780 64.740 183.920 ;
        RECT 54.865 183.440 57.930 183.580 ;
        RECT 54.865 183.395 55.155 183.440 ;
        RECT 57.610 183.380 57.930 183.440 ;
        RECT 59.465 183.395 59.755 183.625 ;
        RECT 60.385 183.580 60.675 183.625 ;
        RECT 60.830 183.580 61.150 183.640 ;
        RECT 60.385 183.440 61.150 183.580 ;
        RECT 60.385 183.395 60.675 183.440 ;
        RECT 60.830 183.380 61.150 183.440 ;
        RECT 61.305 183.395 61.595 183.625 ;
        RECT 61.765 183.590 62.055 183.625 ;
        RECT 62.760 183.590 62.900 183.780 ;
        RECT 61.765 183.450 62.900 183.590 ;
        RECT 63.590 183.580 63.910 183.640 ;
        RECT 64.065 183.580 64.355 183.625 ;
        RECT 61.765 183.395 62.055 183.450 ;
        RECT 63.590 183.440 64.355 183.580 ;
        RECT 64.600 183.580 64.740 183.780 ;
        RECT 64.970 183.720 65.290 183.980 ;
        RECT 72.815 183.920 73.105 183.965 ;
        RECT 75.335 183.920 75.625 183.965 ;
        RECT 76.525 183.920 76.815 183.965 ;
        RECT 72.815 183.780 76.815 183.920 ;
        RECT 72.815 183.735 73.105 183.780 ;
        RECT 75.335 183.735 75.625 183.780 ;
        RECT 76.525 183.735 76.815 183.780 ;
        RECT 77.390 183.720 77.710 183.980 ;
        RECT 64.600 183.440 65.200 183.580 ;
        RECT 43.350 183.240 43.670 183.300 ;
        RECT 47.965 183.240 48.255 183.285 ;
        RECT 43.350 183.100 48.255 183.240 ;
        RECT 43.350 183.040 43.670 183.100 ;
        RECT 47.965 183.055 48.255 183.100 ;
        RECT 50.710 183.240 51.030 183.300 ;
        RECT 54.405 183.240 54.695 183.285 ;
        RECT 50.710 183.100 54.695 183.240 ;
        RECT 61.380 183.240 61.520 183.395 ;
        RECT 63.590 183.380 63.910 183.440 ;
        RECT 64.065 183.395 64.355 183.440 ;
        RECT 64.510 183.240 64.830 183.300 ;
        RECT 61.380 183.100 64.830 183.240 ;
        RECT 65.060 183.240 65.200 183.440 ;
        RECT 65.430 183.380 65.750 183.640 ;
        RECT 67.285 183.580 67.575 183.625 ;
        RECT 73.250 183.580 73.570 183.640 ;
        RECT 67.285 183.440 73.570 183.580 ;
        RECT 67.285 183.395 67.575 183.440 ;
        RECT 73.250 183.380 73.570 183.440 ;
        RECT 65.905 183.240 66.195 183.285 ;
        RECT 65.060 183.100 66.195 183.240 ;
        RECT 50.710 183.040 51.030 183.100 ;
        RECT 54.405 183.055 54.695 183.100 ;
        RECT 64.510 183.040 64.830 183.100 ;
        RECT 65.905 183.055 66.195 183.100 ;
        RECT 71.870 183.240 72.190 183.300 ;
        RECT 76.070 183.240 76.360 183.285 ;
        RECT 71.870 183.100 76.360 183.240 ;
        RECT 71.870 183.040 72.190 183.100 ;
        RECT 76.070 183.055 76.360 183.100 ;
        RECT 32.770 182.760 39.440 182.900 ;
        RECT 45.190 182.900 45.510 182.960 ;
        RECT 47.505 182.900 47.795 182.945 ;
        RECT 48.870 182.900 49.190 182.960 ;
        RECT 45.190 182.760 49.190 182.900 ;
        RECT 32.770 182.700 33.090 182.760 ;
        RECT 34.610 182.700 34.930 182.760 ;
        RECT 35.085 182.715 35.375 182.760 ;
        RECT 45.190 182.700 45.510 182.760 ;
        RECT 47.505 182.715 47.795 182.760 ;
        RECT 48.870 182.700 49.190 182.760 ;
        RECT 52.565 182.900 52.855 182.945 ;
        RECT 53.010 182.900 53.330 182.960 ;
        RECT 52.565 182.760 53.330 182.900 ;
        RECT 52.565 182.715 52.855 182.760 ;
        RECT 53.010 182.700 53.330 182.760 ;
        RECT 60.830 182.900 61.150 182.960 ;
        RECT 62.685 182.900 62.975 182.945 ;
        RECT 60.830 182.760 62.975 182.900 ;
        RECT 60.830 182.700 61.150 182.760 ;
        RECT 62.685 182.715 62.975 182.760 ;
        RECT 63.130 182.700 63.450 182.960 ;
        RECT 69.110 182.700 69.430 182.960 ;
        RECT 70.030 182.700 70.350 182.960 ;
        RECT 13.380 182.080 92.040 182.560 ;
        RECT 100.970 182.410 102.630 184.070 ;
        RECT 112.120 183.415 112.600 219.295 ;
        RECT 113.420 207.865 113.680 208.185 ;
        RECT 112.755 206.960 112.985 207.250 ;
        RECT 112.800 205.425 112.940 206.960 ;
        RECT 112.740 205.105 113.000 205.425 ;
        RECT 112.755 204.660 112.985 204.950 ;
        RECT 112.800 202.665 112.940 204.660 ;
        RECT 113.435 203.955 113.665 204.030 ;
        RECT 113.435 203.815 114.640 203.955 ;
        RECT 113.435 203.740 113.665 203.815 ;
        RECT 113.435 203.280 113.665 203.570 ;
        RECT 113.480 203.125 113.620 203.280 ;
        RECT 113.420 202.805 113.680 203.125 ;
        RECT 114.115 202.795 114.345 203.085 ;
        RECT 112.740 202.345 113.000 202.665 ;
        RECT 113.775 202.400 114.005 202.690 ;
        RECT 113.095 201.945 113.325 202.235 ;
        RECT 113.140 200.825 113.280 201.945 ;
        RECT 113.820 201.500 113.960 202.400 ;
        RECT 113.775 201.210 114.005 201.500 ;
        RECT 113.080 200.505 113.340 200.825 ;
        RECT 113.820 198.980 113.960 201.210 ;
        RECT 114.160 200.985 114.300 202.795 ;
        RECT 114.115 200.695 114.345 200.985 ;
        RECT 114.160 199.415 114.300 200.695 ;
        RECT 114.115 199.125 114.345 199.415 ;
        RECT 113.775 198.690 114.005 198.980 ;
        RECT 112.740 198.435 113.000 198.525 ;
        RECT 112.740 198.295 113.280 198.435 ;
        RECT 112.740 198.205 113.000 198.295 ;
        RECT 112.755 195.675 112.985 195.750 ;
        RECT 113.140 195.675 113.280 198.295 ;
        RECT 114.500 198.065 114.640 203.815 ;
        RECT 114.440 197.745 114.700 198.065 ;
        RECT 114.115 196.380 114.345 196.670 ;
        RECT 112.755 195.535 113.280 195.675 ;
        RECT 112.755 195.460 112.985 195.535 ;
        RECT 114.160 194.845 114.300 196.380 ;
        RECT 113.420 194.525 113.680 194.845 ;
        RECT 114.100 194.525 114.360 194.845 ;
        RECT 112.740 192.225 113.000 192.545 ;
        RECT 112.800 191.150 112.940 192.225 ;
        RECT 113.420 191.765 113.680 192.085 ;
        RECT 112.755 190.860 112.985 191.150 ;
        RECT 114.455 189.940 114.685 190.230 ;
        RECT 113.760 189.465 114.020 189.785 ;
        RECT 113.420 189.005 113.680 189.325 ;
        RECT 113.820 187.930 113.960 189.465 ;
        RECT 114.100 188.545 114.360 188.865 ;
        RECT 113.775 187.640 114.005 187.930 ;
        RECT 114.160 186.550 114.300 188.545 ;
        RECT 114.500 188.405 114.640 189.940 ;
        RECT 114.440 188.085 114.700 188.405 ;
        RECT 114.115 186.260 114.345 186.550 ;
        RECT 114.440 185.785 114.700 186.105 ;
        RECT 114.500 185.630 114.640 185.785 ;
        RECT 114.455 185.340 114.685 185.630 ;
        RECT 114.840 183.415 115.320 219.295 ;
        RECT 115.860 217.370 116.000 220.285 ;
        RECT 148.630 220.050 148.950 220.310 ;
        RECT 148.140 219.570 148.400 219.890 ;
        RECT 116.480 217.525 116.740 217.845 ;
        RECT 115.815 217.080 116.045 217.370 ;
        RECT 116.540 216.450 116.680 217.525 ;
        RECT 116.495 216.160 116.725 216.450 ;
        RECT 117.160 214.765 117.420 215.085 ;
        RECT 117.160 212.925 117.420 213.245 ;
        RECT 117.160 212.465 117.420 212.785 ;
        RECT 116.155 211.560 116.385 211.850 ;
        RECT 116.200 206.345 116.340 211.560 ;
        RECT 117.160 210.165 117.420 210.485 ;
        RECT 117.220 208.185 117.360 210.165 ;
        RECT 117.160 207.865 117.420 208.185 ;
        RECT 116.140 206.025 116.400 206.345 ;
        RECT 117.220 205.870 117.360 207.865 ;
        RECT 117.175 205.580 117.405 205.870 ;
        RECT 116.155 203.270 116.385 203.560 ;
        RECT 115.815 202.835 116.045 203.125 ;
        RECT 115.860 201.555 116.000 202.835 ;
        RECT 115.815 201.265 116.045 201.555 ;
        RECT 115.460 200.505 115.720 200.825 ;
        RECT 115.520 198.510 115.660 200.505 ;
        RECT 115.860 199.455 116.000 201.265 ;
        RECT 116.200 201.040 116.340 203.270 ;
        RECT 117.160 201.655 117.420 201.745 ;
        RECT 116.540 201.515 117.420 201.655 ;
        RECT 116.155 200.750 116.385 201.040 ;
        RECT 116.200 199.850 116.340 200.750 ;
        RECT 116.540 200.305 116.680 201.515 ;
        RECT 117.160 201.425 117.420 201.515 ;
        RECT 116.820 200.505 117.080 200.825 ;
        RECT 116.495 200.015 116.725 200.305 ;
        RECT 116.155 199.560 116.385 199.850 ;
        RECT 115.815 199.165 116.045 199.455 ;
        RECT 116.495 198.895 116.725 198.970 ;
        RECT 116.880 198.895 117.020 200.505 ;
        RECT 116.495 198.755 117.020 198.895 ;
        RECT 116.495 198.680 116.725 198.755 ;
        RECT 115.475 198.220 115.705 198.510 ;
        RECT 116.495 196.380 116.725 196.670 ;
        RECT 116.140 194.985 116.400 195.305 ;
        RECT 116.140 194.525 116.400 194.845 ;
        RECT 116.200 190.230 116.340 194.525 ;
        RECT 116.540 192.990 116.680 196.380 ;
        RECT 117.160 195.905 117.420 196.225 ;
        RECT 116.495 192.700 116.725 192.990 ;
        RECT 116.155 189.940 116.385 190.230 ;
        RECT 116.140 189.465 116.400 189.785 ;
        RECT 116.200 188.390 116.340 189.465 ;
        RECT 116.480 189.005 116.740 189.325 ;
        RECT 116.155 188.100 116.385 188.390 ;
        RECT 116.155 187.640 116.385 187.930 ;
        RECT 116.200 185.185 116.340 187.640 ;
        RECT 116.540 187.010 116.680 189.005 ;
        RECT 116.495 186.720 116.725 187.010 ;
        RECT 117.160 186.245 117.420 186.565 ;
        RECT 117.220 186.090 117.360 186.245 ;
        RECT 117.175 185.800 117.405 186.090 ;
        RECT 116.140 184.865 116.400 185.185 ;
        RECT 117.560 183.415 118.040 219.295 ;
        RECT 119.880 217.525 120.140 217.845 ;
        RECT 119.215 215.230 119.445 215.520 ;
        RECT 118.520 214.765 118.780 215.085 ;
        RECT 118.580 212.265 118.720 214.765 ;
        RECT 119.260 213.000 119.400 215.230 ;
        RECT 119.555 214.795 119.785 215.085 ;
        RECT 119.600 213.515 119.740 214.795 ;
        RECT 119.555 213.225 119.785 213.515 ;
        RECT 119.215 212.710 119.445 213.000 ;
        RECT 118.535 211.975 118.765 212.265 ;
        RECT 119.260 211.810 119.400 212.710 ;
        RECT 119.215 211.520 119.445 211.810 ;
        RECT 119.600 211.415 119.740 213.225 ;
        RECT 119.555 211.125 119.785 211.415 ;
        RECT 119.200 210.625 119.460 210.945 ;
        RECT 118.875 205.580 119.105 205.870 ;
        RECT 118.920 201.285 119.060 205.580 ;
        RECT 118.860 200.965 119.120 201.285 ;
        RECT 119.880 200.505 120.140 200.825 ;
        RECT 119.940 199.430 120.080 200.505 ;
        RECT 119.895 199.140 120.125 199.430 ;
        RECT 118.875 195.215 119.105 195.290 ;
        RECT 118.875 195.075 119.400 195.215 ;
        RECT 118.875 195.000 119.105 195.075 ;
        RECT 118.860 193.605 119.120 193.925 ;
        RECT 118.195 192.915 118.425 192.990 ;
        RECT 118.195 192.775 118.720 192.915 ;
        RECT 118.195 192.700 118.425 192.775 ;
        RECT 118.195 189.940 118.425 190.230 ;
        RECT 118.240 189.785 118.380 189.940 ;
        RECT 118.180 189.465 118.440 189.785 ;
        RECT 118.580 189.695 118.720 192.775 ;
        RECT 118.860 192.225 119.120 192.545 ;
        RECT 118.860 190.845 119.120 191.165 ;
        RECT 118.875 189.695 119.105 189.770 ;
        RECT 118.580 189.555 119.105 189.695 ;
        RECT 118.180 189.005 118.440 189.325 ;
        RECT 118.580 187.395 118.720 189.555 ;
        RECT 118.875 189.480 119.105 189.555 ;
        RECT 118.875 188.560 119.105 188.850 ;
        RECT 118.920 188.405 119.060 188.560 ;
        RECT 118.860 188.085 119.120 188.405 ;
        RECT 118.860 187.395 119.120 187.485 ;
        RECT 118.580 187.255 119.120 187.395 ;
        RECT 118.860 187.165 119.120 187.255 ;
        RECT 118.860 185.785 119.120 186.105 ;
        RECT 119.260 185.645 119.400 195.075 ;
        RECT 119.555 194.080 119.785 194.370 ;
        RECT 119.600 188.865 119.740 194.080 ;
        RECT 119.895 191.320 120.125 191.610 ;
        RECT 119.940 189.325 120.080 191.320 ;
        RECT 119.880 189.005 120.140 189.325 ;
        RECT 119.540 188.545 119.800 188.865 ;
        RECT 119.895 188.100 120.125 188.390 ;
        RECT 119.940 187.945 120.080 188.100 ;
        RECT 119.880 187.625 120.140 187.945 ;
        RECT 119.200 185.325 119.460 185.645 ;
        RECT 118.860 184.865 119.120 185.185 ;
        RECT 120.280 183.415 120.760 219.295 ;
        RECT 121.240 217.985 121.500 218.305 ;
        RECT 121.300 217.370 121.440 217.985 ;
        RECT 121.580 217.525 121.840 217.845 ;
        RECT 121.255 217.080 121.485 217.370 ;
        RECT 121.640 215.070 121.780 217.525 ;
        RECT 121.935 216.160 122.165 216.450 ;
        RECT 121.595 214.780 121.825 215.070 ;
        RECT 120.900 212.925 121.160 213.245 ;
        RECT 120.960 211.850 121.100 212.925 ;
        RECT 121.240 212.465 121.500 212.785 ;
        RECT 120.915 211.560 121.145 211.850 ;
        RECT 120.915 202.820 121.145 203.110 ;
        RECT 120.960 201.745 121.100 202.820 ;
        RECT 120.900 201.425 121.160 201.745 ;
        RECT 121.300 200.735 121.440 212.465 ;
        RECT 121.580 210.165 121.840 210.485 ;
        RECT 121.980 210.025 122.120 216.160 ;
        RECT 121.920 209.705 122.180 210.025 ;
        RECT 121.935 206.960 122.165 207.250 ;
        RECT 121.580 206.025 121.840 206.345 ;
        RECT 121.595 205.120 121.825 205.410 ;
        RECT 121.640 201.195 121.780 205.120 ;
        RECT 121.980 204.950 122.120 206.960 ;
        RECT 121.935 204.660 122.165 204.950 ;
        RECT 121.640 201.055 122.460 201.195 ;
        RECT 120.960 200.595 121.440 200.735 ;
        RECT 120.960 194.385 121.100 200.595 ;
        RECT 121.920 200.505 122.180 200.825 ;
        RECT 121.255 200.035 121.485 200.325 ;
        RECT 121.300 198.225 121.440 200.035 ;
        RECT 121.595 199.640 121.825 199.930 ;
        RECT 121.640 198.740 121.780 199.640 ;
        RECT 121.935 199.185 122.165 199.475 ;
        RECT 121.595 198.450 121.825 198.740 ;
        RECT 121.255 197.935 121.485 198.225 ;
        RECT 121.300 196.655 121.440 197.935 ;
        RECT 121.255 196.365 121.485 196.655 ;
        RECT 121.640 196.220 121.780 198.450 ;
        RECT 121.595 195.930 121.825 196.220 ;
        RECT 121.980 195.675 122.120 199.185 ;
        RECT 122.320 196.225 122.460 201.055 ;
        RECT 122.260 195.905 122.520 196.225 ;
        RECT 121.300 195.535 122.120 195.675 ;
        RECT 120.900 194.065 121.160 194.385 ;
        RECT 120.915 193.620 121.145 193.910 ;
        RECT 120.960 192.085 121.100 193.620 ;
        RECT 121.300 192.990 121.440 195.535 ;
        RECT 121.920 194.985 122.180 195.305 ;
        RECT 121.580 194.065 121.840 194.385 ;
        RECT 121.255 192.700 121.485 192.990 ;
        RECT 120.900 191.765 121.160 192.085 ;
        RECT 121.640 190.690 121.780 194.065 ;
        RECT 121.595 190.400 121.825 190.690 ;
        RECT 121.595 190.155 121.825 190.230 ;
        RECT 121.980 190.155 122.120 194.985 ;
        RECT 122.600 190.845 122.860 191.165 ;
        RECT 121.595 190.015 122.120 190.155 ;
        RECT 121.595 189.940 121.825 190.015 ;
        RECT 121.580 189.005 121.840 189.325 ;
        RECT 120.900 188.085 121.160 188.405 ;
        RECT 120.960 186.550 121.100 188.085 ;
        RECT 121.255 187.640 121.485 187.930 ;
        RECT 120.915 186.260 121.145 186.550 ;
        RECT 121.300 185.185 121.440 187.640 ;
        RECT 121.640 186.105 121.780 189.005 ;
        RECT 121.920 188.545 122.180 188.865 ;
        RECT 121.920 187.165 122.180 187.485 ;
        RECT 122.600 187.165 122.860 187.485 ;
        RECT 121.980 186.550 122.120 187.165 ;
        RECT 122.260 186.705 122.520 187.025 ;
        RECT 121.935 186.260 122.165 186.550 ;
        RECT 121.580 185.785 121.840 186.105 ;
        RECT 121.240 184.865 121.500 185.185 ;
        RECT 122.320 185.170 122.460 186.705 ;
        RECT 122.275 184.880 122.505 185.170 ;
        RECT 123.000 183.415 123.480 219.295 ;
        RECT 124.640 217.755 124.900 217.845 ;
        RECT 124.360 217.615 124.900 217.755 ;
        RECT 123.975 216.205 124.205 216.495 ;
        RECT 124.020 215.545 124.160 216.205 ;
        RECT 123.960 215.225 124.220 215.545 ;
        RECT 124.360 210.945 124.500 217.615 ;
        RECT 124.640 217.525 124.900 217.615 ;
        RECT 124.995 217.055 125.225 217.345 ;
        RECT 124.655 216.660 124.885 216.950 ;
        RECT 124.700 215.760 124.840 216.660 ;
        RECT 124.655 215.470 124.885 215.760 ;
        RECT 124.700 213.240 124.840 215.470 ;
        RECT 125.040 215.245 125.180 217.055 ;
        RECT 124.995 214.955 125.225 215.245 ;
        RECT 125.040 213.675 125.180 214.955 ;
        RECT 124.995 213.385 125.225 213.675 ;
        RECT 124.655 212.950 124.885 213.240 ;
        RECT 124.300 210.625 124.560 210.945 ;
        RECT 125.335 210.640 125.565 210.930 ;
        RECT 124.360 205.870 124.500 210.625 ;
        RECT 125.380 210.025 125.520 210.640 ;
        RECT 125.320 209.705 125.580 210.025 ;
        RECT 124.315 205.795 124.545 205.870 ;
        RECT 123.680 205.655 124.545 205.795 ;
        RECT 123.680 200.825 123.820 205.655 ;
        RECT 124.315 205.580 124.545 205.655 ;
        RECT 124.995 205.095 125.225 205.385 ;
        RECT 123.960 204.645 124.220 204.965 ;
        RECT 124.655 204.700 124.885 204.990 ;
        RECT 124.020 204.415 124.160 204.645 ;
        RECT 124.315 204.415 124.545 204.535 ;
        RECT 124.020 204.275 124.545 204.415 ;
        RECT 124.315 204.245 124.545 204.275 ;
        RECT 124.700 203.800 124.840 204.700 ;
        RECT 124.655 203.510 124.885 203.800 ;
        RECT 124.700 201.280 124.840 203.510 ;
        RECT 125.040 203.285 125.180 205.095 ;
        RECT 124.995 202.995 125.225 203.285 ;
        RECT 125.040 201.715 125.180 202.995 ;
        RECT 124.995 201.425 125.225 201.715 ;
        RECT 124.655 200.990 124.885 201.280 ;
        RECT 123.620 200.505 123.880 200.825 ;
        RECT 123.635 198.680 123.865 198.970 ;
        RECT 123.680 198.065 123.820 198.680 ;
        RECT 124.655 198.220 124.885 198.510 ;
        RECT 123.620 197.745 123.880 198.065 ;
        RECT 124.700 197.605 124.840 198.220 ;
        RECT 124.640 197.285 124.900 197.605 ;
        RECT 124.980 196.365 125.240 196.685 ;
        RECT 125.335 195.920 125.565 196.210 ;
        RECT 125.380 195.305 125.520 195.920 ;
        RECT 125.320 194.985 125.580 195.305 ;
        RECT 124.300 191.765 124.560 192.085 ;
        RECT 123.620 190.845 123.880 191.165 ;
        RECT 123.680 188.850 123.820 190.845 ;
        RECT 124.640 189.465 124.900 189.785 ;
        RECT 124.300 189.005 124.560 189.325 ;
        RECT 123.635 188.560 123.865 188.850 ;
        RECT 124.360 187.470 124.500 189.005 ;
        RECT 124.315 187.180 124.545 187.470 ;
        RECT 124.300 186.705 124.560 187.025 ;
        RECT 124.300 186.245 124.560 186.565 ;
        RECT 124.315 186.015 124.545 186.090 ;
        RECT 124.700 186.015 124.840 189.465 ;
        RECT 125.320 189.005 125.580 189.325 ;
        RECT 125.380 188.390 125.520 189.005 ;
        RECT 125.335 188.100 125.565 188.390 ;
        RECT 124.315 185.875 124.840 186.015 ;
        RECT 124.315 185.800 124.545 185.875 ;
        RECT 125.720 183.415 126.200 219.295 ;
        RECT 128.040 217.985 128.300 218.305 ;
        RECT 126.680 217.525 126.940 217.845 ;
        RECT 127.360 217.525 127.620 217.845 ;
        RECT 126.340 215.225 126.600 215.545 ;
        RECT 126.740 211.315 126.880 217.525 ;
        RECT 127.420 216.450 127.560 217.525 ;
        RECT 128.100 217.370 128.240 217.985 ;
        RECT 128.055 217.080 128.285 217.370 ;
        RECT 127.375 216.160 127.605 216.450 ;
        RECT 128.055 213.400 128.285 213.690 ;
        RECT 127.035 212.940 127.265 213.230 ;
        RECT 127.080 212.785 127.220 212.940 ;
        RECT 128.100 212.785 128.240 213.400 ;
        RECT 127.020 212.465 127.280 212.785 ;
        RECT 128.040 212.465 128.300 212.785 ;
        RECT 127.020 212.005 127.280 212.325 ;
        RECT 127.035 211.315 127.265 211.390 ;
        RECT 126.740 211.175 127.265 211.315 ;
        RECT 127.035 211.100 127.265 211.175 ;
        RECT 126.695 210.615 126.925 210.905 ;
        RECT 126.740 208.805 126.880 210.615 ;
        RECT 127.035 210.220 127.265 210.510 ;
        RECT 127.080 209.320 127.220 210.220 ;
        RECT 127.715 209.765 127.945 210.055 ;
        RECT 127.035 209.030 127.265 209.320 ;
        RECT 126.695 208.515 126.925 208.805 ;
        RECT 126.740 207.235 126.880 208.515 ;
        RECT 126.695 206.945 126.925 207.235 ;
        RECT 127.080 206.800 127.220 209.030 ;
        RECT 127.035 206.510 127.265 206.800 ;
        RECT 127.760 206.345 127.900 209.765 ;
        RECT 127.700 206.025 127.960 206.345 ;
        RECT 127.760 204.965 127.900 206.025 ;
        RECT 126.680 204.645 126.940 204.965 ;
        RECT 127.700 204.645 127.960 204.965 ;
        RECT 126.740 204.030 126.880 204.645 ;
        RECT 128.040 204.185 128.300 204.505 ;
        RECT 126.695 203.740 126.925 204.030 ;
        RECT 127.375 201.900 127.605 202.190 ;
        RECT 127.035 201.655 127.265 201.730 ;
        RECT 126.740 201.515 127.265 201.655 ;
        RECT 126.740 196.225 126.880 201.515 ;
        RECT 127.035 201.440 127.265 201.515 ;
        RECT 127.035 200.520 127.265 200.810 ;
        RECT 127.080 198.525 127.220 200.520 ;
        RECT 127.420 199.890 127.560 201.900 ;
        RECT 127.375 199.600 127.605 199.890 ;
        RECT 127.020 198.205 127.280 198.525 ;
        RECT 127.020 197.745 127.280 198.065 ;
        RECT 127.080 197.130 127.220 197.745 ;
        RECT 128.100 197.605 128.240 204.185 ;
        RECT 128.040 197.285 128.300 197.605 ;
        RECT 127.035 196.840 127.265 197.130 ;
        RECT 126.680 195.905 126.940 196.225 ;
        RECT 126.740 190.230 126.880 195.905 ;
        RECT 127.360 193.605 127.620 193.925 ;
        RECT 127.420 192.530 127.560 193.605 ;
        RECT 127.375 192.240 127.605 192.530 ;
        RECT 127.375 191.995 127.605 192.070 ;
        RECT 127.375 191.855 127.900 191.995 ;
        RECT 127.375 191.780 127.605 191.855 ;
        RECT 127.360 191.305 127.620 191.625 ;
        RECT 127.035 190.860 127.265 191.150 ;
        RECT 126.695 189.940 126.925 190.230 ;
        RECT 127.080 187.485 127.220 190.860 ;
        RECT 127.760 189.785 127.900 191.855 ;
        RECT 127.700 189.465 127.960 189.785 ;
        RECT 127.375 188.560 127.605 188.850 ;
        RECT 127.420 188.405 127.560 188.560 ;
        RECT 127.360 188.085 127.620 188.405 ;
        RECT 127.360 187.625 127.620 187.945 ;
        RECT 128.040 187.625 128.300 187.945 ;
        RECT 127.020 187.165 127.280 187.485 ;
        RECT 127.375 186.260 127.605 186.550 ;
        RECT 127.420 186.105 127.560 186.260 ;
        RECT 127.360 185.785 127.620 186.105 ;
        RECT 128.100 185.630 128.240 187.625 ;
        RECT 128.055 185.340 128.285 185.630 ;
        RECT 128.440 183.415 128.920 219.295 ;
        RECT 130.080 217.525 130.340 217.845 ;
        RECT 130.140 216.450 130.280 217.525 ;
        RECT 130.095 216.160 130.325 216.450 ;
        RECT 130.760 212.925 131.020 213.245 ;
        RECT 129.060 212.465 129.320 212.785 ;
        RECT 129.740 209.705 130.000 210.025 ;
        RECT 129.755 205.795 129.985 205.870 ;
        RECT 129.460 205.655 129.985 205.795 ;
        RECT 129.460 200.350 129.600 205.655 ;
        RECT 129.755 205.580 129.985 205.655 ;
        RECT 129.755 204.875 129.985 204.950 ;
        RECT 129.755 204.735 130.280 204.875 ;
        RECT 129.755 204.660 129.985 204.735 ;
        RECT 129.740 204.185 130.000 204.505 ;
        RECT 130.140 203.495 130.280 204.735 ;
        RECT 130.760 204.645 131.020 204.965 ;
        RECT 130.760 204.185 131.020 204.505 ;
        RECT 130.435 203.495 130.665 203.570 ;
        RECT 130.140 203.355 130.665 203.495 ;
        RECT 130.435 203.280 130.665 203.355 ;
        RECT 130.095 202.820 130.325 203.110 ;
        RECT 129.755 201.900 129.985 202.190 ;
        RECT 129.800 201.745 129.940 201.900 ;
        RECT 129.740 201.425 130.000 201.745 ;
        RECT 129.740 200.505 130.000 200.825 ;
        RECT 129.415 200.060 129.645 200.350 ;
        RECT 130.140 197.515 130.280 202.820 ;
        RECT 130.480 200.365 130.620 203.280 ;
        RECT 130.820 202.650 130.960 204.185 ;
        RECT 130.775 202.360 131.005 202.650 ;
        RECT 130.420 200.045 130.680 200.365 ;
        RECT 130.140 197.375 130.620 197.515 ;
        RECT 130.080 196.825 130.340 197.145 ;
        RECT 130.480 196.225 130.620 197.375 ;
        RECT 130.420 195.905 130.680 196.225 ;
        RECT 129.075 195.000 129.305 195.290 ;
        RECT 129.120 194.385 129.260 195.000 ;
        RECT 129.060 194.065 129.320 194.385 ;
        RECT 129.755 194.295 129.985 194.370 ;
        RECT 129.755 194.155 130.280 194.295 ;
        RECT 129.755 194.080 129.985 194.155 ;
        RECT 129.755 193.160 129.985 193.450 ;
        RECT 129.415 191.780 129.645 192.070 ;
        RECT 129.060 191.305 129.320 191.625 ;
        RECT 129.120 191.150 129.260 191.305 ;
        RECT 129.075 190.860 129.305 191.150 ;
        RECT 129.460 189.785 129.600 191.780 ;
        RECT 129.800 191.610 129.940 193.160 ;
        RECT 129.755 191.320 129.985 191.610 ;
        RECT 129.800 191.165 129.940 191.320 ;
        RECT 129.740 190.845 130.000 191.165 ;
        RECT 129.755 190.615 129.985 190.690 ;
        RECT 130.140 190.615 130.280 194.155 ;
        RECT 130.760 193.605 131.020 193.925 ;
        RECT 129.755 190.475 130.280 190.615 ;
        RECT 129.755 190.400 129.985 190.475 ;
        RECT 129.740 189.925 130.000 190.245 ;
        RECT 129.400 189.465 129.660 189.785 ;
        RECT 129.075 189.235 129.305 189.310 ;
        RECT 129.075 189.095 129.600 189.235 ;
        RECT 129.075 189.020 129.305 189.095 ;
        RECT 129.460 188.775 129.600 189.095 ;
        RECT 129.755 188.775 129.985 188.850 ;
        RECT 129.460 188.635 129.985 188.775 ;
        RECT 129.460 187.025 129.600 188.635 ;
        RECT 129.755 188.560 129.985 188.635 ;
        RECT 129.740 187.625 130.000 187.945 ;
        RECT 130.140 187.855 130.280 190.475 ;
        RECT 130.420 187.855 130.680 187.945 ;
        RECT 130.140 187.715 130.680 187.855 ;
        RECT 130.420 187.625 130.680 187.715 ;
        RECT 129.740 187.165 130.000 187.485 ;
        RECT 129.400 186.705 129.660 187.025 ;
        RECT 129.800 186.550 129.940 187.165 ;
        RECT 129.755 186.260 129.985 186.550 ;
        RECT 130.760 186.245 131.020 186.565 ;
        RECT 130.820 185.630 130.960 186.245 ;
        RECT 130.775 185.340 131.005 185.630 ;
        RECT 131.160 183.415 131.640 219.295 ;
        RECT 131.780 217.525 132.040 217.845 ;
        RECT 133.140 217.525 133.400 217.845 ;
        RECT 132.475 215.230 132.705 215.520 ;
        RECT 132.135 214.795 132.365 215.085 ;
        RECT 132.180 213.515 132.320 214.795 ;
        RECT 132.135 213.225 132.365 213.515 ;
        RECT 132.180 211.415 132.320 213.225 ;
        RECT 132.520 213.000 132.660 215.230 ;
        RECT 132.475 212.710 132.705 213.000 ;
        RECT 132.520 211.810 132.660 212.710 ;
        RECT 133.200 212.265 133.340 217.525 ;
        RECT 133.155 211.975 133.385 212.265 ;
        RECT 132.475 211.520 132.705 211.810 ;
        RECT 132.135 211.125 132.365 211.415 ;
        RECT 132.800 210.625 133.060 210.945 ;
        RECT 133.140 206.945 133.400 207.265 ;
        RECT 131.780 200.965 132.040 201.285 ;
        RECT 131.840 200.810 131.980 200.965 ;
        RECT 131.795 200.520 132.025 200.810 ;
        RECT 132.460 200.505 132.720 200.825 ;
        RECT 131.780 195.905 132.040 196.225 ;
        RECT 131.840 192.990 131.980 195.905 ;
        RECT 132.520 195.290 132.660 200.505 ;
        RECT 133.480 197.745 133.740 198.065 ;
        RECT 133.480 195.445 133.740 195.765 ;
        RECT 132.475 195.000 132.705 195.290 ;
        RECT 131.795 192.700 132.025 192.990 ;
        RECT 132.800 192.685 133.060 193.005 ;
        RECT 132.800 191.765 133.060 192.085 ;
        RECT 133.540 191.150 133.680 195.445 ;
        RECT 133.495 190.860 133.725 191.150 ;
        RECT 131.780 189.465 132.040 189.785 ;
        RECT 131.840 186.550 131.980 189.465 ;
        RECT 132.800 187.395 133.060 187.485 ;
        RECT 132.800 187.255 133.340 187.395 ;
        RECT 132.800 187.165 133.060 187.255 ;
        RECT 131.795 186.260 132.025 186.550 ;
        RECT 132.815 186.260 133.045 186.550 ;
        RECT 132.860 186.105 133.000 186.260 ;
        RECT 132.800 185.785 133.060 186.105 ;
        RECT 133.200 186.015 133.340 187.255 ;
        RECT 133.495 186.015 133.725 186.090 ;
        RECT 133.200 185.875 133.725 186.015 ;
        RECT 133.495 185.800 133.725 185.875 ;
        RECT 132.800 184.865 133.060 185.185 ;
        RECT 133.880 183.415 134.360 219.295 ;
        RECT 134.500 217.525 134.760 217.845 ;
        RECT 134.515 215.700 134.745 215.990 ;
        RECT 134.560 213.245 134.700 215.700 ;
        RECT 135.520 215.225 135.780 215.545 ;
        RECT 135.535 214.320 135.765 214.610 ;
        RECT 135.195 213.400 135.425 213.690 ;
        RECT 135.580 213.615 135.720 214.320 ;
        RECT 135.580 213.475 136.400 213.615 ;
        RECT 134.500 212.925 134.760 213.245 ;
        RECT 134.900 212.355 135.040 212.760 ;
        RECT 134.855 212.325 135.085 212.355 ;
        RECT 134.840 212.005 135.100 212.325 ;
        RECT 134.900 204.875 135.040 212.005 ;
        RECT 135.240 210.945 135.380 213.400 ;
        RECT 135.875 212.915 136.105 213.205 ;
        RECT 135.535 212.520 135.765 212.810 ;
        RECT 135.580 211.620 135.720 212.520 ;
        RECT 135.535 211.330 135.765 211.620 ;
        RECT 135.180 210.625 135.440 210.945 ;
        RECT 135.240 208.185 135.380 210.625 ;
        RECT 135.580 209.100 135.720 211.330 ;
        RECT 135.920 211.105 136.060 212.915 ;
        RECT 135.875 210.815 136.105 211.105 ;
        RECT 135.920 209.535 136.060 210.815 ;
        RECT 135.875 209.245 136.105 209.535 ;
        RECT 135.535 208.810 135.765 209.100 ;
        RECT 135.180 207.865 135.440 208.185 ;
        RECT 135.875 206.715 136.105 206.790 ;
        RECT 134.560 204.735 135.040 204.875 ;
        RECT 135.240 206.575 136.105 206.715 ;
        RECT 134.560 198.525 134.700 204.735 ;
        RECT 134.855 204.245 135.085 204.535 ;
        RECT 134.500 198.205 134.760 198.525 ;
        RECT 134.560 197.590 134.700 198.205 ;
        RECT 134.900 198.065 135.040 204.245 ;
        RECT 134.840 197.745 135.100 198.065 ;
        RECT 135.240 197.605 135.380 206.575 ;
        RECT 135.875 206.500 136.105 206.575 ;
        RECT 135.520 205.565 135.780 205.885 ;
        RECT 135.875 205.095 136.105 205.385 ;
        RECT 135.535 204.700 135.765 204.990 ;
        RECT 135.580 203.800 135.720 204.700 ;
        RECT 135.535 203.510 135.765 203.800 ;
        RECT 135.580 201.280 135.720 203.510 ;
        RECT 135.920 203.285 136.060 205.095 ;
        RECT 136.260 204.965 136.400 213.475 ;
        RECT 136.200 204.645 136.460 204.965 ;
        RECT 135.875 202.995 136.105 203.285 ;
        RECT 135.920 201.715 136.060 202.995 ;
        RECT 135.875 201.425 136.105 201.715 ;
        RECT 135.535 200.990 135.765 201.280 ;
        RECT 136.215 198.680 136.445 198.970 ;
        RECT 136.260 198.525 136.400 198.680 ;
        RECT 136.200 198.205 136.460 198.525 ;
        RECT 134.515 197.300 134.745 197.590 ;
        RECT 135.180 197.285 135.440 197.605 ;
        RECT 134.840 196.595 135.100 196.685 ;
        RECT 135.240 196.595 135.380 197.285 ;
        RECT 135.860 196.825 136.120 197.145 ;
        RECT 134.840 196.455 135.380 196.595 ;
        RECT 134.840 196.365 135.100 196.455 ;
        RECT 134.900 195.290 135.040 196.365 ;
        RECT 134.855 195.000 135.085 195.290 ;
        RECT 134.515 193.620 134.745 193.910 ;
        RECT 134.560 193.005 134.700 193.620 ;
        RECT 134.500 192.685 134.760 193.005 ;
        RECT 135.195 192.915 135.425 192.990 ;
        RECT 134.900 192.775 135.425 192.915 ;
        RECT 134.900 192.455 135.040 192.775 ;
        RECT 135.195 192.700 135.425 192.775 ;
        RECT 134.560 192.315 135.040 192.455 ;
        RECT 135.535 192.455 135.765 192.530 ;
        RECT 135.535 192.315 136.060 192.455 ;
        RECT 134.560 187.855 134.700 192.315 ;
        RECT 135.535 192.240 135.765 192.315 ;
        RECT 135.535 191.780 135.765 192.070 ;
        RECT 135.195 191.535 135.425 191.610 ;
        RECT 134.900 191.395 135.425 191.535 ;
        RECT 134.900 190.230 135.040 191.395 ;
        RECT 135.195 191.320 135.425 191.395 ;
        RECT 135.180 190.845 135.440 191.165 ;
        RECT 135.240 190.690 135.380 190.845 ;
        RECT 135.195 190.400 135.425 190.690 ;
        RECT 134.855 189.940 135.085 190.230 ;
        RECT 135.195 189.480 135.425 189.770 ;
        RECT 135.240 188.405 135.380 189.480 ;
        RECT 135.580 189.325 135.720 191.780 ;
        RECT 135.920 190.245 136.060 192.315 ;
        RECT 135.860 189.925 136.120 190.245 ;
        RECT 135.520 189.005 135.780 189.325 ;
        RECT 135.180 188.085 135.440 188.405 ;
        RECT 135.180 187.855 135.440 187.945 ;
        RECT 134.560 187.715 135.440 187.855 ;
        RECT 135.180 187.625 135.440 187.715 ;
        RECT 135.180 186.245 135.440 186.565 ;
        RECT 135.180 185.785 135.440 186.105 ;
        RECT 135.240 185.630 135.380 185.785 ;
        RECT 135.920 185.645 136.060 189.925 ;
        RECT 136.215 188.560 136.445 188.850 ;
        RECT 136.260 187.025 136.400 188.560 ;
        RECT 136.200 186.705 136.460 187.025 ;
        RECT 135.195 185.340 135.425 185.630 ;
        RECT 135.860 185.325 136.120 185.645 ;
        RECT 136.600 183.415 137.080 219.295 ;
        RECT 138.920 217.985 139.180 218.305 ;
        RECT 138.980 217.370 139.120 217.985 ;
        RECT 138.935 217.080 139.165 217.370 ;
        RECT 138.255 216.160 138.485 216.450 ;
        RECT 137.560 215.225 137.820 215.545 ;
        RECT 137.620 213.615 137.760 215.225 ;
        RECT 137.915 213.615 138.145 213.690 ;
        RECT 137.620 213.475 138.145 213.615 ;
        RECT 137.235 200.980 137.465 201.270 ;
        RECT 137.280 200.825 137.420 200.980 ;
        RECT 137.220 200.505 137.480 200.825 ;
        RECT 137.620 195.765 137.760 213.475 ;
        RECT 137.915 213.400 138.145 213.475 ;
        RECT 137.915 212.480 138.145 212.770 ;
        RECT 137.960 212.325 138.100 212.480 ;
        RECT 137.900 212.005 138.160 212.325 ;
        RECT 138.300 210.945 138.440 216.160 ;
        RECT 138.920 215.685 139.180 216.005 ;
        RECT 138.935 213.860 139.165 214.150 ;
        RECT 138.240 210.625 138.500 210.945 ;
        RECT 138.980 210.485 139.120 213.860 ;
        RECT 138.920 210.165 139.180 210.485 ;
        RECT 138.920 207.865 139.180 208.185 ;
        RECT 138.980 205.885 139.120 207.865 ;
        RECT 138.920 205.565 139.180 205.885 ;
        RECT 138.920 204.645 139.180 204.965 ;
        RECT 138.255 201.440 138.485 201.730 ;
        RECT 138.300 201.285 138.440 201.440 ;
        RECT 138.980 201.285 139.120 204.645 ;
        RECT 138.240 200.965 138.500 201.285 ;
        RECT 138.920 200.965 139.180 201.285 ;
        RECT 137.915 197.760 138.145 198.050 ;
        RECT 137.960 197.605 138.100 197.760 ;
        RECT 137.900 197.285 138.160 197.605 ;
        RECT 138.580 195.905 138.840 196.225 ;
        RECT 137.560 195.445 137.820 195.765 ;
        RECT 137.915 195.000 138.145 195.290 ;
        RECT 137.235 194.755 137.465 194.830 ;
        RECT 137.235 194.615 137.760 194.755 ;
        RECT 137.235 194.540 137.465 194.615 ;
        RECT 137.220 193.605 137.480 193.925 ;
        RECT 137.620 191.165 137.760 194.615 ;
        RECT 137.960 191.995 138.100 195.000 ;
        RECT 138.255 194.755 138.485 194.830 ;
        RECT 138.255 194.615 139.120 194.755 ;
        RECT 138.255 194.540 138.485 194.615 ;
        RECT 138.595 192.700 138.825 192.990 ;
        RECT 138.240 191.995 138.500 192.085 ;
        RECT 137.960 191.855 138.500 191.995 ;
        RECT 138.240 191.765 138.500 191.855 ;
        RECT 138.640 191.625 138.780 192.700 ;
        RECT 138.580 191.305 138.840 191.625 ;
        RECT 137.560 190.845 137.820 191.165 ;
        RECT 138.580 190.845 138.840 191.165 ;
        RECT 138.255 190.615 138.485 190.690 ;
        RECT 137.960 190.475 138.485 190.615 ;
        RECT 137.960 189.310 138.100 190.475 ;
        RECT 138.255 190.400 138.485 190.475 ;
        RECT 138.255 189.695 138.485 189.770 ;
        RECT 138.640 189.695 138.780 190.845 ;
        RECT 138.255 189.555 138.780 189.695 ;
        RECT 138.255 189.480 138.485 189.555 ;
        RECT 137.915 189.020 138.145 189.310 ;
        RECT 138.240 188.085 138.500 188.405 ;
        RECT 138.240 186.705 138.500 187.025 ;
        RECT 138.255 185.800 138.485 186.090 ;
        RECT 138.640 186.015 138.780 189.555 ;
        RECT 138.980 188.405 139.120 194.615 ;
        RECT 138.920 188.085 139.180 188.405 ;
        RECT 138.920 186.015 139.180 186.105 ;
        RECT 138.640 185.875 139.180 186.015 ;
        RECT 138.300 185.645 138.440 185.800 ;
        RECT 138.920 185.785 139.180 185.875 ;
        RECT 138.240 185.325 138.500 185.645 ;
        RECT 139.320 183.415 139.800 219.295 ;
        RECT 140.635 217.540 140.865 217.830 ;
        RECT 140.295 216.205 140.525 216.495 ;
        RECT 140.340 216.005 140.480 216.205 ;
        RECT 140.280 215.685 140.540 216.005 ;
        RECT 139.940 210.855 140.200 210.945 ;
        RECT 139.940 210.715 140.480 210.855 ;
        RECT 139.940 210.625 140.200 210.715 ;
        RECT 139.940 210.165 140.200 210.485 ;
        RECT 140.340 207.635 140.480 210.715 ;
        RECT 140.680 208.185 140.820 217.540 ;
        RECT 141.315 217.055 141.545 217.345 ;
        RECT 140.975 216.660 141.205 216.950 ;
        RECT 141.020 215.760 141.160 216.660 ;
        RECT 140.975 215.470 141.205 215.760 ;
        RECT 141.020 213.240 141.160 215.470 ;
        RECT 141.360 215.245 141.500 217.055 ;
        RECT 141.315 214.955 141.545 215.245 ;
        RECT 141.360 213.675 141.500 214.955 ;
        RECT 141.315 213.385 141.545 213.675 ;
        RECT 140.975 212.950 141.205 213.240 ;
        RECT 140.620 207.865 140.880 208.185 ;
        RECT 140.635 207.635 140.865 207.710 ;
        RECT 140.340 207.495 140.865 207.635 ;
        RECT 140.635 207.420 140.865 207.495 ;
        RECT 141.640 205.565 141.900 205.885 ;
        RECT 140.635 203.740 140.865 204.030 ;
        RECT 140.295 203.280 140.525 203.570 ;
        RECT 139.940 201.425 140.200 201.745 ;
        RECT 140.000 199.430 140.140 201.425 ;
        RECT 139.955 199.140 140.185 199.430 ;
        RECT 140.340 195.765 140.480 203.280 ;
        RECT 140.680 201.745 140.820 203.740 ;
        RECT 140.975 202.575 141.205 202.650 ;
        RECT 140.975 202.435 141.500 202.575 ;
        RECT 140.975 202.360 141.205 202.435 ;
        RECT 140.620 201.425 140.880 201.745 ;
        RECT 140.620 200.965 140.880 201.285 ;
        RECT 140.620 200.045 140.880 200.365 ;
        RECT 140.680 198.525 140.820 200.045 ;
        RECT 140.620 198.205 140.880 198.525 ;
        RECT 140.620 197.745 140.880 198.065 ;
        RECT 140.680 197.145 140.820 197.745 ;
        RECT 140.960 197.285 141.220 197.605 ;
        RECT 141.360 197.515 141.500 202.435 ;
        RECT 141.640 200.505 141.900 200.825 ;
        RECT 141.700 198.510 141.840 200.505 ;
        RECT 141.655 198.220 141.885 198.510 ;
        RECT 141.360 197.375 141.840 197.515 ;
        RECT 140.620 196.825 140.880 197.145 ;
        RECT 141.315 196.815 141.545 197.105 ;
        RECT 140.975 196.420 141.205 196.710 ;
        RECT 140.635 195.965 140.865 196.255 ;
        RECT 140.280 195.445 140.540 195.765 ;
        RECT 140.680 194.845 140.820 195.965 ;
        RECT 141.020 195.520 141.160 196.420 ;
        RECT 140.975 195.230 141.205 195.520 ;
        RECT 140.620 194.525 140.880 194.845 ;
        RECT 141.020 193.000 141.160 195.230 ;
        RECT 141.360 195.005 141.500 196.815 ;
        RECT 141.700 195.765 141.840 197.375 ;
        RECT 141.640 195.445 141.900 195.765 ;
        RECT 141.315 194.715 141.545 195.005 ;
        RECT 141.360 193.435 141.500 194.715 ;
        RECT 141.315 193.145 141.545 193.435 ;
        RECT 140.975 192.710 141.205 193.000 ;
        RECT 141.700 192.455 141.840 195.445 ;
        RECT 140.680 192.315 141.840 192.455 ;
        RECT 140.680 189.770 140.820 192.315 ;
        RECT 141.640 190.385 141.900 190.705 ;
        RECT 140.635 189.480 140.865 189.770 ;
        RECT 140.620 188.545 140.880 188.865 ;
        RECT 141.640 187.625 141.900 187.945 ;
        RECT 140.620 187.165 140.880 187.485 ;
        RECT 139.940 186.245 140.200 186.565 ;
        RECT 139.940 185.785 140.200 186.105 ;
        RECT 140.620 184.865 140.880 185.185 ;
        RECT 142.040 183.415 142.520 219.295 ;
        RECT 144.360 213.385 144.620 213.705 ;
        RECT 143.355 211.090 143.585 211.380 ;
        RECT 143.015 210.655 143.245 210.945 ;
        RECT 143.060 209.375 143.200 210.655 ;
        RECT 143.015 209.085 143.245 209.375 ;
        RECT 142.660 207.865 142.920 208.185 ;
        RECT 142.720 206.255 142.860 207.865 ;
        RECT 143.060 207.275 143.200 209.085 ;
        RECT 143.400 208.860 143.540 211.090 ;
        RECT 143.355 208.570 143.585 208.860 ;
        RECT 144.360 208.785 144.620 209.105 ;
        RECT 143.400 207.670 143.540 208.570 ;
        RECT 143.695 207.780 143.925 208.070 ;
        RECT 143.355 207.380 143.585 207.670 ;
        RECT 143.015 206.985 143.245 207.275 ;
        RECT 143.355 206.500 143.585 206.790 ;
        RECT 143.400 206.330 143.540 206.500 ;
        RECT 143.355 206.255 143.585 206.330 ;
        RECT 142.720 206.115 143.585 206.255 ;
        RECT 142.720 197.605 142.860 206.115 ;
        RECT 143.355 206.040 143.585 206.115 ;
        RECT 143.740 205.885 143.880 207.780 ;
        RECT 144.020 206.485 144.280 206.805 ;
        RECT 143.015 205.555 143.245 205.845 ;
        RECT 143.680 205.565 143.940 205.885 ;
        RECT 143.060 203.745 143.200 205.555 ;
        RECT 143.355 205.160 143.585 205.450 ;
        RECT 143.400 204.260 143.540 205.160 ;
        RECT 144.080 205.105 144.220 206.485 ;
        RECT 144.035 204.815 144.265 205.105 ;
        RECT 143.355 203.970 143.585 204.260 ;
        RECT 143.015 203.455 143.245 203.745 ;
        RECT 143.060 202.175 143.200 203.455 ;
        RECT 143.015 201.885 143.245 202.175 ;
        RECT 143.400 201.740 143.540 203.970 ;
        RECT 144.420 203.955 144.560 208.785 ;
        RECT 144.080 203.815 144.560 203.955 ;
        RECT 143.355 201.450 143.585 201.740 ;
        RECT 143.000 200.965 143.260 201.285 ;
        RECT 142.660 197.285 142.920 197.605 ;
        RECT 143.060 195.750 143.200 200.965 ;
        RECT 143.340 200.045 143.600 200.365 ;
        RECT 143.400 196.595 143.540 200.045 ;
        RECT 144.080 198.970 144.220 203.815 ;
        RECT 144.375 199.140 144.605 199.430 ;
        RECT 144.035 198.680 144.265 198.970 ;
        RECT 144.420 198.525 144.560 199.140 ;
        RECT 144.360 198.205 144.620 198.525 ;
        RECT 144.020 197.745 144.280 198.065 ;
        RECT 143.680 196.825 143.940 197.145 ;
        RECT 143.695 196.595 143.925 196.670 ;
        RECT 143.400 196.455 143.925 196.595 ;
        RECT 143.695 196.380 143.925 196.455 ;
        RECT 143.340 195.905 143.600 196.225 ;
        RECT 143.015 195.460 143.245 195.750 ;
        RECT 142.660 194.525 142.920 194.845 ;
        RECT 142.720 192.990 142.860 194.525 ;
        RECT 143.015 194.080 143.245 194.370 ;
        RECT 142.675 192.700 142.905 192.990 ;
        RECT 143.060 191.610 143.200 194.080 ;
        RECT 143.400 193.835 143.540 195.905 ;
        RECT 143.680 195.445 143.940 195.765 ;
        RECT 143.740 194.830 143.880 195.445 ;
        RECT 143.695 194.540 143.925 194.830 ;
        RECT 143.680 193.835 143.940 193.925 ;
        RECT 143.400 193.695 143.940 193.835 ;
        RECT 143.680 193.605 143.940 193.695 ;
        RECT 143.740 192.070 143.880 193.605 ;
        RECT 143.695 191.780 143.925 192.070 ;
        RECT 143.015 191.320 143.245 191.610 ;
        RECT 143.680 190.845 143.940 191.165 ;
        RECT 143.000 190.385 143.260 190.705 ;
        RECT 143.695 190.400 143.925 190.690 ;
        RECT 143.060 189.695 143.200 190.385 ;
        RECT 143.355 189.695 143.585 189.770 ;
        RECT 143.060 189.555 143.585 189.695 ;
        RECT 143.355 189.480 143.585 189.555 ;
        RECT 142.660 188.545 142.920 188.865 ;
        RECT 142.720 186.550 142.860 188.545 ;
        RECT 143.740 187.945 143.880 190.400 ;
        RECT 143.680 187.625 143.940 187.945 ;
        RECT 143.000 187.165 143.260 187.485 ;
        RECT 142.675 186.260 142.905 186.550 ;
        RECT 143.060 186.090 143.200 187.165 ;
        RECT 143.015 185.800 143.245 186.090 ;
        RECT 143.680 184.865 143.940 185.185 ;
        RECT 144.760 183.415 145.240 219.295 ;
        RECT 146.060 213.385 146.320 213.705 ;
        RECT 146.120 211.390 146.260 213.385 ;
        RECT 146.075 211.315 146.305 211.390 ;
        RECT 146.075 211.175 146.600 211.315 ;
        RECT 146.075 211.100 146.305 211.175 ;
        RECT 146.060 208.785 146.320 209.105 ;
        RECT 146.060 208.325 146.320 208.645 ;
        RECT 146.075 207.420 146.305 207.710 ;
        RECT 145.380 206.485 145.640 206.805 ;
        RECT 145.380 201.425 145.640 201.745 ;
        RECT 146.120 199.355 146.260 207.420 ;
        RECT 146.460 204.950 146.600 211.175 ;
        RECT 147.095 210.180 147.325 210.470 ;
        RECT 146.755 207.880 146.985 208.170 ;
        RECT 146.415 204.660 146.645 204.950 ;
        RECT 146.800 200.825 146.940 207.880 ;
        RECT 147.140 205.425 147.280 210.180 ;
        RECT 147.080 205.105 147.340 205.425 ;
        RECT 146.740 200.505 147.000 200.825 ;
        RECT 147.095 199.600 147.325 199.890 ;
        RECT 146.120 199.215 146.940 199.355 ;
        RECT 146.075 198.680 146.305 198.970 ;
        RECT 146.120 198.525 146.260 198.680 ;
        RECT 146.060 198.205 146.320 198.525 ;
        RECT 145.380 197.745 145.640 198.065 ;
        RECT 145.440 195.290 145.580 197.745 ;
        RECT 146.060 195.445 146.320 195.765 ;
        RECT 145.395 195.000 145.625 195.290 ;
        RECT 146.120 194.830 146.260 195.445 ;
        RECT 146.075 194.540 146.305 194.830 ;
        RECT 146.800 193.925 146.940 199.215 ;
        RECT 147.140 198.985 147.280 199.600 ;
        RECT 147.080 198.665 147.340 198.985 ;
        RECT 146.740 193.605 147.000 193.925 ;
        RECT 147.080 192.225 147.340 192.545 ;
        RECT 145.380 191.765 145.640 192.085 ;
        RECT 145.440 188.850 145.580 191.765 ;
        RECT 147.140 191.610 147.280 192.225 ;
        RECT 147.095 191.320 147.325 191.610 ;
        RECT 146.060 190.385 146.320 190.705 ;
        RECT 145.395 188.560 145.625 188.850 ;
        RECT 145.380 188.085 145.640 188.405 ;
        RECT 145.440 187.470 145.580 188.085 ;
        RECT 146.060 187.625 146.320 187.945 ;
        RECT 145.395 187.180 145.625 187.470 ;
        RECT 146.060 186.245 146.320 186.565 ;
        RECT 145.395 185.800 145.625 186.090 ;
        RECT 145.440 185.645 145.580 185.800 ;
        RECT 145.380 185.325 145.640 185.645 ;
        RECT 146.060 184.865 146.320 185.185 ;
        RECT 147.480 183.415 147.960 219.295 ;
        RECT 148.200 201.290 148.340 219.570 ;
        RECT 148.110 200.960 148.440 201.290 ;
        RECT 148.720 198.955 148.860 220.050 ;
        RECT 148.630 198.695 148.950 198.955 ;
        RECT 149.210 198.060 149.350 220.770 ;
        RECT 149.770 205.430 149.910 221.830 ;
        RECT 149.680 205.100 150.000 205.430 ;
        RECT 148.670 197.920 149.350 198.060 ;
        RECT 148.670 192.550 148.810 197.920 ;
        RECT 148.570 192.220 148.900 192.550 ;
        RECT 22.205 181.880 22.495 181.925 ;
        RECT 22.650 181.880 22.970 181.940 ;
        RECT 22.205 181.740 22.970 181.880 ;
        RECT 22.205 181.695 22.495 181.740 ;
        RECT 22.650 181.680 22.970 181.740 ;
        RECT 31.850 181.880 32.170 181.940 ;
        RECT 34.150 181.880 34.470 181.940 ;
        RECT 35.530 181.880 35.850 181.940 ;
        RECT 31.850 181.740 32.540 181.880 ;
        RECT 31.850 181.680 32.170 181.740 ;
        RECT 24.030 181.540 24.350 181.600 ;
        RECT 30.470 181.540 30.790 181.600 ;
        RECT 32.400 181.585 32.540 181.740 ;
        RECT 34.150 181.740 35.850 181.880 ;
        RECT 34.150 181.680 34.470 181.740 ;
        RECT 35.530 181.680 35.850 181.740 ;
        RECT 43.365 181.880 43.655 181.925 ;
        RECT 49.345 181.880 49.635 181.925 ;
        RECT 43.365 181.740 49.635 181.880 ;
        RECT 43.365 181.695 43.655 181.740 ;
        RECT 49.345 181.695 49.635 181.740 ;
        RECT 50.710 181.680 51.030 181.940 ;
        RECT 52.565 181.880 52.855 181.925 ;
        RECT 53.470 181.880 53.790 181.940 ;
        RECT 52.565 181.740 53.790 181.880 ;
        RECT 52.565 181.695 52.855 181.740 ;
        RECT 53.470 181.680 53.790 181.740 ;
        RECT 57.610 181.680 57.930 181.940 ;
        RECT 58.990 181.880 59.310 181.940 ;
        RECT 64.525 181.880 64.815 181.925 ;
        RECT 65.430 181.880 65.750 181.940 ;
        RECT 58.990 181.740 63.820 181.880 ;
        RECT 58.990 181.680 59.310 181.740 ;
        RECT 31.405 181.540 31.695 181.585 ;
        RECT 24.030 181.400 31.695 181.540 ;
        RECT 24.030 181.340 24.350 181.400 ;
        RECT 30.470 181.340 30.790 181.400 ;
        RECT 31.405 181.355 31.695 181.400 ;
        RECT 32.325 181.540 32.615 181.585 ;
        RECT 44.285 181.540 44.575 181.585 ;
        RECT 49.930 181.540 50.220 181.585 ;
        RECT 32.325 181.400 36.680 181.540 ;
        RECT 32.325 181.355 32.615 181.400 ;
        RECT 36.540 181.260 36.680 181.400 ;
        RECT 44.285 181.400 50.220 181.540 ;
        RECT 50.800 181.540 50.940 181.680 ;
        RECT 59.450 181.540 59.770 181.600 ;
        RECT 63.130 181.540 63.450 181.600 ;
        RECT 50.800 181.400 56.000 181.540 ;
        RECT 44.285 181.355 44.575 181.400 ;
        RECT 49.930 181.355 50.220 181.400 ;
        RECT 18.510 181.200 18.830 181.260 ;
        RECT 23.125 181.200 23.415 181.245 ;
        RECT 18.510 181.060 23.415 181.200 ;
        RECT 18.510 181.000 18.830 181.060 ;
        RECT 23.125 181.015 23.415 181.060 ;
        RECT 23.200 180.860 23.340 181.015 ;
        RECT 31.850 181.000 32.170 181.260 ;
        RECT 35.085 181.015 35.375 181.245 ;
        RECT 33.245 180.860 33.535 180.905 ;
        RECT 34.610 180.860 34.930 180.920 ;
        RECT 23.200 180.720 34.930 180.860 ;
        RECT 35.160 180.860 35.300 181.015 ;
        RECT 35.530 181.000 35.850 181.260 ;
        RECT 35.990 181.000 36.310 181.260 ;
        RECT 36.450 181.000 36.770 181.260 ;
        RECT 41.510 181.000 41.830 181.260 ;
        RECT 43.810 181.000 44.130 181.260 ;
        RECT 44.745 181.200 45.035 181.245 ;
        RECT 45.190 181.200 45.510 181.260 ;
        RECT 44.745 181.060 45.510 181.200 ;
        RECT 44.745 181.015 45.035 181.060 ;
        RECT 45.190 181.000 45.510 181.060 ;
        RECT 46.125 181.015 46.415 181.245 ;
        RECT 47.045 181.200 47.335 181.245 ;
        RECT 48.885 181.200 49.175 181.245 ;
        RECT 47.045 181.060 49.175 181.200 ;
        RECT 47.045 181.015 47.335 181.060 ;
        RECT 48.885 181.015 49.175 181.060 ;
        RECT 51.185 181.200 51.475 181.245 ;
        RECT 51.185 181.060 52.320 181.200 ;
        RECT 51.185 181.015 51.475 181.060 ;
        RECT 37.830 180.860 38.150 180.920 ;
        RECT 41.065 180.860 41.355 180.905 ;
        RECT 35.160 180.720 41.355 180.860 ;
        RECT 43.900 180.860 44.040 181.000 ;
        RECT 46.200 180.860 46.340 181.015 ;
        RECT 43.900 180.720 46.340 180.860 ;
        RECT 33.245 180.675 33.535 180.720 ;
        RECT 34.610 180.660 34.930 180.720 ;
        RECT 37.830 180.660 38.150 180.720 ;
        RECT 41.065 180.675 41.355 180.720 ;
        RECT 28.630 180.180 28.950 180.240 ;
        RECT 30.485 180.180 30.775 180.225 ;
        RECT 31.390 180.180 31.710 180.240 ;
        RECT 28.630 180.040 31.710 180.180 ;
        RECT 28.630 179.980 28.950 180.040 ;
        RECT 30.485 179.995 30.775 180.040 ;
        RECT 31.390 179.980 31.710 180.040 ;
        RECT 34.165 180.180 34.455 180.225 ;
        RECT 34.610 180.180 34.930 180.240 ;
        RECT 34.165 180.040 34.930 180.180 ;
        RECT 46.200 180.180 46.340 180.720 ;
        RECT 47.505 180.860 47.795 180.905 ;
        RECT 47.950 180.860 48.270 180.920 ;
        RECT 47.505 180.720 48.270 180.860 ;
        RECT 48.960 180.860 49.100 181.015 ;
        RECT 51.645 180.860 51.935 180.905 ;
        RECT 48.960 180.720 51.935 180.860 ;
        RECT 47.505 180.675 47.795 180.720 ;
        RECT 47.950 180.660 48.270 180.720 ;
        RECT 51.645 180.675 51.935 180.720 ;
        RECT 47.030 180.520 47.350 180.580 ;
        RECT 52.180 180.520 52.320 181.060 ;
        RECT 53.945 181.015 54.235 181.245 ;
        RECT 54.865 181.200 55.155 181.245 ;
        RECT 55.310 181.200 55.630 181.260 ;
        RECT 55.860 181.245 56.000 181.400 ;
        RECT 59.450 181.400 63.450 181.540 ;
        RECT 63.680 181.540 63.820 181.740 ;
        RECT 64.525 181.740 65.750 181.880 ;
        RECT 64.525 181.695 64.815 181.740 ;
        RECT 65.430 181.680 65.750 181.740 ;
        RECT 73.250 181.880 73.570 181.940 ;
        RECT 77.865 181.880 78.155 181.925 ;
        RECT 73.250 181.740 78.155 181.880 ;
        RECT 73.250 181.680 73.570 181.740 ;
        RECT 77.865 181.695 78.155 181.740 ;
        RECT 64.970 181.540 65.290 181.600 ;
        RECT 66.365 181.540 66.655 181.585 ;
        RECT 63.680 181.400 66.655 181.540 ;
        RECT 59.450 181.340 59.770 181.400 ;
        RECT 63.130 181.340 63.450 181.400 ;
        RECT 64.970 181.340 65.290 181.400 ;
        RECT 66.365 181.355 66.655 181.400 ;
        RECT 68.650 181.340 68.970 181.600 ;
        RECT 69.570 181.585 69.890 181.600 ;
        RECT 69.570 181.355 69.955 181.585 ;
        RECT 70.490 181.540 70.810 181.600 ;
        RECT 72.190 181.540 72.480 181.585 ;
        RECT 70.490 181.400 72.480 181.540 ;
        RECT 69.570 181.340 69.890 181.355 ;
        RECT 70.490 181.340 70.810 181.400 ;
        RECT 72.190 181.355 72.480 181.400 ;
        RECT 54.865 181.060 55.630 181.200 ;
        RECT 54.865 181.015 55.155 181.060 ;
        RECT 52.550 180.660 52.870 180.920 ;
        RECT 54.020 180.860 54.160 181.015 ;
        RECT 55.310 181.000 55.630 181.060 ;
        RECT 55.785 181.015 56.075 181.245 ;
        RECT 57.165 181.200 57.455 181.245 ;
        RECT 57.610 181.200 57.930 181.260 ;
        RECT 57.165 181.060 57.930 181.200 ;
        RECT 57.165 181.015 57.455 181.060 ;
        RECT 57.610 181.000 57.930 181.060 ;
        RECT 58.545 181.015 58.835 181.245 ;
        RECT 56.230 180.860 56.550 180.920 ;
        RECT 54.020 180.720 56.550 180.860 ;
        RECT 47.030 180.380 52.320 180.520 ;
        RECT 47.030 180.320 47.350 180.380 ;
        RECT 48.410 180.180 48.730 180.240 ;
        RECT 46.200 180.040 48.730 180.180 ;
        RECT 34.165 179.995 34.455 180.040 ;
        RECT 34.610 179.980 34.930 180.040 ;
        RECT 48.410 179.980 48.730 180.040 ;
        RECT 48.870 180.180 49.190 180.240 ;
        RECT 54.020 180.180 54.160 180.720 ;
        RECT 56.230 180.660 56.550 180.720 ;
        RECT 56.690 180.860 57.010 180.920 ;
        RECT 58.620 180.860 58.760 181.015 ;
        RECT 58.990 181.000 59.310 181.260 ;
        RECT 60.370 181.000 60.690 181.260 ;
        RECT 60.830 181.000 61.150 181.260 ;
        RECT 61.765 181.200 62.055 181.245 ;
        RECT 68.190 181.200 68.510 181.260 ;
        RECT 61.765 181.060 62.900 181.200 ;
        RECT 61.765 181.015 62.055 181.060 ;
        RECT 62.760 180.920 62.900 181.060 ;
        RECT 63.680 181.060 68.510 181.200 ;
        RECT 56.690 180.720 58.760 180.860 ;
        RECT 56.690 180.660 57.010 180.720 ;
        RECT 62.670 180.660 62.990 180.920 ;
        RECT 63.145 180.675 63.435 180.905 ;
        RECT 62.210 180.520 62.530 180.580 ;
        RECT 63.220 180.520 63.360 180.675 ;
        RECT 62.210 180.380 63.360 180.520 ;
        RECT 62.210 180.320 62.530 180.380 ;
        RECT 48.870 180.040 54.160 180.180 ;
        RECT 48.870 179.980 49.190 180.040 ;
        RECT 57.150 179.980 57.470 180.240 ;
        RECT 63.680 180.225 63.820 181.060 ;
        RECT 68.190 181.000 68.510 181.060 ;
        RECT 70.030 180.860 70.350 180.920 ;
        RECT 66.440 180.720 70.350 180.860 ;
        RECT 64.510 180.520 64.830 180.580 ;
        RECT 65.445 180.520 65.735 180.565 ;
        RECT 64.510 180.380 65.735 180.520 ;
        RECT 64.510 180.320 64.830 180.380 ;
        RECT 65.445 180.335 65.735 180.380 ;
        RECT 66.440 180.225 66.580 180.720 ;
        RECT 70.030 180.660 70.350 180.720 ;
        RECT 70.950 180.660 71.270 180.920 ;
        RECT 71.845 180.860 72.135 180.905 ;
        RECT 73.035 180.860 73.325 180.905 ;
        RECT 75.555 180.860 75.845 180.905 ;
        RECT 71.845 180.720 75.845 180.860 ;
        RECT 71.845 180.675 72.135 180.720 ;
        RECT 73.035 180.675 73.325 180.720 ;
        RECT 75.555 180.675 75.845 180.720 ;
        RECT 71.450 180.520 71.740 180.565 ;
        RECT 73.550 180.520 73.840 180.565 ;
        RECT 75.120 180.520 75.410 180.565 ;
        RECT 71.450 180.380 75.410 180.520 ;
        RECT 71.450 180.335 71.740 180.380 ;
        RECT 73.550 180.335 73.840 180.380 ;
        RECT 75.120 180.335 75.410 180.380 ;
        RECT 63.605 179.995 63.895 180.225 ;
        RECT 66.365 179.995 66.655 180.225 ;
        RECT 69.110 180.180 69.430 180.240 ;
        RECT 69.585 180.180 69.875 180.225 ;
        RECT 69.110 180.040 69.875 180.180 ;
        RECT 69.110 179.980 69.430 180.040 ;
        RECT 69.585 179.995 69.875 180.040 ;
        RECT 70.505 180.180 70.795 180.225 ;
        RECT 71.870 180.180 72.190 180.240 ;
        RECT 70.505 180.040 72.190 180.180 ;
        RECT 70.505 179.995 70.795 180.040 ;
        RECT 71.870 179.980 72.190 180.040 ;
        RECT 13.380 179.360 92.040 179.840 ;
        RECT 18.510 179.160 18.830 179.220 ;
        RECT 18.985 179.160 19.275 179.205 ;
        RECT 18.510 179.020 19.275 179.160 ;
        RECT 18.510 178.960 18.830 179.020 ;
        RECT 18.985 178.975 19.275 179.020 ;
        RECT 28.645 179.160 28.935 179.205 ;
        RECT 30.930 179.160 31.250 179.220 ;
        RECT 28.645 179.020 31.250 179.160 ;
        RECT 28.645 178.975 28.935 179.020 ;
        RECT 30.930 178.960 31.250 179.020 ;
        RECT 36.450 179.160 36.770 179.220 ;
        RECT 36.925 179.160 37.215 179.205 ;
        RECT 36.450 179.020 37.215 179.160 ;
        RECT 36.450 178.960 36.770 179.020 ;
        RECT 36.925 178.975 37.215 179.020 ;
        RECT 37.830 178.960 38.150 179.220 ;
        RECT 47.950 178.960 48.270 179.220 ;
        RECT 49.790 178.960 50.110 179.220 ;
        RECT 50.800 179.020 51.860 179.160 ;
        RECT 21.730 178.820 22.020 178.865 ;
        RECT 23.300 178.820 23.590 178.865 ;
        RECT 25.400 178.820 25.690 178.865 ;
        RECT 21.730 178.680 25.690 178.820 ;
        RECT 21.730 178.635 22.020 178.680 ;
        RECT 23.300 178.635 23.590 178.680 ;
        RECT 25.400 178.635 25.690 178.680 ;
        RECT 26.805 178.820 27.095 178.865 ;
        RECT 28.170 178.820 28.490 178.880 ;
        RECT 26.805 178.680 28.490 178.820 ;
        RECT 26.805 178.635 27.095 178.680 ;
        RECT 28.170 178.620 28.490 178.680 ;
        RECT 30.510 178.820 30.800 178.865 ;
        RECT 32.610 178.820 32.900 178.865 ;
        RECT 34.180 178.820 34.470 178.865 ;
        RECT 30.510 178.680 34.470 178.820 ;
        RECT 30.510 178.635 30.800 178.680 ;
        RECT 32.610 178.635 32.900 178.680 ;
        RECT 34.180 178.635 34.470 178.680 ;
        RECT 37.370 178.820 37.690 178.880 ;
        RECT 38.765 178.820 39.055 178.865 ;
        RECT 41.970 178.820 42.290 178.880 ;
        RECT 37.370 178.680 42.290 178.820 ;
        RECT 37.370 178.620 37.690 178.680 ;
        RECT 38.765 178.635 39.055 178.680 ;
        RECT 41.970 178.620 42.290 178.680 ;
        RECT 21.295 178.480 21.585 178.525 ;
        RECT 23.815 178.480 24.105 178.525 ;
        RECT 25.005 178.480 25.295 178.525 ;
        RECT 21.295 178.340 25.295 178.480 ;
        RECT 21.295 178.295 21.585 178.340 ;
        RECT 23.815 178.295 24.105 178.340 ;
        RECT 25.005 178.295 25.295 178.340 ;
        RECT 30.905 178.480 31.195 178.525 ;
        RECT 32.095 178.480 32.385 178.525 ;
        RECT 34.615 178.480 34.905 178.525 ;
        RECT 30.905 178.340 34.905 178.480 ;
        RECT 30.905 178.295 31.195 178.340 ;
        RECT 32.095 178.295 32.385 178.340 ;
        RECT 34.615 178.295 34.905 178.340 ;
        RECT 25.870 177.940 26.190 178.200 ;
        RECT 30.025 178.140 30.315 178.185 ;
        RECT 38.290 178.140 38.610 178.200 ;
        RECT 30.025 178.000 38.610 178.140 ;
        RECT 30.025 177.955 30.315 178.000 ;
        RECT 38.290 177.940 38.610 178.000 ;
        RECT 45.650 178.140 45.970 178.200 ;
        RECT 46.125 178.140 46.415 178.185 ;
        RECT 45.650 178.000 46.415 178.140 ;
        RECT 45.650 177.940 45.970 178.000 ;
        RECT 46.125 177.955 46.415 178.000 ;
        RECT 47.030 177.940 47.350 178.200 ;
        RECT 48.040 178.140 48.180 178.960 ;
        RECT 48.410 178.480 48.730 178.540 ;
        RECT 49.345 178.480 49.635 178.525 ;
        RECT 48.410 178.340 49.635 178.480 ;
        RECT 48.410 178.280 48.730 178.340 ;
        RECT 49.345 178.295 49.635 178.340 ;
        RECT 48.885 178.140 49.175 178.185 ;
        RECT 48.040 178.000 49.175 178.140 ;
        RECT 48.885 177.955 49.175 178.000 ;
        RECT 50.265 178.140 50.555 178.185 ;
        RECT 50.800 178.140 50.940 179.020 ;
        RECT 51.185 178.635 51.475 178.865 ;
        RECT 51.720 178.820 51.860 179.020 ;
        RECT 52.550 178.960 52.870 179.220 ;
        RECT 56.690 178.960 57.010 179.220 ;
        RECT 57.610 178.960 57.930 179.220 ;
        RECT 58.545 179.160 58.835 179.205 ;
        RECT 58.990 179.160 59.310 179.220 ;
        RECT 62.685 179.160 62.975 179.205 ;
        RECT 58.545 179.020 62.975 179.160 ;
        RECT 58.545 178.975 58.835 179.020 ;
        RECT 58.990 178.960 59.310 179.020 ;
        RECT 62.685 178.975 62.975 179.020 ;
        RECT 69.570 179.160 69.890 179.220 ;
        RECT 69.570 179.020 72.100 179.160 ;
        RECT 69.570 178.960 69.890 179.020 ;
        RECT 54.390 178.820 54.710 178.880 ;
        RECT 59.910 178.820 60.230 178.880 ;
        RECT 51.720 178.680 60.230 178.820 ;
        RECT 50.265 178.000 50.940 178.140 ;
        RECT 51.260 178.140 51.400 178.635 ;
        RECT 54.390 178.620 54.710 178.680 ;
        RECT 59.910 178.620 60.230 178.680 ;
        RECT 60.845 178.820 61.135 178.865 ;
        RECT 61.750 178.820 62.070 178.880 ;
        RECT 60.845 178.680 62.070 178.820 ;
        RECT 60.845 178.635 61.135 178.680 ;
        RECT 61.750 178.620 62.070 178.680 ;
        RECT 54.865 178.480 55.155 178.525 ;
        RECT 57.610 178.480 57.930 178.540 ;
        RECT 69.110 178.480 69.430 178.540 ;
        RECT 71.960 178.525 72.100 179.020 ;
        RECT 54.865 178.340 56.230 178.480 ;
        RECT 54.865 178.295 55.155 178.340 ;
        RECT 56.090 178.200 56.230 178.340 ;
        RECT 57.610 178.340 69.430 178.480 ;
        RECT 57.610 178.280 57.930 178.340 ;
        RECT 69.110 178.280 69.430 178.340 ;
        RECT 70.505 178.480 70.795 178.525 ;
        RECT 70.505 178.340 71.640 178.480 ;
        RECT 70.505 178.295 70.795 178.340 ;
        RECT 53.485 178.140 53.775 178.185 ;
        RECT 51.260 178.000 53.775 178.140 ;
        RECT 50.265 177.955 50.555 178.000 ;
        RECT 53.485 177.955 53.775 178.000 ;
        RECT 53.945 177.955 54.235 178.185 ;
        RECT 23.110 177.800 23.430 177.860 ;
        RECT 24.550 177.800 24.840 177.845 ;
        RECT 31.250 177.800 31.540 177.845 ;
        RECT 23.110 177.660 24.840 177.800 ;
        RECT 23.110 177.600 23.430 177.660 ;
        RECT 24.550 177.615 24.840 177.660 ;
        RECT 29.640 177.660 31.540 177.800 ;
        RECT 28.630 177.260 28.950 177.520 ;
        RECT 29.640 177.505 29.780 177.660 ;
        RECT 31.250 177.615 31.540 177.660 ;
        RECT 35.530 177.800 35.850 177.860 ;
        RECT 40.145 177.800 40.435 177.845 ;
        RECT 35.530 177.660 40.435 177.800 ;
        RECT 35.530 177.600 35.850 177.660 ;
        RECT 40.145 177.615 40.435 177.660 ;
        RECT 41.510 177.800 41.830 177.860 ;
        RECT 49.330 177.800 49.650 177.860 ;
        RECT 54.020 177.800 54.160 177.955 ;
        RECT 55.310 177.940 55.630 178.200 ;
        RECT 56.090 178.000 56.550 178.200 ;
        RECT 56.230 177.940 56.550 178.000 ;
        RECT 57.165 178.140 57.455 178.185 ;
        RECT 60.370 178.140 60.690 178.200 ;
        RECT 61.305 178.140 61.595 178.185 ;
        RECT 57.165 178.000 60.140 178.140 ;
        RECT 57.165 177.955 57.455 178.000 ;
        RECT 41.510 177.660 54.160 177.800 ;
        RECT 56.320 177.800 56.460 177.940 ;
        RECT 60.000 177.860 60.140 178.000 ;
        RECT 60.370 178.000 61.595 178.140 ;
        RECT 60.370 177.940 60.690 178.000 ;
        RECT 61.305 177.955 61.595 178.000 ;
        RECT 64.065 177.955 64.355 178.185 ;
        RECT 58.990 177.800 59.310 177.860 ;
        RECT 56.320 177.660 59.310 177.800 ;
        RECT 41.510 177.600 41.830 177.660 ;
        RECT 49.330 177.600 49.650 177.660 ;
        RECT 58.990 177.600 59.310 177.660 ;
        RECT 59.450 177.600 59.770 177.860 ;
        RECT 59.910 177.600 60.230 177.860 ;
        RECT 29.565 177.275 29.855 177.505 ;
        RECT 58.465 177.460 58.755 177.505 ;
        RECT 61.305 177.460 61.595 177.505 ;
        RECT 58.465 177.320 61.595 177.460 ;
        RECT 64.140 177.460 64.280 177.955 ;
        RECT 64.510 177.940 64.830 178.200 ;
        RECT 64.985 178.140 65.275 178.185 ;
        RECT 65.430 178.140 65.750 178.200 ;
        RECT 64.985 178.000 65.750 178.140 ;
        RECT 64.985 177.955 65.275 178.000 ;
        RECT 65.430 177.940 65.750 178.000 ;
        RECT 65.890 177.940 66.210 178.200 ;
        RECT 71.500 178.185 71.640 178.340 ;
        RECT 71.885 178.295 72.175 178.525 ;
        RECT 70.075 177.955 70.365 178.185 ;
        RECT 70.965 177.955 71.255 178.185 ;
        RECT 71.425 177.955 71.715 178.185 ;
        RECT 72.345 178.140 72.635 178.185 ;
        RECT 72.790 178.140 73.110 178.200 ;
        RECT 72.345 178.000 73.110 178.140 ;
        RECT 101.005 178.120 102.595 182.410 ;
        RECT 100.100 178.100 140.370 178.120 ;
        RECT 100.100 178.080 140.860 178.100 ;
        RECT 72.345 177.955 72.635 178.000 ;
        RECT 68.190 177.800 68.510 177.860 ;
        RECT 70.120 177.800 70.260 177.955 ;
        RECT 68.190 177.660 70.260 177.800 ;
        RECT 68.190 177.600 68.510 177.660 ;
        RECT 70.030 177.460 70.350 177.520 ;
        RECT 64.140 177.320 70.350 177.460 ;
        RECT 71.040 177.460 71.180 177.955 ;
        RECT 72.790 177.940 73.110 178.000 ;
        RECT 71.410 177.460 71.730 177.520 ;
        RECT 71.040 177.320 71.730 177.460 ;
        RECT 58.465 177.275 58.755 177.320 ;
        RECT 61.305 177.275 61.595 177.320 ;
        RECT 70.030 177.260 70.350 177.320 ;
        RECT 71.410 177.260 71.730 177.320 ;
        RECT 13.380 176.640 92.040 177.120 ;
        RECT 99.990 177.050 140.860 178.080 ;
        RECT 99.990 176.770 100.770 177.050 ;
        RECT 23.110 176.240 23.430 176.500 ;
        RECT 49.790 176.440 50.110 176.500 ;
        RECT 63.590 176.440 63.910 176.500 ;
        RECT 49.790 176.300 63.910 176.440 ;
        RECT 49.790 176.240 50.110 176.300 ;
        RECT 63.590 176.240 63.910 176.300 ;
        RECT 18.510 176.100 18.830 176.160 ;
        RECT 20.825 176.100 21.115 176.145 ;
        RECT 18.510 175.960 21.115 176.100 ;
        RECT 18.510 175.900 18.830 175.960 ;
        RECT 20.825 175.915 21.115 175.960 ;
        RECT 61.290 176.100 61.610 176.160 ;
        RECT 64.510 176.100 64.830 176.160 ;
        RECT 72.345 176.100 72.635 176.145 ;
        RECT 73.710 176.100 74.030 176.160 ;
        RECT 61.290 175.960 64.830 176.100 ;
        RECT 61.290 175.900 61.610 175.960 ;
        RECT 64.510 175.900 64.830 175.960 ;
        RECT 71.500 175.960 72.635 176.100 ;
        RECT 71.500 175.820 71.640 175.960 ;
        RECT 72.345 175.915 72.635 175.960 ;
        RECT 72.880 175.960 74.030 176.100 ;
        RECT 44.745 175.760 45.035 175.805 ;
        RECT 45.190 175.760 45.510 175.820 ;
        RECT 44.745 175.620 45.510 175.760 ;
        RECT 44.745 175.575 45.035 175.620 ;
        RECT 45.190 175.560 45.510 175.620 ;
        RECT 45.665 175.760 45.955 175.805 ;
        RECT 48.870 175.760 49.190 175.820 ;
        RECT 45.665 175.620 49.190 175.760 ;
        RECT 45.665 175.575 45.955 175.620 ;
        RECT 48.870 175.560 49.190 175.620 ;
        RECT 69.110 175.560 69.430 175.820 ;
        RECT 70.490 175.560 70.810 175.820 ;
        RECT 71.410 175.560 71.730 175.820 ;
        RECT 71.870 175.560 72.190 175.820 ;
        RECT 72.880 175.805 73.020 175.960 ;
        RECT 73.710 175.900 74.030 175.960 ;
        RECT 72.805 175.575 73.095 175.805 ;
        RECT 73.250 175.560 73.570 175.820 ;
        RECT 74.185 175.760 74.475 175.805 ;
        RECT 74.630 175.760 74.950 175.820 ;
        RECT 74.185 175.620 74.950 175.760 ;
        RECT 74.185 175.575 74.475 175.620 ;
        RECT 74.630 175.560 74.950 175.620 ;
        RECT 68.665 175.420 68.955 175.465 ;
        RECT 70.030 175.420 70.350 175.480 ;
        RECT 68.665 175.280 70.350 175.420 ;
        RECT 68.665 175.235 68.955 175.280 ;
        RECT 22.190 175.080 22.510 175.140 ;
        RECT 28.630 175.080 28.950 175.140 ;
        RECT 22.190 174.940 28.950 175.080 ;
        RECT 22.190 174.880 22.510 174.940 ;
        RECT 28.630 174.880 28.950 174.940 ;
        RECT 44.270 175.080 44.590 175.140 ;
        RECT 51.170 175.080 51.490 175.140 ;
        RECT 53.930 175.080 54.250 175.140 ;
        RECT 44.270 174.940 54.250 175.080 ;
        RECT 69.660 175.080 69.800 175.280 ;
        RECT 70.030 175.220 70.350 175.280 ;
        RECT 70.965 175.420 71.255 175.465 ;
        RECT 72.330 175.420 72.650 175.480 ;
        RECT 70.965 175.280 72.650 175.420 ;
        RECT 70.965 175.235 71.255 175.280 ;
        RECT 72.330 175.220 72.650 175.280 ;
        RECT 99.990 175.260 100.880 176.770 ;
        RECT 106.550 176.380 107.800 176.820 ;
        RECT 117.640 176.640 118.600 176.800 ;
        RECT 120.030 176.750 120.810 177.050 ;
        RECT 140.080 176.800 140.860 177.050 ;
        RECT 104.490 176.370 109.730 176.380 ;
        RECT 101.540 176.270 116.840 176.370 ;
        RECT 101.540 176.260 116.875 176.270 ;
        RECT 101.500 176.140 116.875 176.260 ;
        RECT 101.500 176.030 105.500 176.140 ;
        RECT 106.550 176.060 108.290 176.140 ;
        RECT 108.870 176.060 116.875 176.140 ;
        RECT 106.550 175.980 107.800 176.060 ;
        RECT 108.875 176.040 116.875 176.060 ;
        RECT 71.870 175.080 72.190 175.140 ;
        RECT 69.660 174.940 72.190 175.080 ;
        RECT 44.270 174.880 44.590 174.940 ;
        RECT 51.170 174.880 51.490 174.940 ;
        RECT 53.930 174.880 54.250 174.940 ;
        RECT 71.870 174.880 72.190 174.940 ;
        RECT 43.810 174.740 44.130 174.800 ;
        RECT 44.745 174.740 45.035 174.785 ;
        RECT 43.810 174.600 45.035 174.740 ;
        RECT 43.810 174.540 44.130 174.600 ;
        RECT 44.745 174.555 45.035 174.600 ;
        RECT 53.010 174.740 53.330 174.800 ;
        RECT 69.570 174.740 69.890 174.800 ;
        RECT 53.010 174.600 69.890 174.740 ;
        RECT 53.010 174.540 53.330 174.600 ;
        RECT 69.570 174.540 69.890 174.600 ;
        RECT 71.410 174.740 71.730 174.800 ;
        RECT 72.790 174.740 73.110 174.800 ;
        RECT 71.410 174.600 73.110 174.740 ;
        RECT 71.410 174.540 71.730 174.600 ;
        RECT 72.790 174.540 73.110 174.600 ;
        RECT 100.050 174.670 100.880 175.260 ;
        RECT 101.110 175.730 101.340 175.980 ;
        RECT 105.660 175.840 105.890 175.980 ;
        RECT 108.440 175.840 108.670 175.990 ;
        RECT 105.660 175.730 108.670 175.840 ;
        RECT 117.080 175.730 117.310 175.990 ;
        RECT 101.110 175.290 117.310 175.730 ;
        RECT 101.110 175.020 101.340 175.290 ;
        RECT 105.660 175.260 117.310 175.290 ;
        RECT 105.660 175.170 108.670 175.260 ;
        RECT 105.660 175.020 105.890 175.170 ;
        RECT 108.440 175.030 108.670 175.170 ;
        RECT 117.080 175.030 117.310 175.260 ;
        RECT 101.500 174.740 105.500 174.970 ;
        RECT 108.875 174.760 116.875 174.980 ;
        RECT 117.640 174.760 118.880 176.640 ;
        RECT 108.875 174.750 118.880 174.760 ;
        RECT 101.500 174.670 105.490 174.740 ;
        RECT 100.050 174.560 105.490 174.670 ;
        RECT 108.930 174.620 118.880 174.750 ;
        RECT 119.930 175.260 120.810 176.750 ;
        RECT 126.430 176.330 127.680 176.770 ;
        RECT 137.520 176.620 138.480 176.750 ;
        RECT 124.370 176.320 129.610 176.330 ;
        RECT 121.420 176.220 136.720 176.320 ;
        RECT 121.420 176.210 136.755 176.220 ;
        RECT 121.380 176.090 136.755 176.210 ;
        RECT 121.380 175.980 125.380 176.090 ;
        RECT 126.430 176.010 128.170 176.090 ;
        RECT 128.750 176.010 136.755 176.090 ;
        RECT 126.430 175.930 127.680 176.010 ;
        RECT 128.755 175.990 136.755 176.010 ;
        RECT 120.990 175.680 121.220 175.930 ;
        RECT 125.540 175.790 125.770 175.930 ;
        RECT 128.320 175.790 128.550 175.940 ;
        RECT 125.540 175.680 128.550 175.790 ;
        RECT 136.960 175.680 137.190 175.940 ;
        RECT 119.930 174.620 120.760 175.260 ;
        RECT 120.990 175.240 137.190 175.680 ;
        RECT 120.990 174.970 121.220 175.240 ;
        RECT 125.540 175.210 137.190 175.240 ;
        RECT 125.540 175.120 128.550 175.210 ;
        RECT 125.540 174.970 125.770 175.120 ;
        RECT 128.320 174.980 128.550 175.120 ;
        RECT 136.960 174.980 137.190 175.210 ;
        RECT 121.380 174.690 125.380 174.920 ;
        RECT 128.755 174.710 136.755 174.930 ;
        RECT 137.520 174.710 138.700 176.620 ;
        RECT 128.755 174.700 138.700 174.710 ;
        RECT 121.380 174.620 125.370 174.690 ;
        RECT 108.930 174.590 118.600 174.620 ;
        RECT 100.050 174.470 103.180 174.560 ;
        RECT 116.670 174.540 118.600 174.590 ;
        RECT 13.380 173.920 92.040 174.400 ;
        RECT 30.470 173.720 30.790 173.780 ;
        RECT 30.945 173.720 31.235 173.765 ;
        RECT 30.470 173.580 31.235 173.720 ;
        RECT 30.470 173.520 30.790 173.580 ;
        RECT 30.945 173.535 31.235 173.580 ;
        RECT 33.245 173.720 33.535 173.765 ;
        RECT 37.370 173.720 37.690 173.780 ;
        RECT 33.245 173.580 37.690 173.720 ;
        RECT 33.245 173.535 33.535 173.580 ;
        RECT 28.630 173.380 28.950 173.440 ;
        RECT 32.325 173.380 32.615 173.425 ;
        RECT 28.630 173.240 32.615 173.380 ;
        RECT 28.630 173.180 28.950 173.240 ;
        RECT 32.325 173.195 32.615 173.240 ;
        RECT 30.010 173.040 30.330 173.100 ;
        RECT 33.320 173.040 33.460 173.535 ;
        RECT 37.370 173.520 37.690 173.580 ;
        RECT 43.825 173.720 44.115 173.765 ;
        RECT 44.270 173.720 44.590 173.780 ;
        RECT 43.825 173.580 44.590 173.720 ;
        RECT 43.825 173.535 44.115 173.580 ;
        RECT 44.270 173.520 44.590 173.580 ;
        RECT 46.125 173.720 46.415 173.765 ;
        RECT 47.030 173.720 47.350 173.780 ;
        RECT 46.125 173.580 47.350 173.720 ;
        RECT 46.125 173.535 46.415 173.580 ;
        RECT 47.030 173.520 47.350 173.580 ;
        RECT 48.870 173.520 49.190 173.780 ;
        RECT 59.005 173.720 59.295 173.765 ;
        RECT 59.910 173.720 60.230 173.780 ;
        RECT 59.005 173.580 60.230 173.720 ;
        RECT 59.005 173.535 59.295 173.580 ;
        RECT 59.910 173.520 60.230 173.580 ;
        RECT 70.045 173.720 70.335 173.765 ;
        RECT 70.490 173.720 70.810 173.780 ;
        RECT 70.045 173.580 70.810 173.720 ;
        RECT 70.045 173.535 70.335 173.580 ;
        RECT 70.490 173.520 70.810 173.580 ;
        RECT 73.250 173.720 73.570 173.780 ;
        RECT 76.470 173.720 76.790 173.780 ;
        RECT 73.250 173.580 76.790 173.720 ;
        RECT 73.250 173.520 73.570 173.580 ;
        RECT 76.470 173.520 76.790 173.580 ;
        RECT 44.730 173.380 45.050 173.440 ;
        RECT 47.490 173.380 47.810 173.440 ;
        RECT 53.945 173.380 54.235 173.425 ;
        RECT 44.730 173.240 54.235 173.380 ;
        RECT 44.730 173.180 45.050 173.240 ;
        RECT 47.490 173.180 47.810 173.240 ;
        RECT 53.945 173.195 54.235 173.240 ;
        RECT 58.545 173.195 58.835 173.425 ;
        RECT 66.825 173.380 67.115 173.425 ;
        RECT 71.410 173.380 71.730 173.440 ;
        RECT 66.825 173.240 71.730 173.380 ;
        RECT 66.825 173.195 67.115 173.240 ;
        RECT 30.010 172.900 33.460 173.040 ;
        RECT 30.010 172.840 30.330 172.900 ;
        RECT 38.290 172.840 38.610 173.100 ;
        RECT 58.070 173.040 58.390 173.100 ;
        RECT 42.520 172.900 58.390 173.040 ;
        RECT 58.620 173.040 58.760 173.195 ;
        RECT 71.410 173.180 71.730 173.240 ;
        RECT 72.790 173.380 73.110 173.440 ;
        RECT 74.630 173.380 74.950 173.440 ;
        RECT 72.790 173.240 74.950 173.380 ;
        RECT 72.790 173.180 73.110 173.240 ;
        RECT 74.630 173.180 74.950 173.240 ;
        RECT 78.810 173.380 79.100 173.425 ;
        RECT 80.910 173.380 81.200 173.425 ;
        RECT 82.480 173.380 82.770 173.425 ;
        RECT 78.810 173.240 82.770 173.380 ;
        RECT 78.810 173.195 79.100 173.240 ;
        RECT 80.910 173.195 81.200 173.240 ;
        RECT 82.480 173.195 82.770 173.240 ;
        RECT 69.585 173.040 69.875 173.085 ;
        RECT 70.030 173.040 70.350 173.100 ;
        RECT 77.390 173.040 77.710 173.100 ;
        RECT 78.325 173.040 78.615 173.085 ;
        RECT 58.620 172.900 61.980 173.040 ;
        RECT 29.550 172.700 29.870 172.760 ;
        RECT 31.390 172.700 31.710 172.760 ;
        RECT 42.520 172.745 42.660 172.900 ;
        RECT 58.070 172.840 58.390 172.900 ;
        RECT 29.550 172.560 31.710 172.700 ;
        RECT 29.550 172.500 29.870 172.560 ;
        RECT 31.390 172.500 31.710 172.560 ;
        RECT 42.445 172.515 42.735 172.745 ;
        RECT 42.890 172.700 43.210 172.760 ;
        RECT 47.505 172.700 47.795 172.745 ;
        RECT 42.890 172.560 47.795 172.700 ;
        RECT 42.890 172.500 43.210 172.560 ;
        RECT 27.710 172.360 28.030 172.420 ;
        RECT 30.025 172.360 30.315 172.405 ;
        RECT 27.710 172.220 30.315 172.360 ;
        RECT 31.480 172.360 31.620 172.500 ;
        RECT 33.085 172.360 33.375 172.405 ;
        RECT 31.480 172.220 33.375 172.360 ;
        RECT 27.710 172.160 28.030 172.220 ;
        RECT 30.025 172.175 30.315 172.220 ;
        RECT 33.085 172.175 33.375 172.220 ;
        RECT 34.165 172.360 34.455 172.405 ;
        RECT 35.070 172.360 35.390 172.420 ;
        RECT 43.810 172.405 44.130 172.420 ;
        RECT 34.165 172.220 35.390 172.360 ;
        RECT 34.165 172.175 34.455 172.220 ;
        RECT 35.070 172.160 35.390 172.220 ;
        RECT 43.745 172.175 44.130 172.405 ;
        RECT 43.810 172.160 44.130 172.175 ;
        RECT 44.730 172.160 45.050 172.420 ;
        RECT 46.200 172.405 46.340 172.560 ;
        RECT 47.505 172.515 47.795 172.560 ;
        RECT 47.950 172.700 48.270 172.760 ;
        RECT 48.885 172.700 49.175 172.745 ;
        RECT 47.950 172.560 49.175 172.700 ;
        RECT 47.950 172.500 48.270 172.560 ;
        RECT 48.885 172.515 49.175 172.560 ;
        RECT 53.010 172.500 53.330 172.760 ;
        RECT 55.325 172.700 55.615 172.745 ;
        RECT 57.150 172.700 57.470 172.760 ;
        RECT 55.325 172.560 57.470 172.700 ;
        RECT 55.325 172.515 55.615 172.560 ;
        RECT 57.150 172.500 57.470 172.560 ;
        RECT 57.610 172.500 57.930 172.760 ;
        RECT 58.545 172.515 58.835 172.745 ;
        RECT 46.045 172.220 46.340 172.405 ;
        RECT 46.045 172.175 46.335 172.220 ;
        RECT 47.045 172.175 47.335 172.405 ;
        RECT 53.930 172.360 54.250 172.420 ;
        RECT 54.405 172.360 54.695 172.405 ;
        RECT 53.930 172.220 54.695 172.360 ;
        RECT 58.620 172.360 58.760 172.515 ;
        RECT 59.910 172.500 60.230 172.760 ;
        RECT 61.840 172.745 61.980 172.900 ;
        RECT 64.140 172.900 70.350 173.040 ;
        RECT 64.140 172.760 64.280 172.900 ;
        RECT 69.585 172.855 69.875 172.900 ;
        RECT 70.030 172.840 70.350 172.900 ;
        RECT 71.040 172.900 73.940 173.040 ;
        RECT 61.765 172.515 62.055 172.745 ;
        RECT 63.590 172.700 63.910 172.760 ;
        RECT 63.395 172.560 63.910 172.700 ;
        RECT 63.590 172.500 63.910 172.560 ;
        RECT 64.050 172.500 64.370 172.760 ;
        RECT 68.205 172.700 68.495 172.745 ;
        RECT 69.110 172.700 69.430 172.760 ;
        RECT 71.040 172.745 71.180 172.900 ;
        RECT 73.800 172.760 73.940 172.900 ;
        RECT 77.390 172.900 78.615 173.040 ;
        RECT 77.390 172.840 77.710 172.900 ;
        RECT 78.325 172.855 78.615 172.900 ;
        RECT 79.205 173.040 79.495 173.085 ;
        RECT 80.395 173.040 80.685 173.085 ;
        RECT 82.915 173.040 83.205 173.085 ;
        RECT 79.205 172.900 83.205 173.040 ;
        RECT 79.205 172.855 79.495 172.900 ;
        RECT 80.395 172.855 80.685 172.900 ;
        RECT 82.915 172.855 83.205 172.900 ;
        RECT 68.205 172.560 69.430 172.700 ;
        RECT 68.205 172.515 68.495 172.560 ;
        RECT 69.110 172.500 69.430 172.560 ;
        RECT 70.965 172.515 71.255 172.745 ;
        RECT 71.870 172.500 72.190 172.760 ;
        RECT 73.710 172.500 74.030 172.760 ;
        RECT 75.105 172.700 75.395 172.745 ;
        RECT 79.605 172.700 79.895 172.745 ;
        RECT 75.105 172.560 79.895 172.700 ;
        RECT 75.105 172.515 75.395 172.560 ;
        RECT 79.605 172.515 79.895 172.560 ;
        RECT 60.385 172.360 60.675 172.405 ;
        RECT 58.620 172.220 60.675 172.360 ;
        RECT 30.930 172.065 31.250 172.080 ;
        RECT 30.930 171.835 31.315 172.065 ;
        RECT 30.930 171.820 31.250 171.835 ;
        RECT 31.850 171.820 32.170 172.080 ;
        RECT 42.430 172.020 42.750 172.080 ;
        RECT 42.905 172.020 43.195 172.065 ;
        RECT 42.430 171.880 43.195 172.020 ;
        RECT 42.430 171.820 42.750 171.880 ;
        RECT 42.905 171.835 43.195 171.880 ;
        RECT 45.190 171.820 45.510 172.080 ;
        RECT 47.120 172.020 47.260 172.175 ;
        RECT 53.930 172.160 54.250 172.220 ;
        RECT 54.405 172.175 54.695 172.220 ;
        RECT 60.385 172.175 60.675 172.220 ;
        RECT 60.845 172.360 61.135 172.405 ;
        RECT 62.225 172.360 62.515 172.405 ;
        RECT 60.845 172.220 62.515 172.360 ;
        RECT 60.845 172.175 61.135 172.220 ;
        RECT 62.225 172.175 62.515 172.220 ;
        RECT 67.745 172.360 68.035 172.405 ;
        RECT 69.570 172.360 69.890 172.420 ;
        RECT 72.345 172.360 72.635 172.405 ;
        RECT 74.185 172.360 74.475 172.405 ;
        RECT 75.565 172.360 75.855 172.405 ;
        RECT 67.745 172.220 69.340 172.360 ;
        RECT 67.745 172.175 68.035 172.220 ;
        RECT 47.965 172.020 48.255 172.065 ;
        RECT 48.410 172.020 48.730 172.080 ;
        RECT 47.120 171.880 48.730 172.020 ;
        RECT 60.460 172.020 60.600 172.175 ;
        RECT 67.820 172.020 67.960 172.175 ;
        RECT 60.460 171.880 67.960 172.020 ;
        RECT 68.190 172.020 68.510 172.080 ;
        RECT 68.665 172.020 68.955 172.065 ;
        RECT 68.190 171.880 68.955 172.020 ;
        RECT 69.200 172.020 69.340 172.220 ;
        RECT 69.570 172.220 73.940 172.360 ;
        RECT 69.570 172.160 69.890 172.220 ;
        RECT 72.345 172.175 72.635 172.220 ;
        RECT 73.800 172.080 73.940 172.220 ;
        RECT 74.185 172.220 75.855 172.360 ;
        RECT 74.185 172.175 74.475 172.220 ;
        RECT 75.565 172.175 75.855 172.220 ;
        RECT 76.470 172.160 76.790 172.420 ;
        RECT 77.405 172.175 77.695 172.405 ;
        RECT 72.790 172.020 73.110 172.080 ;
        RECT 69.200 171.880 73.110 172.020 ;
        RECT 47.965 171.835 48.255 171.880 ;
        RECT 48.410 171.820 48.730 171.880 ;
        RECT 68.190 171.820 68.510 171.880 ;
        RECT 68.665 171.835 68.955 171.880 ;
        RECT 72.790 171.820 73.110 171.880 ;
        RECT 73.250 171.820 73.570 172.080 ;
        RECT 73.710 171.820 74.030 172.080 ;
        RECT 74.630 172.020 74.950 172.080 ;
        RECT 77.480 172.020 77.620 172.175 ;
        RECT 85.225 172.020 85.515 172.065 ;
        RECT 74.630 171.880 85.515 172.020 ;
        RECT 74.630 171.820 74.950 171.880 ;
        RECT 85.225 171.835 85.515 171.880 ;
        RECT 13.380 171.200 92.040 171.680 ;
        RECT 100.050 171.200 100.880 174.470 ;
        RECT 104.530 174.010 109.780 174.020 ;
        RECT 104.530 173.900 116.840 174.010 ;
        RECT 101.560 173.840 116.840 173.900 ;
        RECT 101.560 173.830 116.875 173.840 ;
        RECT 101.500 173.700 116.875 173.830 ;
        RECT 101.500 173.690 106.660 173.700 ;
        RECT 101.500 173.600 105.500 173.690 ;
        RECT 108.875 173.610 116.875 173.700 ;
        RECT 108.960 173.600 116.850 173.610 ;
        RECT 101.110 173.240 101.340 173.550 ;
        RECT 101.560 173.240 105.460 173.600 ;
        RECT 105.660 173.240 105.890 173.550 ;
        RECT 101.110 171.900 105.890 173.240 ;
        RECT 101.110 171.590 101.340 171.900 ;
        RECT 105.660 171.590 105.890 171.900 ;
        RECT 108.440 173.020 108.670 173.560 ;
        RECT 109.480 173.020 110.490 173.050 ;
        RECT 117.080 173.020 117.310 173.560 ;
        RECT 108.440 172.120 117.310 173.020 ;
        RECT 108.440 171.600 108.670 172.120 ;
        RECT 109.480 172.050 110.490 172.120 ;
        RECT 117.080 171.600 117.310 172.120 ;
        RECT 101.500 171.310 105.500 171.540 ;
        RECT 108.875 171.320 116.875 171.550 ;
        RECT 100.050 171.160 101.180 171.200 ;
        RECT 100.050 171.080 101.420 171.160 ;
        RECT 101.790 171.090 105.450 171.310 ;
        RECT 101.790 171.080 103.230 171.090 ;
        RECT 30.470 170.800 30.790 171.060 ;
        RECT 57.610 171.000 57.930 171.060 ;
        RECT 61.750 171.000 62.070 171.060 ;
        RECT 42.520 170.860 62.070 171.000 ;
        RECT 25.870 170.660 26.190 170.720 ;
        RECT 30.930 170.660 31.250 170.720 ;
        RECT 38.290 170.660 38.610 170.720 ;
        RECT 22.280 170.520 31.250 170.660 ;
        RECT 22.280 170.365 22.420 170.520 ;
        RECT 25.870 170.460 26.190 170.520 ;
        RECT 30.930 170.460 31.250 170.520 ;
        RECT 31.940 170.520 38.610 170.660 ;
        RECT 22.205 170.135 22.495 170.365 ;
        RECT 22.650 170.320 22.970 170.380 ;
        RECT 23.485 170.320 23.775 170.365 ;
        RECT 22.650 170.180 23.775 170.320 ;
        RECT 22.650 170.120 22.970 170.180 ;
        RECT 23.485 170.135 23.775 170.180 ;
        RECT 29.550 170.120 29.870 170.380 ;
        RECT 30.010 170.320 30.330 170.380 ;
        RECT 30.485 170.320 30.775 170.365 ;
        RECT 31.940 170.320 32.080 170.520 ;
        RECT 38.290 170.460 38.610 170.520 ;
        RECT 32.310 170.365 32.630 170.380 ;
        RECT 30.010 170.180 30.775 170.320 ;
        RECT 30.010 170.120 30.330 170.180 ;
        RECT 30.485 170.135 30.775 170.180 ;
        RECT 31.020 170.180 32.080 170.320 ;
        RECT 32.280 170.320 32.630 170.365 ;
        RECT 41.970 170.320 42.290 170.380 ;
        RECT 42.520 170.365 42.660 170.860 ;
        RECT 57.610 170.800 57.930 170.860 ;
        RECT 61.750 170.800 62.070 170.860 ;
        RECT 65.445 171.000 65.735 171.045 ;
        RECT 65.890 171.000 66.210 171.060 ;
        RECT 65.445 170.860 66.210 171.000 ;
        RECT 65.445 170.815 65.735 170.860 ;
        RECT 65.890 170.800 66.210 170.860 ;
        RECT 66.350 170.800 66.670 171.060 ;
        RECT 100.050 171.040 103.230 171.080 ;
        RECT 100.050 170.950 102.740 171.040 ;
        RECT 108.940 171.030 116.830 171.320 ;
        RECT 100.050 170.890 102.070 170.950 ;
        RECT 100.050 170.840 101.820 170.890 ;
        RECT 58.530 170.660 58.850 170.720 ;
        RECT 70.950 170.660 71.270 170.720 ;
        RECT 50.340 170.520 71.270 170.660 ;
        RECT 50.340 170.380 50.480 170.520 ;
        RECT 58.530 170.460 58.850 170.520 ;
        RECT 70.950 170.460 71.270 170.520 ;
        RECT 42.445 170.320 42.735 170.365 ;
        RECT 32.280 170.180 32.780 170.320 ;
        RECT 41.970 170.180 42.735 170.320 ;
        RECT 31.020 170.025 31.160 170.180 ;
        RECT 32.280 170.135 32.630 170.180 ;
        RECT 32.310 170.120 32.630 170.135 ;
        RECT 41.970 170.120 42.290 170.180 ;
        RECT 42.445 170.135 42.735 170.180 ;
        RECT 46.585 170.320 46.875 170.365 ;
        RECT 49.330 170.320 49.650 170.380 ;
        RECT 46.585 170.180 49.650 170.320 ;
        RECT 46.585 170.135 46.875 170.180 ;
        RECT 49.330 170.120 49.650 170.180 ;
        RECT 49.805 170.320 50.095 170.365 ;
        RECT 50.250 170.320 50.570 170.380 ;
        RECT 51.170 170.365 51.490 170.380 ;
        RECT 49.805 170.180 50.570 170.320 ;
        RECT 49.805 170.135 50.095 170.180 ;
        RECT 50.250 170.120 50.570 170.180 ;
        RECT 51.140 170.135 51.490 170.365 ;
        RECT 57.165 170.320 57.455 170.365 ;
        RECT 51.170 170.120 51.490 170.135 ;
        RECT 56.780 170.180 57.455 170.320 ;
        RECT 23.085 169.980 23.375 170.025 ;
        RECT 24.275 169.980 24.565 170.025 ;
        RECT 26.795 169.980 27.085 170.025 ;
        RECT 23.085 169.840 27.085 169.980 ;
        RECT 23.085 169.795 23.375 169.840 ;
        RECT 24.275 169.795 24.565 169.840 ;
        RECT 26.795 169.795 27.085 169.840 ;
        RECT 30.945 169.795 31.235 170.025 ;
        RECT 31.825 169.980 32.115 170.025 ;
        RECT 33.015 169.980 33.305 170.025 ;
        RECT 35.535 169.980 35.825 170.025 ;
        RECT 31.825 169.840 35.825 169.980 ;
        RECT 31.825 169.795 32.115 169.840 ;
        RECT 33.015 169.795 33.305 169.840 ;
        RECT 35.535 169.795 35.825 169.840 ;
        RECT 40.605 169.980 40.895 170.025 ;
        RECT 45.665 169.980 45.955 170.025 ;
        RECT 40.605 169.840 45.955 169.980 ;
        RECT 40.605 169.795 40.895 169.840 ;
        RECT 45.665 169.795 45.955 169.840 ;
        RECT 50.685 169.980 50.975 170.025 ;
        RECT 51.875 169.980 52.165 170.025 ;
        RECT 54.395 169.980 54.685 170.025 ;
        RECT 50.685 169.840 54.685 169.980 ;
        RECT 50.685 169.795 50.975 169.840 ;
        RECT 51.875 169.795 52.165 169.840 ;
        RECT 54.395 169.795 54.685 169.840 ;
        RECT 22.690 169.640 22.980 169.685 ;
        RECT 24.790 169.640 25.080 169.685 ;
        RECT 26.360 169.640 26.650 169.685 ;
        RECT 22.690 169.500 26.650 169.640 ;
        RECT 22.690 169.455 22.980 169.500 ;
        RECT 24.790 169.455 25.080 169.500 ;
        RECT 26.360 169.455 26.650 169.500 ;
        RECT 31.430 169.640 31.720 169.685 ;
        RECT 33.530 169.640 33.820 169.685 ;
        RECT 35.100 169.640 35.390 169.685 ;
        RECT 31.430 169.500 35.390 169.640 ;
        RECT 31.430 169.455 31.720 169.500 ;
        RECT 33.530 169.455 33.820 169.500 ;
        RECT 35.100 169.455 35.390 169.500 ;
        RECT 46.110 169.440 46.430 169.700 ;
        RECT 50.290 169.640 50.580 169.685 ;
        RECT 52.390 169.640 52.680 169.685 ;
        RECT 53.960 169.640 54.250 169.685 ;
        RECT 50.290 169.500 54.250 169.640 ;
        RECT 50.290 169.455 50.580 169.500 ;
        RECT 52.390 169.455 52.680 169.500 ;
        RECT 53.960 169.455 54.250 169.500 ;
        RECT 27.250 169.300 27.570 169.360 ;
        RECT 29.105 169.300 29.395 169.345 ;
        RECT 27.250 169.160 29.395 169.300 ;
        RECT 27.250 169.100 27.570 169.160 ;
        RECT 29.105 169.115 29.395 169.160 ;
        RECT 29.550 169.300 29.870 169.360 ;
        RECT 31.850 169.300 32.170 169.360 ;
        RECT 29.550 169.160 32.170 169.300 ;
        RECT 29.550 169.100 29.870 169.160 ;
        RECT 31.850 169.100 32.170 169.160 ;
        RECT 37.370 169.300 37.690 169.360 ;
        RECT 37.845 169.300 38.135 169.345 ;
        RECT 37.370 169.160 38.135 169.300 ;
        RECT 37.370 169.100 37.690 169.160 ;
        RECT 37.845 169.115 38.135 169.160 ;
        RECT 51.630 169.300 51.950 169.360 ;
        RECT 55.310 169.300 55.630 169.360 ;
        RECT 56.780 169.345 56.920 170.180 ;
        RECT 57.165 170.135 57.455 170.180 ;
        RECT 57.610 170.320 57.930 170.380 ;
        RECT 59.005 170.320 59.295 170.365 ;
        RECT 57.610 170.180 59.295 170.320 ;
        RECT 57.610 170.120 57.930 170.180 ;
        RECT 59.005 170.135 59.295 170.180 ;
        RECT 61.750 170.120 62.070 170.380 ;
        RECT 66.350 170.320 66.640 170.365 ;
        RECT 67.730 170.320 68.050 170.380 ;
        RECT 66.350 170.180 68.050 170.320 ;
        RECT 66.350 170.135 66.640 170.180 ;
        RECT 67.730 170.120 68.050 170.180 ;
        RECT 68.205 170.320 68.495 170.365 ;
        RECT 69.110 170.320 69.430 170.380 ;
        RECT 71.870 170.320 72.190 170.380 ;
        RECT 76.530 170.320 76.820 170.365 ;
        RECT 68.205 170.180 70.030 170.320 ;
        RECT 68.205 170.135 68.495 170.180 ;
        RECT 69.110 170.120 69.430 170.180 ;
        RECT 58.085 169.980 58.375 170.025 ;
        RECT 64.050 169.980 64.370 170.040 ;
        RECT 58.085 169.840 64.370 169.980 ;
        RECT 58.085 169.795 58.375 169.840 ;
        RECT 64.050 169.780 64.370 169.840 ;
        RECT 68.650 169.780 68.970 170.040 ;
        RECT 57.625 169.640 57.915 169.685 ;
        RECT 59.910 169.640 60.230 169.700 ;
        RECT 57.625 169.500 60.230 169.640 ;
        RECT 69.890 169.640 70.030 170.180 ;
        RECT 71.870 170.180 76.820 170.320 ;
        RECT 71.870 170.120 72.190 170.180 ;
        RECT 76.530 170.135 76.820 170.180 ;
        RECT 77.390 170.320 77.710 170.380 ;
        RECT 77.865 170.320 78.155 170.365 ;
        RECT 77.390 170.180 78.155 170.320 ;
        RECT 77.390 170.120 77.710 170.180 ;
        RECT 77.865 170.135 78.155 170.180 ;
        RECT 73.275 169.980 73.565 170.025 ;
        RECT 75.795 169.980 76.085 170.025 ;
        RECT 76.985 169.980 77.275 170.025 ;
        RECT 73.275 169.840 77.275 169.980 ;
        RECT 73.275 169.795 73.565 169.840 ;
        RECT 75.795 169.795 76.085 169.840 ;
        RECT 76.985 169.795 77.275 169.840 ;
        RECT 70.965 169.640 71.255 169.685 ;
        RECT 69.890 169.500 71.255 169.640 ;
        RECT 57.625 169.455 57.915 169.500 ;
        RECT 59.910 169.440 60.230 169.500 ;
        RECT 70.965 169.455 71.255 169.500 ;
        RECT 73.710 169.640 74.000 169.685 ;
        RECT 75.280 169.640 75.570 169.685 ;
        RECT 77.380 169.640 77.670 169.685 ;
        RECT 73.710 169.500 77.670 169.640 ;
        RECT 73.710 169.455 74.000 169.500 ;
        RECT 75.280 169.455 75.570 169.500 ;
        RECT 77.380 169.455 77.670 169.500 ;
        RECT 56.705 169.300 56.995 169.345 ;
        RECT 51.630 169.160 56.995 169.300 ;
        RECT 51.630 169.100 51.950 169.160 ;
        RECT 55.310 169.100 55.630 169.160 ;
        RECT 56.705 169.115 56.995 169.160 ;
        RECT 58.085 169.300 58.375 169.345 ;
        RECT 60.370 169.300 60.690 169.360 ;
        RECT 58.085 169.160 60.690 169.300 ;
        RECT 58.085 169.115 58.375 169.160 ;
        RECT 60.370 169.100 60.690 169.160 ;
        RECT 60.830 169.100 61.150 169.360 ;
        RECT 61.750 169.300 62.070 169.360 ;
        RECT 71.410 169.300 71.730 169.360 ;
        RECT 61.750 169.160 71.730 169.300 ;
        RECT 61.750 169.100 62.070 169.160 ;
        RECT 71.410 169.100 71.730 169.160 ;
        RECT 13.380 168.480 92.040 168.960 ;
        RECT 22.650 168.080 22.970 168.340 ;
        RECT 23.585 168.280 23.875 168.325 ;
        RECT 26.805 168.280 27.095 168.325 ;
        RECT 41.970 168.280 42.290 168.340 ;
        RECT 23.585 168.140 27.095 168.280 ;
        RECT 23.585 168.095 23.875 168.140 ;
        RECT 26.805 168.095 27.095 168.140 ;
        RECT 36.540 168.140 42.290 168.280 ;
        RECT 25.425 167.940 25.715 167.985 ;
        RECT 28.170 167.940 28.490 168.000 ;
        RECT 25.425 167.800 28.490 167.940 ;
        RECT 25.425 167.755 25.715 167.800 ;
        RECT 28.170 167.740 28.490 167.800 ;
        RECT 31.850 167.600 32.170 167.660 ;
        RECT 29.180 167.460 32.170 167.600 ;
        RECT 29.180 167.320 29.320 167.460 ;
        RECT 31.850 167.400 32.170 167.460 ;
        RECT 27.250 167.260 27.570 167.320 ;
        RECT 27.725 167.260 28.015 167.305 ;
        RECT 27.250 167.120 28.015 167.260 ;
        RECT 27.250 167.060 27.570 167.120 ;
        RECT 27.725 167.075 28.015 167.120 ;
        RECT 27.800 166.920 27.940 167.075 ;
        RECT 29.090 167.060 29.410 167.320 ;
        RECT 30.930 167.060 31.250 167.320 ;
        RECT 35.530 167.060 35.850 167.320 ;
        RECT 36.540 167.305 36.680 168.140 ;
        RECT 41.970 168.080 42.290 168.140 ;
        RECT 47.950 168.080 48.270 168.340 ;
        RECT 51.170 168.280 51.490 168.340 ;
        RECT 51.645 168.280 51.935 168.325 ;
        RECT 51.170 168.140 51.935 168.280 ;
        RECT 51.170 168.080 51.490 168.140 ;
        RECT 51.645 168.095 51.935 168.140 ;
        RECT 54.390 168.280 54.710 168.340 ;
        RECT 57.150 168.280 57.470 168.340 ;
        RECT 54.390 168.140 57.470 168.280 ;
        RECT 54.390 168.080 54.710 168.140 ;
        RECT 57.150 168.080 57.470 168.140 ;
        RECT 71.870 168.080 72.190 168.340 ;
        RECT 72.805 168.280 73.095 168.325 ;
        RECT 73.250 168.280 73.570 168.340 ;
        RECT 72.805 168.140 73.570 168.280 ;
        RECT 72.805 168.095 73.095 168.140 ;
        RECT 41.550 167.940 41.840 167.985 ;
        RECT 43.650 167.940 43.940 167.985 ;
        RECT 45.220 167.940 45.510 167.985 ;
        RECT 41.550 167.800 45.510 167.940 ;
        RECT 41.550 167.755 41.840 167.800 ;
        RECT 43.650 167.755 43.940 167.800 ;
        RECT 45.220 167.755 45.510 167.800 ;
        RECT 49.330 167.940 49.650 168.000 ;
        RECT 54.850 167.940 55.170 168.000 ;
        RECT 56.705 167.940 56.995 167.985 ;
        RECT 49.330 167.800 63.820 167.940 ;
        RECT 49.330 167.740 49.650 167.800 ;
        RECT 54.850 167.740 55.170 167.800 ;
        RECT 56.705 167.755 56.995 167.800 ;
        RECT 63.680 167.660 63.820 167.800 ;
        RECT 41.945 167.600 42.235 167.645 ;
        RECT 43.135 167.600 43.425 167.645 ;
        RECT 45.655 167.600 45.945 167.645 ;
        RECT 41.945 167.460 45.945 167.600 ;
        RECT 41.945 167.415 42.235 167.460 ;
        RECT 43.135 167.415 43.425 167.460 ;
        RECT 45.655 167.415 45.945 167.460 ;
        RECT 48.500 167.460 53.700 167.600 ;
        RECT 36.465 167.075 36.755 167.305 ;
        RECT 37.845 167.260 38.135 167.305 ;
        RECT 38.290 167.260 38.610 167.320 ;
        RECT 40.130 167.260 40.450 167.320 ;
        RECT 42.430 167.305 42.750 167.320 ;
        RECT 41.065 167.260 41.355 167.305 ;
        RECT 42.400 167.260 42.750 167.305 ;
        RECT 37.845 167.120 41.355 167.260 ;
        RECT 42.235 167.120 42.750 167.260 ;
        RECT 37.845 167.075 38.135 167.120 ;
        RECT 38.290 167.060 38.610 167.120 ;
        RECT 40.130 167.060 40.450 167.120 ;
        RECT 41.065 167.075 41.355 167.120 ;
        RECT 42.400 167.075 42.750 167.120 ;
        RECT 42.430 167.060 42.750 167.075 ;
        RECT 44.730 167.260 45.050 167.320 ;
        RECT 48.500 167.305 48.640 167.460 ;
        RECT 48.425 167.260 48.715 167.305 ;
        RECT 44.730 167.120 48.715 167.260 ;
        RECT 44.730 167.060 45.050 167.120 ;
        RECT 48.425 167.075 48.715 167.120 ;
        RECT 49.330 167.060 49.650 167.320 ;
        RECT 49.805 167.075 50.095 167.305 ;
        RECT 50.265 167.260 50.555 167.305 ;
        RECT 51.630 167.260 51.950 167.320 ;
        RECT 50.265 167.120 51.950 167.260 ;
        RECT 50.265 167.075 50.555 167.120 ;
        RECT 29.550 166.920 29.870 166.980 ;
        RECT 27.800 166.780 29.870 166.920 ;
        RECT 29.550 166.720 29.870 166.780 ;
        RECT 37.385 166.920 37.675 166.965 ;
        RECT 42.890 166.920 43.210 166.980 ;
        RECT 37.385 166.780 43.210 166.920 ;
        RECT 37.385 166.735 37.675 166.780 ;
        RECT 42.890 166.720 43.210 166.780 ;
        RECT 45.190 166.920 45.510 166.980 ;
        RECT 49.880 166.920 50.020 167.075 ;
        RECT 51.630 167.060 51.950 167.120 ;
        RECT 52.565 167.260 52.855 167.305 ;
        RECT 53.010 167.260 53.330 167.320 ;
        RECT 53.560 167.305 53.700 167.460 ;
        RECT 57.610 167.400 57.930 167.660 ;
        RECT 58.530 167.600 58.850 167.660 ;
        RECT 61.765 167.600 62.055 167.645 ;
        RECT 62.210 167.600 62.530 167.660 ;
        RECT 58.530 167.460 62.530 167.600 ;
        RECT 58.530 167.400 58.850 167.460 ;
        RECT 61.765 167.415 62.055 167.460 ;
        RECT 62.210 167.400 62.530 167.460 ;
        RECT 63.590 167.400 63.910 167.660 ;
        RECT 65.905 167.600 66.195 167.645 ;
        RECT 68.650 167.600 68.970 167.660 ;
        RECT 72.880 167.600 73.020 168.095 ;
        RECT 73.250 168.080 73.570 168.140 ;
        RECT 65.905 167.460 68.970 167.600 ;
        RECT 65.905 167.415 66.195 167.460 ;
        RECT 68.650 167.400 68.970 167.460 ;
        RECT 69.890 167.460 73.020 167.600 ;
        RECT 100.050 167.500 100.880 170.840 ;
        RECT 108.930 170.540 116.850 170.550 ;
        RECT 105.160 170.530 116.850 170.540 ;
        RECT 101.540 170.410 116.850 170.530 ;
        RECT 101.540 170.400 116.875 170.410 ;
        RECT 101.500 170.280 116.875 170.400 ;
        RECT 101.500 170.170 105.500 170.280 ;
        RECT 101.110 169.830 101.340 170.120 ;
        RECT 101.560 169.830 105.450 170.170 ;
        RECT 105.660 169.830 105.890 170.120 ;
        RECT 101.110 168.460 105.890 169.830 ;
        RECT 101.110 168.160 101.340 168.460 ;
        RECT 105.660 168.160 105.890 168.460 ;
        RECT 101.500 167.880 105.500 168.110 ;
        RECT 101.750 167.650 105.320 167.880 ;
        RECT 101.750 167.500 105.440 167.650 ;
        RECT 52.565 167.120 53.330 167.260 ;
        RECT 52.565 167.075 52.855 167.120 ;
        RECT 45.190 166.780 50.020 166.920 ;
        RECT 50.710 166.920 51.030 166.980 ;
        RECT 52.640 166.920 52.780 167.075 ;
        RECT 53.010 167.060 53.330 167.120 ;
        RECT 53.485 167.075 53.775 167.305 ;
        RECT 53.945 167.075 54.235 167.305 ;
        RECT 54.020 166.920 54.160 167.075 ;
        RECT 58.070 167.060 58.390 167.320 ;
        RECT 60.830 167.260 61.150 167.320 ;
        RECT 64.065 167.260 64.355 167.305 ;
        RECT 59.080 167.120 64.355 167.260 ;
        RECT 59.080 166.980 59.220 167.120 ;
        RECT 60.830 167.060 61.150 167.120 ;
        RECT 64.065 167.075 64.355 167.120 ;
        RECT 55.325 166.920 55.615 166.965 ;
        RECT 58.990 166.920 59.310 166.980 ;
        RECT 50.710 166.780 52.780 166.920 ;
        RECT 53.100 166.780 59.310 166.920 ;
        RECT 45.190 166.720 45.510 166.780 ;
        RECT 50.710 166.720 51.030 166.780 ;
        RECT 23.585 166.580 23.875 166.625 ;
        RECT 25.410 166.580 25.730 166.640 ;
        RECT 27.710 166.580 28.030 166.640 ;
        RECT 23.585 166.440 28.030 166.580 ;
        RECT 23.585 166.395 23.875 166.440 ;
        RECT 25.410 166.380 25.730 166.440 ;
        RECT 27.710 166.380 28.030 166.440 ;
        RECT 28.170 166.580 28.490 166.640 ;
        RECT 28.645 166.580 28.935 166.625 ;
        RECT 36.910 166.580 37.230 166.640 ;
        RECT 28.170 166.440 37.230 166.580 ;
        RECT 28.170 166.380 28.490 166.440 ;
        RECT 28.645 166.395 28.935 166.440 ;
        RECT 36.910 166.380 37.230 166.440 ;
        RECT 39.210 166.580 39.530 166.640 ;
        RECT 53.100 166.580 53.240 166.780 ;
        RECT 55.325 166.735 55.615 166.780 ;
        RECT 58.990 166.720 59.310 166.780 ;
        RECT 39.210 166.440 53.240 166.580 ;
        RECT 39.210 166.380 39.530 166.440 ;
        RECT 53.470 166.380 53.790 166.640 ;
        RECT 53.930 166.580 54.250 166.640 ;
        RECT 69.890 166.580 70.030 167.460 ;
        RECT 70.965 167.260 71.255 167.305 ;
        RECT 77.390 167.260 77.710 167.320 ;
        RECT 70.965 167.120 77.710 167.260 ;
        RECT 100.050 167.240 105.440 167.500 ;
        RECT 106.690 167.330 107.310 170.280 ;
        RECT 108.875 170.180 116.875 170.280 ;
        RECT 108.930 170.170 116.850 170.180 ;
        RECT 108.440 169.470 108.670 170.130 ;
        RECT 109.450 169.470 110.450 169.560 ;
        RECT 117.080 169.470 117.310 170.130 ;
        RECT 108.440 168.650 117.310 169.470 ;
        RECT 108.440 168.170 108.670 168.650 ;
        RECT 109.450 168.560 110.450 168.650 ;
        RECT 117.080 168.170 117.310 168.650 ;
        RECT 108.875 167.890 116.875 168.120 ;
        RECT 70.965 167.075 71.255 167.120 ;
        RECT 77.390 167.060 77.710 167.120 ;
        RECT 100.010 167.220 105.440 167.240 ;
        RECT 72.330 166.965 72.650 166.980 ;
        RECT 72.330 166.735 72.935 166.965 ;
        RECT 72.330 166.720 72.650 166.735 ;
        RECT 73.710 166.720 74.030 166.980 ;
        RECT 100.010 166.760 105.450 167.220 ;
        RECT 53.930 166.440 70.030 166.580 ;
        RECT 53.930 166.380 54.250 166.440 ;
        RECT 13.380 165.760 92.040 166.240 ;
        RECT 27.265 165.560 27.555 165.605 ;
        RECT 29.090 165.560 29.410 165.620 ;
        RECT 27.265 165.420 29.410 165.560 ;
        RECT 27.265 165.375 27.555 165.420 ;
        RECT 29.090 165.360 29.410 165.420 ;
        RECT 33.690 165.560 34.010 165.620 ;
        RECT 46.110 165.560 46.430 165.620 ;
        RECT 60.370 165.560 60.690 165.620 ;
        RECT 33.690 165.420 60.690 165.560 ;
        RECT 33.690 165.360 34.010 165.420 ;
        RECT 46.110 165.360 46.430 165.420 ;
        RECT 60.370 165.360 60.690 165.420 ;
        RECT 64.525 165.560 64.815 165.605 ;
        RECT 66.350 165.560 66.670 165.620 ;
        RECT 64.525 165.420 66.670 165.560 ;
        RECT 64.525 165.375 64.815 165.420 ;
        RECT 66.350 165.360 66.670 165.420 ;
        RECT 100.010 165.410 102.050 166.760 ;
        RECT 103.800 166.750 105.450 166.760 ;
        RECT 102.490 165.480 103.490 166.200 ;
        RECT 103.800 165.940 104.110 166.750 ;
        RECT 104.570 166.470 105.450 166.750 ;
        RECT 105.690 166.930 107.310 167.330 ;
        RECT 108.960 166.980 116.830 167.890 ;
        RECT 104.510 166.240 105.510 166.470 ;
        RECT 105.690 166.280 106.040 166.930 ;
        RECT 106.690 166.920 107.310 166.930 ;
        RECT 108.875 166.750 116.875 166.980 ;
        RECT 108.960 166.740 116.830 166.750 ;
        RECT 104.570 166.030 105.450 166.050 ;
        RECT 103.840 165.650 104.110 165.940 ;
        RECT 104.510 165.800 105.510 166.030 ;
        RECT 105.670 165.990 106.040 166.280 ;
        RECT 105.700 165.930 106.040 165.990 ;
        RECT 106.800 166.600 107.560 166.650 ;
        RECT 108.440 166.600 108.670 166.700 ;
        RECT 106.800 166.390 108.670 166.600 ;
        RECT 117.080 166.390 117.310 166.700 ;
        RECT 106.800 165.970 109.340 166.390 ;
        RECT 116.710 165.970 117.310 166.390 ;
        RECT 104.570 165.650 105.450 165.800 ;
        RECT 104.580 165.480 105.310 165.650 ;
        RECT 24.045 165.220 24.335 165.265 ;
        RECT 28.630 165.220 28.950 165.280 ;
        RECT 24.045 165.080 28.950 165.220 ;
        RECT 24.045 165.035 24.335 165.080 ;
        RECT 28.630 165.020 28.950 165.080 ;
        RECT 36.465 165.220 36.755 165.265 ;
        RECT 39.210 165.220 39.530 165.280 ;
        RECT 36.465 165.080 39.530 165.220 ;
        RECT 36.465 165.035 36.755 165.080 ;
        RECT 39.210 165.020 39.530 165.080 ;
        RECT 58.070 165.220 58.390 165.280 ;
        RECT 67.270 165.220 67.590 165.280 ;
        RECT 68.665 165.220 68.955 165.265 ;
        RECT 58.070 165.080 68.955 165.220 ;
        RECT 58.070 165.020 58.390 165.080 ;
        RECT 67.270 165.020 67.590 165.080 ;
        RECT 68.665 165.035 68.955 165.080 ;
        RECT 72.805 165.220 73.095 165.265 ;
        RECT 77.390 165.220 77.710 165.280 ;
        RECT 72.805 165.080 77.710 165.220 ;
        RECT 72.805 165.035 73.095 165.080 ;
        RECT 77.390 165.020 77.710 165.080 ;
        RECT 24.965 164.695 25.255 164.925 ;
        RECT 25.040 164.540 25.180 164.695 ;
        RECT 27.710 164.680 28.030 164.940 ;
        RECT 28.185 164.880 28.475 164.925 ;
        RECT 29.550 164.880 29.870 164.940 ;
        RECT 28.185 164.740 32.080 164.880 ;
        RECT 28.185 164.695 28.475 164.740 ;
        RECT 29.550 164.680 29.870 164.740 ;
        RECT 30.485 164.540 30.775 164.585 ;
        RECT 30.930 164.540 31.250 164.600 ;
        RECT 25.040 164.400 29.320 164.540 ;
        RECT 29.180 164.245 29.320 164.400 ;
        RECT 30.485 164.400 31.250 164.540 ;
        RECT 31.940 164.540 32.080 164.740 ;
        RECT 34.150 164.680 34.470 164.940 ;
        RECT 35.545 164.695 35.835 164.925 ;
        RECT 36.925 164.880 37.215 164.925 ;
        RECT 37.370 164.880 37.690 164.940 ;
        RECT 36.925 164.740 37.690 164.880 ;
        RECT 36.925 164.695 37.215 164.740 ;
        RECT 35.070 164.540 35.390 164.600 ;
        RECT 35.620 164.540 35.760 164.695 ;
        RECT 37.370 164.680 37.690 164.740 ;
        RECT 58.530 164.680 58.850 164.940 ;
        RECT 58.990 164.880 59.310 164.940 ;
        RECT 63.590 164.925 63.910 164.940 ;
        RECT 62.685 164.880 62.975 164.925 ;
        RECT 58.990 164.740 62.975 164.880 ;
        RECT 58.990 164.680 59.310 164.740 ;
        RECT 62.685 164.695 62.975 164.740 ;
        RECT 63.455 164.695 63.910 164.925 ;
        RECT 63.590 164.680 63.910 164.695 ;
        RECT 64.050 164.880 64.370 164.940 ;
        RECT 65.905 164.880 66.195 164.925 ;
        RECT 64.050 164.740 66.195 164.880 ;
        RECT 64.050 164.680 64.370 164.740 ;
        RECT 65.905 164.695 66.195 164.740 ;
        RECT 37.830 164.540 38.150 164.600 ;
        RECT 31.940 164.400 38.150 164.540 ;
        RECT 30.485 164.355 30.775 164.400 ;
        RECT 30.930 164.340 31.250 164.400 ;
        RECT 35.070 164.340 35.390 164.400 ;
        RECT 37.830 164.340 38.150 164.400 ;
        RECT 29.105 164.200 29.395 164.245 ;
        RECT 31.850 164.200 32.170 164.260 ;
        RECT 29.105 164.060 32.170 164.200 ;
        RECT 29.105 164.015 29.395 164.060 ;
        RECT 31.850 164.000 32.170 164.060 ;
        RECT 25.870 163.660 26.190 163.920 ;
        RECT 26.330 163.660 26.650 163.920 ;
        RECT 32.770 163.860 33.090 163.920 ;
        RECT 34.625 163.860 34.915 163.905 ;
        RECT 32.770 163.720 34.915 163.860 ;
        RECT 63.680 163.860 63.820 164.680 ;
        RECT 64.970 163.860 65.290 163.920 ;
        RECT 66.365 163.860 66.655 163.905 ;
        RECT 63.680 163.720 66.655 163.860 ;
        RECT 32.770 163.660 33.090 163.720 ;
        RECT 34.625 163.675 34.915 163.720 ;
        RECT 64.970 163.660 65.290 163.720 ;
        RECT 66.365 163.675 66.655 163.720 ;
        RECT 13.380 163.040 92.040 163.520 ;
        RECT 25.870 162.840 26.190 162.900 ;
        RECT 28.645 162.840 28.935 162.885 ;
        RECT 25.870 162.700 28.935 162.840 ;
        RECT 25.870 162.640 26.190 162.700 ;
        RECT 28.645 162.655 28.935 162.700 ;
        RECT 31.390 162.840 31.710 162.900 ;
        RECT 31.865 162.840 32.155 162.885 ;
        RECT 37.370 162.840 37.690 162.900 ;
        RECT 31.390 162.700 32.155 162.840 ;
        RECT 31.390 162.640 31.710 162.700 ;
        RECT 31.865 162.655 32.155 162.700 ;
        RECT 32.400 162.700 37.690 162.840 ;
        RECT 26.330 162.500 26.650 162.560 ;
        RECT 26.805 162.500 27.095 162.545 ;
        RECT 26.330 162.360 27.095 162.500 ;
        RECT 26.330 162.300 26.650 162.360 ;
        RECT 26.805 162.315 27.095 162.360 ;
        RECT 32.400 162.160 32.540 162.700 ;
        RECT 37.370 162.640 37.690 162.700 ;
        RECT 42.890 162.840 43.210 162.900 ;
        RECT 42.890 162.700 56.460 162.840 ;
        RECT 42.890 162.640 43.210 162.700 ;
        RECT 33.690 162.500 34.010 162.560 ;
        RECT 35.070 162.500 35.390 162.560 ;
        RECT 36.465 162.500 36.755 162.545 ;
        RECT 33.690 162.360 34.380 162.500 ;
        RECT 33.690 162.300 34.010 162.360 ;
        RECT 29.640 162.020 32.540 162.160 ;
        RECT 22.650 161.820 22.970 161.880 ;
        RECT 22.650 161.680 27.480 161.820 ;
        RECT 22.650 161.620 22.970 161.680 ;
        RECT 27.340 161.480 27.480 161.680 ;
        RECT 28.645 161.480 28.935 161.525 ;
        RECT 27.340 161.340 28.935 161.480 ;
        RECT 29.640 161.480 29.780 162.020 ;
        RECT 30.025 161.820 30.315 161.865 ;
        RECT 32.310 161.820 32.630 161.880 ;
        RECT 30.025 161.680 32.630 161.820 ;
        RECT 30.025 161.635 30.315 161.680 ;
        RECT 32.310 161.620 32.630 161.680 ;
        RECT 32.770 161.620 33.090 161.880 ;
        RECT 34.240 161.865 34.380 162.360 ;
        RECT 35.070 162.360 36.755 162.500 ;
        RECT 35.070 162.300 35.390 162.360 ;
        RECT 36.465 162.315 36.755 162.360 ;
        RECT 38.750 162.500 39.070 162.560 ;
        RECT 38.750 162.360 50.940 162.500 ;
        RECT 38.750 162.300 39.070 162.360 ;
        RECT 34.610 161.960 34.930 162.220 ;
        RECT 36.925 162.160 37.215 162.205 ;
        RECT 35.620 162.020 37.215 162.160 ;
        RECT 35.620 161.865 35.760 162.020 ;
        RECT 36.925 161.975 37.215 162.020 ;
        RECT 37.370 162.160 37.690 162.220 ;
        RECT 37.370 162.020 38.980 162.160 ;
        RECT 37.370 161.960 37.690 162.020 ;
        RECT 33.705 161.820 33.995 161.865 ;
        RECT 33.595 161.680 33.995 161.820 ;
        RECT 33.705 161.635 33.995 161.680 ;
        RECT 34.165 161.820 34.455 161.865 ;
        RECT 34.165 161.680 34.565 161.820 ;
        RECT 34.165 161.635 34.455 161.680 ;
        RECT 35.545 161.635 35.835 161.865 ;
        RECT 30.945 161.480 31.235 161.525 ;
        RECT 29.640 161.340 31.235 161.480 ;
        RECT 28.645 161.295 28.935 161.340 ;
        RECT 30.945 161.295 31.235 161.340 ;
        RECT 31.850 161.480 32.170 161.540 ;
        RECT 33.780 161.480 33.920 161.635 ;
        RECT 31.850 161.340 33.920 161.480 ;
        RECT 34.240 161.480 34.380 161.635 ;
        RECT 37.830 161.620 38.150 161.880 ;
        RECT 38.840 161.865 38.980 162.020 ;
        RECT 42.890 161.960 43.210 162.220 ;
        RECT 50.800 162.205 50.940 162.360 ;
        RECT 50.725 161.975 51.015 162.205 ;
        RECT 38.765 161.635 39.055 161.865 ;
        RECT 39.210 161.620 39.530 161.880 ;
        RECT 42.430 161.620 42.750 161.880 ;
        RECT 49.805 161.820 50.095 161.865 ;
        RECT 42.980 161.680 50.095 161.820 ;
        RECT 34.610 161.480 34.930 161.540 ;
        RECT 34.240 161.340 34.930 161.480 ;
        RECT 31.850 161.280 32.170 161.340 ;
        RECT 34.610 161.280 34.930 161.340 ;
        RECT 41.970 161.480 42.290 161.540 ;
        RECT 42.980 161.480 43.120 161.680 ;
        RECT 49.805 161.635 50.095 161.680 ;
        RECT 50.250 161.620 50.570 161.880 ;
        RECT 51.185 161.820 51.475 161.865 ;
        RECT 54.390 161.820 54.710 161.880 ;
        RECT 56.320 161.865 56.460 162.700 ;
        RECT 60.920 162.360 68.880 162.500 ;
        RECT 59.465 162.160 59.755 162.205 ;
        RECT 59.465 162.020 60.600 162.160 ;
        RECT 59.465 161.975 59.755 162.020 ;
        RECT 54.865 161.820 55.155 161.865 ;
        RECT 51.185 161.680 55.155 161.820 ;
        RECT 51.185 161.635 51.475 161.680 ;
        RECT 54.390 161.620 54.710 161.680 ;
        RECT 54.865 161.635 55.155 161.680 ;
        RECT 56.245 161.635 56.535 161.865 ;
        RECT 58.990 161.620 59.310 161.880 ;
        RECT 60.460 161.865 60.600 162.020 ;
        RECT 59.925 161.820 60.215 161.865 ;
        RECT 59.815 161.680 60.215 161.820 ;
        RECT 60.460 161.680 60.775 161.865 ;
        RECT 59.925 161.635 60.215 161.680 ;
        RECT 60.485 161.635 60.775 161.680 ;
        RECT 41.970 161.340 43.120 161.480 ;
        RECT 47.965 161.480 48.255 161.525 ;
        RECT 47.965 161.340 55.080 161.480 ;
        RECT 41.970 161.280 42.290 161.340 ;
        RECT 47.965 161.295 48.255 161.340 ;
        RECT 54.940 161.200 55.080 161.340 ;
        RECT 55.785 161.295 56.075 161.525 ;
        RECT 60.000 161.480 60.140 161.635 ;
        RECT 60.920 161.480 61.060 162.360 ;
        RECT 63.605 162.160 63.895 162.205 ;
        RECT 61.380 162.020 63.895 162.160 ;
        RECT 61.380 161.865 61.520 162.020 ;
        RECT 63.605 161.975 63.895 162.020 ;
        RECT 68.205 161.975 68.495 162.205 ;
        RECT 61.305 161.635 61.595 161.865 ;
        RECT 61.765 161.635 62.055 161.865 ;
        RECT 62.345 161.820 62.635 161.865 ;
        RECT 64.970 161.820 65.290 161.880 ;
        RECT 62.300 161.635 62.635 161.820 ;
        RECT 64.775 161.680 65.290 161.820 ;
        RECT 61.840 161.480 61.980 161.635 ;
        RECT 60.000 161.340 61.980 161.480 ;
        RECT 29.550 160.940 29.870 161.200 ;
        RECT 40.590 160.940 40.910 161.200 ;
        RECT 47.490 160.940 47.810 161.200 ;
        RECT 48.410 161.140 48.730 161.200 ;
        RECT 48.885 161.140 49.175 161.185 ;
        RECT 48.410 161.000 49.175 161.140 ;
        RECT 48.410 160.940 48.730 161.000 ;
        RECT 48.885 160.955 49.175 161.000 ;
        RECT 53.470 161.140 53.790 161.200 ;
        RECT 53.945 161.140 54.235 161.185 ;
        RECT 53.470 161.000 54.235 161.140 ;
        RECT 53.470 160.940 53.790 161.000 ;
        RECT 53.945 160.955 54.235 161.000 ;
        RECT 54.850 160.940 55.170 161.200 ;
        RECT 55.310 161.140 55.630 161.200 ;
        RECT 55.860 161.140 56.000 161.295 ;
        RECT 57.165 161.140 57.455 161.185 ;
        RECT 62.300 161.140 62.440 161.635 ;
        RECT 64.970 161.620 65.290 161.680 ;
        RECT 65.430 161.820 65.750 161.880 ;
        RECT 68.280 161.820 68.420 161.975 ;
        RECT 68.740 161.865 68.880 162.360 ;
        RECT 70.505 162.160 70.795 162.205 ;
        RECT 73.390 162.160 73.680 162.205 ;
        RECT 70.505 162.020 73.680 162.160 ;
        RECT 70.505 161.975 70.795 162.020 ;
        RECT 73.390 161.975 73.680 162.020 ;
        RECT 65.430 161.680 68.420 161.820 ;
        RECT 68.665 161.820 68.955 161.865 ;
        RECT 70.030 161.820 70.350 161.880 ;
        RECT 68.665 161.680 70.350 161.820 ;
        RECT 65.430 161.620 65.750 161.680 ;
        RECT 68.665 161.635 68.955 161.680 ;
        RECT 70.030 161.620 70.350 161.680 ;
        RECT 70.950 161.620 71.270 161.880 ;
        RECT 72.330 161.620 72.650 161.880 ;
        RECT 72.790 161.620 73.110 161.880 ;
        RECT 100.010 161.770 100.780 165.410 ;
        RECT 102.460 164.360 105.310 165.480 ;
        RECT 105.700 165.180 106.050 165.930 ;
        RECT 106.800 165.810 108.670 165.970 ;
        RECT 106.800 165.760 107.560 165.810 ;
        RECT 108.440 165.740 108.670 165.810 ;
        RECT 117.080 165.740 117.310 165.970 ;
        RECT 108.875 165.460 116.875 165.690 ;
        RECT 105.700 165.120 105.990 165.180 ;
        RECT 105.610 165.000 105.990 165.120 ;
        RECT 108.970 165.060 116.830 165.460 ;
        RECT 117.640 165.060 118.600 174.540 ;
        RECT 119.930 174.510 125.370 174.620 ;
        RECT 128.810 174.600 138.700 174.700 ;
        RECT 139.960 175.280 140.860 176.800 ;
        RECT 146.460 176.380 147.710 176.820 ;
        RECT 144.400 176.370 149.640 176.380 ;
        RECT 141.450 176.270 156.750 176.370 ;
        RECT 141.450 176.260 156.785 176.270 ;
        RECT 141.410 176.140 156.785 176.260 ;
        RECT 141.410 176.030 145.410 176.140 ;
        RECT 146.460 176.060 148.200 176.140 ;
        RECT 148.780 176.060 156.785 176.140 ;
        RECT 146.460 175.980 147.710 176.060 ;
        RECT 148.785 176.040 156.785 176.060 ;
        RECT 141.020 175.730 141.250 175.980 ;
        RECT 145.570 175.840 145.800 175.980 ;
        RECT 148.350 175.840 148.580 175.990 ;
        RECT 145.570 175.730 148.580 175.840 ;
        RECT 156.990 175.730 157.220 175.990 ;
        RECT 141.020 175.290 157.220 175.730 ;
        RECT 139.960 174.670 140.790 175.280 ;
        RECT 141.020 175.020 141.250 175.290 ;
        RECT 145.570 175.260 157.220 175.290 ;
        RECT 145.570 175.170 148.580 175.260 ;
        RECT 145.570 175.020 145.800 175.170 ;
        RECT 148.350 175.030 148.580 175.170 ;
        RECT 156.990 175.030 157.220 175.260 ;
        RECT 141.410 174.740 145.410 174.970 ;
        RECT 148.785 174.760 156.785 174.980 ;
        RECT 157.550 174.760 158.510 176.800 ;
        RECT 148.785 174.750 158.510 174.760 ;
        RECT 141.410 174.670 145.400 174.740 ;
        RECT 128.810 174.540 138.480 174.600 ;
        RECT 119.930 174.420 123.060 174.510 ;
        RECT 136.550 174.490 138.480 174.540 ;
        RECT 119.930 171.150 120.760 174.420 ;
        RECT 124.410 173.960 129.660 173.970 ;
        RECT 124.410 173.850 136.720 173.960 ;
        RECT 121.440 173.790 136.720 173.850 ;
        RECT 121.440 173.780 136.755 173.790 ;
        RECT 121.380 173.650 136.755 173.780 ;
        RECT 121.380 173.640 126.540 173.650 ;
        RECT 121.380 173.550 125.380 173.640 ;
        RECT 128.755 173.560 136.755 173.650 ;
        RECT 128.840 173.550 136.730 173.560 ;
        RECT 120.990 173.190 121.220 173.500 ;
        RECT 121.440 173.190 125.340 173.550 ;
        RECT 125.540 173.190 125.770 173.500 ;
        RECT 120.990 171.850 125.770 173.190 ;
        RECT 120.990 171.540 121.220 171.850 ;
        RECT 125.540 171.540 125.770 171.850 ;
        RECT 128.320 172.970 128.550 173.510 ;
        RECT 129.360 172.970 130.370 173.000 ;
        RECT 136.960 172.970 137.190 173.510 ;
        RECT 128.320 172.070 137.190 172.970 ;
        RECT 128.320 171.550 128.550 172.070 ;
        RECT 129.360 172.000 130.370 172.070 ;
        RECT 136.960 171.550 137.190 172.070 ;
        RECT 121.380 171.260 125.380 171.490 ;
        RECT 128.755 171.270 136.755 171.500 ;
        RECT 119.930 171.110 121.060 171.150 ;
        RECT 119.930 171.030 121.300 171.110 ;
        RECT 121.670 171.040 125.330 171.260 ;
        RECT 121.670 171.030 123.110 171.040 ;
        RECT 119.930 170.990 123.110 171.030 ;
        RECT 119.930 170.900 122.620 170.990 ;
        RECT 128.820 170.980 136.710 171.270 ;
        RECT 119.930 170.840 121.950 170.900 ;
        RECT 119.930 170.790 121.700 170.840 ;
        RECT 119.930 167.450 120.760 170.790 ;
        RECT 128.810 170.490 136.730 170.500 ;
        RECT 125.040 170.480 136.730 170.490 ;
        RECT 121.420 170.360 136.730 170.480 ;
        RECT 121.420 170.350 136.755 170.360 ;
        RECT 121.380 170.230 136.755 170.350 ;
        RECT 121.380 170.120 125.380 170.230 ;
        RECT 120.990 169.780 121.220 170.070 ;
        RECT 121.440 169.780 125.330 170.120 ;
        RECT 125.540 169.780 125.770 170.070 ;
        RECT 120.990 168.410 125.770 169.780 ;
        RECT 120.990 168.110 121.220 168.410 ;
        RECT 125.540 168.110 125.770 168.410 ;
        RECT 121.380 167.830 125.380 168.060 ;
        RECT 121.630 167.600 125.200 167.830 ;
        RECT 121.630 167.450 125.320 167.600 ;
        RECT 119.930 167.170 125.320 167.450 ;
        RECT 126.570 167.280 127.190 170.230 ;
        RECT 128.755 170.130 136.755 170.230 ;
        RECT 128.810 170.120 136.730 170.130 ;
        RECT 128.320 169.420 128.550 170.080 ;
        RECT 129.330 169.420 130.330 169.510 ;
        RECT 136.960 169.420 137.190 170.080 ;
        RECT 128.320 168.600 137.190 169.420 ;
        RECT 128.320 168.120 128.550 168.600 ;
        RECT 129.330 168.510 130.330 168.600 ;
        RECT 136.960 168.120 137.190 168.600 ;
        RECT 128.755 167.840 136.755 168.070 ;
        RECT 119.930 166.710 125.330 167.170 ;
        RECT 119.930 165.370 121.930 166.710 ;
        RECT 123.680 166.700 125.330 166.710 ;
        RECT 122.370 165.430 123.370 166.150 ;
        RECT 123.680 165.890 123.990 166.700 ;
        RECT 124.450 166.420 125.330 166.700 ;
        RECT 125.570 166.880 127.190 167.280 ;
        RECT 128.840 166.930 136.710 167.840 ;
        RECT 124.390 166.190 125.390 166.420 ;
        RECT 125.570 166.230 125.920 166.880 ;
        RECT 126.570 166.870 127.190 166.880 ;
        RECT 128.755 166.700 136.755 166.930 ;
        RECT 128.840 166.690 136.710 166.700 ;
        RECT 124.450 165.980 125.330 166.000 ;
        RECT 123.720 165.600 123.990 165.890 ;
        RECT 124.390 165.750 125.390 165.980 ;
        RECT 125.550 165.940 125.920 166.230 ;
        RECT 125.580 165.880 125.920 165.940 ;
        RECT 126.680 166.550 127.440 166.600 ;
        RECT 128.320 166.550 128.550 166.650 ;
        RECT 126.680 166.340 128.550 166.550 ;
        RECT 136.960 166.340 137.190 166.650 ;
        RECT 126.680 165.920 129.220 166.340 ;
        RECT 136.590 165.920 137.190 166.340 ;
        RECT 124.450 165.600 125.330 165.750 ;
        RECT 124.460 165.430 125.190 165.600 ;
        RECT 102.400 164.130 105.400 164.360 ;
        RECT 105.610 164.170 105.950 165.000 ;
        RECT 107.960 164.990 118.600 165.060 ;
        RECT 102.450 164.100 105.310 164.130 ;
        RECT 102.450 164.080 103.620 164.100 ;
        RECT 104.580 164.090 105.310 164.100 ;
        RECT 102.400 163.690 105.400 163.920 ;
        RECT 105.605 163.880 105.950 164.170 ;
        RECT 106.140 163.950 118.600 164.990 ;
        RECT 120.000 165.360 121.930 165.370 ;
        RECT 106.140 163.930 118.560 163.950 ;
        RECT 105.610 163.770 105.950 163.880 ;
        RECT 106.180 163.920 111.850 163.930 ;
        RECT 112.850 163.920 118.560 163.930 ;
        RECT 102.490 163.520 105.350 163.690 ;
        RECT 106.180 163.520 106.610 163.920 ;
        RECT 102.460 163.150 106.610 163.520 ;
        RECT 55.310 161.000 62.440 161.140 ;
        RECT 55.310 160.940 55.630 161.000 ;
        RECT 57.165 160.955 57.455 161.000 ;
        RECT 63.130 160.940 63.450 161.200 ;
        RECT 74.185 161.140 74.475 161.185 ;
        RECT 74.630 161.140 74.950 161.200 ;
        RECT 74.185 161.000 74.950 161.140 ;
        RECT 74.185 160.955 74.475 161.000 ;
        RECT 74.630 160.940 74.950 161.000 ;
        RECT 13.380 160.320 92.040 160.800 ;
        RECT 24.505 159.935 24.795 160.165 ;
        RECT 24.580 159.440 24.720 159.935 ;
        RECT 31.390 159.920 31.710 160.180 ;
        RECT 31.850 160.120 32.170 160.180 ;
        RECT 32.785 160.120 33.075 160.165 ;
        RECT 31.850 159.980 33.075 160.120 ;
        RECT 31.850 159.920 32.170 159.980 ;
        RECT 32.785 159.935 33.075 159.980 ;
        RECT 38.765 160.120 39.055 160.165 ;
        RECT 42.890 160.120 43.210 160.180 ;
        RECT 47.045 160.120 47.335 160.165 ;
        RECT 50.250 160.120 50.570 160.180 ;
        RECT 38.765 159.980 43.210 160.120 ;
        RECT 46.835 159.980 50.570 160.120 ;
        RECT 38.765 159.935 39.055 159.980 ;
        RECT 42.890 159.920 43.210 159.980 ;
        RECT 47.045 159.935 47.335 159.980 ;
        RECT 29.550 159.780 29.870 159.840 ;
        RECT 30.070 159.780 30.360 159.825 ;
        RECT 29.550 159.640 30.360 159.780 ;
        RECT 29.550 159.580 29.870 159.640 ;
        RECT 30.070 159.595 30.360 159.640 ;
        RECT 31.480 159.440 31.620 159.920 ;
        RECT 41.970 159.780 42.290 159.840 ;
        RECT 37.920 159.640 42.290 159.780 ;
        RECT 33.690 159.440 34.010 159.500 ;
        RECT 37.920 159.485 38.060 159.640 ;
        RECT 41.970 159.580 42.290 159.640 ;
        RECT 42.430 159.780 42.750 159.840 ;
        RECT 47.120 159.780 47.260 159.935 ;
        RECT 50.250 159.920 50.570 159.980 ;
        RECT 54.390 159.920 54.710 160.180 ;
        RECT 62.210 159.780 62.530 159.840 ;
        RECT 73.710 159.780 74.030 159.840 ;
        RECT 74.630 159.825 74.950 159.840 ;
        RECT 42.430 159.640 47.260 159.780 ;
        RECT 47.580 159.640 62.530 159.780 ;
        RECT 42.430 159.580 42.750 159.640 ;
        RECT 24.580 159.300 34.010 159.440 ;
        RECT 33.690 159.240 34.010 159.300 ;
        RECT 37.845 159.255 38.135 159.485 ;
        RECT 38.750 159.440 39.070 159.500 ;
        RECT 39.670 159.440 39.990 159.500 ;
        RECT 38.750 159.300 39.990 159.440 ;
        RECT 38.750 159.240 39.070 159.300 ;
        RECT 39.670 159.240 39.990 159.300 ;
        RECT 40.130 159.240 40.450 159.500 ;
        RECT 41.510 159.485 41.830 159.500 ;
        RECT 47.580 159.485 47.720 159.640 ;
        RECT 62.210 159.580 62.530 159.640 ;
        RECT 69.890 159.640 74.030 159.780 ;
        RECT 48.870 159.485 49.190 159.500 ;
        RECT 41.480 159.255 41.830 159.485 ;
        RECT 47.505 159.255 47.795 159.485 ;
        RECT 48.840 159.255 49.190 159.485 ;
        RECT 41.510 159.240 41.830 159.255 ;
        RECT 48.870 159.240 49.190 159.255 ;
        RECT 53.470 159.440 53.790 159.500 ;
        RECT 57.165 159.440 57.455 159.485 ;
        RECT 53.470 159.300 57.455 159.440 ;
        RECT 53.470 159.240 53.790 159.300 ;
        RECT 57.165 159.255 57.455 159.300 ;
        RECT 57.610 159.440 57.930 159.500 ;
        RECT 58.085 159.440 58.375 159.485 ;
        RECT 57.610 159.300 58.375 159.440 ;
        RECT 57.610 159.240 57.930 159.300 ;
        RECT 58.085 159.255 58.375 159.300 ;
        RECT 58.545 159.440 58.835 159.485 ;
        RECT 65.430 159.440 65.750 159.500 ;
        RECT 69.890 159.440 70.030 159.640 ;
        RECT 73.710 159.580 74.030 159.640 ;
        RECT 74.600 159.595 74.950 159.825 ;
        RECT 74.630 159.580 74.950 159.595 ;
        RECT 75.550 159.580 75.870 159.840 ;
        RECT 100.010 159.670 100.880 161.770 ;
        RECT 106.550 161.380 107.800 161.820 ;
        RECT 117.700 161.800 118.560 163.920 ;
        RECT 120.000 161.800 120.770 165.360 ;
        RECT 122.340 164.310 125.190 165.430 ;
        RECT 125.580 165.130 125.930 165.880 ;
        RECT 126.680 165.760 128.550 165.920 ;
        RECT 126.680 165.710 127.440 165.760 ;
        RECT 128.320 165.690 128.550 165.760 ;
        RECT 136.960 165.690 137.190 165.920 ;
        RECT 128.755 165.410 136.755 165.640 ;
        RECT 125.580 165.070 125.870 165.130 ;
        RECT 125.490 164.950 125.870 165.070 ;
        RECT 128.850 165.010 136.710 165.410 ;
        RECT 137.520 165.010 138.480 174.490 ;
        RECT 139.960 174.560 145.400 174.670 ;
        RECT 148.840 174.590 158.510 174.750 ;
        RECT 139.960 174.470 143.090 174.560 ;
        RECT 156.580 174.540 158.510 174.590 ;
        RECT 139.960 171.200 140.790 174.470 ;
        RECT 144.440 174.010 149.690 174.020 ;
        RECT 144.440 173.900 156.750 174.010 ;
        RECT 141.470 173.840 156.750 173.900 ;
        RECT 141.470 173.830 156.785 173.840 ;
        RECT 141.410 173.700 156.785 173.830 ;
        RECT 141.410 173.690 146.570 173.700 ;
        RECT 141.410 173.600 145.410 173.690 ;
        RECT 148.785 173.610 156.785 173.700 ;
        RECT 148.870 173.600 156.760 173.610 ;
        RECT 141.020 173.240 141.250 173.550 ;
        RECT 141.470 173.240 145.370 173.600 ;
        RECT 145.570 173.240 145.800 173.550 ;
        RECT 141.020 171.900 145.800 173.240 ;
        RECT 141.020 171.590 141.250 171.900 ;
        RECT 145.570 171.590 145.800 171.900 ;
        RECT 148.350 173.020 148.580 173.560 ;
        RECT 149.390 173.020 150.400 173.050 ;
        RECT 156.990 173.020 157.220 173.560 ;
        RECT 148.350 172.120 157.220 173.020 ;
        RECT 148.350 171.600 148.580 172.120 ;
        RECT 149.390 172.050 150.400 172.120 ;
        RECT 156.990 171.600 157.220 172.120 ;
        RECT 141.410 171.310 145.410 171.540 ;
        RECT 148.785 171.320 156.785 171.550 ;
        RECT 139.960 171.160 141.090 171.200 ;
        RECT 139.960 171.080 141.330 171.160 ;
        RECT 141.700 171.090 145.360 171.310 ;
        RECT 141.700 171.080 143.140 171.090 ;
        RECT 139.960 171.040 143.140 171.080 ;
        RECT 139.960 170.950 142.650 171.040 ;
        RECT 148.850 171.030 156.740 171.320 ;
        RECT 139.960 170.890 141.980 170.950 ;
        RECT 139.960 170.840 141.730 170.890 ;
        RECT 139.960 167.500 140.790 170.840 ;
        RECT 148.840 170.540 156.760 170.550 ;
        RECT 145.070 170.530 156.760 170.540 ;
        RECT 141.450 170.410 156.760 170.530 ;
        RECT 141.450 170.400 156.785 170.410 ;
        RECT 141.410 170.280 156.785 170.400 ;
        RECT 141.410 170.170 145.410 170.280 ;
        RECT 141.020 169.830 141.250 170.120 ;
        RECT 141.470 169.830 145.360 170.170 ;
        RECT 145.570 169.830 145.800 170.120 ;
        RECT 141.020 168.460 145.800 169.830 ;
        RECT 141.020 168.160 141.250 168.460 ;
        RECT 145.570 168.160 145.800 168.460 ;
        RECT 141.410 167.880 145.410 168.110 ;
        RECT 141.660 167.650 145.230 167.880 ;
        RECT 141.660 167.500 145.350 167.650 ;
        RECT 139.960 167.270 145.350 167.500 ;
        RECT 146.600 167.330 147.220 170.280 ;
        RECT 148.785 170.180 156.785 170.280 ;
        RECT 148.840 170.170 156.760 170.180 ;
        RECT 148.350 169.470 148.580 170.130 ;
        RECT 149.360 169.470 150.360 169.560 ;
        RECT 156.990 169.470 157.220 170.130 ;
        RECT 148.350 168.650 157.220 169.470 ;
        RECT 148.350 168.170 148.580 168.650 ;
        RECT 149.360 168.560 150.360 168.650 ;
        RECT 156.990 168.170 157.220 168.650 ;
        RECT 148.785 167.890 156.785 168.120 ;
        RECT 122.280 164.080 125.280 164.310 ;
        RECT 125.490 164.120 125.830 164.950 ;
        RECT 127.840 164.940 138.480 165.010 ;
        RECT 122.330 164.050 125.190 164.080 ;
        RECT 122.330 164.030 123.500 164.050 ;
        RECT 124.460 164.040 125.190 164.050 ;
        RECT 122.280 163.640 125.280 163.870 ;
        RECT 125.485 163.830 125.830 164.120 ;
        RECT 126.020 163.900 138.480 164.940 ;
        RECT 139.930 167.220 145.350 167.270 ;
        RECT 139.930 166.760 145.360 167.220 ;
        RECT 139.930 165.410 141.960 166.760 ;
        RECT 143.710 166.750 145.360 166.760 ;
        RECT 142.400 165.480 143.400 166.200 ;
        RECT 143.710 165.940 144.020 166.750 ;
        RECT 144.480 166.470 145.360 166.750 ;
        RECT 145.600 166.930 147.220 167.330 ;
        RECT 148.870 166.980 156.740 167.890 ;
        RECT 144.420 166.240 145.420 166.470 ;
        RECT 145.600 166.280 145.950 166.930 ;
        RECT 146.600 166.920 147.220 166.930 ;
        RECT 148.785 166.750 156.785 166.980 ;
        RECT 148.870 166.740 156.740 166.750 ;
        RECT 144.480 166.030 145.360 166.050 ;
        RECT 143.750 165.650 144.020 165.940 ;
        RECT 144.420 165.800 145.420 166.030 ;
        RECT 145.580 165.990 145.950 166.280 ;
        RECT 145.610 165.930 145.950 165.990 ;
        RECT 146.710 166.600 147.470 166.650 ;
        RECT 148.350 166.600 148.580 166.700 ;
        RECT 146.710 166.390 148.580 166.600 ;
        RECT 156.990 166.390 157.220 166.700 ;
        RECT 146.710 165.970 149.250 166.390 ;
        RECT 156.620 165.970 157.220 166.390 ;
        RECT 144.480 165.650 145.360 165.800 ;
        RECT 144.490 165.480 145.220 165.650 ;
        RECT 126.020 163.880 138.460 163.900 ;
        RECT 125.490 163.720 125.830 163.830 ;
        RECT 126.060 163.870 131.730 163.880 ;
        RECT 132.730 163.870 138.460 163.880 ;
        RECT 122.370 163.470 125.230 163.640 ;
        RECT 126.060 163.470 126.490 163.870 ;
        RECT 122.340 163.100 126.490 163.470 ;
        RECT 104.490 161.370 109.730 161.380 ;
        RECT 101.540 161.270 116.840 161.370 ;
        RECT 101.540 161.260 116.875 161.270 ;
        RECT 101.500 161.140 116.875 161.260 ;
        RECT 101.500 161.030 105.500 161.140 ;
        RECT 106.550 161.060 108.290 161.140 ;
        RECT 108.870 161.060 116.875 161.140 ;
        RECT 106.550 160.980 107.800 161.060 ;
        RECT 108.875 161.040 116.875 161.060 ;
        RECT 101.110 160.730 101.340 160.980 ;
        RECT 105.660 160.840 105.890 160.980 ;
        RECT 108.440 160.840 108.670 160.990 ;
        RECT 105.660 160.730 108.670 160.840 ;
        RECT 117.080 160.730 117.310 160.990 ;
        RECT 101.110 160.290 117.310 160.730 ;
        RECT 101.110 160.020 101.340 160.290 ;
        RECT 105.660 160.260 117.310 160.290 ;
        RECT 105.660 160.170 108.670 160.260 ;
        RECT 105.660 160.020 105.890 160.170 ;
        RECT 108.440 160.030 108.670 160.170 ;
        RECT 117.080 160.030 117.310 160.260 ;
        RECT 101.500 159.740 105.500 159.970 ;
        RECT 108.875 159.760 116.875 159.980 ;
        RECT 117.640 159.760 118.600 161.800 ;
        RECT 108.875 159.750 118.600 159.760 ;
        RECT 101.500 159.670 105.490 159.740 ;
        RECT 75.640 159.440 75.780 159.580 ;
        RECT 58.545 159.300 70.030 159.440 ;
        RECT 72.880 159.300 75.780 159.440 ;
        RECT 100.010 159.560 105.490 159.670 ;
        RECT 108.930 159.590 118.600 159.750 ;
        RECT 100.010 159.470 103.180 159.560 ;
        RECT 116.670 159.540 118.600 159.590 ;
        RECT 58.545 159.255 58.835 159.300 ;
        RECT 65.430 159.240 65.750 159.300 ;
        RECT 72.880 159.160 73.020 159.300 ;
        RECT 26.815 159.100 27.105 159.145 ;
        RECT 29.335 159.100 29.625 159.145 ;
        RECT 30.525 159.100 30.815 159.145 ;
        RECT 26.815 158.960 30.815 159.100 ;
        RECT 26.815 158.915 27.105 158.960 ;
        RECT 29.335 158.915 29.625 158.960 ;
        RECT 30.525 158.915 30.815 158.960 ;
        RECT 31.390 158.900 31.710 159.160 ;
        RECT 35.085 159.100 35.375 159.145 ;
        RECT 35.990 159.100 36.310 159.160 ;
        RECT 35.085 158.960 36.310 159.100 ;
        RECT 35.085 158.915 35.375 158.960 ;
        RECT 35.990 158.900 36.310 158.960 ;
        RECT 41.025 159.100 41.315 159.145 ;
        RECT 42.215 159.100 42.505 159.145 ;
        RECT 44.735 159.100 45.025 159.145 ;
        RECT 41.025 158.960 45.025 159.100 ;
        RECT 41.025 158.915 41.315 158.960 ;
        RECT 42.215 158.915 42.505 158.960 ;
        RECT 44.735 158.915 45.025 158.960 ;
        RECT 48.385 159.100 48.675 159.145 ;
        RECT 49.575 159.100 49.865 159.145 ;
        RECT 52.095 159.100 52.385 159.145 ;
        RECT 48.385 158.960 52.385 159.100 ;
        RECT 48.385 158.915 48.675 158.960 ;
        RECT 49.575 158.915 49.865 158.960 ;
        RECT 52.095 158.915 52.385 158.960 ;
        RECT 54.850 159.100 55.170 159.160 ;
        RECT 72.790 159.100 73.110 159.160 ;
        RECT 54.850 158.960 73.110 159.100 ;
        RECT 54.850 158.900 55.170 158.960 ;
        RECT 72.790 158.900 73.110 158.960 ;
        RECT 73.265 159.100 73.555 159.145 ;
        RECT 74.145 159.100 74.435 159.145 ;
        RECT 75.335 159.100 75.625 159.145 ;
        RECT 77.855 159.100 78.145 159.145 ;
        RECT 73.265 158.915 73.605 159.100 ;
        RECT 74.145 158.960 78.145 159.100 ;
        RECT 74.145 158.915 74.435 158.960 ;
        RECT 75.335 158.915 75.625 158.960 ;
        RECT 77.855 158.915 78.145 158.960 ;
        RECT 27.250 158.760 27.540 158.805 ;
        RECT 28.820 158.760 29.110 158.805 ;
        RECT 30.920 158.760 31.210 158.805 ;
        RECT 27.250 158.620 31.210 158.760 ;
        RECT 27.250 158.575 27.540 158.620 ;
        RECT 28.820 158.575 29.110 158.620 ;
        RECT 30.920 158.575 31.210 158.620 ;
        RECT 40.630 158.760 40.920 158.805 ;
        RECT 42.730 158.760 43.020 158.805 ;
        RECT 44.300 158.760 44.590 158.805 ;
        RECT 40.630 158.620 44.590 158.760 ;
        RECT 40.630 158.575 40.920 158.620 ;
        RECT 42.730 158.575 43.020 158.620 ;
        RECT 44.300 158.575 44.590 158.620 ;
        RECT 47.990 158.760 48.280 158.805 ;
        RECT 50.090 158.760 50.380 158.805 ;
        RECT 51.660 158.760 51.950 158.805 ;
        RECT 47.990 158.620 51.950 158.760 ;
        RECT 47.990 158.575 48.280 158.620 ;
        RECT 50.090 158.575 50.380 158.620 ;
        RECT 51.660 158.575 51.950 158.620 ;
        RECT 52.550 158.760 52.870 158.820 ;
        RECT 70.950 158.760 71.270 158.820 ;
        RECT 71.870 158.760 72.190 158.820 ;
        RECT 52.550 158.620 72.190 158.760 ;
        RECT 52.550 158.560 52.870 158.620 ;
        RECT 70.950 158.560 71.270 158.620 ;
        RECT 71.870 158.560 72.190 158.620 ;
        RECT 34.625 158.420 34.915 158.465 ;
        RECT 35.530 158.420 35.850 158.480 ;
        RECT 34.625 158.280 35.850 158.420 ;
        RECT 34.625 158.235 34.915 158.280 ;
        RECT 35.530 158.220 35.850 158.280 ;
        RECT 56.245 158.420 56.535 158.465 ;
        RECT 61.290 158.420 61.610 158.480 ;
        RECT 56.245 158.280 61.610 158.420 ;
        RECT 56.245 158.235 56.535 158.280 ;
        RECT 61.290 158.220 61.610 158.280 ;
        RECT 61.750 158.420 62.070 158.480 ;
        RECT 72.790 158.420 73.110 158.480 ;
        RECT 61.750 158.280 73.110 158.420 ;
        RECT 73.465 158.420 73.605 158.915 ;
        RECT 73.750 158.760 74.040 158.805 ;
        RECT 75.850 158.760 76.140 158.805 ;
        RECT 77.420 158.760 77.710 158.805 ;
        RECT 73.750 158.620 77.710 158.760 ;
        RECT 73.750 158.575 74.040 158.620 ;
        RECT 75.850 158.575 76.140 158.620 ;
        RECT 77.420 158.575 77.710 158.620 ;
        RECT 78.310 158.420 78.630 158.480 ;
        RECT 73.465 158.280 78.630 158.420 ;
        RECT 61.750 158.220 62.070 158.280 ;
        RECT 72.790 158.220 73.110 158.280 ;
        RECT 78.310 158.220 78.630 158.280 ;
        RECT 80.150 158.220 80.470 158.480 ;
        RECT 13.380 157.600 92.040 158.080 ;
        RECT 40.605 157.400 40.895 157.445 ;
        RECT 41.510 157.400 41.830 157.460 ;
        RECT 40.605 157.260 41.830 157.400 ;
        RECT 40.605 157.215 40.895 157.260 ;
        RECT 41.510 157.200 41.830 157.260 ;
        RECT 48.870 157.200 49.190 157.460 ;
        RECT 54.405 157.400 54.695 157.445 ;
        RECT 54.850 157.400 55.170 157.460 ;
        RECT 54.405 157.260 55.170 157.400 ;
        RECT 54.405 157.215 54.695 157.260 ;
        RECT 54.850 157.200 55.170 157.260 ;
        RECT 60.845 157.400 61.135 157.445 ;
        RECT 63.130 157.400 63.450 157.460 ;
        RECT 60.845 157.260 63.450 157.400 ;
        RECT 60.845 157.215 61.135 157.260 ;
        RECT 63.130 157.200 63.450 157.260 ;
        RECT 71.870 157.400 72.190 157.460 ;
        RECT 74.170 157.400 74.490 157.460 ;
        RECT 71.870 157.260 74.490 157.400 ;
        RECT 71.870 157.200 72.190 157.260 ;
        RECT 74.170 157.200 74.490 157.260 ;
        RECT 52.550 157.060 52.870 157.120 ;
        RECT 45.740 156.920 52.870 157.060 ;
        RECT 26.330 156.720 26.650 156.780 ;
        RECT 33.690 156.720 34.010 156.780 ;
        RECT 35.085 156.720 35.375 156.765 ;
        RECT 26.330 156.580 27.940 156.720 ;
        RECT 26.330 156.520 26.650 156.580 ;
        RECT 26.805 156.380 27.095 156.425 ;
        RECT 27.250 156.380 27.570 156.440 ;
        RECT 27.800 156.425 27.940 156.580 ;
        RECT 33.690 156.580 35.375 156.720 ;
        RECT 33.690 156.520 34.010 156.580 ;
        RECT 35.085 156.535 35.375 156.580 ;
        RECT 40.590 156.720 40.910 156.780 ;
        RECT 45.740 156.765 45.880 156.920 ;
        RECT 52.550 156.860 52.870 156.920 ;
        RECT 57.165 157.060 57.455 157.105 ;
        RECT 58.085 157.060 58.375 157.105 ;
        RECT 61.750 157.060 62.070 157.120 ;
        RECT 68.205 157.060 68.495 157.105 ;
        RECT 57.165 156.920 58.375 157.060 ;
        RECT 57.165 156.875 57.455 156.920 ;
        RECT 58.085 156.875 58.375 156.920 ;
        RECT 58.620 156.920 62.070 157.060 ;
        RECT 41.400 156.720 41.690 156.765 ;
        RECT 40.590 156.580 41.690 156.720 ;
        RECT 40.590 156.520 40.910 156.580 ;
        RECT 41.400 156.535 41.690 156.580 ;
        RECT 43.825 156.720 44.115 156.765 ;
        RECT 45.665 156.720 45.955 156.765 ;
        RECT 58.620 156.720 58.760 156.920 ;
        RECT 61.750 156.860 62.070 156.920 ;
        RECT 64.600 156.920 68.495 157.060 ;
        RECT 43.825 156.580 45.955 156.720 ;
        RECT 43.825 156.535 44.115 156.580 ;
        RECT 45.665 156.535 45.955 156.580 ;
        RECT 51.260 156.580 58.760 156.720 ;
        RECT 59.925 156.720 60.215 156.765 ;
        RECT 63.590 156.720 63.910 156.780 ;
        RECT 59.925 156.580 63.910 156.720 ;
        RECT 26.805 156.240 27.570 156.380 ;
        RECT 26.805 156.195 27.095 156.240 ;
        RECT 27.250 156.180 27.570 156.240 ;
        RECT 27.725 156.195 28.015 156.425 ;
        RECT 34.165 156.380 34.455 156.425 ;
        RECT 34.610 156.380 34.930 156.440 ;
        RECT 34.165 156.240 34.930 156.380 ;
        RECT 34.165 156.195 34.455 156.240 ;
        RECT 34.610 156.180 34.930 156.240 ;
        RECT 47.950 156.425 48.270 156.440 ;
        RECT 47.950 156.195 48.380 156.425 ;
        RECT 47.950 156.180 48.270 156.195 ;
        RECT 42.445 156.040 42.735 156.085 ;
        RECT 47.045 156.040 47.335 156.085 ;
        RECT 49.790 156.040 50.110 156.100 ;
        RECT 42.445 155.900 50.110 156.040 ;
        RECT 42.445 155.855 42.735 155.900 ;
        RECT 47.045 155.855 47.335 155.900 ;
        RECT 49.790 155.840 50.110 155.900 ;
        RECT 23.570 155.700 23.890 155.760 ;
        RECT 26.805 155.700 27.095 155.745 ;
        RECT 23.570 155.560 27.095 155.700 ;
        RECT 23.570 155.500 23.890 155.560 ;
        RECT 26.805 155.515 27.095 155.560 ;
        RECT 31.850 155.700 32.170 155.760 ;
        RECT 33.245 155.700 33.535 155.745 ;
        RECT 31.850 155.560 33.535 155.700 ;
        RECT 31.850 155.500 32.170 155.560 ;
        RECT 33.245 155.515 33.535 155.560 ;
        RECT 41.985 155.700 42.275 155.745 ;
        RECT 42.890 155.700 43.210 155.760 ;
        RECT 47.490 155.700 47.810 155.760 ;
        RECT 51.260 155.700 51.400 156.580 ;
        RECT 59.925 156.535 60.215 156.580 ;
        RECT 63.590 156.520 63.910 156.580 ;
        RECT 64.600 156.440 64.740 156.920 ;
        RECT 68.205 156.875 68.495 156.920 ;
        RECT 72.790 157.060 73.110 157.120 ;
        RECT 75.090 157.060 75.410 157.120 ;
        RECT 72.790 156.920 75.410 157.060 ;
        RECT 72.790 156.860 73.110 156.920 ;
        RECT 75.090 156.860 75.410 156.920 ;
        RECT 78.810 157.060 79.100 157.105 ;
        RECT 80.910 157.060 81.200 157.105 ;
        RECT 82.480 157.060 82.770 157.105 ;
        RECT 78.810 156.920 82.770 157.060 ;
        RECT 78.810 156.875 79.100 156.920 ;
        RECT 80.910 156.875 81.200 156.920 ;
        RECT 82.480 156.875 82.770 156.920 ;
        RECT 66.350 156.520 66.670 156.780 ;
        RECT 68.650 156.720 68.970 156.780 ;
        RECT 70.505 156.720 70.795 156.765 ;
        RECT 77.850 156.720 78.170 156.780 ;
        RECT 68.650 156.580 70.795 156.720 ;
        RECT 68.650 156.520 68.970 156.580 ;
        RECT 70.505 156.535 70.795 156.580 ;
        RECT 72.880 156.580 78.170 156.720 ;
        RECT 54.390 156.380 54.710 156.440 ;
        RECT 55.030 156.380 55.320 156.425 ;
        RECT 54.390 156.240 55.320 156.380 ;
        RECT 54.390 156.180 54.710 156.240 ;
        RECT 55.030 156.195 55.320 156.240 ;
        RECT 57.610 156.180 57.930 156.440 ;
        RECT 58.990 156.180 59.310 156.440 ;
        RECT 61.290 156.180 61.610 156.440 ;
        RECT 62.670 156.180 62.990 156.440 ;
        RECT 63.145 156.195 63.435 156.425 ;
        RECT 64.065 156.380 64.355 156.425 ;
        RECT 63.680 156.240 64.355 156.380 ;
        RECT 63.220 156.040 63.360 156.195 ;
        RECT 56.090 155.900 63.360 156.040 ;
        RECT 41.985 155.560 51.400 155.700 ;
        RECT 54.390 155.700 54.710 155.760 ;
        RECT 55.310 155.700 55.630 155.760 ;
        RECT 56.090 155.700 56.230 155.900 ;
        RECT 54.390 155.560 56.230 155.700 ;
        RECT 41.985 155.515 42.275 155.560 ;
        RECT 42.890 155.500 43.210 155.560 ;
        RECT 47.490 155.500 47.810 155.560 ;
        RECT 54.390 155.500 54.710 155.560 ;
        RECT 55.310 155.500 55.630 155.560 ;
        RECT 61.750 155.500 62.070 155.760 ;
        RECT 63.680 155.700 63.820 156.240 ;
        RECT 64.065 156.195 64.355 156.240 ;
        RECT 64.510 156.180 64.830 156.440 ;
        RECT 66.810 156.180 67.130 156.440 ;
        RECT 70.030 156.180 70.350 156.440 ;
        RECT 71.870 156.180 72.190 156.440 ;
        RECT 72.880 156.425 73.020 156.580 ;
        RECT 77.850 156.520 78.170 156.580 ;
        RECT 78.310 156.520 78.630 156.780 ;
        RECT 79.205 156.720 79.495 156.765 ;
        RECT 80.395 156.720 80.685 156.765 ;
        RECT 82.915 156.720 83.205 156.765 ;
        RECT 79.205 156.580 83.205 156.720 ;
        RECT 79.205 156.535 79.495 156.580 ;
        RECT 80.395 156.535 80.685 156.580 ;
        RECT 82.915 156.535 83.205 156.580 ;
        RECT 72.805 156.195 73.095 156.425 ;
        RECT 73.265 156.380 73.555 156.425 ;
        RECT 74.170 156.380 74.490 156.440 ;
        RECT 73.265 156.240 74.490 156.380 ;
        RECT 73.265 156.195 73.555 156.240 ;
        RECT 74.170 156.180 74.490 156.240 ;
        RECT 75.090 156.180 75.410 156.440 ;
        RECT 100.010 156.200 100.880 159.470 ;
        RECT 104.530 159.010 109.780 159.020 ;
        RECT 104.530 158.900 116.840 159.010 ;
        RECT 101.560 158.840 116.840 158.900 ;
        RECT 101.560 158.830 116.875 158.840 ;
        RECT 101.500 158.700 116.875 158.830 ;
        RECT 101.500 158.690 106.660 158.700 ;
        RECT 101.500 158.600 105.500 158.690 ;
        RECT 108.875 158.610 116.875 158.700 ;
        RECT 108.960 158.600 116.850 158.610 ;
        RECT 101.110 158.240 101.340 158.550 ;
        RECT 101.560 158.240 105.460 158.600 ;
        RECT 105.660 158.240 105.890 158.550 ;
        RECT 101.110 156.900 105.890 158.240 ;
        RECT 101.110 156.590 101.340 156.900 ;
        RECT 105.660 156.590 105.890 156.900 ;
        RECT 108.440 158.020 108.670 158.560 ;
        RECT 109.480 158.020 110.490 158.050 ;
        RECT 117.080 158.020 117.310 158.560 ;
        RECT 108.440 157.120 117.310 158.020 ;
        RECT 108.440 156.600 108.670 157.120 ;
        RECT 109.480 157.050 110.490 157.120 ;
        RECT 117.080 156.600 117.310 157.120 ;
        RECT 101.500 156.310 105.500 156.540 ;
        RECT 108.875 156.320 116.875 156.550 ;
        RECT 100.010 156.160 101.180 156.200 ;
        RECT 72.345 156.040 72.635 156.085 ;
        RECT 75.690 156.040 75.980 156.085 ;
        RECT 79.550 156.040 79.840 156.085 ;
        RECT 72.345 155.900 75.980 156.040 ;
        RECT 72.345 155.855 72.635 155.900 ;
        RECT 75.690 155.855 75.980 155.900 ;
        RECT 76.560 155.900 79.840 156.040 ;
        RECT 64.050 155.700 64.370 155.760 ;
        RECT 64.985 155.700 65.275 155.745 ;
        RECT 63.680 155.560 65.275 155.700 ;
        RECT 64.050 155.500 64.370 155.560 ;
        RECT 64.985 155.515 65.275 155.560 ;
        RECT 73.250 155.700 73.570 155.760 ;
        RECT 76.560 155.745 76.700 155.900 ;
        RECT 79.550 155.855 79.840 155.900 ;
        RECT 100.010 156.080 101.420 156.160 ;
        RECT 101.790 156.090 105.450 156.310 ;
        RECT 101.790 156.080 103.230 156.090 ;
        RECT 100.010 156.040 103.230 156.080 ;
        RECT 100.010 155.950 102.740 156.040 ;
        RECT 108.940 156.030 116.830 156.320 ;
        RECT 100.010 155.890 102.070 155.950 ;
        RECT 100.010 155.840 101.820 155.890 ;
        RECT 74.645 155.700 74.935 155.745 ;
        RECT 73.250 155.560 74.935 155.700 ;
        RECT 73.250 155.500 73.570 155.560 ;
        RECT 74.645 155.515 74.935 155.560 ;
        RECT 76.485 155.515 76.775 155.745 ;
        RECT 78.310 155.700 78.630 155.760 ;
        RECT 85.225 155.700 85.515 155.745 ;
        RECT 78.310 155.560 85.515 155.700 ;
        RECT 78.310 155.500 78.630 155.560 ;
        RECT 85.225 155.515 85.515 155.560 ;
        RECT 13.380 154.880 92.040 155.360 ;
        RECT 27.250 154.680 27.570 154.740 ;
        RECT 25.960 154.540 27.570 154.680 ;
        RECT 22.650 154.140 22.970 154.400 ;
        RECT 25.960 154.385 26.100 154.540 ;
        RECT 27.250 154.480 27.570 154.540 ;
        RECT 34.165 154.680 34.455 154.725 ;
        RECT 34.610 154.680 34.930 154.740 ;
        RECT 35.530 154.680 35.850 154.740 ;
        RECT 34.165 154.540 35.850 154.680 ;
        RECT 34.165 154.495 34.455 154.540 ;
        RECT 34.610 154.480 34.930 154.540 ;
        RECT 35.530 154.480 35.850 154.540 ;
        RECT 50.250 154.680 50.570 154.740 ;
        RECT 57.610 154.680 57.930 154.740 ;
        RECT 62.225 154.680 62.515 154.725 ;
        RECT 71.870 154.680 72.190 154.740 ;
        RECT 74.630 154.680 74.950 154.740 ;
        RECT 50.250 154.540 53.240 154.680 ;
        RECT 50.250 154.480 50.570 154.540 ;
        RECT 23.745 154.340 24.035 154.385 ;
        RECT 24.965 154.340 25.255 154.385 ;
        RECT 23.745 154.200 25.255 154.340 ;
        RECT 23.745 154.155 24.035 154.200 ;
        RECT 24.965 154.155 25.255 154.200 ;
        RECT 25.885 154.155 26.175 154.385 ;
        RECT 26.330 154.340 26.650 154.400 ;
        RECT 26.805 154.340 27.095 154.385 ;
        RECT 31.390 154.340 31.710 154.400 ;
        RECT 26.330 154.200 27.095 154.340 ;
        RECT 26.330 154.140 26.650 154.200 ;
        RECT 26.805 154.155 27.095 154.200 ;
        RECT 27.340 154.200 31.710 154.340 ;
        RECT 27.340 154.045 27.480 154.200 ;
        RECT 31.390 154.140 31.710 154.200 ;
        RECT 39.670 154.340 39.990 154.400 ;
        RECT 39.670 154.200 51.400 154.340 ;
        RECT 39.670 154.140 39.990 154.200 ;
        RECT 27.265 153.815 27.555 154.045 ;
        RECT 28.545 154.000 28.835 154.045 ;
        RECT 27.800 153.860 28.835 154.000 ;
        RECT 27.800 153.660 27.940 153.860 ;
        RECT 28.545 153.815 28.835 153.860 ;
        RECT 49.330 154.000 49.650 154.060 ;
        RECT 51.260 154.045 51.400 154.200 ;
        RECT 53.100 154.045 53.240 154.540 ;
        RECT 57.610 154.540 62.515 154.680 ;
        RECT 57.610 154.480 57.930 154.540 ;
        RECT 62.225 154.495 62.515 154.540 ;
        RECT 70.580 154.540 71.640 154.680 ;
        RECT 70.580 154.385 70.720 154.540 ;
        RECT 70.505 154.155 70.795 154.385 ;
        RECT 70.950 154.140 71.270 154.400 ;
        RECT 71.500 154.340 71.640 154.540 ;
        RECT 71.870 154.540 74.950 154.680 ;
        RECT 71.870 154.480 72.190 154.540 ;
        RECT 74.630 154.480 74.950 154.540 ;
        RECT 73.710 154.340 74.030 154.400 ;
        RECT 75.405 154.340 75.695 154.385 ;
        RECT 71.500 154.200 75.695 154.340 ;
        RECT 73.710 154.140 74.030 154.200 ;
        RECT 75.405 154.155 75.695 154.200 ;
        RECT 76.485 154.340 76.775 154.385 ;
        RECT 78.310 154.340 78.630 154.400 ;
        RECT 76.485 154.200 78.630 154.340 ;
        RECT 76.485 154.155 76.775 154.200 ;
        RECT 50.265 154.000 50.555 154.045 ;
        RECT 49.330 153.860 50.555 154.000 ;
        RECT 49.330 153.800 49.650 153.860 ;
        RECT 50.265 153.815 50.555 153.860 ;
        RECT 51.185 154.000 51.475 154.045 ;
        RECT 52.565 154.000 52.855 154.045 ;
        RECT 51.185 153.860 52.855 154.000 ;
        RECT 51.185 153.815 51.475 153.860 ;
        RECT 52.565 153.815 52.855 153.860 ;
        RECT 53.025 153.815 53.315 154.045 ;
        RECT 53.470 154.000 53.790 154.060 ;
        RECT 53.945 154.000 54.235 154.045 ;
        RECT 53.470 153.860 54.235 154.000 ;
        RECT 24.580 153.520 27.940 153.660 ;
        RECT 28.145 153.660 28.435 153.705 ;
        RECT 29.335 153.660 29.625 153.705 ;
        RECT 31.855 153.660 32.145 153.705 ;
        RECT 28.145 153.520 32.145 153.660 ;
        RECT 50.340 153.660 50.480 153.815 ;
        RECT 53.100 153.660 53.240 153.815 ;
        RECT 53.470 153.800 53.790 153.860 ;
        RECT 53.945 153.815 54.235 153.860 ;
        RECT 54.850 153.800 55.170 154.060 ;
        RECT 56.245 154.000 56.535 154.045 ;
        RECT 57.150 154.000 57.470 154.060 ;
        RECT 56.245 153.860 57.470 154.000 ;
        RECT 56.245 153.815 56.535 153.860 ;
        RECT 57.150 153.800 57.470 153.860 ;
        RECT 63.130 153.800 63.450 154.060 ;
        RECT 64.065 154.000 64.355 154.045 ;
        RECT 64.510 154.000 64.830 154.060 ;
        RECT 64.065 153.860 64.830 154.000 ;
        RECT 64.065 153.815 64.355 153.860 ;
        RECT 64.510 153.800 64.830 153.860 ;
        RECT 66.810 154.000 67.130 154.060 ;
        RECT 67.285 154.000 67.575 154.045 ;
        RECT 66.810 153.860 67.575 154.000 ;
        RECT 66.810 153.800 67.130 153.860 ;
        RECT 67.285 153.815 67.575 153.860 ;
        RECT 68.205 154.000 68.495 154.045 ;
        RECT 68.650 154.000 68.970 154.060 ;
        RECT 68.205 153.860 68.970 154.000 ;
        RECT 68.205 153.815 68.495 153.860 ;
        RECT 55.325 153.660 55.615 153.705 ;
        RECT 50.340 153.520 52.780 153.660 ;
        RECT 53.100 153.520 55.615 153.660 ;
        RECT 67.360 153.660 67.500 153.815 ;
        RECT 68.650 153.800 68.970 153.860 ;
        RECT 70.030 154.000 70.350 154.060 ;
        RECT 71.425 154.000 71.715 154.045 ;
        RECT 76.560 154.000 76.700 154.155 ;
        RECT 78.310 154.140 78.630 154.200 ;
        RECT 70.030 153.860 76.700 154.000 ;
        RECT 70.030 153.800 70.350 153.860 ;
        RECT 71.425 153.815 71.715 153.860 ;
        RECT 76.945 153.815 77.235 154.045 ;
        RECT 77.405 154.000 77.695 154.045 ;
        RECT 80.150 154.000 80.470 154.060 ;
        RECT 77.405 153.860 80.470 154.000 ;
        RECT 77.405 153.815 77.695 153.860 ;
        RECT 73.710 153.660 74.030 153.720 ;
        RECT 76.470 153.660 76.790 153.720 ;
        RECT 77.020 153.660 77.160 153.815 ;
        RECT 67.360 153.520 72.560 153.660 ;
        RECT 24.580 153.365 24.720 153.520 ;
        RECT 28.145 153.475 28.435 153.520 ;
        RECT 29.335 153.475 29.625 153.520 ;
        RECT 31.855 153.475 32.145 153.520 ;
        RECT 24.505 153.135 24.795 153.365 ;
        RECT 27.750 153.320 28.040 153.365 ;
        RECT 29.850 153.320 30.140 153.365 ;
        RECT 31.420 153.320 31.710 153.365 ;
        RECT 27.750 153.180 31.710 153.320 ;
        RECT 27.750 153.135 28.040 153.180 ;
        RECT 29.850 153.135 30.140 153.180 ;
        RECT 31.420 153.135 31.710 153.180 ;
        RECT 35.990 153.320 36.310 153.380 ;
        RECT 39.210 153.320 39.530 153.380 ;
        RECT 52.640 153.320 52.780 153.520 ;
        RECT 55.325 153.475 55.615 153.520 ;
        RECT 53.485 153.320 53.775 153.365 ;
        RECT 54.390 153.320 54.710 153.380 ;
        RECT 55.770 153.320 56.090 153.380 ;
        RECT 70.030 153.320 70.350 153.380 ;
        RECT 72.420 153.365 72.560 153.520 ;
        RECT 73.710 153.520 77.160 153.660 ;
        RECT 73.710 153.460 74.030 153.520 ;
        RECT 76.470 153.460 76.790 153.520 ;
        RECT 35.990 153.180 52.320 153.320 ;
        RECT 52.640 153.180 54.710 153.320 ;
        RECT 35.990 153.120 36.310 153.180 ;
        RECT 39.210 153.120 39.530 153.180 ;
        RECT 23.570 152.780 23.890 153.040 ;
        RECT 50.250 152.780 50.570 153.040 ;
        RECT 51.630 152.780 51.950 153.040 ;
        RECT 52.180 152.980 52.320 153.180 ;
        RECT 53.485 153.135 53.775 153.180 ;
        RECT 54.390 153.120 54.710 153.180 ;
        RECT 54.940 153.180 56.090 153.320 ;
        RECT 54.940 153.025 55.080 153.180 ;
        RECT 55.770 153.120 56.090 153.180 ;
        RECT 68.280 153.180 70.350 153.320 ;
        RECT 54.865 152.980 55.155 153.025 ;
        RECT 52.180 152.840 55.155 152.980 ;
        RECT 54.865 152.795 55.155 152.840 ;
        RECT 55.310 152.980 55.630 153.040 ;
        RECT 57.165 152.980 57.455 153.025 ;
        RECT 55.310 152.840 57.455 152.980 ;
        RECT 55.310 152.780 55.630 152.840 ;
        RECT 57.165 152.795 57.455 152.840 ;
        RECT 64.050 152.780 64.370 153.040 ;
        RECT 64.970 152.980 65.290 153.040 ;
        RECT 68.280 153.025 68.420 153.180 ;
        RECT 70.030 153.120 70.350 153.180 ;
        RECT 72.345 153.320 72.635 153.365 ;
        RECT 76.010 153.320 76.330 153.380 ;
        RECT 72.345 153.180 76.330 153.320 ;
        RECT 72.345 153.135 72.635 153.180 ;
        RECT 76.010 153.120 76.330 153.180 ;
        RECT 66.365 152.980 66.655 153.025 ;
        RECT 64.970 152.840 66.655 152.980 ;
        RECT 64.970 152.780 65.290 152.840 ;
        RECT 66.365 152.795 66.655 152.840 ;
        RECT 68.205 152.795 68.495 153.025 ;
        RECT 69.570 152.780 69.890 153.040 ;
        RECT 70.950 152.980 71.270 153.040 ;
        RECT 75.565 152.980 75.855 153.025 ;
        RECT 77.480 152.980 77.620 153.815 ;
        RECT 80.150 153.800 80.470 153.860 ;
        RECT 77.850 153.320 78.170 153.380 ;
        RECT 78.325 153.320 78.615 153.365 ;
        RECT 77.850 153.180 78.615 153.320 ;
        RECT 77.850 153.120 78.170 153.180 ;
        RECT 78.325 153.135 78.615 153.180 ;
        RECT 70.950 152.840 77.620 152.980 ;
        RECT 70.950 152.780 71.270 152.840 ;
        RECT 75.565 152.795 75.855 152.840 ;
        RECT 13.380 152.160 92.040 152.640 ;
        RECT 100.010 152.500 100.880 155.840 ;
        RECT 108.930 155.540 116.850 155.550 ;
        RECT 105.160 155.530 116.850 155.540 ;
        RECT 101.540 155.410 116.850 155.530 ;
        RECT 101.540 155.400 116.875 155.410 ;
        RECT 101.500 155.280 116.875 155.400 ;
        RECT 101.500 155.170 105.500 155.280 ;
        RECT 101.110 154.830 101.340 155.120 ;
        RECT 101.560 154.830 105.450 155.170 ;
        RECT 105.660 154.830 105.890 155.120 ;
        RECT 101.110 153.460 105.890 154.830 ;
        RECT 101.110 153.160 101.340 153.460 ;
        RECT 105.660 153.160 105.890 153.460 ;
        RECT 101.500 152.880 105.500 153.110 ;
        RECT 101.750 152.650 105.320 152.880 ;
        RECT 101.750 152.500 105.440 152.650 ;
        RECT 100.010 152.220 105.440 152.500 ;
        RECT 106.690 152.330 107.310 155.280 ;
        RECT 108.875 155.180 116.875 155.280 ;
        RECT 108.930 155.170 116.850 155.180 ;
        RECT 108.440 154.470 108.670 155.130 ;
        RECT 109.450 154.470 110.450 154.560 ;
        RECT 117.080 154.470 117.310 155.130 ;
        RECT 108.440 153.650 117.310 154.470 ;
        RECT 108.440 153.170 108.670 153.650 ;
        RECT 109.450 153.560 110.450 153.650 ;
        RECT 117.080 153.170 117.310 153.650 ;
        RECT 108.875 152.890 116.875 153.120 ;
        RECT 50.250 151.760 50.570 152.020 ;
        RECT 59.910 151.960 60.230 152.020 ;
        RECT 64.050 151.960 64.370 152.020 ;
        RECT 64.525 151.960 64.815 152.005 ;
        RECT 59.910 151.820 63.820 151.960 ;
        RECT 59.910 151.760 60.230 151.820 ;
        RECT 19.470 151.620 19.760 151.665 ;
        RECT 21.570 151.620 21.860 151.665 ;
        RECT 23.140 151.620 23.430 151.665 ;
        RECT 19.470 151.480 23.430 151.620 ;
        RECT 19.470 151.435 19.760 151.480 ;
        RECT 21.570 151.435 21.860 151.480 ;
        RECT 23.140 151.435 23.430 151.480 ;
        RECT 37.385 151.620 37.675 151.665 ;
        RECT 54.850 151.620 55.170 151.680 ;
        RECT 63.680 151.620 63.820 151.820 ;
        RECT 64.050 151.820 64.815 151.960 ;
        RECT 64.050 151.760 64.370 151.820 ;
        RECT 64.525 151.775 64.815 151.820 ;
        RECT 100.010 151.760 105.450 152.220 ;
        RECT 72.330 151.620 72.650 151.680 ;
        RECT 73.710 151.620 74.030 151.680 ;
        RECT 37.385 151.480 45.420 151.620 ;
        RECT 37.385 151.435 37.675 151.480 ;
        RECT 19.865 151.280 20.155 151.325 ;
        RECT 21.055 151.280 21.345 151.325 ;
        RECT 23.575 151.280 23.865 151.325 ;
        RECT 19.865 151.140 23.865 151.280 ;
        RECT 19.865 151.095 20.155 151.140 ;
        RECT 21.055 151.095 21.345 151.140 ;
        RECT 23.575 151.095 23.865 151.140 ;
        RECT 26.330 151.280 26.650 151.340 ;
        RECT 31.390 151.280 31.710 151.340 ;
        RECT 36.910 151.280 37.230 151.340 ;
        RECT 26.330 151.140 29.320 151.280 ;
        RECT 26.330 151.080 26.650 151.140 ;
        RECT 18.970 150.740 19.290 151.000 ;
        RECT 29.180 150.985 29.320 151.140 ;
        RECT 31.390 151.140 33.005 151.280 ;
        RECT 31.390 151.080 31.710 151.140 ;
        RECT 32.865 150.985 33.005 151.140 ;
        RECT 33.780 151.140 37.230 151.280 ;
        RECT 33.780 150.985 33.920 151.140 ;
        RECT 36.910 151.080 37.230 151.140 ;
        RECT 27.725 150.755 28.015 150.985 ;
        RECT 29.105 150.755 29.395 150.985 ;
        RECT 32.325 150.755 32.615 150.985 ;
        RECT 32.790 150.755 33.080 150.985 ;
        RECT 33.705 150.755 33.995 150.985 ;
        RECT 34.855 150.940 35.145 150.985 ;
        RECT 37.460 150.940 37.600 151.435 ;
        RECT 41.525 151.095 41.815 151.325 ;
        RECT 34.855 150.800 37.600 150.940 ;
        RECT 34.855 150.755 35.145 150.800 ;
        RECT 20.350 150.645 20.670 150.660 ;
        RECT 20.320 150.415 20.670 150.645 ;
        RECT 27.800 150.600 27.940 150.755 ;
        RECT 32.400 150.600 32.540 150.755 ;
        RECT 38.750 150.740 39.070 151.000 ;
        RECT 39.210 150.740 39.530 151.000 ;
        RECT 39.670 150.940 39.990 151.000 ;
        RECT 41.065 150.940 41.355 150.985 ;
        RECT 39.670 150.800 41.355 150.940 ;
        RECT 41.600 150.940 41.740 151.095 ;
        RECT 42.890 151.080 43.210 151.340 ;
        RECT 45.280 151.325 45.420 151.480 ;
        RECT 50.340 151.480 55.170 151.620 ;
        RECT 50.340 151.325 50.480 151.480 ;
        RECT 54.850 151.420 55.170 151.480 ;
        RECT 59.540 151.480 63.360 151.620 ;
        RECT 63.680 151.480 74.030 151.620 ;
        RECT 45.205 151.095 45.495 151.325 ;
        RECT 50.265 151.095 50.555 151.325 ;
        RECT 51.630 151.280 51.950 151.340 ;
        RECT 56.705 151.280 56.995 151.325 ;
        RECT 51.630 151.140 56.995 151.280 ;
        RECT 51.630 151.080 51.950 151.140 ;
        RECT 56.705 151.095 56.995 151.140 ;
        RECT 41.970 150.940 42.290 151.000 ;
        RECT 44.730 150.940 45.050 151.000 ;
        RECT 41.600 150.800 45.050 150.940 ;
        RECT 39.670 150.740 39.990 150.800 ;
        RECT 41.065 150.755 41.355 150.800 ;
        RECT 41.970 150.740 42.290 150.800 ;
        RECT 44.730 150.740 45.050 150.800 ;
        RECT 45.665 150.940 45.955 150.985 ;
        RECT 45.665 150.800 50.480 150.940 ;
        RECT 45.665 150.755 45.955 150.800 ;
        RECT 20.350 150.400 20.670 150.415 ;
        RECT 25.960 150.460 32.540 150.600 ;
        RECT 34.165 150.600 34.455 150.645 ;
        RECT 34.165 150.460 34.840 150.600 ;
        RECT 25.960 150.320 26.100 150.460 ;
        RECT 34.165 150.415 34.455 150.460 ;
        RECT 34.700 150.320 34.840 150.460 ;
        RECT 49.345 150.415 49.635 150.645 ;
        RECT 50.340 150.600 50.480 150.800 ;
        RECT 50.710 150.740 51.030 151.000 ;
        RECT 53.025 150.940 53.315 150.985 ;
        RECT 51.260 150.800 53.315 150.940 ;
        RECT 51.260 150.660 51.400 150.800 ;
        RECT 53.025 150.755 53.315 150.800 ;
        RECT 55.310 150.740 55.630 151.000 ;
        RECT 58.545 150.940 58.835 150.985 ;
        RECT 59.540 150.940 59.680 151.480 ;
        RECT 59.910 151.080 60.230 151.340 ;
        RECT 61.290 150.985 61.610 151.000 ;
        RECT 58.545 150.800 59.680 150.940 ;
        RECT 58.545 150.755 58.835 150.800 ;
        RECT 60.385 150.755 60.675 150.985 ;
        RECT 61.125 150.755 61.610 150.985 ;
        RECT 51.170 150.600 51.490 150.660 ;
        RECT 58.990 150.600 59.310 150.660 ;
        RECT 60.460 150.600 60.600 150.755 ;
        RECT 61.290 150.740 61.610 150.755 ;
        RECT 61.750 150.740 62.070 151.000 ;
        RECT 62.710 150.755 63.000 150.985 ;
        RECT 63.220 150.940 63.360 151.480 ;
        RECT 72.330 151.420 72.650 151.480 ;
        RECT 73.710 151.420 74.030 151.480 ;
        RECT 75.565 151.280 75.855 151.325 ;
        RECT 74.720 151.140 75.855 151.280 ;
        RECT 63.220 150.800 63.820 150.940 ;
        RECT 50.340 150.460 51.490 150.600 ;
        RECT 25.870 150.060 26.190 150.320 ;
        RECT 26.790 150.060 27.110 150.320 ;
        RECT 27.250 150.260 27.570 150.320 ;
        RECT 28.645 150.260 28.935 150.305 ;
        RECT 34.610 150.260 34.930 150.320 ;
        RECT 27.250 150.120 34.930 150.260 ;
        RECT 27.250 150.060 27.570 150.120 ;
        RECT 28.645 150.075 28.935 150.120 ;
        RECT 34.610 150.060 34.930 150.120 ;
        RECT 35.530 150.060 35.850 150.320 ;
        RECT 47.505 150.260 47.795 150.305 ;
        RECT 49.420 150.260 49.560 150.415 ;
        RECT 51.170 150.400 51.490 150.460 ;
        RECT 51.720 150.460 60.600 150.600 ;
        RECT 51.720 150.305 51.860 150.460 ;
        RECT 58.990 150.400 59.310 150.460 ;
        RECT 62.210 150.400 62.530 150.660 ;
        RECT 47.505 150.120 49.560 150.260 ;
        RECT 47.505 150.075 47.795 150.120 ;
        RECT 51.645 150.075 51.935 150.305 ;
        RECT 53.490 150.260 53.780 150.305 ;
        RECT 59.930 150.260 60.220 150.305 ;
        RECT 53.490 150.120 60.220 150.260 ;
        RECT 53.490 150.075 53.780 150.120 ;
        RECT 59.930 150.075 60.220 150.120 ;
        RECT 60.830 150.260 61.150 150.320 ;
        RECT 62.760 150.260 62.900 150.755 ;
        RECT 63.680 150.305 63.820 150.800 ;
        RECT 64.065 150.755 64.355 150.985 ;
        RECT 64.985 150.940 65.275 150.985 ;
        RECT 67.730 150.940 68.050 151.000 ;
        RECT 64.985 150.800 68.050 150.940 ;
        RECT 64.985 150.755 65.275 150.800 ;
        RECT 64.140 150.600 64.280 150.755 ;
        RECT 67.730 150.740 68.050 150.800 ;
        RECT 69.570 150.940 69.890 151.000 ;
        RECT 74.720 150.985 74.860 151.140 ;
        RECT 75.565 151.095 75.855 151.140 ;
        RECT 73.725 150.940 74.015 150.985 ;
        RECT 69.570 150.800 74.015 150.940 ;
        RECT 69.570 150.740 69.890 150.800 ;
        RECT 73.725 150.755 74.015 150.800 ;
        RECT 74.645 150.755 74.935 150.985 ;
        RECT 75.090 150.740 75.410 151.000 ;
        RECT 76.010 150.940 76.330 151.000 ;
        RECT 81.990 150.940 82.310 151.000 ;
        RECT 76.010 150.800 82.310 150.940 ;
        RECT 76.010 150.740 76.330 150.800 ;
        RECT 81.990 150.740 82.310 150.800 ;
        RECT 65.890 150.600 66.210 150.660 ;
        RECT 68.650 150.600 68.970 150.660 ;
        RECT 64.140 150.460 68.970 150.600 ;
        RECT 65.890 150.400 66.210 150.460 ;
        RECT 68.650 150.400 68.970 150.460 ;
        RECT 100.010 150.410 102.050 151.760 ;
        RECT 103.800 151.750 105.450 151.760 ;
        RECT 102.490 150.480 103.490 151.200 ;
        RECT 103.800 150.940 104.110 151.750 ;
        RECT 104.570 151.470 105.450 151.750 ;
        RECT 105.690 151.930 107.310 152.330 ;
        RECT 108.960 151.980 116.830 152.890 ;
        RECT 104.510 151.240 105.510 151.470 ;
        RECT 105.690 151.280 106.040 151.930 ;
        RECT 106.690 151.920 107.310 151.930 ;
        RECT 108.875 151.750 116.875 151.980 ;
        RECT 108.960 151.740 116.830 151.750 ;
        RECT 104.570 151.030 105.450 151.050 ;
        RECT 103.840 150.650 104.110 150.940 ;
        RECT 104.510 150.800 105.510 151.030 ;
        RECT 105.670 150.990 106.040 151.280 ;
        RECT 105.700 150.930 106.040 150.990 ;
        RECT 106.800 151.600 107.560 151.650 ;
        RECT 108.440 151.600 108.670 151.700 ;
        RECT 106.800 151.390 108.670 151.600 ;
        RECT 117.080 151.390 117.310 151.700 ;
        RECT 106.800 150.970 109.340 151.390 ;
        RECT 116.710 150.970 117.310 151.390 ;
        RECT 104.570 150.650 105.450 150.800 ;
        RECT 104.580 150.480 105.310 150.650 ;
        RECT 60.830 150.120 62.900 150.260 ;
        RECT 60.830 150.060 61.150 150.120 ;
        RECT 63.605 150.075 63.895 150.305 ;
        RECT 72.330 150.260 72.650 150.320 ;
        RECT 74.185 150.260 74.475 150.305 ;
        RECT 72.330 150.120 74.475 150.260 ;
        RECT 72.330 150.060 72.650 150.120 ;
        RECT 74.185 150.075 74.475 150.120 ;
        RECT 13.380 149.440 92.040 149.920 ;
        RECT 20.350 149.040 20.670 149.300 ;
        RECT 21.285 149.240 21.575 149.285 ;
        RECT 22.650 149.240 22.970 149.300 ;
        RECT 21.285 149.100 22.970 149.240 ;
        RECT 21.285 149.055 21.575 149.100 ;
        RECT 22.650 149.040 22.970 149.100 ;
        RECT 24.885 149.240 25.175 149.285 ;
        RECT 26.330 149.240 26.650 149.300 ;
        RECT 24.885 149.100 26.650 149.240 ;
        RECT 24.885 149.055 25.175 149.100 ;
        RECT 26.330 149.040 26.650 149.100 ;
        RECT 31.390 149.240 31.710 149.300 ;
        RECT 39.670 149.240 39.990 149.300 ;
        RECT 49.805 149.240 50.095 149.285 ;
        RECT 31.390 149.100 39.440 149.240 ;
        RECT 31.390 149.040 31.710 149.100 ;
        RECT 25.870 148.700 26.190 148.960 ;
        RECT 35.530 148.900 35.850 148.960 ;
        RECT 33.320 148.760 35.850 148.900 ;
        RECT 39.300 148.900 39.440 149.100 ;
        RECT 39.670 149.100 50.095 149.240 ;
        RECT 39.670 149.040 39.990 149.100 ;
        RECT 49.805 149.055 50.095 149.100 ;
        RECT 51.645 149.240 51.935 149.285 ;
        RECT 54.850 149.240 55.170 149.300 ;
        RECT 51.645 149.100 55.170 149.240 ;
        RECT 51.645 149.055 51.935 149.100 ;
        RECT 54.850 149.040 55.170 149.100 ;
        RECT 60.830 149.040 61.150 149.300 ;
        RECT 61.290 149.040 61.610 149.300 ;
        RECT 72.790 149.240 73.110 149.300 ;
        RECT 73.265 149.240 73.555 149.285 ;
        RECT 72.790 149.100 73.555 149.240 ;
        RECT 72.790 149.040 73.110 149.100 ;
        RECT 73.265 149.055 73.555 149.100 ;
        RECT 74.645 149.055 74.935 149.285 ;
        RECT 64.970 148.900 65.290 148.960 ;
        RECT 39.300 148.760 49.100 148.900 ;
        RECT 31.850 148.360 32.170 148.620 ;
        RECT 32.310 148.560 32.630 148.620 ;
        RECT 33.320 148.605 33.460 148.760 ;
        RECT 35.530 148.700 35.850 148.760 ;
        RECT 32.785 148.560 33.075 148.605 ;
        RECT 32.310 148.420 33.075 148.560 ;
        RECT 32.310 148.360 32.630 148.420 ;
        RECT 32.785 148.375 33.075 148.420 ;
        RECT 33.245 148.375 33.535 148.605 ;
        RECT 34.610 148.360 34.930 148.620 ;
        RECT 43.810 148.560 44.130 148.620 ;
        RECT 45.250 148.560 45.540 148.605 ;
        RECT 43.810 148.420 45.540 148.560 ;
        RECT 48.960 148.560 49.100 148.760 ;
        RECT 63.680 148.760 65.290 148.900 ;
        RECT 49.330 148.560 49.650 148.620 ;
        RECT 48.960 148.420 49.650 148.560 ;
        RECT 43.810 148.360 44.130 148.420 ;
        RECT 45.250 148.375 45.540 148.420 ;
        RECT 49.330 148.360 49.650 148.420 ;
        RECT 50.250 148.560 50.570 148.620 ;
        RECT 50.725 148.560 51.015 148.605 ;
        RECT 50.250 148.420 51.015 148.560 ;
        RECT 50.250 148.360 50.570 148.420 ;
        RECT 50.725 148.375 51.015 148.420 ;
        RECT 58.990 148.360 59.310 148.620 ;
        RECT 59.925 148.560 60.215 148.605 ;
        RECT 60.830 148.560 61.150 148.620 ;
        RECT 63.680 148.605 63.820 148.760 ;
        RECT 64.970 148.700 65.290 148.760 ;
        RECT 65.445 148.715 65.735 148.945 ;
        RECT 66.350 148.900 66.670 148.960 ;
        RECT 69.125 148.900 69.415 148.945 ;
        RECT 71.410 148.900 71.730 148.960 ;
        RECT 66.350 148.760 67.500 148.900 ;
        RECT 62.685 148.560 62.975 148.605 ;
        RECT 59.925 148.420 62.975 148.560 ;
        RECT 59.925 148.375 60.215 148.420 ;
        RECT 60.830 148.360 61.150 148.420 ;
        RECT 62.685 148.375 62.975 148.420 ;
        RECT 63.145 148.375 63.435 148.605 ;
        RECT 63.605 148.375 63.895 148.605 ;
        RECT 64.525 148.560 64.815 148.605 ;
        RECT 65.520 148.560 65.660 148.715 ;
        RECT 66.350 148.700 66.670 148.760 ;
        RECT 64.525 148.420 65.660 148.560 ;
        RECT 64.525 148.375 64.815 148.420 ;
        RECT 33.800 148.220 34.090 148.265 ;
        RECT 35.070 148.220 35.390 148.280 ;
        RECT 33.800 148.080 35.390 148.220 ;
        RECT 33.800 148.035 34.090 148.080 ;
        RECT 35.070 148.020 35.390 148.080 ;
        RECT 41.995 148.220 42.285 148.265 ;
        RECT 44.515 148.220 44.805 148.265 ;
        RECT 45.705 148.220 45.995 148.265 ;
        RECT 41.995 148.080 45.995 148.220 ;
        RECT 41.995 148.035 42.285 148.080 ;
        RECT 44.515 148.035 44.805 148.080 ;
        RECT 45.705 148.035 45.995 148.080 ;
        RECT 46.570 148.020 46.890 148.280 ;
        RECT 59.080 148.220 59.220 148.360 ;
        RECT 63.220 148.220 63.360 148.375 ;
        RECT 66.810 148.360 67.130 148.620 ;
        RECT 67.360 148.605 67.500 148.760 ;
        RECT 67.820 148.760 69.415 148.900 ;
        RECT 67.820 148.620 67.960 148.760 ;
        RECT 69.125 148.715 69.415 148.760 ;
        RECT 70.580 148.760 71.730 148.900 ;
        RECT 74.720 148.900 74.860 149.055 ;
        RECT 81.990 149.040 82.310 149.300 ;
        RECT 76.330 148.900 76.620 148.945 ;
        RECT 74.720 148.760 76.620 148.900 ;
        RECT 67.285 148.375 67.575 148.605 ;
        RECT 67.730 148.360 68.050 148.620 ;
        RECT 68.650 148.360 68.970 148.620 ;
        RECT 70.580 148.605 70.720 148.760 ;
        RECT 71.410 148.700 71.730 148.760 ;
        RECT 76.330 148.715 76.620 148.760 ;
        RECT 70.500 148.375 70.790 148.605 ;
        RECT 70.965 148.375 71.255 148.605 ;
        RECT 71.870 148.560 72.190 148.620 ;
        RECT 72.805 148.560 73.095 148.605 ;
        RECT 73.250 148.560 73.570 148.620 ;
        RECT 71.870 148.420 73.570 148.560 ;
        RECT 59.080 148.080 63.360 148.220 ;
        RECT 68.190 148.220 68.510 148.280 ;
        RECT 71.040 148.220 71.180 148.375 ;
        RECT 71.870 148.360 72.190 148.420 ;
        RECT 72.805 148.375 73.095 148.420 ;
        RECT 73.250 148.360 73.570 148.420 ;
        RECT 68.190 148.080 71.180 148.220 ;
        RECT 68.190 148.020 68.510 148.080 ;
        RECT 71.410 148.020 71.730 148.280 ;
        RECT 72.330 148.220 72.650 148.280 ;
        RECT 73.850 148.220 74.140 148.265 ;
        RECT 72.330 148.080 74.140 148.220 ;
        RECT 72.330 148.020 72.650 148.080 ;
        RECT 73.850 148.035 74.140 148.080 ;
        RECT 75.090 148.020 75.410 148.280 ;
        RECT 75.985 148.220 76.275 148.265 ;
        RECT 77.175 148.220 77.465 148.265 ;
        RECT 79.695 148.220 79.985 148.265 ;
        RECT 75.985 148.080 79.985 148.220 ;
        RECT 75.985 148.035 76.275 148.080 ;
        RECT 77.175 148.035 77.465 148.080 ;
        RECT 79.695 148.035 79.985 148.080 ;
        RECT 23.125 147.880 23.415 147.925 ;
        RECT 24.030 147.880 24.350 147.940 ;
        RECT 26.790 147.880 27.110 147.940 ;
        RECT 23.125 147.740 24.350 147.880 ;
        RECT 23.125 147.695 23.415 147.740 ;
        RECT 24.030 147.680 24.350 147.740 ;
        RECT 24.580 147.740 27.110 147.880 ;
        RECT 21.285 147.540 21.575 147.585 ;
        RECT 24.580 147.540 24.720 147.740 ;
        RECT 26.790 147.680 27.110 147.740 ;
        RECT 32.325 147.880 32.615 147.925 ;
        RECT 41.510 147.880 41.830 147.940 ;
        RECT 32.325 147.740 41.830 147.880 ;
        RECT 32.325 147.695 32.615 147.740 ;
        RECT 41.510 147.680 41.830 147.740 ;
        RECT 42.430 147.880 42.720 147.925 ;
        RECT 44.000 147.880 44.290 147.925 ;
        RECT 46.100 147.880 46.390 147.925 ;
        RECT 42.430 147.740 46.390 147.880 ;
        RECT 42.430 147.695 42.720 147.740 ;
        RECT 44.000 147.695 44.290 147.740 ;
        RECT 46.100 147.695 46.390 147.740 ;
        RECT 75.590 147.880 75.880 147.925 ;
        RECT 77.690 147.880 77.980 147.925 ;
        RECT 79.260 147.880 79.550 147.925 ;
        RECT 75.590 147.740 79.550 147.880 ;
        RECT 75.590 147.695 75.880 147.740 ;
        RECT 77.690 147.695 77.980 147.740 ;
        RECT 79.260 147.695 79.550 147.740 ;
        RECT 21.285 147.400 24.720 147.540 ;
        RECT 24.965 147.540 25.255 147.585 ;
        RECT 27.250 147.540 27.570 147.600 ;
        RECT 24.965 147.400 27.570 147.540 ;
        RECT 21.285 147.355 21.575 147.400 ;
        RECT 24.965 147.355 25.255 147.400 ;
        RECT 27.250 147.340 27.570 147.400 ;
        RECT 13.380 146.720 92.040 147.200 ;
        RECT 100.010 146.720 100.780 150.410 ;
        RECT 102.460 149.360 105.310 150.480 ;
        RECT 105.700 150.180 106.050 150.930 ;
        RECT 106.800 150.810 108.670 150.970 ;
        RECT 106.800 150.760 107.560 150.810 ;
        RECT 108.440 150.740 108.670 150.810 ;
        RECT 117.080 150.740 117.310 150.970 ;
        RECT 108.875 150.460 116.875 150.690 ;
        RECT 105.700 150.120 105.990 150.180 ;
        RECT 105.610 150.000 105.990 150.120 ;
        RECT 108.970 150.060 116.830 150.460 ;
        RECT 117.640 150.060 118.600 159.540 ;
        RECT 119.930 159.670 120.770 161.800 ;
        RECT 126.430 161.380 127.680 161.820 ;
        RECT 137.600 161.800 138.460 163.870 ;
        RECT 124.370 161.370 129.610 161.380 ;
        RECT 121.420 161.270 136.720 161.370 ;
        RECT 121.420 161.260 136.755 161.270 ;
        RECT 121.380 161.140 136.755 161.260 ;
        RECT 121.380 161.030 125.380 161.140 ;
        RECT 126.430 161.060 128.170 161.140 ;
        RECT 128.750 161.060 136.755 161.140 ;
        RECT 126.430 160.980 127.680 161.060 ;
        RECT 128.755 161.040 136.755 161.060 ;
        RECT 120.990 160.730 121.220 160.980 ;
        RECT 125.540 160.840 125.770 160.980 ;
        RECT 128.320 160.840 128.550 160.990 ;
        RECT 125.540 160.730 128.550 160.840 ;
        RECT 136.960 160.730 137.190 160.990 ;
        RECT 120.990 160.290 137.190 160.730 ;
        RECT 120.990 160.020 121.220 160.290 ;
        RECT 125.540 160.260 137.190 160.290 ;
        RECT 125.540 160.170 128.550 160.260 ;
        RECT 125.540 160.020 125.770 160.170 ;
        RECT 128.320 160.030 128.550 160.170 ;
        RECT 136.960 160.030 137.190 160.260 ;
        RECT 121.380 159.740 125.380 159.970 ;
        RECT 128.755 159.760 136.755 159.980 ;
        RECT 137.520 159.760 138.480 161.800 ;
        RECT 128.755 159.750 138.480 159.760 ;
        RECT 121.380 159.670 125.370 159.740 ;
        RECT 119.930 159.560 125.370 159.670 ;
        RECT 128.810 159.590 138.480 159.750 ;
        RECT 119.930 159.470 123.060 159.560 ;
        RECT 136.550 159.540 138.480 159.590 ;
        RECT 119.930 156.200 120.770 159.470 ;
        RECT 124.410 159.010 129.660 159.020 ;
        RECT 124.410 158.900 136.720 159.010 ;
        RECT 121.440 158.840 136.720 158.900 ;
        RECT 121.440 158.830 136.755 158.840 ;
        RECT 121.380 158.700 136.755 158.830 ;
        RECT 121.380 158.690 126.540 158.700 ;
        RECT 121.380 158.600 125.380 158.690 ;
        RECT 128.755 158.610 136.755 158.700 ;
        RECT 128.840 158.600 136.730 158.610 ;
        RECT 120.990 158.240 121.220 158.550 ;
        RECT 121.440 158.240 125.340 158.600 ;
        RECT 125.540 158.240 125.770 158.550 ;
        RECT 120.990 156.900 125.770 158.240 ;
        RECT 120.990 156.590 121.220 156.900 ;
        RECT 125.540 156.590 125.770 156.900 ;
        RECT 128.320 158.020 128.550 158.560 ;
        RECT 129.360 158.020 130.370 158.050 ;
        RECT 136.960 158.020 137.190 158.560 ;
        RECT 128.320 157.120 137.190 158.020 ;
        RECT 128.320 156.600 128.550 157.120 ;
        RECT 129.360 157.050 130.370 157.120 ;
        RECT 136.960 156.600 137.190 157.120 ;
        RECT 121.380 156.310 125.380 156.540 ;
        RECT 128.755 156.320 136.755 156.550 ;
        RECT 119.930 156.160 121.060 156.200 ;
        RECT 119.930 156.080 121.300 156.160 ;
        RECT 121.670 156.090 125.330 156.310 ;
        RECT 121.670 156.080 123.110 156.090 ;
        RECT 119.930 156.040 123.110 156.080 ;
        RECT 119.930 155.950 122.620 156.040 ;
        RECT 128.820 156.030 136.710 156.320 ;
        RECT 119.930 155.890 121.950 155.950 ;
        RECT 119.930 155.840 121.700 155.890 ;
        RECT 119.930 152.500 120.770 155.840 ;
        RECT 128.810 155.540 136.730 155.550 ;
        RECT 125.040 155.530 136.730 155.540 ;
        RECT 121.420 155.410 136.730 155.530 ;
        RECT 121.420 155.400 136.755 155.410 ;
        RECT 121.380 155.280 136.755 155.400 ;
        RECT 121.380 155.170 125.380 155.280 ;
        RECT 120.990 154.830 121.220 155.120 ;
        RECT 121.440 154.830 125.330 155.170 ;
        RECT 125.540 154.830 125.770 155.120 ;
        RECT 120.990 153.460 125.770 154.830 ;
        RECT 120.990 153.160 121.220 153.460 ;
        RECT 125.540 153.160 125.770 153.460 ;
        RECT 121.380 152.880 125.380 153.110 ;
        RECT 121.630 152.650 125.200 152.880 ;
        RECT 121.630 152.500 125.320 152.650 ;
        RECT 119.930 152.220 125.320 152.500 ;
        RECT 126.570 152.330 127.190 155.280 ;
        RECT 128.755 155.180 136.755 155.280 ;
        RECT 128.810 155.170 136.730 155.180 ;
        RECT 128.320 154.470 128.550 155.130 ;
        RECT 129.330 154.470 130.330 154.560 ;
        RECT 136.960 154.470 137.190 155.130 ;
        RECT 128.320 153.650 137.190 154.470 ;
        RECT 128.320 153.170 128.550 153.650 ;
        RECT 129.330 153.560 130.330 153.650 ;
        RECT 136.960 153.170 137.190 153.650 ;
        RECT 128.755 152.890 136.755 153.120 ;
        RECT 119.930 151.760 125.330 152.220 ;
        RECT 119.930 150.420 121.930 151.760 ;
        RECT 123.680 151.750 125.330 151.760 ;
        RECT 122.370 150.480 123.370 151.200 ;
        RECT 123.680 150.940 123.990 151.750 ;
        RECT 124.450 151.470 125.330 151.750 ;
        RECT 125.570 151.930 127.190 152.330 ;
        RECT 128.840 151.980 136.710 152.890 ;
        RECT 124.390 151.240 125.390 151.470 ;
        RECT 125.570 151.280 125.920 151.930 ;
        RECT 126.570 151.920 127.190 151.930 ;
        RECT 128.755 151.750 136.755 151.980 ;
        RECT 128.840 151.740 136.710 151.750 ;
        RECT 124.450 151.030 125.330 151.050 ;
        RECT 123.720 150.650 123.990 150.940 ;
        RECT 124.390 150.800 125.390 151.030 ;
        RECT 125.550 150.990 125.920 151.280 ;
        RECT 125.580 150.930 125.920 150.990 ;
        RECT 126.680 151.600 127.440 151.650 ;
        RECT 128.320 151.600 128.550 151.700 ;
        RECT 126.680 151.390 128.550 151.600 ;
        RECT 136.960 151.390 137.190 151.700 ;
        RECT 126.680 150.970 129.220 151.390 ;
        RECT 136.590 150.970 137.190 151.390 ;
        RECT 124.450 150.650 125.330 150.800 ;
        RECT 124.460 150.480 125.190 150.650 ;
        RECT 102.400 149.130 105.400 149.360 ;
        RECT 105.610 149.170 105.950 150.000 ;
        RECT 107.960 149.990 118.600 150.060 ;
        RECT 102.450 149.100 105.310 149.130 ;
        RECT 102.450 149.080 103.620 149.100 ;
        RECT 104.580 149.090 105.310 149.100 ;
        RECT 102.400 148.690 105.400 148.920 ;
        RECT 105.605 148.880 105.950 149.170 ;
        RECT 106.140 148.950 118.600 149.990 ;
        RECT 120.000 150.410 121.930 150.420 ;
        RECT 106.140 148.930 118.560 148.950 ;
        RECT 105.610 148.770 105.950 148.880 ;
        RECT 106.180 148.920 111.850 148.930 ;
        RECT 112.850 148.920 118.560 148.930 ;
        RECT 102.490 148.520 105.350 148.690 ;
        RECT 106.180 148.520 106.610 148.920 ;
        RECT 102.460 148.150 106.610 148.520 ;
        RECT 30.485 146.520 30.775 146.565 ;
        RECT 31.850 146.520 32.170 146.580 ;
        RECT 30.485 146.380 32.170 146.520 ;
        RECT 30.485 146.335 30.775 146.380 ;
        RECT 31.850 146.320 32.170 146.380 ;
        RECT 36.910 146.520 37.230 146.580 ;
        RECT 38.765 146.520 39.055 146.565 ;
        RECT 36.910 146.380 39.055 146.520 ;
        RECT 36.910 146.320 37.230 146.380 ;
        RECT 38.765 146.335 39.055 146.380 ;
        RECT 43.810 146.320 44.130 146.580 ;
        RECT 58.990 146.520 59.310 146.580 ;
        RECT 60.385 146.520 60.675 146.565 ;
        RECT 61.305 146.520 61.595 146.565 ;
        RECT 58.990 146.380 61.595 146.520 ;
        RECT 58.990 146.320 59.310 146.380 ;
        RECT 60.385 146.335 60.675 146.380 ;
        RECT 61.305 146.335 61.595 146.380 ;
        RECT 63.130 146.520 63.450 146.580 ;
        RECT 63.605 146.520 63.895 146.565 ;
        RECT 63.130 146.380 63.895 146.520 ;
        RECT 63.130 146.320 63.450 146.380 ;
        RECT 63.605 146.335 63.895 146.380 ;
        RECT 29.090 146.180 29.410 146.240 ;
        RECT 34.610 146.180 34.930 146.240 ;
        RECT 47.030 146.180 47.350 146.240 ;
        RECT 29.090 146.040 34.930 146.180 ;
        RECT 29.090 145.980 29.410 146.040 ;
        RECT 34.610 145.980 34.930 146.040 ;
        RECT 42.520 146.040 47.350 146.180 ;
        RECT 42.520 145.900 42.660 146.040 ;
        RECT 47.030 145.980 47.350 146.040 ;
        RECT 74.630 146.180 74.950 146.240 ;
        RECT 76.025 146.180 76.315 146.225 ;
        RECT 78.325 146.180 78.615 146.225 ;
        RECT 74.630 146.040 78.615 146.180 ;
        RECT 74.630 145.980 74.950 146.040 ;
        RECT 76.025 145.995 76.315 146.040 ;
        RECT 78.325 145.995 78.615 146.040 ;
        RECT 27.710 145.840 28.030 145.900 ;
        RECT 27.710 145.700 33.920 145.840 ;
        RECT 27.710 145.640 28.030 145.700 ;
        RECT 28.170 145.300 28.490 145.560 ;
        RECT 29.090 145.300 29.410 145.560 ;
        RECT 29.550 145.500 29.870 145.560 ;
        RECT 31.390 145.500 31.710 145.560 ;
        RECT 32.860 145.545 33.000 145.700 ;
        RECT 29.550 145.360 31.710 145.500 ;
        RECT 29.550 145.300 29.870 145.360 ;
        RECT 31.390 145.300 31.710 145.360 ;
        RECT 32.785 145.315 33.075 145.545 ;
        RECT 33.245 145.315 33.535 145.545 ;
        RECT 33.320 145.160 33.460 145.315 ;
        RECT 32.400 145.020 33.460 145.160 ;
        RECT 33.780 145.160 33.920 145.700 ;
        RECT 42.430 145.640 42.750 145.900 ;
        RECT 42.890 145.885 43.210 145.900 ;
        RECT 42.890 145.655 43.320 145.885 ;
        RECT 71.425 145.840 71.715 145.885 ;
        RECT 75.090 145.840 75.410 145.900 ;
        RECT 71.425 145.700 75.410 145.840 ;
        RECT 71.425 145.655 71.715 145.700 ;
        RECT 42.890 145.640 43.210 145.655 ;
        RECT 36.465 145.500 36.755 145.545 ;
        RECT 39.225 145.500 39.515 145.545 ;
        RECT 36.465 145.360 39.515 145.500 ;
        RECT 36.465 145.315 36.755 145.360 ;
        RECT 39.225 145.315 39.515 145.360 ;
        RECT 40.605 145.500 40.895 145.545 ;
        RECT 48.870 145.500 49.190 145.560 ;
        RECT 40.605 145.360 49.190 145.500 ;
        RECT 40.605 145.315 40.895 145.360 ;
        RECT 48.870 145.300 49.190 145.360 ;
        RECT 59.005 145.315 59.295 145.545 ;
        RECT 59.465 145.500 59.755 145.545 ;
        RECT 60.370 145.500 60.690 145.560 ;
        RECT 59.465 145.360 60.690 145.500 ;
        RECT 59.465 145.315 59.755 145.360 ;
        RECT 36.925 145.160 37.215 145.205 ;
        RECT 33.780 145.020 37.215 145.160 ;
        RECT 26.330 144.820 26.650 144.880 ;
        RECT 28.645 144.820 28.935 144.865 ;
        RECT 26.330 144.680 28.935 144.820 ;
        RECT 26.330 144.620 26.650 144.680 ;
        RECT 28.645 144.635 28.935 144.680 ;
        RECT 31.850 144.820 32.170 144.880 ;
        RECT 32.400 144.865 32.540 145.020 ;
        RECT 36.925 144.975 37.215 145.020 ;
        RECT 37.845 144.975 38.135 145.205 ;
        RECT 41.985 145.160 42.275 145.205 ;
        RECT 47.490 145.160 47.810 145.220 ;
        RECT 49.790 145.160 50.110 145.220 ;
        RECT 41.985 145.020 50.110 145.160 ;
        RECT 59.080 145.160 59.220 145.315 ;
        RECT 60.370 145.300 60.690 145.360 ;
        RECT 60.830 145.300 61.150 145.560 ;
        RECT 62.685 145.500 62.975 145.545 ;
        RECT 65.430 145.500 65.750 145.560 ;
        RECT 62.685 145.360 65.750 145.500 ;
        RECT 62.685 145.315 62.975 145.360 ;
        RECT 65.430 145.300 65.750 145.360 ;
        RECT 66.825 145.500 67.115 145.545 ;
        RECT 71.500 145.500 71.640 145.655 ;
        RECT 75.090 145.640 75.410 145.700 ;
        RECT 66.825 145.360 70.030 145.500 ;
        RECT 66.825 145.315 67.115 145.360 ;
        RECT 69.890 145.220 70.030 145.360 ;
        RECT 61.290 145.160 61.610 145.220 ;
        RECT 59.080 145.020 61.610 145.160 ;
        RECT 41.985 144.975 42.275 145.020 ;
        RECT 32.325 144.820 32.615 144.865 ;
        RECT 37.920 144.820 38.060 144.975 ;
        RECT 47.490 144.960 47.810 145.020 ;
        RECT 49.790 144.960 50.110 145.020 ;
        RECT 61.290 144.960 61.610 145.020 ;
        RECT 64.970 145.160 65.290 145.220 ;
        RECT 67.270 145.160 67.590 145.220 ;
        RECT 64.970 145.020 67.590 145.160 ;
        RECT 64.970 144.960 65.290 145.020 ;
        RECT 67.270 144.960 67.590 145.020 ;
        RECT 69.570 145.160 70.030 145.220 ;
        RECT 70.580 145.360 71.640 145.500 ;
        RECT 70.580 145.160 70.720 145.360 ;
        RECT 73.710 145.300 74.030 145.560 ;
        RECT 76.930 145.500 77.250 145.560 ;
        RECT 79.245 145.500 79.535 145.545 ;
        RECT 76.930 145.360 79.535 145.500 ;
        RECT 76.930 145.300 77.250 145.360 ;
        RECT 79.245 145.315 79.535 145.360 ;
        RECT 69.570 145.020 70.720 145.160 ;
        RECT 70.950 145.160 71.270 145.220 ;
        RECT 73.265 145.160 73.555 145.205 ;
        RECT 75.550 145.160 75.870 145.220 ;
        RECT 70.950 145.020 75.870 145.160 ;
        RECT 69.570 144.960 69.890 145.020 ;
        RECT 70.950 144.960 71.270 145.020 ;
        RECT 73.265 144.975 73.555 145.020 ;
        RECT 75.550 144.960 75.870 145.020 ;
        RECT 76.025 145.160 76.315 145.205 ;
        RECT 76.470 145.160 76.790 145.220 ;
        RECT 76.025 145.020 76.790 145.160 ;
        RECT 76.025 144.975 76.315 145.020 ;
        RECT 76.470 144.960 76.790 145.020 ;
        RECT 31.850 144.680 38.060 144.820 ;
        RECT 39.210 144.820 39.530 144.880 ;
        RECT 39.685 144.820 39.975 144.865 ;
        RECT 39.210 144.680 39.975 144.820 ;
        RECT 31.850 144.620 32.170 144.680 ;
        RECT 32.325 144.635 32.615 144.680 ;
        RECT 39.210 144.620 39.530 144.680 ;
        RECT 39.685 144.635 39.975 144.680 ;
        RECT 72.330 144.620 72.650 144.880 ;
        RECT 100.010 144.620 100.880 146.720 ;
        RECT 106.550 146.330 107.800 146.770 ;
        RECT 117.700 146.750 118.560 148.920 ;
        RECT 120.000 146.750 120.770 150.410 ;
        RECT 122.340 149.360 125.190 150.480 ;
        RECT 125.580 150.180 125.930 150.930 ;
        RECT 126.680 150.810 128.550 150.970 ;
        RECT 126.680 150.760 127.440 150.810 ;
        RECT 128.320 150.740 128.550 150.810 ;
        RECT 136.960 150.740 137.190 150.970 ;
        RECT 128.755 150.460 136.755 150.690 ;
        RECT 125.580 150.120 125.870 150.180 ;
        RECT 125.490 150.000 125.870 150.120 ;
        RECT 128.850 150.060 136.710 150.460 ;
        RECT 137.520 150.060 138.480 159.540 ;
        RECT 122.280 149.130 125.280 149.360 ;
        RECT 125.490 149.170 125.830 150.000 ;
        RECT 127.840 149.990 138.480 150.060 ;
        RECT 122.330 149.100 125.190 149.130 ;
        RECT 122.330 149.080 123.500 149.100 ;
        RECT 124.460 149.090 125.190 149.100 ;
        RECT 122.280 148.690 125.280 148.920 ;
        RECT 125.485 148.880 125.830 149.170 ;
        RECT 126.020 148.950 138.480 149.990 ;
        RECT 139.930 161.720 140.700 165.410 ;
        RECT 142.370 164.360 145.220 165.480 ;
        RECT 145.610 165.180 145.960 165.930 ;
        RECT 146.710 165.810 148.580 165.970 ;
        RECT 146.710 165.760 147.470 165.810 ;
        RECT 148.350 165.740 148.580 165.810 ;
        RECT 156.990 165.740 157.220 165.970 ;
        RECT 148.785 165.460 156.785 165.690 ;
        RECT 145.610 165.120 145.900 165.180 ;
        RECT 145.520 165.000 145.900 165.120 ;
        RECT 148.880 165.060 156.740 165.460 ;
        RECT 157.550 165.060 158.510 174.540 ;
        RECT 142.310 164.130 145.310 164.360 ;
        RECT 145.520 164.170 145.860 165.000 ;
        RECT 147.870 164.990 158.510 165.060 ;
        RECT 142.360 164.100 145.220 164.130 ;
        RECT 142.360 164.080 143.530 164.100 ;
        RECT 144.490 164.090 145.220 164.100 ;
        RECT 142.310 163.690 145.310 163.920 ;
        RECT 145.515 163.880 145.860 164.170 ;
        RECT 146.050 163.950 158.510 164.990 ;
        RECT 146.050 163.930 158.500 163.950 ;
        RECT 145.520 163.770 145.860 163.880 ;
        RECT 146.090 163.920 151.760 163.930 ;
        RECT 152.760 163.920 158.500 163.930 ;
        RECT 142.400 163.520 145.260 163.690 ;
        RECT 146.090 163.520 146.520 163.920 ;
        RECT 142.370 163.150 146.520 163.520 ;
        RECT 139.930 159.620 140.840 161.720 ;
        RECT 146.510 161.330 147.760 161.770 ;
        RECT 157.640 161.750 158.500 163.920 ;
        RECT 144.450 161.320 149.690 161.330 ;
        RECT 141.500 161.220 156.800 161.320 ;
        RECT 141.500 161.210 156.835 161.220 ;
        RECT 141.460 161.090 156.835 161.210 ;
        RECT 141.460 160.980 145.460 161.090 ;
        RECT 146.510 161.010 148.250 161.090 ;
        RECT 148.830 161.010 156.835 161.090 ;
        RECT 146.510 160.930 147.760 161.010 ;
        RECT 148.835 160.990 156.835 161.010 ;
        RECT 141.070 160.680 141.300 160.930 ;
        RECT 145.620 160.790 145.850 160.930 ;
        RECT 148.400 160.790 148.630 160.940 ;
        RECT 145.620 160.680 148.630 160.790 ;
        RECT 157.040 160.680 157.270 160.940 ;
        RECT 141.070 160.240 157.270 160.680 ;
        RECT 141.070 159.970 141.300 160.240 ;
        RECT 145.620 160.210 157.270 160.240 ;
        RECT 145.620 160.120 148.630 160.210 ;
        RECT 145.620 159.970 145.850 160.120 ;
        RECT 148.400 159.980 148.630 160.120 ;
        RECT 157.040 159.980 157.270 160.210 ;
        RECT 141.460 159.690 145.460 159.920 ;
        RECT 148.835 159.710 156.835 159.930 ;
        RECT 157.600 159.710 158.560 161.750 ;
        RECT 148.835 159.700 158.560 159.710 ;
        RECT 141.460 159.620 145.450 159.690 ;
        RECT 139.930 159.510 145.450 159.620 ;
        RECT 148.890 159.540 158.560 159.700 ;
        RECT 139.930 159.420 143.140 159.510 ;
        RECT 156.630 159.490 158.560 159.540 ;
        RECT 139.930 156.150 140.840 159.420 ;
        RECT 144.490 158.960 149.740 158.970 ;
        RECT 144.490 158.850 156.800 158.960 ;
        RECT 141.520 158.790 156.800 158.850 ;
        RECT 141.520 158.780 156.835 158.790 ;
        RECT 141.460 158.650 156.835 158.780 ;
        RECT 141.460 158.640 146.620 158.650 ;
        RECT 141.460 158.550 145.460 158.640 ;
        RECT 148.835 158.560 156.835 158.650 ;
        RECT 148.920 158.550 156.810 158.560 ;
        RECT 141.070 158.190 141.300 158.500 ;
        RECT 141.520 158.190 145.420 158.550 ;
        RECT 145.620 158.190 145.850 158.500 ;
        RECT 141.070 156.850 145.850 158.190 ;
        RECT 141.070 156.540 141.300 156.850 ;
        RECT 145.620 156.540 145.850 156.850 ;
        RECT 148.400 157.970 148.630 158.510 ;
        RECT 149.440 157.970 150.450 158.000 ;
        RECT 157.040 157.970 157.270 158.510 ;
        RECT 148.400 157.070 157.270 157.970 ;
        RECT 148.400 156.550 148.630 157.070 ;
        RECT 149.440 157.000 150.450 157.070 ;
        RECT 157.040 156.550 157.270 157.070 ;
        RECT 141.460 156.260 145.460 156.490 ;
        RECT 148.835 156.270 156.835 156.500 ;
        RECT 139.930 156.110 141.140 156.150 ;
        RECT 139.930 156.030 141.380 156.110 ;
        RECT 141.750 156.040 145.410 156.260 ;
        RECT 141.750 156.030 143.190 156.040 ;
        RECT 139.930 155.990 143.190 156.030 ;
        RECT 139.930 155.900 142.700 155.990 ;
        RECT 148.900 155.980 156.790 156.270 ;
        RECT 139.930 155.840 142.030 155.900 ;
        RECT 139.930 155.790 141.780 155.840 ;
        RECT 139.930 152.450 140.840 155.790 ;
        RECT 148.890 155.490 156.810 155.500 ;
        RECT 145.120 155.480 156.810 155.490 ;
        RECT 141.500 155.360 156.810 155.480 ;
        RECT 141.500 155.350 156.835 155.360 ;
        RECT 141.460 155.230 156.835 155.350 ;
        RECT 141.460 155.120 145.460 155.230 ;
        RECT 141.070 154.780 141.300 155.070 ;
        RECT 141.520 154.780 145.410 155.120 ;
        RECT 145.620 154.780 145.850 155.070 ;
        RECT 141.070 153.410 145.850 154.780 ;
        RECT 141.070 153.110 141.300 153.410 ;
        RECT 145.620 153.110 145.850 153.410 ;
        RECT 141.460 152.830 145.460 153.060 ;
        RECT 141.710 152.600 145.280 152.830 ;
        RECT 141.710 152.450 145.400 152.600 ;
        RECT 139.930 152.170 145.400 152.450 ;
        RECT 146.650 152.280 147.270 155.230 ;
        RECT 148.835 155.130 156.835 155.230 ;
        RECT 148.890 155.120 156.810 155.130 ;
        RECT 148.400 154.420 148.630 155.080 ;
        RECT 149.410 154.420 150.410 154.510 ;
        RECT 157.040 154.420 157.270 155.080 ;
        RECT 148.400 153.600 157.270 154.420 ;
        RECT 148.400 153.120 148.630 153.600 ;
        RECT 149.410 153.510 150.410 153.600 ;
        RECT 157.040 153.120 157.270 153.600 ;
        RECT 148.835 152.840 156.835 153.070 ;
        RECT 139.930 151.710 145.410 152.170 ;
        RECT 139.930 150.360 142.010 151.710 ;
        RECT 143.760 151.700 145.410 151.710 ;
        RECT 142.450 150.430 143.450 151.150 ;
        RECT 143.760 150.890 144.070 151.700 ;
        RECT 144.530 151.420 145.410 151.700 ;
        RECT 145.650 151.880 147.270 152.280 ;
        RECT 148.920 151.930 156.790 152.840 ;
        RECT 144.470 151.190 145.470 151.420 ;
        RECT 145.650 151.230 146.000 151.880 ;
        RECT 146.650 151.870 147.270 151.880 ;
        RECT 148.835 151.700 156.835 151.930 ;
        RECT 148.920 151.690 156.790 151.700 ;
        RECT 144.530 150.980 145.410 151.000 ;
        RECT 143.800 150.600 144.070 150.890 ;
        RECT 144.470 150.750 145.470 150.980 ;
        RECT 145.630 150.940 146.000 151.230 ;
        RECT 145.660 150.880 146.000 150.940 ;
        RECT 146.760 151.550 147.520 151.600 ;
        RECT 148.400 151.550 148.630 151.650 ;
        RECT 146.760 151.340 148.630 151.550 ;
        RECT 157.040 151.340 157.270 151.650 ;
        RECT 146.760 150.920 149.300 151.340 ;
        RECT 156.670 150.920 157.270 151.340 ;
        RECT 144.530 150.600 145.410 150.750 ;
        RECT 144.540 150.430 145.270 150.600 ;
        RECT 126.020 148.930 138.460 148.950 ;
        RECT 125.490 148.770 125.830 148.880 ;
        RECT 126.060 148.920 131.730 148.930 ;
        RECT 132.730 148.920 138.460 148.930 ;
        RECT 122.370 148.520 125.230 148.690 ;
        RECT 126.060 148.520 126.490 148.920 ;
        RECT 122.340 148.150 126.490 148.520 ;
        RECT 104.490 146.320 109.730 146.330 ;
        RECT 101.540 146.220 116.840 146.320 ;
        RECT 101.540 146.210 116.875 146.220 ;
        RECT 101.500 146.090 116.875 146.210 ;
        RECT 101.500 145.980 105.500 146.090 ;
        RECT 106.550 146.010 108.290 146.090 ;
        RECT 108.870 146.010 116.875 146.090 ;
        RECT 106.550 145.930 107.800 146.010 ;
        RECT 108.875 145.990 116.875 146.010 ;
        RECT 101.110 145.680 101.340 145.930 ;
        RECT 105.660 145.790 105.890 145.930 ;
        RECT 108.440 145.790 108.670 145.940 ;
        RECT 105.660 145.680 108.670 145.790 ;
        RECT 117.080 145.680 117.310 145.940 ;
        RECT 101.110 145.240 117.310 145.680 ;
        RECT 101.110 144.970 101.340 145.240 ;
        RECT 105.660 145.210 117.310 145.240 ;
        RECT 105.660 145.120 108.670 145.210 ;
        RECT 105.660 144.970 105.890 145.120 ;
        RECT 108.440 144.980 108.670 145.120 ;
        RECT 117.080 144.980 117.310 145.210 ;
        RECT 101.500 144.690 105.500 144.920 ;
        RECT 108.875 144.710 116.875 144.930 ;
        RECT 117.640 144.710 118.600 146.750 ;
        RECT 108.875 144.700 118.600 144.710 ;
        RECT 101.500 144.620 105.490 144.690 ;
        RECT 100.010 144.510 105.490 144.620 ;
        RECT 108.930 144.540 118.600 144.700 ;
        RECT 13.380 144.000 92.040 144.480 ;
        RECT 100.010 144.420 103.180 144.510 ;
        RECT 116.670 144.490 118.600 144.540 ;
        RECT 23.125 143.800 23.415 143.845 ;
        RECT 25.870 143.800 26.190 143.860 ;
        RECT 28.170 143.800 28.490 143.860 ;
        RECT 23.125 143.660 28.490 143.800 ;
        RECT 23.125 143.615 23.415 143.660 ;
        RECT 25.870 143.600 26.190 143.660 ;
        RECT 28.170 143.600 28.490 143.660 ;
        RECT 51.170 143.800 51.490 143.860 ;
        RECT 51.645 143.800 51.935 143.845 ;
        RECT 51.170 143.660 51.935 143.800 ;
        RECT 51.170 143.600 51.490 143.660 ;
        RECT 51.645 143.615 51.935 143.660 ;
        RECT 59.925 143.800 60.215 143.845 ;
        RECT 60.830 143.800 61.150 143.860 ;
        RECT 59.925 143.660 61.150 143.800 ;
        RECT 59.925 143.615 60.215 143.660 ;
        RECT 60.830 143.600 61.150 143.660 ;
        RECT 65.430 143.600 65.750 143.860 ;
        RECT 76.470 143.800 76.790 143.860 ;
        RECT 76.945 143.800 77.235 143.845 ;
        RECT 76.470 143.660 77.235 143.800 ;
        RECT 76.470 143.600 76.790 143.660 ;
        RECT 76.945 143.615 77.235 143.660 ;
        RECT 29.090 143.460 29.410 143.520 ;
        RECT 27.800 143.320 29.410 143.460 ;
        RECT 24.030 143.120 24.350 143.180 ;
        RECT 25.425 143.120 25.715 143.165 ;
        RECT 24.030 142.980 25.715 143.120 ;
        RECT 24.030 142.920 24.350 142.980 ;
        RECT 25.425 142.935 25.715 142.980 ;
        RECT 26.345 143.120 26.635 143.165 ;
        RECT 27.250 143.120 27.570 143.180 ;
        RECT 27.800 143.165 27.940 143.320 ;
        RECT 29.090 143.260 29.410 143.320 ;
        RECT 31.405 143.460 31.695 143.505 ;
        RECT 34.150 143.460 34.470 143.520 ;
        RECT 39.210 143.460 39.530 143.520 ;
        RECT 46.570 143.460 46.890 143.520 ;
        RECT 50.250 143.460 50.570 143.520 ;
        RECT 31.405 143.320 34.470 143.460 ;
        RECT 31.405 143.275 31.695 143.320 ;
        RECT 34.150 143.260 34.470 143.320 ;
        RECT 38.380 143.320 39.530 143.460 ;
        RECT 26.345 142.980 27.570 143.120 ;
        RECT 26.345 142.935 26.635 142.980 ;
        RECT 24.965 142.780 25.255 142.825 ;
        RECT 26.420 142.780 26.560 142.935 ;
        RECT 27.250 142.920 27.570 142.980 ;
        RECT 27.725 142.935 28.015 143.165 ;
        RECT 24.965 142.640 26.560 142.780 ;
        RECT 26.790 142.780 27.110 142.840 ;
        RECT 27.800 142.780 27.940 142.935 ;
        RECT 29.550 142.920 29.870 143.180 ;
        RECT 38.380 143.165 38.520 143.320 ;
        RECT 39.210 143.260 39.530 143.320 ;
        RECT 39.760 143.320 46.890 143.460 ;
        RECT 39.760 143.180 39.900 143.320 ;
        RECT 46.570 143.260 46.890 143.320 ;
        RECT 48.500 143.320 50.570 143.460 ;
        RECT 30.025 143.120 30.315 143.165 ;
        RECT 38.305 143.120 38.595 143.165 ;
        RECT 30.025 142.980 38.595 143.120 ;
        RECT 30.025 142.935 30.315 142.980 ;
        RECT 38.305 142.935 38.595 142.980 ;
        RECT 38.765 142.935 39.055 143.165 ;
        RECT 26.790 142.640 27.940 142.780 ;
        RECT 30.930 142.780 31.250 142.840 ;
        RECT 35.085 142.780 35.375 142.825 ;
        RECT 30.930 142.640 35.375 142.780 ;
        RECT 24.965 142.595 25.255 142.640 ;
        RECT 26.790 142.580 27.110 142.640 ;
        RECT 30.930 142.580 31.250 142.640 ;
        RECT 35.085 142.595 35.375 142.640 ;
        RECT 36.450 142.580 36.770 142.840 ;
        RECT 26.330 142.440 26.650 142.500 ;
        RECT 38.840 142.440 38.980 142.935 ;
        RECT 39.670 142.920 39.990 143.180 ;
        RECT 41.510 143.120 41.830 143.180 ;
        RECT 43.365 143.120 43.655 143.165 ;
        RECT 41.510 142.980 43.655 143.120 ;
        RECT 41.510 142.920 41.830 142.980 ;
        RECT 43.365 142.935 43.655 142.980 ;
        RECT 44.730 143.120 45.050 143.180 ;
        RECT 48.500 143.165 48.640 143.320 ;
        RECT 50.250 143.260 50.570 143.320 ;
        RECT 50.725 143.460 51.015 143.505 ;
        RECT 59.450 143.460 59.770 143.520 ;
        RECT 71.380 143.460 71.670 143.505 ;
        RECT 72.330 143.460 72.650 143.520 ;
        RECT 50.725 143.320 59.220 143.460 ;
        RECT 50.725 143.275 51.015 143.320 ;
        RECT 44.730 142.980 45.420 143.120 ;
        RECT 44.730 142.920 45.050 142.980 ;
        RECT 26.330 142.300 38.980 142.440 ;
        RECT 45.280 142.440 45.420 142.980 ;
        RECT 45.665 142.935 45.955 143.165 ;
        RECT 48.425 142.935 48.715 143.165 ;
        RECT 45.740 142.780 45.880 142.935 ;
        RECT 49.330 142.920 49.650 143.180 ;
        RECT 57.150 143.165 57.470 143.180 ;
        RECT 57.150 142.935 57.500 143.165 ;
        RECT 59.080 143.120 59.220 143.320 ;
        RECT 59.450 143.320 67.040 143.460 ;
        RECT 59.450 143.260 59.770 143.320 ;
        RECT 59.910 143.120 60.230 143.180 ;
        RECT 59.080 142.980 60.230 143.120 ;
        RECT 57.150 142.920 57.470 142.935 ;
        RECT 59.910 142.920 60.230 142.980 ;
        RECT 60.370 143.120 60.690 143.180 ;
        RECT 60.845 143.120 61.135 143.165 ;
        RECT 60.370 142.980 61.135 143.120 ;
        RECT 60.370 142.920 60.690 142.980 ;
        RECT 60.845 142.935 61.135 142.980 ;
        RECT 61.290 142.920 61.610 143.180 ;
        RECT 62.760 143.165 62.900 143.320 ;
        RECT 62.685 142.935 62.975 143.165 ;
        RECT 66.350 142.920 66.670 143.180 ;
        RECT 48.885 142.780 49.175 142.825 ;
        RECT 45.740 142.640 49.175 142.780 ;
        RECT 48.885 142.595 49.175 142.640 ;
        RECT 53.955 142.780 54.245 142.825 ;
        RECT 56.475 142.780 56.765 142.825 ;
        RECT 57.665 142.780 57.955 142.825 ;
        RECT 53.955 142.640 57.955 142.780 ;
        RECT 53.955 142.595 54.245 142.640 ;
        RECT 56.475 142.595 56.765 142.640 ;
        RECT 57.665 142.595 57.955 142.640 ;
        RECT 58.530 142.580 58.850 142.840 ;
        RECT 62.225 142.780 62.515 142.825 ;
        RECT 66.440 142.780 66.580 142.920 ;
        RECT 62.225 142.640 66.580 142.780 ;
        RECT 66.900 142.780 67.040 143.320 ;
        RECT 71.380 143.320 72.650 143.460 ;
        RECT 71.380 143.275 71.670 143.320 ;
        RECT 72.330 143.260 72.650 143.320 ;
        RECT 67.285 143.120 67.575 143.165 ;
        RECT 68.190 143.120 68.510 143.180 ;
        RECT 67.285 142.980 68.510 143.120 ;
        RECT 67.285 142.935 67.575 142.980 ;
        RECT 68.190 142.920 68.510 142.980 ;
        RECT 67.745 142.780 68.035 142.825 ;
        RECT 66.900 142.640 68.035 142.780 ;
        RECT 62.225 142.595 62.515 142.640 ;
        RECT 67.745 142.595 68.035 142.640 ;
        RECT 69.570 142.780 69.890 142.840 ;
        RECT 70.045 142.780 70.335 142.825 ;
        RECT 69.570 142.640 70.335 142.780 ;
        RECT 69.570 142.580 69.890 142.640 ;
        RECT 70.045 142.595 70.335 142.640 ;
        RECT 70.925 142.780 71.215 142.825 ;
        RECT 72.115 142.780 72.405 142.825 ;
        RECT 74.635 142.780 74.925 142.825 ;
        RECT 70.925 142.640 74.925 142.780 ;
        RECT 70.925 142.595 71.215 142.640 ;
        RECT 72.115 142.595 72.405 142.640 ;
        RECT 74.635 142.595 74.925 142.640 ;
        RECT 49.790 142.440 50.110 142.500 ;
        RECT 45.280 142.300 50.110 142.440 ;
        RECT 26.330 142.240 26.650 142.300 ;
        RECT 49.790 142.240 50.110 142.300 ;
        RECT 54.390 142.440 54.680 142.485 ;
        RECT 55.960 142.440 56.250 142.485 ;
        RECT 58.060 142.440 58.350 142.485 ;
        RECT 54.390 142.300 58.350 142.440 ;
        RECT 54.390 142.255 54.680 142.300 ;
        RECT 55.960 142.255 56.250 142.300 ;
        RECT 58.060 142.255 58.350 142.300 ;
        RECT 70.530 142.440 70.820 142.485 ;
        RECT 72.630 142.440 72.920 142.485 ;
        RECT 74.200 142.440 74.490 142.485 ;
        RECT 70.530 142.300 74.490 142.440 ;
        RECT 70.530 142.255 70.820 142.300 ;
        RECT 72.630 142.255 72.920 142.300 ;
        RECT 74.200 142.255 74.490 142.300 ;
        RECT 27.250 141.900 27.570 142.160 ;
        RECT 27.710 142.100 28.030 142.160 ;
        RECT 28.185 142.100 28.475 142.145 ;
        RECT 27.710 141.960 28.475 142.100 ;
        RECT 27.710 141.900 28.030 141.960 ;
        RECT 28.185 141.915 28.475 141.960 ;
        RECT 30.945 142.100 31.235 142.145 ;
        RECT 31.390 142.100 31.710 142.160 ;
        RECT 30.945 141.960 31.710 142.100 ;
        RECT 30.945 141.915 31.235 141.960 ;
        RECT 31.390 141.900 31.710 141.960 ;
        RECT 37.385 142.100 37.675 142.145 ;
        RECT 39.210 142.100 39.530 142.160 ;
        RECT 37.385 141.960 39.530 142.100 ;
        RECT 37.385 141.915 37.675 141.960 ;
        RECT 39.210 141.900 39.530 141.960 ;
        RECT 42.430 141.900 42.750 142.160 ;
        RECT 45.650 141.900 45.970 142.160 ;
        RECT 47.490 142.100 47.810 142.160 ;
        RECT 50.265 142.100 50.555 142.145 ;
        RECT 53.470 142.100 53.790 142.160 ;
        RECT 47.490 141.960 53.790 142.100 ;
        RECT 47.490 141.900 47.810 141.960 ;
        RECT 50.265 141.915 50.555 141.960 ;
        RECT 53.470 141.900 53.790 141.960 ;
        RECT 13.380 141.280 92.040 141.760 ;
        RECT 100.010 141.150 100.880 144.420 ;
        RECT 104.530 143.960 109.780 143.970 ;
        RECT 104.530 143.850 116.840 143.960 ;
        RECT 101.560 143.790 116.840 143.850 ;
        RECT 101.560 143.780 116.875 143.790 ;
        RECT 101.500 143.650 116.875 143.780 ;
        RECT 101.500 143.640 106.660 143.650 ;
        RECT 101.500 143.550 105.500 143.640 ;
        RECT 108.875 143.560 116.875 143.650 ;
        RECT 108.960 143.550 116.850 143.560 ;
        RECT 101.110 143.190 101.340 143.500 ;
        RECT 101.560 143.190 105.460 143.550 ;
        RECT 105.660 143.190 105.890 143.500 ;
        RECT 101.110 141.850 105.890 143.190 ;
        RECT 101.110 141.540 101.340 141.850 ;
        RECT 105.660 141.540 105.890 141.850 ;
        RECT 108.440 142.970 108.670 143.510 ;
        RECT 109.480 142.970 110.490 143.000 ;
        RECT 117.080 142.970 117.310 143.510 ;
        RECT 108.440 142.070 117.310 142.970 ;
        RECT 108.440 141.550 108.670 142.070 ;
        RECT 109.480 142.000 110.490 142.070 ;
        RECT 117.080 141.550 117.310 142.070 ;
        RECT 101.500 141.260 105.500 141.490 ;
        RECT 108.875 141.270 116.875 141.500 ;
        RECT 25.885 141.080 26.175 141.125 ;
        RECT 27.710 141.080 28.030 141.140 ;
        RECT 36.450 141.080 36.770 141.140 ;
        RECT 25.885 140.940 28.030 141.080 ;
        RECT 25.885 140.895 26.175 140.940 ;
        RECT 27.710 140.880 28.030 140.940 ;
        RECT 28.260 140.940 36.770 141.080 ;
        RECT 28.260 140.800 28.400 140.940 ;
        RECT 36.450 140.880 36.770 140.940 ;
        RECT 48.885 141.080 49.175 141.125 ;
        RECT 50.250 141.080 50.570 141.140 ;
        RECT 48.885 140.940 50.570 141.080 ;
        RECT 48.885 140.895 49.175 140.940 ;
        RECT 50.250 140.880 50.570 140.940 ;
        RECT 50.725 141.080 51.015 141.125 ;
        RECT 55.310 141.080 55.630 141.140 ;
        RECT 57.150 141.080 57.470 141.140 ;
        RECT 50.725 140.940 55.630 141.080 ;
        RECT 50.725 140.895 51.015 140.940 ;
        RECT 55.310 140.880 55.630 140.940 ;
        RECT 55.860 140.940 57.470 141.080 ;
        RECT 19.470 140.740 19.760 140.785 ;
        RECT 21.570 140.740 21.860 140.785 ;
        RECT 23.140 140.740 23.430 140.785 ;
        RECT 19.470 140.600 23.430 140.740 ;
        RECT 19.470 140.555 19.760 140.600 ;
        RECT 21.570 140.555 21.860 140.600 ;
        RECT 23.140 140.555 23.430 140.600 ;
        RECT 28.170 140.540 28.490 140.800 ;
        RECT 31.850 140.740 32.140 140.785 ;
        RECT 33.420 140.740 33.710 140.785 ;
        RECT 35.520 140.740 35.810 140.785 ;
        RECT 31.850 140.600 35.810 140.740 ;
        RECT 31.850 140.555 32.140 140.600 ;
        RECT 33.420 140.555 33.710 140.600 ;
        RECT 35.520 140.555 35.810 140.600 ;
        RECT 42.470 140.740 42.760 140.785 ;
        RECT 44.570 140.740 44.860 140.785 ;
        RECT 46.140 140.740 46.430 140.785 ;
        RECT 42.470 140.600 46.430 140.740 ;
        RECT 42.470 140.555 42.760 140.600 ;
        RECT 44.570 140.555 44.860 140.600 ;
        RECT 46.140 140.555 46.430 140.600 ;
        RECT 49.330 140.740 49.650 140.800 ;
        RECT 51.645 140.740 51.935 140.785 ;
        RECT 52.550 140.740 52.870 140.800 ;
        RECT 55.860 140.785 56.000 140.940 ;
        RECT 57.150 140.880 57.470 140.940 ;
        RECT 100.010 141.110 101.180 141.150 ;
        RECT 100.010 141.030 101.420 141.110 ;
        RECT 101.790 141.040 105.450 141.260 ;
        RECT 101.790 141.030 103.230 141.040 ;
        RECT 100.010 140.990 103.230 141.030 ;
        RECT 100.010 140.900 102.740 140.990 ;
        RECT 108.940 140.980 116.830 141.270 ;
        RECT 100.010 140.840 102.070 140.900 ;
        RECT 49.330 140.600 52.870 140.740 ;
        RECT 49.330 140.540 49.650 140.600 ;
        RECT 51.645 140.555 51.935 140.600 ;
        RECT 52.550 140.540 52.870 140.600 ;
        RECT 53.100 140.600 55.540 140.740 ;
        RECT 18.970 140.200 19.290 140.460 ;
        RECT 19.865 140.400 20.155 140.445 ;
        RECT 21.055 140.400 21.345 140.445 ;
        RECT 23.575 140.400 23.865 140.445 ;
        RECT 19.865 140.260 23.865 140.400 ;
        RECT 19.865 140.215 20.155 140.260 ;
        RECT 21.055 140.215 21.345 140.260 ;
        RECT 23.575 140.215 23.865 140.260 ;
        RECT 31.415 140.400 31.705 140.445 ;
        RECT 33.935 140.400 34.225 140.445 ;
        RECT 35.125 140.400 35.415 140.445 ;
        RECT 39.670 140.400 39.990 140.460 ;
        RECT 41.985 140.400 42.275 140.445 ;
        RECT 31.415 140.260 35.415 140.400 ;
        RECT 31.415 140.215 31.705 140.260 ;
        RECT 33.935 140.215 34.225 140.260 ;
        RECT 35.125 140.215 35.415 140.260 ;
        RECT 37.000 140.260 42.275 140.400 ;
        RECT 19.060 140.060 19.200 140.200 ;
        RECT 37.000 140.120 37.140 140.260 ;
        RECT 39.670 140.200 39.990 140.260 ;
        RECT 41.985 140.215 42.275 140.260 ;
        RECT 42.865 140.400 43.155 140.445 ;
        RECT 44.055 140.400 44.345 140.445 ;
        RECT 46.575 140.400 46.865 140.445 ;
        RECT 51.170 140.400 51.490 140.460 ;
        RECT 53.100 140.400 53.240 140.600 ;
        RECT 42.865 140.260 46.865 140.400 ;
        RECT 42.865 140.215 43.155 140.260 ;
        RECT 44.055 140.215 44.345 140.260 ;
        RECT 46.575 140.215 46.865 140.260 ;
        RECT 49.880 140.260 51.490 140.400 ;
        RECT 23.110 140.060 23.430 140.120 ;
        RECT 30.930 140.060 31.250 140.120 ;
        RECT 19.060 139.920 31.250 140.060 ;
        RECT 23.110 139.860 23.430 139.920 ;
        RECT 30.930 139.860 31.250 139.920 ;
        RECT 36.005 140.060 36.295 140.105 ;
        RECT 36.910 140.060 37.230 140.120 ;
        RECT 36.005 139.920 37.230 140.060 ;
        RECT 36.005 139.875 36.295 139.920 ;
        RECT 36.910 139.860 37.230 139.920 ;
        RECT 39.210 139.860 39.530 140.120 ;
        RECT 20.320 139.720 20.610 139.765 ;
        RECT 21.270 139.720 21.590 139.780 ;
        RECT 20.320 139.580 21.590 139.720 ;
        RECT 20.320 139.535 20.610 139.580 ;
        RECT 21.270 139.520 21.590 139.580 ;
        RECT 25.410 139.720 25.730 139.780 ;
        RECT 27.725 139.720 28.015 139.765 ;
        RECT 25.410 139.580 28.015 139.720 ;
        RECT 25.410 139.520 25.730 139.580 ;
        RECT 27.725 139.535 28.015 139.580 ;
        RECT 34.780 139.720 35.070 139.765 ;
        RECT 36.465 139.720 36.755 139.765 ;
        RECT 34.780 139.580 36.755 139.720 ;
        RECT 34.780 139.535 35.070 139.580 ;
        RECT 36.465 139.535 36.755 139.580 ;
        RECT 43.320 139.720 43.610 139.765 ;
        RECT 45.190 139.720 45.510 139.780 ;
        RECT 49.880 139.765 50.020 140.260 ;
        RECT 51.170 140.200 51.490 140.260 ;
        RECT 52.180 140.260 53.240 140.400 ;
        RECT 55.400 140.400 55.540 140.600 ;
        RECT 55.785 140.555 56.075 140.785 ;
        RECT 56.230 140.540 56.550 140.800 ;
        RECT 100.010 140.790 101.820 140.840 ;
        RECT 55.400 140.260 57.840 140.400 ;
        RECT 50.710 139.765 51.030 139.780 ;
        RECT 43.320 139.580 45.510 139.720 ;
        RECT 43.320 139.535 43.610 139.580 ;
        RECT 45.190 139.520 45.510 139.580 ;
        RECT 49.805 139.535 50.095 139.765 ;
        RECT 50.710 139.720 51.175 139.765 ;
        RECT 52.180 139.720 52.320 140.260 ;
        RECT 52.565 139.875 52.855 140.105 ;
        RECT 53.470 140.060 53.790 140.120 ;
        RECT 53.945 140.060 54.235 140.105 ;
        RECT 54.390 140.060 54.710 140.120 ;
        RECT 57.700 140.105 57.840 140.260 ;
        RECT 58.530 140.200 58.850 140.460 ;
        RECT 61.750 140.400 62.070 140.460 ;
        RECT 64.525 140.400 64.815 140.445 ;
        RECT 59.080 140.260 64.815 140.400 ;
        RECT 53.470 139.920 54.710 140.060 ;
        RECT 50.710 139.580 52.320 139.720 ;
        RECT 50.710 139.535 51.175 139.580 ;
        RECT 50.710 139.520 51.030 139.535 ;
        RECT 22.650 139.380 22.970 139.440 ;
        RECT 28.170 139.380 28.490 139.440 ;
        RECT 22.650 139.240 28.490 139.380 ;
        RECT 22.650 139.180 22.970 139.240 ;
        RECT 28.170 139.180 28.490 139.240 ;
        RECT 29.105 139.380 29.395 139.425 ;
        RECT 31.850 139.380 32.170 139.440 ;
        RECT 29.105 139.240 32.170 139.380 ;
        RECT 29.105 139.195 29.395 139.240 ;
        RECT 31.850 139.180 32.170 139.240 ;
        RECT 48.870 139.380 49.190 139.440 ;
        RECT 52.640 139.380 52.780 139.875 ;
        RECT 53.470 139.860 53.790 139.920 ;
        RECT 53.945 139.875 54.235 139.920 ;
        RECT 54.390 139.860 54.710 139.920 ;
        RECT 57.625 140.060 57.915 140.105 ;
        RECT 59.080 140.060 59.220 140.260 ;
        RECT 61.750 140.200 62.070 140.260 ;
        RECT 64.525 140.215 64.815 140.260 ;
        RECT 57.625 139.920 59.220 140.060 ;
        RECT 63.590 140.060 63.910 140.120 ;
        RECT 66.350 140.060 66.670 140.120 ;
        RECT 67.285 140.060 67.575 140.105 ;
        RECT 63.590 139.920 67.575 140.060 ;
        RECT 57.625 139.875 57.915 139.920 ;
        RECT 63.590 139.860 63.910 139.920 ;
        RECT 66.350 139.860 66.670 139.920 ;
        RECT 67.285 139.875 67.575 139.920 ;
        RECT 53.010 139.720 53.330 139.780 ;
        RECT 54.990 139.720 55.280 139.765 ;
        RECT 53.010 139.580 55.280 139.720 ;
        RECT 53.010 139.520 53.330 139.580 ;
        RECT 54.990 139.535 55.280 139.580 ;
        RECT 55.770 139.720 56.090 139.780 ;
        RECT 56.245 139.720 56.535 139.765 ;
        RECT 55.770 139.580 56.535 139.720 ;
        RECT 55.770 139.520 56.090 139.580 ;
        RECT 56.245 139.535 56.535 139.580 ;
        RECT 58.990 139.720 59.310 139.780 ;
        RECT 62.685 139.720 62.975 139.765 ;
        RECT 64.970 139.720 65.290 139.780 ;
        RECT 58.990 139.580 65.290 139.720 ;
        RECT 58.990 139.520 59.310 139.580 ;
        RECT 62.685 139.535 62.975 139.580 ;
        RECT 64.970 139.520 65.290 139.580 ;
        RECT 65.445 139.720 65.735 139.765 ;
        RECT 66.810 139.720 67.130 139.780 ;
        RECT 69.110 139.720 69.430 139.780 ;
        RECT 65.445 139.580 69.430 139.720 ;
        RECT 65.445 139.535 65.735 139.580 ;
        RECT 66.810 139.520 67.130 139.580 ;
        RECT 69.110 139.520 69.430 139.580 ;
        RECT 48.870 139.240 52.780 139.380 ;
        RECT 48.870 139.180 49.190 139.240 ;
        RECT 54.390 139.180 54.710 139.440 ;
        RECT 56.690 139.380 57.010 139.440 ;
        RECT 57.165 139.380 57.455 139.425 ;
        RECT 60.830 139.380 61.150 139.440 ;
        RECT 56.690 139.240 61.150 139.380 ;
        RECT 56.690 139.180 57.010 139.240 ;
        RECT 57.165 139.195 57.455 139.240 ;
        RECT 60.830 139.180 61.150 139.240 ;
        RECT 65.890 139.180 66.210 139.440 ;
        RECT 66.365 139.380 66.655 139.425 ;
        RECT 68.190 139.380 68.510 139.440 ;
        RECT 66.365 139.240 68.510 139.380 ;
        RECT 66.365 139.195 66.655 139.240 ;
        RECT 68.190 139.180 68.510 139.240 ;
        RECT 13.380 138.560 92.040 139.040 ;
        RECT 21.270 138.160 21.590 138.420 ;
        RECT 22.205 138.360 22.495 138.405 ;
        RECT 22.650 138.360 22.970 138.420 ;
        RECT 22.205 138.220 22.970 138.360 ;
        RECT 22.205 138.175 22.495 138.220 ;
        RECT 22.650 138.160 22.970 138.220 ;
        RECT 27.725 138.360 28.015 138.405 ;
        RECT 29.185 138.360 29.475 138.405 ;
        RECT 27.725 138.220 29.475 138.360 ;
        RECT 27.725 138.175 28.015 138.220 ;
        RECT 29.185 138.175 29.475 138.220 ;
        RECT 30.025 138.175 30.315 138.405 ;
        RECT 45.190 138.360 45.510 138.420 ;
        RECT 45.665 138.360 45.955 138.405 ;
        RECT 45.190 138.220 45.955 138.360 ;
        RECT 25.870 138.020 26.190 138.080 ;
        RECT 24.120 137.880 26.190 138.020 ;
        RECT 24.120 137.725 24.260 137.880 ;
        RECT 25.870 137.820 26.190 137.880 ;
        RECT 28.170 137.820 28.490 138.080 ;
        RECT 30.100 138.020 30.240 138.175 ;
        RECT 45.190 138.160 45.510 138.220 ;
        RECT 45.665 138.175 45.955 138.220 ;
        RECT 47.030 138.160 47.350 138.420 ;
        RECT 47.490 138.160 47.810 138.420 ;
        RECT 49.345 138.360 49.635 138.405 ;
        RECT 49.790 138.360 50.110 138.420 ;
        RECT 49.345 138.220 50.110 138.360 ;
        RECT 49.345 138.175 49.635 138.220 ;
        RECT 49.790 138.160 50.110 138.220 ;
        RECT 50.250 138.360 50.570 138.420 ;
        RECT 51.185 138.360 51.475 138.405 ;
        RECT 50.250 138.220 51.475 138.360 ;
        RECT 50.250 138.160 50.570 138.220 ;
        RECT 51.185 138.175 51.475 138.220 ;
        RECT 53.010 138.160 53.330 138.420 ;
        RECT 59.910 138.360 60.230 138.420 ;
        RECT 70.950 138.360 71.270 138.420 ;
        RECT 71.885 138.360 72.175 138.405 ;
        RECT 59.910 138.220 72.175 138.360 ;
        RECT 59.910 138.160 60.230 138.220 ;
        RECT 70.950 138.160 71.270 138.220 ;
        RECT 71.885 138.175 72.175 138.220 ;
        RECT 73.265 138.175 73.555 138.405 ;
        RECT 31.710 138.020 32.000 138.065 ;
        RECT 30.100 137.880 32.000 138.020 ;
        RECT 31.710 137.835 32.000 137.880 ;
        RECT 35.530 138.020 35.850 138.080 ;
        RECT 40.605 138.020 40.895 138.065 ;
        RECT 58.990 138.020 59.310 138.080 ;
        RECT 35.530 137.880 59.310 138.020 ;
        RECT 35.530 137.820 35.850 137.880 ;
        RECT 40.605 137.835 40.895 137.880 ;
        RECT 58.990 137.820 59.310 137.880 ;
        RECT 61.290 138.020 61.610 138.080 ;
        RECT 70.030 138.020 70.350 138.080 ;
        RECT 71.410 138.020 71.730 138.080 ;
        RECT 61.290 137.880 71.730 138.020 ;
        RECT 73.340 138.020 73.480 138.175 ;
        RECT 79.290 138.020 79.580 138.065 ;
        RECT 73.340 137.880 79.580 138.020 ;
        RECT 61.290 137.820 61.610 137.880 ;
        RECT 70.030 137.820 70.350 137.880 ;
        RECT 71.410 137.820 71.730 137.880 ;
        RECT 79.290 137.835 79.580 137.880 ;
        RECT 16.225 137.680 16.515 137.725 ;
        RECT 16.225 137.540 21.730 137.680 ;
        RECT 16.225 137.495 16.515 137.540 ;
        RECT 21.590 137.340 21.730 137.540 ;
        RECT 24.045 137.495 24.335 137.725 ;
        RECT 26.790 137.680 27.110 137.740 ;
        RECT 30.485 137.680 30.775 137.725 ;
        RECT 30.930 137.680 31.250 137.740 ;
        RECT 26.790 137.540 30.240 137.680 ;
        RECT 26.790 137.480 27.110 137.540 ;
        RECT 28.170 137.340 28.490 137.400 ;
        RECT 21.590 137.200 28.490 137.340 ;
        RECT 28.170 137.140 28.490 137.200 ;
        RECT 26.330 137.000 26.650 137.060 ;
        RECT 26.330 136.860 29.320 137.000 ;
        RECT 26.330 136.800 26.650 136.860 ;
        RECT 12.070 136.660 12.390 136.720 ;
        RECT 15.305 136.660 15.595 136.705 ;
        RECT 12.070 136.520 15.595 136.660 ;
        RECT 12.070 136.460 12.390 136.520 ;
        RECT 15.305 136.475 15.595 136.520 ;
        RECT 22.205 136.660 22.495 136.705 ;
        RECT 27.250 136.660 27.570 136.720 ;
        RECT 29.180 136.705 29.320 136.860 ;
        RECT 22.205 136.520 27.570 136.660 ;
        RECT 22.205 136.475 22.495 136.520 ;
        RECT 27.250 136.460 27.570 136.520 ;
        RECT 29.105 136.475 29.395 136.705 ;
        RECT 30.100 136.660 30.240 137.540 ;
        RECT 30.485 137.540 31.250 137.680 ;
        RECT 30.485 137.495 30.775 137.540 ;
        RECT 30.930 137.480 31.250 137.540 ;
        RECT 45.650 137.680 45.970 137.740 ;
        RECT 46.460 137.680 46.750 137.725 ;
        RECT 45.650 137.540 46.750 137.680 ;
        RECT 45.650 137.480 45.970 137.540 ;
        RECT 46.460 137.495 46.750 137.540 ;
        RECT 50.250 137.480 50.570 137.740 ;
        RECT 50.725 137.495 51.015 137.725 ;
        RECT 51.170 137.680 51.490 137.740 ;
        RECT 52.105 137.680 52.395 137.725 ;
        RECT 51.170 137.540 52.395 137.680 ;
        RECT 31.365 137.340 31.655 137.385 ;
        RECT 32.555 137.340 32.845 137.385 ;
        RECT 35.075 137.340 35.365 137.385 ;
        RECT 31.365 137.200 35.365 137.340 ;
        RECT 31.365 137.155 31.655 137.200 ;
        RECT 32.555 137.155 32.845 137.200 ;
        RECT 35.075 137.155 35.365 137.200 ;
        RECT 36.910 137.340 37.230 137.400 ;
        RECT 44.285 137.340 44.575 137.385 ;
        RECT 36.910 137.200 44.575 137.340 ;
        RECT 36.910 137.140 37.230 137.200 ;
        RECT 44.285 137.155 44.575 137.200 ;
        RECT 48.870 137.140 49.190 137.400 ;
        RECT 50.800 137.340 50.940 137.495 ;
        RECT 51.170 137.480 51.490 137.540 ;
        RECT 52.105 137.495 52.395 137.540 ;
        RECT 52.180 137.340 52.320 137.495 ;
        RECT 52.550 137.480 52.870 137.740 ;
        RECT 53.485 137.680 53.775 137.725 ;
        RECT 56.230 137.680 56.550 137.740 ;
        RECT 53.485 137.540 56.550 137.680 ;
        RECT 53.485 137.495 53.775 137.540 ;
        RECT 56.230 137.480 56.550 137.540 ;
        RECT 58.530 137.480 58.850 137.740 ;
        RECT 65.890 137.680 66.210 137.740 ;
        RECT 67.285 137.680 67.575 137.725 ;
        RECT 65.890 137.540 67.575 137.680 ;
        RECT 65.890 137.480 66.210 137.540 ;
        RECT 67.285 137.495 67.575 137.540 ;
        RECT 68.190 137.480 68.510 137.740 ;
        RECT 76.930 137.680 77.250 137.740 ;
        RECT 68.740 137.540 77.250 137.680 ;
        RECT 55.770 137.340 56.090 137.400 ;
        RECT 68.740 137.340 68.880 137.540 ;
        RECT 76.930 137.480 77.250 137.540 ;
        RECT 77.390 137.680 77.710 137.740 ;
        RECT 80.625 137.680 80.915 137.725 ;
        RECT 77.390 137.540 80.915 137.680 ;
        RECT 77.390 137.480 77.710 137.540 ;
        RECT 80.625 137.495 80.915 137.540 ;
        RECT 100.010 137.450 100.880 140.790 ;
        RECT 108.930 140.490 116.850 140.500 ;
        RECT 105.160 140.480 116.850 140.490 ;
        RECT 101.540 140.360 116.850 140.480 ;
        RECT 101.540 140.350 116.875 140.360 ;
        RECT 101.500 140.230 116.875 140.350 ;
        RECT 101.500 140.120 105.500 140.230 ;
        RECT 101.110 139.780 101.340 140.070 ;
        RECT 101.560 139.780 105.450 140.120 ;
        RECT 105.660 139.780 105.890 140.070 ;
        RECT 101.110 138.410 105.890 139.780 ;
        RECT 101.110 138.110 101.340 138.410 ;
        RECT 105.660 138.110 105.890 138.410 ;
        RECT 101.500 137.830 105.500 138.060 ;
        RECT 101.750 137.600 105.320 137.830 ;
        RECT 101.750 137.450 105.440 137.600 ;
        RECT 50.800 137.200 51.400 137.340 ;
        RECT 52.180 137.200 56.090 137.340 ;
        RECT 30.970 137.000 31.260 137.045 ;
        RECT 33.070 137.000 33.360 137.045 ;
        RECT 34.640 137.000 34.930 137.045 ;
        RECT 30.970 136.860 34.930 137.000 ;
        RECT 30.970 136.815 31.260 136.860 ;
        RECT 33.070 136.815 33.360 136.860 ;
        RECT 34.640 136.815 34.930 136.860 ;
        RECT 37.385 136.660 37.675 136.705 ;
        RECT 30.100 136.520 37.675 136.660 ;
        RECT 37.385 136.475 37.675 136.520 ;
        RECT 49.790 136.660 50.110 136.720 ;
        RECT 51.260 136.660 51.400 137.200 ;
        RECT 55.770 137.140 56.090 137.200 ;
        RECT 56.320 137.200 68.880 137.340 ;
        RECT 53.470 137.000 53.790 137.060 ;
        RECT 56.320 137.000 56.460 137.200 ;
        RECT 70.030 137.140 70.350 137.400 ;
        RECT 71.410 137.140 71.730 137.400 ;
        RECT 72.470 137.340 72.760 137.385 ;
        RECT 73.250 137.340 73.570 137.400 ;
        RECT 72.470 137.200 73.570 137.340 ;
        RECT 72.470 137.155 72.760 137.200 ;
        RECT 73.250 137.140 73.570 137.200 ;
        RECT 76.035 137.340 76.325 137.385 ;
        RECT 78.555 137.340 78.845 137.385 ;
        RECT 79.745 137.340 80.035 137.385 ;
        RECT 76.035 137.200 80.035 137.340 ;
        RECT 76.035 137.155 76.325 137.200 ;
        RECT 78.555 137.155 78.845 137.200 ;
        RECT 79.745 137.155 80.035 137.200 ;
        RECT 100.010 137.170 105.440 137.450 ;
        RECT 106.690 137.280 107.310 140.230 ;
        RECT 108.875 140.130 116.875 140.230 ;
        RECT 108.930 140.120 116.850 140.130 ;
        RECT 108.440 139.420 108.670 140.080 ;
        RECT 109.450 139.420 110.450 139.510 ;
        RECT 117.080 139.420 117.310 140.080 ;
        RECT 108.440 138.600 117.310 139.420 ;
        RECT 108.440 138.120 108.670 138.600 ;
        RECT 109.450 138.510 110.450 138.600 ;
        RECT 117.080 138.120 117.310 138.600 ;
        RECT 108.875 137.840 116.875 138.070 ;
        RECT 53.470 136.860 56.460 137.000 ;
        RECT 66.350 137.000 66.670 137.060 ;
        RECT 73.725 137.000 74.015 137.045 ;
        RECT 66.350 136.860 74.015 137.000 ;
        RECT 53.470 136.800 53.790 136.860 ;
        RECT 66.350 136.800 66.670 136.860 ;
        RECT 73.725 136.815 74.015 136.860 ;
        RECT 76.470 137.000 76.760 137.045 ;
        RECT 78.040 137.000 78.330 137.045 ;
        RECT 80.140 137.000 80.430 137.045 ;
        RECT 76.470 136.860 80.430 137.000 ;
        RECT 76.470 136.815 76.760 136.860 ;
        RECT 78.040 136.815 78.330 136.860 ;
        RECT 80.140 136.815 80.430 136.860 ;
        RECT 56.690 136.660 57.010 136.720 ;
        RECT 49.790 136.520 57.010 136.660 ;
        RECT 49.790 136.460 50.110 136.520 ;
        RECT 56.690 136.460 57.010 136.520 ;
        RECT 68.205 136.660 68.495 136.705 ;
        RECT 68.650 136.660 68.970 136.720 ;
        RECT 68.205 136.520 68.970 136.660 ;
        RECT 68.205 136.475 68.495 136.520 ;
        RECT 68.650 136.460 68.970 136.520 ;
        RECT 100.010 136.710 105.450 137.170 ;
        RECT 13.380 135.840 92.040 136.320 ;
        RECT 42.890 135.640 43.210 135.700 ;
        RECT 47.030 135.640 47.350 135.700 ;
        RECT 54.390 135.640 54.710 135.700 ;
        RECT 42.890 135.500 54.710 135.640 ;
        RECT 42.890 135.440 43.210 135.500 ;
        RECT 47.030 135.440 47.350 135.500 ;
        RECT 54.390 135.440 54.710 135.500 ;
        RECT 65.890 135.440 66.210 135.700 ;
        RECT 66.350 135.640 66.670 135.700 ;
        RECT 66.825 135.640 67.115 135.685 ;
        RECT 66.350 135.500 67.115 135.640 ;
        RECT 66.350 135.440 66.670 135.500 ;
        RECT 66.825 135.455 67.115 135.500 ;
        RECT 34.150 135.100 34.470 135.360 ;
        RECT 38.790 135.300 39.080 135.345 ;
        RECT 40.890 135.300 41.180 135.345 ;
        RECT 42.460 135.300 42.750 135.345 ;
        RECT 64.970 135.300 65.290 135.360 ;
        RECT 38.790 135.160 42.750 135.300 ;
        RECT 38.790 135.115 39.080 135.160 ;
        RECT 40.890 135.115 41.180 135.160 ;
        RECT 42.460 135.115 42.750 135.160 ;
        RECT 59.540 135.160 65.290 135.300 ;
        RECT 59.540 135.020 59.680 135.160 ;
        RECT 64.970 135.100 65.290 135.160 ;
        RECT 39.185 134.960 39.475 135.005 ;
        RECT 40.375 134.960 40.665 135.005 ;
        RECT 42.895 134.960 43.185 135.005 ;
        RECT 39.185 134.820 43.185 134.960 ;
        RECT 39.185 134.775 39.475 134.820 ;
        RECT 40.375 134.775 40.665 134.820 ;
        RECT 42.895 134.775 43.185 134.820 ;
        RECT 48.870 134.960 49.190 135.020 ;
        RECT 52.565 134.960 52.855 135.005 ;
        RECT 48.870 134.820 58.300 134.960 ;
        RECT 48.870 134.760 49.190 134.820 ;
        RECT 52.565 134.775 52.855 134.820 ;
        RECT 30.930 134.620 31.250 134.680 ;
        RECT 31.405 134.620 31.695 134.665 ;
        RECT 30.930 134.480 31.695 134.620 ;
        RECT 30.930 134.420 31.250 134.480 ;
        RECT 31.405 134.435 31.695 134.480 ;
        RECT 31.850 134.620 32.170 134.680 ;
        RECT 35.545 134.620 35.835 134.665 ;
        RECT 31.850 134.480 35.835 134.620 ;
        RECT 31.850 134.420 32.170 134.480 ;
        RECT 35.545 134.435 35.835 134.480 ;
        RECT 36.910 134.620 37.230 134.680 ;
        RECT 38.305 134.620 38.595 134.665 ;
        RECT 42.430 134.620 42.750 134.680 ;
        RECT 36.910 134.480 38.595 134.620 ;
        RECT 36.910 134.420 37.230 134.480 ;
        RECT 38.305 134.435 38.595 134.480 ;
        RECT 38.840 134.480 42.750 134.620 ;
        RECT 34.165 134.280 34.455 134.325 ;
        RECT 34.610 134.280 34.930 134.340 ;
        RECT 34.165 134.140 34.930 134.280 ;
        RECT 34.165 134.095 34.455 134.140 ;
        RECT 34.610 134.080 34.930 134.140 ;
        RECT 35.085 134.280 35.375 134.325 ;
        RECT 38.840 134.280 38.980 134.480 ;
        RECT 42.430 134.420 42.750 134.480 ;
        RECT 53.470 134.420 53.790 134.680 ;
        RECT 58.160 134.665 58.300 134.820 ;
        RECT 59.450 134.760 59.770 135.020 ;
        RECT 59.910 134.760 60.230 135.020 ;
        RECT 58.085 134.620 58.375 134.665 ;
        RECT 61.290 134.620 61.610 134.680 ;
        RECT 58.085 134.480 61.610 134.620 ;
        RECT 58.085 134.435 58.375 134.480 ;
        RECT 61.290 134.420 61.610 134.480 ;
        RECT 61.750 134.420 62.070 134.680 ;
        RECT 62.685 134.435 62.975 134.665 ;
        RECT 39.670 134.325 39.990 134.340 ;
        RECT 35.085 134.140 38.980 134.280 ;
        RECT 35.085 134.095 35.375 134.140 ;
        RECT 39.640 134.095 39.990 134.325 ;
        RECT 60.510 134.280 60.800 134.325 ;
        RECT 62.225 134.280 62.515 134.325 ;
        RECT 60.510 134.140 62.515 134.280 ;
        RECT 62.760 134.280 62.900 134.435 ;
        RECT 63.590 134.420 63.910 134.680 ;
        RECT 64.525 134.620 64.815 134.665 ;
        RECT 65.980 134.620 66.120 135.440 ;
        RECT 66.900 134.960 67.040 135.455 ;
        RECT 68.190 135.440 68.510 135.700 ;
        RECT 69.110 135.640 69.430 135.700 ;
        RECT 73.250 135.640 73.570 135.700 ;
        RECT 73.725 135.640 74.015 135.685 ;
        RECT 69.110 135.500 70.030 135.640 ;
        RECT 69.110 135.440 69.430 135.500 ;
        RECT 69.890 134.960 70.030 135.500 ;
        RECT 73.250 135.500 74.015 135.640 ;
        RECT 73.250 135.440 73.570 135.500 ;
        RECT 73.725 135.455 74.015 135.500 ;
        RECT 100.010 135.360 102.050 136.710 ;
        RECT 103.800 136.700 105.450 136.710 ;
        RECT 102.490 135.430 103.490 136.150 ;
        RECT 103.800 135.890 104.110 136.700 ;
        RECT 104.570 136.420 105.450 136.700 ;
        RECT 105.690 136.880 107.310 137.280 ;
        RECT 108.960 136.930 116.830 137.840 ;
        RECT 104.510 136.190 105.510 136.420 ;
        RECT 105.690 136.230 106.040 136.880 ;
        RECT 106.690 136.870 107.310 136.880 ;
        RECT 108.875 136.700 116.875 136.930 ;
        RECT 108.960 136.690 116.830 136.700 ;
        RECT 104.570 135.980 105.450 136.000 ;
        RECT 103.840 135.600 104.110 135.890 ;
        RECT 104.510 135.750 105.510 135.980 ;
        RECT 105.670 135.940 106.040 136.230 ;
        RECT 105.700 135.880 106.040 135.940 ;
        RECT 106.800 136.550 107.560 136.600 ;
        RECT 108.440 136.550 108.670 136.650 ;
        RECT 106.800 136.340 108.670 136.550 ;
        RECT 117.080 136.340 117.310 136.650 ;
        RECT 106.800 135.920 109.340 136.340 ;
        RECT 116.710 135.920 117.310 136.340 ;
        RECT 104.570 135.600 105.450 135.750 ;
        RECT 104.580 135.430 105.310 135.600 ;
        RECT 71.425 134.960 71.715 135.005 ;
        RECT 66.900 134.820 68.880 134.960 ;
        RECT 64.525 134.480 66.120 134.620 ;
        RECT 68.740 134.620 68.880 134.820 ;
        RECT 69.660 134.820 71.715 134.960 ;
        RECT 69.660 134.665 69.800 134.820 ;
        RECT 71.425 134.775 71.715 134.820 ;
        RECT 69.125 134.620 69.415 134.665 ;
        RECT 68.740 134.480 69.415 134.620 ;
        RECT 64.525 134.435 64.815 134.480 ;
        RECT 69.125 134.435 69.415 134.480 ;
        RECT 69.585 134.435 69.875 134.665 ;
        RECT 71.885 134.435 72.175 134.665 ;
        RECT 66.810 134.325 67.130 134.340 ;
        RECT 64.065 134.280 64.355 134.325 ;
        RECT 62.760 134.140 64.355 134.280 ;
        RECT 60.510 134.095 60.800 134.140 ;
        RECT 62.225 134.095 62.515 134.140 ;
        RECT 64.065 134.095 64.355 134.140 ;
        RECT 66.745 134.095 67.130 134.325 ;
        RECT 29.090 133.940 29.410 134.000 ;
        RECT 35.160 133.940 35.300 134.095 ;
        RECT 39.670 134.080 39.990 134.095 ;
        RECT 66.810 134.080 67.130 134.095 ;
        RECT 67.730 134.280 68.050 134.340 ;
        RECT 68.205 134.280 68.495 134.325 ;
        RECT 67.730 134.140 68.495 134.280 ;
        RECT 69.200 134.280 69.340 134.435 ;
        RECT 71.960 134.280 72.100 134.435 ;
        RECT 69.200 134.140 72.100 134.280 ;
        RECT 67.730 134.080 68.050 134.140 ;
        RECT 68.205 134.095 68.495 134.140 ;
        RECT 29.090 133.800 35.300 133.940 ;
        RECT 45.205 133.940 45.495 133.985 ;
        RECT 47.490 133.940 47.810 134.000 ;
        RECT 45.205 133.800 47.810 133.940 ;
        RECT 29.090 133.740 29.410 133.800 ;
        RECT 45.205 133.755 45.495 133.800 ;
        RECT 47.490 133.740 47.810 133.800 ;
        RECT 61.290 133.740 61.610 134.000 ;
        RECT 13.380 133.120 92.040 133.600 ;
        RECT 25.410 132.920 25.730 132.980 ;
        RECT 27.265 132.920 27.555 132.965 ;
        RECT 25.410 132.780 27.555 132.920 ;
        RECT 25.410 132.720 25.730 132.780 ;
        RECT 27.265 132.735 27.555 132.780 ;
        RECT 28.185 132.920 28.475 132.965 ;
        RECT 31.390 132.920 31.710 132.980 ;
        RECT 28.185 132.780 31.710 132.920 ;
        RECT 28.185 132.735 28.475 132.780 ;
        RECT 31.390 132.720 31.710 132.780 ;
        RECT 40.605 132.920 40.895 132.965 ;
        RECT 53.945 132.920 54.235 132.965 ;
        RECT 54.390 132.920 54.710 132.980 ;
        RECT 40.605 132.780 50.020 132.920 ;
        RECT 40.605 132.735 40.895 132.780 ;
        RECT 39.685 132.580 39.975 132.625 ;
        RECT 48.870 132.580 49.190 132.640 ;
        RECT 39.685 132.440 49.190 132.580 ;
        RECT 49.880 132.580 50.020 132.780 ;
        RECT 53.945 132.780 54.710 132.920 ;
        RECT 53.945 132.735 54.235 132.780 ;
        RECT 54.390 132.720 54.710 132.780 ;
        RECT 63.590 132.920 63.910 132.980 ;
        RECT 64.525 132.920 64.815 132.965 ;
        RECT 63.590 132.780 64.815 132.920 ;
        RECT 63.590 132.720 63.910 132.780 ;
        RECT 64.525 132.735 64.815 132.780 ;
        RECT 67.730 132.920 68.050 132.980 ;
        RECT 73.265 132.920 73.555 132.965 ;
        RECT 67.730 132.780 73.555 132.920 ;
        RECT 67.730 132.720 68.050 132.780 ;
        RECT 73.265 132.735 73.555 132.780 ;
        RECT 53.010 132.580 53.330 132.640 ;
        RECT 53.485 132.580 53.775 132.625 ;
        RECT 49.880 132.440 53.775 132.580 ;
        RECT 39.685 132.395 39.975 132.440 ;
        RECT 48.870 132.380 49.190 132.440 ;
        RECT 53.010 132.380 53.330 132.440 ;
        RECT 53.485 132.395 53.775 132.440 ;
        RECT 58.960 132.580 59.250 132.625 ;
        RECT 61.290 132.580 61.610 132.640 ;
        RECT 69.570 132.580 69.890 132.640 ;
        RECT 74.170 132.580 74.490 132.640 ;
        RECT 76.470 132.580 76.790 132.640 ;
        RECT 58.960 132.440 61.610 132.580 ;
        RECT 58.960 132.395 59.250 132.440 ;
        RECT 61.290 132.380 61.610 132.440 ;
        RECT 66.440 132.440 76.790 132.580 ;
        RECT 41.065 132.240 41.355 132.285 ;
        RECT 42.890 132.240 43.210 132.300 ;
        RECT 41.065 132.100 43.210 132.240 ;
        RECT 41.065 132.055 41.355 132.100 ;
        RECT 42.890 132.040 43.210 132.100 ;
        RECT 46.585 132.240 46.875 132.285 ;
        RECT 47.030 132.240 47.350 132.300 ;
        RECT 46.585 132.100 47.350 132.240 ;
        RECT 46.585 132.055 46.875 132.100 ;
        RECT 47.030 132.040 47.350 132.100 ;
        RECT 47.490 132.040 47.810 132.300 ;
        RECT 49.790 132.040 50.110 132.300 ;
        RECT 54.530 132.240 54.820 132.285 ;
        RECT 51.720 132.100 54.820 132.240 ;
        RECT 30.025 131.900 30.315 131.945 ;
        RECT 30.930 131.900 31.250 131.960 ;
        RECT 30.025 131.760 31.250 131.900 ;
        RECT 30.025 131.715 30.315 131.760 ;
        RECT 30.930 131.700 31.250 131.760 ;
        RECT 35.990 131.700 36.310 131.960 ;
        RECT 46.125 131.900 46.415 131.945 ;
        RECT 47.580 131.900 47.720 132.040 ;
        RECT 46.125 131.760 47.720 131.900 ;
        RECT 46.125 131.715 46.415 131.760 ;
        RECT 50.250 131.700 50.570 131.960 ;
        RECT 51.720 131.945 51.860 132.100 ;
        RECT 54.530 132.055 54.820 132.100 ;
        RECT 57.625 132.240 57.915 132.285 ;
        RECT 58.070 132.240 58.390 132.300 ;
        RECT 66.440 132.285 66.580 132.440 ;
        RECT 69.570 132.380 69.890 132.440 ;
        RECT 74.170 132.380 74.490 132.440 ;
        RECT 76.470 132.380 76.790 132.440 ;
        RECT 67.730 132.285 68.050 132.300 ;
        RECT 57.625 132.100 58.390 132.240 ;
        RECT 57.625 132.055 57.915 132.100 ;
        RECT 58.070 132.040 58.390 132.100 ;
        RECT 66.365 132.055 66.655 132.285 ;
        RECT 67.700 132.055 68.050 132.285 ;
        RECT 67.730 132.040 68.050 132.055 ;
        RECT 51.645 131.715 51.935 131.945 ;
        RECT 52.105 131.715 52.395 131.945 ;
        RECT 58.505 131.900 58.795 131.945 ;
        RECT 59.695 131.900 59.985 131.945 ;
        RECT 62.215 131.900 62.505 131.945 ;
        RECT 58.505 131.760 62.505 131.900 ;
        RECT 58.505 131.715 58.795 131.760 ;
        RECT 59.695 131.715 59.985 131.760 ;
        RECT 62.215 131.715 62.505 131.760 ;
        RECT 67.245 131.900 67.535 131.945 ;
        RECT 68.435 131.900 68.725 131.945 ;
        RECT 70.955 131.900 71.245 131.945 ;
        RECT 67.245 131.760 71.245 131.900 ;
        RECT 67.245 131.715 67.535 131.760 ;
        RECT 68.435 131.715 68.725 131.760 ;
        RECT 70.955 131.715 71.245 131.760 ;
        RECT 100.010 131.720 100.780 135.360 ;
        RECT 102.460 134.310 105.310 135.430 ;
        RECT 105.700 135.130 106.050 135.880 ;
        RECT 106.800 135.760 108.670 135.920 ;
        RECT 106.800 135.710 107.560 135.760 ;
        RECT 108.440 135.690 108.670 135.760 ;
        RECT 117.080 135.690 117.310 135.920 ;
        RECT 108.875 135.410 116.875 135.640 ;
        RECT 105.700 135.070 105.990 135.130 ;
        RECT 105.610 134.950 105.990 135.070 ;
        RECT 108.970 135.010 116.830 135.410 ;
        RECT 117.640 135.010 118.600 144.490 ;
        RECT 119.930 144.620 120.770 146.750 ;
        RECT 126.430 146.330 127.680 146.770 ;
        RECT 137.600 146.750 138.460 148.920 ;
        RECT 124.370 146.320 129.610 146.330 ;
        RECT 121.420 146.220 136.720 146.320 ;
        RECT 121.420 146.210 136.755 146.220 ;
        RECT 121.380 146.090 136.755 146.210 ;
        RECT 121.380 145.980 125.380 146.090 ;
        RECT 126.430 146.010 128.170 146.090 ;
        RECT 128.750 146.010 136.755 146.090 ;
        RECT 126.430 145.930 127.680 146.010 ;
        RECT 128.755 145.990 136.755 146.010 ;
        RECT 120.990 145.680 121.220 145.930 ;
        RECT 125.540 145.790 125.770 145.930 ;
        RECT 128.320 145.790 128.550 145.940 ;
        RECT 125.540 145.680 128.550 145.790 ;
        RECT 136.960 145.680 137.190 145.940 ;
        RECT 120.990 145.240 137.190 145.680 ;
        RECT 120.990 144.970 121.220 145.240 ;
        RECT 125.540 145.210 137.190 145.240 ;
        RECT 125.540 145.120 128.550 145.210 ;
        RECT 125.540 144.970 125.770 145.120 ;
        RECT 128.320 144.980 128.550 145.120 ;
        RECT 136.960 144.980 137.190 145.210 ;
        RECT 121.380 144.690 125.380 144.920 ;
        RECT 128.755 144.710 136.755 144.930 ;
        RECT 137.520 144.710 138.480 146.750 ;
        RECT 128.755 144.700 138.480 144.710 ;
        RECT 121.380 144.620 125.370 144.690 ;
        RECT 119.930 144.510 125.370 144.620 ;
        RECT 128.810 144.540 138.480 144.700 ;
        RECT 119.930 144.420 123.060 144.510 ;
        RECT 136.550 144.490 138.480 144.540 ;
        RECT 119.930 141.150 120.770 144.420 ;
        RECT 124.410 143.960 129.660 143.970 ;
        RECT 124.410 143.850 136.720 143.960 ;
        RECT 121.440 143.790 136.720 143.850 ;
        RECT 121.440 143.780 136.755 143.790 ;
        RECT 121.380 143.650 136.755 143.780 ;
        RECT 121.380 143.640 126.540 143.650 ;
        RECT 121.380 143.550 125.380 143.640 ;
        RECT 128.755 143.560 136.755 143.650 ;
        RECT 128.840 143.550 136.730 143.560 ;
        RECT 120.990 143.190 121.220 143.500 ;
        RECT 121.440 143.190 125.340 143.550 ;
        RECT 125.540 143.190 125.770 143.500 ;
        RECT 120.990 141.850 125.770 143.190 ;
        RECT 120.990 141.540 121.220 141.850 ;
        RECT 125.540 141.540 125.770 141.850 ;
        RECT 128.320 142.970 128.550 143.510 ;
        RECT 129.360 142.970 130.370 143.000 ;
        RECT 136.960 142.970 137.190 143.510 ;
        RECT 128.320 142.070 137.190 142.970 ;
        RECT 128.320 141.550 128.550 142.070 ;
        RECT 129.360 142.000 130.370 142.070 ;
        RECT 136.960 141.550 137.190 142.070 ;
        RECT 121.380 141.260 125.380 141.490 ;
        RECT 128.755 141.270 136.755 141.500 ;
        RECT 119.930 141.110 121.060 141.150 ;
        RECT 119.930 141.030 121.300 141.110 ;
        RECT 121.670 141.040 125.330 141.260 ;
        RECT 121.670 141.030 123.110 141.040 ;
        RECT 119.930 140.990 123.110 141.030 ;
        RECT 119.930 140.900 122.620 140.990 ;
        RECT 128.820 140.980 136.710 141.270 ;
        RECT 119.930 140.840 121.950 140.900 ;
        RECT 119.930 140.790 121.700 140.840 ;
        RECT 119.930 137.450 120.770 140.790 ;
        RECT 128.810 140.490 136.730 140.500 ;
        RECT 125.040 140.480 136.730 140.490 ;
        RECT 121.420 140.360 136.730 140.480 ;
        RECT 121.420 140.350 136.755 140.360 ;
        RECT 121.380 140.230 136.755 140.350 ;
        RECT 121.380 140.120 125.380 140.230 ;
        RECT 120.990 139.780 121.220 140.070 ;
        RECT 121.440 139.780 125.330 140.120 ;
        RECT 125.540 139.780 125.770 140.070 ;
        RECT 120.990 138.410 125.770 139.780 ;
        RECT 120.990 138.110 121.220 138.410 ;
        RECT 125.540 138.110 125.770 138.410 ;
        RECT 121.380 137.830 125.380 138.060 ;
        RECT 121.630 137.600 125.200 137.830 ;
        RECT 121.630 137.450 125.320 137.600 ;
        RECT 119.930 137.170 125.320 137.450 ;
        RECT 126.570 137.280 127.190 140.230 ;
        RECT 128.755 140.130 136.755 140.230 ;
        RECT 128.810 140.120 136.730 140.130 ;
        RECT 128.320 139.420 128.550 140.080 ;
        RECT 129.330 139.420 130.330 139.510 ;
        RECT 136.960 139.420 137.190 140.080 ;
        RECT 128.320 138.600 137.190 139.420 ;
        RECT 128.320 138.120 128.550 138.600 ;
        RECT 129.330 138.510 130.330 138.600 ;
        RECT 136.960 138.120 137.190 138.600 ;
        RECT 128.755 137.840 136.755 138.070 ;
        RECT 119.930 136.710 125.330 137.170 ;
        RECT 119.930 135.370 121.930 136.710 ;
        RECT 123.680 136.700 125.330 136.710 ;
        RECT 122.370 135.430 123.370 136.150 ;
        RECT 123.680 135.890 123.990 136.700 ;
        RECT 124.450 136.420 125.330 136.700 ;
        RECT 125.570 136.880 127.190 137.280 ;
        RECT 128.840 136.930 136.710 137.840 ;
        RECT 124.390 136.190 125.390 136.420 ;
        RECT 125.570 136.230 125.920 136.880 ;
        RECT 126.570 136.870 127.190 136.880 ;
        RECT 128.755 136.700 136.755 136.930 ;
        RECT 128.840 136.690 136.710 136.700 ;
        RECT 124.450 135.980 125.330 136.000 ;
        RECT 123.720 135.600 123.990 135.890 ;
        RECT 124.390 135.750 125.390 135.980 ;
        RECT 125.550 135.940 125.920 136.230 ;
        RECT 125.580 135.880 125.920 135.940 ;
        RECT 126.680 136.550 127.440 136.600 ;
        RECT 128.320 136.550 128.550 136.650 ;
        RECT 126.680 136.340 128.550 136.550 ;
        RECT 136.960 136.340 137.190 136.650 ;
        RECT 126.680 135.920 129.220 136.340 ;
        RECT 136.590 135.920 137.190 136.340 ;
        RECT 124.450 135.600 125.330 135.750 ;
        RECT 124.460 135.430 125.190 135.600 ;
        RECT 102.400 134.080 105.400 134.310 ;
        RECT 105.610 134.120 105.950 134.950 ;
        RECT 107.960 134.940 118.600 135.010 ;
        RECT 102.450 134.050 105.310 134.080 ;
        RECT 102.450 134.030 103.620 134.050 ;
        RECT 104.580 134.040 105.310 134.050 ;
        RECT 102.400 133.640 105.400 133.870 ;
        RECT 105.605 133.830 105.950 134.120 ;
        RECT 106.140 133.900 118.600 134.940 ;
        RECT 120.000 135.360 121.930 135.370 ;
        RECT 106.140 133.880 118.560 133.900 ;
        RECT 105.610 133.720 105.950 133.830 ;
        RECT 106.180 133.870 111.850 133.880 ;
        RECT 112.850 133.870 118.560 133.880 ;
        RECT 102.490 133.470 105.350 133.640 ;
        RECT 106.180 133.470 106.610 133.870 ;
        RECT 102.460 133.100 106.610 133.470 ;
        RECT 39.670 131.360 39.990 131.620 ;
        RECT 48.870 131.560 49.190 131.620 ;
        RECT 52.180 131.560 52.320 131.715 ;
        RECT 48.870 131.420 52.320 131.560 ;
        RECT 58.110 131.560 58.400 131.605 ;
        RECT 60.210 131.560 60.500 131.605 ;
        RECT 61.780 131.560 62.070 131.605 ;
        RECT 58.110 131.420 62.070 131.560 ;
        RECT 48.870 131.360 49.190 131.420 ;
        RECT 58.110 131.375 58.400 131.420 ;
        RECT 60.210 131.375 60.500 131.420 ;
        RECT 61.780 131.375 62.070 131.420 ;
        RECT 66.850 131.560 67.140 131.605 ;
        RECT 68.950 131.560 69.240 131.605 ;
        RECT 70.520 131.560 70.810 131.605 ;
        RECT 66.850 131.420 70.810 131.560 ;
        RECT 66.850 131.375 67.140 131.420 ;
        RECT 68.950 131.375 69.240 131.420 ;
        RECT 70.520 131.375 70.810 131.420 ;
        RECT 28.185 131.220 28.475 131.265 ;
        RECT 29.090 131.220 29.410 131.280 ;
        RECT 28.185 131.080 29.410 131.220 ;
        RECT 28.185 131.035 28.475 131.080 ;
        RECT 29.090 131.020 29.410 131.080 ;
        RECT 31.390 131.220 31.710 131.280 ;
        RECT 34.165 131.220 34.455 131.265 ;
        RECT 34.610 131.220 34.930 131.280 ;
        RECT 31.390 131.080 34.930 131.220 ;
        RECT 31.390 131.020 31.710 131.080 ;
        RECT 34.165 131.035 34.455 131.080 ;
        RECT 34.610 131.020 34.930 131.080 ;
        RECT 37.830 131.220 38.150 131.280 ;
        RECT 38.765 131.220 39.055 131.265 ;
        RECT 37.830 131.080 39.055 131.220 ;
        RECT 37.830 131.020 38.150 131.080 ;
        RECT 38.765 131.035 39.055 131.080 ;
        RECT 42.890 131.020 43.210 131.280 ;
        RECT 45.650 131.220 45.970 131.280 ;
        RECT 47.045 131.220 47.335 131.265 ;
        RECT 45.650 131.080 47.335 131.220 ;
        RECT 45.650 131.020 45.970 131.080 ;
        RECT 47.045 131.035 47.335 131.080 ;
        RECT 55.310 131.020 55.630 131.280 ;
        RECT 13.380 130.400 92.040 130.880 ;
        RECT 60.830 130.000 61.150 130.260 ;
        RECT 67.730 130.200 68.050 130.260 ;
        RECT 68.665 130.200 68.955 130.245 ;
        RECT 67.730 130.060 68.955 130.200 ;
        RECT 67.730 130.000 68.050 130.060 ;
        RECT 68.665 130.015 68.955 130.060 ;
        RECT 29.550 129.860 29.840 129.905 ;
        RECT 31.120 129.860 31.410 129.905 ;
        RECT 33.220 129.860 33.510 129.905 ;
        RECT 29.550 129.720 33.510 129.860 ;
        RECT 29.550 129.675 29.840 129.720 ;
        RECT 31.120 129.675 31.410 129.720 ;
        RECT 33.220 129.675 33.510 129.720 ;
        RECT 36.950 129.860 37.240 129.905 ;
        RECT 39.050 129.860 39.340 129.905 ;
        RECT 40.620 129.860 40.910 129.905 ;
        RECT 36.950 129.720 40.910 129.860 ;
        RECT 36.950 129.675 37.240 129.720 ;
        RECT 39.050 129.675 39.340 129.720 ;
        RECT 40.620 129.675 40.910 129.720 ;
        RECT 42.430 129.860 42.750 129.920 ;
        RECT 47.045 129.860 47.335 129.905 ;
        RECT 42.430 129.720 47.335 129.860 ;
        RECT 42.430 129.660 42.750 129.720 ;
        RECT 47.045 129.675 47.335 129.720 ;
        RECT 54.430 129.860 54.720 129.905 ;
        RECT 56.530 129.860 56.820 129.905 ;
        RECT 58.100 129.860 58.390 129.905 ;
        RECT 70.030 129.860 70.350 129.920 ;
        RECT 54.430 129.720 58.390 129.860 ;
        RECT 54.430 129.675 54.720 129.720 ;
        RECT 56.530 129.675 56.820 129.720 ;
        RECT 58.100 129.675 58.390 129.720 ;
        RECT 65.520 129.720 70.350 129.860 ;
        RECT 29.115 129.520 29.405 129.565 ;
        RECT 31.635 129.520 31.925 129.565 ;
        RECT 32.825 129.520 33.115 129.565 ;
        RECT 34.150 129.520 34.470 129.580 ;
        RECT 29.115 129.380 33.115 129.520 ;
        RECT 29.115 129.335 29.405 129.380 ;
        RECT 31.635 129.335 31.925 129.380 ;
        RECT 32.825 129.335 33.115 129.380 ;
        RECT 33.320 129.380 34.470 129.520 ;
        RECT 32.425 129.180 32.715 129.225 ;
        RECT 33.320 129.180 33.460 129.380 ;
        RECT 34.150 129.320 34.470 129.380 ;
        RECT 37.345 129.520 37.635 129.565 ;
        RECT 38.535 129.520 38.825 129.565 ;
        RECT 41.055 129.520 41.345 129.565 ;
        RECT 46.125 129.520 46.415 129.565 ;
        RECT 37.345 129.380 41.345 129.520 ;
        RECT 37.345 129.335 37.635 129.380 ;
        RECT 38.535 129.335 38.825 129.380 ;
        RECT 41.055 129.335 41.345 129.380 ;
        RECT 44.820 129.380 46.415 129.520 ;
        RECT 32.425 129.040 33.460 129.180 ;
        RECT 33.705 129.180 33.995 129.225 ;
        RECT 36.465 129.180 36.755 129.225 ;
        RECT 36.910 129.180 37.230 129.240 ;
        RECT 37.830 129.225 38.150 129.240 ;
        RECT 37.800 129.180 38.150 129.225 ;
        RECT 40.590 129.180 40.910 129.240 ;
        RECT 33.705 129.040 37.230 129.180 ;
        RECT 37.635 129.040 38.150 129.180 ;
        RECT 32.425 128.995 32.715 129.040 ;
        RECT 33.705 128.995 33.995 129.040 ;
        RECT 36.465 128.995 36.755 129.040 ;
        RECT 36.910 128.980 37.230 129.040 ;
        RECT 37.800 128.995 38.150 129.040 ;
        RECT 37.830 128.980 38.150 128.995 ;
        RECT 38.840 129.040 40.910 129.180 ;
        RECT 28.630 128.840 28.950 128.900 ;
        RECT 35.085 128.840 35.375 128.885 ;
        RECT 28.630 128.700 35.375 128.840 ;
        RECT 28.630 128.640 28.950 128.700 ;
        RECT 35.085 128.655 35.375 128.700 ;
        RECT 36.005 128.840 36.295 128.885 ;
        RECT 38.840 128.840 38.980 129.040 ;
        RECT 40.590 128.980 40.910 129.040 ;
        RECT 43.350 129.180 43.670 129.240 ;
        RECT 44.285 129.180 44.575 129.225 ;
        RECT 43.350 129.040 44.575 129.180 ;
        RECT 43.350 128.980 43.670 129.040 ;
        RECT 44.285 128.995 44.575 129.040 ;
        RECT 43.825 128.840 44.115 128.885 ;
        RECT 36.005 128.700 38.980 128.840 ;
        RECT 39.300 128.700 44.115 128.840 ;
        RECT 36.005 128.655 36.295 128.700 ;
        RECT 26.790 128.300 27.110 128.560 ;
        RECT 34.165 128.500 34.455 128.545 ;
        RECT 39.300 128.500 39.440 128.700 ;
        RECT 43.825 128.655 44.115 128.700 ;
        RECT 34.165 128.360 39.440 128.500 ;
        RECT 40.590 128.500 40.910 128.560 ;
        RECT 43.365 128.500 43.655 128.545 ;
        RECT 44.820 128.500 44.960 129.380 ;
        RECT 46.125 129.335 46.415 129.380 ;
        RECT 47.490 129.520 47.810 129.580 ;
        RECT 65.520 129.565 65.660 129.720 ;
        RECT 70.030 129.660 70.350 129.720 ;
        RECT 100.010 129.620 100.880 131.720 ;
        RECT 106.550 131.330 107.800 131.770 ;
        RECT 117.700 131.750 118.560 133.870 ;
        RECT 120.000 131.810 120.770 135.360 ;
        RECT 122.340 134.310 125.190 135.430 ;
        RECT 125.580 135.130 125.930 135.880 ;
        RECT 126.680 135.760 128.550 135.920 ;
        RECT 126.680 135.710 127.440 135.760 ;
        RECT 128.320 135.690 128.550 135.760 ;
        RECT 136.960 135.690 137.190 135.920 ;
        RECT 128.755 135.410 136.755 135.640 ;
        RECT 125.580 135.070 125.870 135.130 ;
        RECT 125.490 134.950 125.870 135.070 ;
        RECT 128.850 135.010 136.710 135.410 ;
        RECT 137.520 135.010 138.480 144.490 ;
        RECT 122.280 134.080 125.280 134.310 ;
        RECT 125.490 134.120 125.830 134.950 ;
        RECT 127.840 134.940 138.480 135.010 ;
        RECT 122.330 134.050 125.190 134.080 ;
        RECT 122.330 134.030 123.500 134.050 ;
        RECT 124.460 134.040 125.190 134.050 ;
        RECT 122.280 133.640 125.280 133.870 ;
        RECT 125.485 133.830 125.830 134.120 ;
        RECT 126.020 133.900 138.480 134.940 ;
        RECT 139.930 146.720 140.700 150.360 ;
        RECT 142.420 149.310 145.270 150.430 ;
        RECT 145.660 150.130 146.010 150.880 ;
        RECT 146.760 150.760 148.630 150.920 ;
        RECT 146.760 150.710 147.520 150.760 ;
        RECT 148.400 150.690 148.630 150.760 ;
        RECT 157.040 150.690 157.270 150.920 ;
        RECT 148.835 150.410 156.835 150.640 ;
        RECT 145.660 150.070 145.950 150.130 ;
        RECT 145.570 149.950 145.950 150.070 ;
        RECT 148.930 150.010 156.790 150.410 ;
        RECT 157.600 150.010 158.560 159.490 ;
        RECT 142.360 149.080 145.360 149.310 ;
        RECT 145.570 149.120 145.910 149.950 ;
        RECT 147.920 149.940 158.560 150.010 ;
        RECT 142.410 149.050 145.270 149.080 ;
        RECT 142.410 149.030 143.580 149.050 ;
        RECT 144.540 149.040 145.270 149.050 ;
        RECT 142.360 148.640 145.360 148.870 ;
        RECT 145.565 148.830 145.910 149.120 ;
        RECT 146.100 148.900 158.560 149.940 ;
        RECT 146.100 148.880 158.500 148.900 ;
        RECT 145.570 148.720 145.910 148.830 ;
        RECT 146.140 148.870 151.810 148.880 ;
        RECT 152.810 148.870 158.500 148.880 ;
        RECT 142.450 148.470 145.310 148.640 ;
        RECT 146.140 148.470 146.570 148.870 ;
        RECT 142.420 148.100 146.570 148.470 ;
        RECT 139.930 144.620 140.790 146.720 ;
        RECT 146.460 146.330 147.710 146.770 ;
        RECT 157.640 146.750 158.500 148.870 ;
        RECT 144.400 146.320 149.640 146.330 ;
        RECT 141.450 146.220 156.750 146.320 ;
        RECT 141.450 146.210 156.785 146.220 ;
        RECT 141.410 146.090 156.785 146.210 ;
        RECT 141.410 145.980 145.410 146.090 ;
        RECT 146.460 146.010 148.200 146.090 ;
        RECT 148.780 146.010 156.785 146.090 ;
        RECT 146.460 145.930 147.710 146.010 ;
        RECT 148.785 145.990 156.785 146.010 ;
        RECT 141.020 145.680 141.250 145.930 ;
        RECT 145.570 145.790 145.800 145.930 ;
        RECT 148.350 145.790 148.580 145.940 ;
        RECT 145.570 145.680 148.580 145.790 ;
        RECT 156.990 145.680 157.220 145.940 ;
        RECT 141.020 145.240 157.220 145.680 ;
        RECT 141.020 144.970 141.250 145.240 ;
        RECT 145.570 145.210 157.220 145.240 ;
        RECT 145.570 145.120 148.580 145.210 ;
        RECT 145.570 144.970 145.800 145.120 ;
        RECT 148.350 144.980 148.580 145.120 ;
        RECT 156.990 144.980 157.220 145.210 ;
        RECT 141.410 144.690 145.410 144.920 ;
        RECT 148.785 144.710 156.785 144.930 ;
        RECT 157.550 144.710 158.510 146.750 ;
        RECT 148.785 144.700 158.510 144.710 ;
        RECT 141.410 144.620 145.400 144.690 ;
        RECT 139.930 144.510 145.400 144.620 ;
        RECT 148.840 144.540 158.510 144.700 ;
        RECT 139.930 144.420 143.090 144.510 ;
        RECT 156.580 144.490 158.510 144.540 ;
        RECT 139.930 141.150 140.790 144.420 ;
        RECT 144.440 143.960 149.690 143.970 ;
        RECT 144.440 143.850 156.750 143.960 ;
        RECT 141.470 143.790 156.750 143.850 ;
        RECT 141.470 143.780 156.785 143.790 ;
        RECT 141.410 143.650 156.785 143.780 ;
        RECT 141.410 143.640 146.570 143.650 ;
        RECT 141.410 143.550 145.410 143.640 ;
        RECT 148.785 143.560 156.785 143.650 ;
        RECT 148.870 143.550 156.760 143.560 ;
        RECT 141.020 143.190 141.250 143.500 ;
        RECT 141.470 143.190 145.370 143.550 ;
        RECT 145.570 143.190 145.800 143.500 ;
        RECT 141.020 141.850 145.800 143.190 ;
        RECT 141.020 141.540 141.250 141.850 ;
        RECT 145.570 141.540 145.800 141.850 ;
        RECT 148.350 142.970 148.580 143.510 ;
        RECT 149.390 142.970 150.400 143.000 ;
        RECT 156.990 142.970 157.220 143.510 ;
        RECT 148.350 142.070 157.220 142.970 ;
        RECT 148.350 141.550 148.580 142.070 ;
        RECT 149.390 142.000 150.400 142.070 ;
        RECT 156.990 141.550 157.220 142.070 ;
        RECT 141.410 141.260 145.410 141.490 ;
        RECT 148.785 141.270 156.785 141.500 ;
        RECT 139.930 141.110 141.090 141.150 ;
        RECT 139.930 141.030 141.330 141.110 ;
        RECT 141.700 141.040 145.360 141.260 ;
        RECT 141.700 141.030 143.140 141.040 ;
        RECT 139.930 140.990 143.140 141.030 ;
        RECT 139.930 140.900 142.650 140.990 ;
        RECT 148.850 140.980 156.740 141.270 ;
        RECT 139.930 140.840 141.980 140.900 ;
        RECT 139.930 140.790 141.730 140.840 ;
        RECT 139.930 137.450 140.790 140.790 ;
        RECT 148.840 140.490 156.760 140.500 ;
        RECT 145.070 140.480 156.760 140.490 ;
        RECT 141.450 140.360 156.760 140.480 ;
        RECT 141.450 140.350 156.785 140.360 ;
        RECT 141.410 140.230 156.785 140.350 ;
        RECT 141.410 140.120 145.410 140.230 ;
        RECT 141.020 139.780 141.250 140.070 ;
        RECT 141.470 139.780 145.360 140.120 ;
        RECT 145.570 139.780 145.800 140.070 ;
        RECT 141.020 138.410 145.800 139.780 ;
        RECT 141.020 138.110 141.250 138.410 ;
        RECT 145.570 138.110 145.800 138.410 ;
        RECT 141.410 137.830 145.410 138.060 ;
        RECT 141.660 137.600 145.230 137.830 ;
        RECT 141.660 137.450 145.350 137.600 ;
        RECT 139.930 137.170 145.350 137.450 ;
        RECT 146.600 137.280 147.220 140.230 ;
        RECT 148.785 140.130 156.785 140.230 ;
        RECT 148.840 140.120 156.760 140.130 ;
        RECT 148.350 139.420 148.580 140.080 ;
        RECT 149.360 139.420 150.360 139.510 ;
        RECT 156.990 139.420 157.220 140.080 ;
        RECT 148.350 138.600 157.220 139.420 ;
        RECT 148.350 138.120 148.580 138.600 ;
        RECT 149.360 138.510 150.360 138.600 ;
        RECT 156.990 138.120 157.220 138.600 ;
        RECT 148.785 137.840 156.785 138.070 ;
        RECT 139.930 136.710 145.360 137.170 ;
        RECT 139.930 135.360 141.960 136.710 ;
        RECT 143.710 136.700 145.360 136.710 ;
        RECT 142.400 135.430 143.400 136.150 ;
        RECT 143.710 135.890 144.020 136.700 ;
        RECT 144.480 136.420 145.360 136.700 ;
        RECT 145.600 136.880 147.220 137.280 ;
        RECT 148.870 136.930 156.740 137.840 ;
        RECT 144.420 136.190 145.420 136.420 ;
        RECT 145.600 136.230 145.950 136.880 ;
        RECT 146.600 136.870 147.220 136.880 ;
        RECT 148.785 136.700 156.785 136.930 ;
        RECT 148.870 136.690 156.740 136.700 ;
        RECT 144.480 135.980 145.360 136.000 ;
        RECT 143.750 135.600 144.020 135.890 ;
        RECT 144.420 135.750 145.420 135.980 ;
        RECT 145.580 135.940 145.950 136.230 ;
        RECT 145.610 135.880 145.950 135.940 ;
        RECT 146.710 136.550 147.470 136.600 ;
        RECT 148.350 136.550 148.580 136.650 ;
        RECT 146.710 136.340 148.580 136.550 ;
        RECT 156.990 136.340 157.220 136.650 ;
        RECT 146.710 135.920 149.250 136.340 ;
        RECT 156.620 135.920 157.220 136.340 ;
        RECT 144.480 135.600 145.360 135.750 ;
        RECT 144.490 135.430 145.220 135.600 ;
        RECT 126.020 133.880 138.460 133.900 ;
        RECT 125.490 133.720 125.830 133.830 ;
        RECT 126.060 133.870 131.730 133.880 ;
        RECT 132.730 133.870 138.460 133.880 ;
        RECT 122.370 133.470 125.230 133.640 ;
        RECT 126.060 133.470 126.490 133.870 ;
        RECT 122.340 133.100 126.490 133.470 ;
        RECT 104.490 131.320 109.730 131.330 ;
        RECT 101.540 131.220 116.840 131.320 ;
        RECT 101.540 131.210 116.875 131.220 ;
        RECT 101.500 131.090 116.875 131.210 ;
        RECT 101.500 130.980 105.500 131.090 ;
        RECT 106.550 131.010 108.290 131.090 ;
        RECT 108.870 131.010 116.875 131.090 ;
        RECT 106.550 130.930 107.800 131.010 ;
        RECT 108.875 130.990 116.875 131.010 ;
        RECT 101.110 130.680 101.340 130.930 ;
        RECT 105.660 130.790 105.890 130.930 ;
        RECT 108.440 130.790 108.670 130.940 ;
        RECT 105.660 130.680 108.670 130.790 ;
        RECT 117.080 130.680 117.310 130.940 ;
        RECT 101.110 130.240 117.310 130.680 ;
        RECT 101.110 129.970 101.340 130.240 ;
        RECT 105.660 130.210 117.310 130.240 ;
        RECT 105.660 130.120 108.670 130.210 ;
        RECT 105.660 129.970 105.890 130.120 ;
        RECT 108.440 129.980 108.670 130.120 ;
        RECT 117.080 129.980 117.310 130.210 ;
        RECT 101.500 129.690 105.500 129.920 ;
        RECT 108.875 129.710 116.875 129.930 ;
        RECT 117.640 129.710 118.600 131.750 ;
        RECT 108.875 129.700 118.600 129.710 ;
        RECT 101.500 129.620 105.490 129.690 ;
        RECT 54.825 129.520 55.115 129.565 ;
        RECT 56.015 129.520 56.305 129.565 ;
        RECT 58.535 129.520 58.825 129.565 ;
        RECT 47.490 129.380 53.700 129.520 ;
        RECT 45.650 128.980 45.970 129.240 ;
        RECT 46.200 129.180 46.340 129.335 ;
        RECT 47.490 129.320 47.810 129.380 ;
        RECT 49.330 129.180 49.650 129.240 ;
        RECT 53.560 129.225 53.700 129.380 ;
        RECT 54.825 129.380 58.825 129.520 ;
        RECT 54.825 129.335 55.115 129.380 ;
        RECT 56.015 129.335 56.305 129.380 ;
        RECT 58.535 129.335 58.825 129.380 ;
        RECT 65.445 129.335 65.735 129.565 ;
        RECT 67.870 129.520 68.160 129.565 ;
        RECT 68.650 129.520 68.970 129.580 ;
        RECT 67.870 129.380 68.970 129.520 ;
        RECT 67.870 129.335 68.160 129.380 ;
        RECT 68.650 129.320 68.970 129.380 ;
        RECT 100.010 129.510 105.490 129.620 ;
        RECT 108.930 129.540 118.600 129.700 ;
        RECT 100.010 129.420 103.180 129.510 ;
        RECT 116.670 129.490 118.600 129.540 ;
        RECT 50.265 129.180 50.555 129.225 ;
        RECT 52.565 129.180 52.855 129.225 ;
        RECT 46.200 129.040 52.855 129.180 ;
        RECT 49.330 128.980 49.650 129.040 ;
        RECT 50.265 128.995 50.555 129.040 ;
        RECT 52.565 128.995 52.855 129.040 ;
        RECT 53.485 128.995 53.775 129.225 ;
        RECT 53.945 129.180 54.235 129.225 ;
        RECT 58.070 129.180 58.390 129.240 ;
        RECT 53.945 129.040 58.390 129.180 ;
        RECT 53.945 128.995 54.235 129.040 ;
        RECT 58.070 128.980 58.390 129.040 ;
        RECT 64.970 129.180 65.290 129.240 ;
        RECT 66.825 129.180 67.115 129.225 ;
        RECT 64.970 129.040 67.115 129.180 ;
        RECT 64.970 128.980 65.290 129.040 ;
        RECT 66.825 128.995 67.115 129.040 ;
        RECT 45.190 128.840 45.510 128.900 ;
        RECT 55.310 128.885 55.630 128.900 ;
        RECT 47.505 128.840 47.795 128.885 ;
        RECT 55.280 128.840 55.630 128.885 ;
        RECT 45.190 128.700 47.795 128.840 ;
        RECT 55.115 128.700 55.630 128.840 ;
        RECT 45.190 128.640 45.510 128.700 ;
        RECT 47.505 128.655 47.795 128.700 ;
        RECT 55.280 128.655 55.630 128.700 ;
        RECT 55.310 128.640 55.630 128.655 ;
        RECT 40.590 128.360 44.960 128.500 ;
        RECT 46.110 128.500 46.430 128.560 ;
        RECT 49.790 128.500 50.110 128.560 ;
        RECT 52.565 128.500 52.855 128.545 ;
        RECT 46.110 128.360 52.855 128.500 ;
        RECT 34.165 128.315 34.455 128.360 ;
        RECT 40.590 128.300 40.910 128.360 ;
        RECT 43.365 128.315 43.655 128.360 ;
        RECT 46.110 128.300 46.430 128.360 ;
        RECT 49.790 128.300 50.110 128.360 ;
        RECT 52.565 128.315 52.855 128.360 ;
        RECT 54.390 128.500 54.710 128.560 ;
        RECT 67.285 128.500 67.575 128.545 ;
        RECT 54.390 128.360 67.575 128.500 ;
        RECT 54.390 128.300 54.710 128.360 ;
        RECT 67.285 128.315 67.575 128.360 ;
        RECT 13.380 127.680 92.040 128.160 ;
        RECT 28.630 127.280 28.950 127.540 ;
        RECT 35.990 127.280 36.310 127.540 ;
        RECT 47.505 127.295 47.795 127.525 ;
        RECT 45.650 127.140 45.970 127.200 ;
        RECT 37.460 127.000 45.970 127.140 ;
        RECT 34.265 126.800 34.555 126.845 ;
        RECT 35.070 126.800 35.390 126.860 ;
        RECT 34.265 126.660 35.390 126.800 ;
        RECT 34.265 126.615 34.555 126.660 ;
        RECT 35.070 126.600 35.390 126.660 ;
        RECT 37.460 126.520 37.600 127.000 ;
        RECT 45.650 126.940 45.970 127.000 ;
        RECT 37.845 126.800 38.135 126.845 ;
        RECT 45.190 126.800 45.510 126.860 ;
        RECT 37.845 126.660 45.510 126.800 ;
        RECT 37.845 126.615 38.135 126.660 ;
        RECT 45.190 126.600 45.510 126.660 ;
        RECT 46.110 126.600 46.430 126.860 ;
        RECT 47.580 126.800 47.720 127.295 ;
        RECT 49.245 126.800 49.535 126.845 ;
        RECT 47.580 126.660 49.535 126.800 ;
        RECT 49.245 126.615 49.535 126.660 ;
        RECT 30.955 126.460 31.245 126.505 ;
        RECT 33.475 126.460 33.765 126.505 ;
        RECT 34.665 126.460 34.955 126.505 ;
        RECT 30.955 126.320 34.955 126.460 ;
        RECT 30.955 126.275 31.245 126.320 ;
        RECT 33.475 126.275 33.765 126.320 ;
        RECT 34.665 126.275 34.955 126.320 ;
        RECT 35.545 126.275 35.835 126.505 ;
        RECT 31.390 126.120 31.680 126.165 ;
        RECT 32.960 126.120 33.250 126.165 ;
        RECT 35.060 126.120 35.350 126.165 ;
        RECT 31.390 125.980 35.350 126.120 ;
        RECT 35.620 126.120 35.760 126.275 ;
        RECT 37.370 126.260 37.690 126.520 ;
        RECT 40.130 126.460 40.450 126.520 ;
        RECT 40.605 126.460 40.895 126.505 ;
        RECT 40.130 126.320 40.895 126.460 ;
        RECT 40.130 126.260 40.450 126.320 ;
        RECT 40.605 126.275 40.895 126.320 ;
        RECT 41.970 126.460 42.290 126.520 ;
        RECT 44.270 126.460 44.590 126.520 ;
        RECT 41.970 126.320 44.590 126.460 ;
        RECT 41.970 126.260 42.290 126.320 ;
        RECT 44.270 126.260 44.590 126.320 ;
        RECT 44.745 126.460 45.035 126.505 ;
        RECT 45.650 126.460 45.970 126.520 ;
        RECT 44.745 126.320 45.970 126.460 ;
        RECT 44.745 126.275 45.035 126.320 ;
        RECT 45.650 126.260 45.970 126.320 ;
        RECT 46.570 126.260 46.890 126.520 ;
        RECT 47.965 126.275 48.255 126.505 ;
        RECT 48.845 126.460 49.135 126.505 ;
        RECT 50.035 126.460 50.325 126.505 ;
        RECT 52.555 126.460 52.845 126.505 ;
        RECT 48.845 126.320 52.845 126.460 ;
        RECT 48.845 126.275 49.135 126.320 ;
        RECT 50.035 126.275 50.325 126.320 ;
        RECT 52.555 126.275 52.845 126.320 ;
        RECT 36.910 126.120 37.230 126.180 ;
        RECT 48.040 126.120 48.180 126.275 ;
        RECT 35.620 125.980 48.180 126.120 ;
        RECT 48.450 126.120 48.740 126.165 ;
        RECT 50.550 126.120 50.840 126.165 ;
        RECT 52.120 126.120 52.410 126.165 ;
        RECT 48.450 125.980 52.410 126.120 ;
        RECT 31.390 125.935 31.680 125.980 ;
        RECT 32.960 125.935 33.250 125.980 ;
        RECT 35.060 125.935 35.350 125.980 ;
        RECT 36.910 125.920 37.230 125.980 ;
        RECT 44.820 125.840 44.960 125.980 ;
        RECT 48.450 125.935 48.740 125.980 ;
        RECT 50.550 125.935 50.840 125.980 ;
        RECT 52.120 125.935 52.410 125.980 ;
        RECT 53.470 126.120 53.790 126.180 ;
        RECT 54.865 126.120 55.155 126.165 ;
        RECT 53.470 125.980 55.155 126.120 ;
        RECT 53.470 125.920 53.790 125.980 ;
        RECT 54.865 125.935 55.155 125.980 ;
        RECT 100.010 126.150 100.880 129.420 ;
        RECT 104.530 128.960 109.780 128.970 ;
        RECT 104.530 128.850 116.840 128.960 ;
        RECT 101.560 128.790 116.840 128.850 ;
        RECT 101.560 128.780 116.875 128.790 ;
        RECT 101.500 128.650 116.875 128.780 ;
        RECT 101.500 128.640 106.660 128.650 ;
        RECT 101.500 128.550 105.500 128.640 ;
        RECT 108.875 128.560 116.875 128.650 ;
        RECT 108.960 128.550 116.850 128.560 ;
        RECT 101.110 128.190 101.340 128.500 ;
        RECT 101.560 128.190 105.460 128.550 ;
        RECT 105.660 128.190 105.890 128.500 ;
        RECT 101.110 126.850 105.890 128.190 ;
        RECT 101.110 126.540 101.340 126.850 ;
        RECT 105.660 126.540 105.890 126.850 ;
        RECT 108.440 127.970 108.670 128.510 ;
        RECT 109.480 127.970 110.490 128.000 ;
        RECT 117.080 127.970 117.310 128.510 ;
        RECT 108.440 127.070 117.310 127.970 ;
        RECT 108.440 126.550 108.670 127.070 ;
        RECT 109.480 127.000 110.490 127.070 ;
        RECT 117.080 126.550 117.310 127.070 ;
        RECT 101.500 126.260 105.500 126.490 ;
        RECT 108.875 126.270 116.875 126.500 ;
        RECT 100.010 126.110 101.180 126.150 ;
        RECT 100.010 126.030 101.420 126.110 ;
        RECT 101.790 126.040 105.450 126.260 ;
        RECT 101.790 126.030 103.230 126.040 ;
        RECT 100.010 125.990 103.230 126.030 ;
        RECT 100.010 125.900 102.740 125.990 ;
        RECT 108.940 125.980 116.830 126.270 ;
        RECT 100.010 125.840 102.070 125.900 ;
        RECT 39.670 125.780 39.990 125.840 ;
        RECT 41.970 125.780 42.290 125.840 ;
        RECT 39.670 125.640 42.290 125.780 ;
        RECT 39.670 125.580 39.990 125.640 ;
        RECT 41.970 125.580 42.290 125.640 ;
        RECT 43.810 125.580 44.130 125.840 ;
        RECT 44.730 125.580 45.050 125.840 ;
        RECT 45.650 125.780 45.970 125.840 ;
        RECT 48.870 125.780 49.190 125.840 ;
        RECT 45.650 125.640 49.190 125.780 ;
        RECT 45.650 125.580 45.970 125.640 ;
        RECT 48.870 125.580 49.190 125.640 ;
        RECT 100.010 125.790 101.820 125.840 ;
        RECT 13.380 124.960 92.040 125.440 ;
        RECT 35.070 124.560 35.390 124.820 ;
        RECT 40.130 124.560 40.450 124.820 ;
        RECT 40.605 124.760 40.895 124.805 ;
        RECT 42.890 124.760 43.210 124.820 ;
        RECT 40.605 124.620 43.210 124.760 ;
        RECT 40.605 124.575 40.895 124.620 ;
        RECT 42.890 124.560 43.210 124.620 ;
        RECT 45.190 124.760 45.510 124.820 ;
        RECT 47.030 124.760 47.350 124.820 ;
        RECT 48.410 124.760 48.730 124.820 ;
        RECT 48.885 124.760 49.175 124.805 ;
        RECT 45.190 124.620 46.295 124.760 ;
        RECT 45.190 124.560 45.510 124.620 ;
        RECT 36.465 124.420 36.755 124.465 ;
        RECT 37.370 124.420 37.690 124.480 ;
        RECT 36.465 124.280 37.690 124.420 ;
        RECT 36.465 124.235 36.755 124.280 ;
        RECT 37.370 124.220 37.690 124.280 ;
        RECT 41.510 124.220 41.830 124.480 ;
        RECT 42.010 124.420 42.300 124.465 ;
        RECT 44.110 124.420 44.400 124.465 ;
        RECT 45.680 124.420 45.970 124.465 ;
        RECT 42.010 124.280 45.970 124.420 ;
        RECT 46.155 124.420 46.295 124.620 ;
        RECT 47.030 124.620 49.175 124.760 ;
        RECT 47.030 124.560 47.350 124.620 ;
        RECT 48.410 124.560 48.730 124.620 ;
        RECT 48.885 124.575 49.175 124.620 ;
        RECT 53.945 124.420 54.235 124.465 ;
        RECT 46.155 124.280 54.235 124.420 ;
        RECT 42.010 124.235 42.300 124.280 ;
        RECT 44.110 124.235 44.400 124.280 ;
        RECT 45.680 124.235 45.970 124.280 ;
        RECT 53.945 124.235 54.235 124.280 ;
        RECT 26.790 124.080 27.110 124.140 ;
        RECT 28.185 124.080 28.475 124.125 ;
        RECT 26.790 123.940 28.475 124.080 ;
        RECT 26.790 123.880 27.110 123.940 ;
        RECT 28.185 123.895 28.475 123.940 ;
        RECT 36.910 123.880 37.230 124.140 ;
        RECT 41.600 124.080 41.740 124.220 ;
        RECT 38.380 123.940 41.740 124.080 ;
        RECT 42.405 124.080 42.695 124.125 ;
        RECT 43.595 124.080 43.885 124.125 ;
        RECT 46.115 124.080 46.405 124.125 ;
        RECT 42.405 123.940 46.405 124.080 ;
        RECT 36.005 123.555 36.295 123.785 ;
        RECT 37.385 123.740 37.675 123.785 ;
        RECT 37.830 123.740 38.150 123.800 ;
        RECT 38.380 123.785 38.520 123.940 ;
        RECT 42.405 123.895 42.695 123.940 ;
        RECT 43.595 123.895 43.885 123.940 ;
        RECT 46.115 123.895 46.405 123.940 ;
        RECT 49.330 123.880 49.650 124.140 ;
        RECT 65.905 124.080 66.195 124.125 ;
        RECT 66.365 124.080 66.655 124.125 ;
        RECT 65.905 123.940 66.655 124.080 ;
        RECT 65.905 123.895 66.195 123.940 ;
        RECT 66.365 123.895 66.655 123.940 ;
        RECT 37.385 123.600 38.150 123.740 ;
        RECT 37.385 123.555 37.675 123.600 ;
        RECT 36.080 123.400 36.220 123.555 ;
        RECT 37.830 123.540 38.150 123.600 ;
        RECT 38.305 123.555 38.595 123.785 ;
        RECT 39.210 123.540 39.530 123.800 ;
        RECT 39.670 123.540 39.990 123.800 ;
        RECT 41.065 123.555 41.355 123.785 ;
        RECT 41.525 123.740 41.815 123.785 ;
        RECT 44.730 123.740 45.050 123.800 ;
        RECT 41.525 123.600 45.050 123.740 ;
        RECT 41.525 123.555 41.815 123.600 ;
        RECT 40.590 123.400 40.910 123.460 ;
        RECT 36.080 123.260 40.910 123.400 ;
        RECT 40.590 123.200 40.910 123.260 ;
        RECT 31.405 123.060 31.695 123.105 ;
        RECT 31.850 123.060 32.170 123.120 ;
        RECT 31.405 122.920 32.170 123.060 ;
        RECT 41.140 123.060 41.280 123.555 ;
        RECT 44.730 123.540 45.050 123.600 ;
        RECT 48.870 123.540 49.190 123.800 ;
        RECT 59.910 123.540 60.230 123.800 ;
        RECT 67.730 123.540 68.050 123.800 ;
        RECT 68.190 123.540 68.510 123.800 ;
        RECT 68.665 123.555 68.955 123.785 ;
        RECT 69.110 123.740 69.430 123.800 ;
        RECT 69.585 123.740 69.875 123.785 ;
        RECT 69.110 123.600 69.875 123.740 ;
        RECT 42.860 123.400 43.150 123.445 ;
        RECT 43.810 123.400 44.130 123.460 ;
        RECT 42.860 123.260 44.130 123.400 ;
        RECT 42.860 123.215 43.150 123.260 ;
        RECT 43.810 123.200 44.130 123.260 ;
        RECT 53.025 123.215 53.315 123.445 ;
        RECT 65.890 123.400 66.210 123.460 ;
        RECT 68.740 123.400 68.880 123.555 ;
        RECT 69.110 123.540 69.430 123.600 ;
        RECT 69.585 123.555 69.875 123.600 ;
        RECT 65.890 123.260 68.880 123.400 ;
        RECT 46.570 123.060 46.890 123.120 ;
        RECT 41.140 122.920 46.890 123.060 ;
        RECT 31.405 122.875 31.695 122.920 ;
        RECT 31.850 122.860 32.170 122.920 ;
        RECT 46.570 122.860 46.890 122.920 ;
        RECT 50.725 123.060 51.015 123.105 ;
        RECT 51.170 123.060 51.490 123.120 ;
        RECT 53.100 123.060 53.240 123.215 ;
        RECT 65.890 123.200 66.210 123.260 ;
        RECT 50.725 122.920 53.240 123.060 ;
        RECT 56.690 123.060 57.010 123.120 ;
        RECT 57.165 123.060 57.455 123.105 ;
        RECT 56.690 122.920 57.455 123.060 ;
        RECT 50.725 122.875 51.015 122.920 ;
        RECT 51.170 122.860 51.490 122.920 ;
        RECT 56.690 122.860 57.010 122.920 ;
        RECT 57.165 122.875 57.455 122.920 ;
        RECT 61.750 123.060 62.070 123.120 ;
        RECT 62.685 123.060 62.975 123.105 ;
        RECT 61.750 122.920 62.975 123.060 ;
        RECT 61.750 122.860 62.070 122.920 ;
        RECT 62.685 122.875 62.975 122.920 ;
        RECT 13.380 122.240 92.040 122.720 ;
        RECT 100.010 122.450 100.880 125.790 ;
        RECT 108.930 125.490 116.850 125.500 ;
        RECT 105.160 125.480 116.850 125.490 ;
        RECT 101.540 125.360 116.850 125.480 ;
        RECT 101.540 125.350 116.875 125.360 ;
        RECT 101.500 125.230 116.875 125.350 ;
        RECT 101.500 125.120 105.500 125.230 ;
        RECT 101.110 124.780 101.340 125.070 ;
        RECT 101.560 124.780 105.450 125.120 ;
        RECT 105.660 124.780 105.890 125.070 ;
        RECT 101.110 123.410 105.890 124.780 ;
        RECT 101.110 123.110 101.340 123.410 ;
        RECT 105.660 123.110 105.890 123.410 ;
        RECT 101.500 122.830 105.500 123.060 ;
        RECT 101.750 122.600 105.320 122.830 ;
        RECT 101.750 122.450 105.440 122.600 ;
        RECT 100.010 122.170 105.440 122.450 ;
        RECT 106.690 122.280 107.310 125.230 ;
        RECT 108.875 125.130 116.875 125.230 ;
        RECT 108.930 125.120 116.850 125.130 ;
        RECT 108.440 124.420 108.670 125.080 ;
        RECT 109.450 124.420 110.450 124.510 ;
        RECT 117.080 124.420 117.310 125.080 ;
        RECT 108.440 123.600 117.310 124.420 ;
        RECT 108.440 123.120 108.670 123.600 ;
        RECT 109.450 123.510 110.450 123.600 ;
        RECT 117.080 123.120 117.310 123.600 ;
        RECT 108.875 122.840 116.875 123.070 ;
        RECT 30.025 122.040 30.315 122.085 ;
        RECT 30.930 122.040 31.250 122.100 ;
        RECT 30.025 121.900 31.250 122.040 ;
        RECT 30.025 121.855 30.315 121.900 ;
        RECT 30.930 121.840 31.250 121.900 ;
        RECT 46.570 122.040 46.890 122.100 ;
        RECT 47.965 122.040 48.255 122.085 ;
        RECT 46.570 121.900 48.255 122.040 ;
        RECT 46.570 121.840 46.890 121.900 ;
        RECT 47.965 121.855 48.255 121.900 ;
        RECT 48.870 122.040 49.190 122.100 ;
        RECT 63.145 122.040 63.435 122.085 ;
        RECT 48.870 121.900 63.435 122.040 ;
        RECT 48.870 121.840 49.190 121.900 ;
        RECT 63.145 121.855 63.435 121.900 ;
        RECT 46.125 121.700 46.415 121.745 ;
        RECT 58.070 121.700 58.390 121.760 ;
        RECT 46.125 121.560 48.640 121.700 ;
        RECT 46.125 121.515 46.415 121.560 ;
        RECT 48.500 121.420 48.640 121.560 ;
        RECT 55.400 121.560 58.390 121.700 ;
        RECT 23.110 121.160 23.430 121.420 ;
        RECT 23.570 121.360 23.890 121.420 ;
        RECT 24.405 121.360 24.695 121.405 ;
        RECT 23.570 121.220 24.695 121.360 ;
        RECT 23.570 121.160 23.890 121.220 ;
        RECT 24.405 121.175 24.695 121.220 ;
        RECT 47.045 121.175 47.335 121.405 ;
        RECT 48.410 121.360 48.730 121.420 ;
        RECT 48.885 121.360 49.175 121.405 ;
        RECT 48.410 121.220 49.175 121.360 ;
        RECT 24.005 121.020 24.295 121.065 ;
        RECT 25.195 121.020 25.485 121.065 ;
        RECT 27.715 121.020 28.005 121.065 ;
        RECT 24.005 120.880 28.005 121.020 ;
        RECT 47.120 121.020 47.260 121.175 ;
        RECT 48.410 121.160 48.730 121.220 ;
        RECT 48.885 121.175 49.175 121.220 ;
        RECT 49.790 121.160 50.110 121.420 ;
        RECT 55.400 121.405 55.540 121.560 ;
        RECT 58.070 121.500 58.390 121.560 ;
        RECT 100.010 121.710 105.450 122.170 ;
        RECT 56.690 121.405 57.010 121.420 ;
        RECT 55.325 121.175 55.615 121.405 ;
        RECT 56.660 121.360 57.010 121.405 ;
        RECT 62.685 121.360 62.975 121.405 ;
        RECT 56.495 121.220 57.010 121.360 ;
        RECT 56.660 121.175 57.010 121.220 ;
        RECT 56.690 121.160 57.010 121.175 ;
        RECT 62.300 121.220 62.975 121.360 ;
        RECT 49.880 121.020 50.020 121.160 ;
        RECT 47.120 120.880 50.020 121.020 ;
        RECT 56.205 121.020 56.495 121.065 ;
        RECT 57.395 121.020 57.685 121.065 ;
        RECT 59.915 121.020 60.205 121.065 ;
        RECT 56.205 120.880 60.205 121.020 ;
        RECT 24.005 120.835 24.295 120.880 ;
        RECT 25.195 120.835 25.485 120.880 ;
        RECT 27.715 120.835 28.005 120.880 ;
        RECT 56.205 120.835 56.495 120.880 ;
        RECT 57.395 120.835 57.685 120.880 ;
        RECT 59.915 120.835 60.205 120.880 ;
        RECT 23.610 120.680 23.900 120.725 ;
        RECT 25.710 120.680 26.000 120.725 ;
        RECT 27.280 120.680 27.570 120.725 ;
        RECT 23.610 120.540 27.570 120.680 ;
        RECT 23.610 120.495 23.900 120.540 ;
        RECT 25.710 120.495 26.000 120.540 ;
        RECT 27.280 120.495 27.570 120.540 ;
        RECT 41.050 120.680 41.370 120.740 ;
        RECT 62.300 120.725 62.440 121.220 ;
        RECT 62.685 121.175 62.975 121.220 ;
        RECT 63.605 121.360 63.895 121.405 ;
        RECT 67.270 121.360 67.590 121.420 ;
        RECT 63.605 121.220 67.590 121.360 ;
        RECT 63.605 121.175 63.895 121.220 ;
        RECT 67.270 121.160 67.590 121.220 ;
        RECT 72.905 121.360 73.195 121.405 ;
        RECT 73.710 121.360 74.030 121.420 ;
        RECT 72.905 121.220 74.030 121.360 ;
        RECT 72.905 121.175 73.195 121.220 ;
        RECT 73.710 121.160 74.030 121.220 ;
        RECT 74.170 121.360 74.490 121.420 ;
        RECT 76.930 121.360 77.250 121.420 ;
        RECT 74.170 121.220 77.250 121.360 ;
        RECT 74.170 121.160 74.490 121.220 ;
        RECT 76.930 121.160 77.250 121.220 ;
        RECT 69.595 121.020 69.885 121.065 ;
        RECT 72.115 121.020 72.405 121.065 ;
        RECT 73.305 121.020 73.595 121.065 ;
        RECT 69.595 120.880 73.595 121.020 ;
        RECT 69.595 120.835 69.885 120.880 ;
        RECT 72.115 120.835 72.405 120.880 ;
        RECT 73.305 120.835 73.595 120.880 ;
        RECT 49.805 120.680 50.095 120.725 ;
        RECT 41.050 120.540 50.095 120.680 ;
        RECT 41.050 120.480 41.370 120.540 ;
        RECT 49.805 120.495 50.095 120.540 ;
        RECT 55.810 120.680 56.100 120.725 ;
        RECT 57.910 120.680 58.200 120.725 ;
        RECT 59.480 120.680 59.770 120.725 ;
        RECT 55.810 120.540 59.770 120.680 ;
        RECT 55.810 120.495 56.100 120.540 ;
        RECT 57.910 120.495 58.200 120.540 ;
        RECT 59.480 120.495 59.770 120.540 ;
        RECT 62.225 120.495 62.515 120.725 ;
        RECT 70.030 120.680 70.320 120.725 ;
        RECT 71.600 120.680 71.890 120.725 ;
        RECT 73.700 120.680 73.990 120.725 ;
        RECT 70.030 120.540 73.990 120.680 ;
        RECT 70.030 120.495 70.320 120.540 ;
        RECT 71.600 120.495 71.890 120.540 ;
        RECT 73.700 120.495 73.990 120.540 ;
        RECT 45.190 120.140 45.510 120.400 ;
        RECT 67.285 120.340 67.575 120.385 ;
        RECT 68.650 120.340 68.970 120.400 ;
        RECT 67.285 120.200 68.970 120.340 ;
        RECT 67.285 120.155 67.575 120.200 ;
        RECT 68.650 120.140 68.970 120.200 ;
        RECT 100.010 120.360 102.050 121.710 ;
        RECT 103.800 121.700 105.450 121.710 ;
        RECT 102.490 120.430 103.490 121.150 ;
        RECT 103.800 120.890 104.110 121.700 ;
        RECT 104.570 121.420 105.450 121.700 ;
        RECT 105.690 121.880 107.310 122.280 ;
        RECT 108.960 121.930 116.830 122.840 ;
        RECT 104.510 121.190 105.510 121.420 ;
        RECT 105.690 121.230 106.040 121.880 ;
        RECT 106.690 121.870 107.310 121.880 ;
        RECT 108.875 121.700 116.875 121.930 ;
        RECT 108.960 121.690 116.830 121.700 ;
        RECT 104.570 120.980 105.450 121.000 ;
        RECT 103.840 120.600 104.110 120.890 ;
        RECT 104.510 120.750 105.510 120.980 ;
        RECT 105.670 120.940 106.040 121.230 ;
        RECT 105.700 120.880 106.040 120.940 ;
        RECT 106.800 121.550 107.560 121.600 ;
        RECT 108.440 121.550 108.670 121.650 ;
        RECT 106.800 121.340 108.670 121.550 ;
        RECT 117.080 121.340 117.310 121.650 ;
        RECT 106.800 120.920 109.340 121.340 ;
        RECT 116.710 120.920 117.310 121.340 ;
        RECT 104.570 120.600 105.450 120.750 ;
        RECT 104.580 120.430 105.310 120.600 ;
        RECT 13.380 119.520 92.040 120.000 ;
        RECT 23.570 119.120 23.890 119.380 ;
        RECT 24.490 119.320 24.810 119.380 ;
        RECT 31.390 119.320 31.710 119.380 ;
        RECT 24.490 119.180 31.710 119.320 ;
        RECT 24.490 119.120 24.810 119.180 ;
        RECT 31.390 119.120 31.710 119.180 ;
        RECT 67.270 119.120 67.590 119.380 ;
        RECT 67.730 119.120 68.050 119.380 ;
        RECT 73.710 119.320 74.030 119.380 ;
        RECT 74.185 119.320 74.475 119.365 ;
        RECT 73.710 119.180 74.475 119.320 ;
        RECT 73.710 119.120 74.030 119.180 ;
        RECT 74.185 119.135 74.475 119.180 ;
        RECT 18.970 118.980 19.260 119.025 ;
        RECT 20.540 118.980 20.830 119.025 ;
        RECT 22.640 118.980 22.930 119.025 ;
        RECT 27.290 118.980 27.580 119.025 ;
        RECT 29.390 118.980 29.680 119.025 ;
        RECT 30.960 118.980 31.250 119.025 ;
        RECT 18.970 118.840 22.930 118.980 ;
        RECT 18.970 118.795 19.260 118.840 ;
        RECT 20.540 118.795 20.830 118.840 ;
        RECT 22.640 118.795 22.930 118.840 ;
        RECT 23.200 118.840 27.020 118.980 ;
        RECT 23.200 118.700 23.340 118.840 ;
        RECT 18.535 118.640 18.825 118.685 ;
        RECT 21.055 118.640 21.345 118.685 ;
        RECT 22.245 118.640 22.535 118.685 ;
        RECT 18.535 118.500 22.535 118.640 ;
        RECT 18.535 118.455 18.825 118.500 ;
        RECT 21.055 118.455 21.345 118.500 ;
        RECT 22.245 118.455 22.535 118.500 ;
        RECT 23.110 118.440 23.430 118.700 ;
        RECT 26.880 118.685 27.020 118.840 ;
        RECT 27.290 118.840 31.250 118.980 ;
        RECT 27.290 118.795 27.580 118.840 ;
        RECT 29.390 118.795 29.680 118.840 ;
        RECT 30.960 118.795 31.250 118.840 ;
        RECT 53.050 118.980 53.340 119.025 ;
        RECT 55.150 118.980 55.440 119.025 ;
        RECT 56.720 118.980 57.010 119.025 ;
        RECT 53.050 118.840 57.010 118.980 ;
        RECT 53.050 118.795 53.340 118.840 ;
        RECT 55.150 118.795 55.440 118.840 ;
        RECT 56.720 118.795 57.010 118.840 ;
        RECT 60.870 118.980 61.160 119.025 ;
        RECT 62.970 118.980 63.260 119.025 ;
        RECT 64.540 118.980 64.830 119.025 ;
        RECT 60.870 118.840 64.830 118.980 ;
        RECT 60.870 118.795 61.160 118.840 ;
        RECT 62.970 118.795 63.260 118.840 ;
        RECT 64.540 118.795 64.830 118.840 ;
        RECT 26.805 118.455 27.095 118.685 ;
        RECT 27.685 118.640 27.975 118.685 ;
        RECT 28.875 118.640 29.165 118.685 ;
        RECT 31.395 118.640 31.685 118.685 ;
        RECT 27.685 118.500 31.685 118.640 ;
        RECT 27.685 118.455 27.975 118.500 ;
        RECT 28.875 118.455 29.165 118.500 ;
        RECT 31.395 118.455 31.685 118.500 ;
        RECT 53.445 118.640 53.735 118.685 ;
        RECT 54.635 118.640 54.925 118.685 ;
        RECT 57.155 118.640 57.445 118.685 ;
        RECT 53.445 118.500 57.445 118.640 ;
        RECT 53.445 118.455 53.735 118.500 ;
        RECT 54.635 118.455 54.925 118.500 ;
        RECT 57.155 118.455 57.445 118.500 ;
        RECT 61.265 118.640 61.555 118.685 ;
        RECT 62.455 118.640 62.745 118.685 ;
        RECT 64.975 118.640 65.265 118.685 ;
        RECT 61.265 118.500 65.265 118.640 ;
        RECT 67.360 118.640 67.500 119.120 ;
        RECT 70.505 118.640 70.795 118.685 ;
        RECT 67.360 118.500 70.795 118.640 ;
        RECT 61.265 118.455 61.555 118.500 ;
        RECT 62.455 118.455 62.745 118.500 ;
        RECT 64.975 118.455 65.265 118.500 ;
        RECT 70.505 118.455 70.795 118.500 ;
        RECT 24.490 118.100 24.810 118.360 ;
        RECT 24.950 118.300 25.270 118.360 ;
        RECT 25.425 118.300 25.715 118.345 ;
        RECT 24.950 118.160 25.715 118.300 ;
        RECT 24.950 118.100 25.270 118.160 ;
        RECT 25.425 118.115 25.715 118.160 ;
        RECT 25.885 118.115 26.175 118.345 ;
        RECT 36.925 118.300 37.215 118.345 ;
        RECT 33.780 118.160 37.215 118.300 ;
        RECT 21.900 117.960 22.190 118.005 ;
        RECT 24.030 117.960 24.350 118.020 ;
        RECT 21.900 117.820 24.350 117.960 ;
        RECT 21.900 117.775 22.190 117.820 ;
        RECT 24.030 117.760 24.350 117.820 ;
        RECT 16.225 117.620 16.515 117.665 ;
        RECT 18.050 117.620 18.370 117.680 ;
        RECT 16.225 117.480 18.370 117.620 ;
        RECT 16.225 117.435 16.515 117.480 ;
        RECT 18.050 117.420 18.370 117.480 ;
        RECT 24.490 117.620 24.810 117.680 ;
        RECT 25.960 117.620 26.100 118.115 ;
        RECT 26.330 117.960 26.650 118.020 ;
        RECT 28.030 117.960 28.320 118.005 ;
        RECT 26.330 117.820 28.320 117.960 ;
        RECT 26.330 117.760 26.650 117.820 ;
        RECT 28.030 117.775 28.320 117.820 ;
        RECT 24.490 117.480 26.100 117.620 ;
        RECT 30.930 117.620 31.250 117.680 ;
        RECT 33.780 117.665 33.920 118.160 ;
        RECT 36.925 118.115 37.215 118.160 ;
        RECT 41.050 118.100 41.370 118.360 ;
        RECT 50.250 118.300 50.570 118.360 ;
        RECT 52.565 118.300 52.855 118.345 ;
        RECT 58.070 118.300 58.390 118.360 ;
        RECT 61.750 118.345 62.070 118.360 ;
        RECT 60.385 118.300 60.675 118.345 ;
        RECT 61.720 118.300 62.070 118.345 ;
        RECT 50.250 118.160 60.675 118.300 ;
        RECT 61.555 118.160 62.070 118.300 ;
        RECT 50.250 118.100 50.570 118.160 ;
        RECT 52.565 118.115 52.855 118.160 ;
        RECT 58.070 118.100 58.390 118.160 ;
        RECT 60.385 118.115 60.675 118.160 ;
        RECT 61.720 118.115 62.070 118.160 ;
        RECT 61.750 118.100 62.070 118.115 ;
        RECT 68.650 118.300 68.970 118.360 ;
        RECT 71.425 118.300 71.715 118.345 ;
        RECT 71.870 118.300 72.190 118.360 ;
        RECT 68.650 118.160 72.190 118.300 ;
        RECT 68.650 118.100 68.970 118.160 ;
        RECT 71.425 118.115 71.715 118.160 ;
        RECT 71.870 118.100 72.190 118.160 ;
        RECT 73.250 118.100 73.570 118.360 ;
        RECT 53.930 118.005 54.250 118.020 ;
        RECT 53.900 117.775 54.250 118.005 ;
        RECT 53.930 117.760 54.250 117.775 ;
        RECT 66.350 117.960 66.670 118.020 ;
        RECT 72.345 117.960 72.635 118.005 ;
        RECT 66.350 117.820 72.635 117.960 ;
        RECT 66.350 117.760 66.670 117.820 ;
        RECT 72.345 117.775 72.635 117.820 ;
        RECT 72.790 117.760 73.110 118.020 ;
        RECT 33.705 117.620 33.995 117.665 ;
        RECT 30.930 117.480 33.995 117.620 ;
        RECT 24.490 117.420 24.810 117.480 ;
        RECT 30.930 117.420 31.250 117.480 ;
        RECT 33.705 117.435 33.995 117.480 ;
        RECT 34.150 117.420 34.470 117.680 ;
        RECT 37.830 117.620 38.150 117.680 ;
        RECT 38.305 117.620 38.595 117.665 ;
        RECT 37.830 117.480 38.595 117.620 ;
        RECT 37.830 117.420 38.150 117.480 ;
        RECT 38.305 117.435 38.595 117.480 ;
        RECT 57.150 117.620 57.470 117.680 ;
        RECT 59.465 117.620 59.755 117.665 ;
        RECT 57.150 117.480 59.755 117.620 ;
        RECT 57.150 117.420 57.470 117.480 ;
        RECT 59.465 117.435 59.755 117.480 ;
        RECT 13.380 116.800 92.040 117.280 ;
        RECT 100.010 116.810 100.780 120.360 ;
        RECT 102.460 119.310 105.310 120.430 ;
        RECT 105.700 120.130 106.050 120.880 ;
        RECT 106.800 120.760 108.670 120.920 ;
        RECT 106.800 120.710 107.560 120.760 ;
        RECT 108.440 120.690 108.670 120.760 ;
        RECT 117.080 120.690 117.310 120.920 ;
        RECT 108.875 120.410 116.875 120.640 ;
        RECT 105.700 120.070 105.990 120.130 ;
        RECT 105.610 119.950 105.990 120.070 ;
        RECT 108.970 120.010 116.830 120.410 ;
        RECT 117.640 120.010 118.600 129.490 ;
        RECT 119.930 129.680 120.770 131.810 ;
        RECT 126.430 131.390 127.680 131.830 ;
        RECT 137.600 131.810 138.460 133.870 ;
        RECT 124.370 131.380 129.610 131.390 ;
        RECT 121.420 131.280 136.720 131.380 ;
        RECT 121.420 131.270 136.755 131.280 ;
        RECT 121.380 131.150 136.755 131.270 ;
        RECT 121.380 131.040 125.380 131.150 ;
        RECT 126.430 131.070 128.170 131.150 ;
        RECT 128.750 131.070 136.755 131.150 ;
        RECT 126.430 130.990 127.680 131.070 ;
        RECT 128.755 131.050 136.755 131.070 ;
        RECT 120.990 130.740 121.220 130.990 ;
        RECT 125.540 130.850 125.770 130.990 ;
        RECT 128.320 130.850 128.550 131.000 ;
        RECT 125.540 130.740 128.550 130.850 ;
        RECT 136.960 130.740 137.190 131.000 ;
        RECT 120.990 130.300 137.190 130.740 ;
        RECT 120.990 130.030 121.220 130.300 ;
        RECT 125.540 130.270 137.190 130.300 ;
        RECT 125.540 130.180 128.550 130.270 ;
        RECT 125.540 130.030 125.770 130.180 ;
        RECT 128.320 130.040 128.550 130.180 ;
        RECT 136.960 130.040 137.190 130.270 ;
        RECT 121.380 129.750 125.380 129.980 ;
        RECT 128.755 129.770 136.755 129.990 ;
        RECT 137.520 129.770 138.480 131.810 ;
        RECT 128.755 129.760 138.480 129.770 ;
        RECT 121.380 129.680 125.370 129.750 ;
        RECT 119.930 129.570 125.370 129.680 ;
        RECT 128.810 129.600 138.480 129.760 ;
        RECT 119.930 129.480 123.060 129.570 ;
        RECT 136.550 129.550 138.480 129.600 ;
        RECT 119.930 126.210 120.770 129.480 ;
        RECT 124.410 129.020 129.660 129.030 ;
        RECT 124.410 128.910 136.720 129.020 ;
        RECT 121.440 128.850 136.720 128.910 ;
        RECT 121.440 128.840 136.755 128.850 ;
        RECT 121.380 128.710 136.755 128.840 ;
        RECT 121.380 128.700 126.540 128.710 ;
        RECT 121.380 128.610 125.380 128.700 ;
        RECT 128.755 128.620 136.755 128.710 ;
        RECT 128.840 128.610 136.730 128.620 ;
        RECT 120.990 128.250 121.220 128.560 ;
        RECT 121.440 128.250 125.340 128.610 ;
        RECT 125.540 128.250 125.770 128.560 ;
        RECT 120.990 126.910 125.770 128.250 ;
        RECT 120.990 126.600 121.220 126.910 ;
        RECT 125.540 126.600 125.770 126.910 ;
        RECT 128.320 128.030 128.550 128.570 ;
        RECT 129.360 128.030 130.370 128.060 ;
        RECT 136.960 128.030 137.190 128.570 ;
        RECT 128.320 127.130 137.190 128.030 ;
        RECT 128.320 126.610 128.550 127.130 ;
        RECT 129.360 127.060 130.370 127.130 ;
        RECT 136.960 126.610 137.190 127.130 ;
        RECT 121.380 126.320 125.380 126.550 ;
        RECT 128.755 126.330 136.755 126.560 ;
        RECT 119.930 126.170 121.060 126.210 ;
        RECT 119.930 126.090 121.300 126.170 ;
        RECT 121.670 126.100 125.330 126.320 ;
        RECT 121.670 126.090 123.110 126.100 ;
        RECT 119.930 126.050 123.110 126.090 ;
        RECT 119.930 125.960 122.620 126.050 ;
        RECT 128.820 126.040 136.710 126.330 ;
        RECT 119.930 125.900 121.950 125.960 ;
        RECT 119.930 125.850 121.700 125.900 ;
        RECT 119.930 122.510 120.770 125.850 ;
        RECT 128.810 125.550 136.730 125.560 ;
        RECT 125.040 125.540 136.730 125.550 ;
        RECT 121.420 125.420 136.730 125.540 ;
        RECT 121.420 125.410 136.755 125.420 ;
        RECT 121.380 125.290 136.755 125.410 ;
        RECT 121.380 125.180 125.380 125.290 ;
        RECT 120.990 124.840 121.220 125.130 ;
        RECT 121.440 124.840 125.330 125.180 ;
        RECT 125.540 124.840 125.770 125.130 ;
        RECT 120.990 123.470 125.770 124.840 ;
        RECT 120.990 123.170 121.220 123.470 ;
        RECT 125.540 123.170 125.770 123.470 ;
        RECT 121.380 122.890 125.380 123.120 ;
        RECT 121.630 122.660 125.200 122.890 ;
        RECT 121.630 122.510 125.320 122.660 ;
        RECT 119.930 122.230 125.320 122.510 ;
        RECT 126.570 122.340 127.190 125.290 ;
        RECT 128.755 125.190 136.755 125.290 ;
        RECT 128.810 125.180 136.730 125.190 ;
        RECT 128.320 124.480 128.550 125.140 ;
        RECT 129.330 124.480 130.330 124.570 ;
        RECT 136.960 124.480 137.190 125.140 ;
        RECT 128.320 123.660 137.190 124.480 ;
        RECT 128.320 123.180 128.550 123.660 ;
        RECT 129.330 123.570 130.330 123.660 ;
        RECT 136.960 123.180 137.190 123.660 ;
        RECT 128.755 122.900 136.755 123.130 ;
        RECT 119.930 121.770 125.330 122.230 ;
        RECT 119.930 120.430 121.930 121.770 ;
        RECT 123.680 121.760 125.330 121.770 ;
        RECT 122.370 120.490 123.370 121.210 ;
        RECT 123.680 120.950 123.990 121.760 ;
        RECT 124.450 121.480 125.330 121.760 ;
        RECT 125.570 121.940 127.190 122.340 ;
        RECT 128.840 121.990 136.710 122.900 ;
        RECT 124.390 121.250 125.390 121.480 ;
        RECT 125.570 121.290 125.920 121.940 ;
        RECT 126.570 121.930 127.190 121.940 ;
        RECT 128.755 121.760 136.755 121.990 ;
        RECT 128.840 121.750 136.710 121.760 ;
        RECT 124.450 121.040 125.330 121.060 ;
        RECT 123.720 120.660 123.990 120.950 ;
        RECT 124.390 120.810 125.390 121.040 ;
        RECT 125.550 121.000 125.920 121.290 ;
        RECT 125.580 120.940 125.920 121.000 ;
        RECT 126.680 121.610 127.440 121.660 ;
        RECT 128.320 121.610 128.550 121.710 ;
        RECT 126.680 121.400 128.550 121.610 ;
        RECT 136.960 121.400 137.190 121.710 ;
        RECT 126.680 120.980 129.220 121.400 ;
        RECT 136.590 120.980 137.190 121.400 ;
        RECT 124.450 120.660 125.330 120.810 ;
        RECT 124.460 120.490 125.190 120.660 ;
        RECT 102.400 119.080 105.400 119.310 ;
        RECT 105.610 119.120 105.950 119.950 ;
        RECT 107.960 119.940 118.600 120.010 ;
        RECT 102.450 119.050 105.310 119.080 ;
        RECT 102.450 119.030 103.620 119.050 ;
        RECT 104.580 119.040 105.310 119.050 ;
        RECT 102.400 118.640 105.400 118.870 ;
        RECT 105.605 118.830 105.950 119.120 ;
        RECT 106.140 118.900 118.600 119.940 ;
        RECT 120.000 120.420 121.930 120.430 ;
        RECT 106.140 118.880 118.560 118.900 ;
        RECT 105.610 118.720 105.950 118.830 ;
        RECT 106.180 118.870 111.850 118.880 ;
        RECT 112.850 118.870 118.560 118.880 ;
        RECT 102.490 118.470 105.350 118.640 ;
        RECT 106.180 118.470 106.610 118.870 ;
        RECT 102.460 118.100 106.610 118.470 ;
        RECT 100.000 116.780 100.780 116.810 ;
        RECT 25.885 116.415 26.175 116.645 ;
        RECT 39.210 116.600 39.530 116.660 ;
        RECT 40.145 116.600 40.435 116.645 ;
        RECT 39.210 116.460 40.435 116.600 ;
        RECT 24.030 116.260 24.350 116.320 ;
        RECT 25.960 116.260 26.100 116.415 ;
        RECT 39.210 116.400 39.530 116.460 ;
        RECT 40.145 116.415 40.435 116.460 ;
        RECT 57.165 116.600 57.455 116.645 ;
        RECT 59.910 116.600 60.230 116.660 ;
        RECT 57.165 116.460 60.230 116.600 ;
        RECT 57.165 116.415 57.455 116.460 ;
        RECT 59.910 116.400 60.230 116.460 ;
        RECT 66.350 116.400 66.670 116.660 ;
        RECT 68.190 116.600 68.510 116.660 ;
        RECT 69.125 116.600 69.415 116.645 ;
        RECT 68.190 116.460 69.415 116.600 ;
        RECT 68.190 116.400 68.510 116.460 ;
        RECT 69.125 116.415 69.415 116.460 ;
        RECT 24.030 116.120 26.100 116.260 ;
        RECT 26.725 116.260 27.015 116.305 ;
        RECT 27.250 116.260 27.570 116.320 ;
        RECT 26.725 116.120 27.570 116.260 ;
        RECT 24.030 116.060 24.350 116.120 ;
        RECT 26.725 116.075 27.015 116.120 ;
        RECT 27.250 116.060 27.570 116.120 ;
        RECT 27.725 116.260 28.015 116.305 ;
        RECT 34.150 116.260 34.470 116.320 ;
        RECT 39.300 116.260 39.440 116.400 ;
        RECT 27.725 116.120 34.470 116.260 ;
        RECT 27.725 116.075 28.015 116.120 ;
        RECT 34.150 116.060 34.470 116.120 ;
        RECT 37.460 116.120 39.440 116.260 ;
        RECT 12.070 115.920 12.390 115.980 ;
        RECT 15.305 115.920 15.595 115.965 ;
        RECT 12.070 115.780 15.595 115.920 ;
        RECT 12.070 115.720 12.390 115.780 ;
        RECT 15.305 115.735 15.595 115.780 ;
        RECT 24.950 115.720 25.270 115.980 ;
        RECT 25.425 115.920 25.715 115.965 ;
        RECT 28.185 115.920 28.475 115.965 ;
        RECT 25.425 115.780 28.475 115.920 ;
        RECT 25.425 115.735 25.715 115.780 ;
        RECT 28.185 115.735 28.475 115.780 ;
        RECT 31.850 115.720 32.170 115.980 ;
        RECT 37.460 115.965 37.600 116.120 ;
        RECT 32.785 115.735 33.075 115.965 ;
        RECT 37.385 115.735 37.675 115.965 ;
        RECT 25.040 115.580 25.180 115.720 ;
        RECT 27.250 115.580 27.570 115.640 ;
        RECT 25.040 115.440 27.570 115.580 ;
        RECT 27.250 115.380 27.570 115.440 ;
        RECT 31.405 115.580 31.695 115.625 ;
        RECT 32.325 115.580 32.615 115.625 ;
        RECT 31.405 115.440 32.615 115.580 ;
        RECT 31.405 115.395 31.695 115.440 ;
        RECT 32.325 115.395 32.615 115.440 ;
        RECT 16.225 115.240 16.515 115.285 ;
        RECT 16.670 115.240 16.990 115.300 ;
        RECT 16.225 115.100 16.990 115.240 ;
        RECT 16.225 115.055 16.515 115.100 ;
        RECT 16.670 115.040 16.990 115.100 ;
        RECT 24.045 115.240 24.335 115.285 ;
        RECT 26.330 115.240 26.650 115.300 ;
        RECT 24.045 115.100 26.650 115.240 ;
        RECT 24.045 115.055 24.335 115.100 ;
        RECT 26.330 115.040 26.650 115.100 ;
        RECT 30.930 115.240 31.250 115.300 ;
        RECT 32.860 115.240 33.000 115.735 ;
        RECT 36.910 115.380 37.230 115.640 ;
        RECT 30.930 115.100 33.000 115.240 ;
        RECT 30.930 115.040 31.250 115.100 ;
        RECT 37.460 114.960 37.600 115.735 ;
        RECT 37.830 115.720 38.150 115.980 ;
        RECT 40.145 115.735 40.435 115.965 ;
        RECT 40.590 115.920 40.910 115.980 ;
        RECT 41.065 115.920 41.355 115.965 ;
        RECT 41.970 115.920 42.290 115.980 ;
        RECT 40.590 115.780 42.290 115.920 ;
        RECT 38.305 115.395 38.595 115.625 ;
        RECT 40.220 115.580 40.360 115.735 ;
        RECT 40.590 115.720 40.910 115.780 ;
        RECT 41.065 115.735 41.355 115.780 ;
        RECT 41.970 115.720 42.290 115.780 ;
        RECT 44.270 115.920 44.590 115.980 ;
        RECT 45.190 115.920 45.510 115.980 ;
        RECT 44.270 115.780 45.510 115.920 ;
        RECT 44.270 115.720 44.590 115.780 ;
        RECT 45.190 115.720 45.510 115.780 ;
        RECT 46.125 115.735 46.415 115.965 ;
        RECT 41.510 115.580 41.830 115.640 ;
        RECT 40.220 115.440 41.830 115.580 ;
        RECT 38.380 115.240 38.520 115.395 ;
        RECT 41.510 115.380 41.830 115.440 ;
        RECT 42.890 115.240 43.210 115.300 ;
        RECT 38.380 115.100 43.210 115.240 ;
        RECT 42.890 115.040 43.210 115.100 ;
        RECT 45.190 115.240 45.510 115.300 ;
        RECT 46.200 115.240 46.340 115.735 ;
        RECT 50.250 115.720 50.570 115.980 ;
        RECT 51.630 115.965 51.950 115.980 ;
        RECT 51.600 115.735 51.950 115.965 ;
        RECT 51.630 115.720 51.950 115.735 ;
        RECT 65.890 115.720 66.210 115.980 ;
        RECT 66.825 115.920 67.115 115.965 ;
        RECT 68.280 115.920 68.420 116.400 ;
        RECT 66.825 115.780 68.420 115.920 ;
        RECT 66.825 115.735 67.115 115.780 ;
        RECT 49.790 115.380 50.110 115.640 ;
        RECT 51.145 115.580 51.435 115.625 ;
        RECT 52.335 115.580 52.625 115.625 ;
        RECT 54.855 115.580 55.145 115.625 ;
        RECT 51.145 115.440 55.145 115.580 ;
        RECT 51.145 115.395 51.435 115.440 ;
        RECT 52.335 115.395 52.625 115.440 ;
        RECT 54.855 115.395 55.145 115.440 ;
        RECT 46.585 115.240 46.875 115.285 ;
        RECT 45.190 115.100 46.875 115.240 ;
        RECT 45.190 115.040 45.510 115.100 ;
        RECT 46.585 115.055 46.875 115.100 ;
        RECT 50.750 115.240 51.040 115.285 ;
        RECT 52.850 115.240 53.140 115.285 ;
        RECT 54.420 115.240 54.710 115.285 ;
        RECT 50.750 115.100 54.710 115.240 ;
        RECT 68.280 115.240 68.420 115.780 ;
        RECT 68.650 115.720 68.970 115.980 ;
        RECT 69.585 115.920 69.875 115.965 ;
        RECT 70.030 115.920 70.350 115.980 ;
        RECT 69.585 115.780 70.350 115.920 ;
        RECT 69.585 115.735 69.875 115.780 ;
        RECT 70.030 115.720 70.350 115.780 ;
        RECT 88.430 115.920 88.750 115.980 ;
        RECT 88.905 115.920 89.195 115.965 ;
        RECT 88.430 115.780 89.195 115.920 ;
        RECT 88.430 115.720 88.750 115.780 ;
        RECT 88.905 115.735 89.195 115.780 ;
        RECT 71.870 115.580 72.190 115.640 ;
        RECT 72.345 115.580 72.635 115.625 ;
        RECT 71.870 115.440 72.635 115.580 ;
        RECT 71.870 115.380 72.190 115.440 ;
        RECT 72.345 115.395 72.635 115.440 ;
        RECT 73.725 115.240 74.015 115.285 ;
        RECT 68.280 115.100 74.015 115.240 ;
        RECT 50.750 115.055 51.040 115.100 ;
        RECT 52.850 115.055 53.140 115.100 ;
        RECT 54.420 115.055 54.710 115.100 ;
        RECT 73.725 115.055 74.015 115.100 ;
        RECT 89.810 115.040 90.130 115.300 ;
        RECT 26.805 114.900 27.095 114.945 ;
        RECT 31.850 114.900 32.170 114.960 ;
        RECT 26.805 114.760 32.170 114.900 ;
        RECT 26.805 114.715 27.095 114.760 ;
        RECT 31.850 114.700 32.170 114.760 ;
        RECT 35.990 114.700 36.310 114.960 ;
        RECT 37.370 114.700 37.690 114.960 ;
        RECT 43.810 114.900 44.130 114.960 ;
        RECT 44.745 114.900 45.035 114.945 ;
        RECT 43.810 114.760 45.035 114.900 ;
        RECT 43.810 114.700 44.130 114.760 ;
        RECT 44.745 114.715 45.035 114.760 ;
        RECT 45.650 114.700 45.970 114.960 ;
        RECT 74.645 114.900 74.935 114.945 ;
        RECT 79.230 114.900 79.550 114.960 ;
        RECT 74.645 114.760 79.550 114.900 ;
        RECT 74.645 114.715 74.935 114.760 ;
        RECT 79.230 114.700 79.550 114.760 ;
        RECT 100.000 114.680 100.830 116.780 ;
        RECT 106.500 116.390 107.750 116.830 ;
        RECT 117.700 116.810 118.560 118.870 ;
        RECT 120.000 116.810 120.770 120.420 ;
        RECT 122.340 119.370 125.190 120.490 ;
        RECT 125.580 120.190 125.930 120.940 ;
        RECT 126.680 120.820 128.550 120.980 ;
        RECT 126.680 120.770 127.440 120.820 ;
        RECT 128.320 120.750 128.550 120.820 ;
        RECT 136.960 120.750 137.190 120.980 ;
        RECT 128.755 120.470 136.755 120.700 ;
        RECT 125.580 120.130 125.870 120.190 ;
        RECT 125.490 120.010 125.870 120.130 ;
        RECT 128.850 120.070 136.710 120.470 ;
        RECT 137.520 120.070 138.480 129.550 ;
        RECT 122.280 119.140 125.280 119.370 ;
        RECT 125.490 119.180 125.830 120.010 ;
        RECT 127.840 120.000 138.480 120.070 ;
        RECT 122.330 119.110 125.190 119.140 ;
        RECT 122.330 119.090 123.500 119.110 ;
        RECT 124.460 119.100 125.190 119.110 ;
        RECT 122.280 118.700 125.280 118.930 ;
        RECT 125.485 118.890 125.830 119.180 ;
        RECT 126.020 118.960 138.480 120.000 ;
        RECT 139.930 131.780 140.700 135.360 ;
        RECT 142.370 134.310 145.220 135.430 ;
        RECT 145.610 135.130 145.960 135.880 ;
        RECT 146.710 135.760 148.580 135.920 ;
        RECT 146.710 135.710 147.470 135.760 ;
        RECT 148.350 135.690 148.580 135.760 ;
        RECT 156.990 135.690 157.220 135.920 ;
        RECT 148.785 135.410 156.785 135.640 ;
        RECT 145.610 135.070 145.900 135.130 ;
        RECT 145.520 134.950 145.900 135.070 ;
        RECT 148.880 135.010 156.740 135.410 ;
        RECT 157.550 135.010 158.510 144.490 ;
        RECT 142.310 134.080 145.310 134.310 ;
        RECT 145.520 134.120 145.860 134.950 ;
        RECT 147.870 134.940 158.510 135.010 ;
        RECT 142.360 134.050 145.220 134.080 ;
        RECT 142.360 134.030 143.530 134.050 ;
        RECT 144.490 134.040 145.220 134.050 ;
        RECT 142.310 133.640 145.310 133.870 ;
        RECT 145.515 133.830 145.860 134.120 ;
        RECT 146.050 133.900 158.510 134.940 ;
        RECT 146.050 133.880 158.500 133.900 ;
        RECT 145.520 133.720 145.860 133.830 ;
        RECT 146.090 133.870 151.760 133.880 ;
        RECT 152.760 133.870 158.500 133.880 ;
        RECT 142.400 133.470 145.260 133.640 ;
        RECT 146.090 133.470 146.520 133.870 ;
        RECT 142.370 133.100 146.520 133.470 ;
        RECT 139.930 129.680 140.790 131.780 ;
        RECT 146.460 131.390 147.710 131.830 ;
        RECT 157.640 131.810 158.500 133.870 ;
        RECT 144.400 131.380 149.640 131.390 ;
        RECT 141.450 131.280 156.750 131.380 ;
        RECT 141.450 131.270 156.785 131.280 ;
        RECT 141.410 131.150 156.785 131.270 ;
        RECT 141.410 131.040 145.410 131.150 ;
        RECT 146.460 131.070 148.200 131.150 ;
        RECT 148.780 131.070 156.785 131.150 ;
        RECT 146.460 130.990 147.710 131.070 ;
        RECT 148.785 131.050 156.785 131.070 ;
        RECT 141.020 130.740 141.250 130.990 ;
        RECT 145.570 130.850 145.800 130.990 ;
        RECT 148.350 130.850 148.580 131.000 ;
        RECT 145.570 130.740 148.580 130.850 ;
        RECT 156.990 130.740 157.220 131.000 ;
        RECT 141.020 130.300 157.220 130.740 ;
        RECT 141.020 130.030 141.250 130.300 ;
        RECT 145.570 130.270 157.220 130.300 ;
        RECT 145.570 130.180 148.580 130.270 ;
        RECT 145.570 130.030 145.800 130.180 ;
        RECT 148.350 130.040 148.580 130.180 ;
        RECT 156.990 130.040 157.220 130.270 ;
        RECT 141.410 129.750 145.410 129.980 ;
        RECT 148.785 129.770 156.785 129.990 ;
        RECT 157.550 129.770 158.510 131.810 ;
        RECT 148.785 129.760 158.510 129.770 ;
        RECT 141.410 129.680 145.400 129.750 ;
        RECT 139.930 129.570 145.400 129.680 ;
        RECT 148.840 129.600 158.510 129.760 ;
        RECT 139.930 129.480 143.090 129.570 ;
        RECT 156.580 129.550 158.510 129.600 ;
        RECT 139.930 126.210 140.790 129.480 ;
        RECT 144.440 129.020 149.690 129.030 ;
        RECT 144.440 128.910 156.750 129.020 ;
        RECT 141.470 128.850 156.750 128.910 ;
        RECT 141.470 128.840 156.785 128.850 ;
        RECT 141.410 128.710 156.785 128.840 ;
        RECT 141.410 128.700 146.570 128.710 ;
        RECT 141.410 128.610 145.410 128.700 ;
        RECT 148.785 128.620 156.785 128.710 ;
        RECT 148.870 128.610 156.760 128.620 ;
        RECT 141.020 128.250 141.250 128.560 ;
        RECT 141.470 128.250 145.370 128.610 ;
        RECT 145.570 128.250 145.800 128.560 ;
        RECT 141.020 126.910 145.800 128.250 ;
        RECT 141.020 126.600 141.250 126.910 ;
        RECT 145.570 126.600 145.800 126.910 ;
        RECT 148.350 128.030 148.580 128.570 ;
        RECT 149.390 128.030 150.400 128.060 ;
        RECT 156.990 128.030 157.220 128.570 ;
        RECT 148.350 127.130 157.220 128.030 ;
        RECT 148.350 126.610 148.580 127.130 ;
        RECT 149.390 127.060 150.400 127.130 ;
        RECT 156.990 126.610 157.220 127.130 ;
        RECT 141.410 126.320 145.410 126.550 ;
        RECT 148.785 126.330 156.785 126.560 ;
        RECT 139.930 126.170 141.090 126.210 ;
        RECT 139.930 126.090 141.330 126.170 ;
        RECT 141.700 126.100 145.360 126.320 ;
        RECT 141.700 126.090 143.140 126.100 ;
        RECT 139.930 126.050 143.140 126.090 ;
        RECT 139.930 125.960 142.650 126.050 ;
        RECT 148.850 126.040 156.740 126.330 ;
        RECT 139.930 125.900 141.980 125.960 ;
        RECT 139.930 125.850 141.730 125.900 ;
        RECT 139.930 122.510 140.790 125.850 ;
        RECT 148.840 125.550 156.760 125.560 ;
        RECT 145.070 125.540 156.760 125.550 ;
        RECT 141.450 125.420 156.760 125.540 ;
        RECT 141.450 125.410 156.785 125.420 ;
        RECT 141.410 125.290 156.785 125.410 ;
        RECT 141.410 125.180 145.410 125.290 ;
        RECT 141.020 124.840 141.250 125.130 ;
        RECT 141.470 124.840 145.360 125.180 ;
        RECT 145.570 124.840 145.800 125.130 ;
        RECT 141.020 123.470 145.800 124.840 ;
        RECT 141.020 123.170 141.250 123.470 ;
        RECT 145.570 123.170 145.800 123.470 ;
        RECT 141.410 122.890 145.410 123.120 ;
        RECT 141.660 122.660 145.230 122.890 ;
        RECT 141.660 122.510 145.350 122.660 ;
        RECT 139.930 122.230 145.350 122.510 ;
        RECT 146.600 122.340 147.220 125.290 ;
        RECT 148.785 125.190 156.785 125.290 ;
        RECT 148.840 125.180 156.760 125.190 ;
        RECT 148.350 124.480 148.580 125.140 ;
        RECT 149.360 124.480 150.360 124.570 ;
        RECT 156.990 124.480 157.220 125.140 ;
        RECT 148.350 123.660 157.220 124.480 ;
        RECT 148.350 123.180 148.580 123.660 ;
        RECT 149.360 123.570 150.360 123.660 ;
        RECT 156.990 123.180 157.220 123.660 ;
        RECT 148.785 122.900 156.785 123.130 ;
        RECT 139.930 121.770 145.360 122.230 ;
        RECT 139.930 120.420 141.960 121.770 ;
        RECT 143.710 121.760 145.360 121.770 ;
        RECT 142.400 120.490 143.400 121.210 ;
        RECT 143.710 120.950 144.020 121.760 ;
        RECT 144.480 121.480 145.360 121.760 ;
        RECT 145.600 121.940 147.220 122.340 ;
        RECT 148.870 121.990 156.740 122.900 ;
        RECT 144.420 121.250 145.420 121.480 ;
        RECT 145.600 121.290 145.950 121.940 ;
        RECT 146.600 121.930 147.220 121.940 ;
        RECT 148.785 121.760 156.785 121.990 ;
        RECT 148.870 121.750 156.740 121.760 ;
        RECT 144.480 121.040 145.360 121.060 ;
        RECT 143.750 120.660 144.020 120.950 ;
        RECT 144.420 120.810 145.420 121.040 ;
        RECT 145.580 121.000 145.950 121.290 ;
        RECT 145.610 120.940 145.950 121.000 ;
        RECT 146.710 121.610 147.470 121.660 ;
        RECT 148.350 121.610 148.580 121.710 ;
        RECT 146.710 121.400 148.580 121.610 ;
        RECT 156.990 121.400 157.220 121.710 ;
        RECT 146.710 120.980 149.250 121.400 ;
        RECT 156.620 120.980 157.220 121.400 ;
        RECT 144.480 120.660 145.360 120.810 ;
        RECT 144.490 120.490 145.220 120.660 ;
        RECT 126.020 118.940 138.460 118.960 ;
        RECT 125.490 118.780 125.830 118.890 ;
        RECT 126.060 118.930 131.730 118.940 ;
        RECT 132.730 118.930 138.460 118.940 ;
        RECT 122.370 118.530 125.230 118.700 ;
        RECT 126.060 118.530 126.490 118.930 ;
        RECT 122.340 118.160 126.490 118.530 ;
        RECT 104.440 116.380 109.680 116.390 ;
        RECT 101.490 116.280 116.790 116.380 ;
        RECT 101.490 116.270 116.825 116.280 ;
        RECT 101.450 116.150 116.825 116.270 ;
        RECT 101.450 116.040 105.450 116.150 ;
        RECT 106.500 116.070 108.240 116.150 ;
        RECT 108.820 116.070 116.825 116.150 ;
        RECT 106.500 115.990 107.750 116.070 ;
        RECT 108.825 116.050 116.825 116.070 ;
        RECT 101.060 115.740 101.290 115.990 ;
        RECT 105.610 115.850 105.840 115.990 ;
        RECT 108.390 115.850 108.620 116.000 ;
        RECT 105.610 115.740 108.620 115.850 ;
        RECT 117.030 115.740 117.260 116.000 ;
        RECT 101.060 115.300 117.260 115.740 ;
        RECT 101.060 115.030 101.290 115.300 ;
        RECT 105.610 115.270 117.260 115.300 ;
        RECT 105.610 115.180 108.620 115.270 ;
        RECT 105.610 115.030 105.840 115.180 ;
        RECT 108.390 115.040 108.620 115.180 ;
        RECT 117.030 115.040 117.260 115.270 ;
        RECT 101.450 114.750 105.450 114.980 ;
        RECT 108.825 114.770 116.825 114.990 ;
        RECT 117.590 114.770 118.560 116.810 ;
        RECT 108.825 114.760 118.560 114.770 ;
        RECT 101.450 114.680 105.440 114.750 ;
        RECT 100.000 114.570 105.440 114.680 ;
        RECT 108.880 114.600 118.560 114.760 ;
        RECT 13.380 114.080 92.040 114.560 ;
        RECT 100.000 114.480 103.130 114.570 ;
        RECT 116.620 114.550 118.560 114.600 ;
        RECT 57.165 113.880 57.455 113.925 ;
        RECT 57.610 113.880 57.930 113.940 ;
        RECT 57.165 113.740 57.930 113.880 ;
        RECT 57.165 113.695 57.455 113.740 ;
        RECT 57.610 113.680 57.930 113.740 ;
        RECT 88.430 113.680 88.750 113.940 ;
        RECT 35.110 113.540 35.400 113.585 ;
        RECT 37.210 113.540 37.500 113.585 ;
        RECT 38.780 113.540 39.070 113.585 ;
        RECT 35.110 113.400 39.070 113.540 ;
        RECT 35.110 113.355 35.400 113.400 ;
        RECT 37.210 113.355 37.500 113.400 ;
        RECT 38.780 113.355 39.070 113.400 ;
        RECT 45.230 113.540 45.520 113.585 ;
        RECT 47.330 113.540 47.620 113.585 ;
        RECT 48.900 113.540 49.190 113.585 ;
        RECT 45.230 113.400 49.190 113.540 ;
        RECT 45.230 113.355 45.520 113.400 ;
        RECT 47.330 113.355 47.620 113.400 ;
        RECT 48.900 113.355 49.190 113.400 ;
        RECT 49.790 113.540 50.110 113.600 ;
        RECT 51.645 113.540 51.935 113.585 ;
        RECT 49.790 113.400 51.935 113.540 ;
        RECT 49.790 113.340 50.110 113.400 ;
        RECT 51.645 113.355 51.935 113.400 ;
        RECT 59.030 113.540 59.320 113.585 ;
        RECT 61.130 113.540 61.420 113.585 ;
        RECT 62.700 113.540 62.990 113.585 ;
        RECT 59.030 113.400 62.990 113.540 ;
        RECT 59.030 113.355 59.320 113.400 ;
        RECT 61.130 113.355 61.420 113.400 ;
        RECT 62.700 113.355 62.990 113.400 ;
        RECT 70.030 113.340 70.350 113.600 ;
        RECT 72.790 113.540 73.080 113.585 ;
        RECT 74.360 113.540 74.650 113.585 ;
        RECT 76.460 113.540 76.750 113.585 ;
        RECT 72.790 113.400 76.750 113.540 ;
        RECT 72.790 113.355 73.080 113.400 ;
        RECT 74.360 113.355 74.650 113.400 ;
        RECT 76.460 113.355 76.750 113.400 ;
        RECT 35.505 113.200 35.795 113.245 ;
        RECT 36.695 113.200 36.985 113.245 ;
        RECT 39.215 113.200 39.505 113.245 ;
        RECT 35.505 113.060 39.505 113.200 ;
        RECT 35.505 113.015 35.795 113.060 ;
        RECT 36.695 113.015 36.985 113.060 ;
        RECT 39.215 113.015 39.505 113.060 ;
        RECT 44.730 113.000 45.050 113.260 ;
        RECT 45.625 113.200 45.915 113.245 ;
        RECT 46.815 113.200 47.105 113.245 ;
        RECT 49.335 113.200 49.625 113.245 ;
        RECT 45.625 113.060 49.625 113.200 ;
        RECT 45.625 113.015 45.915 113.060 ;
        RECT 46.815 113.015 47.105 113.060 ;
        RECT 49.335 113.015 49.625 113.060 ;
        RECT 12.070 112.860 12.390 112.920 ;
        RECT 14.845 112.860 15.135 112.905 ;
        RECT 12.070 112.720 15.135 112.860 ;
        RECT 12.070 112.660 12.390 112.720 ;
        RECT 14.845 112.675 15.135 112.720 ;
        RECT 16.225 112.860 16.515 112.905 ;
        RECT 17.130 112.860 17.450 112.920 ;
        RECT 21.730 112.860 22.050 112.920 ;
        RECT 22.205 112.860 22.495 112.905 ;
        RECT 16.225 112.720 20.580 112.860 ;
        RECT 16.225 112.675 16.515 112.720 ;
        RECT 17.130 112.660 17.450 112.720 ;
        RECT 8.390 112.520 8.710 112.580 ;
        RECT 20.440 112.520 20.580 112.720 ;
        RECT 21.730 112.720 22.495 112.860 ;
        RECT 21.730 112.660 22.050 112.720 ;
        RECT 22.205 112.675 22.495 112.720 ;
        RECT 23.110 112.860 23.430 112.920 ;
        RECT 31.390 112.860 31.710 112.920 ;
        RECT 34.625 112.860 34.915 112.905 ;
        RECT 23.110 112.720 34.915 112.860 ;
        RECT 23.110 112.660 23.430 112.720 ;
        RECT 31.390 112.660 31.710 112.720 ;
        RECT 34.625 112.675 34.915 112.720 ;
        RECT 35.620 112.720 42.660 112.860 ;
        RECT 26.790 112.520 27.110 112.580 ;
        RECT 35.620 112.520 35.760 112.720 ;
        RECT 8.390 112.380 20.120 112.520 ;
        RECT 20.440 112.380 35.760 112.520 ;
        RECT 35.960 112.520 36.250 112.565 ;
        RECT 41.985 112.520 42.275 112.565 ;
        RECT 35.960 112.380 42.275 112.520 ;
        RECT 8.390 112.320 8.710 112.380 ;
        RECT 19.430 111.980 19.750 112.240 ;
        RECT 19.980 112.180 20.120 112.380 ;
        RECT 26.790 112.320 27.110 112.380 ;
        RECT 35.960 112.335 36.250 112.380 ;
        RECT 41.985 112.335 42.275 112.380 ;
        RECT 36.910 112.180 37.230 112.240 ;
        RECT 19.980 112.040 37.230 112.180 ;
        RECT 36.910 111.980 37.230 112.040 ;
        RECT 40.590 112.180 40.910 112.240 ;
        RECT 41.510 112.180 41.830 112.240 ;
        RECT 40.590 112.040 41.830 112.180 ;
        RECT 42.520 112.180 42.660 112.720 ;
        RECT 42.890 112.660 43.210 112.920 ;
        RECT 43.810 112.660 44.130 112.920 ;
        RECT 44.270 112.860 44.590 112.920 ;
        RECT 49.880 112.860 50.020 113.340 ;
        RECT 58.070 113.200 58.390 113.260 ;
        RECT 58.545 113.200 58.835 113.245 ;
        RECT 58.070 113.060 58.835 113.200 ;
        RECT 58.070 113.000 58.390 113.060 ;
        RECT 58.545 113.015 58.835 113.060 ;
        RECT 59.425 113.200 59.715 113.245 ;
        RECT 60.615 113.200 60.905 113.245 ;
        RECT 63.135 113.200 63.425 113.245 ;
        RECT 59.425 113.060 63.425 113.200 ;
        RECT 59.425 113.015 59.715 113.060 ;
        RECT 60.615 113.015 60.905 113.060 ;
        RECT 63.135 113.015 63.425 113.060 ;
        RECT 72.355 113.200 72.645 113.245 ;
        RECT 74.875 113.200 75.165 113.245 ;
        RECT 76.065 113.200 76.355 113.245 ;
        RECT 72.355 113.060 76.355 113.200 ;
        RECT 72.355 113.015 72.645 113.060 ;
        RECT 74.875 113.015 75.165 113.060 ;
        RECT 76.065 113.015 76.355 113.060 ;
        RECT 44.270 112.720 44.770 112.860 ;
        RECT 45.740 112.720 50.020 112.860 ;
        RECT 44.270 112.660 44.590 112.720 ;
        RECT 44.730 112.520 45.050 112.580 ;
        RECT 45.740 112.520 45.880 112.720 ;
        RECT 55.325 112.675 55.615 112.905 ;
        RECT 64.510 112.860 64.830 112.920 ;
        RECT 65.905 112.860 66.195 112.905 ;
        RECT 64.510 112.720 66.195 112.860 ;
        RECT 46.110 112.565 46.430 112.580 ;
        RECT 44.730 112.380 45.880 112.520 ;
        RECT 44.730 112.320 45.050 112.380 ;
        RECT 46.080 112.335 46.430 112.565 ;
        RECT 46.110 112.320 46.430 112.335 ;
        RECT 55.400 112.180 55.540 112.675 ;
        RECT 64.510 112.660 64.830 112.720 ;
        RECT 65.905 112.675 66.195 112.720 ;
        RECT 66.825 112.675 67.115 112.905 ;
        RECT 69.585 112.860 69.875 112.905 ;
        RECT 70.490 112.860 70.810 112.920 ;
        RECT 72.790 112.860 73.110 112.920 ;
        RECT 69.585 112.720 73.110 112.860 ;
        RECT 69.585 112.675 69.875 112.720 ;
        RECT 57.150 112.320 57.470 112.580 ;
        RECT 59.880 112.520 60.170 112.565 ;
        RECT 66.365 112.520 66.655 112.565 ;
        RECT 59.880 112.380 66.655 112.520 ;
        RECT 66.900 112.520 67.040 112.675 ;
        RECT 70.490 112.660 70.810 112.720 ;
        RECT 72.790 112.660 73.110 112.720 ;
        RECT 76.930 112.860 77.250 112.920 ;
        RECT 79.690 112.860 80.010 112.920 ;
        RECT 76.930 112.720 80.010 112.860 ;
        RECT 76.930 112.660 77.250 112.720 ;
        RECT 79.690 112.660 80.010 112.720 ;
        RECT 87.510 112.660 87.830 112.920 ;
        RECT 88.430 112.860 88.750 112.920 ;
        RECT 88.905 112.860 89.195 112.905 ;
        RECT 88.430 112.720 89.195 112.860 ;
        RECT 88.430 112.660 88.750 112.720 ;
        RECT 88.905 112.675 89.195 112.720 ;
        RECT 70.950 112.520 71.270 112.580 ;
        RECT 66.900 112.380 71.270 112.520 ;
        RECT 59.880 112.335 60.170 112.380 ;
        RECT 66.365 112.335 66.655 112.380 ;
        RECT 70.950 112.320 71.270 112.380 ;
        RECT 74.630 112.520 74.950 112.580 ;
        RECT 75.610 112.520 75.900 112.565 ;
        RECT 74.630 112.380 75.900 112.520 ;
        RECT 74.630 112.320 74.950 112.380 ;
        RECT 75.610 112.335 75.900 112.380 ;
        RECT 56.230 112.180 56.550 112.240 ;
        RECT 42.520 112.040 56.550 112.180 ;
        RECT 40.590 111.980 40.910 112.040 ;
        RECT 41.510 111.980 41.830 112.040 ;
        RECT 56.230 111.980 56.550 112.040 ;
        RECT 58.085 112.180 58.375 112.225 ;
        RECT 64.970 112.180 65.290 112.240 ;
        RECT 58.085 112.040 65.290 112.180 ;
        RECT 58.085 111.995 58.375 112.040 ;
        RECT 64.970 111.980 65.290 112.040 ;
        RECT 65.445 112.180 65.735 112.225 ;
        RECT 66.810 112.180 67.130 112.240 ;
        RECT 68.650 112.180 68.970 112.240 ;
        RECT 65.445 112.040 68.970 112.180 ;
        RECT 65.445 111.995 65.735 112.040 ;
        RECT 66.810 111.980 67.130 112.040 ;
        RECT 68.650 111.980 68.970 112.040 ;
        RECT 69.110 112.180 69.430 112.240 ;
        RECT 74.170 112.180 74.490 112.240 ;
        RECT 69.110 112.040 74.490 112.180 ;
        RECT 69.110 111.980 69.430 112.040 ;
        RECT 74.170 111.980 74.490 112.040 ;
        RECT 89.810 111.980 90.130 112.240 ;
        RECT 13.380 111.360 92.040 111.840 ;
        RECT 21.285 111.160 21.575 111.205 ;
        RECT 22.190 111.160 22.510 111.220 ;
        RECT 21.285 111.020 22.510 111.160 ;
        RECT 21.285 110.975 21.575 111.020 ;
        RECT 22.190 110.960 22.510 111.020 ;
        RECT 23.110 110.960 23.430 111.220 ;
        RECT 38.305 111.160 38.595 111.205 ;
        RECT 42.890 111.160 43.210 111.220 ;
        RECT 38.305 111.020 40.820 111.160 ;
        RECT 38.305 110.975 38.595 111.020 ;
        RECT 23.200 110.820 23.340 110.960 ;
        RECT 21.820 110.680 23.340 110.820 ;
        RECT 32.740 110.820 33.030 110.865 ;
        RECT 35.990 110.820 36.310 110.880 ;
        RECT 32.740 110.680 36.310 110.820 ;
        RECT 21.820 110.540 21.960 110.680 ;
        RECT 32.740 110.635 33.030 110.680 ;
        RECT 35.990 110.620 36.310 110.680 ;
        RECT 16.225 110.480 16.515 110.525 ;
        RECT 16.670 110.480 16.990 110.540 ;
        RECT 16.225 110.340 16.990 110.480 ;
        RECT 16.225 110.295 16.515 110.340 ;
        RECT 16.670 110.280 16.990 110.340 ;
        RECT 18.050 110.280 18.370 110.540 ;
        RECT 21.730 110.280 22.050 110.540 ;
        RECT 23.110 110.525 23.430 110.540 ;
        RECT 23.080 110.295 23.430 110.525 ;
        RECT 23.110 110.280 23.430 110.295 ;
        RECT 27.250 110.480 27.570 110.540 ;
        RECT 29.105 110.480 29.395 110.525 ;
        RECT 27.250 110.340 29.395 110.480 ;
        RECT 27.250 110.280 27.570 110.340 ;
        RECT 29.105 110.295 29.395 110.340 ;
        RECT 30.025 110.480 30.315 110.525 ;
        RECT 30.930 110.480 31.250 110.540 ;
        RECT 30.025 110.340 31.250 110.480 ;
        RECT 30.025 110.295 30.315 110.340 ;
        RECT 30.930 110.280 31.250 110.340 ;
        RECT 31.390 110.280 31.710 110.540 ;
        RECT 36.450 110.480 36.770 110.540 ;
        RECT 40.680 110.525 40.820 111.020 ;
        RECT 42.890 111.020 44.040 111.160 ;
        RECT 42.890 110.960 43.210 111.020 ;
        RECT 41.510 110.820 41.830 110.880 ;
        RECT 43.365 110.820 43.655 110.865 ;
        RECT 41.510 110.680 43.655 110.820 ;
        RECT 43.900 110.820 44.040 111.020 ;
        RECT 46.110 110.960 46.430 111.220 ;
        RECT 64.510 110.960 64.830 111.220 ;
        RECT 64.970 111.160 65.290 111.220 ;
        RECT 67.285 111.160 67.575 111.205 ;
        RECT 64.970 111.020 67.575 111.160 ;
        RECT 64.970 110.960 65.290 111.020 ;
        RECT 67.285 110.975 67.575 111.020 ;
        RECT 68.665 110.975 68.955 111.205 ;
        RECT 70.045 111.160 70.335 111.205 ;
        RECT 70.490 111.160 70.810 111.220 ;
        RECT 70.045 111.020 70.810 111.160 ;
        RECT 70.045 110.975 70.335 111.020 ;
        RECT 47.045 110.820 47.335 110.865 ;
        RECT 43.900 110.680 47.335 110.820 ;
        RECT 41.510 110.620 41.830 110.680 ;
        RECT 43.365 110.635 43.655 110.680 ;
        RECT 47.045 110.635 47.335 110.680 ;
        RECT 39.685 110.480 39.975 110.525 ;
        RECT 36.450 110.340 39.975 110.480 ;
        RECT 36.450 110.280 36.770 110.340 ;
        RECT 39.685 110.295 39.975 110.340 ;
        RECT 40.605 110.480 40.895 110.525 ;
        RECT 41.050 110.480 41.370 110.540 ;
        RECT 40.605 110.340 41.370 110.480 ;
        RECT 40.605 110.295 40.895 110.340 ;
        RECT 41.050 110.280 41.370 110.340 ;
        RECT 42.430 110.480 42.750 110.540 ;
        RECT 44.270 110.480 44.590 110.540 ;
        RECT 42.430 110.340 44.590 110.480 ;
        RECT 42.430 110.280 42.750 110.340 ;
        RECT 44.270 110.280 44.590 110.340 ;
        RECT 44.745 110.480 45.035 110.525 ;
        RECT 45.190 110.480 45.510 110.540 ;
        RECT 44.745 110.340 45.510 110.480 ;
        RECT 44.745 110.295 45.035 110.340 ;
        RECT 45.190 110.280 45.510 110.340 ;
        RECT 46.585 110.295 46.875 110.525 ;
        RECT 17.590 109.940 17.910 110.200 ;
        RECT 22.625 110.140 22.915 110.185 ;
        RECT 23.815 110.140 24.105 110.185 ;
        RECT 26.335 110.140 26.625 110.185 ;
        RECT 22.625 110.000 26.625 110.140 ;
        RECT 22.625 109.955 22.915 110.000 ;
        RECT 23.815 109.955 24.105 110.000 ;
        RECT 26.335 109.955 26.625 110.000 ;
        RECT 32.285 110.140 32.575 110.185 ;
        RECT 33.475 110.140 33.765 110.185 ;
        RECT 35.995 110.140 36.285 110.185 ;
        RECT 32.285 110.000 36.285 110.140 ;
        RECT 32.285 109.955 32.575 110.000 ;
        RECT 33.475 109.955 33.765 110.000 ;
        RECT 35.995 109.955 36.285 110.000 ;
        RECT 45.650 110.140 45.970 110.200 ;
        RECT 46.125 110.140 46.415 110.185 ;
        RECT 45.650 110.000 46.415 110.140 ;
        RECT 45.650 109.940 45.970 110.000 ;
        RECT 46.125 109.955 46.415 110.000 ;
        RECT 16.685 109.800 16.975 109.845 ;
        RECT 22.230 109.800 22.520 109.845 ;
        RECT 24.330 109.800 24.620 109.845 ;
        RECT 25.900 109.800 26.190 109.845 ;
        RECT 16.685 109.660 21.730 109.800 ;
        RECT 16.685 109.615 16.975 109.660 ;
        RECT 17.145 109.460 17.435 109.505 ;
        RECT 18.510 109.460 18.830 109.520 ;
        RECT 17.145 109.320 18.830 109.460 ;
        RECT 21.590 109.460 21.730 109.660 ;
        RECT 22.230 109.660 26.190 109.800 ;
        RECT 22.230 109.615 22.520 109.660 ;
        RECT 24.330 109.615 24.620 109.660 ;
        RECT 25.900 109.615 26.190 109.660 ;
        RECT 31.890 109.800 32.180 109.845 ;
        RECT 33.990 109.800 34.280 109.845 ;
        RECT 35.560 109.800 35.850 109.845 ;
        RECT 31.890 109.660 35.850 109.800 ;
        RECT 31.890 109.615 32.180 109.660 ;
        RECT 33.990 109.615 34.280 109.660 ;
        RECT 35.560 109.615 35.850 109.660 ;
        RECT 41.525 109.800 41.815 109.845 ;
        RECT 46.660 109.800 46.800 110.295 ;
        RECT 56.230 110.280 56.550 110.540 ;
        RECT 57.150 110.280 57.470 110.540 ;
        RECT 57.610 110.280 57.930 110.540 ;
        RECT 63.590 110.280 63.910 110.540 ;
        RECT 67.360 110.480 67.500 110.975 ;
        RECT 68.740 110.820 68.880 110.975 ;
        RECT 70.490 110.960 70.810 111.020 ;
        RECT 100.000 111.210 100.830 114.480 ;
        RECT 104.480 114.020 109.730 114.030 ;
        RECT 104.480 113.910 116.790 114.020 ;
        RECT 101.510 113.850 116.790 113.910 ;
        RECT 101.510 113.840 116.825 113.850 ;
        RECT 101.450 113.710 116.825 113.840 ;
        RECT 101.450 113.700 106.610 113.710 ;
        RECT 101.450 113.610 105.450 113.700 ;
        RECT 108.825 113.620 116.825 113.710 ;
        RECT 108.910 113.610 116.800 113.620 ;
        RECT 101.060 113.250 101.290 113.560 ;
        RECT 101.510 113.250 105.410 113.610 ;
        RECT 105.610 113.250 105.840 113.560 ;
        RECT 101.060 111.910 105.840 113.250 ;
        RECT 101.060 111.600 101.290 111.910 ;
        RECT 105.610 111.600 105.840 111.910 ;
        RECT 108.390 113.030 108.620 113.570 ;
        RECT 109.430 113.030 110.440 113.060 ;
        RECT 117.030 113.030 117.260 113.570 ;
        RECT 108.390 112.130 117.260 113.030 ;
        RECT 108.390 111.610 108.620 112.130 ;
        RECT 109.430 112.060 110.440 112.130 ;
        RECT 117.030 111.610 117.260 112.130 ;
        RECT 101.450 111.320 105.450 111.550 ;
        RECT 108.825 111.330 116.825 111.560 ;
        RECT 100.000 111.170 101.130 111.210 ;
        RECT 100.000 111.090 101.370 111.170 ;
        RECT 101.740 111.100 105.400 111.320 ;
        RECT 101.740 111.090 103.180 111.100 ;
        RECT 100.000 111.050 103.180 111.090 ;
        RECT 100.000 110.960 102.690 111.050 ;
        RECT 108.890 111.040 116.780 111.330 ;
        RECT 100.000 110.900 102.020 110.960 ;
        RECT 70.950 110.820 71.270 110.880 ;
        RECT 73.250 110.820 73.570 110.880 ;
        RECT 73.725 110.820 74.015 110.865 ;
        RECT 68.740 110.680 74.015 110.820 ;
        RECT 70.950 110.620 71.270 110.680 ;
        RECT 73.250 110.620 73.570 110.680 ;
        RECT 73.725 110.635 74.015 110.680 ;
        RECT 100.000 110.850 101.770 110.900 ;
        RECT 69.570 110.480 69.890 110.540 ;
        RECT 67.360 110.340 69.890 110.480 ;
        RECT 69.570 110.280 69.890 110.340 ;
        RECT 75.090 110.480 75.410 110.540 ;
        RECT 75.565 110.480 75.855 110.525 ;
        RECT 75.090 110.340 75.855 110.480 ;
        RECT 75.090 110.280 75.410 110.340 ;
        RECT 75.565 110.295 75.855 110.340 ;
        RECT 79.690 110.280 80.010 110.540 ;
        RECT 81.070 110.525 81.390 110.540 ;
        RECT 81.040 110.295 81.390 110.525 ;
        RECT 81.070 110.280 81.390 110.295 ;
        RECT 56.690 110.140 57.010 110.200 ;
        RECT 57.700 110.140 57.840 110.280 ;
        RECT 56.690 110.000 57.840 110.140 ;
        RECT 62.225 110.140 62.515 110.185 ;
        RECT 65.445 110.140 65.735 110.185 ;
        RECT 62.225 110.000 65.735 110.140 ;
        RECT 56.690 109.940 57.010 110.000 ;
        RECT 62.225 109.955 62.515 110.000 ;
        RECT 65.445 109.955 65.735 110.000 ;
        RECT 41.525 109.660 46.800 109.800 ;
        RECT 59.465 109.800 59.755 109.845 ;
        RECT 62.685 109.800 62.975 109.845 ;
        RECT 64.050 109.800 64.370 109.860 ;
        RECT 59.465 109.660 64.370 109.800 ;
        RECT 65.520 109.800 65.660 109.955 ;
        RECT 66.810 109.940 67.130 110.200 ;
        RECT 67.730 110.185 68.050 110.200 ;
        RECT 67.730 109.955 68.160 110.185 ;
        RECT 72.805 109.955 73.095 110.185 ;
        RECT 74.170 110.140 74.490 110.200 ;
        RECT 74.645 110.140 74.935 110.185 ;
        RECT 74.170 110.000 74.935 110.140 ;
        RECT 67.730 109.940 68.050 109.955 ;
        RECT 68.650 109.800 68.970 109.860 ;
        RECT 65.520 109.660 68.970 109.800 ;
        RECT 41.525 109.615 41.815 109.660 ;
        RECT 59.465 109.615 59.755 109.660 ;
        RECT 62.685 109.615 62.975 109.660 ;
        RECT 64.050 109.600 64.370 109.660 ;
        RECT 68.650 109.600 68.970 109.660 ;
        RECT 70.490 109.800 70.810 109.860 ;
        RECT 72.330 109.800 72.650 109.860 ;
        RECT 72.880 109.800 73.020 109.955 ;
        RECT 74.170 109.940 74.490 110.000 ;
        RECT 74.645 109.955 74.935 110.000 ;
        RECT 80.585 110.140 80.875 110.185 ;
        RECT 81.775 110.140 82.065 110.185 ;
        RECT 84.295 110.140 84.585 110.185 ;
        RECT 87.510 110.140 87.830 110.200 ;
        RECT 89.825 110.140 90.115 110.185 ;
        RECT 80.585 110.000 84.585 110.140 ;
        RECT 80.585 109.955 80.875 110.000 ;
        RECT 81.775 109.955 82.065 110.000 ;
        RECT 84.295 109.955 84.585 110.000 ;
        RECT 86.680 110.000 90.115 110.140 ;
        RECT 75.105 109.800 75.395 109.845 ;
        RECT 78.770 109.800 79.090 109.860 ;
        RECT 86.680 109.845 86.820 110.000 ;
        RECT 87.510 109.940 87.830 110.000 ;
        RECT 89.825 109.955 90.115 110.000 ;
        RECT 70.490 109.660 73.020 109.800 ;
        RECT 74.260 109.660 79.090 109.800 ;
        RECT 70.490 109.600 70.810 109.660 ;
        RECT 72.330 109.600 72.650 109.660 ;
        RECT 27.710 109.460 28.030 109.520 ;
        RECT 21.590 109.320 28.030 109.460 ;
        RECT 17.145 109.275 17.435 109.320 ;
        RECT 18.510 109.260 18.830 109.320 ;
        RECT 27.710 109.260 28.030 109.320 ;
        RECT 28.170 109.460 28.490 109.520 ;
        RECT 28.645 109.460 28.935 109.505 ;
        RECT 28.170 109.320 28.935 109.460 ;
        RECT 28.170 109.260 28.490 109.320 ;
        RECT 28.645 109.275 28.935 109.320 ;
        RECT 29.105 109.460 29.395 109.505 ;
        RECT 40.130 109.460 40.450 109.520 ;
        RECT 29.105 109.320 40.450 109.460 ;
        RECT 29.105 109.275 29.395 109.320 ;
        RECT 40.130 109.260 40.450 109.320 ;
        RECT 40.590 109.260 40.910 109.520 ;
        RECT 44.285 109.460 44.575 109.505 ;
        RECT 44.730 109.460 45.050 109.520 ;
        RECT 45.205 109.460 45.495 109.505 ;
        RECT 44.285 109.320 45.495 109.460 ;
        RECT 44.285 109.275 44.575 109.320 ;
        RECT 44.730 109.260 45.050 109.320 ;
        RECT 45.205 109.275 45.495 109.320 ;
        RECT 65.890 109.460 66.210 109.520 ;
        RECT 74.260 109.460 74.400 109.660 ;
        RECT 75.105 109.615 75.395 109.660 ;
        RECT 78.770 109.600 79.090 109.660 ;
        RECT 80.190 109.800 80.480 109.845 ;
        RECT 82.290 109.800 82.580 109.845 ;
        RECT 83.860 109.800 84.150 109.845 ;
        RECT 80.190 109.660 84.150 109.800 ;
        RECT 80.190 109.615 80.480 109.660 ;
        RECT 82.290 109.615 82.580 109.660 ;
        RECT 83.860 109.615 84.150 109.660 ;
        RECT 86.605 109.615 86.895 109.845 ;
        RECT 65.890 109.320 74.400 109.460 ;
        RECT 65.890 109.260 66.210 109.320 ;
        RECT 74.630 109.260 74.950 109.520 ;
        RECT 87.050 109.260 87.370 109.520 ;
        RECT 13.380 108.640 92.040 109.120 ;
        RECT 21.270 108.440 21.590 108.500 ;
        RECT 21.745 108.440 22.035 108.485 ;
        RECT 21.270 108.300 22.035 108.440 ;
        RECT 21.270 108.240 21.590 108.300 ;
        RECT 21.745 108.255 22.035 108.300 ;
        RECT 23.110 108.240 23.430 108.500 ;
        RECT 24.045 108.440 24.335 108.485 ;
        RECT 27.250 108.440 27.570 108.500 ;
        RECT 24.045 108.300 27.570 108.440 ;
        RECT 24.045 108.255 24.335 108.300 ;
        RECT 15.330 108.100 15.620 108.145 ;
        RECT 17.430 108.100 17.720 108.145 ;
        RECT 19.000 108.100 19.290 108.145 ;
        RECT 15.330 107.960 19.290 108.100 ;
        RECT 15.330 107.915 15.620 107.960 ;
        RECT 17.430 107.915 17.720 107.960 ;
        RECT 19.000 107.915 19.290 107.960 ;
        RECT 22.665 108.100 22.955 108.145 ;
        RECT 24.120 108.100 24.260 108.255 ;
        RECT 27.250 108.240 27.570 108.300 ;
        RECT 27.710 108.440 28.030 108.500 ;
        RECT 30.945 108.440 31.235 108.485 ;
        RECT 27.710 108.300 31.235 108.440 ;
        RECT 27.710 108.240 28.030 108.300 ;
        RECT 30.945 108.255 31.235 108.300 ;
        RECT 31.865 108.255 32.155 108.485 ;
        RECT 36.450 108.440 36.770 108.500 ;
        RECT 36.925 108.440 37.215 108.485 ;
        RECT 36.450 108.300 37.215 108.440 ;
        RECT 26.330 108.100 26.650 108.160 ;
        RECT 28.170 108.100 28.490 108.160 ;
        RECT 31.940 108.100 32.080 108.255 ;
        RECT 36.450 108.240 36.770 108.300 ;
        RECT 36.925 108.255 37.215 108.300 ;
        RECT 39.225 108.440 39.515 108.485 ;
        RECT 42.430 108.440 42.750 108.500 ;
        RECT 39.225 108.300 42.750 108.440 ;
        RECT 39.225 108.255 39.515 108.300 ;
        RECT 42.430 108.240 42.750 108.300 ;
        RECT 50.725 108.255 51.015 108.485 ;
        RECT 22.665 107.960 24.260 108.100 ;
        RECT 25.500 107.960 32.080 108.100 ;
        RECT 22.665 107.915 22.955 107.960 ;
        RECT 15.725 107.760 16.015 107.805 ;
        RECT 16.915 107.760 17.205 107.805 ;
        RECT 19.435 107.760 19.725 107.805 ;
        RECT 15.725 107.620 19.725 107.760 ;
        RECT 15.725 107.575 16.015 107.620 ;
        RECT 16.915 107.575 17.205 107.620 ;
        RECT 19.435 107.575 19.725 107.620 ;
        RECT 23.570 107.560 23.890 107.820 ;
        RECT 14.845 107.420 15.135 107.465 ;
        RECT 21.730 107.420 22.050 107.480 ;
        RECT 14.845 107.280 22.050 107.420 ;
        RECT 14.845 107.235 15.135 107.280 ;
        RECT 21.730 107.220 22.050 107.280 ;
        RECT 22.205 107.420 22.495 107.465 ;
        RECT 22.650 107.420 22.970 107.480 ;
        RECT 24.490 107.420 24.810 107.480 ;
        RECT 22.205 107.280 24.810 107.420 ;
        RECT 22.205 107.235 22.495 107.280 ;
        RECT 22.650 107.220 22.970 107.280 ;
        RECT 24.490 107.220 24.810 107.280 ;
        RECT 24.965 107.430 25.255 107.465 ;
        RECT 25.500 107.430 25.640 107.960 ;
        RECT 26.330 107.900 26.650 107.960 ;
        RECT 28.170 107.900 28.490 107.960 ;
        RECT 36.540 107.760 36.680 108.240 ;
        RECT 39.670 108.100 39.990 108.160 ;
        RECT 40.145 108.100 40.435 108.145 ;
        RECT 39.670 107.960 40.435 108.100 ;
        RECT 39.670 107.900 39.990 107.960 ;
        RECT 40.145 107.915 40.435 107.960 ;
        RECT 40.590 108.100 40.910 108.160 ;
        RECT 50.800 108.100 50.940 108.255 ;
        RECT 58.990 108.240 59.310 108.500 ;
        RECT 63.590 108.440 63.910 108.500 ;
        RECT 65.430 108.440 65.750 108.500 ;
        RECT 66.825 108.440 67.115 108.485 ;
        RECT 63.590 108.300 67.115 108.440 ;
        RECT 63.590 108.240 63.910 108.300 ;
        RECT 65.430 108.240 65.750 108.300 ;
        RECT 66.825 108.255 67.115 108.300 ;
        RECT 69.110 108.440 69.430 108.500 ;
        RECT 70.045 108.440 70.335 108.485 ;
        RECT 69.110 108.300 70.335 108.440 ;
        RECT 57.150 108.100 57.470 108.160 ;
        RECT 40.590 107.960 57.470 108.100 ;
        RECT 40.590 107.900 40.910 107.960 ;
        RECT 57.150 107.900 57.470 107.960 ;
        RECT 25.960 107.620 33.000 107.760 ;
        RECT 25.960 107.480 26.100 107.620 ;
        RECT 24.965 107.290 25.640 107.430 ;
        RECT 24.965 107.235 25.255 107.290 ;
        RECT 25.870 107.220 26.190 107.480 ;
        RECT 28.645 107.420 28.935 107.465 ;
        RECT 30.485 107.420 30.775 107.465 ;
        RECT 26.420 107.280 28.935 107.420 ;
        RECT 15.290 107.080 15.610 107.140 ;
        RECT 16.070 107.080 16.360 107.125 ;
        RECT 15.290 106.940 16.360 107.080 ;
        RECT 15.290 106.880 15.610 106.940 ;
        RECT 16.070 106.895 16.360 106.940 ;
        RECT 16.670 107.080 16.990 107.140 ;
        RECT 26.420 107.080 26.560 107.280 ;
        RECT 28.645 107.235 28.935 107.280 ;
        RECT 29.180 107.280 30.775 107.420 ;
        RECT 16.670 106.940 26.560 107.080 ;
        RECT 16.670 106.880 16.990 106.940 ;
        RECT 26.420 106.740 26.560 106.940 ;
        RECT 26.790 107.080 27.110 107.140 ;
        RECT 29.180 107.080 29.320 107.280 ;
        RECT 30.485 107.235 30.775 107.280 ;
        RECT 30.930 107.420 31.250 107.480 ;
        RECT 32.860 107.465 33.000 107.620 ;
        RECT 35.620 107.620 36.680 107.760 ;
        RECT 36.910 107.760 37.230 107.820 ;
        RECT 66.900 107.760 67.040 108.255 ;
        RECT 69.110 108.240 69.430 108.300 ;
        RECT 70.045 108.255 70.335 108.300 ;
        RECT 72.330 108.240 72.650 108.500 ;
        RECT 73.250 108.440 73.570 108.500 ;
        RECT 75.090 108.440 75.410 108.500 ;
        RECT 73.250 108.300 75.410 108.440 ;
        RECT 73.250 108.240 73.570 108.300 ;
        RECT 75.090 108.240 75.410 108.300 ;
        RECT 81.070 108.440 81.390 108.500 ;
        RECT 82.005 108.440 82.295 108.485 ;
        RECT 81.070 108.300 82.295 108.440 ;
        RECT 81.070 108.240 81.390 108.300 ;
        RECT 82.005 108.255 82.295 108.300 ;
        RECT 88.430 108.240 88.750 108.500 ;
        RECT 68.650 108.100 68.970 108.160 ;
        RECT 71.870 108.100 72.190 108.160 ;
        RECT 74.185 108.100 74.475 108.145 ;
        RECT 75.550 108.100 75.870 108.160 ;
        RECT 68.650 107.960 73.020 108.100 ;
        RECT 68.650 107.900 68.970 107.960 ;
        RECT 71.870 107.900 72.190 107.960 ;
        RECT 72.880 107.805 73.020 107.960 ;
        RECT 74.185 107.960 78.540 108.100 ;
        RECT 74.185 107.915 74.475 107.960 ;
        RECT 75.550 107.900 75.870 107.960 ;
        RECT 36.910 107.620 52.780 107.760 ;
        RECT 66.900 107.620 72.560 107.760 ;
        RECT 35.620 107.465 35.760 107.620 ;
        RECT 36.910 107.560 37.230 107.620 ;
        RECT 31.865 107.420 32.155 107.465 ;
        RECT 30.930 107.280 32.155 107.420 ;
        RECT 30.930 107.220 31.250 107.280 ;
        RECT 31.865 107.235 32.155 107.280 ;
        RECT 32.785 107.235 33.075 107.465 ;
        RECT 35.545 107.235 35.835 107.465 ;
        RECT 36.465 107.420 36.755 107.465 ;
        RECT 37.370 107.420 37.690 107.480 ;
        RECT 36.465 107.280 37.690 107.420 ;
        RECT 36.465 107.235 36.755 107.280 ;
        RECT 37.370 107.220 37.690 107.280 ;
        RECT 38.305 107.235 38.595 107.465 ;
        RECT 39.685 107.420 39.975 107.465 ;
        RECT 41.970 107.420 42.290 107.480 ;
        RECT 39.685 107.280 42.290 107.420 ;
        RECT 39.685 107.235 39.975 107.280 ;
        RECT 26.790 106.940 29.320 107.080 ;
        RECT 29.695 107.080 29.985 107.125 ;
        RECT 31.390 107.080 31.710 107.140 ;
        RECT 38.380 107.080 38.520 107.235 ;
        RECT 41.970 107.220 42.290 107.280 ;
        RECT 42.905 107.235 43.195 107.465 ;
        RECT 38.750 107.080 39.070 107.140 ;
        RECT 42.980 107.080 43.120 107.235 ;
        RECT 44.270 107.220 44.590 107.480 ;
        RECT 44.745 107.420 45.035 107.465 ;
        RECT 45.190 107.420 45.510 107.480 ;
        RECT 44.745 107.280 45.510 107.420 ;
        RECT 44.745 107.235 45.035 107.280 ;
        RECT 45.190 107.220 45.510 107.280 ;
        RECT 45.650 107.220 45.970 107.480 ;
        RECT 52.640 107.465 52.780 107.620 ;
        RECT 52.565 107.235 52.855 107.465 ;
        RECT 66.365 107.420 66.655 107.465 ;
        RECT 66.810 107.420 67.130 107.480 ;
        RECT 68.650 107.420 68.970 107.480 ;
        RECT 72.420 107.465 72.560 107.620 ;
        RECT 72.805 107.575 73.095 107.805 ;
        RECT 73.340 107.620 75.780 107.760 ;
        RECT 66.365 107.280 72.100 107.420 ;
        RECT 66.365 107.235 66.655 107.280 ;
        RECT 66.810 107.220 67.130 107.280 ;
        RECT 68.650 107.220 68.970 107.280 ;
        RECT 47.030 107.080 47.350 107.140 ;
        RECT 29.695 106.940 31.710 107.080 ;
        RECT 26.790 106.880 27.110 106.940 ;
        RECT 29.695 106.895 29.985 106.940 ;
        RECT 31.390 106.880 31.710 106.940 ;
        RECT 36.080 106.940 38.060 107.080 ;
        RECT 38.380 106.940 47.350 107.080 ;
        RECT 36.080 106.740 36.220 106.940 ;
        RECT 26.420 106.600 36.220 106.740 ;
        RECT 36.450 106.540 36.770 106.800 ;
        RECT 37.920 106.740 38.060 106.940 ;
        RECT 38.750 106.880 39.070 106.940 ;
        RECT 47.030 106.880 47.350 106.940 ;
        RECT 49.790 106.880 50.110 107.140 ;
        RECT 56.690 107.080 57.010 107.140 ;
        RECT 71.960 107.080 72.100 107.280 ;
        RECT 72.345 107.235 72.635 107.465 ;
        RECT 73.340 107.420 73.480 107.620 ;
        RECT 75.640 107.465 75.780 107.620 ;
        RECT 78.400 107.465 78.540 107.960 ;
        RECT 84.750 107.560 85.070 107.820 ;
        RECT 100.000 107.510 100.830 110.850 ;
        RECT 108.880 110.550 116.800 110.560 ;
        RECT 105.110 110.540 116.800 110.550 ;
        RECT 101.490 110.420 116.800 110.540 ;
        RECT 101.490 110.410 116.825 110.420 ;
        RECT 101.450 110.290 116.825 110.410 ;
        RECT 101.450 110.180 105.450 110.290 ;
        RECT 101.060 109.840 101.290 110.130 ;
        RECT 101.510 109.840 105.400 110.180 ;
        RECT 105.610 109.840 105.840 110.130 ;
        RECT 101.060 108.470 105.840 109.840 ;
        RECT 101.060 108.170 101.290 108.470 ;
        RECT 105.610 108.170 105.840 108.470 ;
        RECT 101.450 107.890 105.450 108.120 ;
        RECT 101.700 107.660 105.270 107.890 ;
        RECT 101.700 107.510 105.390 107.660 ;
        RECT 74.645 107.420 74.935 107.465 ;
        RECT 72.880 107.280 73.480 107.420 ;
        RECT 73.800 107.280 74.935 107.420 ;
        RECT 72.880 107.080 73.020 107.280 ;
        RECT 50.340 106.940 57.010 107.080 ;
        RECT 50.340 106.740 50.480 106.940 ;
        RECT 56.690 106.880 57.010 106.940 ;
        RECT 69.200 106.940 71.640 107.080 ;
        RECT 71.960 106.940 73.020 107.080 ;
        RECT 69.200 106.800 69.340 106.940 ;
        RECT 37.920 106.600 50.480 106.740 ;
        RECT 50.710 106.785 51.030 106.800 ;
        RECT 50.710 106.555 51.095 106.785 ;
        RECT 50.710 106.540 51.030 106.555 ;
        RECT 51.630 106.540 51.950 106.800 ;
        RECT 69.110 106.540 69.430 106.800 ;
        RECT 70.030 106.540 70.350 106.800 ;
        RECT 71.500 106.740 71.640 106.940 ;
        RECT 73.800 106.740 73.940 107.280 ;
        RECT 74.645 107.235 74.935 107.280 ;
        RECT 75.565 107.235 75.855 107.465 ;
        RECT 78.325 107.235 78.615 107.465 ;
        RECT 78.770 107.420 79.090 107.480 ;
        RECT 83.845 107.420 84.135 107.465 ;
        RECT 87.050 107.420 87.370 107.480 ;
        RECT 78.770 107.280 79.285 107.420 ;
        RECT 83.845 107.280 87.370 107.420 ;
        RECT 78.770 107.220 79.090 107.280 ;
        RECT 83.845 107.235 84.135 107.280 ;
        RECT 87.050 107.220 87.370 107.280 ;
        RECT 87.510 107.220 87.830 107.480 ;
        RECT 100.000 107.230 105.390 107.510 ;
        RECT 106.640 107.340 107.260 110.290 ;
        RECT 108.825 110.190 116.825 110.290 ;
        RECT 108.880 110.180 116.800 110.190 ;
        RECT 108.390 109.480 108.620 110.140 ;
        RECT 109.400 109.480 110.400 109.570 ;
        RECT 117.030 109.480 117.260 110.140 ;
        RECT 108.390 108.660 117.260 109.480 ;
        RECT 108.390 108.180 108.620 108.660 ;
        RECT 109.400 108.570 110.400 108.660 ;
        RECT 117.030 108.180 117.260 108.660 ;
        RECT 108.825 107.900 116.825 108.130 ;
        RECT 71.500 106.600 73.940 106.740 ;
        RECT 76.930 106.740 77.250 106.800 ;
        RECT 80.165 106.740 80.455 106.785 ;
        RECT 76.930 106.600 80.455 106.740 ;
        RECT 76.930 106.540 77.250 106.600 ;
        RECT 80.165 106.555 80.455 106.600 ;
        RECT 82.910 106.740 83.230 106.800 ;
        RECT 84.305 106.740 84.595 106.785 ;
        RECT 82.910 106.600 84.595 106.740 ;
        RECT 82.910 106.540 83.230 106.600 ;
        RECT 84.305 106.555 84.595 106.600 ;
        RECT 100.000 106.770 105.400 107.230 ;
        RECT 13.380 105.920 92.040 106.400 ;
        RECT 15.290 105.520 15.610 105.780 ;
        RECT 23.570 105.720 23.890 105.780 ;
        RECT 24.965 105.720 25.255 105.765 ;
        RECT 23.570 105.580 25.255 105.720 ;
        RECT 23.570 105.520 23.890 105.580 ;
        RECT 24.965 105.535 25.255 105.580 ;
        RECT 38.750 105.520 39.070 105.780 ;
        RECT 39.670 105.720 39.990 105.780 ;
        RECT 40.145 105.720 40.435 105.765 ;
        RECT 39.670 105.580 40.435 105.720 ;
        RECT 39.670 105.520 39.990 105.580 ;
        RECT 40.145 105.535 40.435 105.580 ;
        RECT 41.970 105.720 42.290 105.780 ;
        RECT 42.905 105.720 43.195 105.765 ;
        RECT 45.190 105.720 45.510 105.780 ;
        RECT 57.150 105.765 57.470 105.780 ;
        RECT 50.725 105.720 51.015 105.765 ;
        RECT 41.970 105.580 43.195 105.720 ;
        RECT 41.970 105.520 42.290 105.580 ;
        RECT 42.905 105.535 43.195 105.580 ;
        RECT 43.440 105.580 51.015 105.720 ;
        RECT 16.670 105.180 16.990 105.440 ;
        RECT 17.130 105.180 17.450 105.440 ;
        RECT 17.835 105.380 18.125 105.425 ;
        RECT 19.430 105.380 19.750 105.440 ;
        RECT 22.190 105.380 22.510 105.440 ;
        RECT 25.410 105.380 25.730 105.440 ;
        RECT 36.450 105.380 36.770 105.440 ;
        RECT 17.835 105.240 19.750 105.380 ;
        RECT 17.835 105.195 18.125 105.240 ;
        RECT 19.430 105.180 19.750 105.240 ;
        RECT 21.820 105.240 22.510 105.380 ;
        RECT 16.225 104.855 16.515 105.085 ;
        RECT 16.300 104.700 16.440 104.855 ;
        RECT 18.510 104.840 18.830 105.100 ;
        RECT 20.365 105.040 20.655 105.085 ;
        RECT 21.270 105.040 21.590 105.100 ;
        RECT 21.820 105.085 21.960 105.240 ;
        RECT 22.190 105.180 22.510 105.240 ;
        RECT 22.740 105.240 26.560 105.380 ;
        RECT 22.740 105.085 22.880 105.240 ;
        RECT 25.410 105.180 25.730 105.240 ;
        RECT 26.420 105.100 26.560 105.240 ;
        RECT 36.450 105.240 41.280 105.380 ;
        RECT 36.450 105.180 36.770 105.240 ;
        RECT 20.365 104.900 21.590 105.040 ;
        RECT 20.365 104.855 20.655 104.900 ;
        RECT 21.270 104.840 21.590 104.900 ;
        RECT 21.745 104.855 22.035 105.085 ;
        RECT 22.665 104.855 22.955 105.085 ;
        RECT 23.110 104.840 23.430 105.100 ;
        RECT 26.330 104.840 26.650 105.100 ;
        RECT 26.790 105.040 27.110 105.100 ;
        RECT 31.865 105.040 32.155 105.085 ;
        RECT 26.790 104.900 32.155 105.040 ;
        RECT 26.790 104.840 27.110 104.900 ;
        RECT 31.865 104.855 32.155 104.900 ;
        RECT 33.200 105.040 33.490 105.085 ;
        RECT 33.200 104.900 37.600 105.040 ;
        RECT 33.200 104.855 33.490 104.900 ;
        RECT 17.590 104.700 17.910 104.760 ;
        RECT 22.205 104.700 22.495 104.745 ;
        RECT 23.570 104.700 23.890 104.760 ;
        RECT 24.965 104.700 25.255 104.745 ;
        RECT 16.300 104.560 20.120 104.700 ;
        RECT 17.590 104.500 17.910 104.560 ;
        RECT 14.370 104.360 14.690 104.420 ;
        RECT 19.445 104.360 19.735 104.405 ;
        RECT 14.370 104.220 19.735 104.360 ;
        RECT 19.980 104.360 20.120 104.560 ;
        RECT 22.205 104.560 25.255 104.700 ;
        RECT 22.205 104.515 22.495 104.560 ;
        RECT 23.570 104.500 23.890 104.560 ;
        RECT 24.965 104.515 25.255 104.560 ;
        RECT 25.870 104.700 26.190 104.760 ;
        RECT 30.945 104.700 31.235 104.745 ;
        RECT 25.870 104.560 31.235 104.700 ;
        RECT 25.870 104.500 26.190 104.560 ;
        RECT 30.945 104.515 31.235 104.560 ;
        RECT 32.745 104.700 33.035 104.745 ;
        RECT 33.935 104.700 34.225 104.745 ;
        RECT 36.455 104.700 36.745 104.745 ;
        RECT 32.745 104.560 36.745 104.700 ;
        RECT 37.460 104.700 37.600 104.900 ;
        RECT 39.670 104.840 39.990 105.100 ;
        RECT 41.140 105.085 41.280 105.240 ;
        RECT 41.065 104.855 41.355 105.085 ;
        RECT 42.445 105.040 42.735 105.085 ;
        RECT 42.890 105.040 43.210 105.100 ;
        RECT 43.440 105.085 43.580 105.580 ;
        RECT 45.190 105.520 45.510 105.580 ;
        RECT 50.725 105.535 51.015 105.580 ;
        RECT 57.150 105.535 57.535 105.765 ;
        RECT 64.050 105.720 64.370 105.780 ;
        RECT 67.270 105.720 67.590 105.780 ;
        RECT 76.010 105.720 76.330 105.780 ;
        RECT 78.785 105.720 79.075 105.765 ;
        RECT 84.750 105.720 85.070 105.780 ;
        RECT 64.050 105.580 77.620 105.720 ;
        RECT 57.150 105.520 57.470 105.535 ;
        RECT 64.050 105.520 64.370 105.580 ;
        RECT 67.270 105.520 67.590 105.580 ;
        RECT 76.010 105.520 76.330 105.580 ;
        RECT 56.230 105.180 56.550 105.440 ;
        RECT 66.810 105.380 67.130 105.440 ;
        RECT 67.730 105.380 68.050 105.440 ;
        RECT 66.810 105.240 77.160 105.380 ;
        RECT 66.810 105.180 67.130 105.240 ;
        RECT 67.730 105.180 68.050 105.240 ;
        RECT 77.020 105.100 77.160 105.240 ;
        RECT 42.445 104.900 43.210 105.040 ;
        RECT 42.445 104.855 42.735 104.900 ;
        RECT 42.890 104.840 43.210 104.900 ;
        RECT 43.365 104.855 43.655 105.085 ;
        RECT 45.160 105.040 45.450 105.085 ;
        RECT 46.570 105.040 46.890 105.100 ;
        RECT 45.160 104.900 46.890 105.040 ;
        RECT 45.160 104.855 45.450 104.900 ;
        RECT 46.570 104.840 46.890 104.900 ;
        RECT 65.430 104.840 65.750 105.100 ;
        RECT 69.110 105.040 69.430 105.100 ;
        RECT 73.265 105.040 73.555 105.085 ;
        RECT 69.110 104.900 73.555 105.040 ;
        RECT 69.110 104.840 69.430 104.900 ;
        RECT 73.265 104.855 73.555 104.900 ;
        RECT 74.185 105.040 74.475 105.085 ;
        RECT 75.090 105.040 75.410 105.100 ;
        RECT 74.185 104.900 75.410 105.040 ;
        RECT 74.185 104.855 74.475 104.900 ;
        RECT 75.090 104.840 75.410 104.900 ;
        RECT 75.565 104.855 75.855 105.085 ;
        RECT 41.985 104.700 42.275 104.745 ;
        RECT 37.460 104.560 42.275 104.700 ;
        RECT 32.745 104.515 33.035 104.560 ;
        RECT 33.935 104.515 34.225 104.560 ;
        RECT 36.455 104.515 36.745 104.560 ;
        RECT 41.985 104.515 42.275 104.560 ;
        RECT 43.810 104.500 44.130 104.760 ;
        RECT 44.705 104.700 44.995 104.745 ;
        RECT 45.895 104.700 46.185 104.745 ;
        RECT 48.415 104.700 48.705 104.745 ;
        RECT 44.705 104.560 48.705 104.700 ;
        RECT 44.705 104.515 44.995 104.560 ;
        RECT 45.895 104.515 46.185 104.560 ;
        RECT 48.415 104.515 48.705 104.560 ;
        RECT 53.930 104.700 54.250 104.760 ;
        RECT 54.865 104.700 55.155 104.745 ;
        RECT 53.930 104.560 55.155 104.700 ;
        RECT 53.930 104.500 54.250 104.560 ;
        RECT 54.865 104.515 55.155 104.560 ;
        RECT 55.310 104.700 55.630 104.760 ;
        RECT 58.545 104.700 58.835 104.745 ;
        RECT 55.310 104.560 58.835 104.700 ;
        RECT 55.310 104.500 55.630 104.560 ;
        RECT 58.545 104.515 58.835 104.560 ;
        RECT 66.825 104.700 67.115 104.745 ;
        RECT 69.200 104.700 69.340 104.840 ;
        RECT 66.825 104.560 69.340 104.700 ;
        RECT 73.710 104.700 74.030 104.760 ;
        RECT 75.640 104.700 75.780 104.855 ;
        RECT 76.470 104.840 76.790 105.100 ;
        RECT 76.930 104.840 77.250 105.100 ;
        RECT 77.480 105.085 77.620 105.580 ;
        RECT 78.785 105.580 85.070 105.720 ;
        RECT 78.785 105.535 79.075 105.580 ;
        RECT 84.750 105.520 85.070 105.580 ;
        RECT 100.000 105.430 102.000 106.770 ;
        RECT 103.750 106.760 105.400 106.770 ;
        RECT 102.440 105.490 103.440 106.210 ;
        RECT 103.750 105.950 104.060 106.760 ;
        RECT 104.520 106.480 105.400 106.760 ;
        RECT 105.640 106.940 107.260 107.340 ;
        RECT 108.910 106.990 116.780 107.900 ;
        RECT 104.460 106.250 105.460 106.480 ;
        RECT 105.640 106.290 105.990 106.940 ;
        RECT 106.640 106.930 107.260 106.940 ;
        RECT 108.825 106.760 116.825 106.990 ;
        RECT 108.910 106.750 116.780 106.760 ;
        RECT 104.520 106.040 105.400 106.060 ;
        RECT 103.790 105.660 104.060 105.950 ;
        RECT 104.460 105.810 105.460 106.040 ;
        RECT 105.620 106.000 105.990 106.290 ;
        RECT 105.650 105.940 105.990 106.000 ;
        RECT 106.750 106.610 107.510 106.660 ;
        RECT 108.390 106.610 108.620 106.710 ;
        RECT 106.750 106.400 108.620 106.610 ;
        RECT 117.030 106.400 117.260 106.710 ;
        RECT 106.750 105.980 109.290 106.400 ;
        RECT 116.660 105.980 117.260 106.400 ;
        RECT 104.520 105.660 105.400 105.810 ;
        RECT 104.530 105.490 105.260 105.660 ;
        RECT 100.080 105.420 102.000 105.430 ;
        RECT 77.405 104.855 77.695 105.085 ;
        RECT 80.625 104.855 80.915 105.085 ;
        RECT 73.710 104.560 75.780 104.700 ;
        RECT 66.825 104.515 67.115 104.560 ;
        RECT 73.710 104.500 74.030 104.560 ;
        RECT 24.045 104.360 24.335 104.405 ;
        RECT 24.490 104.360 24.810 104.420 ;
        RECT 32.350 104.360 32.640 104.405 ;
        RECT 34.450 104.360 34.740 104.405 ;
        RECT 36.020 104.360 36.310 104.405 ;
        RECT 19.980 104.220 28.860 104.360 ;
        RECT 14.370 104.160 14.690 104.220 ;
        RECT 19.445 104.175 19.735 104.220 ;
        RECT 24.045 104.175 24.335 104.220 ;
        RECT 24.490 104.160 24.810 104.220 ;
        RECT 25.870 103.820 26.190 104.080 ;
        RECT 26.330 104.020 26.650 104.080 ;
        RECT 28.185 104.020 28.475 104.065 ;
        RECT 26.330 103.880 28.475 104.020 ;
        RECT 28.720 104.020 28.860 104.220 ;
        RECT 32.350 104.220 36.310 104.360 ;
        RECT 32.350 104.175 32.640 104.220 ;
        RECT 34.450 104.175 34.740 104.220 ;
        RECT 36.020 104.175 36.310 104.220 ;
        RECT 44.310 104.360 44.600 104.405 ;
        RECT 46.410 104.360 46.700 104.405 ;
        RECT 47.980 104.360 48.270 104.405 ;
        RECT 44.310 104.220 48.270 104.360 ;
        RECT 44.310 104.175 44.600 104.220 ;
        RECT 46.410 104.175 46.700 104.220 ;
        RECT 47.980 104.175 48.270 104.220 ;
        RECT 58.085 104.360 58.375 104.405 ;
        RECT 80.150 104.360 80.470 104.420 ;
        RECT 80.700 104.360 80.840 104.855 ;
        RECT 87.510 104.700 87.830 104.760 ;
        RECT 88.905 104.700 89.195 104.745 ;
        RECT 87.510 104.560 89.195 104.700 ;
        RECT 87.510 104.500 87.830 104.560 ;
        RECT 88.905 104.515 89.195 104.560 ;
        RECT 102.410 104.370 105.260 105.490 ;
        RECT 105.650 105.190 106.000 105.940 ;
        RECT 106.750 105.820 108.620 105.980 ;
        RECT 106.750 105.770 107.510 105.820 ;
        RECT 108.390 105.750 108.620 105.820 ;
        RECT 117.030 105.750 117.260 105.980 ;
        RECT 108.825 105.470 116.825 105.700 ;
        RECT 105.650 105.130 105.940 105.190 ;
        RECT 105.560 105.010 105.940 105.130 ;
        RECT 108.920 105.070 116.780 105.470 ;
        RECT 117.590 105.070 118.560 114.550 ;
        RECT 119.930 114.680 120.770 116.810 ;
        RECT 126.430 116.390 127.680 116.830 ;
        RECT 137.600 116.810 138.460 118.930 ;
        RECT 124.370 116.380 129.610 116.390 ;
        RECT 121.420 116.280 136.720 116.380 ;
        RECT 121.420 116.270 136.755 116.280 ;
        RECT 121.380 116.150 136.755 116.270 ;
        RECT 121.380 116.040 125.380 116.150 ;
        RECT 126.430 116.070 128.170 116.150 ;
        RECT 128.750 116.070 136.755 116.150 ;
        RECT 126.430 115.990 127.680 116.070 ;
        RECT 128.755 116.050 136.755 116.070 ;
        RECT 120.990 115.740 121.220 115.990 ;
        RECT 125.540 115.850 125.770 115.990 ;
        RECT 128.320 115.850 128.550 116.000 ;
        RECT 125.540 115.740 128.550 115.850 ;
        RECT 136.960 115.740 137.190 116.000 ;
        RECT 120.990 115.300 137.190 115.740 ;
        RECT 120.990 115.030 121.220 115.300 ;
        RECT 125.540 115.270 137.190 115.300 ;
        RECT 125.540 115.180 128.550 115.270 ;
        RECT 125.540 115.030 125.770 115.180 ;
        RECT 128.320 115.040 128.550 115.180 ;
        RECT 136.960 115.040 137.190 115.270 ;
        RECT 121.380 114.750 125.380 114.980 ;
        RECT 128.755 114.770 136.755 114.990 ;
        RECT 137.520 114.770 138.480 116.810 ;
        RECT 128.755 114.760 138.480 114.770 ;
        RECT 121.380 114.680 125.370 114.750 ;
        RECT 119.930 114.570 125.370 114.680 ;
        RECT 128.810 114.600 138.480 114.760 ;
        RECT 119.930 114.480 123.060 114.570 ;
        RECT 136.550 114.550 138.480 114.600 ;
        RECT 119.930 111.210 120.770 114.480 ;
        RECT 124.410 114.020 129.660 114.030 ;
        RECT 124.410 113.910 136.720 114.020 ;
        RECT 121.440 113.850 136.720 113.910 ;
        RECT 121.440 113.840 136.755 113.850 ;
        RECT 121.380 113.710 136.755 113.840 ;
        RECT 121.380 113.700 126.540 113.710 ;
        RECT 121.380 113.610 125.380 113.700 ;
        RECT 128.755 113.620 136.755 113.710 ;
        RECT 128.840 113.610 136.730 113.620 ;
        RECT 120.990 113.250 121.220 113.560 ;
        RECT 121.440 113.250 125.340 113.610 ;
        RECT 125.540 113.250 125.770 113.560 ;
        RECT 120.990 111.910 125.770 113.250 ;
        RECT 120.990 111.600 121.220 111.910 ;
        RECT 125.540 111.600 125.770 111.910 ;
        RECT 128.320 113.030 128.550 113.570 ;
        RECT 129.360 113.030 130.370 113.060 ;
        RECT 136.960 113.030 137.190 113.570 ;
        RECT 128.320 112.130 137.190 113.030 ;
        RECT 128.320 111.610 128.550 112.130 ;
        RECT 129.360 112.060 130.370 112.130 ;
        RECT 136.960 111.610 137.190 112.130 ;
        RECT 121.380 111.320 125.380 111.550 ;
        RECT 128.755 111.330 136.755 111.560 ;
        RECT 119.930 111.170 121.060 111.210 ;
        RECT 119.930 111.090 121.300 111.170 ;
        RECT 121.670 111.100 125.330 111.320 ;
        RECT 121.670 111.090 123.110 111.100 ;
        RECT 119.930 111.050 123.110 111.090 ;
        RECT 119.930 110.960 122.620 111.050 ;
        RECT 128.820 111.040 136.710 111.330 ;
        RECT 119.930 110.900 121.950 110.960 ;
        RECT 119.930 110.850 121.700 110.900 ;
        RECT 119.930 107.510 120.770 110.850 ;
        RECT 128.810 110.550 136.730 110.560 ;
        RECT 125.040 110.540 136.730 110.550 ;
        RECT 121.420 110.420 136.730 110.540 ;
        RECT 121.420 110.410 136.755 110.420 ;
        RECT 121.380 110.290 136.755 110.410 ;
        RECT 121.380 110.180 125.380 110.290 ;
        RECT 120.990 109.840 121.220 110.130 ;
        RECT 121.440 109.840 125.330 110.180 ;
        RECT 125.540 109.840 125.770 110.130 ;
        RECT 120.990 108.470 125.770 109.840 ;
        RECT 120.990 108.170 121.220 108.470 ;
        RECT 125.540 108.170 125.770 108.470 ;
        RECT 121.380 107.890 125.380 108.120 ;
        RECT 121.630 107.660 125.200 107.890 ;
        RECT 121.630 107.510 125.320 107.660 ;
        RECT 119.930 107.230 125.320 107.510 ;
        RECT 126.570 107.340 127.190 110.290 ;
        RECT 128.755 110.190 136.755 110.290 ;
        RECT 128.810 110.180 136.730 110.190 ;
        RECT 128.320 109.480 128.550 110.140 ;
        RECT 129.330 109.480 130.330 109.570 ;
        RECT 136.960 109.480 137.190 110.140 ;
        RECT 128.320 108.660 137.190 109.480 ;
        RECT 128.320 108.180 128.550 108.660 ;
        RECT 129.330 108.570 130.330 108.660 ;
        RECT 136.960 108.180 137.190 108.660 ;
        RECT 128.755 107.900 136.755 108.130 ;
        RECT 119.930 106.770 125.330 107.230 ;
        RECT 119.930 105.880 121.930 106.770 ;
        RECT 123.680 106.760 125.330 106.770 ;
        RECT 58.085 104.220 80.840 104.360 ;
        RECT 58.085 104.175 58.375 104.220 ;
        RECT 80.150 104.160 80.470 104.220 ;
        RECT 102.350 104.140 105.350 104.370 ;
        RECT 105.560 104.180 105.900 105.010 ;
        RECT 107.910 105.000 118.560 105.070 ;
        RECT 102.400 104.110 105.260 104.140 ;
        RECT 102.400 104.090 103.570 104.110 ;
        RECT 104.530 104.100 105.260 104.110 ;
        RECT 49.790 104.020 50.110 104.080 ;
        RECT 28.720 103.880 50.110 104.020 ;
        RECT 26.330 103.820 26.650 103.880 ;
        RECT 28.185 103.835 28.475 103.880 ;
        RECT 49.790 103.820 50.110 103.880 ;
        RECT 52.090 103.820 52.410 104.080 ;
        RECT 56.690 104.020 57.010 104.080 ;
        RECT 57.165 104.020 57.455 104.065 ;
        RECT 56.690 103.880 57.455 104.020 ;
        RECT 56.690 103.820 57.010 103.880 ;
        RECT 57.165 103.835 57.455 103.880 ;
        RECT 61.750 103.820 62.070 104.080 ;
        RECT 65.430 104.020 65.750 104.080 ;
        RECT 65.905 104.020 66.195 104.065 ;
        RECT 65.430 103.880 66.195 104.020 ;
        RECT 65.430 103.820 65.750 103.880 ;
        RECT 65.905 103.835 66.195 103.880 ;
        RECT 66.365 104.020 66.655 104.065 ;
        RECT 67.730 104.020 68.050 104.080 ;
        RECT 66.365 103.880 68.050 104.020 ;
        RECT 66.365 103.835 66.655 103.880 ;
        RECT 67.730 103.820 68.050 103.880 ;
        RECT 73.710 104.020 74.030 104.080 ;
        RECT 74.645 104.020 74.935 104.065 ;
        RECT 73.710 103.880 74.935 104.020 ;
        RECT 73.710 103.820 74.030 103.880 ;
        RECT 74.645 103.835 74.935 103.880 ;
        RECT 75.090 104.020 75.410 104.080 ;
        RECT 76.930 104.020 77.250 104.080 ;
        RECT 79.705 104.020 79.995 104.065 ;
        RECT 75.090 103.880 79.995 104.020 ;
        RECT 75.090 103.820 75.410 103.880 ;
        RECT 76.930 103.820 77.250 103.880 ;
        RECT 79.705 103.835 79.995 103.880 ;
        RECT 84.290 104.020 84.610 104.080 ;
        RECT 86.145 104.020 86.435 104.065 ;
        RECT 84.290 103.880 86.435 104.020 ;
        RECT 84.290 103.820 84.610 103.880 ;
        RECT 86.145 103.835 86.435 103.880 ;
        RECT 102.350 103.700 105.350 103.930 ;
        RECT 105.555 103.890 105.900 104.180 ;
        RECT 106.090 104.040 118.560 105.000 ;
        RECT 119.900 105.420 121.930 105.880 ;
        RECT 122.370 105.490 123.370 106.210 ;
        RECT 123.680 105.950 123.990 106.760 ;
        RECT 124.450 106.480 125.330 106.760 ;
        RECT 125.570 106.940 127.190 107.340 ;
        RECT 128.840 106.990 136.710 107.900 ;
        RECT 124.390 106.250 125.390 106.480 ;
        RECT 125.570 106.290 125.920 106.940 ;
        RECT 126.570 106.930 127.190 106.940 ;
        RECT 128.755 106.760 136.755 106.990 ;
        RECT 128.840 106.750 136.710 106.760 ;
        RECT 124.450 106.040 125.330 106.060 ;
        RECT 123.720 105.660 123.990 105.950 ;
        RECT 124.390 105.810 125.390 106.040 ;
        RECT 125.550 106.000 125.920 106.290 ;
        RECT 125.580 105.940 125.920 106.000 ;
        RECT 126.680 106.610 127.440 106.660 ;
        RECT 128.320 106.610 128.550 106.710 ;
        RECT 126.680 106.400 128.550 106.610 ;
        RECT 136.960 106.400 137.190 106.710 ;
        RECT 126.680 105.980 129.220 106.400 ;
        RECT 136.590 105.980 137.190 106.400 ;
        RECT 124.450 105.660 125.330 105.810 ;
        RECT 124.460 105.490 125.190 105.660 ;
        RECT 106.090 103.960 118.550 104.040 ;
        RECT 106.090 103.940 118.420 103.960 ;
        RECT 105.560 103.780 105.900 103.890 ;
        RECT 106.130 103.930 111.800 103.940 ;
        RECT 112.800 103.930 118.420 103.940 ;
        RECT 13.380 103.200 92.040 103.680 ;
        RECT 102.440 103.530 105.300 103.700 ;
        RECT 106.130 103.530 107.465 103.930 ;
        RECT 102.410 103.160 107.465 103.530 ;
        RECT 15.765 103.000 16.055 103.045 ;
        RECT 21.730 103.000 22.050 103.060 ;
        RECT 22.650 103.000 22.970 103.060 ;
        RECT 33.705 103.000 33.995 103.045 ;
        RECT 15.765 102.860 22.970 103.000 ;
        RECT 15.765 102.815 16.055 102.860 ;
        RECT 21.730 102.800 22.050 102.860 ;
        RECT 22.650 102.800 22.970 102.860 ;
        RECT 24.120 102.860 33.995 103.000 ;
        RECT 24.120 102.720 24.260 102.860 ;
        RECT 33.705 102.815 33.995 102.860 ;
        RECT 38.765 103.000 39.055 103.045 ;
        RECT 39.670 103.000 39.990 103.060 ;
        RECT 38.765 102.860 39.990 103.000 ;
        RECT 38.765 102.815 39.055 102.860 ;
        RECT 39.670 102.800 39.990 102.860 ;
        RECT 40.145 103.000 40.435 103.045 ;
        RECT 43.350 103.000 43.670 103.060 ;
        RECT 40.145 102.860 43.670 103.000 ;
        RECT 40.145 102.815 40.435 102.860 ;
        RECT 43.350 102.800 43.670 102.860 ;
        RECT 46.570 102.800 46.890 103.060 ;
        RECT 50.710 103.000 51.030 103.060 ;
        RECT 51.185 103.000 51.475 103.045 ;
        RECT 50.710 102.860 51.475 103.000 ;
        RECT 50.710 102.800 51.030 102.860 ;
        RECT 51.185 102.815 51.475 102.860 ;
        RECT 53.485 103.000 53.775 103.045 ;
        RECT 55.310 103.000 55.630 103.060 ;
        RECT 53.485 102.860 55.630 103.000 ;
        RECT 53.485 102.815 53.775 102.860 ;
        RECT 55.310 102.800 55.630 102.860 ;
        RECT 87.510 102.800 87.830 103.060 ;
        RECT 106.195 102.975 107.465 103.160 ;
        RECT 24.030 102.660 24.350 102.720 ;
        RECT 18.600 102.520 24.350 102.660 ;
        RECT 12.070 101.980 12.390 102.040 ;
        RECT 15.305 101.980 15.595 102.025 ;
        RECT 12.070 101.840 15.595 101.980 ;
        RECT 12.070 101.780 12.390 101.840 ;
        RECT 15.305 101.795 15.595 101.840 ;
        RECT 17.605 101.980 17.895 102.025 ;
        RECT 18.050 101.980 18.370 102.040 ;
        RECT 18.600 102.025 18.740 102.520 ;
        RECT 24.030 102.460 24.350 102.520 ;
        RECT 27.290 102.660 27.580 102.705 ;
        RECT 29.390 102.660 29.680 102.705 ;
        RECT 30.960 102.660 31.250 102.705 ;
        RECT 45.205 102.660 45.495 102.705 ;
        RECT 27.290 102.520 31.250 102.660 ;
        RECT 27.290 102.475 27.580 102.520 ;
        RECT 29.390 102.475 29.680 102.520 ;
        RECT 30.960 102.475 31.250 102.520 ;
        RECT 41.600 102.520 45.495 102.660 ;
        RECT 23.570 102.120 23.890 102.380 ;
        RECT 26.790 102.120 27.110 102.380 ;
        RECT 27.685 102.320 27.975 102.365 ;
        RECT 28.875 102.320 29.165 102.365 ;
        RECT 31.395 102.320 31.685 102.365 ;
        RECT 41.600 102.320 41.740 102.520 ;
        RECT 45.205 102.475 45.495 102.520 ;
        RECT 56.230 102.660 56.520 102.705 ;
        RECT 57.800 102.660 58.090 102.705 ;
        RECT 59.900 102.660 60.190 102.705 ;
        RECT 56.230 102.520 60.190 102.660 ;
        RECT 56.230 102.475 56.520 102.520 ;
        RECT 57.800 102.475 58.090 102.520 ;
        RECT 59.900 102.475 60.190 102.520 ;
        RECT 65.905 102.660 66.195 102.705 ;
        RECT 68.190 102.660 68.510 102.720 ;
        RECT 77.390 102.660 77.710 102.720 ;
        RECT 65.905 102.520 68.510 102.660 ;
        RECT 65.905 102.475 66.195 102.520 ;
        RECT 68.190 102.460 68.510 102.520 ;
        RECT 74.260 102.520 77.710 102.660 ;
        RECT 44.730 102.320 45.050 102.380 ;
        RECT 27.685 102.180 31.685 102.320 ;
        RECT 27.685 102.135 27.975 102.180 ;
        RECT 28.875 102.135 29.165 102.180 ;
        RECT 31.395 102.135 31.685 102.180 ;
        RECT 39.300 102.180 41.740 102.320 ;
        RECT 17.605 101.840 18.370 101.980 ;
        RECT 17.605 101.795 17.895 101.840 ;
        RECT 18.050 101.780 18.370 101.840 ;
        RECT 18.525 101.795 18.815 102.025 ;
        RECT 19.430 101.780 19.750 102.040 ;
        RECT 24.045 101.980 24.335 102.025 ;
        RECT 26.330 101.980 26.650 102.040 ;
        RECT 39.300 102.025 39.440 102.180 ;
        RECT 24.045 101.840 26.650 101.980 ;
        RECT 24.045 101.795 24.335 101.840 ;
        RECT 26.330 101.780 26.650 101.840 ;
        RECT 38.305 101.795 38.595 102.025 ;
        RECT 39.225 101.795 39.515 102.025 ;
        RECT 18.140 101.640 18.280 101.780 ;
        RECT 23.570 101.640 23.890 101.700 ;
        RECT 28.030 101.640 28.320 101.685 ;
        RECT 18.140 101.500 23.890 101.640 ;
        RECT 23.570 101.440 23.890 101.500 ;
        RECT 25.960 101.500 28.320 101.640 ;
        RECT 38.380 101.640 38.520 101.795 ;
        RECT 41.050 101.780 41.370 102.040 ;
        RECT 41.600 102.025 41.740 102.180 ;
        RECT 42.520 102.180 45.050 102.320 ;
        RECT 41.525 101.980 41.815 102.025 ;
        RECT 41.970 101.980 42.290 102.040 ;
        RECT 42.520 102.025 42.660 102.180 ;
        RECT 44.730 102.120 45.050 102.180 ;
        RECT 55.795 102.320 56.085 102.365 ;
        RECT 58.315 102.320 58.605 102.365 ;
        RECT 59.505 102.320 59.795 102.365 ;
        RECT 55.795 102.180 59.795 102.320 ;
        RECT 55.795 102.135 56.085 102.180 ;
        RECT 58.315 102.135 58.605 102.180 ;
        RECT 59.505 102.135 59.795 102.180 ;
        RECT 61.750 102.320 62.070 102.380 ;
        RECT 63.145 102.320 63.435 102.365 ;
        RECT 61.750 102.180 63.435 102.320 ;
        RECT 61.750 102.120 62.070 102.180 ;
        RECT 63.145 102.135 63.435 102.180 ;
        RECT 64.065 102.320 64.355 102.365 ;
        RECT 73.265 102.320 73.555 102.365 ;
        RECT 64.065 102.180 73.555 102.320 ;
        RECT 64.065 102.135 64.355 102.180 ;
        RECT 73.265 102.135 73.555 102.180 ;
        RECT 41.525 101.840 42.290 101.980 ;
        RECT 41.525 101.795 41.815 101.840 ;
        RECT 41.970 101.780 42.290 101.840 ;
        RECT 42.445 101.795 42.735 102.025 ;
        RECT 42.890 101.780 43.210 102.040 ;
        RECT 43.365 101.795 43.655 102.025 ;
        RECT 44.285 101.980 44.575 102.025 ;
        RECT 45.190 101.980 45.510 102.040 ;
        RECT 44.285 101.840 45.510 101.980 ;
        RECT 44.285 101.795 44.575 101.840 ;
        RECT 43.440 101.640 43.580 101.795 ;
        RECT 45.190 101.780 45.510 101.840 ;
        RECT 45.650 101.780 45.970 102.040 ;
        RECT 51.645 101.980 51.935 102.025 ;
        RECT 57.150 101.980 57.470 102.040 ;
        RECT 60.385 101.980 60.675 102.025 ;
        RECT 51.645 101.840 56.000 101.980 ;
        RECT 51.645 101.795 51.935 101.840 ;
        RECT 55.860 101.700 56.000 101.840 ;
        RECT 57.150 101.840 60.675 101.980 ;
        RECT 57.150 101.780 57.470 101.840 ;
        RECT 60.385 101.795 60.675 101.840 ;
        RECT 64.970 101.780 65.290 102.040 ;
        RECT 66.810 101.780 67.130 102.040 ;
        RECT 67.270 101.980 67.590 102.040 ;
        RECT 74.260 102.025 74.400 102.520 ;
        RECT 77.390 102.460 77.710 102.520 ;
        RECT 81.110 102.660 81.400 102.705 ;
        RECT 83.210 102.660 83.500 102.705 ;
        RECT 84.780 102.660 85.070 102.705 ;
        RECT 81.110 102.520 85.070 102.660 ;
        RECT 81.110 102.475 81.400 102.520 ;
        RECT 83.210 102.475 83.500 102.520 ;
        RECT 84.780 102.475 85.070 102.520 ;
        RECT 74.645 102.320 74.935 102.365 ;
        RECT 75.090 102.320 75.410 102.380 ;
        RECT 76.930 102.320 77.250 102.380 ;
        RECT 74.645 102.180 75.410 102.320 ;
        RECT 74.645 102.135 74.935 102.180 ;
        RECT 75.090 102.120 75.410 102.180 ;
        RECT 75.640 102.180 77.250 102.320 ;
        RECT 75.640 102.025 75.780 102.180 ;
        RECT 76.930 102.120 77.250 102.180 ;
        RECT 81.505 102.320 81.795 102.365 ;
        RECT 82.695 102.320 82.985 102.365 ;
        RECT 85.215 102.320 85.505 102.365 ;
        RECT 81.505 102.180 85.505 102.320 ;
        RECT 81.505 102.135 81.795 102.180 ;
        RECT 82.695 102.135 82.985 102.180 ;
        RECT 85.215 102.135 85.505 102.180 ;
        RECT 67.745 101.980 68.035 102.025 ;
        RECT 67.270 101.840 68.035 101.980 ;
        RECT 67.270 101.780 67.590 101.840 ;
        RECT 67.745 101.795 68.035 101.840 ;
        RECT 72.805 101.795 73.095 102.025 ;
        RECT 73.725 101.795 74.015 102.025 ;
        RECT 74.185 101.795 74.475 102.025 ;
        RECT 75.565 101.795 75.855 102.025 ;
        RECT 76.025 101.795 76.315 102.025 ;
        RECT 38.380 101.500 43.580 101.640 ;
        RECT 18.510 101.100 18.830 101.360 ;
        RECT 22.190 101.100 22.510 101.360 ;
        RECT 25.960 101.345 26.100 101.500 ;
        RECT 28.030 101.455 28.320 101.500 ;
        RECT 41.600 101.360 41.740 101.500 ;
        RECT 55.770 101.440 56.090 101.700 ;
        RECT 59.160 101.640 59.450 101.685 ;
        RECT 62.685 101.640 62.975 101.685 ;
        RECT 66.900 101.640 67.040 101.780 ;
        RECT 59.160 101.500 61.060 101.640 ;
        RECT 59.160 101.455 59.450 101.500 ;
        RECT 25.885 101.115 26.175 101.345 ;
        RECT 41.510 101.100 41.830 101.360 ;
        RECT 60.920 101.345 61.060 101.500 ;
        RECT 62.685 101.500 67.040 101.640 ;
        RECT 62.685 101.455 62.975 101.500 ;
        RECT 60.845 101.115 61.135 101.345 ;
        RECT 66.350 101.300 66.670 101.360 ;
        RECT 67.285 101.300 67.575 101.345 ;
        RECT 66.350 101.160 67.575 101.300 ;
        RECT 72.880 101.300 73.020 101.795 ;
        RECT 73.800 101.640 73.940 101.795 ;
        RECT 74.630 101.640 74.950 101.700 ;
        RECT 76.100 101.640 76.240 101.795 ;
        RECT 80.610 101.780 80.930 102.040 ;
        RECT 73.800 101.500 76.240 101.640 ;
        RECT 81.960 101.640 82.250 101.685 ;
        RECT 82.450 101.640 82.770 101.700 ;
        RECT 81.960 101.500 82.770 101.640 ;
        RECT 74.630 101.440 74.950 101.500 ;
        RECT 81.960 101.455 82.250 101.500 ;
        RECT 82.450 101.440 82.770 101.500 ;
        RECT 75.090 101.300 75.410 101.360 ;
        RECT 72.880 101.160 75.410 101.300 ;
        RECT 66.350 101.100 66.670 101.160 ;
        RECT 67.285 101.115 67.575 101.160 ;
        RECT 75.090 101.100 75.410 101.160 ;
        RECT 76.945 101.300 77.235 101.345 ;
        RECT 85.210 101.300 85.530 101.360 ;
        RECT 76.945 101.160 85.530 101.300 ;
        RECT 76.945 101.115 77.235 101.160 ;
        RECT 85.210 101.100 85.530 101.160 ;
        RECT 106.195 101.085 107.455 102.975 ;
        RECT 119.900 102.760 120.990 105.420 ;
        RECT 122.340 104.370 125.190 105.490 ;
        RECT 125.580 105.190 125.930 105.940 ;
        RECT 126.680 105.820 128.550 105.980 ;
        RECT 126.680 105.770 127.440 105.820 ;
        RECT 128.320 105.750 128.550 105.820 ;
        RECT 136.960 105.750 137.190 105.980 ;
        RECT 128.755 105.470 136.755 105.700 ;
        RECT 125.580 105.130 125.870 105.190 ;
        RECT 125.490 105.010 125.870 105.130 ;
        RECT 128.850 105.070 136.710 105.470 ;
        RECT 137.520 105.070 138.480 114.550 ;
        RECT 139.930 116.780 140.700 120.420 ;
        RECT 142.370 119.370 145.220 120.490 ;
        RECT 145.610 120.190 145.960 120.940 ;
        RECT 146.710 120.820 148.580 120.980 ;
        RECT 146.710 120.770 147.470 120.820 ;
        RECT 148.350 120.750 148.580 120.820 ;
        RECT 156.990 120.750 157.220 120.980 ;
        RECT 148.785 120.470 156.785 120.700 ;
        RECT 145.610 120.130 145.900 120.190 ;
        RECT 145.520 120.010 145.900 120.130 ;
        RECT 148.880 120.070 156.740 120.470 ;
        RECT 157.550 120.070 158.510 129.550 ;
        RECT 142.310 119.140 145.310 119.370 ;
        RECT 145.520 119.180 145.860 120.010 ;
        RECT 147.870 120.000 158.510 120.070 ;
        RECT 142.360 119.110 145.220 119.140 ;
        RECT 142.360 119.090 143.530 119.110 ;
        RECT 144.490 119.100 145.220 119.110 ;
        RECT 142.310 118.700 145.310 118.930 ;
        RECT 145.515 118.890 145.860 119.180 ;
        RECT 146.050 118.960 158.510 120.000 ;
        RECT 146.050 118.940 158.500 118.960 ;
        RECT 145.520 118.780 145.860 118.890 ;
        RECT 146.090 118.930 151.760 118.940 ;
        RECT 152.760 118.930 158.500 118.940 ;
        RECT 142.400 118.530 145.260 118.700 ;
        RECT 146.090 118.530 146.520 118.930 ;
        RECT 142.370 118.160 146.520 118.530 ;
        RECT 139.930 114.680 140.790 116.780 ;
        RECT 146.460 116.390 147.710 116.830 ;
        RECT 157.640 116.810 158.500 118.930 ;
        RECT 144.400 116.380 149.640 116.390 ;
        RECT 141.450 116.280 156.750 116.380 ;
        RECT 141.450 116.270 156.785 116.280 ;
        RECT 141.410 116.150 156.785 116.270 ;
        RECT 141.410 116.040 145.410 116.150 ;
        RECT 146.460 116.070 148.200 116.150 ;
        RECT 148.780 116.070 156.785 116.150 ;
        RECT 146.460 115.990 147.710 116.070 ;
        RECT 148.785 116.050 156.785 116.070 ;
        RECT 141.020 115.740 141.250 115.990 ;
        RECT 145.570 115.850 145.800 115.990 ;
        RECT 148.350 115.850 148.580 116.000 ;
        RECT 145.570 115.740 148.580 115.850 ;
        RECT 156.990 115.740 157.220 116.000 ;
        RECT 141.020 115.300 157.220 115.740 ;
        RECT 141.020 115.030 141.250 115.300 ;
        RECT 145.570 115.270 157.220 115.300 ;
        RECT 145.570 115.180 148.580 115.270 ;
        RECT 145.570 115.030 145.800 115.180 ;
        RECT 148.350 115.040 148.580 115.180 ;
        RECT 156.990 115.040 157.220 115.270 ;
        RECT 141.410 114.750 145.410 114.980 ;
        RECT 148.785 114.770 156.785 114.990 ;
        RECT 157.550 114.770 158.510 116.810 ;
        RECT 148.785 114.760 158.510 114.770 ;
        RECT 141.410 114.680 145.400 114.750 ;
        RECT 139.930 114.570 145.400 114.680 ;
        RECT 148.840 114.600 158.510 114.760 ;
        RECT 139.930 114.480 143.090 114.570 ;
        RECT 156.580 114.550 158.510 114.600 ;
        RECT 139.930 111.210 140.790 114.480 ;
        RECT 144.440 114.020 149.690 114.030 ;
        RECT 144.440 113.910 156.750 114.020 ;
        RECT 141.470 113.850 156.750 113.910 ;
        RECT 141.470 113.840 156.785 113.850 ;
        RECT 141.410 113.710 156.785 113.840 ;
        RECT 141.410 113.700 146.570 113.710 ;
        RECT 141.410 113.610 145.410 113.700 ;
        RECT 148.785 113.620 156.785 113.710 ;
        RECT 148.870 113.610 156.760 113.620 ;
        RECT 141.020 113.250 141.250 113.560 ;
        RECT 141.470 113.250 145.370 113.610 ;
        RECT 145.570 113.250 145.800 113.560 ;
        RECT 141.020 111.910 145.800 113.250 ;
        RECT 141.020 111.600 141.250 111.910 ;
        RECT 145.570 111.600 145.800 111.910 ;
        RECT 148.350 113.030 148.580 113.570 ;
        RECT 149.390 113.030 150.400 113.060 ;
        RECT 156.990 113.030 157.220 113.570 ;
        RECT 148.350 112.130 157.220 113.030 ;
        RECT 148.350 111.610 148.580 112.130 ;
        RECT 149.390 112.060 150.400 112.130 ;
        RECT 156.990 111.610 157.220 112.130 ;
        RECT 141.410 111.320 145.410 111.550 ;
        RECT 148.785 111.330 156.785 111.560 ;
        RECT 139.930 111.170 141.090 111.210 ;
        RECT 139.930 111.090 141.330 111.170 ;
        RECT 141.700 111.100 145.360 111.320 ;
        RECT 141.700 111.090 143.140 111.100 ;
        RECT 139.930 111.050 143.140 111.090 ;
        RECT 139.930 110.960 142.650 111.050 ;
        RECT 148.850 111.040 156.740 111.330 ;
        RECT 139.930 110.900 141.980 110.960 ;
        RECT 139.930 110.850 141.730 110.900 ;
        RECT 139.930 107.510 140.790 110.850 ;
        RECT 148.840 110.550 156.760 110.560 ;
        RECT 145.070 110.540 156.760 110.550 ;
        RECT 141.450 110.420 156.760 110.540 ;
        RECT 141.450 110.410 156.785 110.420 ;
        RECT 141.410 110.290 156.785 110.410 ;
        RECT 141.410 110.180 145.410 110.290 ;
        RECT 141.020 109.840 141.250 110.130 ;
        RECT 141.470 109.840 145.360 110.180 ;
        RECT 145.570 109.840 145.800 110.130 ;
        RECT 141.020 108.470 145.800 109.840 ;
        RECT 141.020 108.170 141.250 108.470 ;
        RECT 145.570 108.170 145.800 108.470 ;
        RECT 141.410 107.890 145.410 108.120 ;
        RECT 141.660 107.660 145.230 107.890 ;
        RECT 141.660 107.510 145.350 107.660 ;
        RECT 139.930 107.230 145.350 107.510 ;
        RECT 146.600 107.340 147.220 110.290 ;
        RECT 148.785 110.190 156.785 110.290 ;
        RECT 148.840 110.180 156.760 110.190 ;
        RECT 148.350 109.480 148.580 110.140 ;
        RECT 149.360 109.480 150.360 109.570 ;
        RECT 156.990 109.480 157.220 110.140 ;
        RECT 148.350 108.660 157.220 109.480 ;
        RECT 148.350 108.180 148.580 108.660 ;
        RECT 149.360 108.570 150.360 108.660 ;
        RECT 156.990 108.180 157.220 108.660 ;
        RECT 148.785 107.900 156.785 108.130 ;
        RECT 139.930 106.770 145.360 107.230 ;
        RECT 139.930 106.630 141.960 106.770 ;
        RECT 139.960 105.430 141.960 106.630 ;
        RECT 143.710 106.760 145.360 106.770 ;
        RECT 142.400 105.490 143.400 106.210 ;
        RECT 143.710 105.950 144.020 106.760 ;
        RECT 144.480 106.480 145.360 106.760 ;
        RECT 145.600 106.940 147.220 107.340 ;
        RECT 148.870 106.990 156.740 107.900 ;
        RECT 144.420 106.250 145.420 106.480 ;
        RECT 145.600 106.290 145.950 106.940 ;
        RECT 146.600 106.930 147.220 106.940 ;
        RECT 148.785 106.760 156.785 106.990 ;
        RECT 148.870 106.750 156.740 106.760 ;
        RECT 144.480 106.040 145.360 106.060 ;
        RECT 143.750 105.660 144.020 105.950 ;
        RECT 144.420 105.810 145.420 106.040 ;
        RECT 145.580 106.000 145.950 106.290 ;
        RECT 145.610 105.940 145.950 106.000 ;
        RECT 146.710 106.610 147.470 106.660 ;
        RECT 148.350 106.610 148.580 106.710 ;
        RECT 146.710 106.400 148.580 106.610 ;
        RECT 156.990 106.400 157.220 106.710 ;
        RECT 146.710 105.980 149.250 106.400 ;
        RECT 156.620 105.980 157.220 106.400 ;
        RECT 144.480 105.660 145.360 105.810 ;
        RECT 144.490 105.490 145.220 105.660 ;
        RECT 140.040 105.420 141.960 105.430 ;
        RECT 122.280 104.140 125.280 104.370 ;
        RECT 125.490 104.180 125.830 105.010 ;
        RECT 127.840 105.000 138.480 105.070 ;
        RECT 122.330 104.110 125.190 104.140 ;
        RECT 122.330 104.090 123.500 104.110 ;
        RECT 124.460 104.100 125.190 104.110 ;
        RECT 122.280 103.700 125.280 103.930 ;
        RECT 125.485 103.890 125.830 104.180 ;
        RECT 126.020 103.960 138.480 105.000 ;
        RECT 142.370 104.370 145.220 105.490 ;
        RECT 145.610 105.190 145.960 105.940 ;
        RECT 146.710 105.820 148.580 105.980 ;
        RECT 146.710 105.770 147.470 105.820 ;
        RECT 148.350 105.750 148.580 105.820 ;
        RECT 156.990 105.750 157.220 105.980 ;
        RECT 148.785 105.470 156.785 105.700 ;
        RECT 145.610 105.130 145.900 105.190 ;
        RECT 145.520 105.010 145.900 105.130 ;
        RECT 148.880 105.070 156.740 105.470 ;
        RECT 157.550 105.070 158.510 114.550 ;
        RECT 142.310 104.140 145.310 104.370 ;
        RECT 145.520 104.180 145.860 105.010 ;
        RECT 147.870 105.000 158.510 105.070 ;
        RECT 142.360 104.110 145.220 104.140 ;
        RECT 142.360 104.090 143.530 104.110 ;
        RECT 144.490 104.100 145.220 104.110 ;
        RECT 126.020 103.940 138.350 103.960 ;
        RECT 125.490 103.780 125.830 103.890 ;
        RECT 126.060 103.930 131.730 103.940 ;
        RECT 132.730 103.930 138.350 103.940 ;
        RECT 122.370 103.530 125.230 103.700 ;
        RECT 126.060 103.530 126.490 103.930 ;
        RECT 142.310 103.700 145.310 103.930 ;
        RECT 145.515 103.890 145.860 104.180 ;
        RECT 146.050 103.960 158.510 105.000 ;
        RECT 146.050 103.940 158.460 103.960 ;
        RECT 145.520 103.780 145.860 103.890 ;
        RECT 146.090 103.930 151.760 103.940 ;
        RECT 152.760 103.930 158.460 103.940 ;
        RECT 142.400 103.530 145.260 103.700 ;
        RECT 146.090 103.530 146.520 103.930 ;
        RECT 122.340 103.160 126.490 103.530 ;
        RECT 142.370 103.160 146.520 103.530 ;
        RECT 113.040 102.695 116.730 102.710 ;
        RECT 119.900 102.695 135.450 102.760 ;
        RECT 113.040 101.710 135.450 102.695 ;
        RECT 113.040 101.690 132.370 101.710 ;
        RECT 113.040 101.675 123.360 101.690 ;
        RECT 113.040 101.660 116.730 101.675 ;
        RECT 99.990 101.065 112.800 101.085 ;
        RECT 13.380 100.480 92.040 100.960 ;
        RECT 23.570 100.080 23.890 100.340 ;
        RECT 24.030 100.080 24.350 100.340 ;
        RECT 41.050 100.280 41.370 100.340 ;
        RECT 42.905 100.280 43.195 100.325 ;
        RECT 41.050 100.140 43.195 100.280 ;
        RECT 41.050 100.080 41.370 100.140 ;
        RECT 42.905 100.095 43.195 100.140 ;
        RECT 44.745 100.280 45.035 100.325 ;
        RECT 53.930 100.280 54.250 100.340 ;
        RECT 44.745 100.140 54.250 100.280 ;
        RECT 44.745 100.095 45.035 100.140 ;
        RECT 53.930 100.080 54.250 100.140 ;
        RECT 64.525 100.280 64.815 100.325 ;
        RECT 64.970 100.280 65.290 100.340 ;
        RECT 64.525 100.140 65.290 100.280 ;
        RECT 64.525 100.095 64.815 100.140 ;
        RECT 64.970 100.080 65.290 100.140 ;
        RECT 65.445 100.095 65.735 100.325 ;
        RECT 65.890 100.280 66.210 100.340 ;
        RECT 67.730 100.280 68.050 100.340 ;
        RECT 65.890 100.140 68.050 100.280 ;
        RECT 16.180 99.940 16.470 99.985 ;
        RECT 26.345 99.940 26.635 99.985 ;
        RECT 16.180 99.800 26.635 99.940 ;
        RECT 16.180 99.755 16.470 99.800 ;
        RECT 26.345 99.755 26.635 99.800 ;
        RECT 43.810 99.940 44.130 100.000 ;
        RECT 48.870 99.940 49.190 100.000 ;
        RECT 43.810 99.800 49.190 99.940 ;
        RECT 43.810 99.740 44.130 99.800 ;
        RECT 14.830 99.400 15.150 99.660 ;
        RECT 22.190 99.600 22.510 99.660 ;
        RECT 25.885 99.600 26.175 99.645 ;
        RECT 22.190 99.460 26.175 99.600 ;
        RECT 22.190 99.400 22.510 99.460 ;
        RECT 25.885 99.415 26.175 99.460 ;
        RECT 26.805 99.415 27.095 99.645 ;
        RECT 45.205 99.600 45.495 99.645 ;
        RECT 46.110 99.600 46.430 99.660 ;
        RECT 47.120 99.645 47.260 99.800 ;
        RECT 48.870 99.740 49.190 99.800 ;
        RECT 56.690 99.940 57.010 100.000 ;
        RECT 57.165 99.940 57.455 99.985 ;
        RECT 56.690 99.800 57.455 99.940 ;
        RECT 56.690 99.740 57.010 99.800 ;
        RECT 57.165 99.755 57.455 99.800 ;
        RECT 58.960 99.940 59.250 99.985 ;
        RECT 65.520 99.940 65.660 100.095 ;
        RECT 65.890 100.080 66.210 100.140 ;
        RECT 67.730 100.080 68.050 100.140 ;
        RECT 74.630 100.080 74.950 100.340 ;
        RECT 76.470 100.280 76.790 100.340 ;
        RECT 77.405 100.280 77.695 100.325 ;
        RECT 76.470 100.140 77.695 100.280 ;
        RECT 76.470 100.080 76.790 100.140 ;
        RECT 77.405 100.095 77.695 100.140 ;
        RECT 82.450 100.080 82.770 100.340 ;
        RECT 84.290 100.080 84.610 100.340 ;
        RECT 99.970 100.255 112.810 101.065 ;
        RECT 99.990 100.195 112.800 100.255 ;
        RECT 80.625 99.940 80.915 99.985 ;
        RECT 58.960 99.800 65.660 99.940 ;
        RECT 76.560 99.800 80.915 99.940 ;
        RECT 100.990 99.835 101.430 100.195 ;
        RECT 102.570 100.085 103.730 100.195 ;
        RECT 102.570 99.835 103.010 100.085 ;
        RECT 104.160 99.835 104.600 100.195 ;
        RECT 105.750 99.835 106.190 100.195 ;
        RECT 58.960 99.755 59.250 99.800 ;
        RECT 48.410 99.645 48.730 99.660 ;
        RECT 45.205 99.460 46.430 99.600 ;
        RECT 45.205 99.415 45.495 99.460 ;
        RECT 15.725 99.260 16.015 99.305 ;
        RECT 16.915 99.260 17.205 99.305 ;
        RECT 19.435 99.260 19.725 99.305 ;
        RECT 23.000 99.260 23.290 99.305 ;
        RECT 15.725 99.120 19.725 99.260 ;
        RECT 15.725 99.075 16.015 99.120 ;
        RECT 16.915 99.075 17.205 99.120 ;
        RECT 19.435 99.075 19.725 99.120 ;
        RECT 21.820 99.120 23.290 99.260 ;
        RECT 15.330 98.920 15.620 98.965 ;
        RECT 17.430 98.920 17.720 98.965 ;
        RECT 19.000 98.920 19.290 98.965 ;
        RECT 15.330 98.780 19.290 98.920 ;
        RECT 15.330 98.735 15.620 98.780 ;
        RECT 17.430 98.735 17.720 98.780 ;
        RECT 19.000 98.735 19.290 98.780 ;
        RECT 21.820 98.640 21.960 99.120 ;
        RECT 23.000 99.075 23.290 99.120 ;
        RECT 25.410 99.060 25.730 99.320 ;
        RECT 26.330 99.260 26.650 99.320 ;
        RECT 26.880 99.260 27.020 99.415 ;
        RECT 46.110 99.400 46.430 99.460 ;
        RECT 47.045 99.415 47.335 99.645 ;
        RECT 48.380 99.415 48.730 99.645 ;
        RECT 48.410 99.400 48.730 99.415 ;
        RECT 56.230 99.400 56.550 99.660 ;
        RECT 66.350 99.600 66.670 99.660 ;
        RECT 67.285 99.600 67.575 99.645 ;
        RECT 66.350 99.460 67.575 99.600 ;
        RECT 66.350 99.400 66.670 99.460 ;
        RECT 67.285 99.415 67.575 99.460 ;
        RECT 69.110 99.600 69.430 99.660 ;
        RECT 72.345 99.600 72.635 99.645 ;
        RECT 69.110 99.460 72.635 99.600 ;
        RECT 69.110 99.400 69.430 99.460 ;
        RECT 72.345 99.415 72.635 99.460 ;
        RECT 73.725 99.600 74.015 99.645 ;
        RECT 74.170 99.600 74.490 99.660 ;
        RECT 73.725 99.460 74.490 99.600 ;
        RECT 73.725 99.415 74.015 99.460 ;
        RECT 74.170 99.400 74.490 99.460 ;
        RECT 75.550 99.400 75.870 99.660 ;
        RECT 76.010 99.600 76.330 99.660 ;
        RECT 76.560 99.645 76.700 99.800 ;
        RECT 80.625 99.755 80.915 99.800 ;
        RECT 100.130 99.785 100.360 99.815 ;
        RECT 100.520 99.785 100.750 99.835 ;
        RECT 76.485 99.600 76.775 99.645 ;
        RECT 79.245 99.600 79.535 99.645 ;
        RECT 76.010 99.460 76.775 99.600 ;
        RECT 76.010 99.400 76.330 99.460 ;
        RECT 76.485 99.415 76.775 99.460 ;
        RECT 77.020 99.460 79.535 99.600 ;
        RECT 26.330 99.120 27.020 99.260 ;
        RECT 26.330 99.060 26.650 99.120 ;
        RECT 45.665 99.075 45.955 99.305 ;
        RECT 47.925 99.260 48.215 99.305 ;
        RECT 49.115 99.260 49.405 99.305 ;
        RECT 51.635 99.260 51.925 99.305 ;
        RECT 57.625 99.260 57.915 99.305 ;
        RECT 47.925 99.120 51.925 99.260 ;
        RECT 47.925 99.075 48.215 99.120 ;
        RECT 49.115 99.075 49.405 99.120 ;
        RECT 51.635 99.075 51.925 99.120 ;
        RECT 57.240 99.120 57.915 99.260 ;
        RECT 45.740 98.920 45.880 99.075 ;
        RECT 57.240 98.980 57.380 99.120 ;
        RECT 57.625 99.075 57.915 99.120 ;
        RECT 58.505 99.260 58.795 99.305 ;
        RECT 59.695 99.260 59.985 99.305 ;
        RECT 62.215 99.260 62.505 99.305 ;
        RECT 58.505 99.120 62.505 99.260 ;
        RECT 58.505 99.075 58.795 99.120 ;
        RECT 59.695 99.075 59.985 99.120 ;
        RECT 62.215 99.075 62.505 99.120 ;
        RECT 68.190 99.260 68.510 99.320 ;
        RECT 70.490 99.260 70.810 99.320 ;
        RECT 68.190 99.120 70.810 99.260 ;
        RECT 68.190 99.060 68.510 99.120 ;
        RECT 70.490 99.060 70.810 99.120 ;
        RECT 73.265 99.260 73.555 99.305 ;
        RECT 74.630 99.260 74.950 99.320 ;
        RECT 75.640 99.260 75.780 99.400 ;
        RECT 73.265 99.120 75.780 99.260 ;
        RECT 73.265 99.075 73.555 99.120 ;
        RECT 74.630 99.060 74.950 99.120 ;
        RECT 47.030 98.920 47.350 98.980 ;
        RECT 45.740 98.780 47.350 98.920 ;
        RECT 47.030 98.720 47.350 98.780 ;
        RECT 47.530 98.920 47.820 98.965 ;
        RECT 49.630 98.920 49.920 98.965 ;
        RECT 51.200 98.920 51.490 98.965 ;
        RECT 47.530 98.780 51.490 98.920 ;
        RECT 47.530 98.735 47.820 98.780 ;
        RECT 49.630 98.735 49.920 98.780 ;
        RECT 51.200 98.735 51.490 98.780 ;
        RECT 51.720 98.780 56.460 98.920 ;
        RECT 21.730 98.380 22.050 98.640 ;
        RECT 22.190 98.380 22.510 98.640 ;
        RECT 34.150 98.580 34.470 98.640 ;
        RECT 51.720 98.580 51.860 98.780 ;
        RECT 34.150 98.440 51.860 98.580 ;
        RECT 34.150 98.380 34.470 98.440 ;
        RECT 55.770 98.380 56.090 98.640 ;
        RECT 56.320 98.580 56.460 98.780 ;
        RECT 57.150 98.720 57.470 98.980 ;
        RECT 58.110 98.920 58.400 98.965 ;
        RECT 60.210 98.920 60.500 98.965 ;
        RECT 61.780 98.920 62.070 98.965 ;
        RECT 58.110 98.780 62.070 98.920 ;
        RECT 58.110 98.735 58.400 98.780 ;
        RECT 60.210 98.735 60.500 98.780 ;
        RECT 61.780 98.735 62.070 98.780 ;
        RECT 72.790 98.720 73.110 98.980 ;
        RECT 75.550 98.720 75.870 98.980 ;
        RECT 76.470 98.920 76.790 98.980 ;
        RECT 77.020 98.920 77.160 99.460 ;
        RECT 79.245 99.415 79.535 99.460 ;
        RECT 79.690 99.400 80.010 99.660 ;
        RECT 78.310 99.260 78.630 99.320 ;
        RECT 78.785 99.260 79.075 99.305 ;
        RECT 78.310 99.120 79.075 99.260 ;
        RECT 78.310 99.060 78.630 99.120 ;
        RECT 78.785 99.075 79.075 99.120 ;
        RECT 84.750 99.060 85.070 99.320 ;
        RECT 85.210 99.060 85.530 99.320 ;
        RECT 76.470 98.780 77.160 98.920 ;
        RECT 77.390 98.920 77.710 98.980 ;
        RECT 81.530 98.920 81.850 98.980 ;
        RECT 77.390 98.780 81.850 98.920 ;
        RECT 76.470 98.720 76.790 98.780 ;
        RECT 77.390 98.720 77.710 98.780 ;
        RECT 81.530 98.720 81.850 98.780 ;
        RECT 77.850 98.580 78.170 98.640 ;
        RECT 56.320 98.440 78.170 98.580 ;
        RECT 77.850 98.380 78.170 98.440 ;
        RECT 79.230 98.380 79.550 98.640 ;
        RECT 13.380 97.760 92.040 98.240 ;
        RECT 18.510 97.560 18.830 97.620 ;
        RECT 18.985 97.560 19.275 97.605 ;
        RECT 18.510 97.420 19.275 97.560 ;
        RECT 18.510 97.360 18.830 97.420 ;
        RECT 18.985 97.375 19.275 97.420 ;
        RECT 19.430 97.360 19.750 97.620 ;
        RECT 37.830 97.560 38.150 97.620 ;
        RECT 41.525 97.560 41.815 97.605 ;
        RECT 37.830 97.420 41.815 97.560 ;
        RECT 37.830 97.360 38.150 97.420 ;
        RECT 41.525 97.375 41.815 97.420 ;
        RECT 47.965 97.560 48.255 97.605 ;
        RECT 48.410 97.560 48.730 97.620 ;
        RECT 47.965 97.420 48.730 97.560 ;
        RECT 47.965 97.375 48.255 97.420 ;
        RECT 48.410 97.360 48.730 97.420 ;
        RECT 68.205 97.560 68.495 97.605 ;
        RECT 69.110 97.560 69.430 97.620 ;
        RECT 68.205 97.420 69.430 97.560 ;
        RECT 68.205 97.375 68.495 97.420 ;
        RECT 69.110 97.360 69.430 97.420 ;
        RECT 74.630 97.360 74.950 97.620 ;
        RECT 75.090 97.560 75.410 97.620 ;
        RECT 76.025 97.560 76.315 97.605 ;
        RECT 78.310 97.560 78.630 97.620 ;
        RECT 75.090 97.420 76.315 97.560 ;
        RECT 75.090 97.360 75.410 97.420 ;
        RECT 76.025 97.375 76.315 97.420 ;
        RECT 77.480 97.420 78.630 97.560 ;
        RECT 34.650 97.220 34.940 97.265 ;
        RECT 36.750 97.220 37.040 97.265 ;
        RECT 38.320 97.220 38.610 97.265 ;
        RECT 34.650 97.080 38.610 97.220 ;
        RECT 34.650 97.035 34.940 97.080 ;
        RECT 36.750 97.035 37.040 97.080 ;
        RECT 38.320 97.035 38.610 97.080 ;
        RECT 41.065 97.220 41.355 97.265 ;
        RECT 50.710 97.220 51.030 97.280 ;
        RECT 74.170 97.220 74.490 97.280 ;
        RECT 77.480 97.220 77.620 97.420 ;
        RECT 78.310 97.360 78.630 97.420 ;
        RECT 82.925 97.560 83.215 97.605 ;
        RECT 84.750 97.560 85.070 97.620 ;
        RECT 82.925 97.420 85.070 97.560 ;
        RECT 82.925 97.375 83.215 97.420 ;
        RECT 84.750 97.360 85.070 97.420 ;
        RECT 41.065 97.080 44.500 97.220 ;
        RECT 41.065 97.035 41.355 97.080 ;
        RECT 19.905 96.880 20.195 96.925 ;
        RECT 20.365 96.880 20.655 96.925 ;
        RECT 19.905 96.740 20.655 96.880 ;
        RECT 19.905 96.695 20.195 96.740 ;
        RECT 20.365 96.695 20.655 96.740 ;
        RECT 26.790 96.880 27.110 96.940 ;
        RECT 44.360 96.925 44.500 97.080 ;
        RECT 50.710 97.080 54.620 97.220 ;
        RECT 50.710 97.020 51.030 97.080 ;
        RECT 34.165 96.880 34.455 96.925 ;
        RECT 26.790 96.740 34.455 96.880 ;
        RECT 26.790 96.680 27.110 96.740 ;
        RECT 34.165 96.695 34.455 96.740 ;
        RECT 35.045 96.880 35.335 96.925 ;
        RECT 36.235 96.880 36.525 96.925 ;
        RECT 38.755 96.880 39.045 96.925 ;
        RECT 35.045 96.740 39.045 96.880 ;
        RECT 35.045 96.695 35.335 96.740 ;
        RECT 36.235 96.695 36.525 96.740 ;
        RECT 38.755 96.695 39.045 96.740 ;
        RECT 44.285 96.880 44.575 96.925 ;
        RECT 45.190 96.880 45.510 96.940 ;
        RECT 44.285 96.740 45.510 96.880 ;
        RECT 44.285 96.695 44.575 96.740 ;
        RECT 45.190 96.680 45.510 96.740 ;
        RECT 51.170 96.680 51.490 96.940 ;
        RECT 18.525 96.355 18.815 96.585 ;
        RECT 21.730 96.540 22.050 96.600 ;
        RECT 23.125 96.540 23.415 96.585 ;
        RECT 21.730 96.400 23.415 96.540 ;
        RECT 18.600 96.200 18.740 96.355 ;
        RECT 21.730 96.340 22.050 96.400 ;
        RECT 23.125 96.355 23.415 96.400 ;
        RECT 50.265 96.540 50.555 96.585 ;
        RECT 52.090 96.540 52.410 96.600 ;
        RECT 54.480 96.585 54.620 97.080 ;
        RECT 74.170 97.080 77.620 97.220 ;
        RECT 77.850 97.220 78.170 97.280 ;
        RECT 77.850 97.080 80.840 97.220 ;
        RECT 74.170 97.020 74.490 97.080 ;
        RECT 77.850 97.020 78.170 97.080 ;
        RECT 55.770 96.880 56.090 96.940 ;
        RECT 58.530 96.880 58.850 96.940 ;
        RECT 55.770 96.740 58.850 96.880 ;
        RECT 55.770 96.680 56.090 96.740 ;
        RECT 58.530 96.680 58.850 96.740 ;
        RECT 65.430 96.880 65.750 96.940 ;
        RECT 65.430 96.740 69.800 96.880 ;
        RECT 65.430 96.680 65.750 96.740 ;
        RECT 69.660 96.600 69.800 96.740 ;
        RECT 80.150 96.680 80.470 96.940 ;
        RECT 80.700 96.925 80.840 97.080 ;
        RECT 80.625 96.695 80.915 96.925 ;
        RECT 50.265 96.400 52.410 96.540 ;
        RECT 50.265 96.355 50.555 96.400 ;
        RECT 52.090 96.340 52.410 96.400 ;
        RECT 54.405 96.355 54.695 96.585 ;
        RECT 61.750 96.340 62.070 96.600 ;
        RECT 64.985 96.540 65.275 96.585 ;
        RECT 68.190 96.540 68.510 96.600 ;
        RECT 64.985 96.400 68.510 96.540 ;
        RECT 64.985 96.355 65.275 96.400 ;
        RECT 68.190 96.340 68.510 96.400 ;
        RECT 69.570 96.340 69.890 96.600 ;
        RECT 70.490 96.340 70.810 96.600 ;
        RECT 72.790 96.540 73.110 96.600 ;
        RECT 74.185 96.540 74.475 96.585 ;
        RECT 72.790 96.400 74.475 96.540 ;
        RECT 72.790 96.340 73.110 96.400 ;
        RECT 74.185 96.355 74.475 96.400 ;
        RECT 74.630 96.340 74.950 96.600 ;
        RECT 22.650 96.200 22.970 96.260 ;
        RECT 25.410 96.200 25.730 96.260 ;
        RECT 35.530 96.245 35.850 96.260 ;
        RECT 18.600 96.060 25.730 96.200 ;
        RECT 22.650 96.000 22.970 96.060 ;
        RECT 25.410 96.000 25.730 96.060 ;
        RECT 35.500 96.015 35.850 96.245 ;
        RECT 49.805 96.200 50.095 96.245 ;
        RECT 54.865 96.200 55.155 96.245 ;
        RECT 55.310 96.200 55.630 96.260 ;
        RECT 49.805 96.060 52.780 96.200 ;
        RECT 49.805 96.015 50.095 96.060 ;
        RECT 35.530 96.000 35.850 96.015 ;
        RECT 52.640 95.905 52.780 96.060 ;
        RECT 54.865 96.060 55.630 96.200 ;
        RECT 54.865 96.015 55.155 96.060 ;
        RECT 55.310 96.000 55.630 96.060 ;
        RECT 68.650 96.200 68.970 96.260 ;
        RECT 69.125 96.200 69.415 96.245 ;
        RECT 72.330 96.200 72.650 96.260 ;
        RECT 68.650 96.060 69.415 96.200 ;
        RECT 68.650 96.000 68.970 96.060 ;
        RECT 69.125 96.015 69.415 96.060 ;
        RECT 69.660 96.060 72.650 96.200 ;
        RECT 52.565 95.675 52.855 95.905 ;
        RECT 67.270 95.660 67.590 95.920 ;
        RECT 68.125 95.860 68.415 95.905 ;
        RECT 69.660 95.860 69.800 96.060 ;
        RECT 72.330 96.000 72.650 96.060 ;
        RECT 68.125 95.720 69.800 95.860 ;
        RECT 70.030 95.860 70.350 95.920 ;
        RECT 76.470 95.860 76.790 95.920 ;
        RECT 70.030 95.720 76.790 95.860 ;
        RECT 68.125 95.675 68.415 95.720 ;
        RECT 70.030 95.660 70.350 95.720 ;
        RECT 76.470 95.660 76.790 95.720 ;
        RECT 81.070 95.660 81.390 95.920 ;
        RECT 13.380 95.040 92.040 95.520 ;
        RECT 22.665 94.840 22.955 94.885 ;
        RECT 23.110 94.840 23.430 94.900 ;
        RECT 26.330 94.840 26.650 94.900 ;
        RECT 22.665 94.700 26.650 94.840 ;
        RECT 22.665 94.655 22.955 94.700 ;
        RECT 23.110 94.640 23.430 94.700 ;
        RECT 26.330 94.640 26.650 94.700 ;
        RECT 33.245 94.840 33.535 94.885 ;
        RECT 34.150 94.840 34.470 94.900 ;
        RECT 33.245 94.700 34.470 94.840 ;
        RECT 33.245 94.655 33.535 94.700 ;
        RECT 34.150 94.640 34.470 94.700 ;
        RECT 35.085 94.840 35.375 94.885 ;
        RECT 35.530 94.840 35.850 94.900 ;
        RECT 45.190 94.885 45.510 94.900 ;
        RECT 35.085 94.700 35.850 94.840 ;
        RECT 35.085 94.655 35.375 94.700 ;
        RECT 35.530 94.640 35.850 94.700 ;
        RECT 36.925 94.840 37.215 94.885 ;
        RECT 40.145 94.840 40.435 94.885 ;
        RECT 36.925 94.700 40.435 94.840 ;
        RECT 36.925 94.655 37.215 94.700 ;
        RECT 40.145 94.655 40.435 94.700 ;
        RECT 45.190 94.655 45.575 94.885 ;
        RECT 55.325 94.840 55.615 94.885 ;
        RECT 61.750 94.840 62.070 94.900 ;
        RECT 55.325 94.700 62.070 94.840 ;
        RECT 55.325 94.655 55.615 94.700 ;
        RECT 45.190 94.640 45.510 94.655 ;
        RECT 18.510 94.500 18.830 94.560 ;
        RECT 37.385 94.500 37.675 94.545 ;
        RECT 37.830 94.500 38.150 94.560 ;
        RECT 18.510 94.360 21.040 94.500 ;
        RECT 18.510 94.300 18.830 94.360 ;
        RECT 20.900 94.205 21.040 94.360 ;
        RECT 37.385 94.360 38.150 94.500 ;
        RECT 37.385 94.315 37.675 94.360 ;
        RECT 37.830 94.300 38.150 94.360 ;
        RECT 44.270 94.300 44.590 94.560 ;
        RECT 18.065 94.160 18.355 94.205 ;
        RECT 18.065 94.020 20.580 94.160 ;
        RECT 18.065 93.975 18.355 94.020 ;
        RECT 18.525 93.635 18.815 93.865 ;
        RECT 18.600 93.480 18.740 93.635 ;
        RECT 18.970 93.620 19.290 93.880 ;
        RECT 20.440 93.820 20.580 94.020 ;
        RECT 20.825 93.975 21.115 94.205 ;
        RECT 21.745 94.160 22.035 94.205 ;
        RECT 22.650 94.160 22.970 94.220 ;
        RECT 21.745 94.020 22.970 94.160 ;
        RECT 21.745 93.975 22.035 94.020 ;
        RECT 22.650 93.960 22.970 94.020 ;
        RECT 26.345 94.160 26.635 94.205 ;
        RECT 26.790 94.160 27.110 94.220 ;
        RECT 27.710 94.205 28.030 94.220 ;
        RECT 26.345 94.020 27.110 94.160 ;
        RECT 26.345 93.975 26.635 94.020 ;
        RECT 26.790 93.960 27.110 94.020 ;
        RECT 27.680 93.975 28.030 94.205 ;
        RECT 27.710 93.960 28.030 93.975 ;
        RECT 41.970 93.960 42.290 94.220 ;
        RECT 42.445 94.160 42.735 94.205 ;
        RECT 55.400 94.160 55.540 94.655 ;
        RECT 61.750 94.640 62.070 94.700 ;
        RECT 65.445 94.655 65.735 94.885 ;
        RECT 76.025 94.840 76.315 94.885 ;
        RECT 81.070 94.840 81.390 94.900 ;
        RECT 76.025 94.700 81.390 94.840 ;
        RECT 76.025 94.655 76.315 94.700 ;
        RECT 61.000 94.500 61.290 94.545 ;
        RECT 65.520 94.500 65.660 94.655 ;
        RECT 81.070 94.640 81.390 94.700 ;
        RECT 82.465 94.840 82.755 94.885 ;
        RECT 82.910 94.840 83.230 94.900 ;
        RECT 82.465 94.700 83.230 94.840 ;
        RECT 82.465 94.655 82.755 94.700 ;
        RECT 82.910 94.640 83.230 94.700 ;
        RECT 61.000 94.360 65.660 94.500 ;
        RECT 61.000 94.315 61.290 94.360 ;
        RECT 66.810 94.300 67.130 94.560 ;
        RECT 67.285 94.500 67.575 94.545 ;
        RECT 69.125 94.500 69.415 94.545 ;
        RECT 67.285 94.360 69.415 94.500 ;
        RECT 67.285 94.315 67.575 94.360 ;
        RECT 69.125 94.315 69.415 94.360 ;
        RECT 71.040 94.360 81.300 94.500 ;
        RECT 42.445 94.020 55.540 94.160 ;
        RECT 56.320 94.020 62.900 94.160 ;
        RECT 42.445 93.975 42.735 94.020 ;
        RECT 21.270 93.820 21.590 93.880 ;
        RECT 25.410 93.820 25.730 93.880 ;
        RECT 20.440 93.680 25.730 93.820 ;
        RECT 21.270 93.620 21.590 93.680 ;
        RECT 25.410 93.620 25.730 93.680 ;
        RECT 27.225 93.820 27.515 93.865 ;
        RECT 28.415 93.820 28.705 93.865 ;
        RECT 30.935 93.820 31.225 93.865 ;
        RECT 27.225 93.680 31.225 93.820 ;
        RECT 27.225 93.635 27.515 93.680 ;
        RECT 28.415 93.635 28.705 93.680 ;
        RECT 30.935 93.635 31.225 93.680 ;
        RECT 38.290 93.620 38.610 93.880 ;
        RECT 43.365 93.820 43.655 93.865 ;
        RECT 55.770 93.820 56.090 93.880 ;
        RECT 43.365 93.680 56.090 93.820 ;
        RECT 43.365 93.635 43.655 93.680 ;
        RECT 55.770 93.620 56.090 93.680 ;
        RECT 22.650 93.480 22.970 93.540 ;
        RECT 24.950 93.480 25.270 93.540 ;
        RECT 26.830 93.480 27.120 93.525 ;
        RECT 28.930 93.480 29.220 93.525 ;
        RECT 30.500 93.480 30.790 93.525 ;
        RECT 56.320 93.480 56.460 94.020 ;
        RECT 57.635 93.820 57.925 93.865 ;
        RECT 60.155 93.820 60.445 93.865 ;
        RECT 61.345 93.820 61.635 93.865 ;
        RECT 57.635 93.680 61.635 93.820 ;
        RECT 57.635 93.635 57.925 93.680 ;
        RECT 60.155 93.635 60.445 93.680 ;
        RECT 61.345 93.635 61.635 93.680 ;
        RECT 62.225 93.635 62.515 93.865 ;
        RECT 18.600 93.340 26.560 93.480 ;
        RECT 22.650 93.280 22.970 93.340 ;
        RECT 24.950 93.280 25.270 93.340 ;
        RECT 16.210 92.940 16.530 93.200 ;
        RECT 21.730 92.940 22.050 93.200 ;
        RECT 26.420 93.140 26.560 93.340 ;
        RECT 26.830 93.340 30.790 93.480 ;
        RECT 26.830 93.295 27.120 93.340 ;
        RECT 28.930 93.295 29.220 93.340 ;
        RECT 30.500 93.295 30.790 93.340 ;
        RECT 31.480 93.340 56.460 93.480 ;
        RECT 58.070 93.480 58.360 93.525 ;
        RECT 59.640 93.480 59.930 93.525 ;
        RECT 61.740 93.480 62.030 93.525 ;
        RECT 58.070 93.340 62.030 93.480 ;
        RECT 31.480 93.140 31.620 93.340 ;
        RECT 58.070 93.295 58.360 93.340 ;
        RECT 59.640 93.295 59.930 93.340 ;
        RECT 61.740 93.295 62.030 93.340 ;
        RECT 26.420 93.000 31.620 93.140 ;
        RECT 45.190 92.940 45.510 93.200 ;
        RECT 46.125 93.140 46.415 93.185 ;
        RECT 48.410 93.140 48.730 93.200 ;
        RECT 46.125 93.000 48.730 93.140 ;
        RECT 46.125 92.955 46.415 93.000 ;
        RECT 48.410 92.940 48.730 93.000 ;
        RECT 57.150 93.140 57.470 93.200 ;
        RECT 62.300 93.140 62.440 93.635 ;
        RECT 62.760 93.480 62.900 94.020 ;
        RECT 66.365 93.975 66.655 94.205 ;
        RECT 66.440 93.820 66.580 93.975 ;
        RECT 68.190 93.960 68.510 94.220 ;
        RECT 70.030 93.960 70.350 94.220 ;
        RECT 70.490 93.960 70.810 94.220 ;
        RECT 69.110 93.820 69.430 93.880 ;
        RECT 66.440 93.680 69.430 93.820 ;
        RECT 69.110 93.620 69.430 93.680 ;
        RECT 71.040 93.480 71.180 94.360 ;
        RECT 71.425 93.975 71.715 94.205 ;
        RECT 71.500 93.820 71.640 93.975 ;
        RECT 71.870 93.960 72.190 94.220 ;
        RECT 72.790 94.160 73.110 94.220 ;
        RECT 74.185 94.160 74.475 94.205 ;
        RECT 72.790 94.020 74.475 94.160 ;
        RECT 72.790 93.960 73.110 94.020 ;
        RECT 74.185 93.975 74.475 94.020 ;
        RECT 76.470 93.960 76.790 94.220 ;
        RECT 77.405 94.160 77.695 94.205 ;
        RECT 77.850 94.160 78.170 94.220 ;
        RECT 77.405 94.020 78.170 94.160 ;
        RECT 77.405 93.975 77.695 94.020 ;
        RECT 77.850 93.960 78.170 94.020 ;
        RECT 78.325 94.160 78.615 94.205 ;
        RECT 79.705 94.160 79.995 94.205 ;
        RECT 78.325 94.020 79.995 94.160 ;
        RECT 78.325 93.975 78.615 94.020 ;
        RECT 79.705 93.975 79.995 94.020 ;
        RECT 80.150 94.160 80.470 94.220 ;
        RECT 81.160 94.205 81.300 94.360 ;
        RECT 80.625 94.160 80.915 94.205 ;
        RECT 80.150 94.020 80.915 94.160 ;
        RECT 80.150 93.960 80.470 94.020 ;
        RECT 80.625 93.975 80.915 94.020 ;
        RECT 81.085 93.975 81.375 94.205 ;
        RECT 81.545 93.975 81.835 94.205 ;
        RECT 73.250 93.820 73.570 93.880 ;
        RECT 71.500 93.680 73.570 93.820 ;
        RECT 73.250 93.620 73.570 93.680 ;
        RECT 74.645 93.635 74.935 93.865 ;
        RECT 76.930 93.820 77.250 93.880 ;
        RECT 79.230 93.820 79.550 93.880 ;
        RECT 81.620 93.820 81.760 93.975 ;
        RECT 76.930 93.680 81.760 93.820 ;
        RECT 100.130 93.895 100.750 99.785 ;
        RECT 62.760 93.340 71.180 93.480 ;
        RECT 74.720 93.480 74.860 93.635 ;
        RECT 76.930 93.620 77.250 93.680 ;
        RECT 79.230 93.620 79.550 93.680 ;
        RECT 100.130 93.615 100.370 93.895 ;
        RECT 100.520 93.835 100.750 93.895 ;
        RECT 100.960 93.895 101.430 99.835 ;
        RECT 102.100 99.765 102.330 99.835 ;
        RECT 101.800 93.915 102.330 99.765 ;
        RECT 101.800 93.895 101.960 93.915 ;
        RECT 100.960 93.835 101.190 93.895 ;
        RECT 101.810 93.655 101.960 93.895 ;
        RECT 102.100 93.835 102.330 93.915 ;
        RECT 102.540 93.915 103.010 99.835 ;
        RECT 103.680 99.765 103.910 99.835 ;
        RECT 103.310 95.175 103.920 99.765 ;
        RECT 102.540 93.835 102.770 93.915 ;
        RECT 103.290 93.885 103.920 95.175 ;
        RECT 104.120 93.925 104.600 99.835 ;
        RECT 105.260 99.785 105.490 99.835 ;
        RECT 77.850 93.480 78.170 93.540 ;
        RECT 74.720 93.340 78.170 93.480 ;
        RECT 77.850 93.280 78.170 93.340 ;
        RECT 57.150 93.000 62.440 93.140 ;
        RECT 67.270 93.140 67.590 93.200 ;
        RECT 69.570 93.140 69.890 93.200 ;
        RECT 71.870 93.140 72.190 93.200 ;
        RECT 67.270 93.000 72.190 93.140 ;
        RECT 57.150 92.940 57.470 93.000 ;
        RECT 67.270 92.940 67.590 93.000 ;
        RECT 69.570 92.940 69.890 93.000 ;
        RECT 71.870 92.940 72.190 93.000 ;
        RECT 75.105 93.140 75.395 93.185 ;
        RECT 78.770 93.140 79.090 93.200 ;
        RECT 75.105 93.000 79.090 93.140 ;
        RECT 75.105 92.955 75.395 93.000 ;
        RECT 78.770 92.940 79.090 93.000 ;
        RECT 13.380 92.320 92.040 92.800 ;
        RECT 21.745 92.120 22.035 92.165 ;
        RECT 22.650 92.120 22.970 92.180 ;
        RECT 21.745 91.980 22.970 92.120 ;
        RECT 21.745 91.935 22.035 91.980 ;
        RECT 22.650 91.920 22.970 91.980 ;
        RECT 24.490 91.920 24.810 92.180 ;
        RECT 25.425 92.120 25.715 92.165 ;
        RECT 25.870 92.120 26.190 92.180 ;
        RECT 25.425 91.980 26.190 92.120 ;
        RECT 25.425 91.935 25.715 91.980 ;
        RECT 25.870 91.920 26.190 91.980 ;
        RECT 27.265 92.120 27.555 92.165 ;
        RECT 27.710 92.120 28.030 92.180 ;
        RECT 27.265 91.980 28.030 92.120 ;
        RECT 27.265 91.935 27.555 91.980 ;
        RECT 27.710 91.920 28.030 91.980 ;
        RECT 48.885 92.120 49.175 92.165 ;
        RECT 49.330 92.120 49.650 92.180 ;
        RECT 48.885 91.980 49.650 92.120 ;
        RECT 48.885 91.935 49.175 91.980 ;
        RECT 49.330 91.920 49.650 91.980 ;
        RECT 72.345 91.935 72.635 92.165 ;
        RECT 72.790 92.120 73.110 92.180 ;
        RECT 73.265 92.120 73.555 92.165 ;
        RECT 72.790 91.980 73.555 92.120 ;
        RECT 15.330 91.780 15.620 91.825 ;
        RECT 17.430 91.780 17.720 91.825 ;
        RECT 19.000 91.780 19.290 91.825 ;
        RECT 15.330 91.640 19.290 91.780 ;
        RECT 15.330 91.595 15.620 91.640 ;
        RECT 17.430 91.595 17.720 91.640 ;
        RECT 19.000 91.595 19.290 91.640 ;
        RECT 14.830 91.240 15.150 91.500 ;
        RECT 15.725 91.440 16.015 91.485 ;
        RECT 16.915 91.440 17.205 91.485 ;
        RECT 19.435 91.440 19.725 91.485 ;
        RECT 23.110 91.440 23.430 91.500 ;
        RECT 15.725 91.300 19.725 91.440 ;
        RECT 15.725 91.255 16.015 91.300 ;
        RECT 16.915 91.255 17.205 91.300 ;
        RECT 19.435 91.255 19.725 91.300 ;
        RECT 22.280 91.300 23.430 91.440 ;
        RECT 25.960 91.440 26.100 91.920 ;
        RECT 30.025 91.440 30.315 91.485 ;
        RECT 25.960 91.300 30.315 91.440 ;
        RECT 14.920 91.100 15.060 91.240 ;
        RECT 21.730 91.100 22.050 91.160 ;
        RECT 14.920 90.960 22.050 91.100 ;
        RECT 21.730 90.900 22.050 90.960 ;
        RECT 16.210 90.805 16.530 90.820 ;
        RECT 16.180 90.760 16.530 90.805 ;
        RECT 16.015 90.620 16.530 90.760 ;
        RECT 16.180 90.575 16.530 90.620 ;
        RECT 16.210 90.560 16.530 90.575 ;
        RECT 18.970 90.760 19.290 90.820 ;
        RECT 22.280 90.760 22.420 91.300 ;
        RECT 23.110 91.240 23.430 91.300 ;
        RECT 30.025 91.255 30.315 91.300 ;
        RECT 38.750 91.440 39.070 91.500 ;
        RECT 41.065 91.440 41.355 91.485 ;
        RECT 41.970 91.440 42.290 91.500 ;
        RECT 68.650 91.440 68.970 91.500 ;
        RECT 72.420 91.440 72.560 91.935 ;
        RECT 72.790 91.920 73.110 91.980 ;
        RECT 73.265 91.935 73.555 91.980 ;
        RECT 38.750 91.300 42.290 91.440 ;
        RECT 38.750 91.240 39.070 91.300 ;
        RECT 41.065 91.255 41.355 91.300 ;
        RECT 41.970 91.240 42.290 91.300 ;
        RECT 68.280 91.300 72.560 91.440 ;
        RECT 25.410 91.100 25.730 91.160 ;
        RECT 27.710 91.100 28.030 91.160 ;
        RECT 29.565 91.100 29.855 91.145 ;
        RECT 25.410 90.960 29.855 91.100 ;
        RECT 25.410 90.900 25.730 90.960 ;
        RECT 27.710 90.900 28.030 90.960 ;
        RECT 29.565 90.915 29.855 90.960 ;
        RECT 47.965 90.915 48.255 91.145 ;
        RECT 48.410 91.100 48.730 91.160 ;
        RECT 68.280 91.145 68.420 91.300 ;
        RECT 68.650 91.240 68.970 91.300 ;
        RECT 80.150 91.240 80.470 91.500 ;
        RECT 100.130 91.185 100.510 93.615 ;
        RECT 100.710 93.605 101.000 93.630 ;
        RECT 100.700 92.905 101.020 93.605 ;
        RECT 100.650 91.875 101.650 92.905 ;
        RECT 100.700 91.185 101.020 91.875 ;
        RECT 48.885 91.100 49.175 91.145 ;
        RECT 48.410 90.960 49.175 91.100 ;
        RECT 18.970 90.620 22.420 90.760 ;
        RECT 23.110 90.760 23.430 90.820 ;
        RECT 23.585 90.760 23.875 90.805 ;
        RECT 23.110 90.620 23.875 90.760 ;
        RECT 18.970 90.560 19.290 90.620 ;
        RECT 23.110 90.560 23.430 90.620 ;
        RECT 23.585 90.575 23.875 90.620 ;
        RECT 29.105 90.760 29.395 90.805 ;
        RECT 34.150 90.760 34.470 90.820 ;
        RECT 29.105 90.620 34.470 90.760 ;
        RECT 29.105 90.575 29.395 90.620 ;
        RECT 34.150 90.560 34.470 90.620 ;
        RECT 46.585 90.760 46.875 90.805 ;
        RECT 47.030 90.760 47.350 90.820 ;
        RECT 46.585 90.620 47.350 90.760 ;
        RECT 48.040 90.760 48.180 90.915 ;
        RECT 48.410 90.900 48.730 90.960 ;
        RECT 48.885 90.915 49.175 90.960 ;
        RECT 68.205 90.915 68.495 91.145 ;
        RECT 69.125 91.100 69.415 91.145 ;
        RECT 72.790 91.100 73.110 91.160 ;
        RECT 69.125 90.960 73.110 91.100 ;
        RECT 69.125 90.915 69.415 90.960 ;
        RECT 72.500 90.900 73.110 90.960 ;
        RECT 78.770 90.900 79.090 91.160 ;
        RECT 79.230 90.900 79.550 91.160 ;
        RECT 81.545 91.100 81.835 91.145 ;
        RECT 81.990 91.100 82.310 91.160 ;
        RECT 81.545 90.960 82.310 91.100 ;
        RECT 81.545 90.915 81.835 90.960 ;
        RECT 81.990 90.900 82.310 90.960 ;
        RECT 89.810 90.900 90.130 91.160 ;
        RECT 52.550 90.760 52.870 90.820 ;
        RECT 48.040 90.620 52.870 90.760 ;
        RECT 46.585 90.575 46.875 90.620 ;
        RECT 47.030 90.560 47.350 90.620 ;
        RECT 52.550 90.560 52.870 90.620 ;
        RECT 67.270 90.560 67.590 90.820 ;
        RECT 70.490 90.760 70.810 90.820 ;
        RECT 71.425 90.760 71.715 90.805 ;
        RECT 72.500 90.790 72.865 90.900 ;
        RECT 100.130 90.875 100.370 91.185 ;
        RECT 100.720 91.145 101.020 91.185 ;
        RECT 100.720 91.135 101.010 91.145 ;
        RECT 101.810 91.125 102.010 93.655 ;
        RECT 102.290 93.625 102.580 93.630 ;
        RECT 102.280 92.955 102.620 93.625 ;
        RECT 102.150 91.925 103.150 92.955 ;
        RECT 102.280 91.155 102.620 91.925 ;
        RECT 102.300 91.135 102.590 91.155 ;
        RECT 100.530 90.875 100.760 90.975 ;
        RECT 100.130 90.865 100.760 90.875 ;
        RECT 70.490 90.620 71.715 90.760 ;
        RECT 72.575 90.745 72.865 90.790 ;
        RECT 70.490 90.560 70.810 90.620 ;
        RECT 71.425 90.575 71.715 90.620 ;
        RECT 22.190 90.420 22.510 90.480 ;
        RECT 24.585 90.420 24.875 90.465 ;
        RECT 22.190 90.280 24.875 90.420 ;
        RECT 22.190 90.220 22.510 90.280 ;
        RECT 24.585 90.235 24.875 90.280 ;
        RECT 41.510 90.420 41.830 90.480 ;
        RECT 43.825 90.420 44.115 90.465 ;
        RECT 41.510 90.280 44.115 90.420 ;
        RECT 41.510 90.220 41.830 90.280 ;
        RECT 43.825 90.235 44.115 90.280 ;
        RECT 49.790 90.220 50.110 90.480 ;
        RECT 70.030 90.420 70.350 90.480 ;
        RECT 77.850 90.420 78.170 90.480 ;
        RECT 81.085 90.420 81.375 90.465 ;
        RECT 70.030 90.280 81.375 90.420 ;
        RECT 70.030 90.220 70.350 90.280 ;
        RECT 77.850 90.220 78.170 90.280 ;
        RECT 81.085 90.235 81.375 90.280 ;
        RECT 87.050 90.220 87.370 90.480 ;
        RECT 13.380 89.600 92.040 90.080 ;
        RECT 17.145 89.400 17.435 89.445 ;
        RECT 18.510 89.400 18.830 89.460 ;
        RECT 24.490 89.400 24.810 89.460 ;
        RECT 17.145 89.260 18.830 89.400 ;
        RECT 17.145 89.215 17.435 89.260 ;
        RECT 18.510 89.200 18.830 89.260 ;
        RECT 19.060 89.260 24.810 89.400 ;
        RECT 19.060 89.060 19.200 89.260 ;
        RECT 24.490 89.200 24.810 89.260 ;
        RECT 26.330 89.400 26.650 89.460 ;
        RECT 26.330 89.260 27.020 89.400 ;
        RECT 26.330 89.200 26.650 89.260 ;
        RECT 21.730 89.060 22.050 89.120 ;
        RECT 26.880 89.105 27.020 89.260 ;
        RECT 38.750 89.200 39.070 89.460 ;
        RECT 39.685 89.215 39.975 89.445 ;
        RECT 18.140 88.920 19.200 89.060 ;
        RECT 19.520 88.920 26.560 89.060 ;
        RECT 18.140 87.745 18.280 88.920 ;
        RECT 18.970 88.520 19.290 88.780 ;
        RECT 19.520 88.765 19.660 88.920 ;
        RECT 21.730 88.860 22.050 88.920 ;
        RECT 19.445 88.535 19.735 88.765 ;
        RECT 20.780 88.720 21.070 88.765 ;
        RECT 22.190 88.720 22.510 88.780 ;
        RECT 20.780 88.580 22.510 88.720 ;
        RECT 26.420 88.720 26.560 88.920 ;
        RECT 26.805 88.875 27.095 89.105 ;
        RECT 27.250 89.060 27.570 89.120 ;
        RECT 27.805 89.060 28.095 89.105 ;
        RECT 27.250 88.920 28.095 89.060 ;
        RECT 27.250 88.860 27.570 88.920 ;
        RECT 27.805 88.875 28.095 88.920 ;
        RECT 33.200 89.060 33.490 89.105 ;
        RECT 39.760 89.060 39.900 89.215 ;
        RECT 41.510 89.200 41.830 89.460 ;
        RECT 42.890 89.400 43.210 89.460 ;
        RECT 45.665 89.400 45.955 89.445 ;
        RECT 42.890 89.260 45.955 89.400 ;
        RECT 42.890 89.200 43.210 89.260 ;
        RECT 45.665 89.215 45.955 89.260 ;
        RECT 49.330 89.200 49.650 89.460 ;
        RECT 52.090 89.400 52.410 89.460 ;
        RECT 49.880 89.260 52.410 89.400 ;
        RECT 49.880 89.060 50.020 89.260 ;
        RECT 52.090 89.200 52.410 89.260 ;
        RECT 52.550 89.200 52.870 89.460 ;
        RECT 64.065 89.400 64.355 89.445 ;
        RECT 68.650 89.400 68.970 89.460 ;
        RECT 64.065 89.260 68.970 89.400 ;
        RECT 64.065 89.215 64.355 89.260 ;
        RECT 68.650 89.200 68.970 89.260 ;
        RECT 72.330 89.200 72.650 89.460 ;
        RECT 74.185 89.400 74.475 89.445 ;
        RECT 74.630 89.400 74.950 89.460 ;
        RECT 74.185 89.260 74.950 89.400 ;
        RECT 74.185 89.215 74.475 89.260 ;
        RECT 74.630 89.200 74.950 89.260 ;
        RECT 87.510 89.400 87.830 89.460 ;
        RECT 88.445 89.400 88.735 89.445 ;
        RECT 89.810 89.400 90.130 89.460 ;
        RECT 87.510 89.260 90.130 89.400 ;
        RECT 87.510 89.200 87.830 89.260 ;
        RECT 88.445 89.215 88.735 89.260 ;
        RECT 89.810 89.200 90.130 89.260 ;
        RECT 33.200 88.920 39.900 89.060 ;
        RECT 47.120 88.920 50.020 89.060 ;
        RECT 50.265 89.060 50.555 89.105 ;
        RECT 56.690 89.060 57.010 89.120 ;
        RECT 50.265 88.920 57.010 89.060 ;
        RECT 33.200 88.875 33.490 88.920 ;
        RECT 44.270 88.720 44.590 88.780 ;
        RECT 47.120 88.765 47.260 88.920 ;
        RECT 50.265 88.875 50.555 88.920 ;
        RECT 56.690 88.860 57.010 88.920 ;
        RECT 67.285 89.060 67.575 89.105 ;
        RECT 69.570 89.060 69.890 89.120 ;
        RECT 67.285 88.920 73.480 89.060 ;
        RECT 67.285 88.875 67.575 88.920 ;
        RECT 69.570 88.860 69.890 88.920 ;
        RECT 47.045 88.720 47.335 88.765 ;
        RECT 26.420 88.580 27.020 88.720 ;
        RECT 20.780 88.535 21.070 88.580 ;
        RECT 22.190 88.520 22.510 88.580 ;
        RECT 26.880 88.440 27.020 88.580 ;
        RECT 44.270 88.580 47.335 88.720 ;
        RECT 44.270 88.520 44.590 88.580 ;
        RECT 47.045 88.535 47.335 88.580 ;
        RECT 47.505 88.535 47.795 88.765 ;
        RECT 18.525 88.195 18.815 88.425 ;
        RECT 20.325 88.380 20.615 88.425 ;
        RECT 21.515 88.380 21.805 88.425 ;
        RECT 24.035 88.380 24.325 88.425 ;
        RECT 20.325 88.240 24.325 88.380 ;
        RECT 20.325 88.195 20.615 88.240 ;
        RECT 21.515 88.195 21.805 88.240 ;
        RECT 24.035 88.195 24.325 88.240 ;
        RECT 26.790 88.380 27.110 88.440 ;
        RECT 31.865 88.380 32.155 88.425 ;
        RECT 26.790 88.240 32.155 88.380 ;
        RECT 18.065 87.515 18.355 87.745 ;
        RECT 18.600 87.700 18.740 88.195 ;
        RECT 26.790 88.180 27.110 88.240 ;
        RECT 31.865 88.195 32.155 88.240 ;
        RECT 32.745 88.380 33.035 88.425 ;
        RECT 33.935 88.380 34.225 88.425 ;
        RECT 36.455 88.380 36.745 88.425 ;
        RECT 32.745 88.240 36.745 88.380 ;
        RECT 32.745 88.195 33.035 88.240 ;
        RECT 33.935 88.195 34.225 88.240 ;
        RECT 36.455 88.195 36.745 88.240 ;
        RECT 36.910 88.380 37.230 88.440 ;
        RECT 41.985 88.380 42.275 88.425 ;
        RECT 36.910 88.240 42.275 88.380 ;
        RECT 36.910 88.180 37.230 88.240 ;
        RECT 41.985 88.195 42.275 88.240 ;
        RECT 42.905 88.195 43.195 88.425 ;
        RECT 47.580 88.380 47.720 88.535 ;
        RECT 47.950 88.520 48.270 88.780 ;
        RECT 48.885 88.720 49.175 88.765 ;
        RECT 49.790 88.720 50.110 88.780 ;
        RECT 48.885 88.580 50.110 88.720 ;
        RECT 48.885 88.535 49.175 88.580 ;
        RECT 49.790 88.520 50.110 88.580 ;
        RECT 52.090 88.520 52.410 88.780 ;
        RECT 58.500 88.720 58.790 88.765 ;
        RECT 65.445 88.720 65.735 88.765 ;
        RECT 58.500 88.580 65.735 88.720 ;
        RECT 58.500 88.535 58.790 88.580 ;
        RECT 65.445 88.535 65.735 88.580 ;
        RECT 66.350 88.520 66.670 88.780 ;
        RECT 66.810 88.520 67.130 88.780 ;
        RECT 67.875 88.720 68.165 88.765 ;
        RECT 67.360 88.580 68.165 88.720 ;
        RECT 54.865 88.380 55.155 88.425 ;
        RECT 47.580 88.240 55.155 88.380 ;
        RECT 19.930 88.040 20.220 88.085 ;
        RECT 22.030 88.040 22.320 88.085 ;
        RECT 23.600 88.040 23.890 88.085 ;
        RECT 19.930 87.900 23.890 88.040 ;
        RECT 19.930 87.855 20.220 87.900 ;
        RECT 22.030 87.855 22.320 87.900 ;
        RECT 23.600 87.855 23.890 87.900 ;
        RECT 24.490 88.040 24.810 88.100 ;
        RECT 32.350 88.040 32.640 88.085 ;
        RECT 34.450 88.040 34.740 88.085 ;
        RECT 36.020 88.040 36.310 88.085 ;
        RECT 24.490 87.900 27.940 88.040 ;
        RECT 24.490 87.840 24.810 87.900 ;
        RECT 23.110 87.700 23.430 87.760 ;
        RECT 26.330 87.700 26.650 87.760 ;
        RECT 27.800 87.745 27.940 87.900 ;
        RECT 32.350 87.900 36.310 88.040 ;
        RECT 42.980 88.040 43.120 88.195 ;
        RECT 49.330 88.040 49.650 88.100 ;
        RECT 42.980 87.900 49.650 88.040 ;
        RECT 32.350 87.855 32.640 87.900 ;
        RECT 34.450 87.855 34.740 87.900 ;
        RECT 36.020 87.855 36.310 87.900 ;
        RECT 49.330 87.840 49.650 87.900 ;
        RECT 50.340 87.760 50.480 88.240 ;
        RECT 54.865 88.195 55.155 88.240 ;
        RECT 57.150 88.180 57.470 88.440 ;
        RECT 58.045 88.380 58.335 88.425 ;
        RECT 59.235 88.380 59.525 88.425 ;
        RECT 61.755 88.380 62.045 88.425 ;
        RECT 58.045 88.240 62.045 88.380 ;
        RECT 58.045 88.195 58.335 88.240 ;
        RECT 59.235 88.195 59.525 88.240 ;
        RECT 61.755 88.195 62.045 88.240 ;
        RECT 65.890 88.380 66.210 88.440 ;
        RECT 67.360 88.380 67.500 88.580 ;
        RECT 67.875 88.535 68.165 88.580 ;
        RECT 68.650 88.720 68.970 88.780 ;
        RECT 70.045 88.720 70.335 88.765 ;
        RECT 70.490 88.720 70.810 88.780 ;
        RECT 68.650 88.580 70.810 88.720 ;
        RECT 68.650 88.520 68.970 88.580 ;
        RECT 70.045 88.535 70.335 88.580 ;
        RECT 70.490 88.520 70.810 88.580 ;
        RECT 72.790 88.520 73.110 88.780 ;
        RECT 73.340 88.765 73.480 88.920 ;
        RECT 73.265 88.535 73.555 88.765 ;
        RECT 74.720 88.720 74.860 89.200 ;
        RECT 78.770 89.060 79.090 89.120 ;
        RECT 80.150 89.060 80.470 89.120 ;
        RECT 100.100 89.065 100.760 90.865 ;
        RECT 78.770 88.920 80.470 89.060 ;
        RECT 100.130 89.045 100.360 89.065 ;
        RECT 100.530 88.975 100.760 89.065 ;
        RECT 100.970 90.905 101.200 90.975 ;
        RECT 100.970 89.095 101.530 90.905 ;
        RECT 101.810 90.865 101.960 91.125 ;
        RECT 102.110 90.865 102.340 90.975 ;
        RECT 101.810 90.855 102.340 90.865 ;
        RECT 100.970 88.975 101.200 89.095 ;
        RECT 78.770 88.860 79.090 88.920 ;
        RECT 80.150 88.860 80.470 88.920 ;
        RECT 77.865 88.720 78.155 88.765 ;
        RECT 74.720 88.580 78.155 88.720 ;
        RECT 77.865 88.535 78.155 88.580 ;
        RECT 79.230 88.520 79.550 88.780 ;
        RECT 79.690 88.520 80.010 88.780 ;
        RECT 80.610 88.720 80.930 88.780 ;
        RECT 82.910 88.765 83.230 88.780 ;
        RECT 81.545 88.720 81.835 88.765 ;
        RECT 80.610 88.580 81.835 88.720 ;
        RECT 80.610 88.520 80.930 88.580 ;
        RECT 81.545 88.535 81.835 88.580 ;
        RECT 82.880 88.535 83.230 88.765 ;
        RECT 82.910 88.520 83.230 88.535 ;
        RECT 88.890 88.520 89.210 88.780 ;
        RECT 101.360 88.775 101.530 89.095 ;
        RECT 101.770 89.055 102.340 90.855 ;
        RECT 101.820 89.045 102.340 89.055 ;
        RECT 102.110 88.975 102.340 89.045 ;
        RECT 102.550 90.925 102.780 90.975 ;
        RECT 102.550 90.895 103.060 90.925 ;
        RECT 102.550 89.085 103.090 90.895 ;
        RECT 103.290 90.875 103.480 93.885 ;
        RECT 103.680 93.835 103.910 93.885 ;
        RECT 104.120 93.835 104.350 93.925 ;
        RECT 104.870 93.885 105.490 99.785 ;
        RECT 103.840 92.955 104.200 93.635 ;
        RECT 103.660 91.925 104.660 92.955 ;
        RECT 103.840 91.135 104.200 91.925 ;
        RECT 103.690 90.875 103.920 90.975 ;
        RECT 103.290 90.205 103.920 90.875 ;
        RECT 102.550 88.975 102.780 89.085 ;
        RECT 102.920 88.855 103.090 89.085 ;
        RECT 103.310 89.005 103.920 90.205 ;
        RECT 103.690 88.975 103.920 89.005 ;
        RECT 104.130 90.925 104.360 90.975 ;
        RECT 104.130 89.045 104.670 90.925 ;
        RECT 104.890 90.905 105.060 93.885 ;
        RECT 105.260 93.835 105.490 93.885 ;
        RECT 105.700 93.915 106.190 99.835 ;
        RECT 106.840 99.755 107.070 99.835 ;
        RECT 105.700 93.835 105.930 93.915 ;
        RECT 106.430 93.875 107.070 99.755 ;
        RECT 105.450 93.625 105.740 93.630 ;
        RECT 105.440 92.985 105.780 93.625 ;
        RECT 105.270 91.955 106.270 92.985 ;
        RECT 105.440 91.145 105.780 91.955 ;
        RECT 105.460 91.135 105.750 91.145 ;
        RECT 105.270 90.905 105.500 90.975 ;
        RECT 104.890 90.865 105.500 90.905 ;
        RECT 104.870 89.065 105.500 90.865 ;
        RECT 104.900 89.045 105.500 89.065 ;
        RECT 104.130 88.975 104.360 89.045 ;
        RECT 100.000 88.635 101.000 88.645 ;
        RECT 101.280 88.635 101.530 88.775 ;
        RECT 102.910 88.635 103.090 88.855 ;
        RECT 104.500 88.805 104.670 89.045 ;
        RECT 105.270 88.975 105.500 89.045 ;
        RECT 105.710 90.905 105.940 90.975 ;
        RECT 105.710 89.025 106.250 90.905 ;
        RECT 106.440 90.895 106.630 93.875 ;
        RECT 106.840 93.835 107.070 93.875 ;
        RECT 107.270 93.865 107.710 100.195 ;
        RECT 108.890 99.835 109.330 100.195 ;
        RECT 110.480 99.835 110.920 100.195 ;
        RECT 112.060 99.835 112.500 100.195 ;
        RECT 108.420 99.815 108.650 99.835 ;
        RECT 107.970 93.885 108.650 99.815 ;
        RECT 107.280 93.835 107.510 93.865 ;
        RECT 107.030 93.625 107.320 93.630 ;
        RECT 107.010 92.955 107.370 93.625 ;
        RECT 106.820 91.925 107.820 92.955 ;
        RECT 107.010 91.135 107.370 91.925 ;
        RECT 106.850 90.895 107.080 90.975 ;
        RECT 106.440 89.045 107.080 90.895 ;
        RECT 105.710 88.975 105.940 89.025 ;
        RECT 104.490 88.635 104.670 88.805 ;
        RECT 106.080 88.635 106.250 89.025 ;
        RECT 106.850 88.975 107.080 89.045 ;
        RECT 107.290 90.925 107.520 90.975 ;
        RECT 107.980 90.935 108.240 93.885 ;
        RECT 108.420 93.835 108.650 93.885 ;
        RECT 108.860 93.895 109.330 99.835 ;
        RECT 110.000 99.795 110.230 99.835 ;
        RECT 108.860 93.835 109.090 93.895 ;
        RECT 109.550 93.885 110.230 99.795 ;
        RECT 108.610 93.625 108.900 93.630 ;
        RECT 108.580 92.985 108.920 93.625 ;
        RECT 108.440 91.955 109.440 92.985 ;
        RECT 108.580 91.135 108.920 91.955 ;
        RECT 108.430 90.935 108.660 90.975 ;
        RECT 107.290 89.045 107.830 90.925 ;
        RECT 107.290 88.975 107.520 89.045 ;
        RECT 107.660 88.635 107.830 89.045 ;
        RECT 107.980 89.015 108.660 90.935 ;
        RECT 108.430 88.975 108.660 89.015 ;
        RECT 108.870 90.915 109.100 90.975 ;
        RECT 108.870 89.035 109.420 90.915 ;
        RECT 109.600 90.895 109.860 93.885 ;
        RECT 110.000 93.835 110.230 93.885 ;
        RECT 110.440 93.875 110.920 99.835 ;
        RECT 111.580 99.795 111.810 99.835 ;
        RECT 111.150 93.905 111.810 99.795 ;
        RECT 111.150 93.885 111.410 93.905 ;
        RECT 110.440 93.835 110.670 93.875 ;
        RECT 111.160 93.675 111.410 93.885 ;
        RECT 111.580 93.835 111.810 93.905 ;
        RECT 112.020 93.925 112.500 99.835 ;
        RECT 112.020 93.835 112.250 93.925 ;
        RECT 110.190 93.625 110.480 93.630 ;
        RECT 110.180 92.955 110.510 93.625 ;
        RECT 110.010 91.925 111.010 92.955 ;
        RECT 110.180 91.135 110.510 91.925 ;
        RECT 111.160 91.575 111.460 93.675 ;
        RECT 111.770 93.625 112.060 93.630 ;
        RECT 111.750 92.975 112.110 93.625 ;
        RECT 111.670 91.945 112.670 92.975 ;
        RECT 111.240 91.125 111.460 91.575 ;
        RECT 111.750 91.135 112.110 91.945 ;
        RECT 110.010 90.895 110.240 90.975 ;
        RECT 109.580 89.045 110.240 90.895 ;
        RECT 108.870 88.975 109.100 89.035 ;
        RECT 109.260 88.635 109.420 89.035 ;
        RECT 110.010 88.975 110.240 89.045 ;
        RECT 110.450 90.915 110.680 90.975 ;
        RECT 110.450 89.025 111.000 90.915 ;
        RECT 111.240 90.885 111.420 91.125 ;
        RECT 111.590 90.885 111.820 90.975 ;
        RECT 111.240 90.735 111.820 90.885 ;
        RECT 111.210 89.065 111.820 90.735 ;
        RECT 111.220 89.035 111.820 89.065 ;
        RECT 110.450 88.975 110.680 89.025 ;
        RECT 110.830 88.635 111.000 89.025 ;
        RECT 111.590 88.975 111.820 89.035 ;
        RECT 112.030 90.915 112.260 90.975 ;
        RECT 112.030 89.065 112.720 90.915 ;
        RECT 112.030 88.975 112.260 89.065 ;
        RECT 112.410 88.815 112.720 89.065 ;
        RECT 112.390 88.775 112.720 88.815 ;
        RECT 112.390 88.635 112.880 88.775 ;
        RECT 100.000 88.605 112.880 88.635 ;
        RECT 99.980 88.550 112.880 88.605 ;
        RECT 113.070 88.550 113.700 101.660 ;
        RECT 119.900 101.650 120.990 101.675 ;
        RECT 134.480 99.950 135.430 101.710 ;
        RECT 136.630 99.960 138.450 102.060 ;
        RECT 139.570 99.960 141.390 102.060 ;
        RECT 142.470 99.960 144.300 102.090 ;
        RECT 145.440 99.960 147.270 102.090 ;
        RECT 148.420 99.970 150.250 102.100 ;
        RECT 136.630 99.955 136.880 99.960 ;
        RECT 138.110 99.955 138.360 99.960 ;
        RECT 139.590 99.955 139.840 99.960 ;
        RECT 141.070 99.955 141.320 99.960 ;
        RECT 142.550 99.955 142.800 99.960 ;
        RECT 144.030 99.955 144.280 99.960 ;
        RECT 145.510 99.955 145.760 99.960 ;
        RECT 146.990 99.955 147.240 99.960 ;
        RECT 148.470 99.955 148.720 99.970 ;
        RECT 149.950 99.955 150.200 99.970 ;
        RECT 151.370 99.960 153.200 102.090 ;
        RECT 151.430 99.955 151.680 99.960 ;
        RECT 152.910 99.955 153.160 99.960 ;
        RECT 154.340 99.950 156.170 102.080 ;
        RECT 157.270 99.980 158.460 103.930 ;
        RECT 157.350 99.955 157.600 99.980 ;
        RECT 135.150 99.340 135.400 99.365 ;
        RECT 136.630 99.340 136.880 99.365 ;
        RECT 135.100 99.300 136.910 99.340 ;
        RECT 135.100 97.270 136.940 99.300 ;
        RECT 138.090 97.270 139.910 99.370 ;
        RECT 141.030 97.280 142.850 99.380 ;
        RECT 144.030 99.360 144.280 99.365 ;
        RECT 145.510 99.360 145.760 99.365 ;
        RECT 135.100 97.240 136.910 97.270 ;
        RECT 138.110 97.260 138.360 97.270 ;
        RECT 139.590 97.260 139.840 97.270 ;
        RECT 141.070 97.260 141.320 97.280 ;
        RECT 142.550 97.260 142.800 97.280 ;
        RECT 143.960 97.230 145.790 99.360 ;
        RECT 146.940 97.240 148.770 99.370 ;
        RECT 149.930 97.240 151.760 99.370 ;
        RECT 152.910 99.360 153.160 99.365 ;
        RECT 154.390 99.360 154.640 99.365 ;
        RECT 152.850 97.230 154.680 99.360 ;
        RECT 155.820 97.240 157.650 99.370 ;
        RECT 117.600 93.110 130.450 93.240 ;
        RECT 117.600 92.280 130.480 93.110 ;
        RECT 118.410 91.720 119.370 91.950 ;
        RECT 118.130 91.480 118.360 91.515 ;
        RECT 65.890 88.240 67.500 88.380 ;
        RECT 65.890 88.180 66.210 88.240 ;
        RECT 53.470 87.840 53.790 88.100 ;
        RECT 57.650 88.040 57.940 88.085 ;
        RECT 59.750 88.040 60.040 88.085 ;
        RECT 61.320 88.040 61.610 88.085 ;
        RECT 57.650 87.900 61.610 88.040 ;
        RECT 57.650 87.855 57.940 87.900 ;
        RECT 59.750 87.855 60.040 87.900 ;
        RECT 61.320 87.855 61.610 87.900 ;
        RECT 71.885 88.040 72.175 88.085 ;
        RECT 72.880 88.040 73.020 88.520 ;
        RECT 74.170 88.380 74.490 88.440 ;
        RECT 75.090 88.380 75.410 88.440 ;
        RECT 74.170 88.240 75.410 88.380 ;
        RECT 74.170 88.180 74.490 88.240 ;
        RECT 75.090 88.180 75.410 88.240 ;
        RECT 82.425 88.380 82.715 88.425 ;
        RECT 83.615 88.380 83.905 88.425 ;
        RECT 86.135 88.380 86.425 88.425 ;
        RECT 82.425 88.240 86.425 88.380 ;
        RECT 82.425 88.195 82.715 88.240 ;
        RECT 83.615 88.195 83.905 88.240 ;
        RECT 86.135 88.195 86.425 88.240 ;
        RECT 71.885 87.900 73.020 88.040 ;
        RECT 82.030 88.040 82.320 88.085 ;
        RECT 84.130 88.040 84.420 88.085 ;
        RECT 85.700 88.040 85.990 88.085 ;
        RECT 82.030 87.900 85.990 88.040 ;
        RECT 71.885 87.855 72.175 87.900 ;
        RECT 82.030 87.855 82.320 87.900 ;
        RECT 84.130 87.855 84.420 87.900 ;
        RECT 85.700 87.855 85.990 87.900 ;
        RECT 89.810 87.840 90.130 88.100 ;
        RECT 18.600 87.560 26.650 87.700 ;
        RECT 23.110 87.500 23.430 87.560 ;
        RECT 26.330 87.500 26.650 87.560 ;
        RECT 27.725 87.515 28.015 87.745 ;
        RECT 28.645 87.700 28.935 87.745 ;
        RECT 30.930 87.700 31.250 87.760 ;
        RECT 28.645 87.560 31.250 87.700 ;
        RECT 28.645 87.515 28.935 87.560 ;
        RECT 30.930 87.500 31.250 87.560 ;
        RECT 50.250 87.500 50.570 87.760 ;
        RECT 64.970 87.700 65.290 87.760 ;
        RECT 68.650 87.700 68.970 87.760 ;
        RECT 64.970 87.560 68.970 87.700 ;
        RECT 64.970 87.500 65.290 87.560 ;
        RECT 68.650 87.500 68.970 87.560 ;
        RECT 74.170 87.700 74.490 87.760 ;
        RECT 75.550 87.700 75.870 87.760 ;
        RECT 74.170 87.560 75.870 87.700 ;
        RECT 74.170 87.500 74.490 87.560 ;
        RECT 75.550 87.500 75.870 87.560 ;
        RECT 80.625 87.700 80.915 87.745 ;
        RECT 84.750 87.700 85.070 87.760 ;
        RECT 80.625 87.560 85.070 87.700 ;
        RECT 99.980 87.645 117.170 88.550 ;
        RECT 99.980 87.615 112.880 87.645 ;
        RECT 100.000 87.575 112.880 87.615 ;
        RECT 80.625 87.515 80.915 87.560 ;
        RECT 84.750 87.500 85.070 87.560 ;
        RECT 13.380 86.880 92.040 87.360 ;
        RECT 22.190 86.480 22.510 86.740 ;
        RECT 25.425 86.680 25.715 86.725 ;
        RECT 27.250 86.680 27.570 86.740 ;
        RECT 25.425 86.540 27.570 86.680 ;
        RECT 25.425 86.495 25.715 86.540 ;
        RECT 27.250 86.480 27.570 86.540 ;
        RECT 45.190 86.680 45.510 86.740 ;
        RECT 45.665 86.680 45.955 86.725 ;
        RECT 50.250 86.680 50.570 86.740 ;
        RECT 45.190 86.540 50.570 86.680 ;
        RECT 45.190 86.480 45.510 86.540 ;
        RECT 45.665 86.495 45.955 86.540 ;
        RECT 50.250 86.480 50.570 86.540 ;
        RECT 67.745 86.680 68.035 86.725 ;
        RECT 68.190 86.680 68.510 86.740 ;
        RECT 69.570 86.680 69.890 86.740 ;
        RECT 73.265 86.680 73.555 86.725 ;
        RECT 75.550 86.680 75.870 86.740 ;
        RECT 82.910 86.680 83.230 86.740 ;
        RECT 83.385 86.680 83.675 86.725 ;
        RECT 67.745 86.540 73.555 86.680 ;
        RECT 67.745 86.495 68.035 86.540 ;
        RECT 68.190 86.480 68.510 86.540 ;
        RECT 69.570 86.480 69.890 86.540 ;
        RECT 73.265 86.495 73.555 86.540 ;
        RECT 73.900 86.540 80.840 86.680 ;
        RECT 23.570 86.140 23.890 86.400 ;
        RECT 28.210 86.340 28.500 86.385 ;
        RECT 30.310 86.340 30.600 86.385 ;
        RECT 31.880 86.340 32.170 86.385 ;
        RECT 28.210 86.200 32.170 86.340 ;
        RECT 28.210 86.155 28.500 86.200 ;
        RECT 30.310 86.155 30.600 86.200 ;
        RECT 31.880 86.155 32.170 86.200 ;
        RECT 43.825 86.340 44.115 86.385 ;
        RECT 44.270 86.340 44.590 86.400 ;
        RECT 43.825 86.200 44.590 86.340 ;
        RECT 43.825 86.155 44.115 86.200 ;
        RECT 44.270 86.140 44.590 86.200 ;
        RECT 48.410 86.140 48.730 86.400 ;
        RECT 49.330 86.340 49.650 86.400 ;
        RECT 51.170 86.340 51.490 86.400 ;
        RECT 49.330 86.200 51.490 86.340 ;
        RECT 49.330 86.140 49.650 86.200 ;
        RECT 51.170 86.140 51.490 86.200 ;
        RECT 57.650 86.340 57.940 86.385 ;
        RECT 59.750 86.340 60.040 86.385 ;
        RECT 61.320 86.340 61.610 86.385 ;
        RECT 57.650 86.200 61.610 86.340 ;
        RECT 57.650 86.155 57.940 86.200 ;
        RECT 59.750 86.155 60.040 86.200 ;
        RECT 61.320 86.155 61.610 86.200 ;
        RECT 64.065 86.340 64.355 86.385 ;
        RECT 73.900 86.340 74.040 86.540 ;
        RECT 75.550 86.480 75.870 86.540 ;
        RECT 77.850 86.340 78.170 86.400 ;
        RECT 64.065 86.200 66.120 86.340 ;
        RECT 64.065 86.155 64.355 86.200 ;
        RECT 21.745 86.000 22.035 86.045 ;
        RECT 23.660 86.000 23.800 86.140 ;
        RECT 25.410 86.000 25.730 86.060 ;
        RECT 21.745 85.860 23.340 86.000 ;
        RECT 23.660 85.860 25.730 86.000 ;
        RECT 21.745 85.815 22.035 85.860 ;
        RECT 23.200 85.705 23.340 85.860 ;
        RECT 23.125 85.475 23.415 85.705 ;
        RECT 23.570 85.460 23.890 85.720 ;
        RECT 25.040 85.705 25.180 85.860 ;
        RECT 25.410 85.800 25.730 85.860 ;
        RECT 26.790 86.000 27.110 86.060 ;
        RECT 27.725 86.000 28.015 86.045 ;
        RECT 26.790 85.860 28.015 86.000 ;
        RECT 26.790 85.800 27.110 85.860 ;
        RECT 27.725 85.815 28.015 85.860 ;
        RECT 28.605 86.000 28.895 86.045 ;
        RECT 29.795 86.000 30.085 86.045 ;
        RECT 32.315 86.000 32.605 86.045 ;
        RECT 28.605 85.860 32.605 86.000 ;
        RECT 28.605 85.815 28.895 85.860 ;
        RECT 29.795 85.815 30.085 85.860 ;
        RECT 32.315 85.815 32.605 85.860 ;
        RECT 55.770 85.800 56.090 86.060 ;
        RECT 57.150 85.800 57.470 86.060 ;
        RECT 58.045 86.000 58.335 86.045 ;
        RECT 59.235 86.000 59.525 86.045 ;
        RECT 61.755 86.000 62.045 86.045 ;
        RECT 64.525 86.000 64.815 86.045 ;
        RECT 58.045 85.860 62.045 86.000 ;
        RECT 58.045 85.815 58.335 85.860 ;
        RECT 59.235 85.815 59.525 85.860 ;
        RECT 61.755 85.815 62.045 85.860 ;
        RECT 62.300 85.860 64.815 86.000 ;
        RECT 24.965 85.475 25.255 85.705 ;
        RECT 43.365 85.475 43.655 85.705 ;
        RECT 58.500 85.660 58.790 85.705 ;
        RECT 62.300 85.660 62.440 85.860 ;
        RECT 64.525 85.815 64.815 85.860 ;
        RECT 58.500 85.520 62.440 85.660 ;
        RECT 58.500 85.475 58.790 85.520 ;
        RECT 19.905 85.320 20.195 85.365 ;
        RECT 20.825 85.320 21.115 85.365 ;
        RECT 22.190 85.320 22.510 85.380 ;
        RECT 19.905 85.180 20.580 85.320 ;
        RECT 19.905 85.135 20.195 85.180 ;
        RECT 20.440 85.040 20.580 85.180 ;
        RECT 20.825 85.180 22.510 85.320 ;
        RECT 20.825 85.135 21.115 85.180 ;
        RECT 22.190 85.120 22.510 85.180 ;
        RECT 28.170 85.320 28.490 85.380 ;
        RECT 28.950 85.320 29.240 85.365 ;
        RECT 28.170 85.180 29.240 85.320 ;
        RECT 43.440 85.320 43.580 85.475 ;
        RECT 65.430 85.460 65.750 85.720 ;
        RECT 65.980 85.705 66.120 86.200 ;
        RECT 73.340 86.200 74.040 86.340 ;
        RECT 74.260 86.200 78.170 86.340 ;
        RECT 73.340 86.060 73.480 86.200 ;
        RECT 69.660 85.860 70.720 86.000 ;
        RECT 65.905 85.660 66.195 85.705 ;
        RECT 66.350 85.660 66.670 85.720 ;
        RECT 65.905 85.520 66.670 85.660 ;
        RECT 65.905 85.475 66.195 85.520 ;
        RECT 66.350 85.460 66.670 85.520 ;
        RECT 66.825 85.475 67.115 85.705 ;
        RECT 67.285 85.660 67.575 85.705 ;
        RECT 67.730 85.660 68.050 85.720 ;
        RECT 67.285 85.520 68.050 85.660 ;
        RECT 67.285 85.475 67.575 85.520 ;
        RECT 45.650 85.320 45.970 85.380 ;
        RECT 43.440 85.180 45.970 85.320 ;
        RECT 28.170 85.120 28.490 85.180 ;
        RECT 28.950 85.135 29.240 85.180 ;
        RECT 45.650 85.120 45.970 85.180 ;
        RECT 50.250 85.320 50.570 85.380 ;
        RECT 53.010 85.320 53.330 85.380 ;
        RECT 50.250 85.180 53.330 85.320 ;
        RECT 50.250 85.120 50.570 85.180 ;
        RECT 53.010 85.120 53.330 85.180 ;
        RECT 20.350 84.980 20.670 85.040 ;
        RECT 22.650 84.980 22.970 85.040 ;
        RECT 20.350 84.840 22.970 84.980 ;
        RECT 20.350 84.780 20.670 84.840 ;
        RECT 22.650 84.780 22.970 84.840 ;
        RECT 34.610 84.780 34.930 85.040 ;
        RECT 40.130 84.780 40.450 85.040 ;
        RECT 46.570 84.780 46.890 85.040 ;
        RECT 47.965 84.980 48.255 85.025 ;
        RECT 49.330 84.980 49.650 85.040 ;
        RECT 47.965 84.840 49.650 84.980 ;
        RECT 47.965 84.795 48.255 84.840 ;
        RECT 49.330 84.780 49.650 84.840 ;
        RECT 52.550 84.780 52.870 85.040 ;
        RECT 54.390 84.780 54.710 85.040 ;
        RECT 54.865 84.980 55.155 85.025 ;
        RECT 57.610 84.980 57.930 85.040 ;
        RECT 54.865 84.840 57.930 84.980 ;
        RECT 54.865 84.795 55.155 84.840 ;
        RECT 57.610 84.780 57.930 84.840 ;
        RECT 65.890 84.980 66.210 85.040 ;
        RECT 66.900 84.980 67.040 85.475 ;
        RECT 67.730 85.460 68.050 85.520 ;
        RECT 68.650 85.460 68.970 85.720 ;
        RECT 69.660 85.705 69.800 85.860 ;
        RECT 70.580 85.720 70.720 85.860 ;
        RECT 73.250 85.800 73.570 86.060 ;
        RECT 74.260 86.045 74.400 86.200 ;
        RECT 77.850 86.140 78.170 86.200 ;
        RECT 74.185 85.815 74.475 86.045 ;
        RECT 76.930 86.000 77.250 86.060 ;
        RECT 77.405 86.000 77.695 86.045 ;
        RECT 80.165 86.000 80.455 86.045 ;
        RECT 76.930 85.860 80.455 86.000 ;
        RECT 76.930 85.800 77.250 85.860 ;
        RECT 77.405 85.815 77.695 85.860 ;
        RECT 80.165 85.815 80.455 85.860 ;
        RECT 69.585 85.475 69.875 85.705 ;
        RECT 70.045 85.475 70.335 85.705 ;
        RECT 70.490 85.660 70.810 85.720 ;
        RECT 70.965 85.660 71.255 85.705 ;
        RECT 70.490 85.520 71.255 85.660 ;
        RECT 65.890 84.840 67.040 84.980 ;
        RECT 68.740 84.980 68.880 85.460 ;
        RECT 70.120 84.980 70.260 85.475 ;
        RECT 70.490 85.460 70.810 85.520 ;
        RECT 70.965 85.475 71.255 85.520 ;
        RECT 72.790 85.460 73.110 85.720 ;
        RECT 74.630 85.660 74.950 85.720 ;
        RECT 75.565 85.660 75.855 85.705 ;
        RECT 74.630 85.520 75.855 85.660 ;
        RECT 74.630 85.460 74.950 85.520 ;
        RECT 75.565 85.475 75.855 85.520 ;
        RECT 78.325 85.475 78.615 85.705 ;
        RECT 79.245 85.475 79.535 85.705 ;
        RECT 79.705 85.660 79.995 85.705 ;
        RECT 80.700 85.660 80.840 86.540 ;
        RECT 82.910 86.540 83.675 86.680 ;
        RECT 82.910 86.480 83.230 86.540 ;
        RECT 83.385 86.495 83.675 86.540 ;
        RECT 88.445 86.680 88.735 86.725 ;
        RECT 88.890 86.680 89.210 86.740 ;
        RECT 88.445 86.540 89.210 86.680 ;
        RECT 88.445 86.495 88.735 86.540 ;
        RECT 88.890 86.480 89.210 86.540 ;
        RECT 82.005 86.000 82.295 86.045 ;
        RECT 86.145 86.000 86.435 86.045 ;
        RECT 82.005 85.860 86.435 86.000 ;
        RECT 82.005 85.815 82.295 85.860 ;
        RECT 86.145 85.815 86.435 85.860 ;
        RECT 79.705 85.520 80.840 85.660 ;
        RECT 81.085 85.660 81.375 85.705 ;
        RECT 81.530 85.660 81.850 85.720 ;
        RECT 81.085 85.520 81.850 85.660 ;
        RECT 79.705 85.475 79.995 85.520 ;
        RECT 81.085 85.475 81.375 85.520 ;
        RECT 76.470 85.120 76.790 85.380 ;
        RECT 77.390 85.320 77.710 85.380 ;
        RECT 78.400 85.320 78.540 85.475 ;
        RECT 77.390 85.180 78.540 85.320 ;
        RECT 77.390 85.120 77.710 85.180 ;
        RECT 68.740 84.840 70.260 84.980 ;
        RECT 65.890 84.780 66.210 84.840 ;
        RECT 70.490 84.780 70.810 85.040 ;
        RECT 74.185 84.980 74.475 85.025 ;
        RECT 76.010 84.980 76.330 85.040 ;
        RECT 79.320 84.980 79.460 85.475 ;
        RECT 81.530 85.460 81.850 85.520 ;
        RECT 85.225 85.660 85.515 85.705 ;
        RECT 87.050 85.660 87.370 85.720 ;
        RECT 85.225 85.520 87.370 85.660 ;
        RECT 85.225 85.475 85.515 85.520 ;
        RECT 87.050 85.460 87.370 85.520 ;
        RECT 87.510 85.460 87.830 85.720 ;
        RECT 84.750 85.320 85.070 85.380 ;
        RECT 85.685 85.320 85.975 85.365 ;
        RECT 84.750 85.180 85.975 85.320 ;
        RECT 84.750 85.120 85.070 85.180 ;
        RECT 85.685 85.135 85.975 85.180 ;
        RECT 74.185 84.840 79.460 84.980 ;
        RECT 100.540 84.895 101.150 87.235 ;
        RECT 101.980 87.045 102.640 87.365 ;
        RECT 102.030 84.925 102.640 87.045 ;
        RECT 102.480 84.895 102.640 84.925 ;
        RECT 103.500 84.885 104.050 87.235 ;
        RECT 105.010 84.865 105.560 87.215 ;
        RECT 106.470 84.895 107.020 87.245 ;
        RECT 107.950 84.925 108.500 87.275 ;
        RECT 109.400 84.915 109.950 87.265 ;
        RECT 110.900 84.925 111.450 87.275 ;
        RECT 112.320 87.135 112.880 87.575 ;
        RECT 112.320 84.975 112.890 87.135 ;
        RECT 112.320 84.965 112.880 84.975 ;
        RECT 74.185 84.795 74.475 84.840 ;
        RECT 76.010 84.780 76.330 84.840 ;
        RECT 13.380 84.160 92.040 84.640 ;
        RECT 28.170 83.760 28.490 84.020 ;
        RECT 45.650 83.960 45.970 84.020 ;
        RECT 46.585 83.960 46.875 84.005 ;
        RECT 45.650 83.820 46.875 83.960 ;
        RECT 45.650 83.760 45.970 83.820 ;
        RECT 46.585 83.775 46.875 83.820 ;
        RECT 47.045 83.960 47.335 84.005 ;
        RECT 47.950 83.960 48.270 84.020 ;
        RECT 47.045 83.820 48.270 83.960 ;
        RECT 47.045 83.775 47.335 83.820 ;
        RECT 47.950 83.760 48.270 83.820 ;
        RECT 56.690 83.960 57.010 84.020 ;
        RECT 57.165 83.960 57.455 84.005 ;
        RECT 56.690 83.820 57.455 83.960 ;
        RECT 56.690 83.760 57.010 83.820 ;
        RECT 57.165 83.775 57.455 83.820 ;
        RECT 27.710 83.620 28.030 83.680 ;
        RECT 30.485 83.620 30.775 83.665 ;
        RECT 42.430 83.620 42.750 83.680 ;
        RECT 48.870 83.620 49.190 83.680 ;
        RECT 27.710 83.480 30.775 83.620 ;
        RECT 27.710 83.420 28.030 83.480 ;
        RECT 30.485 83.435 30.775 83.480 ;
        RECT 39.760 83.480 49.190 83.620 ;
        RECT 30.025 83.280 30.315 83.325 ;
        RECT 31.390 83.280 31.710 83.340 ;
        RECT 34.610 83.280 34.930 83.340 ;
        RECT 39.760 83.325 39.900 83.480 ;
        RECT 42.430 83.420 42.750 83.480 ;
        RECT 48.870 83.420 49.190 83.480 ;
        RECT 49.330 83.420 49.650 83.680 ;
        RECT 51.600 83.620 51.890 83.665 ;
        RECT 52.550 83.620 52.870 83.680 ;
        RECT 51.600 83.480 52.870 83.620 ;
        RECT 51.600 83.435 51.890 83.480 ;
        RECT 52.550 83.420 52.870 83.480 ;
        RECT 41.050 83.325 41.370 83.340 ;
        RECT 30.025 83.140 34.930 83.280 ;
        RECT 30.025 83.095 30.315 83.140 ;
        RECT 31.390 83.080 31.710 83.140 ;
        RECT 34.610 83.080 34.930 83.140 ;
        RECT 39.685 83.095 39.975 83.325 ;
        RECT 41.020 83.095 41.370 83.325 ;
        RECT 41.050 83.080 41.370 83.095 ;
        RECT 47.030 83.280 47.350 83.340 ;
        RECT 47.965 83.280 48.255 83.325 ;
        RECT 47.030 83.140 48.255 83.280 ;
        RECT 57.240 83.280 57.380 83.775 ;
        RECT 57.610 83.760 57.930 84.020 ;
        RECT 66.810 83.960 67.130 84.020 ;
        RECT 68.205 83.960 68.495 84.005 ;
        RECT 69.110 83.960 69.430 84.020 ;
        RECT 70.490 83.960 70.810 84.020 ;
        RECT 66.810 83.820 70.810 83.960 ;
        RECT 66.810 83.760 67.130 83.820 ;
        RECT 68.205 83.775 68.495 83.820 ;
        RECT 69.110 83.760 69.430 83.820 ;
        RECT 70.490 83.760 70.810 83.820 ;
        RECT 71.410 83.960 71.730 84.020 ;
        RECT 74.170 83.960 74.490 84.020 ;
        RECT 75.895 83.960 76.185 84.005 ;
        RECT 71.410 83.820 76.185 83.960 ;
        RECT 71.410 83.760 71.730 83.820 ;
        RECT 74.170 83.760 74.490 83.820 ;
        RECT 75.895 83.775 76.185 83.820 ;
        RECT 99.980 83.715 100.370 83.725 ;
        RECT 71.885 83.620 72.175 83.665 ;
        RECT 72.790 83.620 73.110 83.680 ;
        RECT 66.485 83.480 73.110 83.620 ;
        RECT 66.485 83.340 66.625 83.480 ;
        RECT 71.885 83.435 72.175 83.480 ;
        RECT 72.790 83.420 73.110 83.480 ;
        RECT 76.930 83.420 77.250 83.680 ;
        RECT 60.385 83.280 60.675 83.325 ;
        RECT 57.240 83.140 60.675 83.280 ;
        RECT 47.030 83.080 47.350 83.140 ;
        RECT 47.965 83.095 48.255 83.140 ;
        RECT 60.385 83.095 60.675 83.140 ;
        RECT 66.350 83.080 66.670 83.340 ;
        RECT 79.230 83.280 79.550 83.340 ;
        RECT 66.900 83.140 79.550 83.280 ;
        RECT 30.930 82.740 31.250 83.000 ;
        RECT 40.565 82.940 40.855 82.985 ;
        RECT 41.755 82.940 42.045 82.985 ;
        RECT 44.275 82.940 44.565 82.985 ;
        RECT 40.565 82.800 44.565 82.940 ;
        RECT 40.565 82.755 40.855 82.800 ;
        RECT 41.755 82.755 42.045 82.800 ;
        RECT 44.275 82.755 44.565 82.800 ;
        RECT 46.570 82.940 46.890 83.000 ;
        RECT 48.425 82.940 48.715 82.985 ;
        RECT 46.570 82.800 48.715 82.940 ;
        RECT 46.570 82.740 46.890 82.800 ;
        RECT 48.425 82.755 48.715 82.800 ;
        RECT 48.870 82.940 49.190 83.000 ;
        RECT 50.265 82.940 50.555 82.985 ;
        RECT 48.870 82.800 50.555 82.940 ;
        RECT 48.870 82.740 49.190 82.800 ;
        RECT 50.265 82.755 50.555 82.800 ;
        RECT 51.145 82.940 51.435 82.985 ;
        RECT 52.335 82.940 52.625 82.985 ;
        RECT 54.855 82.940 55.145 82.985 ;
        RECT 51.145 82.800 55.145 82.940 ;
        RECT 51.145 82.755 51.435 82.800 ;
        RECT 52.335 82.755 52.625 82.800 ;
        RECT 54.855 82.755 55.145 82.800 ;
        RECT 40.170 82.600 40.460 82.645 ;
        RECT 42.270 82.600 42.560 82.645 ;
        RECT 43.840 82.600 44.130 82.645 ;
        RECT 50.750 82.600 51.040 82.645 ;
        RECT 52.850 82.600 53.140 82.645 ;
        RECT 54.420 82.600 54.710 82.645 ;
        RECT 40.170 82.460 44.130 82.600 ;
        RECT 40.170 82.415 40.460 82.460 ;
        RECT 42.270 82.415 42.560 82.460 ;
        RECT 43.840 82.415 44.130 82.460 ;
        RECT 44.360 82.460 49.975 82.600 ;
        RECT 34.610 82.260 34.930 82.320 ;
        RECT 44.360 82.260 44.500 82.460 ;
        RECT 34.610 82.120 44.500 82.260 ;
        RECT 34.610 82.060 34.930 82.120 ;
        RECT 49.330 82.060 49.650 82.320 ;
        RECT 49.835 82.260 49.975 82.460 ;
        RECT 50.750 82.460 54.710 82.600 ;
        RECT 50.750 82.415 51.040 82.460 ;
        RECT 52.850 82.415 53.140 82.460 ;
        RECT 54.420 82.415 54.710 82.460 ;
        RECT 66.900 82.260 67.040 83.140 ;
        RECT 79.230 83.080 79.550 83.140 ;
        RECT 85.685 83.280 85.975 83.325 ;
        RECT 88.430 83.280 88.750 83.340 ;
        RECT 89.825 83.280 90.115 83.325 ;
        RECT 85.685 83.140 90.115 83.280 ;
        RECT 85.685 83.095 85.975 83.140 ;
        RECT 88.430 83.080 88.750 83.140 ;
        RECT 89.825 83.095 90.115 83.140 ;
        RECT 72.330 82.940 72.650 83.000 ;
        RECT 69.200 82.800 72.650 82.940 ;
        RECT 69.200 82.645 69.340 82.800 ;
        RECT 72.330 82.740 72.650 82.800 ;
        RECT 99.980 82.780 101.000 83.715 ;
        RECT 69.125 82.415 69.415 82.645 ;
        RECT 70.030 82.400 70.350 82.660 ;
        RECT 74.630 82.600 74.950 82.660 ;
        RECT 72.500 82.460 74.950 82.600 ;
        RECT 49.835 82.120 67.040 82.260 ;
        RECT 68.190 82.060 68.510 82.320 ;
        RECT 69.585 82.260 69.875 82.305 ;
        RECT 72.500 82.260 72.640 82.460 ;
        RECT 74.630 82.400 74.950 82.460 ;
        RECT 69.585 82.120 72.640 82.260 ;
        RECT 72.790 82.260 73.110 82.320 ;
        RECT 75.105 82.260 75.395 82.305 ;
        RECT 72.790 82.120 75.395 82.260 ;
        RECT 69.585 82.075 69.875 82.120 ;
        RECT 72.790 82.060 73.110 82.120 ;
        RECT 75.105 82.075 75.395 82.120 ;
        RECT 76.010 82.060 76.330 82.320 ;
        RECT 86.590 82.060 86.910 82.320 ;
        RECT 87.050 82.060 87.370 82.320 ;
        RECT 13.380 81.440 92.040 81.920 ;
        RECT 99.980 81.760 101.030 82.780 ;
        RECT 99.980 81.555 101.000 81.760 ;
        RECT 22.650 81.240 22.970 81.300 ;
        RECT 23.585 81.240 23.875 81.285 ;
        RECT 24.490 81.240 24.810 81.300 ;
        RECT 19.060 81.100 24.810 81.240 ;
        RECT 19.060 80.605 19.200 81.100 ;
        RECT 22.650 81.040 22.970 81.100 ;
        RECT 23.585 81.055 23.875 81.100 ;
        RECT 24.490 81.040 24.810 81.100 ;
        RECT 41.050 81.240 41.370 81.300 ;
        RECT 42.445 81.240 42.735 81.285 ;
        RECT 41.050 81.100 42.735 81.240 ;
        RECT 41.050 81.040 41.370 81.100 ;
        RECT 42.445 81.055 42.735 81.100 ;
        RECT 49.330 81.240 49.650 81.300 ;
        RECT 52.565 81.240 52.855 81.285 ;
        RECT 49.330 81.100 52.855 81.240 ;
        RECT 49.330 81.040 49.650 81.100 ;
        RECT 52.565 81.055 52.855 81.100 ;
        RECT 53.010 81.240 53.330 81.300 ;
        RECT 53.485 81.240 53.775 81.285 ;
        RECT 53.010 81.100 53.775 81.240 ;
        RECT 53.010 81.040 53.330 81.100 ;
        RECT 53.485 81.055 53.775 81.100 ;
        RECT 54.390 81.240 54.710 81.300 ;
        RECT 54.865 81.240 55.155 81.285 ;
        RECT 54.390 81.100 55.155 81.240 ;
        RECT 54.390 81.040 54.710 81.100 ;
        RECT 54.865 81.055 55.155 81.100 ;
        RECT 68.190 81.240 68.510 81.300 ;
        RECT 69.125 81.240 69.415 81.285 ;
        RECT 68.190 81.100 69.415 81.240 ;
        RECT 68.190 81.040 68.510 81.100 ;
        RECT 69.125 81.055 69.415 81.100 ;
        RECT 77.405 81.240 77.695 81.285 ;
        RECT 86.130 81.240 86.450 81.300 ;
        RECT 77.405 81.100 86.450 81.240 ;
        RECT 77.405 81.055 77.695 81.100 ;
        RECT 86.130 81.040 86.450 81.100 ;
        RECT 88.430 81.040 88.750 81.300 ;
        RECT 89.810 81.040 90.130 81.300 ;
        RECT 22.190 80.900 22.510 80.960 ;
        RECT 25.885 80.900 26.175 80.945 ;
        RECT 35.530 80.900 35.850 80.960 ;
        RECT 73.710 80.900 74.030 80.960 ;
        RECT 76.930 80.900 77.250 80.960 ;
        RECT 19.520 80.760 24.720 80.900 ;
        RECT 18.985 80.375 19.275 80.605 ;
        RECT 19.520 80.265 19.660 80.760 ;
        RECT 22.190 80.700 22.510 80.760 ;
        RECT 19.905 80.560 20.195 80.605 ;
        RECT 23.570 80.560 23.890 80.620 ;
        RECT 19.905 80.420 23.890 80.560 ;
        RECT 19.905 80.375 20.195 80.420 ;
        RECT 18.065 80.035 18.355 80.265 ;
        RECT 19.445 80.035 19.735 80.265 ;
        RECT 18.140 79.880 18.280 80.035 ;
        RECT 20.350 80.020 20.670 80.280 ;
        RECT 20.900 80.265 21.040 80.420 ;
        RECT 23.570 80.360 23.890 80.420 ;
        RECT 20.825 80.035 21.115 80.265 ;
        RECT 21.745 80.220 22.035 80.265 ;
        RECT 22.650 80.220 22.970 80.280 ;
        RECT 24.580 80.265 24.720 80.760 ;
        RECT 25.885 80.760 31.160 80.900 ;
        RECT 25.885 80.715 26.175 80.760 ;
        RECT 31.020 80.605 31.160 80.760 ;
        RECT 35.530 80.760 70.030 80.900 ;
        RECT 35.530 80.700 35.850 80.760 ;
        RECT 30.945 80.375 31.235 80.605 ;
        RECT 38.290 80.560 38.610 80.620 ;
        RECT 39.225 80.560 39.515 80.605 ;
        RECT 38.290 80.420 39.515 80.560 ;
        RECT 38.290 80.360 38.610 80.420 ;
        RECT 39.225 80.375 39.515 80.420 ;
        RECT 21.745 80.080 22.970 80.220 ;
        RECT 21.745 80.035 22.035 80.080 ;
        RECT 20.900 79.880 21.040 80.035 ;
        RECT 22.650 80.020 22.970 80.080 ;
        RECT 23.125 80.035 23.415 80.265 ;
        RECT 24.505 80.035 24.795 80.265 ;
        RECT 27.710 80.220 28.030 80.280 ;
        RECT 30.025 80.220 30.315 80.265 ;
        RECT 27.710 80.080 30.315 80.220 ;
        RECT 39.300 80.220 39.440 80.375 ;
        RECT 40.130 80.360 40.450 80.620 ;
        RECT 46.110 80.560 46.430 80.620 ;
        RECT 47.505 80.560 47.795 80.605 ;
        RECT 46.110 80.420 47.795 80.560 ;
        RECT 46.110 80.360 46.430 80.420 ;
        RECT 47.505 80.375 47.795 80.420 ;
        RECT 48.410 80.360 48.730 80.620 ;
        RECT 57.625 80.560 57.915 80.605 ;
        RECT 58.530 80.560 58.850 80.620 ;
        RECT 57.625 80.420 58.850 80.560 ;
        RECT 69.890 80.560 70.030 80.760 ;
        RECT 73.710 80.760 77.250 80.900 ;
        RECT 73.710 80.700 74.030 80.760 ;
        RECT 76.930 80.700 77.250 80.760 ;
        RECT 82.030 80.900 82.320 80.945 ;
        RECT 84.130 80.900 84.420 80.945 ;
        RECT 85.700 80.900 85.990 80.945 ;
        RECT 82.030 80.760 85.990 80.900 ;
        RECT 82.030 80.715 82.320 80.760 ;
        RECT 84.130 80.715 84.420 80.760 ;
        RECT 85.700 80.715 85.990 80.760 ;
        RECT 80.610 80.560 80.930 80.620 ;
        RECT 81.545 80.560 81.835 80.605 ;
        RECT 69.890 80.420 79.920 80.560 ;
        RECT 57.625 80.375 57.915 80.420 ;
        RECT 58.530 80.360 58.850 80.420 ;
        RECT 41.970 80.220 42.290 80.280 ;
        RECT 39.300 80.080 42.290 80.220 ;
        RECT 18.140 79.740 21.040 79.880 ;
        RECT 21.270 79.680 21.590 79.940 ;
        RECT 17.145 79.540 17.435 79.585 ;
        RECT 18.510 79.540 18.830 79.600 ;
        RECT 17.145 79.400 18.830 79.540 ;
        RECT 17.145 79.355 17.435 79.400 ;
        RECT 18.510 79.340 18.830 79.400 ;
        RECT 20.810 79.540 21.130 79.600 ;
        RECT 23.200 79.540 23.340 80.035 ;
        RECT 23.570 79.880 23.890 79.940 ;
        RECT 24.580 79.880 24.720 80.035 ;
        RECT 27.710 80.020 28.030 80.080 ;
        RECT 30.025 80.035 30.315 80.080 ;
        RECT 41.970 80.020 42.290 80.080 ;
        RECT 57.165 80.220 57.455 80.265 ;
        RECT 58.070 80.220 58.390 80.280 ;
        RECT 64.525 80.220 64.815 80.265 ;
        RECT 57.165 80.080 64.815 80.220 ;
        RECT 57.165 80.035 57.455 80.080 ;
        RECT 58.070 80.020 58.390 80.080 ;
        RECT 64.525 80.035 64.815 80.080 ;
        RECT 67.745 80.220 68.035 80.265 ;
        RECT 70.950 80.220 71.270 80.280 ;
        RECT 67.745 80.080 71.270 80.220 ;
        RECT 67.745 80.035 68.035 80.080 ;
        RECT 70.950 80.020 71.270 80.080 ;
        RECT 73.710 80.020 74.030 80.280 ;
        RECT 74.645 80.035 74.935 80.265 ;
        RECT 75.105 80.035 75.395 80.265 ;
        RECT 23.570 79.740 24.720 79.880 ;
        RECT 52.090 79.880 52.410 79.940 ;
        RECT 54.405 79.880 54.695 79.925 ;
        RECT 52.090 79.740 54.695 79.880 ;
        RECT 23.570 79.680 23.890 79.740 ;
        RECT 52.090 79.680 52.410 79.740 ;
        RECT 54.405 79.695 54.695 79.740 ;
        RECT 66.350 79.880 66.670 79.940 ;
        RECT 69.110 79.925 69.430 79.940 ;
        RECT 68.205 79.880 68.495 79.925 ;
        RECT 66.350 79.740 68.495 79.880 ;
        RECT 66.350 79.680 66.670 79.740 ;
        RECT 68.205 79.695 68.495 79.740 ;
        RECT 69.110 79.695 69.495 79.925 ;
        RECT 69.110 79.680 69.430 79.695 ;
        RECT 20.810 79.400 23.340 79.540 ;
        RECT 28.185 79.540 28.475 79.585 ;
        RECT 29.090 79.540 29.410 79.600 ;
        RECT 28.185 79.400 29.410 79.540 ;
        RECT 20.810 79.340 21.130 79.400 ;
        RECT 28.185 79.355 28.475 79.400 ;
        RECT 29.090 79.340 29.410 79.400 ;
        RECT 30.485 79.540 30.775 79.585 ;
        RECT 35.530 79.540 35.850 79.600 ;
        RECT 30.485 79.400 35.850 79.540 ;
        RECT 30.485 79.355 30.775 79.400 ;
        RECT 35.530 79.340 35.850 79.400 ;
        RECT 40.605 79.540 40.895 79.585 ;
        RECT 42.890 79.540 43.210 79.600 ;
        RECT 40.605 79.400 43.210 79.540 ;
        RECT 40.605 79.355 40.895 79.400 ;
        RECT 42.890 79.340 43.210 79.400 ;
        RECT 44.730 79.340 45.050 79.600 ;
        RECT 51.630 79.340 51.950 79.600 ;
        RECT 53.405 79.540 53.695 79.585 ;
        RECT 55.310 79.540 55.630 79.600 ;
        RECT 53.405 79.400 55.630 79.540 ;
        RECT 53.405 79.355 53.695 79.400 ;
        RECT 55.310 79.340 55.630 79.400 ;
        RECT 56.705 79.540 56.995 79.585 ;
        RECT 59.450 79.540 59.770 79.600 ;
        RECT 56.705 79.400 59.770 79.540 ;
        RECT 56.705 79.355 56.995 79.400 ;
        RECT 59.450 79.340 59.770 79.400 ;
        RECT 70.030 79.540 70.350 79.600 ;
        RECT 74.720 79.540 74.860 80.035 ;
        RECT 75.180 79.880 75.320 80.035 ;
        RECT 75.550 80.020 75.870 80.280 ;
        RECT 76.010 80.220 76.330 80.280 ;
        RECT 76.485 80.220 76.775 80.265 ;
        RECT 76.010 80.080 76.775 80.220 ;
        RECT 76.010 80.020 76.330 80.080 ;
        RECT 76.485 80.035 76.775 80.080 ;
        RECT 78.310 80.020 78.630 80.280 ;
        RECT 78.770 80.220 79.090 80.280 ;
        RECT 79.780 80.265 79.920 80.420 ;
        RECT 80.610 80.420 81.835 80.560 ;
        RECT 80.610 80.360 80.930 80.420 ;
        RECT 81.545 80.375 81.835 80.420 ;
        RECT 82.425 80.560 82.715 80.605 ;
        RECT 83.615 80.560 83.905 80.605 ;
        RECT 86.135 80.560 86.425 80.605 ;
        RECT 82.425 80.420 86.425 80.560 ;
        RECT 82.425 80.375 82.715 80.420 ;
        RECT 83.615 80.375 83.905 80.420 ;
        RECT 86.135 80.375 86.425 80.420 ;
        RECT 79.245 80.220 79.535 80.265 ;
        RECT 78.770 80.080 79.535 80.220 ;
        RECT 78.770 80.020 79.090 80.080 ;
        RECT 79.245 80.035 79.535 80.080 ;
        RECT 79.705 80.035 79.995 80.265 ;
        RECT 80.150 80.020 80.470 80.280 ;
        RECT 86.590 80.220 86.910 80.280 ;
        RECT 88.905 80.220 89.195 80.265 ;
        RECT 86.590 80.080 89.195 80.220 ;
        RECT 86.590 80.020 86.910 80.080 ;
        RECT 88.905 80.035 89.195 80.080 ;
        RECT 81.530 79.880 81.850 79.940 ;
        RECT 75.180 79.740 81.850 79.880 ;
        RECT 79.320 79.600 79.460 79.740 ;
        RECT 81.530 79.680 81.850 79.740 ;
        RECT 82.880 79.880 83.170 79.925 ;
        RECT 83.370 79.880 83.690 79.940 ;
        RECT 82.880 79.740 83.690 79.880 ;
        RECT 82.880 79.695 83.170 79.740 ;
        RECT 83.370 79.680 83.690 79.740 ;
        RECT 70.030 79.400 74.860 79.540 ;
        RECT 70.030 79.340 70.350 79.400 ;
        RECT 79.230 79.340 79.550 79.600 ;
        RECT 81.085 79.540 81.375 79.585 ;
        RECT 85.670 79.540 85.990 79.600 ;
        RECT 81.085 79.400 85.990 79.540 ;
        RECT 81.085 79.355 81.375 79.400 ;
        RECT 85.670 79.340 85.990 79.400 ;
        RECT 13.380 78.720 92.040 79.200 ;
        RECT 22.650 78.320 22.970 78.580 ;
        RECT 35.530 78.320 35.850 78.580 ;
        RECT 46.110 78.520 46.430 78.580 ;
        RECT 46.585 78.520 46.875 78.565 ;
        RECT 46.110 78.380 46.875 78.520 ;
        RECT 46.110 78.320 46.430 78.380 ;
        RECT 46.585 78.335 46.875 78.380 ;
        RECT 47.505 78.520 47.795 78.565 ;
        RECT 48.410 78.520 48.730 78.580 ;
        RECT 47.505 78.380 48.730 78.520 ;
        RECT 47.505 78.335 47.795 78.380 ;
        RECT 48.410 78.320 48.730 78.380 ;
        RECT 57.625 78.520 57.915 78.565 ;
        RECT 58.070 78.520 58.390 78.580 ;
        RECT 70.490 78.520 70.810 78.580 ;
        RECT 73.250 78.520 73.570 78.580 ;
        RECT 77.865 78.520 78.155 78.565 ;
        RECT 78.310 78.520 78.630 78.580 ;
        RECT 57.625 78.380 58.390 78.520 ;
        RECT 57.625 78.335 57.915 78.380 ;
        RECT 58.070 78.320 58.390 78.380 ;
        RECT 66.440 78.380 75.780 78.520 ;
        RECT 21.730 78.180 22.050 78.240 ;
        RECT 15.840 78.040 22.050 78.180 ;
        RECT 22.740 78.180 22.880 78.320 ;
        RECT 42.430 78.180 42.750 78.240 ;
        RECT 22.740 78.040 26.560 78.180 ;
        RECT 15.840 77.885 15.980 78.040 ;
        RECT 21.730 77.980 22.050 78.040 ;
        RECT 17.130 77.885 17.450 77.900 ;
        RECT 15.765 77.655 16.055 77.885 ;
        RECT 17.100 77.655 17.450 77.885 ;
        RECT 17.130 77.640 17.450 77.655 ;
        RECT 23.570 77.840 23.890 77.900 ;
        RECT 26.420 77.885 26.560 78.040 ;
        RECT 28.720 78.040 42.750 78.180 ;
        RECT 28.720 77.885 28.860 78.040 ;
        RECT 24.965 77.840 25.255 77.885 ;
        RECT 23.570 77.700 25.255 77.840 ;
        RECT 23.570 77.640 23.890 77.700 ;
        RECT 24.965 77.655 25.255 77.700 ;
        RECT 26.345 77.655 26.635 77.885 ;
        RECT 28.645 77.655 28.935 77.885 ;
        RECT 29.090 77.840 29.410 77.900 ;
        RECT 39.760 77.885 39.900 78.040 ;
        RECT 42.430 77.980 42.750 78.040 ;
        RECT 52.090 78.180 52.410 78.240 ;
        RECT 55.770 78.180 56.090 78.240 ;
        RECT 52.090 78.040 56.090 78.180 ;
        RECT 52.090 77.980 52.410 78.040 ;
        RECT 55.770 77.980 56.090 78.040 ;
        RECT 63.300 78.180 63.590 78.225 ;
        RECT 65.445 78.180 65.735 78.225 ;
        RECT 63.300 78.040 65.735 78.180 ;
        RECT 63.300 77.995 63.590 78.040 ;
        RECT 65.445 77.995 65.735 78.040 ;
        RECT 41.050 77.885 41.370 77.900 ;
        RECT 29.925 77.840 30.215 77.885 ;
        RECT 29.090 77.700 30.215 77.840 ;
        RECT 29.090 77.640 29.410 77.700 ;
        RECT 29.925 77.655 30.215 77.700 ;
        RECT 39.685 77.655 39.975 77.885 ;
        RECT 41.020 77.655 41.370 77.885 ;
        RECT 41.050 77.640 41.370 77.655 ;
        RECT 53.010 77.885 53.330 77.900 ;
        RECT 53.010 77.655 53.360 77.885 ;
        RECT 64.050 77.840 64.370 77.900 ;
        RECT 66.440 77.885 66.580 78.380 ;
        RECT 70.490 78.320 70.810 78.380 ;
        RECT 73.250 78.320 73.570 78.380 ;
        RECT 70.030 78.180 70.350 78.240 ;
        RECT 73.710 78.180 74.030 78.240 ;
        RECT 75.105 78.180 75.395 78.225 ;
        RECT 69.660 78.040 70.350 78.180 ;
        RECT 64.525 77.840 64.815 77.885 ;
        RECT 64.050 77.700 64.815 77.840 ;
        RECT 53.010 77.640 53.330 77.655 ;
        RECT 64.050 77.640 64.370 77.700 ;
        RECT 64.525 77.655 64.815 77.700 ;
        RECT 66.365 77.655 66.655 77.885 ;
        RECT 66.825 77.840 67.115 77.885 ;
        RECT 67.270 77.840 67.590 77.900 ;
        RECT 69.660 77.885 69.800 78.040 ;
        RECT 70.030 77.980 70.350 78.040 ;
        RECT 70.580 78.040 75.395 78.180 ;
        RECT 75.640 78.180 75.780 78.380 ;
        RECT 77.865 78.380 78.630 78.520 ;
        RECT 77.865 78.335 78.155 78.380 ;
        RECT 78.310 78.320 78.630 78.380 ;
        RECT 83.370 78.320 83.690 78.580 ;
        RECT 85.225 78.520 85.515 78.565 ;
        RECT 87.050 78.520 87.370 78.580 ;
        RECT 85.225 78.380 87.370 78.520 ;
        RECT 85.225 78.335 85.515 78.380 ;
        RECT 87.050 78.320 87.370 78.380 ;
        RECT 76.025 78.180 76.315 78.225 ;
        RECT 75.640 78.040 76.315 78.180 ;
        RECT 66.825 77.700 67.590 77.840 ;
        RECT 66.825 77.655 67.115 77.700 ;
        RECT 67.270 77.640 67.590 77.700 ;
        RECT 67.745 77.655 68.035 77.885 ;
        RECT 69.585 77.655 69.875 77.885 ;
        RECT 70.580 77.840 70.720 78.040 ;
        RECT 73.710 77.980 74.030 78.040 ;
        RECT 75.105 77.995 75.395 78.040 ;
        RECT 76.025 77.995 76.315 78.040 ;
        RECT 85.670 77.980 85.990 78.240 ;
        RECT 70.120 77.700 70.720 77.840 ;
        RECT 16.645 77.500 16.935 77.545 ;
        RECT 17.835 77.500 18.125 77.545 ;
        RECT 20.355 77.500 20.645 77.545 ;
        RECT 16.645 77.360 20.645 77.500 ;
        RECT 16.645 77.315 16.935 77.360 ;
        RECT 17.835 77.315 18.125 77.360 ;
        RECT 20.355 77.315 20.645 77.360 ;
        RECT 29.525 77.500 29.815 77.545 ;
        RECT 30.715 77.500 31.005 77.545 ;
        RECT 33.235 77.500 33.525 77.545 ;
        RECT 29.525 77.360 33.525 77.500 ;
        RECT 29.525 77.315 29.815 77.360 ;
        RECT 30.715 77.315 31.005 77.360 ;
        RECT 33.235 77.315 33.525 77.360 ;
        RECT 40.565 77.500 40.855 77.545 ;
        RECT 41.755 77.500 42.045 77.545 ;
        RECT 44.275 77.500 44.565 77.545 ;
        RECT 40.565 77.360 44.565 77.500 ;
        RECT 40.565 77.315 40.855 77.360 ;
        RECT 41.755 77.315 42.045 77.360 ;
        RECT 44.275 77.315 44.565 77.360 ;
        RECT 49.815 77.500 50.105 77.545 ;
        RECT 52.335 77.500 52.625 77.545 ;
        RECT 53.525 77.500 53.815 77.545 ;
        RECT 49.815 77.360 53.815 77.500 ;
        RECT 49.815 77.315 50.105 77.360 ;
        RECT 52.335 77.315 52.625 77.360 ;
        RECT 53.525 77.315 53.815 77.360 ;
        RECT 54.405 77.315 54.695 77.545 ;
        RECT 59.935 77.500 60.225 77.545 ;
        RECT 62.455 77.500 62.745 77.545 ;
        RECT 63.645 77.500 63.935 77.545 ;
        RECT 59.935 77.360 63.935 77.500 ;
        RECT 67.820 77.500 67.960 77.655 ;
        RECT 70.120 77.545 70.260 77.700 ;
        RECT 70.950 77.640 71.270 77.900 ;
        RECT 71.870 77.840 72.190 77.900 ;
        RECT 72.805 77.840 73.095 77.885 ;
        RECT 71.870 77.700 73.095 77.840 ;
        RECT 71.870 77.640 72.190 77.700 ;
        RECT 72.805 77.655 73.095 77.700 ;
        RECT 68.665 77.500 68.955 77.545 ;
        RECT 67.820 77.360 68.955 77.500 ;
        RECT 59.935 77.315 60.225 77.360 ;
        RECT 62.455 77.315 62.745 77.360 ;
        RECT 63.645 77.315 63.935 77.360 ;
        RECT 68.665 77.315 68.955 77.360 ;
        RECT 70.045 77.315 70.335 77.545 ;
        RECT 70.490 77.500 70.810 77.560 ;
        RECT 71.410 77.500 71.730 77.560 ;
        RECT 70.490 77.360 71.730 77.500 ;
        RECT 72.880 77.500 73.020 77.655 ;
        RECT 74.170 77.640 74.490 77.900 ;
        RECT 75.565 77.655 75.855 77.885 ;
        RECT 76.945 77.840 77.235 77.885 ;
        RECT 78.310 77.840 78.630 77.900 ;
        RECT 76.945 77.700 78.630 77.840 ;
        RECT 76.945 77.655 77.235 77.700 ;
        RECT 75.640 77.500 75.780 77.655 ;
        RECT 78.310 77.640 78.630 77.700 ;
        RECT 87.525 77.840 87.815 77.885 ;
        RECT 88.430 77.840 88.750 77.900 ;
        RECT 87.525 77.700 88.750 77.840 ;
        RECT 87.525 77.655 87.815 77.700 ;
        RECT 88.430 77.640 88.750 77.700 ;
        RECT 99.980 77.735 100.370 81.555 ;
        RECT 101.460 81.315 102.460 83.715 ;
        RECT 102.950 81.585 103.950 83.735 ;
        RECT 101.210 81.085 102.460 81.315 ;
        RECT 100.650 80.925 102.460 81.085 ;
        RECT 102.720 80.945 103.950 81.585 ;
        RECT 104.430 81.575 105.430 83.725 ;
        RECT 105.890 81.575 106.890 83.715 ;
        RECT 100.650 80.625 101.930 80.925 ;
        RECT 100.650 78.745 101.650 80.625 ;
        RECT 102.720 80.475 103.400 80.945 ;
        RECT 104.210 80.935 105.430 81.575 ;
        RECT 104.210 80.475 104.890 80.935 ;
        RECT 105.700 80.925 106.890 81.575 ;
        RECT 107.390 81.545 108.390 83.735 ;
        RECT 110.330 83.715 112.640 83.725 ;
        RECT 107.150 80.945 108.390 81.545 ;
        RECT 108.900 81.535 109.900 83.715 ;
        RECT 110.330 81.545 112.810 83.715 ;
        RECT 105.700 80.475 106.380 80.925 ;
        RECT 107.150 80.475 107.830 80.945 ;
        RECT 102.100 80.005 103.400 80.475 ;
        RECT 102.100 78.835 103.140 80.005 ;
        RECT 103.610 79.995 104.890 80.475 ;
        RECT 105.080 79.995 106.380 80.475 ;
        RECT 103.610 78.835 104.650 79.995 ;
        RECT 105.080 78.835 106.120 79.995 ;
        RECT 106.570 79.965 107.830 80.475 ;
        RECT 108.650 80.925 109.900 81.535 ;
        RECT 110.160 80.935 112.810 81.545 ;
        RECT 108.650 80.465 109.330 80.925 ;
        RECT 110.160 80.475 110.840 80.935 ;
        RECT 111.810 80.925 112.810 80.935 ;
        RECT 100.650 78.295 101.880 78.745 ;
        RECT 102.100 78.295 103.430 78.835 ;
        RECT 103.610 78.295 104.920 78.835 ;
        RECT 105.080 78.295 106.410 78.835 ;
        RECT 106.570 78.825 107.610 79.965 ;
        RECT 108.050 79.955 109.330 80.465 ;
        RECT 109.530 79.965 110.840 80.475 ;
        RECT 108.050 78.825 109.090 79.955 ;
        RECT 106.570 78.295 107.840 78.825 ;
        RECT 101.200 77.735 101.880 78.295 ;
        RECT 102.750 77.745 103.430 78.295 ;
        RECT 104.240 77.755 104.920 78.295 ;
        RECT 105.730 77.755 106.410 78.295 ;
        RECT 107.160 77.755 107.840 78.295 ;
        RECT 108.050 78.285 109.350 78.825 ;
        RECT 109.530 78.295 110.570 79.965 ;
        RECT 108.670 77.755 109.350 78.285 ;
        RECT 79.690 77.500 80.010 77.560 ;
        RECT 72.880 77.360 80.010 77.500 ;
        RECT 16.250 77.160 16.540 77.205 ;
        RECT 18.350 77.160 18.640 77.205 ;
        RECT 19.920 77.160 20.210 77.205 ;
        RECT 16.250 77.020 20.210 77.160 ;
        RECT 16.250 76.975 16.540 77.020 ;
        RECT 18.350 76.975 18.640 77.020 ;
        RECT 19.920 76.975 20.210 77.020 ;
        RECT 24.950 77.160 25.270 77.220 ;
        RECT 27.725 77.160 28.015 77.205 ;
        RECT 24.950 77.020 28.015 77.160 ;
        RECT 24.950 76.960 25.270 77.020 ;
        RECT 27.725 76.975 28.015 77.020 ;
        RECT 29.130 77.160 29.420 77.205 ;
        RECT 31.230 77.160 31.520 77.205 ;
        RECT 32.800 77.160 33.090 77.205 ;
        RECT 29.130 77.020 33.090 77.160 ;
        RECT 29.130 76.975 29.420 77.020 ;
        RECT 31.230 76.975 31.520 77.020 ;
        RECT 32.800 76.975 33.090 77.020 ;
        RECT 40.170 77.160 40.460 77.205 ;
        RECT 42.270 77.160 42.560 77.205 ;
        RECT 43.840 77.160 44.130 77.205 ;
        RECT 40.170 77.020 44.130 77.160 ;
        RECT 40.170 76.975 40.460 77.020 ;
        RECT 42.270 76.975 42.560 77.020 ;
        RECT 43.840 76.975 44.130 77.020 ;
        RECT 50.250 77.160 50.540 77.205 ;
        RECT 51.820 77.160 52.110 77.205 ;
        RECT 53.920 77.160 54.210 77.205 ;
        RECT 50.250 77.020 54.210 77.160 ;
        RECT 50.250 76.975 50.540 77.020 ;
        RECT 51.820 76.975 52.110 77.020 ;
        RECT 53.920 76.975 54.210 77.020 ;
        RECT 25.410 76.620 25.730 76.880 ;
        RECT 52.550 76.820 52.870 76.880 ;
        RECT 54.480 76.820 54.620 77.315 ;
        RECT 70.490 77.300 70.810 77.360 ;
        RECT 71.410 77.300 71.730 77.360 ;
        RECT 79.690 77.300 80.010 77.360 ;
        RECT 86.130 77.300 86.450 77.560 ;
        RECT 60.370 77.160 60.660 77.205 ;
        RECT 61.940 77.160 62.230 77.205 ;
        RECT 64.040 77.160 64.330 77.205 ;
        RECT 60.370 77.020 64.330 77.160 ;
        RECT 60.370 76.975 60.660 77.020 ;
        RECT 61.940 76.975 62.230 77.020 ;
        RECT 64.040 76.975 64.330 77.020 ;
        RECT 67.270 76.960 67.590 77.220 ;
        RECT 74.170 77.160 74.490 77.220 ;
        RECT 75.550 77.160 75.870 77.220 ;
        RECT 74.170 77.020 75.870 77.160 ;
        RECT 74.170 76.960 74.490 77.020 ;
        RECT 75.550 76.960 75.870 77.020 ;
        RECT 52.550 76.680 54.620 76.820 ;
        RECT 88.445 76.820 88.735 76.865 ;
        RECT 88.890 76.820 89.210 76.880 ;
        RECT 88.445 76.680 89.210 76.820 ;
        RECT 52.550 76.620 52.870 76.680 ;
        RECT 88.445 76.635 88.735 76.680 ;
        RECT 88.890 76.620 89.210 76.680 ;
        RECT 13.380 76.000 92.040 76.480 ;
        RECT 16.685 75.800 16.975 75.845 ;
        RECT 17.130 75.800 17.450 75.860 ;
        RECT 16.685 75.660 17.450 75.800 ;
        RECT 16.685 75.615 16.975 75.660 ;
        RECT 17.130 75.600 17.450 75.660 ;
        RECT 21.285 75.800 21.575 75.845 ;
        RECT 22.650 75.800 22.970 75.860 ;
        RECT 21.285 75.660 22.970 75.800 ;
        RECT 21.285 75.615 21.575 75.660 ;
        RECT 22.650 75.600 22.970 75.660 ;
        RECT 23.570 75.600 23.890 75.860 ;
        RECT 41.050 75.800 41.370 75.860 ;
        RECT 42.445 75.800 42.735 75.845 ;
        RECT 52.090 75.800 52.410 75.860 ;
        RECT 41.050 75.660 42.735 75.800 ;
        RECT 41.050 75.600 41.370 75.660 ;
        RECT 42.445 75.615 42.735 75.660 ;
        RECT 45.280 75.660 52.410 75.800 ;
        RECT 19.445 75.460 19.735 75.505 ;
        RECT 23.660 75.460 23.800 75.600 ;
        RECT 19.445 75.320 23.800 75.460 ;
        RECT 29.590 75.460 29.880 75.505 ;
        RECT 31.690 75.460 31.980 75.505 ;
        RECT 33.260 75.460 33.550 75.505 ;
        RECT 29.590 75.320 33.550 75.460 ;
        RECT 19.445 75.275 19.735 75.320 ;
        RECT 29.590 75.275 29.880 75.320 ;
        RECT 31.690 75.275 31.980 75.320 ;
        RECT 33.260 75.275 33.550 75.320 ;
        RECT 41.970 75.460 42.290 75.520 ;
        RECT 45.280 75.460 45.420 75.660 ;
        RECT 52.090 75.600 52.410 75.660 ;
        RECT 52.565 75.800 52.855 75.845 ;
        RECT 53.010 75.800 53.330 75.860 ;
        RECT 52.565 75.660 53.330 75.800 ;
        RECT 52.565 75.615 52.855 75.660 ;
        RECT 53.010 75.600 53.330 75.660 ;
        RECT 57.165 75.800 57.455 75.845 ;
        RECT 72.790 75.800 73.110 75.860 ;
        RECT 73.265 75.800 73.555 75.845 ;
        RECT 76.470 75.800 76.790 75.860 ;
        RECT 57.165 75.660 64.740 75.800 ;
        RECT 57.165 75.615 57.455 75.660 ;
        RECT 57.240 75.460 57.380 75.615 ;
        RECT 41.970 75.320 45.420 75.460 ;
        RECT 41.970 75.260 42.290 75.320 ;
        RECT 18.050 75.120 18.370 75.180 ;
        RECT 21.270 75.120 21.590 75.180 ;
        RECT 17.680 74.980 21.590 75.120 ;
        RECT 17.680 74.825 17.820 74.980 ;
        RECT 18.050 74.920 18.370 74.980 ;
        RECT 21.270 74.920 21.590 74.980 ;
        RECT 29.985 75.120 30.275 75.165 ;
        RECT 31.175 75.120 31.465 75.165 ;
        RECT 33.695 75.120 33.985 75.165 ;
        RECT 29.985 74.980 33.985 75.120 ;
        RECT 29.985 74.935 30.275 74.980 ;
        RECT 31.175 74.935 31.465 74.980 ;
        RECT 33.695 74.935 33.985 74.980 ;
        RECT 44.730 74.920 45.050 75.180 ;
        RECT 45.280 75.165 45.420 75.320 ;
        RECT 48.960 75.320 57.380 75.460 ;
        RECT 59.910 75.460 60.200 75.505 ;
        RECT 61.480 75.460 61.770 75.505 ;
        RECT 63.580 75.460 63.870 75.505 ;
        RECT 59.910 75.320 63.870 75.460 ;
        RECT 48.960 75.165 49.100 75.320 ;
        RECT 59.910 75.275 60.200 75.320 ;
        RECT 61.480 75.275 61.770 75.320 ;
        RECT 63.580 75.275 63.870 75.320 ;
        RECT 45.205 74.935 45.495 75.165 ;
        RECT 48.885 74.935 49.175 75.165 ;
        RECT 49.345 74.935 49.635 75.165 ;
        RECT 51.630 75.120 51.950 75.180 ;
        RECT 54.865 75.120 55.155 75.165 ;
        RECT 51.630 74.980 55.155 75.120 ;
        RECT 17.605 74.595 17.895 74.825 ;
        RECT 18.510 74.580 18.830 74.840 ;
        RECT 22.650 74.780 22.970 74.840 ;
        RECT 23.125 74.780 23.415 74.825 ;
        RECT 22.650 74.640 23.415 74.780 ;
        RECT 22.650 74.580 22.970 74.640 ;
        RECT 23.125 74.595 23.415 74.640 ;
        RECT 24.965 74.780 25.255 74.825 ;
        RECT 25.410 74.780 25.730 74.840 ;
        RECT 24.965 74.640 25.730 74.780 ;
        RECT 24.965 74.595 25.255 74.640 ;
        RECT 25.410 74.580 25.730 74.640 ;
        RECT 29.105 74.780 29.395 74.825 ;
        RECT 41.525 74.780 41.815 74.825 ;
        RECT 42.430 74.780 42.750 74.840 ;
        RECT 29.105 74.640 42.750 74.780 ;
        RECT 29.105 74.595 29.395 74.640 ;
        RECT 41.525 74.595 41.815 74.640 ;
        RECT 42.430 74.580 42.750 74.640 ;
        RECT 47.490 74.780 47.810 74.840 ;
        RECT 49.420 74.780 49.560 74.935 ;
        RECT 51.630 74.920 51.950 74.980 ;
        RECT 54.865 74.935 55.155 74.980 ;
        RECT 55.770 74.920 56.090 75.180 ;
        RECT 64.600 75.165 64.740 75.660 ;
        RECT 72.790 75.660 76.790 75.800 ;
        RECT 72.790 75.600 73.110 75.660 ;
        RECT 73.265 75.615 73.555 75.660 ;
        RECT 76.470 75.600 76.790 75.660 ;
        RECT 88.430 75.600 88.750 75.860 ;
        RECT 99.980 75.585 101.000 77.735 ;
        RECT 101.200 77.165 102.510 77.735 ;
        RECT 102.750 77.255 103.960 77.745 ;
        RECT 104.240 77.255 105.470 77.755 ;
        RECT 105.730 77.255 106.940 77.755 ;
        RECT 101.470 75.575 102.510 77.165 ;
        RECT 102.920 75.565 103.960 77.255 ;
        RECT 104.430 75.575 105.470 77.255 ;
        RECT 105.900 75.575 106.940 77.255 ;
        RECT 107.160 77.245 108.430 77.755 ;
        RECT 108.670 77.245 109.900 77.755 ;
        RECT 107.390 75.575 108.430 77.245 ;
        RECT 108.860 75.575 109.900 77.245 ;
        RECT 116.265 75.625 117.170 87.645 ;
        RECT 118.030 84.370 118.360 91.480 ;
        RECT 118.020 83.515 118.360 84.370 ;
        RECT 118.020 83.510 118.340 83.515 ;
        RECT 118.020 82.930 118.260 83.510 ;
        RECT 118.670 83.310 119.140 91.720 ;
        RECT 119.640 91.515 119.860 92.280 ;
        RECT 120.840 91.720 122.800 91.950 ;
        RECT 124.270 91.720 126.230 91.950 ;
        RECT 127.700 91.720 128.660 91.950 ;
        RECT 119.420 91.310 119.860 91.515 ;
        RECT 120.560 91.490 120.790 91.515 ;
        RECT 120.560 91.480 120.800 91.490 ;
        RECT 119.420 83.570 119.810 91.310 ;
        RECT 120.390 84.420 120.800 91.480 ;
        RECT 121.380 85.130 122.280 91.720 ;
        RECT 122.850 91.470 123.080 91.515 ;
        RECT 123.990 91.490 124.220 91.515 ;
        RECT 120.380 83.600 120.800 84.420 ;
        RECT 121.350 84.120 122.350 85.130 ;
        RECT 119.420 83.515 119.650 83.570 ;
        RECT 120.380 83.515 120.790 83.600 ;
        RECT 118.410 83.080 119.370 83.310 ;
        RECT 118.020 82.440 118.340 82.930 ;
        RECT 117.580 81.190 118.420 82.440 ;
        RECT 118.020 80.140 118.260 81.190 ;
        RECT 118.560 80.530 119.230 83.080 ;
        RECT 120.380 81.300 120.700 83.515 ;
        RECT 121.380 83.310 122.280 84.120 ;
        RECT 122.850 83.580 123.370 91.470 ;
        RECT 122.850 83.515 123.080 83.580 ;
        RECT 123.850 83.570 124.230 91.490 ;
        RECT 124.930 85.090 125.750 91.720 ;
        RECT 126.280 91.470 126.510 91.515 ;
        RECT 127.420 91.470 127.650 91.515 ;
        RECT 124.840 84.090 125.840 85.090 ;
        RECT 123.860 83.515 124.220 83.570 ;
        RECT 120.840 83.080 122.800 83.310 ;
        RECT 123.860 81.950 124.120 83.515 ;
        RECT 124.930 83.310 125.750 84.090 ;
        RECT 126.280 83.600 127.660 91.470 ;
        RECT 128.010 91.350 128.430 91.720 ;
        RECT 128.710 91.470 128.940 91.515 ;
        RECT 129.340 91.470 130.480 92.280 ;
        RECT 128.710 87.490 130.480 91.470 ;
        RECT 128.710 86.490 130.470 87.490 ;
        RECT 128.710 85.550 130.480 86.490 ;
        RECT 134.410 85.550 139.730 85.560 ;
        RECT 128.710 84.950 139.730 85.550 ;
        RECT 128.710 84.870 136.330 84.950 ;
        RECT 128.710 84.550 136.160 84.870 ;
        RECT 126.280 83.515 126.510 83.600 ;
        RECT 127.420 83.515 127.650 83.600 ;
        RECT 128.010 83.310 128.430 83.980 ;
        RECT 128.710 83.610 130.480 84.550 ;
        RECT 128.710 83.515 128.940 83.610 ;
        RECT 124.270 83.080 126.230 83.310 ;
        RECT 127.700 83.080 128.660 83.310 ;
        RECT 127.800 82.200 128.590 83.080 ;
        RECT 129.340 82.600 130.480 83.610 ;
        RECT 123.860 81.330 127.480 81.950 ;
        RECT 127.750 81.440 128.640 82.200 ;
        RECT 118.420 80.300 119.380 80.530 ;
        RECT 118.020 79.130 118.370 80.140 ;
        RECT 118.030 76.180 118.370 79.130 ;
        RECT 118.140 76.140 118.370 76.180 ;
        RECT 118.670 75.980 119.110 80.300 ;
        RECT 120.380 80.140 120.710 81.300 ;
        RECT 120.850 80.300 122.810 80.530 ;
        RECT 119.430 80.130 119.660 80.140 ;
        RECT 119.430 77.820 119.840 80.130 ;
        RECT 120.380 80.100 120.800 80.140 ;
        RECT 121.160 80.100 122.500 80.300 ;
        RECT 123.860 80.140 124.120 81.330 ;
        RECT 127.070 80.680 127.470 81.330 ;
        RECT 129.410 81.250 130.480 82.600 ;
        RECT 134.410 84.540 136.160 84.550 ;
        RECT 134.410 83.750 134.760 84.540 ;
        RECT 136.910 84.520 139.710 84.770 ;
        RECT 135.150 84.300 135.440 84.330 ;
        RECT 135.140 84.050 135.460 84.300 ;
        RECT 136.910 83.895 137.070 84.520 ;
        RECT 137.210 84.050 137.540 84.380 ;
        RECT 137.820 84.250 138.030 84.520 ;
        RECT 137.890 83.910 138.030 84.250 ;
        RECT 138.170 84.050 138.500 84.380 ;
        RECT 138.970 84.040 139.710 84.520 ;
        RECT 137.890 83.895 138.180 83.910 ;
        RECT 138.970 83.895 139.140 84.040 ;
        RECT 139.320 83.960 139.710 84.040 ;
        RECT 134.960 83.750 135.190 83.895 ;
        RECT 129.410 80.820 131.250 81.250 ;
        RECT 129.410 80.780 130.470 80.820 ;
        RECT 128.470 80.680 129.220 80.690 ;
        RECT 127.070 80.630 129.220 80.680 ;
        RECT 127.070 80.590 129.400 80.630 ;
        RECT 124.280 80.300 126.240 80.530 ;
        RECT 127.070 80.340 130.630 80.590 ;
        RECT 127.070 80.330 128.410 80.340 ;
        RECT 128.120 80.310 128.410 80.330 ;
        RECT 120.380 79.170 122.500 80.100 ;
        RECT 119.430 76.140 119.930 77.820 ;
        RECT 120.500 76.200 122.500 79.170 ;
        RECT 120.570 76.140 120.800 76.200 ;
        RECT 118.420 75.750 119.380 75.980 ;
        RECT 116.265 75.520 118.010 75.625 ;
        RECT 119.730 75.520 119.930 76.140 ;
        RECT 121.160 75.980 122.500 76.200 ;
        RECT 122.860 80.090 123.090 80.140 ;
        RECT 123.860 80.090 124.230 80.140 ;
        RECT 124.570 80.090 125.940 80.300 ;
        RECT 129.280 80.250 130.630 80.340 ;
        RECT 130.230 80.245 130.520 80.250 ;
        RECT 122.860 77.870 123.310 80.090 ;
        RECT 123.860 79.800 125.940 80.090 ;
        RECT 122.860 77.380 123.360 77.870 ;
        RECT 122.860 76.710 123.450 77.380 ;
        RECT 122.860 76.460 123.510 76.710 ;
        RECT 122.860 76.430 123.560 76.460 ;
        RECT 122.860 76.140 123.090 76.430 ;
        RECT 123.320 76.060 123.560 76.430 ;
        RECT 123.870 76.200 125.940 79.800 ;
        RECT 123.870 76.180 124.230 76.200 ;
        RECT 124.000 76.140 124.230 76.180 ;
        RECT 120.850 75.750 122.810 75.980 ;
        RECT 123.240 75.820 123.560 76.060 ;
        RECT 124.570 75.980 125.940 76.200 ;
        RECT 126.290 79.960 126.520 80.140 ;
        RECT 127.930 80.090 128.160 80.150 ;
        RECT 128.370 80.090 128.600 80.150 ;
        RECT 127.180 80.080 128.160 80.090 ;
        RECT 126.750 79.960 128.160 80.080 ;
        RECT 126.290 79.210 128.160 79.960 ;
        RECT 128.350 79.950 128.750 80.090 ;
        RECT 130.040 79.950 130.270 80.040 ;
        RECT 130.480 79.990 130.710 80.040 ;
        RECT 130.880 79.990 131.250 80.820 ;
        RECT 128.350 79.220 130.310 79.950 ;
        RECT 128.350 79.210 128.750 79.220 ;
        RECT 126.290 78.750 127.650 79.210 ;
        RECT 127.930 79.150 128.160 79.210 ;
        RECT 128.370 79.150 128.600 79.210 ;
        RECT 126.290 78.480 128.750 78.750 ;
        RECT 126.290 78.440 128.460 78.480 ;
        RECT 126.290 76.690 127.640 78.440 ;
        RECT 128.920 78.260 130.300 79.220 ;
        RECT 128.920 78.130 130.320 78.260 ;
        RECT 128.200 77.130 130.320 78.130 ;
        RECT 128.920 77.100 130.320 77.130 ;
        RECT 130.040 77.090 130.320 77.100 ;
        RECT 130.480 77.130 131.250 79.990 ;
        RECT 134.410 79.895 135.190 83.750 ;
        RECT 135.400 83.840 135.630 83.895 ;
        RECT 135.400 80.660 136.040 83.840 ;
        RECT 135.400 79.950 136.050 80.660 ;
        RECT 136.540 80.130 136.770 83.895 ;
        RECT 136.910 83.750 137.250 83.895 ;
        RECT 135.400 79.895 135.630 79.950 ;
        RECT 134.410 79.880 135.160 79.895 ;
        RECT 134.410 79.870 134.760 79.880 ;
        RECT 135.150 79.590 135.440 79.690 ;
        RECT 134.910 79.080 135.590 79.590 ;
        RECT 134.410 78.080 135.590 79.080 ;
        RECT 134.910 77.590 135.590 78.080 ;
        RECT 135.140 77.550 135.430 77.590 ;
        RECT 134.950 77.340 135.180 77.390 ;
        RECT 130.040 77.040 130.270 77.090 ;
        RECT 130.480 77.040 130.710 77.130 ;
        RECT 130.880 77.100 131.250 77.130 ;
        RECT 126.290 76.390 128.990 76.690 ;
        RECT 126.290 76.140 126.520 76.390 ;
        RECT 123.200 75.520 123.560 75.820 ;
        RECT 124.280 75.750 126.240 75.980 ;
        RECT 126.900 75.550 128.990 76.390 ;
        RECT 134.410 76.460 135.180 77.340 ;
        RECT 134.410 76.240 134.810 76.460 ;
        RECT 134.950 76.390 135.180 76.460 ;
        RECT 135.390 77.330 135.620 77.390 ;
        RECT 135.830 77.330 136.050 79.950 ;
        RECT 136.330 79.895 136.770 80.130 ;
        RECT 137.020 79.895 137.250 83.750 ;
        RECT 137.500 80.070 137.730 83.895 ;
        RECT 137.890 83.760 138.210 83.895 ;
        RECT 137.390 79.895 137.730 80.070 ;
        RECT 137.980 79.895 138.210 83.760 ;
        RECT 138.460 80.090 138.690 83.895 ;
        RECT 138.380 80.040 138.690 80.090 ;
        RECT 138.350 79.895 138.690 80.040 ;
        RECT 138.940 79.895 139.170 83.895 ;
        RECT 136.330 79.880 136.620 79.895 ;
        RECT 137.390 79.890 137.600 79.895 ;
        RECT 138.350 79.890 138.550 79.895 ;
        RECT 136.330 79.200 136.590 79.880 ;
        RECT 136.730 79.410 137.060 79.740 ;
        RECT 137.390 79.230 137.550 79.890 ;
        RECT 137.690 79.410 138.020 79.740 ;
        RECT 138.350 79.260 138.510 79.890 ;
        RECT 138.650 79.410 138.980 79.740 ;
        RECT 136.330 79.190 136.620 79.200 ;
        RECT 137.390 79.190 137.600 79.230 ;
        RECT 138.350 79.190 138.550 79.260 ;
        RECT 136.330 79.050 138.550 79.190 ;
        RECT 139.410 79.140 139.700 83.960 ;
        RECT 135.390 77.050 136.050 77.330 ;
        RECT 136.320 79.020 138.550 79.050 ;
        RECT 136.320 78.540 138.520 79.020 ;
        RECT 136.320 78.190 138.790 78.540 ;
        RECT 136.320 78.100 138.800 78.190 ;
        RECT 138.940 78.140 139.940 79.140 ;
        RECT 136.320 77.390 136.730 78.100 ;
        RECT 137.200 77.550 137.530 77.880 ;
        RECT 137.680 77.530 137.850 78.100 ;
        RECT 138.470 78.090 138.800 78.100 ;
        RECT 138.160 77.550 138.490 77.880 ;
        RECT 138.650 77.530 138.800 78.090 ;
        RECT 137.680 77.390 137.820 77.530 ;
        RECT 138.650 77.390 138.790 77.530 ;
        RECT 136.320 77.150 136.760 77.390 ;
        RECT 135.390 76.450 136.020 77.050 ;
        RECT 135.390 76.390 135.620 76.450 ;
        RECT 136.530 76.390 136.760 77.150 ;
        RECT 137.010 76.560 137.240 77.390 ;
        RECT 137.490 77.160 137.820 77.390 ;
        RECT 137.010 76.390 137.340 76.560 ;
        RECT 137.490 76.390 137.720 77.160 ;
        RECT 137.970 76.620 138.200 77.390 ;
        RECT 138.450 77.170 138.790 77.390 ;
        RECT 138.930 77.310 139.160 77.390 ;
        RECT 139.410 77.310 139.700 78.140 ;
        RECT 137.970 76.390 138.310 76.620 ;
        RECT 138.450 76.390 138.680 77.170 ;
        RECT 138.930 76.390 139.700 77.310 ;
        RECT 134.410 75.700 134.900 76.240 ;
        RECT 135.110 76.020 135.460 76.230 ;
        RECT 135.120 75.960 135.460 76.020 ;
        RECT 136.720 75.910 137.050 76.240 ;
        RECT 137.200 75.750 137.340 76.390 ;
        RECT 138.150 76.240 138.310 76.390 ;
        RECT 137.680 75.910 138.010 76.240 ;
        RECT 138.150 75.750 138.320 76.240 ;
        RECT 138.640 75.910 138.970 76.240 ;
        RECT 139.110 75.750 139.700 76.390 ;
        RECT 134.410 75.680 135.410 75.700 ;
        RECT 134.410 75.550 136.210 75.680 ;
        RECT 126.900 75.520 136.210 75.550 ;
        RECT 67.270 75.460 67.590 75.520 ;
        RECT 82.030 75.460 82.320 75.505 ;
        RECT 84.130 75.460 84.420 75.505 ;
        RECT 85.700 75.460 85.990 75.505 ;
        RECT 67.270 75.320 71.180 75.460 ;
        RECT 67.270 75.260 67.590 75.320 ;
        RECT 59.475 75.120 59.765 75.165 ;
        RECT 61.995 75.120 62.285 75.165 ;
        RECT 63.185 75.120 63.475 75.165 ;
        RECT 59.475 74.980 63.475 75.120 ;
        RECT 59.475 74.935 59.765 74.980 ;
        RECT 61.995 74.935 62.285 74.980 ;
        RECT 63.185 74.935 63.475 74.980 ;
        RECT 64.525 74.935 64.815 75.165 ;
        RECT 67.745 75.120 68.035 75.165 ;
        RECT 67.745 74.980 69.800 75.120 ;
        RECT 67.745 74.935 68.035 74.980 ;
        RECT 47.490 74.640 49.560 74.780 ;
        RECT 52.550 74.780 52.870 74.840 ;
        RECT 57.150 74.780 57.470 74.840 ;
        RECT 64.050 74.780 64.370 74.840 ;
        RECT 52.550 74.640 64.370 74.780 ;
        RECT 47.490 74.580 47.810 74.640 ;
        RECT 52.550 74.580 52.870 74.640 ;
        RECT 57.150 74.580 57.470 74.640 ;
        RECT 64.050 74.580 64.370 74.640 ;
        RECT 65.890 74.780 66.210 74.840 ;
        RECT 69.110 74.780 69.430 74.840 ;
        RECT 69.660 74.825 69.800 74.980 ;
        RECT 70.490 74.920 70.810 75.180 ;
        RECT 71.040 74.825 71.180 75.320 ;
        RECT 82.030 75.320 85.990 75.460 ;
        RECT 82.030 75.275 82.320 75.320 ;
        RECT 84.130 75.275 84.420 75.320 ;
        RECT 85.700 75.275 85.990 75.320 ;
        RECT 116.265 75.250 136.210 75.520 ;
        RECT 136.430 75.550 139.700 75.750 ;
        RECT 136.430 75.540 139.260 75.550 ;
        RECT 136.430 75.390 139.180 75.540 ;
        RECT 139.440 75.250 139.700 75.290 ;
        RECT 71.410 75.120 71.730 75.180 ;
        RECT 73.250 75.120 73.570 75.180 ;
        RECT 71.410 74.980 73.570 75.120 ;
        RECT 71.410 74.920 71.730 74.980 ;
        RECT 73.250 74.920 73.570 74.980 ;
        RECT 76.930 75.120 77.250 75.180 ;
        RECT 78.770 75.120 79.090 75.180 ;
        RECT 76.930 74.980 79.090 75.120 ;
        RECT 76.930 74.920 77.250 74.980 ;
        RECT 78.770 74.920 79.090 74.980 ;
        RECT 80.610 75.120 80.930 75.180 ;
        RECT 81.530 75.120 81.850 75.180 ;
        RECT 80.610 74.980 81.850 75.120 ;
        RECT 80.610 74.920 80.930 74.980 ;
        RECT 81.530 74.920 81.850 74.980 ;
        RECT 82.425 75.120 82.715 75.165 ;
        RECT 83.615 75.120 83.905 75.165 ;
        RECT 86.135 75.120 86.425 75.165 ;
        RECT 82.425 74.980 86.425 75.120 ;
        RECT 82.425 74.935 82.715 74.980 ;
        RECT 83.615 74.935 83.905 74.980 ;
        RECT 86.135 74.935 86.425 74.980 ;
        RECT 65.890 74.640 69.430 74.780 ;
        RECT 65.890 74.580 66.210 74.640 ;
        RECT 69.110 74.580 69.430 74.640 ;
        RECT 69.585 74.595 69.875 74.825 ;
        RECT 70.965 74.595 71.255 74.825 ;
        RECT 72.330 74.580 72.650 74.840 ;
        RECT 73.340 74.780 73.480 74.920 ;
        RECT 116.265 74.910 139.700 75.250 ;
        RECT 73.725 74.780 74.015 74.825 ;
        RECT 73.340 74.640 74.015 74.780 ;
        RECT 73.725 74.595 74.015 74.640 ;
        RECT 74.630 74.580 74.950 74.840 ;
        RECT 75.090 74.780 75.410 74.840 ;
        RECT 75.565 74.780 75.855 74.825 ;
        RECT 87.970 74.780 88.290 74.840 ;
        RECT 75.090 74.640 88.290 74.780 ;
        RECT 75.090 74.580 75.410 74.640 ;
        RECT 75.565 74.595 75.855 74.640 ;
        RECT 87.970 74.580 88.290 74.640 ;
        RECT 88.890 74.580 89.210 74.840 ;
        RECT 116.265 74.770 128.990 74.910 ;
        RECT 116.265 74.720 128.980 74.770 ;
        RECT 117.600 74.690 128.980 74.720 ;
        RECT 134.410 74.700 139.700 74.910 ;
        RECT 134.420 74.690 139.700 74.700 ;
        RECT 20.810 74.440 21.130 74.500 ;
        RECT 21.285 74.440 21.575 74.485 ;
        RECT 20.810 74.300 21.575 74.440 ;
        RECT 20.810 74.240 21.130 74.300 ;
        RECT 21.285 74.255 21.575 74.300 ;
        RECT 28.170 74.440 28.490 74.500 ;
        RECT 30.330 74.440 30.620 74.485 ;
        RECT 37.830 74.440 38.150 74.500 ;
        RECT 62.840 74.440 63.130 74.485 ;
        RECT 68.205 74.440 68.495 74.485 ;
        RECT 28.170 74.300 30.620 74.440 ;
        RECT 28.170 74.240 28.490 74.300 ;
        RECT 30.330 74.255 30.620 74.300 ;
        RECT 36.080 74.300 56.230 74.440 ;
        RECT 22.190 73.900 22.510 74.160 ;
        RECT 25.870 73.900 26.190 74.160 ;
        RECT 36.080 74.145 36.220 74.300 ;
        RECT 37.830 74.240 38.150 74.300 ;
        RECT 36.005 73.915 36.295 74.145 ;
        RECT 44.285 74.100 44.575 74.145 ;
        RECT 46.585 74.100 46.875 74.145 ;
        RECT 44.285 73.960 46.875 74.100 ;
        RECT 44.285 73.915 44.575 73.960 ;
        RECT 46.585 73.915 46.875 73.960 ;
        RECT 48.410 73.900 48.730 74.160 ;
        RECT 54.390 73.900 54.710 74.160 ;
        RECT 56.090 74.100 56.230 74.300 ;
        RECT 62.840 74.300 68.495 74.440 ;
        RECT 62.840 74.255 63.130 74.300 ;
        RECT 68.205 74.255 68.495 74.300 ;
        RECT 70.490 74.440 70.810 74.500 ;
        RECT 73.250 74.440 73.570 74.500 ;
        RECT 81.070 74.440 81.390 74.500 ;
        RECT 82.910 74.485 83.230 74.500 ;
        RECT 70.490 74.300 73.570 74.440 ;
        RECT 70.490 74.240 70.810 74.300 ;
        RECT 73.250 74.240 73.570 74.300 ;
        RECT 74.260 74.300 81.390 74.440 ;
        RECT 74.260 74.160 74.400 74.300 ;
        RECT 81.070 74.240 81.390 74.300 ;
        RECT 82.880 74.255 83.230 74.485 ;
        RECT 82.910 74.240 83.230 74.255 ;
        RECT 73.710 74.100 74.030 74.160 ;
        RECT 56.090 73.960 74.030 74.100 ;
        RECT 73.710 73.900 74.030 73.960 ;
        RECT 74.170 73.900 74.490 74.160 ;
        RECT 75.550 74.100 75.870 74.160 ;
        RECT 76.485 74.100 76.775 74.145 ;
        RECT 81.990 74.100 82.310 74.160 ;
        RECT 75.550 73.960 82.310 74.100 ;
        RECT 75.550 73.900 75.870 73.960 ;
        RECT 76.485 73.915 76.775 73.960 ;
        RECT 81.990 73.900 82.310 73.960 ;
        RECT 89.810 73.900 90.130 74.160 ;
        RECT 13.380 73.280 92.040 73.760 ;
        RECT 17.605 73.080 17.895 73.125 ;
        RECT 22.650 73.080 22.970 73.140 ;
        RECT 26.345 73.080 26.635 73.125 ;
        RECT 27.710 73.080 28.030 73.140 ;
        RECT 17.605 72.940 28.030 73.080 ;
        RECT 17.605 72.895 17.895 72.940 ;
        RECT 22.650 72.880 22.970 72.940 ;
        RECT 26.345 72.895 26.635 72.940 ;
        RECT 27.710 72.880 28.030 72.940 ;
        RECT 28.170 72.880 28.490 73.140 ;
        RECT 58.990 73.080 59.310 73.140 ;
        RECT 40.680 72.940 59.310 73.080 ;
        RECT 21.730 72.740 22.050 72.800 ;
        RECT 26.790 72.740 27.110 72.800 ;
        RECT 32.325 72.740 32.615 72.785 ;
        RECT 21.730 72.600 32.615 72.740 ;
        RECT 21.730 72.540 22.050 72.600 ;
        RECT 26.790 72.540 27.110 72.600 ;
        RECT 32.325 72.555 32.615 72.600 ;
        RECT 39.670 72.740 39.990 72.800 ;
        RECT 40.680 72.785 40.820 72.940 ;
        RECT 58.990 72.880 59.310 72.940 ;
        RECT 67.270 73.080 67.590 73.140 ;
        RECT 68.665 73.080 68.955 73.125 ;
        RECT 67.270 72.940 68.955 73.080 ;
        RECT 67.270 72.880 67.590 72.940 ;
        RECT 68.665 72.895 68.955 72.940 ;
        RECT 70.030 72.880 70.350 73.140 ;
        RECT 70.490 72.880 70.810 73.140 ;
        RECT 70.950 72.880 71.270 73.140 ;
        RECT 73.710 73.080 74.030 73.140 ;
        RECT 73.710 72.940 74.400 73.080 ;
        RECT 73.710 72.880 74.030 72.940 ;
        RECT 40.605 72.740 40.895 72.785 ;
        RECT 39.670 72.600 40.895 72.740 ;
        RECT 39.670 72.540 39.990 72.600 ;
        RECT 40.605 72.555 40.895 72.600 ;
        RECT 41.050 72.740 41.370 72.800 ;
        RECT 42.430 72.740 42.750 72.800 ;
        RECT 44.285 72.740 44.575 72.785 ;
        RECT 41.050 72.600 44.575 72.740 ;
        RECT 41.050 72.540 41.370 72.600 ;
        RECT 42.430 72.540 42.750 72.600 ;
        RECT 44.285 72.555 44.575 72.600 ;
        RECT 53.470 72.740 53.790 72.800 ;
        RECT 66.350 72.740 66.670 72.800 ;
        RECT 70.120 72.740 70.260 72.880 ;
        RECT 53.470 72.600 63.360 72.740 ;
        RECT 17.145 72.215 17.435 72.445 ;
        RECT 17.220 71.720 17.360 72.215 ;
        RECT 21.270 72.200 21.590 72.460 ;
        RECT 22.650 72.400 22.970 72.460 ;
        RECT 21.820 72.260 22.970 72.400 ;
        RECT 18.050 71.860 18.370 72.120 ;
        RECT 21.820 72.105 21.960 72.260 ;
        RECT 22.650 72.200 22.970 72.260 ;
        RECT 28.645 72.400 28.935 72.445 ;
        RECT 39.760 72.400 39.900 72.540 ;
        RECT 28.645 72.260 39.900 72.400 ;
        RECT 44.360 72.400 44.500 72.555 ;
        RECT 53.470 72.540 53.790 72.600 ;
        RECT 48.425 72.400 48.715 72.445 ;
        RECT 44.360 72.260 48.715 72.400 ;
        RECT 28.645 72.215 28.935 72.260 ;
        RECT 48.425 72.215 48.715 72.260 ;
        RECT 49.760 72.400 50.050 72.445 ;
        RECT 49.760 72.260 56.000 72.400 ;
        RECT 49.760 72.215 50.050 72.260 ;
        RECT 21.745 71.875 22.035 72.105 ;
        RECT 22.190 71.860 22.510 72.120 ;
        RECT 24.950 71.860 25.270 72.120 ;
        RECT 25.885 72.060 26.175 72.105 ;
        RECT 37.830 72.060 38.150 72.120 ;
        RECT 25.885 71.920 38.150 72.060 ;
        RECT 25.885 71.875 26.175 71.920 ;
        RECT 37.830 71.860 38.150 71.920 ;
        RECT 49.305 72.060 49.595 72.105 ;
        RECT 50.495 72.060 50.785 72.105 ;
        RECT 53.015 72.060 53.305 72.105 ;
        RECT 49.305 71.920 53.305 72.060 ;
        RECT 49.305 71.875 49.595 71.920 ;
        RECT 50.495 71.875 50.785 71.920 ;
        RECT 53.015 71.875 53.305 71.920 ;
        RECT 53.470 72.060 53.790 72.120 ;
        RECT 53.470 71.920 55.540 72.060 ;
        RECT 53.470 71.860 53.790 71.920 ;
        RECT 20.810 71.720 21.130 71.780 ;
        RECT 55.400 71.765 55.540 71.920 ;
        RECT 55.860 71.765 56.000 72.260 ;
        RECT 57.610 72.200 57.930 72.460 ;
        RECT 63.220 72.445 63.360 72.600 ;
        RECT 66.350 72.600 70.260 72.740 ;
        RECT 66.350 72.540 66.670 72.600 ;
        RECT 58.085 72.400 58.375 72.445 ;
        RECT 59.925 72.400 60.215 72.445 ;
        RECT 58.085 72.260 60.215 72.400 ;
        RECT 58.085 72.215 58.375 72.260 ;
        RECT 59.925 72.215 60.215 72.260 ;
        RECT 63.145 72.215 63.435 72.445 ;
        RECT 64.050 72.400 64.370 72.460 ;
        RECT 65.905 72.400 66.195 72.445 ;
        RECT 64.050 72.260 66.195 72.400 ;
        RECT 64.050 72.200 64.370 72.260 ;
        RECT 65.905 72.215 66.195 72.260 ;
        RECT 68.650 72.200 68.970 72.460 ;
        RECT 69.660 72.445 69.800 72.600 ;
        RECT 69.585 72.215 69.875 72.445 ;
        RECT 70.030 72.200 70.350 72.460 ;
        RECT 71.040 72.445 71.180 72.880 ;
        RECT 72.390 72.600 73.020 72.740 ;
        RECT 72.390 72.445 72.530 72.600 ;
        RECT 70.965 72.400 71.255 72.445 ;
        RECT 70.580 72.260 71.255 72.400 ;
        RECT 58.545 71.875 58.835 72.105 ;
        RECT 48.910 71.720 49.200 71.765 ;
        RECT 51.010 71.720 51.300 71.765 ;
        RECT 52.580 71.720 52.870 71.765 ;
        RECT 17.220 71.580 21.730 71.720 ;
        RECT 20.810 71.520 21.130 71.580 ;
        RECT 15.290 71.180 15.610 71.440 ;
        RECT 18.970 71.380 19.290 71.440 ;
        RECT 19.445 71.380 19.735 71.425 ;
        RECT 18.970 71.240 19.735 71.380 ;
        RECT 21.590 71.380 21.730 71.580 ;
        RECT 48.910 71.580 52.870 71.720 ;
        RECT 48.910 71.535 49.200 71.580 ;
        RECT 51.010 71.535 51.300 71.580 ;
        RECT 52.580 71.535 52.870 71.580 ;
        RECT 55.325 71.535 55.615 71.765 ;
        RECT 55.785 71.535 56.075 71.765 ;
        RECT 56.230 71.720 56.550 71.780 ;
        RECT 58.620 71.720 58.760 71.875 ;
        RECT 70.580 71.780 70.720 72.260 ;
        RECT 70.965 72.215 71.255 72.260 ;
        RECT 71.455 72.215 71.745 72.445 ;
        RECT 72.315 72.215 72.605 72.445 ;
        RECT 56.230 71.580 58.760 71.720 ;
        RECT 56.230 71.520 56.550 71.580 ;
        RECT 70.490 71.520 70.810 71.780 ;
        RECT 71.505 71.720 71.645 72.215 ;
        RECT 72.880 72.060 73.020 72.600 ;
        RECT 73.710 72.200 74.030 72.460 ;
        RECT 74.260 72.415 74.400 72.940 ;
        RECT 76.485 72.895 76.775 73.125 ;
        RECT 76.930 73.080 77.250 73.140 ;
        RECT 80.150 73.080 80.470 73.140 ;
        RECT 76.930 72.940 80.470 73.080 ;
        RECT 74.645 72.740 74.935 72.785 ;
        RECT 76.010 72.740 76.330 72.800 ;
        RECT 74.645 72.600 76.330 72.740 ;
        RECT 76.560 72.740 76.700 72.895 ;
        RECT 76.930 72.880 77.250 72.940 ;
        RECT 80.150 72.880 80.470 72.940 ;
        RECT 82.910 72.880 83.230 73.140 ;
        RECT 85.225 72.740 85.515 72.785 ;
        RECT 76.560 72.600 85.515 72.740 ;
        RECT 74.645 72.555 74.935 72.600 ;
        RECT 76.010 72.540 76.330 72.600 ;
        RECT 85.225 72.555 85.515 72.600 ;
        RECT 74.260 72.400 74.860 72.415 ;
        RECT 75.105 72.400 75.395 72.445 ;
        RECT 74.260 72.275 75.395 72.400 ;
        RECT 74.720 72.260 75.395 72.275 ;
        RECT 75.105 72.215 75.395 72.260 ;
        RECT 75.565 72.215 75.855 72.445 ;
        RECT 76.945 72.400 77.235 72.445 ;
        RECT 77.390 72.400 77.710 72.460 ;
        RECT 76.945 72.260 77.710 72.400 ;
        RECT 76.945 72.215 77.235 72.260 ;
        RECT 74.170 72.060 74.490 72.120 ;
        RECT 72.880 71.920 74.490 72.060 ;
        RECT 75.640 72.060 75.780 72.215 ;
        RECT 77.390 72.200 77.710 72.260 ;
        RECT 77.850 72.200 78.170 72.460 ;
        RECT 78.325 72.215 78.615 72.445 ;
        RECT 78.785 72.400 79.075 72.445 ;
        RECT 79.230 72.400 79.550 72.460 ;
        RECT 78.785 72.260 79.550 72.400 ;
        RECT 78.785 72.215 79.075 72.260 ;
        RECT 76.010 72.060 76.330 72.120 ;
        RECT 75.640 71.920 76.330 72.060 ;
        RECT 78.400 72.060 78.540 72.215 ;
        RECT 79.230 72.200 79.550 72.260 ;
        RECT 84.765 72.400 85.055 72.445 ;
        RECT 87.065 72.400 87.355 72.445 ;
        RECT 84.765 72.260 87.355 72.400 ;
        RECT 84.765 72.215 85.055 72.260 ;
        RECT 87.065 72.215 87.355 72.260 ;
        RECT 88.430 72.400 88.750 72.460 ;
        RECT 89.825 72.400 90.115 72.445 ;
        RECT 88.430 72.260 90.115 72.400 ;
        RECT 88.430 72.200 88.750 72.260 ;
        RECT 89.825 72.215 90.115 72.260 ;
        RECT 79.690 72.060 80.010 72.120 ;
        RECT 78.400 71.920 80.010 72.060 ;
        RECT 74.170 71.860 74.490 71.920 ;
        RECT 76.010 71.860 76.330 71.920 ;
        RECT 79.690 71.860 80.010 71.920 ;
        RECT 85.685 71.875 85.975 72.105 ;
        RECT 80.165 71.720 80.455 71.765 ;
        RECT 85.760 71.720 85.900 71.875 ;
        RECT 71.505 71.580 73.020 71.720 ;
        RECT 66.810 71.380 67.130 71.440 ;
        RECT 21.590 71.240 67.130 71.380 ;
        RECT 18.970 71.180 19.290 71.240 ;
        RECT 19.445 71.195 19.735 71.240 ;
        RECT 66.810 71.180 67.130 71.240 ;
        RECT 72.330 71.180 72.650 71.440 ;
        RECT 72.880 71.380 73.020 71.580 ;
        RECT 80.165 71.580 85.900 71.720 ;
        RECT 80.165 71.535 80.455 71.580 ;
        RECT 75.550 71.380 75.870 71.440 ;
        RECT 72.880 71.240 75.870 71.380 ;
        RECT 75.550 71.180 75.870 71.240 ;
        RECT 13.380 70.560 92.040 71.040 ;
        RECT 19.430 70.360 19.750 70.420 ;
        RECT 20.810 70.360 21.130 70.420 ;
        RECT 21.745 70.360 22.035 70.405 ;
        RECT 19.430 70.220 22.035 70.360 ;
        RECT 19.430 70.160 19.750 70.220 ;
        RECT 20.810 70.160 21.130 70.220 ;
        RECT 21.745 70.175 22.035 70.220 ;
        RECT 73.710 70.160 74.030 70.420 ;
        RECT 75.550 70.160 75.870 70.420 ;
        RECT 76.485 70.360 76.775 70.405 ;
        RECT 77.850 70.360 78.170 70.420 ;
        RECT 76.485 70.220 78.170 70.360 ;
        RECT 76.485 70.175 76.775 70.220 ;
        RECT 77.850 70.160 78.170 70.220 ;
        RECT 15.330 70.020 15.620 70.065 ;
        RECT 17.430 70.020 17.720 70.065 ;
        RECT 19.000 70.020 19.290 70.065 ;
        RECT 15.330 69.880 19.290 70.020 ;
        RECT 15.330 69.835 15.620 69.880 ;
        RECT 17.430 69.835 17.720 69.880 ;
        RECT 19.000 69.835 19.290 69.880 ;
        RECT 21.270 70.020 21.590 70.080 ;
        RECT 24.950 70.020 25.270 70.080 ;
        RECT 21.270 69.880 25.270 70.020 ;
        RECT 21.270 69.820 21.590 69.880 ;
        RECT 24.950 69.820 25.270 69.880 ;
        RECT 27.290 70.020 27.580 70.065 ;
        RECT 29.390 70.020 29.680 70.065 ;
        RECT 30.960 70.020 31.250 70.065 ;
        RECT 27.290 69.880 31.250 70.020 ;
        RECT 27.290 69.835 27.580 69.880 ;
        RECT 29.390 69.835 29.680 69.880 ;
        RECT 30.960 69.835 31.250 69.880 ;
        RECT 41.090 70.020 41.380 70.065 ;
        RECT 43.190 70.020 43.480 70.065 ;
        RECT 44.760 70.020 45.050 70.065 ;
        RECT 41.090 69.880 45.050 70.020 ;
        RECT 41.090 69.835 41.380 69.880 ;
        RECT 43.190 69.835 43.480 69.880 ;
        RECT 44.760 69.835 45.050 69.880 ;
        RECT 47.505 70.020 47.795 70.065 ;
        RECT 72.330 70.020 72.650 70.080 ;
        RECT 74.170 70.020 74.490 70.080 ;
        RECT 75.640 70.020 75.780 70.160 ;
        RECT 47.505 69.880 55.540 70.020 ;
        RECT 47.505 69.835 47.795 69.880 ;
        RECT 55.400 69.740 55.540 69.880 ;
        RECT 72.330 69.880 75.780 70.020 ;
        RECT 76.930 70.020 77.250 70.080 ;
        RECT 79.230 70.020 79.550 70.080 ;
        RECT 76.930 69.880 79.550 70.020 ;
        RECT 72.330 69.820 72.650 69.880 ;
        RECT 74.170 69.820 74.490 69.880 ;
        RECT 76.930 69.820 77.250 69.880 ;
        RECT 79.230 69.820 79.550 69.880 ;
        RECT 15.725 69.680 16.015 69.725 ;
        RECT 16.915 69.680 17.205 69.725 ;
        RECT 19.435 69.680 19.725 69.725 ;
        RECT 15.725 69.540 19.725 69.680 ;
        RECT 15.725 69.495 16.015 69.540 ;
        RECT 16.915 69.495 17.205 69.540 ;
        RECT 19.435 69.495 19.725 69.540 ;
        RECT 26.790 69.480 27.110 69.740 ;
        RECT 27.685 69.680 27.975 69.725 ;
        RECT 28.875 69.680 29.165 69.725 ;
        RECT 31.395 69.680 31.685 69.725 ;
        RECT 27.685 69.540 31.685 69.680 ;
        RECT 27.685 69.495 27.975 69.540 ;
        RECT 28.875 69.495 29.165 69.540 ;
        RECT 31.395 69.495 31.685 69.540 ;
        RECT 39.685 69.680 39.975 69.725 ;
        RECT 41.485 69.680 41.775 69.725 ;
        RECT 42.675 69.680 42.965 69.725 ;
        RECT 45.195 69.680 45.485 69.725 ;
        RECT 39.685 69.540 40.360 69.680 ;
        RECT 39.685 69.495 39.975 69.540 ;
        RECT 14.845 69.340 15.135 69.385 ;
        RECT 21.730 69.340 22.050 69.400 ;
        RECT 14.845 69.200 22.050 69.340 ;
        RECT 14.845 69.155 15.135 69.200 ;
        RECT 21.730 69.140 22.050 69.200 ;
        RECT 15.290 69.000 15.610 69.060 ;
        RECT 16.070 69.000 16.360 69.045 ;
        RECT 15.290 68.860 16.360 69.000 ;
        RECT 15.290 68.800 15.610 68.860 ;
        RECT 16.070 68.815 16.360 68.860 ;
        RECT 28.140 69.000 28.430 69.045 ;
        RECT 29.090 69.000 29.410 69.060 ;
        RECT 28.140 68.860 29.410 69.000 ;
        RECT 40.220 69.000 40.360 69.540 ;
        RECT 41.485 69.540 45.485 69.680 ;
        RECT 41.485 69.495 41.775 69.540 ;
        RECT 42.675 69.495 42.965 69.540 ;
        RECT 45.195 69.495 45.485 69.540 ;
        RECT 51.185 69.680 51.475 69.725 ;
        RECT 52.090 69.680 52.410 69.740 ;
        RECT 51.185 69.540 52.410 69.680 ;
        RECT 51.185 69.495 51.475 69.540 ;
        RECT 52.090 69.480 52.410 69.540 ;
        RECT 55.310 69.480 55.630 69.740 ;
        RECT 64.050 69.680 64.370 69.740 ;
        RECT 64.525 69.680 64.815 69.725 ;
        RECT 64.050 69.540 64.815 69.680 ;
        RECT 64.050 69.480 64.370 69.540 ;
        RECT 64.525 69.495 64.815 69.540 ;
        RECT 68.190 69.680 68.510 69.740 ;
        RECT 69.585 69.680 69.875 69.725 ;
        RECT 68.190 69.540 74.860 69.680 ;
        RECT 68.190 69.480 68.510 69.540 ;
        RECT 69.585 69.495 69.875 69.540 ;
        RECT 40.605 69.340 40.895 69.385 ;
        RECT 41.050 69.340 41.370 69.400 ;
        RECT 48.870 69.340 49.190 69.400 ;
        RECT 40.605 69.200 41.370 69.340 ;
        RECT 40.605 69.155 40.895 69.200 ;
        RECT 41.050 69.140 41.370 69.200 ;
        RECT 41.600 69.200 49.190 69.340 ;
        RECT 41.600 69.000 41.740 69.200 ;
        RECT 48.870 69.140 49.190 69.200 ;
        RECT 58.990 69.340 59.310 69.400 ;
        RECT 60.845 69.340 61.135 69.385 ;
        RECT 65.430 69.340 65.750 69.400 ;
        RECT 58.990 69.200 65.750 69.340 ;
        RECT 58.990 69.140 59.310 69.200 ;
        RECT 60.845 69.155 61.135 69.200 ;
        RECT 65.430 69.140 65.750 69.200 ;
        RECT 65.905 69.155 66.195 69.385 ;
        RECT 40.220 68.860 41.740 69.000 ;
        RECT 41.940 69.000 42.230 69.045 ;
        RECT 57.150 69.000 57.470 69.060 ;
        RECT 65.980 69.000 66.120 69.155 ;
        RECT 70.490 69.140 70.810 69.400 ;
        RECT 70.950 69.340 71.270 69.400 ;
        RECT 72.345 69.340 72.635 69.385 ;
        RECT 70.950 69.200 72.635 69.340 ;
        RECT 70.950 69.140 71.270 69.200 ;
        RECT 72.345 69.155 72.635 69.200 ;
        RECT 72.805 69.155 73.095 69.385 ;
        RECT 41.940 68.860 48.180 69.000 ;
        RECT 28.140 68.815 28.430 68.860 ;
        RECT 29.090 68.800 29.410 68.860 ;
        RECT 41.940 68.815 42.230 68.860 ;
        RECT 33.705 68.660 33.995 68.705 ;
        RECT 34.150 68.660 34.470 68.720 ;
        RECT 33.705 68.520 34.470 68.660 ;
        RECT 33.705 68.475 33.995 68.520 ;
        RECT 34.150 68.460 34.470 68.520 ;
        RECT 36.450 68.460 36.770 68.720 ;
        RECT 38.290 68.460 38.610 68.720 ;
        RECT 38.750 68.460 39.070 68.720 ;
        RECT 48.040 68.705 48.180 68.860 ;
        RECT 57.150 68.860 66.120 69.000 ;
        RECT 66.810 69.000 67.130 69.060 ;
        RECT 71.410 69.000 71.730 69.060 ;
        RECT 72.880 69.000 73.020 69.155 ;
        RECT 73.250 69.140 73.570 69.400 ;
        RECT 74.720 69.385 74.860 69.540 ;
        RECT 75.090 69.480 75.410 69.740 ;
        RECT 80.150 69.680 80.470 69.740 ;
        RECT 80.150 69.540 81.300 69.680 ;
        RECT 80.150 69.480 80.470 69.540 ;
        RECT 74.185 69.155 74.475 69.385 ;
        RECT 74.645 69.155 74.935 69.385 ;
        RECT 66.810 68.860 70.030 69.000 ;
        RECT 57.150 68.800 57.470 68.860 ;
        RECT 66.810 68.800 67.130 68.860 ;
        RECT 47.965 68.475 48.255 68.705 ;
        RECT 49.790 68.460 50.110 68.720 ;
        RECT 50.265 68.660 50.555 68.705 ;
        RECT 52.565 68.660 52.855 68.705 ;
        RECT 50.265 68.520 52.855 68.660 ;
        RECT 50.265 68.475 50.555 68.520 ;
        RECT 52.565 68.475 52.855 68.520 ;
        RECT 67.270 68.660 67.590 68.720 ;
        RECT 69.125 68.660 69.415 68.705 ;
        RECT 67.270 68.520 69.415 68.660 ;
        RECT 69.890 68.660 70.030 68.860 ;
        RECT 71.410 68.860 73.020 69.000 ;
        RECT 73.710 69.000 74.030 69.060 ;
        RECT 74.260 69.000 74.400 69.155 ;
        RECT 75.180 69.000 75.320 69.480 ;
        RECT 79.230 69.140 79.550 69.400 ;
        RECT 81.160 69.385 81.300 69.540 ;
        RECT 81.085 69.155 81.375 69.385 ;
        RECT 86.605 69.340 86.895 69.385 ;
        RECT 87.510 69.340 87.830 69.400 ;
        RECT 86.605 69.200 87.830 69.340 ;
        RECT 86.605 69.155 86.895 69.200 ;
        RECT 87.510 69.140 87.830 69.200 ;
        RECT 89.810 69.140 90.130 69.400 ;
        RECT 73.710 68.860 75.320 69.000 ;
        RECT 78.770 69.000 79.090 69.060 ;
        RECT 79.690 69.000 80.010 69.060 ;
        RECT 80.165 69.000 80.455 69.045 ;
        RECT 78.770 68.860 80.455 69.000 ;
        RECT 71.410 68.800 71.730 68.860 ;
        RECT 73.710 68.800 74.030 68.860 ;
        RECT 78.770 68.800 79.090 68.860 ;
        RECT 79.690 68.800 80.010 68.860 ;
        RECT 80.165 68.815 80.455 68.860 ;
        RECT 80.625 69.000 80.915 69.045 ;
        RECT 82.910 69.000 83.230 69.060 ;
        RECT 80.625 68.860 83.230 69.000 ;
        RECT 80.625 68.815 80.915 68.860 ;
        RECT 80.700 68.660 80.840 68.815 ;
        RECT 82.910 68.800 83.230 68.860 ;
        RECT 69.890 68.520 80.840 68.660 ;
        RECT 82.005 68.660 82.295 68.705 ;
        RECT 84.750 68.660 85.070 68.720 ;
        RECT 82.005 68.520 85.070 68.660 ;
        RECT 67.270 68.460 67.590 68.520 ;
        RECT 69.125 68.475 69.415 68.520 ;
        RECT 82.005 68.475 82.295 68.520 ;
        RECT 84.750 68.460 85.070 68.520 ;
        RECT 85.670 68.460 85.990 68.720 ;
        RECT 87.050 68.460 87.370 68.720 ;
        RECT 13.380 67.840 92.040 68.320 ;
        RECT 14.370 67.640 14.690 67.700 ;
        RECT 15.305 67.640 15.595 67.685 ;
        RECT 14.370 67.500 15.595 67.640 ;
        RECT 14.370 67.440 14.690 67.500 ;
        RECT 15.305 67.455 15.595 67.500 ;
        RECT 16.300 67.500 23.800 67.640 ;
        RECT 16.300 67.005 16.440 67.500 ;
        RECT 21.730 67.300 22.050 67.360 ;
        RECT 17.680 67.160 22.050 67.300 ;
        RECT 17.680 67.005 17.820 67.160 ;
        RECT 21.730 67.100 22.050 67.160 ;
        RECT 18.970 67.005 19.290 67.020 ;
        RECT 16.225 66.775 16.515 67.005 ;
        RECT 17.605 66.775 17.895 67.005 ;
        RECT 18.940 66.960 19.290 67.005 ;
        RECT 18.775 66.820 19.290 66.960 ;
        RECT 23.660 66.960 23.800 67.500 ;
        RECT 24.505 67.455 24.795 67.685 ;
        RECT 27.265 67.640 27.555 67.685 ;
        RECT 27.710 67.640 28.030 67.700 ;
        RECT 27.265 67.500 28.030 67.640 ;
        RECT 27.265 67.455 27.555 67.500 ;
        RECT 24.580 67.300 24.720 67.455 ;
        RECT 27.710 67.440 28.030 67.500 ;
        RECT 29.090 67.440 29.410 67.700 ;
        RECT 38.290 67.640 38.610 67.700 ;
        RECT 40.145 67.640 40.435 67.685 ;
        RECT 38.290 67.500 40.435 67.640 ;
        RECT 38.290 67.440 38.610 67.500 ;
        RECT 40.145 67.455 40.435 67.500 ;
        RECT 43.350 67.640 43.670 67.700 ;
        RECT 48.410 67.640 48.730 67.700 ;
        RECT 43.350 67.500 48.730 67.640 ;
        RECT 43.350 67.440 43.670 67.500 ;
        RECT 48.410 67.440 48.730 67.500 ;
        RECT 53.025 67.640 53.315 67.685 ;
        RECT 54.390 67.640 54.710 67.700 ;
        RECT 53.025 67.500 54.710 67.640 ;
        RECT 53.025 67.455 53.315 67.500 ;
        RECT 54.390 67.440 54.710 67.500 ;
        RECT 55.325 67.640 55.615 67.685 ;
        RECT 57.150 67.640 57.470 67.700 ;
        RECT 55.325 67.500 57.470 67.640 ;
        RECT 55.325 67.455 55.615 67.500 ;
        RECT 57.150 67.440 57.470 67.500 ;
        RECT 65.445 67.455 65.735 67.685 ;
        RECT 24.950 67.300 25.270 67.360 ;
        RECT 62.840 67.300 63.130 67.345 ;
        RECT 65.520 67.300 65.660 67.455 ;
        RECT 67.270 67.440 67.590 67.700 ;
        RECT 74.645 67.455 74.935 67.685 ;
        RECT 78.325 67.640 78.615 67.685 ;
        RECT 86.590 67.640 86.910 67.700 ;
        RECT 78.325 67.500 86.910 67.640 ;
        RECT 78.325 67.455 78.615 67.500 ;
        RECT 24.580 67.160 59.680 67.300 ;
        RECT 24.950 67.100 25.270 67.160 ;
        RECT 23.660 66.820 31.160 66.960 ;
        RECT 18.940 66.775 19.290 66.820 ;
        RECT 18.970 66.760 19.290 66.775 ;
        RECT 18.485 66.620 18.775 66.665 ;
        RECT 19.675 66.620 19.965 66.665 ;
        RECT 22.195 66.620 22.485 66.665 ;
        RECT 18.485 66.480 22.485 66.620 ;
        RECT 18.485 66.435 18.775 66.480 ;
        RECT 19.675 66.435 19.965 66.480 ;
        RECT 22.195 66.435 22.485 66.480 ;
        RECT 25.870 66.420 26.190 66.680 ;
        RECT 26.805 66.620 27.095 66.665 ;
        RECT 28.170 66.620 28.490 66.680 ;
        RECT 26.805 66.480 28.490 66.620 ;
        RECT 31.020 66.620 31.160 66.820 ;
        RECT 43.350 66.760 43.670 67.020 ;
        RECT 43.810 66.760 44.130 67.020 ;
        RECT 44.285 66.960 44.575 67.005 ;
        RECT 44.730 66.960 45.050 67.020 ;
        RECT 44.285 66.820 45.050 66.960 ;
        RECT 44.285 66.775 44.575 66.820 ;
        RECT 44.730 66.760 45.050 66.820 ;
        RECT 45.205 66.775 45.495 67.005 ;
        RECT 45.665 66.960 45.955 67.005 ;
        RECT 49.330 66.960 49.650 67.020 ;
        RECT 45.665 66.820 49.650 66.960 ;
        RECT 45.665 66.775 45.955 66.820 ;
        RECT 31.390 66.620 31.710 66.680 ;
        RECT 45.280 66.620 45.420 66.775 ;
        RECT 49.330 66.760 49.650 66.820 ;
        RECT 54.865 66.960 55.155 67.005 ;
        RECT 58.990 66.960 59.310 67.020 ;
        RECT 54.865 66.820 59.310 66.960 ;
        RECT 59.540 66.960 59.680 67.160 ;
        RECT 62.840 67.160 65.660 67.300 ;
        RECT 65.980 67.160 74.400 67.300 ;
        RECT 62.840 67.115 63.130 67.160 ;
        RECT 65.980 66.960 66.120 67.160 ;
        RECT 59.540 66.820 66.120 66.960 ;
        RECT 67.745 66.960 68.035 67.005 ;
        RECT 68.650 66.960 68.970 67.020 ;
        RECT 70.950 66.960 71.270 67.020 ;
        RECT 67.745 66.820 71.270 66.960 ;
        RECT 54.865 66.775 55.155 66.820 ;
        RECT 58.990 66.760 59.310 66.820 ;
        RECT 67.745 66.775 68.035 66.820 ;
        RECT 68.650 66.760 68.970 66.820 ;
        RECT 70.950 66.760 71.270 66.820 ;
        RECT 72.330 66.960 72.650 67.020 ;
        RECT 72.805 66.960 73.095 67.005 ;
        RECT 72.330 66.820 73.095 66.960 ;
        RECT 72.330 66.760 72.650 66.820 ;
        RECT 72.805 66.775 73.095 66.820 ;
        RECT 73.710 66.760 74.030 67.020 ;
        RECT 31.020 66.480 45.420 66.620 ;
        RECT 26.805 66.435 27.095 66.480 ;
        RECT 28.170 66.420 28.490 66.480 ;
        RECT 31.390 66.420 31.710 66.480 ;
        RECT 48.410 66.420 48.730 66.680 ;
        RECT 51.170 66.420 51.490 66.680 ;
        RECT 55.785 66.435 56.075 66.665 ;
        RECT 59.475 66.620 59.765 66.665 ;
        RECT 61.995 66.620 62.285 66.665 ;
        RECT 63.185 66.620 63.475 66.665 ;
        RECT 59.475 66.480 63.475 66.620 ;
        RECT 59.475 66.435 59.765 66.480 ;
        RECT 61.995 66.435 62.285 66.480 ;
        RECT 63.185 66.435 63.475 66.480 ;
        RECT 64.065 66.620 64.355 66.665 ;
        RECT 64.510 66.620 64.830 66.680 ;
        RECT 64.065 66.480 64.830 66.620 ;
        RECT 64.065 66.435 64.355 66.480 ;
        RECT 18.090 66.280 18.380 66.325 ;
        RECT 20.190 66.280 20.480 66.325 ;
        RECT 21.760 66.280 22.050 66.325 ;
        RECT 18.090 66.140 22.050 66.280 ;
        RECT 18.090 66.095 18.380 66.140 ;
        RECT 20.190 66.095 20.480 66.140 ;
        RECT 21.760 66.095 22.050 66.140 ;
        RECT 46.585 66.280 46.875 66.325 ;
        RECT 53.010 66.280 53.330 66.340 ;
        RECT 46.585 66.140 53.330 66.280 ;
        RECT 46.585 66.095 46.875 66.140 ;
        RECT 53.010 66.080 53.330 66.140 ;
        RECT 19.430 65.940 19.750 66.000 ;
        RECT 21.270 65.940 21.590 66.000 ;
        RECT 19.430 65.800 21.590 65.940 ;
        RECT 19.430 65.740 19.750 65.800 ;
        RECT 21.270 65.740 21.590 65.800 ;
        RECT 47.490 65.940 47.810 66.000 ;
        RECT 55.860 65.940 56.000 66.435 ;
        RECT 64.510 66.420 64.830 66.480 ;
        RECT 68.205 66.620 68.495 66.665 ;
        RECT 69.570 66.620 69.890 66.680 ;
        RECT 68.205 66.480 69.890 66.620 ;
        RECT 74.260 66.620 74.400 67.160 ;
        RECT 74.720 66.960 74.860 67.455 ;
        RECT 86.590 67.440 86.910 67.500 ;
        RECT 88.430 67.640 88.750 67.700 ;
        RECT 88.905 67.640 89.195 67.685 ;
        RECT 89.810 67.640 90.130 67.700 ;
        RECT 88.430 67.500 90.130 67.640 ;
        RECT 88.430 67.440 88.750 67.500 ;
        RECT 88.905 67.455 89.195 67.500 ;
        RECT 89.810 67.440 90.130 67.500 ;
        RECT 77.390 67.300 77.710 67.360 ;
        RECT 76.100 67.160 77.710 67.300 ;
        RECT 76.100 67.005 76.240 67.160 ;
        RECT 77.390 67.100 77.710 67.160 ;
        RECT 79.690 67.100 80.010 67.360 ;
        RECT 83.340 67.300 83.630 67.345 ;
        RECT 83.830 67.300 84.150 67.360 ;
        RECT 83.340 67.160 84.150 67.300 ;
        RECT 83.340 67.115 83.630 67.160 ;
        RECT 83.830 67.100 84.150 67.160 ;
        RECT 75.105 66.960 75.395 67.005 ;
        RECT 74.720 66.820 75.395 66.960 ;
        RECT 75.105 66.775 75.395 66.820 ;
        RECT 76.025 66.775 76.315 67.005 ;
        RECT 76.470 66.760 76.790 67.020 ;
        RECT 76.930 66.760 77.250 67.020 ;
        RECT 78.770 66.760 79.090 67.020 ;
        RECT 80.165 66.775 80.455 67.005 ;
        RECT 80.240 66.620 80.380 66.775 ;
        RECT 80.610 66.760 80.930 67.020 ;
        RECT 81.530 66.960 81.850 67.020 ;
        RECT 82.005 66.960 82.295 67.005 ;
        RECT 81.530 66.820 82.295 66.960 ;
        RECT 81.530 66.760 81.850 66.820 ;
        RECT 82.005 66.775 82.295 66.820 ;
        RECT 82.450 66.760 82.770 67.020 ;
        RECT 90.270 66.760 90.590 67.020 ;
        RECT 82.540 66.620 82.680 66.760 ;
        RECT 74.260 66.480 82.680 66.620 ;
        RECT 82.885 66.620 83.175 66.665 ;
        RECT 84.075 66.620 84.365 66.665 ;
        RECT 86.595 66.620 86.885 66.665 ;
        RECT 82.885 66.480 86.885 66.620 ;
        RECT 68.205 66.435 68.495 66.480 ;
        RECT 69.570 66.420 69.890 66.480 ;
        RECT 82.885 66.435 83.175 66.480 ;
        RECT 84.075 66.435 84.365 66.480 ;
        RECT 86.595 66.435 86.885 66.480 ;
        RECT 59.910 66.280 60.200 66.325 ;
        RECT 61.480 66.280 61.770 66.325 ;
        RECT 63.580 66.280 63.870 66.325 ;
        RECT 59.910 66.140 63.870 66.280 ;
        RECT 59.910 66.095 60.200 66.140 ;
        RECT 61.480 66.095 61.770 66.140 ;
        RECT 63.580 66.095 63.870 66.140 ;
        RECT 71.870 66.280 72.190 66.340 ;
        RECT 76.470 66.280 76.790 66.340 ;
        RECT 71.870 66.140 76.790 66.280 ;
        RECT 71.870 66.080 72.190 66.140 ;
        RECT 76.470 66.080 76.790 66.140 ;
        RECT 77.390 66.280 77.710 66.340 ;
        RECT 80.610 66.280 80.930 66.340 ;
        RECT 77.390 66.140 80.930 66.280 ;
        RECT 77.390 66.080 77.710 66.140 ;
        RECT 80.610 66.080 80.930 66.140 ;
        RECT 82.490 66.280 82.780 66.325 ;
        RECT 84.590 66.280 84.880 66.325 ;
        RECT 86.160 66.280 86.450 66.325 ;
        RECT 82.490 66.140 86.450 66.280 ;
        RECT 82.490 66.095 82.780 66.140 ;
        RECT 84.590 66.095 84.880 66.140 ;
        RECT 86.160 66.095 86.450 66.140 ;
        RECT 87.970 66.280 88.290 66.340 ;
        RECT 89.365 66.280 89.655 66.325 ;
        RECT 87.970 66.140 89.655 66.280 ;
        RECT 87.970 66.080 88.290 66.140 ;
        RECT 89.365 66.095 89.655 66.140 ;
        RECT 58.530 65.940 58.850 66.000 ;
        RECT 60.370 65.940 60.690 66.000 ;
        RECT 47.490 65.800 60.690 65.940 ;
        RECT 47.490 65.740 47.810 65.800 ;
        RECT 58.530 65.740 58.850 65.800 ;
        RECT 60.370 65.740 60.690 65.800 ;
        RECT 72.790 65.740 73.110 66.000 ;
        RECT 81.545 65.940 81.835 65.985 ;
        RECT 85.670 65.940 85.990 66.000 ;
        RECT 81.545 65.800 85.990 65.940 ;
        RECT 81.545 65.755 81.835 65.800 ;
        RECT 85.670 65.740 85.990 65.800 ;
        RECT 13.380 65.120 92.040 65.600 ;
        RECT 28.170 64.920 28.490 64.980 ;
        RECT 34.150 64.920 34.470 64.980 ;
        RECT 40.590 64.920 40.910 64.980 ;
        RECT 28.170 64.780 40.910 64.920 ;
        RECT 28.170 64.720 28.490 64.780 ;
        RECT 34.150 64.720 34.470 64.780 ;
        RECT 40.590 64.720 40.910 64.780 ;
        RECT 41.525 64.920 41.815 64.965 ;
        RECT 43.350 64.920 43.670 64.980 ;
        RECT 41.525 64.780 43.670 64.920 ;
        RECT 41.525 64.735 41.815 64.780 ;
        RECT 43.350 64.720 43.670 64.780 ;
        RECT 49.330 64.920 49.650 64.980 ;
        RECT 50.250 64.920 50.570 64.980 ;
        RECT 49.330 64.780 50.570 64.920 ;
        RECT 49.330 64.720 49.650 64.780 ;
        RECT 50.250 64.720 50.570 64.780 ;
        RECT 59.450 64.720 59.770 64.980 ;
        RECT 77.405 64.920 77.695 64.965 ;
        RECT 78.770 64.920 79.090 64.980 ;
        RECT 77.405 64.780 79.090 64.920 ;
        RECT 77.405 64.735 77.695 64.780 ;
        RECT 78.770 64.720 79.090 64.780 ;
        RECT 83.830 64.720 84.150 64.980 ;
        RECT 34.610 64.580 34.930 64.640 ;
        RECT 18.140 64.440 34.930 64.580 ;
        RECT 16.210 63.700 16.530 63.960 ;
        RECT 18.140 63.945 18.280 64.440 ;
        RECT 34.610 64.380 34.930 64.440 ;
        RECT 35.110 64.580 35.400 64.625 ;
        RECT 37.210 64.580 37.500 64.625 ;
        RECT 38.780 64.580 39.070 64.625 ;
        RECT 35.110 64.440 39.070 64.580 ;
        RECT 35.110 64.395 35.400 64.440 ;
        RECT 37.210 64.395 37.500 64.440 ;
        RECT 38.780 64.395 39.070 64.440 ;
        RECT 53.050 64.580 53.340 64.625 ;
        RECT 55.150 64.580 55.440 64.625 ;
        RECT 56.720 64.580 57.010 64.625 ;
        RECT 53.050 64.440 57.010 64.580 ;
        RECT 53.050 64.395 53.340 64.440 ;
        RECT 55.150 64.395 55.440 64.440 ;
        RECT 56.720 64.395 57.010 64.440 ;
        RECT 27.250 64.240 27.570 64.300 ;
        RECT 35.505 64.240 35.795 64.285 ;
        RECT 36.695 64.240 36.985 64.285 ;
        RECT 39.215 64.240 39.505 64.285 ;
        RECT 27.250 64.100 28.400 64.240 ;
        RECT 27.250 64.040 27.570 64.100 ;
        RECT 18.065 63.715 18.355 63.945 ;
        RECT 21.285 63.900 21.575 63.945 ;
        RECT 22.650 63.900 22.970 63.960 ;
        RECT 28.260 63.945 28.400 64.100 ;
        RECT 35.505 64.100 39.505 64.240 ;
        RECT 35.505 64.055 35.795 64.100 ;
        RECT 36.695 64.055 36.985 64.100 ;
        RECT 39.215 64.055 39.505 64.100 ;
        RECT 47.965 64.240 48.255 64.285 ;
        RECT 48.870 64.240 49.190 64.300 ;
        RECT 47.965 64.100 49.190 64.240 ;
        RECT 47.965 64.055 48.255 64.100 ;
        RECT 48.870 64.040 49.190 64.100 ;
        RECT 52.550 64.040 52.870 64.300 ;
        RECT 53.445 64.240 53.735 64.285 ;
        RECT 54.635 64.240 54.925 64.285 ;
        RECT 57.155 64.240 57.445 64.285 ;
        RECT 53.445 64.100 57.445 64.240 ;
        RECT 59.540 64.240 59.680 64.720 ;
        RECT 89.810 64.380 90.130 64.640 ;
        RECT 62.685 64.240 62.975 64.285 ;
        RECT 59.540 64.100 62.975 64.240 ;
        RECT 53.445 64.055 53.735 64.100 ;
        RECT 54.635 64.055 54.925 64.100 ;
        RECT 57.155 64.055 57.445 64.100 ;
        RECT 62.685 64.055 62.975 64.100 ;
        RECT 67.285 64.240 67.575 64.285 ;
        RECT 67.730 64.240 68.050 64.300 ;
        RECT 70.490 64.240 70.810 64.300 ;
        RECT 73.710 64.240 74.030 64.300 ;
        RECT 67.285 64.100 68.050 64.240 ;
        RECT 67.285 64.055 67.575 64.100 ;
        RECT 67.730 64.040 68.050 64.100 ;
        RECT 68.740 64.100 74.030 64.240 ;
        RECT 21.285 63.760 22.970 63.900 ;
        RECT 21.285 63.715 21.575 63.760 ;
        RECT 22.650 63.700 22.970 63.760 ;
        RECT 28.185 63.715 28.475 63.945 ;
        RECT 28.645 63.715 28.935 63.945 ;
        RECT 29.105 63.715 29.395 63.945 ;
        RECT 27.250 63.560 27.570 63.620 ;
        RECT 28.720 63.560 28.860 63.715 ;
        RECT 27.250 63.420 28.860 63.560 ;
        RECT 27.250 63.360 27.570 63.420 ;
        RECT 12.070 63.220 12.390 63.280 ;
        RECT 15.305 63.220 15.595 63.265 ;
        RECT 12.070 63.080 15.595 63.220 ;
        RECT 12.070 63.020 12.390 63.080 ;
        RECT 15.305 63.035 15.595 63.080 ;
        RECT 17.130 63.020 17.450 63.280 ;
        RECT 20.365 63.220 20.655 63.265 ;
        RECT 23.110 63.220 23.430 63.280 ;
        RECT 20.365 63.080 23.430 63.220 ;
        RECT 20.365 63.035 20.655 63.080 ;
        RECT 23.110 63.020 23.430 63.080 ;
        RECT 25.870 63.220 26.190 63.280 ;
        RECT 26.805 63.220 27.095 63.265 ;
        RECT 25.870 63.080 27.095 63.220 ;
        RECT 25.870 63.020 26.190 63.080 ;
        RECT 26.805 63.035 27.095 63.080 ;
        RECT 28.170 63.220 28.490 63.280 ;
        RECT 29.180 63.220 29.320 63.715 ;
        RECT 30.010 63.700 30.330 63.960 ;
        RECT 31.390 63.700 31.710 63.960 ;
        RECT 34.625 63.900 34.915 63.945 ;
        RECT 41.050 63.900 41.370 63.960 ;
        RECT 34.625 63.760 41.370 63.900 ;
        RECT 34.625 63.715 34.915 63.760 ;
        RECT 41.050 63.700 41.370 63.760 ;
        RECT 46.585 63.900 46.875 63.945 ;
        RECT 48.410 63.900 48.730 63.960 ;
        RECT 46.585 63.760 48.730 63.900 ;
        RECT 46.585 63.715 46.875 63.760 ;
        RECT 48.410 63.700 48.730 63.760 ;
        RECT 51.185 63.900 51.475 63.945 ;
        RECT 51.630 63.900 51.950 63.960 ;
        RECT 51.185 63.760 51.950 63.900 ;
        RECT 51.185 63.715 51.475 63.760 ;
        RECT 51.630 63.700 51.950 63.760 ;
        RECT 58.070 63.900 58.390 63.960 ;
        RECT 63.605 63.900 63.895 63.945 ;
        RECT 58.070 63.760 63.895 63.900 ;
        RECT 58.070 63.700 58.390 63.760 ;
        RECT 63.605 63.715 63.895 63.760 ;
        RECT 65.890 63.900 66.210 63.960 ;
        RECT 68.190 63.900 68.510 63.960 ;
        RECT 68.740 63.945 68.880 64.100 ;
        RECT 70.490 64.040 70.810 64.100 ;
        RECT 73.710 64.040 74.030 64.100 ;
        RECT 74.185 64.240 74.475 64.285 ;
        RECT 76.930 64.240 77.250 64.300 ;
        RECT 81.530 64.240 81.850 64.300 ;
        RECT 74.185 64.100 81.850 64.240 ;
        RECT 74.185 64.055 74.475 64.100 ;
        RECT 76.930 64.040 77.250 64.100 ;
        RECT 81.530 64.040 81.850 64.100 ;
        RECT 85.670 64.240 85.990 64.300 ;
        RECT 86.145 64.240 86.435 64.285 ;
        RECT 85.670 64.100 86.435 64.240 ;
        RECT 85.670 64.040 85.990 64.100 ;
        RECT 86.145 64.055 86.435 64.100 ;
        RECT 86.590 64.040 86.910 64.300 ;
        RECT 65.890 63.760 68.510 63.900 ;
        RECT 65.890 63.700 66.210 63.760 ;
        RECT 68.190 63.700 68.510 63.760 ;
        RECT 68.665 63.715 68.955 63.945 ;
        RECT 72.790 63.900 73.110 63.960 ;
        RECT 75.565 63.900 75.855 63.945 ;
        RECT 72.790 63.760 75.855 63.900 ;
        RECT 72.790 63.700 73.110 63.760 ;
        RECT 75.565 63.715 75.855 63.760 ;
        RECT 76.485 63.900 76.775 63.945 ;
        RECT 77.850 63.900 78.170 63.960 ;
        RECT 79.690 63.900 80.010 63.960 ;
        RECT 76.485 63.760 80.010 63.900 ;
        RECT 76.485 63.715 76.775 63.760 ;
        RECT 77.850 63.700 78.170 63.760 ;
        RECT 79.690 63.700 80.010 63.760 ;
        RECT 80.625 63.900 80.915 63.945 ;
        RECT 87.970 63.900 88.290 63.960 ;
        RECT 80.625 63.760 88.290 63.900 ;
        RECT 80.625 63.715 80.915 63.760 ;
        RECT 87.970 63.700 88.290 63.760 ;
        RECT 88.905 63.900 89.195 63.945 ;
        RECT 89.350 63.900 89.670 63.960 ;
        RECT 88.905 63.760 89.670 63.900 ;
        RECT 88.905 63.715 89.195 63.760 ;
        RECT 89.350 63.700 89.670 63.760 ;
        RECT 30.485 63.375 30.775 63.605 ;
        RECT 35.960 63.560 36.250 63.605 ;
        RECT 36.450 63.560 36.770 63.620 ;
        RECT 35.960 63.420 36.770 63.560 ;
        RECT 35.960 63.375 36.250 63.420 ;
        RECT 28.170 63.080 29.320 63.220 ;
        RECT 29.550 63.220 29.870 63.280 ;
        RECT 30.560 63.220 30.700 63.375 ;
        RECT 36.450 63.360 36.770 63.420 ;
        RECT 53.900 63.560 54.190 63.605 ;
        RECT 55.310 63.560 55.630 63.620 ;
        RECT 53.900 63.420 55.630 63.560 ;
        RECT 53.900 63.375 54.190 63.420 ;
        RECT 55.310 63.360 55.630 63.420 ;
        RECT 65.430 63.560 65.750 63.620 ;
        RECT 67.730 63.560 68.050 63.620 ;
        RECT 70.045 63.560 70.335 63.605 ;
        RECT 65.430 63.420 70.335 63.560 ;
        RECT 65.430 63.360 65.750 63.420 ;
        RECT 67.730 63.360 68.050 63.420 ;
        RECT 70.045 63.375 70.335 63.420 ;
        RECT 85.685 63.560 85.975 63.605 ;
        RECT 87.050 63.560 87.370 63.620 ;
        RECT 85.685 63.420 87.370 63.560 ;
        RECT 85.685 63.375 85.975 63.420 ;
        RECT 87.050 63.360 87.370 63.420 ;
        RECT 29.550 63.080 30.700 63.220 ;
        RECT 31.850 63.220 32.170 63.280 ;
        RECT 32.325 63.220 32.615 63.265 ;
        RECT 31.850 63.080 32.615 63.220 ;
        RECT 28.170 63.020 28.490 63.080 ;
        RECT 29.550 63.020 29.870 63.080 ;
        RECT 31.850 63.020 32.170 63.080 ;
        RECT 32.325 63.035 32.615 63.080 ;
        RECT 44.730 63.020 45.050 63.280 ;
        RECT 47.030 63.020 47.350 63.280 ;
        RECT 49.330 63.220 49.650 63.280 ;
        RECT 50.725 63.220 51.015 63.265 ;
        RECT 52.550 63.220 52.870 63.280 ;
        RECT 49.330 63.080 52.870 63.220 ;
        RECT 49.330 63.020 49.650 63.080 ;
        RECT 50.725 63.035 51.015 63.080 ;
        RECT 52.550 63.020 52.870 63.080 ;
        RECT 59.910 63.020 60.230 63.280 ;
        RECT 66.810 63.020 67.130 63.280 ;
        RECT 67.270 63.020 67.590 63.280 ;
        RECT 83.385 63.220 83.675 63.265 ;
        RECT 85.210 63.220 85.530 63.280 ;
        RECT 83.385 63.080 85.530 63.220 ;
        RECT 83.385 63.035 83.675 63.080 ;
        RECT 85.210 63.020 85.530 63.080 ;
        RECT 13.380 62.400 92.040 62.880 ;
        RECT 26.790 62.200 27.110 62.260 ;
        RECT 29.550 62.200 29.870 62.260 ;
        RECT 16.300 62.060 29.870 62.200 ;
        RECT 16.300 61.905 16.440 62.060 ;
        RECT 26.790 62.000 27.110 62.060 ;
        RECT 29.550 62.000 29.870 62.060 ;
        RECT 31.390 62.200 31.710 62.260 ;
        RECT 38.765 62.200 39.055 62.245 ;
        RECT 31.390 62.060 39.055 62.200 ;
        RECT 31.390 62.000 31.710 62.060 ;
        RECT 38.765 62.015 39.055 62.060 ;
        RECT 49.345 62.200 49.635 62.245 ;
        RECT 51.170 62.200 51.490 62.260 ;
        RECT 49.345 62.060 51.490 62.200 ;
        RECT 49.345 62.015 49.635 62.060 ;
        RECT 51.170 62.000 51.490 62.060 ;
        RECT 53.010 62.000 53.330 62.260 ;
        RECT 55.310 62.000 55.630 62.260 ;
        RECT 57.625 62.200 57.915 62.245 ;
        RECT 58.070 62.200 58.390 62.260 ;
        RECT 57.625 62.060 58.390 62.200 ;
        RECT 57.625 62.015 57.915 62.060 ;
        RECT 58.070 62.000 58.390 62.060 ;
        RECT 65.445 62.015 65.735 62.245 ;
        RECT 66.810 62.200 67.130 62.260 ;
        RECT 66.810 62.060 68.420 62.200 ;
        RECT 16.225 61.675 16.515 61.905 ;
        RECT 17.145 61.860 17.435 61.905 ;
        RECT 22.190 61.860 22.510 61.920 ;
        RECT 32.310 61.860 32.630 61.920 ;
        RECT 35.530 61.860 35.850 61.920 ;
        RECT 17.145 61.720 22.510 61.860 ;
        RECT 17.145 61.675 17.435 61.720 ;
        RECT 22.190 61.660 22.510 61.720 ;
        RECT 24.580 61.720 32.080 61.860 ;
        RECT 21.730 61.520 22.050 61.580 ;
        RECT 24.580 61.565 24.720 61.720 ;
        RECT 25.870 61.565 26.190 61.580 ;
        RECT 31.940 61.565 32.080 61.720 ;
        RECT 32.310 61.720 35.850 61.860 ;
        RECT 32.310 61.660 32.630 61.720 ;
        RECT 35.530 61.660 35.850 61.720 ;
        RECT 43.780 61.860 44.070 61.905 ;
        RECT 44.730 61.860 45.050 61.920 ;
        RECT 43.780 61.720 45.050 61.860 ;
        RECT 43.780 61.675 44.070 61.720 ;
        RECT 44.730 61.660 45.050 61.720 ;
        RECT 53.485 61.860 53.775 61.905 ;
        RECT 59.910 61.860 60.230 61.920 ;
        RECT 53.485 61.720 60.230 61.860 ;
        RECT 53.485 61.675 53.775 61.720 ;
        RECT 59.910 61.660 60.230 61.720 ;
        RECT 63.300 61.860 63.590 61.905 ;
        RECT 65.520 61.860 65.660 62.015 ;
        RECT 66.810 62.000 67.130 62.060 ;
        RECT 63.300 61.720 65.660 61.860 ;
        RECT 63.300 61.675 63.590 61.720 ;
        RECT 67.270 61.660 67.590 61.920 ;
        RECT 33.230 61.565 33.550 61.580 ;
        RECT 24.505 61.520 24.795 61.565 ;
        RECT 25.840 61.520 26.190 61.565 ;
        RECT 21.730 61.380 24.795 61.520 ;
        RECT 25.675 61.380 26.190 61.520 ;
        RECT 21.730 61.320 22.050 61.380 ;
        RECT 24.505 61.335 24.795 61.380 ;
        RECT 25.840 61.335 26.190 61.380 ;
        RECT 31.865 61.335 32.155 61.565 ;
        RECT 33.200 61.335 33.550 61.565 ;
        RECT 25.870 61.320 26.190 61.335 ;
        RECT 33.230 61.320 33.550 61.335 ;
        RECT 41.050 61.520 41.370 61.580 ;
        RECT 42.445 61.520 42.735 61.565 ;
        RECT 41.050 61.380 42.735 61.520 ;
        RECT 41.050 61.320 41.370 61.380 ;
        RECT 42.445 61.335 42.735 61.380 ;
        RECT 64.510 61.320 64.830 61.580 ;
        RECT 65.890 61.520 66.210 61.580 ;
        RECT 66.365 61.520 66.655 61.565 ;
        RECT 65.890 61.380 66.655 61.520 ;
        RECT 65.890 61.320 66.210 61.380 ;
        RECT 66.365 61.335 66.655 61.380 ;
        RECT 66.810 61.320 67.130 61.580 ;
        RECT 68.280 61.565 68.420 62.060 ;
        RECT 70.950 62.000 71.270 62.260 ;
        RECT 79.230 62.200 79.550 62.260 ;
        RECT 81.545 62.200 81.835 62.245 ;
        RECT 79.230 62.060 81.835 62.200 ;
        RECT 79.230 62.000 79.550 62.060 ;
        RECT 81.545 62.015 81.835 62.060 ;
        RECT 85.210 62.000 85.530 62.260 ;
        RECT 87.510 62.000 87.830 62.260 ;
        RECT 71.040 61.860 71.180 62.000 ;
        RECT 74.630 61.860 74.950 61.920 ;
        RECT 69.660 61.720 74.950 61.860 ;
        RECT 68.205 61.335 68.495 61.565 ;
        RECT 68.650 61.320 68.970 61.580 ;
        RECT 69.660 61.565 69.800 61.720 ;
        RECT 74.630 61.660 74.950 61.720 ;
        RECT 69.585 61.335 69.875 61.565 ;
        RECT 70.965 61.520 71.255 61.565 ;
        RECT 76.930 61.520 77.250 61.580 ;
        RECT 70.965 61.380 77.250 61.520 ;
        RECT 70.965 61.335 71.255 61.380 ;
        RECT 22.650 60.980 22.970 61.240 ;
        RECT 24.030 60.980 24.350 61.240 ;
        RECT 25.385 61.180 25.675 61.225 ;
        RECT 26.575 61.180 26.865 61.225 ;
        RECT 29.095 61.180 29.385 61.225 ;
        RECT 25.385 61.040 29.385 61.180 ;
        RECT 25.385 60.995 25.675 61.040 ;
        RECT 26.575 60.995 26.865 61.040 ;
        RECT 29.095 60.995 29.385 61.040 ;
        RECT 32.745 61.180 33.035 61.225 ;
        RECT 33.935 61.180 34.225 61.225 ;
        RECT 36.455 61.180 36.745 61.225 ;
        RECT 32.745 61.040 36.745 61.180 ;
        RECT 32.745 60.995 33.035 61.040 ;
        RECT 33.935 60.995 34.225 61.040 ;
        RECT 36.455 60.995 36.745 61.040 ;
        RECT 43.325 61.180 43.615 61.225 ;
        RECT 44.515 61.180 44.805 61.225 ;
        RECT 47.035 61.180 47.325 61.225 ;
        RECT 43.325 61.040 47.325 61.180 ;
        RECT 43.325 60.995 43.615 61.040 ;
        RECT 44.515 60.995 44.805 61.040 ;
        RECT 47.035 60.995 47.325 61.040 ;
        RECT 52.550 61.180 52.870 61.240 ;
        RECT 55.770 61.180 56.090 61.240 ;
        RECT 52.550 61.040 56.090 61.180 ;
        RECT 52.550 60.980 52.870 61.040 ;
        RECT 55.770 60.980 56.090 61.040 ;
        RECT 59.935 61.180 60.225 61.225 ;
        RECT 62.455 61.180 62.745 61.225 ;
        RECT 63.645 61.180 63.935 61.225 ;
        RECT 59.935 61.040 63.935 61.180 ;
        RECT 64.600 61.180 64.740 61.320 ;
        RECT 71.040 61.180 71.180 61.335 ;
        RECT 76.930 61.320 77.250 61.380 ;
        RECT 77.850 61.520 78.170 61.580 ;
        RECT 81.070 61.520 81.390 61.580 ;
        RECT 77.850 61.380 81.390 61.520 ;
        RECT 77.850 61.320 78.170 61.380 ;
        RECT 81.070 61.320 81.390 61.380 ;
        RECT 82.005 61.335 82.295 61.565 ;
        RECT 64.600 61.040 71.180 61.180 ;
        RECT 73.710 61.180 74.030 61.240 ;
        RECT 82.080 61.180 82.220 61.335 ;
        RECT 88.430 61.320 88.750 61.580 ;
        RECT 88.890 61.320 89.210 61.580 ;
        RECT 73.710 61.040 82.220 61.180 ;
        RECT 59.935 60.995 60.225 61.040 ;
        RECT 62.455 60.995 62.745 61.040 ;
        RECT 63.645 60.995 63.935 61.040 ;
        RECT 73.710 60.980 74.030 61.040 ;
        RECT 85.670 60.980 85.990 61.240 ;
        RECT 86.145 60.995 86.435 61.225 ;
        RECT 16.210 60.840 16.530 60.900 ;
        RECT 24.990 60.840 25.280 60.885 ;
        RECT 27.090 60.840 27.380 60.885 ;
        RECT 28.660 60.840 28.950 60.885 ;
        RECT 16.210 60.700 21.730 60.840 ;
        RECT 16.210 60.640 16.530 60.700 ;
        RECT 18.065 60.500 18.355 60.545 ;
        RECT 18.510 60.500 18.830 60.560 ;
        RECT 18.065 60.360 18.830 60.500 ;
        RECT 21.590 60.500 21.730 60.700 ;
        RECT 24.990 60.700 28.950 60.840 ;
        RECT 24.990 60.655 25.280 60.700 ;
        RECT 27.090 60.655 27.380 60.700 ;
        RECT 28.660 60.655 28.950 60.700 ;
        RECT 32.350 60.840 32.640 60.885 ;
        RECT 34.450 60.840 34.740 60.885 ;
        RECT 36.020 60.840 36.310 60.885 ;
        RECT 32.350 60.700 36.310 60.840 ;
        RECT 32.350 60.655 32.640 60.700 ;
        RECT 34.450 60.655 34.740 60.700 ;
        RECT 36.020 60.655 36.310 60.700 ;
        RECT 42.930 60.840 43.220 60.885 ;
        RECT 45.030 60.840 45.320 60.885 ;
        RECT 46.600 60.840 46.890 60.885 ;
        RECT 42.930 60.700 46.890 60.840 ;
        RECT 42.930 60.655 43.220 60.700 ;
        RECT 45.030 60.655 45.320 60.700 ;
        RECT 46.600 60.655 46.890 60.700 ;
        RECT 60.370 60.840 60.660 60.885 ;
        RECT 61.940 60.840 62.230 60.885 ;
        RECT 64.040 60.840 64.330 60.885 ;
        RECT 60.370 60.700 64.330 60.840 ;
        RECT 60.370 60.655 60.660 60.700 ;
        RECT 61.940 60.655 62.230 60.700 ;
        RECT 64.040 60.655 64.330 60.700 ;
        RECT 77.390 60.840 77.710 60.900 ;
        RECT 86.220 60.840 86.360 60.995 ;
        RECT 77.390 60.700 86.360 60.840 ;
        RECT 77.390 60.640 77.710 60.700 ;
        RECT 89.810 60.640 90.130 60.900 ;
        RECT 27.710 60.500 28.030 60.560 ;
        RECT 31.405 60.500 31.695 60.545 ;
        RECT 35.530 60.500 35.850 60.560 ;
        RECT 21.590 60.360 35.850 60.500 ;
        RECT 18.065 60.315 18.355 60.360 ;
        RECT 18.510 60.300 18.830 60.360 ;
        RECT 27.710 60.300 28.030 60.360 ;
        RECT 31.405 60.315 31.695 60.360 ;
        RECT 35.530 60.300 35.850 60.360 ;
        RECT 69.125 60.500 69.415 60.545 ;
        RECT 70.030 60.500 70.350 60.560 ;
        RECT 69.125 60.360 70.350 60.500 ;
        RECT 69.125 60.315 69.415 60.360 ;
        RECT 70.030 60.300 70.350 60.360 ;
        RECT 73.710 60.500 74.030 60.560 ;
        RECT 80.610 60.500 80.930 60.560 ;
        RECT 73.710 60.360 80.930 60.500 ;
        RECT 73.710 60.300 74.030 60.360 ;
        RECT 80.610 60.300 80.930 60.360 ;
        RECT 83.370 60.300 83.690 60.560 ;
        RECT 13.380 59.680 92.040 60.160 ;
        RECT 13.450 59.480 13.770 59.540 ;
        RECT 15.305 59.480 15.595 59.525 ;
        RECT 13.450 59.340 15.595 59.480 ;
        RECT 13.450 59.280 13.770 59.340 ;
        RECT 15.305 59.295 15.595 59.340 ;
        RECT 22.650 59.480 22.970 59.540 ;
        RECT 26.330 59.480 26.650 59.540 ;
        RECT 22.650 59.340 26.650 59.480 ;
        RECT 22.650 59.280 22.970 59.340 ;
        RECT 26.330 59.280 26.650 59.340 ;
        RECT 28.170 59.480 28.490 59.540 ;
        RECT 28.645 59.480 28.935 59.525 ;
        RECT 28.170 59.340 28.935 59.480 ;
        RECT 28.170 59.280 28.490 59.340 ;
        RECT 28.645 59.295 28.935 59.340 ;
        RECT 32.785 59.480 33.075 59.525 ;
        RECT 33.230 59.480 33.550 59.540 ;
        RECT 32.785 59.340 33.550 59.480 ;
        RECT 32.785 59.295 33.075 59.340 ;
        RECT 33.230 59.280 33.550 59.340 ;
        RECT 42.445 59.480 42.735 59.525 ;
        RECT 42.890 59.480 43.210 59.540 ;
        RECT 42.445 59.340 43.210 59.480 ;
        RECT 42.445 59.295 42.735 59.340 ;
        RECT 42.890 59.280 43.210 59.340 ;
        RECT 49.790 59.480 50.110 59.540 ;
        RECT 50.725 59.480 51.015 59.525 ;
        RECT 49.790 59.340 51.015 59.480 ;
        RECT 49.790 59.280 50.110 59.340 ;
        RECT 50.725 59.295 51.015 59.340 ;
        RECT 56.245 59.480 56.535 59.525 ;
        RECT 57.610 59.480 57.930 59.540 ;
        RECT 56.245 59.340 57.930 59.480 ;
        RECT 56.245 59.295 56.535 59.340 ;
        RECT 57.610 59.280 57.930 59.340 ;
        RECT 66.810 59.480 67.130 59.540 ;
        RECT 72.330 59.480 72.650 59.540 ;
        RECT 66.810 59.340 72.650 59.480 ;
        RECT 66.810 59.280 67.130 59.340 ;
        RECT 72.330 59.280 72.650 59.340 ;
        RECT 72.790 59.480 73.110 59.540 ;
        RECT 76.930 59.480 77.250 59.540 ;
        RECT 72.790 59.340 77.250 59.480 ;
        RECT 72.790 59.280 73.110 59.340 ;
        RECT 76.930 59.280 77.250 59.340 ;
        RECT 77.390 59.280 77.710 59.540 ;
        RECT 81.085 59.480 81.375 59.525 ;
        RECT 85.670 59.480 85.990 59.540 ;
        RECT 81.085 59.340 85.990 59.480 ;
        RECT 81.085 59.295 81.375 59.340 ;
        RECT 85.670 59.280 85.990 59.340 ;
        RECT 87.970 59.480 88.290 59.540 ;
        RECT 88.905 59.480 89.195 59.525 ;
        RECT 87.970 59.340 89.195 59.480 ;
        RECT 87.970 59.280 88.290 59.340 ;
        RECT 88.905 59.295 89.195 59.340 ;
        RECT 17.170 59.140 17.460 59.185 ;
        RECT 19.270 59.140 19.560 59.185 ;
        RECT 20.840 59.140 21.130 59.185 ;
        RECT 17.170 59.000 21.130 59.140 ;
        RECT 17.170 58.955 17.460 59.000 ;
        RECT 19.270 58.955 19.560 59.000 ;
        RECT 20.840 58.955 21.130 59.000 ;
        RECT 22.190 59.140 22.510 59.200 ;
        RECT 23.585 59.140 23.875 59.185 ;
        RECT 24.950 59.140 25.270 59.200 ;
        RECT 30.930 59.140 31.250 59.200 ;
        RECT 22.190 59.000 25.270 59.140 ;
        RECT 22.190 58.940 22.510 59.000 ;
        RECT 23.585 58.955 23.875 59.000 ;
        RECT 24.950 58.940 25.270 59.000 ;
        RECT 30.000 59.000 31.250 59.140 ;
        RECT 17.565 58.800 17.855 58.845 ;
        RECT 18.755 58.800 19.045 58.845 ;
        RECT 21.275 58.800 21.565 58.845 ;
        RECT 17.565 58.660 21.565 58.800 ;
        RECT 17.565 58.615 17.855 58.660 ;
        RECT 18.755 58.615 19.045 58.660 ;
        RECT 21.275 58.615 21.565 58.660 ;
        RECT 16.225 58.275 16.515 58.505 ;
        RECT 16.300 58.120 16.440 58.275 ;
        RECT 16.670 58.260 16.990 58.520 ;
        RECT 22.190 58.460 22.510 58.520 ;
        RECT 17.680 58.320 22.510 58.460 ;
        RECT 17.680 58.120 17.820 58.320 ;
        RECT 22.190 58.260 22.510 58.320 ;
        RECT 26.790 58.260 27.110 58.520 ;
        RECT 27.710 58.260 28.030 58.520 ;
        RECT 29.565 58.460 29.855 58.505 ;
        RECT 30.000 58.460 30.140 59.000 ;
        RECT 30.930 58.940 31.250 59.000 ;
        RECT 35.570 59.140 35.860 59.185 ;
        RECT 37.670 59.140 37.960 59.185 ;
        RECT 39.240 59.140 39.530 59.185 ;
        RECT 35.570 59.000 39.530 59.140 ;
        RECT 35.570 58.955 35.860 59.000 ;
        RECT 37.670 58.955 37.960 59.000 ;
        RECT 39.240 58.955 39.530 59.000 ;
        RECT 40.590 59.140 40.910 59.200 ;
        RECT 65.430 59.140 65.750 59.200 ;
        RECT 73.250 59.140 73.570 59.200 ;
        RECT 82.490 59.140 82.780 59.185 ;
        RECT 84.590 59.140 84.880 59.185 ;
        RECT 86.160 59.140 86.450 59.185 ;
        RECT 40.590 59.000 68.420 59.140 ;
        RECT 40.590 58.940 40.910 59.000 ;
        RECT 65.430 58.940 65.750 59.000 ;
        RECT 31.850 58.800 32.170 58.860 ;
        RECT 30.560 58.660 32.170 58.800 ;
        RECT 30.560 58.505 30.700 58.660 ;
        RECT 31.850 58.600 32.170 58.660 ;
        RECT 35.965 58.800 36.255 58.845 ;
        RECT 37.155 58.800 37.445 58.845 ;
        RECT 39.675 58.800 39.965 58.845 ;
        RECT 35.965 58.660 39.965 58.800 ;
        RECT 35.965 58.615 36.255 58.660 ;
        RECT 37.155 58.615 37.445 58.660 ;
        RECT 39.675 58.615 39.965 58.660 ;
        RECT 45.665 58.800 45.955 58.845 ;
        RECT 47.490 58.800 47.810 58.860 ;
        RECT 45.665 58.660 47.810 58.800 ;
        RECT 45.665 58.615 45.955 58.660 ;
        RECT 47.490 58.600 47.810 58.660 ;
        RECT 48.425 58.800 48.715 58.845 ;
        RECT 58.070 58.800 58.390 58.860 ;
        RECT 58.545 58.800 58.835 58.845 ;
        RECT 48.425 58.660 57.840 58.800 ;
        RECT 48.425 58.615 48.715 58.660 ;
        RECT 28.215 58.320 30.140 58.460 ;
        RECT 18.050 58.165 18.370 58.180 ;
        RECT 16.300 57.980 17.820 58.120 ;
        RECT 18.020 57.935 18.370 58.165 ;
        RECT 18.050 57.920 18.370 57.935 ;
        RECT 18.970 58.120 19.290 58.180 ;
        RECT 23.110 58.120 23.430 58.180 ;
        RECT 28.215 58.120 28.355 58.320 ;
        RECT 29.565 58.275 29.855 58.320 ;
        RECT 30.485 58.275 30.775 58.505 ;
        RECT 30.945 58.275 31.235 58.505 ;
        RECT 31.405 58.460 31.695 58.505 ;
        RECT 32.310 58.460 32.630 58.520 ;
        RECT 31.405 58.320 32.630 58.460 ;
        RECT 31.405 58.275 31.695 58.320 ;
        RECT 18.970 57.980 28.355 58.120 ;
        RECT 29.090 58.120 29.410 58.180 ;
        RECT 31.020 58.120 31.160 58.275 ;
        RECT 32.310 58.260 32.630 58.320 ;
        RECT 35.085 58.460 35.375 58.505 ;
        RECT 41.050 58.460 41.370 58.520 ;
        RECT 35.085 58.320 41.370 58.460 ;
        RECT 35.085 58.275 35.375 58.320 ;
        RECT 41.050 58.260 41.370 58.320 ;
        RECT 48.885 58.460 49.175 58.505 ;
        RECT 51.170 58.460 51.490 58.520 ;
        RECT 48.885 58.320 51.490 58.460 ;
        RECT 57.700 58.460 57.840 58.660 ;
        RECT 58.070 58.660 58.835 58.800 ;
        RECT 58.070 58.600 58.390 58.660 ;
        RECT 58.545 58.615 58.835 58.660 ;
        RECT 59.465 58.800 59.755 58.845 ;
        RECT 60.370 58.800 60.690 58.860 ;
        RECT 67.730 58.800 68.050 58.860 ;
        RECT 59.465 58.660 60.690 58.800 ;
        RECT 59.465 58.615 59.755 58.660 ;
        RECT 60.370 58.600 60.690 58.660 ;
        RECT 67.360 58.660 68.050 58.800 ;
        RECT 68.280 58.800 68.420 59.000 ;
        RECT 69.200 59.000 73.570 59.140 ;
        RECT 69.200 58.800 69.340 59.000 ;
        RECT 73.250 58.940 73.570 59.000 ;
        RECT 73.800 59.000 78.540 59.140 ;
        RECT 68.280 58.660 69.340 58.800 ;
        RECT 69.585 58.800 69.875 58.845 ;
        RECT 73.800 58.800 73.940 59.000 ;
        RECT 69.585 58.660 73.940 58.800 ;
        RECT 74.170 58.800 74.490 58.860 ;
        RECT 75.105 58.800 75.395 58.845 ;
        RECT 74.170 58.660 75.395 58.800 ;
        RECT 64.510 58.460 64.830 58.520 ;
        RECT 57.700 58.320 64.830 58.460 ;
        RECT 48.885 58.275 49.175 58.320 ;
        RECT 51.170 58.260 51.490 58.320 ;
        RECT 64.510 58.260 64.830 58.320 ;
        RECT 66.810 58.260 67.130 58.520 ;
        RECT 67.360 58.505 67.500 58.660 ;
        RECT 67.730 58.600 68.050 58.660 ;
        RECT 69.585 58.615 69.875 58.660 ;
        RECT 74.170 58.600 74.490 58.660 ;
        RECT 75.105 58.615 75.395 58.660 ;
        RECT 75.550 58.600 75.870 58.860 ;
        RECT 67.285 58.275 67.575 58.505 ;
        RECT 68.650 58.260 68.970 58.520 ;
        RECT 69.110 58.260 69.430 58.520 ;
        RECT 70.045 58.460 70.335 58.505 ;
        RECT 70.490 58.460 70.810 58.520 ;
        RECT 70.045 58.320 70.810 58.460 ;
        RECT 70.045 58.275 70.335 58.320 ;
        RECT 29.090 57.980 31.160 58.120 ;
        RECT 36.420 58.120 36.710 58.165 ;
        RECT 39.210 58.120 39.530 58.180 ;
        RECT 36.420 57.980 39.530 58.120 ;
        RECT 18.970 57.920 19.290 57.980 ;
        RECT 23.110 57.920 23.430 57.980 ;
        RECT 29.090 57.920 29.410 57.980 ;
        RECT 36.420 57.935 36.710 57.980 ;
        RECT 39.210 57.920 39.530 57.980 ;
        RECT 44.745 58.120 45.035 58.165 ;
        RECT 55.310 58.120 55.630 58.180 ;
        RECT 44.745 57.980 55.630 58.120 ;
        RECT 44.745 57.935 45.035 57.980 ;
        RECT 55.310 57.920 55.630 57.980 ;
        RECT 67.730 57.920 68.050 58.180 ;
        RECT 19.430 57.780 19.750 57.840 ;
        RECT 21.270 57.780 21.590 57.840 ;
        RECT 19.430 57.640 21.590 57.780 ;
        RECT 19.430 57.580 19.750 57.640 ;
        RECT 21.270 57.580 21.590 57.640 ;
        RECT 28.630 57.780 28.950 57.840 ;
        RECT 31.390 57.780 31.710 57.840 ;
        RECT 28.630 57.640 31.710 57.780 ;
        RECT 28.630 57.580 28.950 57.640 ;
        RECT 31.390 57.580 31.710 57.640 ;
        RECT 41.985 57.780 42.275 57.825 ;
        RECT 44.270 57.780 44.590 57.840 ;
        RECT 41.985 57.640 44.590 57.780 ;
        RECT 41.985 57.595 42.275 57.640 ;
        RECT 44.270 57.580 44.590 57.640 ;
        RECT 58.085 57.780 58.375 57.825 ;
        RECT 60.370 57.780 60.690 57.840 ;
        RECT 58.085 57.640 60.690 57.780 ;
        RECT 58.085 57.595 58.375 57.640 ;
        RECT 60.370 57.580 60.690 57.640 ;
        RECT 65.905 57.780 66.195 57.825 ;
        RECT 66.350 57.780 66.670 57.840 ;
        RECT 65.905 57.640 66.670 57.780 ;
        RECT 65.905 57.595 66.195 57.640 ;
        RECT 66.350 57.580 66.670 57.640 ;
        RECT 69.110 57.780 69.430 57.840 ;
        RECT 70.120 57.780 70.260 58.275 ;
        RECT 70.490 58.260 70.810 58.320 ;
        RECT 70.950 58.260 71.270 58.520 ;
        RECT 71.410 58.260 71.730 58.520 ;
        RECT 71.885 58.275 72.175 58.505 ;
        RECT 71.040 58.120 71.180 58.260 ;
        RECT 71.960 58.120 72.100 58.275 ;
        RECT 72.330 58.260 72.650 58.520 ;
        RECT 72.790 58.260 73.110 58.520 ;
        RECT 73.710 58.260 74.030 58.520 ;
        RECT 74.645 58.460 74.935 58.505 ;
        RECT 76.010 58.460 76.330 58.520 ;
        RECT 74.645 58.320 76.330 58.460 ;
        RECT 74.645 58.275 74.935 58.320 ;
        RECT 76.010 58.260 76.330 58.320 ;
        RECT 76.470 58.260 76.790 58.520 ;
        RECT 78.400 58.505 78.540 59.000 ;
        RECT 82.490 59.000 86.450 59.140 ;
        RECT 82.490 58.955 82.780 59.000 ;
        RECT 84.590 58.955 84.880 59.000 ;
        RECT 86.160 58.955 86.450 59.000 ;
        RECT 81.530 58.800 81.850 58.860 ;
        RECT 82.005 58.800 82.295 58.845 ;
        RECT 81.530 58.660 82.295 58.800 ;
        RECT 81.530 58.600 81.850 58.660 ;
        RECT 82.005 58.615 82.295 58.660 ;
        RECT 82.885 58.800 83.175 58.845 ;
        RECT 84.075 58.800 84.365 58.845 ;
        RECT 86.595 58.800 86.885 58.845 ;
        RECT 82.885 58.660 86.885 58.800 ;
        RECT 82.885 58.615 83.175 58.660 ;
        RECT 84.075 58.615 84.365 58.660 ;
        RECT 86.595 58.615 86.885 58.660 ;
        RECT 78.325 58.275 78.615 58.505 ;
        RECT 78.770 58.460 79.090 58.520 ;
        RECT 79.245 58.460 79.535 58.505 ;
        RECT 78.770 58.320 79.535 58.460 ;
        RECT 78.770 58.260 79.090 58.320 ;
        RECT 79.245 58.275 79.535 58.320 ;
        RECT 80.150 58.260 80.470 58.520 ;
        RECT 83.370 58.505 83.690 58.520 ;
        RECT 83.340 58.460 83.690 58.505 ;
        RECT 83.175 58.320 83.690 58.460 ;
        RECT 88.980 58.460 89.120 59.295 ;
        RECT 89.350 59.280 89.670 59.540 ;
        RECT 90.285 58.460 90.575 58.505 ;
        RECT 88.980 58.320 90.575 58.460 ;
        RECT 83.340 58.275 83.690 58.320 ;
        RECT 90.285 58.275 90.575 58.320 ;
        RECT 83.370 58.260 83.690 58.275 ;
        RECT 71.040 57.980 72.100 58.120 ;
        RECT 73.250 58.120 73.570 58.180 ;
        RECT 79.705 58.120 79.995 58.165 ;
        RECT 73.250 57.980 79.995 58.120 ;
        RECT 73.250 57.920 73.570 57.980 ;
        RECT 79.705 57.935 79.995 57.980 ;
        RECT 69.110 57.640 70.260 57.780 ;
        RECT 70.505 57.780 70.795 57.825 ;
        RECT 70.950 57.780 71.270 57.840 ;
        RECT 70.505 57.640 71.270 57.780 ;
        RECT 69.110 57.580 69.430 57.640 ;
        RECT 70.505 57.595 70.795 57.640 ;
        RECT 70.950 57.580 71.270 57.640 ;
        RECT 71.410 57.780 71.730 57.840 ;
        RECT 76.010 57.780 76.330 57.840 ;
        RECT 71.410 57.640 76.330 57.780 ;
        RECT 71.410 57.580 71.730 57.640 ;
        RECT 76.010 57.580 76.330 57.640 ;
        RECT 13.380 56.960 92.040 57.440 ;
        RECT 16.225 56.760 16.515 56.805 ;
        RECT 18.050 56.760 18.370 56.820 ;
        RECT 16.225 56.620 18.370 56.760 ;
        RECT 16.225 56.575 16.515 56.620 ;
        RECT 18.050 56.560 18.370 56.620 ;
        RECT 21.730 56.760 22.050 56.820 ;
        RECT 26.345 56.760 26.635 56.805 ;
        RECT 36.910 56.760 37.230 56.820 ;
        RECT 21.730 56.620 26.100 56.760 ;
        RECT 21.730 56.560 22.050 56.620 ;
        RECT 20.810 56.420 21.130 56.480 ;
        RECT 18.140 56.280 21.130 56.420 ;
        RECT 25.960 56.420 26.100 56.620 ;
        RECT 26.345 56.620 37.230 56.760 ;
        RECT 26.345 56.575 26.635 56.620 ;
        RECT 36.910 56.560 37.230 56.620 ;
        RECT 39.210 56.760 39.530 56.820 ;
        RECT 39.685 56.760 39.975 56.805 ;
        RECT 39.210 56.620 39.975 56.760 ;
        RECT 39.210 56.560 39.530 56.620 ;
        RECT 39.685 56.575 39.975 56.620 ;
        RECT 47.030 56.760 47.350 56.820 ;
        RECT 47.505 56.760 47.795 56.805 ;
        RECT 47.030 56.620 47.795 56.760 ;
        RECT 47.030 56.560 47.350 56.620 ;
        RECT 47.505 56.575 47.795 56.620 ;
        RECT 68.650 56.560 68.970 56.820 ;
        RECT 72.330 56.760 72.650 56.820 ;
        RECT 69.660 56.620 70.260 56.760 ;
        RECT 27.250 56.420 27.570 56.480 ;
        RECT 29.090 56.420 29.410 56.480 ;
        RECT 25.960 56.280 29.410 56.420 ;
        RECT 18.140 56.125 18.280 56.280 ;
        RECT 20.810 56.220 21.130 56.280 ;
        RECT 27.250 56.220 27.570 56.280 ;
        RECT 17.605 55.895 17.895 56.125 ;
        RECT 18.065 55.895 18.355 56.125 ;
        RECT 17.680 55.400 17.820 55.895 ;
        RECT 18.510 55.880 18.830 56.140 ;
        RECT 18.970 56.080 19.290 56.140 ;
        RECT 19.445 56.080 19.735 56.125 ;
        RECT 18.970 55.940 19.735 56.080 ;
        RECT 18.970 55.880 19.290 55.940 ;
        RECT 19.445 55.895 19.735 55.940 ;
        RECT 19.890 56.080 20.210 56.140 ;
        RECT 19.890 56.030 20.580 56.080 ;
        RECT 21.285 56.030 21.575 56.125 ;
        RECT 19.890 55.940 21.575 56.030 ;
        RECT 19.890 55.880 20.210 55.940 ;
        RECT 20.440 55.895 21.575 55.940 ;
        RECT 20.440 55.890 21.500 55.895 ;
        RECT 21.715 55.880 22.035 56.140 ;
        RECT 22.310 56.110 22.600 56.155 ;
        RECT 22.310 55.970 22.880 56.110 ;
        RECT 22.310 55.925 22.600 55.970 ;
        RECT 22.740 55.460 22.880 55.970 ;
        RECT 23.110 55.880 23.430 56.140 ;
        RECT 23.585 55.895 23.875 56.125 ;
        RECT 24.045 56.080 24.335 56.125 ;
        RECT 24.490 56.080 24.810 56.140 ;
        RECT 24.045 55.940 24.810 56.080 ;
        RECT 24.045 55.895 24.335 55.940 ;
        RECT 17.680 55.260 20.580 55.400 ;
        RECT 20.440 55.120 20.580 55.260 ;
        RECT 22.650 55.200 22.970 55.460 ;
        RECT 23.660 55.400 23.800 55.895 ;
        RECT 24.490 55.880 24.810 55.940 ;
        RECT 24.950 55.880 25.270 56.140 ;
        RECT 25.410 55.880 25.730 56.140 ;
        RECT 26.330 56.080 26.650 56.140 ;
        RECT 28.260 56.125 28.400 56.280 ;
        RECT 29.090 56.220 29.410 56.280 ;
        RECT 30.025 56.420 30.315 56.465 ;
        RECT 31.710 56.420 32.000 56.465 ;
        RECT 30.025 56.280 32.000 56.420 ;
        RECT 30.025 56.235 30.315 56.280 ;
        RECT 31.710 56.235 32.000 56.280 ;
        RECT 35.530 56.420 35.850 56.480 ;
        RECT 55.310 56.420 55.630 56.480 ;
        RECT 69.660 56.465 69.800 56.620 ;
        RECT 35.530 56.280 49.100 56.420 ;
        RECT 35.530 56.220 35.850 56.280 ;
        RECT 26.805 56.080 27.095 56.125 ;
        RECT 26.330 55.940 27.095 56.080 ;
        RECT 26.330 55.880 26.650 55.940 ;
        RECT 26.805 55.895 27.095 55.940 ;
        RECT 27.725 55.895 28.015 56.125 ;
        RECT 28.185 55.895 28.475 56.125 ;
        RECT 24.950 55.400 25.270 55.460 ;
        RECT 23.660 55.260 25.270 55.400 ;
        RECT 24.950 55.200 25.270 55.260 ;
        RECT 19.890 54.860 20.210 55.120 ;
        RECT 20.350 55.060 20.670 55.120 ;
        RECT 24.030 55.060 24.350 55.120 ;
        RECT 20.350 54.920 24.350 55.060 ;
        RECT 27.800 55.060 27.940 55.895 ;
        RECT 28.630 55.880 28.950 56.140 ;
        RECT 30.485 56.080 30.775 56.125 ;
        RECT 30.930 56.080 31.250 56.140 ;
        RECT 30.485 55.940 31.250 56.080 ;
        RECT 30.485 55.895 30.775 55.940 ;
        RECT 30.930 55.880 31.250 55.940 ;
        RECT 41.525 56.080 41.815 56.125 ;
        RECT 43.825 56.080 44.115 56.125 ;
        RECT 41.525 55.940 44.115 56.080 ;
        RECT 41.525 55.895 41.815 55.940 ;
        RECT 43.825 55.895 44.115 55.940 ;
        RECT 44.270 56.080 44.590 56.140 ;
        RECT 46.585 56.080 46.875 56.125 ;
        RECT 44.270 55.940 46.875 56.080 ;
        RECT 44.270 55.880 44.590 55.940 ;
        RECT 46.585 55.895 46.875 55.940 ;
        RECT 48.410 55.880 48.730 56.140 ;
        RECT 48.960 56.125 49.100 56.280 ;
        RECT 55.310 56.280 65.660 56.420 ;
        RECT 55.310 56.220 55.630 56.280 ;
        RECT 48.885 55.895 49.175 56.125 ;
        RECT 49.805 55.895 50.095 56.125 ;
        RECT 31.365 55.740 31.655 55.785 ;
        RECT 32.555 55.740 32.845 55.785 ;
        RECT 35.075 55.740 35.365 55.785 ;
        RECT 31.365 55.600 35.365 55.740 ;
        RECT 31.365 55.555 31.655 55.600 ;
        RECT 32.555 55.555 32.845 55.600 ;
        RECT 35.075 55.555 35.365 55.600 ;
        RECT 41.970 55.540 42.290 55.800 ;
        RECT 42.905 55.740 43.195 55.785 ;
        RECT 49.330 55.740 49.650 55.800 ;
        RECT 42.905 55.600 49.650 55.740 ;
        RECT 49.880 55.740 50.020 55.895 ;
        RECT 50.250 55.880 50.570 56.140 ;
        RECT 65.520 56.125 65.660 56.280 ;
        RECT 69.585 56.235 69.875 56.465 ;
        RECT 54.405 56.080 54.695 56.125 ;
        RECT 56.705 56.080 56.995 56.125 ;
        RECT 54.405 55.940 56.995 56.080 ;
        RECT 54.405 55.895 54.695 55.940 ;
        RECT 56.705 55.895 56.995 55.940 ;
        RECT 65.445 55.895 65.735 56.125 ;
        RECT 69.110 55.880 69.430 56.140 ;
        RECT 70.120 56.080 70.260 56.620 ;
        RECT 70.580 56.620 72.650 56.760 ;
        RECT 70.580 56.465 70.720 56.620 ;
        RECT 72.330 56.560 72.650 56.620 ;
        RECT 77.850 56.560 78.170 56.820 ;
        RECT 70.505 56.235 70.795 56.465 ;
        RECT 70.965 56.420 71.255 56.465 ;
        RECT 71.410 56.420 71.730 56.480 ;
        RECT 74.170 56.420 74.490 56.480 ;
        RECT 76.930 56.420 77.250 56.480 ;
        RECT 79.690 56.420 80.010 56.480 ;
        RECT 70.965 56.280 71.730 56.420 ;
        RECT 70.965 56.235 71.255 56.280 ;
        RECT 71.410 56.220 71.730 56.280 ;
        RECT 72.420 56.280 74.490 56.420 ;
        RECT 71.870 56.080 72.190 56.140 ;
        RECT 72.420 56.125 72.560 56.280 ;
        RECT 74.170 56.220 74.490 56.280 ;
        RECT 75.180 56.280 80.010 56.420 ;
        RECT 70.120 55.940 72.190 56.080 ;
        RECT 71.870 55.880 72.190 55.940 ;
        RECT 72.345 55.895 72.635 56.125 ;
        RECT 72.790 56.080 73.110 56.140 ;
        RECT 73.725 56.080 74.015 56.125 ;
        RECT 72.790 55.940 74.015 56.080 ;
        RECT 72.790 55.880 73.110 55.940 ;
        RECT 73.725 55.895 74.015 55.940 ;
        RECT 53.470 55.740 53.790 55.800 ;
        RECT 49.880 55.600 53.790 55.740 ;
        RECT 42.905 55.555 43.195 55.600 ;
        RECT 49.330 55.540 49.650 55.600 ;
        RECT 53.470 55.540 53.790 55.600 ;
        RECT 54.850 55.540 55.170 55.800 ;
        RECT 55.770 55.540 56.090 55.800 ;
        RECT 58.990 55.740 59.310 55.800 ;
        RECT 59.465 55.740 59.755 55.785 ;
        RECT 58.990 55.600 59.755 55.740 ;
        RECT 58.990 55.540 59.310 55.600 ;
        RECT 59.465 55.555 59.755 55.600 ;
        RECT 60.370 55.740 60.690 55.800 ;
        RECT 63.605 55.740 63.895 55.785 ;
        RECT 60.370 55.600 63.895 55.740 ;
        RECT 60.370 55.540 60.690 55.600 ;
        RECT 63.605 55.555 63.895 55.600 ;
        RECT 65.890 55.740 66.210 55.800 ;
        RECT 65.890 55.600 70.030 55.740 ;
        RECT 65.890 55.540 66.210 55.600 ;
        RECT 30.970 55.400 31.260 55.445 ;
        RECT 33.070 55.400 33.360 55.445 ;
        RECT 34.640 55.400 34.930 55.445 ;
        RECT 30.970 55.260 34.930 55.400 ;
        RECT 30.970 55.215 31.260 55.260 ;
        RECT 33.070 55.215 33.360 55.260 ;
        RECT 34.640 55.215 34.930 55.260 ;
        RECT 67.730 55.400 68.050 55.460 ;
        RECT 69.125 55.400 69.415 55.445 ;
        RECT 67.730 55.260 69.415 55.400 ;
        RECT 69.890 55.400 70.030 55.600 ;
        RECT 70.950 55.540 71.270 55.800 ;
        RECT 74.185 55.740 74.475 55.785 ;
        RECT 75.180 55.740 75.320 56.280 ;
        RECT 76.930 56.220 77.250 56.280 ;
        RECT 79.690 56.220 80.010 56.280 ;
        RECT 75.565 55.895 75.855 56.125 ;
        RECT 76.025 56.080 76.315 56.125 ;
        RECT 76.470 56.080 76.790 56.140 ;
        RECT 77.405 56.080 77.695 56.125 ;
        RECT 76.025 55.940 76.790 56.080 ;
        RECT 76.025 55.895 76.315 55.940 ;
        RECT 74.185 55.600 75.320 55.740 ;
        RECT 74.185 55.555 74.475 55.600 ;
        RECT 75.640 55.400 75.780 55.895 ;
        RECT 76.470 55.880 76.790 55.940 ;
        RECT 77.020 55.940 77.695 56.080 ;
        RECT 77.020 55.445 77.160 55.940 ;
        RECT 77.405 55.895 77.695 55.940 ;
        RECT 80.625 56.080 80.915 56.125 ;
        RECT 81.070 56.080 81.390 56.140 ;
        RECT 81.990 56.125 82.310 56.140 ;
        RECT 80.625 55.940 81.390 56.080 ;
        RECT 80.625 55.895 80.915 55.940 ;
        RECT 81.070 55.880 81.390 55.940 ;
        RECT 81.960 55.895 82.310 56.125 ;
        RECT 81.990 55.880 82.310 55.895 ;
        RECT 83.830 56.080 84.150 56.140 ;
        RECT 88.905 56.080 89.195 56.125 ;
        RECT 83.830 55.940 89.195 56.080 ;
        RECT 83.830 55.880 84.150 55.940 ;
        RECT 88.905 55.895 89.195 55.940 ;
        RECT 79.705 55.740 79.995 55.785 ;
        RECT 80.150 55.740 80.470 55.800 ;
        RECT 79.705 55.600 80.470 55.740 ;
        RECT 79.705 55.555 79.995 55.600 ;
        RECT 80.150 55.540 80.470 55.600 ;
        RECT 81.505 55.740 81.795 55.785 ;
        RECT 82.695 55.740 82.985 55.785 ;
        RECT 85.215 55.740 85.505 55.785 ;
        RECT 81.505 55.600 85.505 55.740 ;
        RECT 81.505 55.555 81.795 55.600 ;
        RECT 82.695 55.555 82.985 55.600 ;
        RECT 85.215 55.555 85.505 55.600 ;
        RECT 69.890 55.260 75.780 55.400 ;
        RECT 67.730 55.200 68.050 55.260 ;
        RECT 69.125 55.215 69.415 55.260 ;
        RECT 76.945 55.215 77.235 55.445 ;
        RECT 81.110 55.400 81.400 55.445 ;
        RECT 83.210 55.400 83.500 55.445 ;
        RECT 84.780 55.400 85.070 55.445 ;
        RECT 81.110 55.260 85.070 55.400 ;
        RECT 81.110 55.215 81.400 55.260 ;
        RECT 83.210 55.215 83.500 55.260 ;
        RECT 84.780 55.215 85.070 55.260 ;
        RECT 31.390 55.060 31.710 55.120 ;
        RECT 27.800 54.920 31.710 55.060 ;
        RECT 20.350 54.860 20.670 54.920 ;
        RECT 24.030 54.860 24.350 54.920 ;
        RECT 31.390 54.860 31.710 54.920 ;
        RECT 35.070 55.060 35.390 55.120 ;
        RECT 37.385 55.060 37.675 55.105 ;
        RECT 35.070 54.920 37.675 55.060 ;
        RECT 35.070 54.860 35.390 54.920 ;
        RECT 37.385 54.875 37.675 54.920 ;
        RECT 52.550 54.860 52.870 55.120 ;
        RECT 60.830 54.860 61.150 55.120 ;
        RECT 70.030 55.060 70.350 55.120 ;
        RECT 71.885 55.060 72.175 55.105 ;
        RECT 75.550 55.060 75.870 55.120 ;
        RECT 70.030 54.920 75.870 55.060 ;
        RECT 70.030 54.860 70.350 54.920 ;
        RECT 71.885 54.875 72.175 54.920 ;
        RECT 75.550 54.860 75.870 54.920 ;
        RECT 78.785 55.060 79.075 55.105 ;
        RECT 85.210 55.060 85.530 55.120 ;
        RECT 78.785 54.920 85.530 55.060 ;
        RECT 78.785 54.875 79.075 54.920 ;
        RECT 85.210 54.860 85.530 54.920 ;
        RECT 87.510 54.860 87.830 55.120 ;
        RECT 89.810 54.860 90.130 55.120 ;
        RECT 13.380 54.240 92.040 54.720 ;
        RECT 16.685 54.040 16.975 54.085 ;
        RECT 22.650 54.040 22.970 54.100 ;
        RECT 34.625 54.040 34.915 54.085 ;
        RECT 41.970 54.040 42.290 54.100 ;
        RECT 16.685 53.900 22.970 54.040 ;
        RECT 16.685 53.855 16.975 53.900 ;
        RECT 22.650 53.840 22.970 53.900 ;
        RECT 31.940 53.900 34.380 54.040 ;
        RECT 17.630 53.700 17.920 53.745 ;
        RECT 19.730 53.700 20.020 53.745 ;
        RECT 21.300 53.700 21.590 53.745 ;
        RECT 17.630 53.560 21.590 53.700 ;
        RECT 17.630 53.515 17.920 53.560 ;
        RECT 19.730 53.515 20.020 53.560 ;
        RECT 21.300 53.515 21.590 53.560 ;
        RECT 16.670 53.360 16.990 53.420 ;
        RECT 17.145 53.360 17.435 53.405 ;
        RECT 16.670 53.220 17.435 53.360 ;
        RECT 16.670 53.160 16.990 53.220 ;
        RECT 17.145 53.175 17.435 53.220 ;
        RECT 18.025 53.360 18.315 53.405 ;
        RECT 19.215 53.360 19.505 53.405 ;
        RECT 21.735 53.360 22.025 53.405 ;
        RECT 18.025 53.220 22.025 53.360 ;
        RECT 18.025 53.175 18.315 53.220 ;
        RECT 19.215 53.175 19.505 53.220 ;
        RECT 21.735 53.175 22.025 53.220 ;
        RECT 17.220 53.020 17.360 53.175 ;
        RECT 25.410 53.020 25.730 53.080 ;
        RECT 31.940 53.065 32.080 53.900 ;
        RECT 34.240 53.360 34.380 53.900 ;
        RECT 34.625 53.900 42.290 54.040 ;
        RECT 34.625 53.855 34.915 53.900 ;
        RECT 41.970 53.840 42.290 53.900 ;
        RECT 48.885 54.040 49.175 54.085 ;
        RECT 54.850 54.040 55.170 54.100 ;
        RECT 48.885 53.900 55.170 54.040 ;
        RECT 48.885 53.855 49.175 53.900 ;
        RECT 54.850 53.840 55.170 53.900 ;
        RECT 55.310 54.040 55.630 54.100 ;
        RECT 55.310 53.900 58.300 54.040 ;
        RECT 55.310 53.840 55.630 53.900 ;
        RECT 53.970 53.700 54.260 53.745 ;
        RECT 56.070 53.700 56.360 53.745 ;
        RECT 57.640 53.700 57.930 53.745 ;
        RECT 53.970 53.560 57.930 53.700 ;
        RECT 58.160 53.700 58.300 53.900 ;
        RECT 60.370 53.840 60.690 54.100 ;
        RECT 64.510 54.040 64.830 54.100 ;
        RECT 68.205 54.040 68.495 54.085 ;
        RECT 81.990 54.040 82.310 54.100 ;
        RECT 82.465 54.040 82.755 54.085 ;
        RECT 64.510 53.900 81.760 54.040 ;
        RECT 64.510 53.840 64.830 53.900 ;
        RECT 68.205 53.855 68.495 53.900 ;
        RECT 60.845 53.700 61.135 53.745 ;
        RECT 58.160 53.560 61.135 53.700 ;
        RECT 53.970 53.515 54.260 53.560 ;
        RECT 56.070 53.515 56.360 53.560 ;
        RECT 57.640 53.515 57.930 53.560 ;
        RECT 60.845 53.515 61.135 53.560 ;
        RECT 63.590 53.700 63.880 53.745 ;
        RECT 65.160 53.700 65.450 53.745 ;
        RECT 67.260 53.700 67.550 53.745 ;
        RECT 63.590 53.560 67.550 53.700 ;
        RECT 63.590 53.515 63.880 53.560 ;
        RECT 65.160 53.515 65.450 53.560 ;
        RECT 67.260 53.515 67.550 53.560 ;
        RECT 70.950 53.700 71.240 53.745 ;
        RECT 72.520 53.700 72.810 53.745 ;
        RECT 74.620 53.700 74.910 53.745 ;
        RECT 70.950 53.560 74.910 53.700 ;
        RECT 70.950 53.515 71.240 53.560 ;
        RECT 72.520 53.515 72.810 53.560 ;
        RECT 74.620 53.515 74.910 53.560 ;
        RECT 76.010 53.500 76.330 53.760 ;
        RECT 81.070 53.500 81.390 53.760 ;
        RECT 54.365 53.360 54.655 53.405 ;
        RECT 55.555 53.360 55.845 53.405 ;
        RECT 58.075 53.360 58.365 53.405 ;
        RECT 32.860 53.220 33.920 53.360 ;
        RECT 34.240 53.220 54.160 53.360 ;
        RECT 17.220 52.880 21.730 53.020 ;
        RECT 14.830 52.480 15.150 52.740 ;
        RECT 15.765 52.495 16.055 52.725 ;
        RECT 18.480 52.680 18.770 52.725 ;
        RECT 19.890 52.680 20.210 52.740 ;
        RECT 18.480 52.540 20.210 52.680 ;
        RECT 21.590 52.680 21.730 52.880 ;
        RECT 25.410 52.880 31.620 53.020 ;
        RECT 25.410 52.820 25.730 52.880 ;
        RECT 26.805 52.680 27.095 52.725 ;
        RECT 28.630 52.680 28.950 52.740 ;
        RECT 21.590 52.540 28.950 52.680 ;
        RECT 31.480 52.680 31.620 52.880 ;
        RECT 31.865 52.835 32.155 53.065 ;
        RECT 32.310 52.820 32.630 53.080 ;
        RECT 32.860 52.680 33.000 53.220 ;
        RECT 33.780 53.065 33.920 53.220 ;
        RECT 33.245 52.835 33.535 53.065 ;
        RECT 33.705 53.020 33.995 53.065 ;
        RECT 48.410 53.020 48.730 53.080 ;
        RECT 49.790 53.020 50.110 53.080 ;
        RECT 33.705 52.880 50.110 53.020 ;
        RECT 33.705 52.835 33.995 52.880 ;
        RECT 31.480 52.540 33.000 52.680 ;
        RECT 18.480 52.495 18.770 52.540 ;
        RECT 15.840 52.340 15.980 52.495 ;
        RECT 19.890 52.480 20.210 52.540 ;
        RECT 26.805 52.495 27.095 52.540 ;
        RECT 28.630 52.480 28.950 52.540 ;
        RECT 16.210 52.340 16.530 52.400 ;
        RECT 24.045 52.340 24.335 52.385 ;
        RECT 33.320 52.340 33.460 52.835 ;
        RECT 48.410 52.820 48.730 52.880 ;
        RECT 49.790 52.820 50.110 52.880 ;
        RECT 50.265 52.835 50.555 53.065 ;
        RECT 51.185 52.835 51.475 53.065 ;
        RECT 34.610 52.680 34.930 52.740 ;
        RECT 50.340 52.680 50.480 52.835 ;
        RECT 34.610 52.540 50.480 52.680 ;
        RECT 34.610 52.480 34.930 52.540 ;
        RECT 15.840 52.200 33.460 52.340 ;
        RECT 51.260 52.340 51.400 52.835 ;
        RECT 51.630 52.820 51.950 53.080 ;
        RECT 53.485 52.835 53.775 53.065 ;
        RECT 54.020 53.020 54.160 53.220 ;
        RECT 54.365 53.220 58.365 53.360 ;
        RECT 54.365 53.175 54.655 53.220 ;
        RECT 55.555 53.175 55.845 53.220 ;
        RECT 58.075 53.175 58.365 53.220 ;
        RECT 63.155 53.360 63.445 53.405 ;
        RECT 65.675 53.360 65.965 53.405 ;
        RECT 66.865 53.360 67.155 53.405 ;
        RECT 63.155 53.220 67.155 53.360 ;
        RECT 63.155 53.175 63.445 53.220 ;
        RECT 65.675 53.175 65.965 53.220 ;
        RECT 66.865 53.175 67.155 53.220 ;
        RECT 70.515 53.360 70.805 53.405 ;
        RECT 73.035 53.360 73.325 53.405 ;
        RECT 74.225 53.360 74.515 53.405 ;
        RECT 70.515 53.220 74.515 53.360 ;
        RECT 70.515 53.175 70.805 53.220 ;
        RECT 73.035 53.175 73.325 53.220 ;
        RECT 74.225 53.175 74.515 53.220 ;
        RECT 75.105 53.360 75.395 53.405 ;
        RECT 81.160 53.360 81.300 53.500 ;
        RECT 81.620 53.405 81.760 53.900 ;
        RECT 81.990 53.900 82.755 54.040 ;
        RECT 81.990 53.840 82.310 53.900 ;
        RECT 82.465 53.855 82.755 53.900 ;
        RECT 75.105 53.220 81.300 53.360 ;
        RECT 75.105 53.175 75.395 53.220 ;
        RECT 81.545 53.175 81.835 53.405 ;
        RECT 61.290 53.020 61.610 53.080 ;
        RECT 54.020 52.880 61.610 53.020 ;
        RECT 53.560 52.680 53.700 52.835 ;
        RECT 61.290 52.820 61.610 52.880 ;
        RECT 66.350 53.065 66.670 53.080 ;
        RECT 66.350 53.020 66.700 53.065 ;
        RECT 67.745 53.020 68.035 53.065 ;
        RECT 75.180 53.020 75.320 53.175 ;
        RECT 84.750 53.160 85.070 53.420 ;
        RECT 85.210 53.160 85.530 53.420 ;
        RECT 87.510 53.360 87.830 53.420 ;
        RECT 89.365 53.360 89.655 53.405 ;
        RECT 90.270 53.360 90.590 53.420 ;
        RECT 87.510 53.220 90.590 53.360 ;
        RECT 87.510 53.160 87.830 53.220 ;
        RECT 89.365 53.175 89.655 53.220 ;
        RECT 90.270 53.160 90.590 53.220 ;
        RECT 66.350 52.880 66.865 53.020 ;
        RECT 67.745 52.880 75.320 53.020 ;
        RECT 66.350 52.835 66.700 52.880 ;
        RECT 67.745 52.835 68.035 52.880 ;
        RECT 66.350 52.820 66.670 52.835 ;
        RECT 75.550 52.820 75.870 53.080 ;
        RECT 76.485 53.020 76.775 53.065 ;
        RECT 76.930 53.020 77.250 53.080 ;
        RECT 76.485 52.880 77.250 53.020 ;
        RECT 76.485 52.835 76.775 52.880 ;
        RECT 76.930 52.820 77.250 52.880 ;
        RECT 53.930 52.680 54.250 52.740 ;
        RECT 53.560 52.540 54.250 52.680 ;
        RECT 53.930 52.480 54.250 52.540 ;
        RECT 54.820 52.680 55.110 52.725 ;
        RECT 58.530 52.680 58.850 52.740 ;
        RECT 54.820 52.540 58.850 52.680 ;
        RECT 54.820 52.495 55.110 52.540 ;
        RECT 58.530 52.480 58.850 52.540 ;
        RECT 71.410 52.680 71.730 52.740 ;
        RECT 73.770 52.680 74.060 52.725 ;
        RECT 71.410 52.540 74.060 52.680 ;
        RECT 71.410 52.480 71.730 52.540 ;
        RECT 73.770 52.495 74.060 52.540 ;
        RECT 62.210 52.340 62.530 52.400 ;
        RECT 51.260 52.200 62.530 52.340 ;
        RECT 16.210 52.140 16.530 52.200 ;
        RECT 24.045 52.155 24.335 52.200 ;
        RECT 62.210 52.140 62.530 52.200 ;
        RECT 78.310 52.140 78.630 52.400 ;
        RECT 84.305 52.340 84.595 52.385 ;
        RECT 86.605 52.340 86.895 52.385 ;
        RECT 84.305 52.200 86.895 52.340 ;
        RECT 84.305 52.155 84.595 52.200 ;
        RECT 86.605 52.155 86.895 52.200 ;
        RECT 13.380 51.520 92.040 52.000 ;
        RECT 28.170 51.320 28.490 51.380 ;
        RECT 33.230 51.320 33.550 51.380 ;
        RECT 28.170 51.180 33.550 51.320 ;
        RECT 28.170 51.120 28.490 51.180 ;
        RECT 33.230 51.120 33.550 51.180 ;
        RECT 33.690 51.320 34.010 51.380 ;
        RECT 35.990 51.320 36.310 51.380 ;
        RECT 33.690 51.180 36.310 51.320 ;
        RECT 33.690 51.120 34.010 51.180 ;
        RECT 35.990 51.120 36.310 51.180 ;
        RECT 58.530 51.120 58.850 51.380 ;
        RECT 60.385 51.320 60.675 51.365 ;
        RECT 60.830 51.320 61.150 51.380 ;
        RECT 60.385 51.180 61.150 51.320 ;
        RECT 60.385 51.135 60.675 51.180 ;
        RECT 60.830 51.120 61.150 51.180 ;
        RECT 61.290 51.320 61.610 51.380 ;
        RECT 77.850 51.320 78.170 51.380 ;
        RECT 61.290 51.180 78.170 51.320 ;
        RECT 61.290 51.120 61.610 51.180 ;
        RECT 77.850 51.120 78.170 51.180 ;
        RECT 24.505 50.980 24.795 51.025 ;
        RECT 26.790 50.980 27.110 51.040 ;
        RECT 24.505 50.840 27.110 50.980 ;
        RECT 24.505 50.795 24.795 50.840 ;
        RECT 26.790 50.780 27.110 50.840 ;
        RECT 31.405 50.980 31.695 51.025 ;
        RECT 39.670 50.980 39.990 51.040 ;
        RECT 52.550 51.025 52.870 51.040 ;
        RECT 52.520 50.980 52.870 51.025 ;
        RECT 31.405 50.840 39.990 50.980 ;
        RECT 52.355 50.840 52.870 50.980 ;
        RECT 31.405 50.795 31.695 50.840 ;
        RECT 39.670 50.780 39.990 50.840 ;
        RECT 52.520 50.795 52.870 50.840 ;
        RECT 52.550 50.780 52.870 50.795 ;
        RECT 77.390 50.980 77.710 51.040 ;
        RECT 78.785 50.980 79.075 51.025 ;
        RECT 77.390 50.840 79.075 50.980 ;
        RECT 77.390 50.780 77.710 50.840 ;
        RECT 78.785 50.795 79.075 50.840 ;
        RECT 16.210 50.440 16.530 50.700 ;
        RECT 18.065 50.640 18.355 50.685 ;
        RECT 20.350 50.640 20.670 50.700 ;
        RECT 18.065 50.500 20.670 50.640 ;
        RECT 18.065 50.455 18.355 50.500 ;
        RECT 20.350 50.440 20.670 50.500 ;
        RECT 25.425 50.455 25.715 50.685 ;
        RECT 26.880 50.640 27.020 50.780 ;
        RECT 31.865 50.640 32.155 50.685 ;
        RECT 26.880 50.500 32.155 50.640 ;
        RECT 31.865 50.455 32.155 50.500 ;
        RECT 32.785 50.640 33.075 50.685 ;
        RECT 34.610 50.640 34.930 50.700 ;
        RECT 32.785 50.500 34.930 50.640 ;
        RECT 32.785 50.455 33.075 50.500 ;
        RECT 12.990 49.960 13.310 50.020 ;
        RECT 17.145 49.960 17.435 50.005 ;
        RECT 25.500 49.960 25.640 50.455 ;
        RECT 34.610 50.440 34.930 50.500 ;
        RECT 38.305 50.455 38.595 50.685 ;
        RECT 27.725 50.300 28.015 50.345 ;
        RECT 28.630 50.300 28.950 50.360 ;
        RECT 30.930 50.300 31.250 50.360 ;
        RECT 27.725 50.160 31.250 50.300 ;
        RECT 27.725 50.115 28.015 50.160 ;
        RECT 28.630 50.100 28.950 50.160 ;
        RECT 30.930 50.100 31.250 50.160 ;
        RECT 31.390 50.300 31.710 50.360 ;
        RECT 33.705 50.300 33.995 50.345 ;
        RECT 31.390 50.160 33.995 50.300 ;
        RECT 38.380 50.300 38.520 50.455 ;
        RECT 41.050 50.440 41.370 50.700 ;
        RECT 41.510 50.440 41.830 50.700 ;
        RECT 42.430 50.440 42.750 50.700 ;
        RECT 42.905 50.640 43.195 50.685 ;
        RECT 44.270 50.640 44.590 50.700 ;
        RECT 45.190 50.685 45.510 50.700 ;
        RECT 42.905 50.500 44.590 50.640 ;
        RECT 42.905 50.455 43.195 50.500 ;
        RECT 44.270 50.440 44.590 50.500 ;
        RECT 45.160 50.455 45.510 50.685 ;
        RECT 51.185 50.640 51.475 50.685 ;
        RECT 53.930 50.640 54.250 50.700 ;
        RECT 51.185 50.500 54.250 50.640 ;
        RECT 51.185 50.455 51.475 50.500 ;
        RECT 45.190 50.440 45.510 50.455 ;
        RECT 53.930 50.440 54.250 50.500 ;
        RECT 78.310 50.440 78.630 50.700 ;
        RECT 90.270 50.440 90.590 50.700 ;
        RECT 38.380 50.160 42.660 50.300 ;
        RECT 31.390 50.100 31.710 50.160 ;
        RECT 33.705 50.115 33.995 50.160 ;
        RECT 42.520 50.020 42.660 50.160 ;
        RECT 43.825 50.115 44.115 50.345 ;
        RECT 44.705 50.300 44.995 50.345 ;
        RECT 45.895 50.300 46.185 50.345 ;
        RECT 48.415 50.300 48.705 50.345 ;
        RECT 44.705 50.160 48.705 50.300 ;
        RECT 44.705 50.115 44.995 50.160 ;
        RECT 45.895 50.115 46.185 50.160 ;
        RECT 48.415 50.115 48.705 50.160 ;
        RECT 52.065 50.300 52.355 50.345 ;
        RECT 53.255 50.300 53.545 50.345 ;
        RECT 55.775 50.300 56.065 50.345 ;
        RECT 52.065 50.160 56.065 50.300 ;
        RECT 52.065 50.115 52.355 50.160 ;
        RECT 53.255 50.115 53.545 50.160 ;
        RECT 55.775 50.115 56.065 50.160 ;
        RECT 41.510 49.960 41.830 50.020 ;
        RECT 12.990 49.820 17.435 49.960 ;
        RECT 12.990 49.760 13.310 49.820 ;
        RECT 17.145 49.775 17.435 49.820 ;
        RECT 21.590 49.820 41.830 49.960 ;
        RECT 14.370 49.620 14.690 49.680 ;
        RECT 15.305 49.620 15.595 49.665 ;
        RECT 14.370 49.480 15.595 49.620 ;
        RECT 14.370 49.420 14.690 49.480 ;
        RECT 15.305 49.435 15.595 49.480 ;
        RECT 16.210 49.620 16.530 49.680 ;
        RECT 21.590 49.620 21.730 49.820 ;
        RECT 41.510 49.760 41.830 49.820 ;
        RECT 42.430 49.960 42.750 50.020 ;
        RECT 43.900 49.960 44.040 50.115 ;
        RECT 60.830 50.100 61.150 50.360 ;
        RECT 61.305 50.115 61.595 50.345 ;
        RECT 42.430 49.820 44.040 49.960 ;
        RECT 44.310 49.960 44.600 50.005 ;
        RECT 46.410 49.960 46.700 50.005 ;
        RECT 47.980 49.960 48.270 50.005 ;
        RECT 44.310 49.820 48.270 49.960 ;
        RECT 42.430 49.760 42.750 49.820 ;
        RECT 44.310 49.775 44.600 49.820 ;
        RECT 46.410 49.775 46.700 49.820 ;
        RECT 47.980 49.775 48.270 49.820 ;
        RECT 50.710 49.760 51.030 50.020 ;
        RECT 51.670 49.960 51.960 50.005 ;
        RECT 53.770 49.960 54.060 50.005 ;
        RECT 55.340 49.960 55.630 50.005 ;
        RECT 51.670 49.820 55.630 49.960 ;
        RECT 51.670 49.775 51.960 49.820 ;
        RECT 53.770 49.775 54.060 49.820 ;
        RECT 55.340 49.775 55.630 49.820 ;
        RECT 58.085 49.960 58.375 50.005 ;
        RECT 58.990 49.960 59.310 50.020 ;
        RECT 58.085 49.820 59.310 49.960 ;
        RECT 58.085 49.775 58.375 49.820 ;
        RECT 58.990 49.760 59.310 49.820 ;
        RECT 16.210 49.480 21.730 49.620 ;
        RECT 26.345 49.620 26.635 49.665 ;
        RECT 28.170 49.620 28.490 49.680 ;
        RECT 26.345 49.480 28.490 49.620 ;
        RECT 16.210 49.420 16.530 49.480 ;
        RECT 26.345 49.435 26.635 49.480 ;
        RECT 28.170 49.420 28.490 49.480 ;
        RECT 40.145 49.620 40.435 49.665 ;
        RECT 47.490 49.620 47.810 49.680 ;
        RECT 40.145 49.480 47.810 49.620 ;
        RECT 40.145 49.435 40.435 49.480 ;
        RECT 47.490 49.420 47.810 49.480 ;
        RECT 49.330 49.620 49.650 49.680 ;
        RECT 55.770 49.620 56.090 49.680 ;
        RECT 61.380 49.620 61.520 50.115 ;
        RECT 88.890 49.960 89.210 50.020 ;
        RECT 89.365 49.960 89.655 50.005 ;
        RECT 88.890 49.820 89.655 49.960 ;
        RECT 88.890 49.760 89.210 49.820 ;
        RECT 89.365 49.775 89.655 49.820 ;
        RECT 49.330 49.480 61.520 49.620 ;
        RECT 49.330 49.420 49.650 49.480 ;
        RECT 55.770 49.420 56.090 49.480 ;
        RECT 13.380 48.800 92.040 49.280 ;
        RECT 30.010 48.600 30.330 48.660 ;
        RECT 37.370 48.600 37.690 48.660 ;
        RECT 30.010 48.460 37.690 48.600 ;
        RECT 30.010 48.400 30.330 48.460 ;
        RECT 37.370 48.400 37.690 48.460 ;
        RECT 37.845 48.600 38.135 48.645 ;
        RECT 41.510 48.600 41.830 48.660 ;
        RECT 37.845 48.460 41.830 48.600 ;
        RECT 37.845 48.415 38.135 48.460 ;
        RECT 41.510 48.400 41.830 48.460 ;
        RECT 45.190 48.600 45.510 48.660 ;
        RECT 45.665 48.600 45.955 48.645 ;
        RECT 45.190 48.460 45.955 48.600 ;
        RECT 45.190 48.400 45.510 48.460 ;
        RECT 45.665 48.415 45.955 48.460 ;
        RECT 53.010 48.600 53.330 48.660 ;
        RECT 57.165 48.600 57.455 48.645 ;
        RECT 53.010 48.460 57.455 48.600 ;
        RECT 53.010 48.400 53.330 48.460 ;
        RECT 57.165 48.415 57.455 48.460 ;
        RECT 62.210 48.400 62.530 48.660 ;
        RECT 63.130 48.600 63.450 48.660 ;
        RECT 71.870 48.600 72.190 48.660 ;
        RECT 63.130 48.460 72.190 48.600 ;
        RECT 63.130 48.400 63.450 48.460 ;
        RECT 71.870 48.400 72.190 48.460 ;
        RECT 12.070 48.260 12.390 48.320 ;
        RECT 15.305 48.260 15.595 48.305 ;
        RECT 21.730 48.260 22.050 48.320 ;
        RECT 25.410 48.260 25.730 48.320 ;
        RECT 12.070 48.120 15.595 48.260 ;
        RECT 12.070 48.060 12.390 48.120 ;
        RECT 15.305 48.075 15.595 48.120 ;
        RECT 17.680 48.120 25.730 48.260 ;
        RECT 16.210 47.380 16.530 47.640 ;
        RECT 17.680 47.625 17.820 48.120 ;
        RECT 21.730 48.060 22.050 48.120 ;
        RECT 25.410 48.060 25.730 48.120 ;
        RECT 31.430 48.260 31.720 48.305 ;
        RECT 33.530 48.260 33.820 48.305 ;
        RECT 35.100 48.260 35.390 48.305 ;
        RECT 31.430 48.120 35.390 48.260 ;
        RECT 31.430 48.075 31.720 48.120 ;
        RECT 33.530 48.075 33.820 48.120 ;
        RECT 35.100 48.075 35.390 48.120 ;
        RECT 38.790 48.260 39.080 48.305 ;
        RECT 40.890 48.260 41.180 48.305 ;
        RECT 42.460 48.260 42.750 48.305 ;
        RECT 38.790 48.120 42.750 48.260 ;
        RECT 38.790 48.075 39.080 48.120 ;
        RECT 40.890 48.075 41.180 48.120 ;
        RECT 42.460 48.075 42.750 48.120 ;
        RECT 44.270 48.260 44.590 48.320 ;
        RECT 72.805 48.260 73.095 48.305 ;
        RECT 44.270 48.120 73.095 48.260 ;
        RECT 44.270 48.060 44.590 48.120 ;
        RECT 72.805 48.075 73.095 48.120 ;
        RECT 20.810 47.920 21.130 47.980 ;
        RECT 29.550 47.920 29.870 47.980 ;
        RECT 19.060 47.780 29.870 47.920 ;
        RECT 17.605 47.395 17.895 47.625 ;
        RECT 18.050 47.580 18.370 47.640 ;
        RECT 19.060 47.625 19.200 47.780 ;
        RECT 20.810 47.720 21.130 47.780 ;
        RECT 18.525 47.580 18.815 47.625 ;
        RECT 18.050 47.440 18.815 47.580 ;
        RECT 18.050 47.380 18.370 47.440 ;
        RECT 18.525 47.395 18.815 47.440 ;
        RECT 18.985 47.395 19.275 47.625 ;
        RECT 19.430 47.380 19.750 47.640 ;
        RECT 22.650 47.380 22.970 47.640 ;
        RECT 26.330 47.580 26.650 47.640 ;
        RECT 27.265 47.580 27.555 47.625 ;
        RECT 26.330 47.440 27.555 47.580 ;
        RECT 26.330 47.380 26.650 47.440 ;
        RECT 27.265 47.395 27.555 47.440 ;
        RECT 20.810 46.700 21.130 46.960 ;
        RECT 21.730 46.700 22.050 46.960 ;
        RECT 27.340 46.900 27.480 47.395 ;
        RECT 28.170 47.380 28.490 47.640 ;
        RECT 28.720 47.625 28.860 47.780 ;
        RECT 29.550 47.720 29.870 47.780 ;
        RECT 30.930 47.720 31.250 47.980 ;
        RECT 31.825 47.920 32.115 47.965 ;
        RECT 33.015 47.920 33.305 47.965 ;
        RECT 35.535 47.920 35.825 47.965 ;
        RECT 31.825 47.780 35.825 47.920 ;
        RECT 31.825 47.735 32.115 47.780 ;
        RECT 33.015 47.735 33.305 47.780 ;
        RECT 35.535 47.735 35.825 47.780 ;
        RECT 39.185 47.920 39.475 47.965 ;
        RECT 40.375 47.920 40.665 47.965 ;
        RECT 42.895 47.920 43.185 47.965 ;
        RECT 39.185 47.780 43.185 47.920 ;
        RECT 39.185 47.735 39.475 47.780 ;
        RECT 40.375 47.735 40.665 47.780 ;
        RECT 42.895 47.735 43.185 47.780 ;
        RECT 47.490 47.920 47.810 47.980 ;
        RECT 47.965 47.920 48.255 47.965 ;
        RECT 47.490 47.780 48.255 47.920 ;
        RECT 47.490 47.720 47.810 47.780 ;
        RECT 47.965 47.735 48.255 47.780 ;
        RECT 48.885 47.920 49.175 47.965 ;
        RECT 49.330 47.920 49.650 47.980 ;
        RECT 48.885 47.780 49.650 47.920 ;
        RECT 48.885 47.735 49.175 47.780 ;
        RECT 49.330 47.720 49.650 47.780 ;
        RECT 50.710 47.920 51.030 47.980 ;
        RECT 55.325 47.920 55.615 47.965 ;
        RECT 50.710 47.780 55.615 47.920 ;
        RECT 50.710 47.720 51.030 47.780 ;
        RECT 55.325 47.735 55.615 47.780 ;
        RECT 55.770 47.920 56.090 47.980 ;
        RECT 74.170 47.920 74.490 47.980 ;
        RECT 55.770 47.780 58.300 47.920 ;
        RECT 55.770 47.720 56.090 47.780 ;
        RECT 28.645 47.395 28.935 47.625 ;
        RECT 29.105 47.580 29.395 47.625 ;
        RECT 31.390 47.580 31.710 47.640 ;
        RECT 35.070 47.580 35.390 47.640 ;
        RECT 29.105 47.440 35.390 47.580 ;
        RECT 29.105 47.395 29.395 47.440 ;
        RECT 31.390 47.380 31.710 47.440 ;
        RECT 35.070 47.380 35.390 47.440 ;
        RECT 38.305 47.580 38.595 47.625 ;
        RECT 42.430 47.580 42.750 47.640 ;
        RECT 38.305 47.440 42.750 47.580 ;
        RECT 38.305 47.395 38.595 47.440 ;
        RECT 42.430 47.380 42.750 47.440 ;
        RECT 42.980 47.440 57.840 47.580 ;
        RECT 30.485 47.240 30.775 47.285 ;
        RECT 32.170 47.240 32.460 47.285 ;
        RECT 30.485 47.100 32.460 47.240 ;
        RECT 30.485 47.055 30.775 47.100 ;
        RECT 32.170 47.055 32.460 47.100 ;
        RECT 33.230 47.240 33.550 47.300 ;
        RECT 34.610 47.240 34.930 47.300 ;
        RECT 33.230 47.100 34.930 47.240 ;
        RECT 33.230 47.040 33.550 47.100 ;
        RECT 34.610 47.040 34.930 47.100 ;
        RECT 39.640 47.240 39.930 47.285 ;
        RECT 40.130 47.240 40.450 47.300 ;
        RECT 42.980 47.240 43.120 47.440 ;
        RECT 39.640 47.100 40.450 47.240 ;
        RECT 39.640 47.055 39.930 47.100 ;
        RECT 40.130 47.040 40.450 47.100 ;
        RECT 40.680 47.100 43.120 47.240 ;
        RECT 47.505 47.240 47.795 47.285 ;
        RECT 52.565 47.240 52.855 47.285 ;
        RECT 47.505 47.100 52.855 47.240 ;
        RECT 40.680 46.900 40.820 47.100 ;
        RECT 47.505 47.055 47.795 47.100 ;
        RECT 52.565 47.055 52.855 47.100 ;
        RECT 56.230 47.040 56.550 47.300 ;
        RECT 27.340 46.760 40.820 46.900 ;
        RECT 41.050 46.900 41.370 46.960 ;
        RECT 45.190 46.900 45.510 46.960 ;
        RECT 41.050 46.760 45.510 46.900 ;
        RECT 41.050 46.700 41.370 46.760 ;
        RECT 45.190 46.700 45.510 46.760 ;
        RECT 57.150 46.700 57.470 46.960 ;
        RECT 57.700 46.900 57.840 47.440 ;
        RECT 58.160 47.240 58.300 47.780 ;
        RECT 63.680 47.780 74.490 47.920 ;
        RECT 58.545 47.580 58.835 47.625 ;
        RECT 63.130 47.580 63.450 47.640 ;
        RECT 63.680 47.625 63.820 47.780 ;
        RECT 74.170 47.720 74.490 47.780 ;
        RECT 58.545 47.440 63.450 47.580 ;
        RECT 58.545 47.395 58.835 47.440 ;
        RECT 63.130 47.380 63.450 47.440 ;
        RECT 63.605 47.395 63.895 47.625 ;
        RECT 64.970 47.380 65.290 47.640 ;
        RECT 65.445 47.580 65.735 47.625 ;
        RECT 66.825 47.580 67.115 47.625 ;
        RECT 68.650 47.580 68.970 47.640 ;
        RECT 65.445 47.440 66.120 47.580 ;
        RECT 65.445 47.395 65.735 47.440 ;
        RECT 59.465 47.240 59.755 47.285 ;
        RECT 58.160 47.100 59.755 47.240 ;
        RECT 59.465 47.055 59.755 47.100 ;
        RECT 60.385 47.240 60.675 47.285 ;
        RECT 62.670 47.240 62.990 47.300 ;
        RECT 64.065 47.240 64.355 47.285 ;
        RECT 60.385 47.100 64.355 47.240 ;
        RECT 60.385 47.055 60.675 47.100 ;
        RECT 62.670 47.040 62.990 47.100 ;
        RECT 64.065 47.055 64.355 47.100 ;
        RECT 65.980 46.900 66.120 47.440 ;
        RECT 66.825 47.440 68.970 47.580 ;
        RECT 66.825 47.395 67.115 47.440 ;
        RECT 68.650 47.380 68.970 47.440 ;
        RECT 70.045 47.580 70.335 47.625 ;
        RECT 70.490 47.580 70.810 47.640 ;
        RECT 70.045 47.440 70.810 47.580 ;
        RECT 70.045 47.395 70.335 47.440 ;
        RECT 70.490 47.380 70.810 47.440 ;
        RECT 71.870 47.380 72.190 47.640 ;
        RECT 78.325 47.580 78.615 47.625 ;
        RECT 73.340 47.440 78.615 47.580 ;
        RECT 66.350 47.240 66.670 47.300 ;
        RECT 70.965 47.240 71.255 47.285 ;
        RECT 66.350 47.100 71.255 47.240 ;
        RECT 66.350 47.040 66.670 47.100 ;
        RECT 70.965 47.055 71.255 47.100 ;
        RECT 71.425 47.240 71.715 47.285 ;
        RECT 72.330 47.240 72.650 47.300 ;
        RECT 73.340 47.240 73.480 47.440 ;
        RECT 78.325 47.395 78.615 47.440 ;
        RECT 71.425 47.100 72.650 47.240 ;
        RECT 71.425 47.055 71.715 47.100 ;
        RECT 72.330 47.040 72.650 47.100 ;
        RECT 72.880 47.100 73.480 47.240 ;
        RECT 57.700 46.760 66.120 46.900 ;
        RECT 68.650 46.900 68.970 46.960 ;
        RECT 72.880 46.900 73.020 47.100 ;
        RECT 74.170 47.040 74.490 47.300 ;
        RECT 75.090 47.040 75.410 47.300 ;
        RECT 78.400 47.240 78.540 47.395 ;
        RECT 79.230 47.380 79.550 47.640 ;
        RECT 79.690 47.380 80.010 47.640 ;
        RECT 80.150 47.380 80.470 47.640 ;
        RECT 84.750 47.240 85.070 47.300 ;
        RECT 78.400 47.100 85.070 47.240 ;
        RECT 84.750 47.040 85.070 47.100 ;
        RECT 68.650 46.760 73.020 46.900 ;
        RECT 68.650 46.700 68.970 46.760 ;
        RECT 73.250 46.700 73.570 46.960 ;
        RECT 81.530 46.700 81.850 46.960 ;
        RECT 13.380 46.080 92.040 46.560 ;
        RECT 18.050 45.680 18.370 45.940 ;
        RECT 23.570 45.880 23.890 45.940 ;
        RECT 25.425 45.880 25.715 45.925 ;
        RECT 38.750 45.880 39.070 45.940 ;
        RECT 19.520 45.740 25.715 45.880 ;
        RECT 14.830 45.540 15.150 45.600 ;
        RECT 16.225 45.540 16.515 45.585 ;
        RECT 14.830 45.400 16.515 45.540 ;
        RECT 14.830 45.340 15.150 45.400 ;
        RECT 16.225 45.355 16.515 45.400 ;
        RECT 17.145 45.540 17.435 45.585 ;
        RECT 19.520 45.540 19.660 45.740 ;
        RECT 23.570 45.680 23.890 45.740 ;
        RECT 25.425 45.695 25.715 45.740 ;
        RECT 27.340 45.740 39.070 45.880 ;
        RECT 17.145 45.400 19.660 45.540 ;
        RECT 19.860 45.540 20.150 45.585 ;
        RECT 20.810 45.540 21.130 45.600 ;
        RECT 19.860 45.400 21.130 45.540 ;
        RECT 17.145 45.355 17.435 45.400 ;
        RECT 19.860 45.355 20.150 45.400 ;
        RECT 16.300 45.200 16.440 45.355 ;
        RECT 20.810 45.340 21.130 45.400 ;
        RECT 22.650 45.540 22.970 45.600 ;
        RECT 26.845 45.540 27.135 45.585 ;
        RECT 27.340 45.540 27.480 45.740 ;
        RECT 38.750 45.680 39.070 45.740 ;
        RECT 74.170 45.880 74.490 45.940 ;
        RECT 81.085 45.880 81.375 45.925 ;
        RECT 83.830 45.880 84.150 45.940 ;
        RECT 74.170 45.740 84.150 45.880 ;
        RECT 74.170 45.680 74.490 45.740 ;
        RECT 81.085 45.695 81.375 45.740 ;
        RECT 83.830 45.680 84.150 45.740 ;
        RECT 22.650 45.400 27.480 45.540 ;
        RECT 27.725 45.540 28.015 45.585 ;
        RECT 27.725 45.400 29.320 45.540 ;
        RECT 22.650 45.340 22.970 45.400 ;
        RECT 26.845 45.355 27.135 45.400 ;
        RECT 27.725 45.355 28.015 45.400 ;
        RECT 25.885 45.200 26.175 45.245 ;
        RECT 27.250 45.200 27.570 45.260 ;
        RECT 29.180 45.245 29.320 45.400 ;
        RECT 31.940 45.400 33.920 45.540 ;
        RECT 16.300 45.060 27.570 45.200 ;
        RECT 25.885 45.015 26.175 45.060 ;
        RECT 27.250 45.000 27.570 45.060 ;
        RECT 28.185 45.015 28.475 45.245 ;
        RECT 29.105 45.015 29.395 45.245 ;
        RECT 16.670 44.860 16.990 44.920 ;
        RECT 18.525 44.860 18.815 44.905 ;
        RECT 16.670 44.720 18.815 44.860 ;
        RECT 16.670 44.660 16.990 44.720 ;
        RECT 18.525 44.675 18.815 44.720 ;
        RECT 19.405 44.860 19.695 44.905 ;
        RECT 20.595 44.860 20.885 44.905 ;
        RECT 23.115 44.860 23.405 44.905 ;
        RECT 19.405 44.720 23.405 44.860 ;
        RECT 19.405 44.675 19.695 44.720 ;
        RECT 20.595 44.675 20.885 44.720 ;
        RECT 23.115 44.675 23.405 44.720 ;
        RECT 25.410 44.860 25.730 44.920 ;
        RECT 26.790 44.860 27.110 44.920 ;
        RECT 28.260 44.860 28.400 45.015 ;
        RECT 29.550 45.000 29.870 45.260 ;
        RECT 30.010 45.000 30.330 45.260 ;
        RECT 31.940 45.245 32.080 45.400 ;
        RECT 31.865 45.015 32.155 45.245 ;
        RECT 33.145 45.200 33.435 45.245 ;
        RECT 32.400 45.060 33.435 45.200 ;
        RECT 33.780 45.200 33.920 45.400 ;
        RECT 39.670 45.340 39.990 45.600 ;
        RECT 41.510 45.540 41.830 45.600 ;
        RECT 44.745 45.540 45.035 45.585 ;
        RECT 54.405 45.540 54.695 45.585 ;
        RECT 55.770 45.540 56.090 45.600 ;
        RECT 41.510 45.400 45.035 45.540 ;
        RECT 41.510 45.340 41.830 45.400 ;
        RECT 44.745 45.355 45.035 45.400 ;
        RECT 49.420 45.400 56.090 45.540 ;
        RECT 42.430 45.200 42.750 45.260 ;
        RECT 45.190 45.200 45.510 45.260 ;
        RECT 47.505 45.200 47.795 45.245 ;
        RECT 48.885 45.200 49.175 45.245 ;
        RECT 33.780 45.060 43.580 45.200 ;
        RECT 25.410 44.720 28.400 44.860 ;
        RECT 29.640 44.860 29.780 45.000 ;
        RECT 30.930 44.860 31.250 44.920 ;
        RECT 29.640 44.720 31.250 44.860 ;
        RECT 25.410 44.660 25.730 44.720 ;
        RECT 26.790 44.660 27.110 44.720 ;
        RECT 30.930 44.660 31.250 44.720 ;
        RECT 31.405 44.860 31.695 44.905 ;
        RECT 32.400 44.860 32.540 45.060 ;
        RECT 33.145 45.015 33.435 45.060 ;
        RECT 42.430 45.000 42.750 45.060 ;
        RECT 43.440 44.905 43.580 45.060 ;
        RECT 45.190 45.060 49.175 45.200 ;
        RECT 45.190 45.000 45.510 45.060 ;
        RECT 47.505 45.015 47.795 45.060 ;
        RECT 48.885 45.015 49.175 45.060 ;
        RECT 31.405 44.720 32.540 44.860 ;
        RECT 32.745 44.860 33.035 44.905 ;
        RECT 33.935 44.860 34.225 44.905 ;
        RECT 36.455 44.860 36.745 44.905 ;
        RECT 32.745 44.720 36.745 44.860 ;
        RECT 31.405 44.675 31.695 44.720 ;
        RECT 32.745 44.675 33.035 44.720 ;
        RECT 33.935 44.675 34.225 44.720 ;
        RECT 36.455 44.675 36.745 44.720 ;
        RECT 43.365 44.860 43.655 44.905 ;
        RECT 44.730 44.860 45.050 44.920 ;
        RECT 43.365 44.720 45.050 44.860 ;
        RECT 43.365 44.675 43.655 44.720 ;
        RECT 44.730 44.660 45.050 44.720 ;
        RECT 19.010 44.520 19.300 44.565 ;
        RECT 21.110 44.520 21.400 44.565 ;
        RECT 22.680 44.520 22.970 44.565 ;
        RECT 19.010 44.380 22.970 44.520 ;
        RECT 19.010 44.335 19.300 44.380 ;
        RECT 21.110 44.335 21.400 44.380 ;
        RECT 22.680 44.335 22.970 44.380 ;
        RECT 32.350 44.520 32.640 44.565 ;
        RECT 34.450 44.520 34.740 44.565 ;
        RECT 36.020 44.520 36.310 44.565 ;
        RECT 32.350 44.380 36.310 44.520 ;
        RECT 32.350 44.335 32.640 44.380 ;
        RECT 34.450 44.335 34.740 44.380 ;
        RECT 36.020 44.335 36.310 44.380 ;
        RECT 38.750 44.320 39.070 44.580 ;
        RECT 23.110 44.180 23.430 44.240 ;
        RECT 49.420 44.180 49.560 45.400 ;
        RECT 54.405 45.355 54.695 45.400 ;
        RECT 55.770 45.340 56.090 45.400 ;
        RECT 67.270 45.540 67.590 45.600 ;
        RECT 73.265 45.540 73.555 45.585 ;
        RECT 78.310 45.540 78.630 45.600 ;
        RECT 67.270 45.400 69.340 45.540 ;
        RECT 67.270 45.340 67.590 45.400 ;
        RECT 69.200 45.260 69.340 45.400 ;
        RECT 73.265 45.400 78.630 45.540 ;
        RECT 73.265 45.355 73.555 45.400 ;
        RECT 49.790 45.200 50.110 45.260 ;
        RECT 50.725 45.200 51.015 45.245 ;
        RECT 51.645 45.200 51.935 45.245 ;
        RECT 52.090 45.200 52.410 45.260 ;
        RECT 49.790 45.060 52.410 45.200 ;
        RECT 49.790 45.000 50.110 45.060 ;
        RECT 50.725 45.015 51.015 45.060 ;
        RECT 51.645 45.015 51.935 45.060 ;
        RECT 52.090 45.000 52.410 45.060 ;
        RECT 53.010 45.000 53.330 45.260 ;
        RECT 53.930 45.200 54.250 45.260 ;
        RECT 56.690 45.200 57.010 45.260 ;
        RECT 53.930 45.060 57.010 45.200 ;
        RECT 53.930 45.000 54.250 45.060 ;
        RECT 56.690 45.000 57.010 45.060 ;
        RECT 61.290 45.000 61.610 45.260 ;
        RECT 62.225 45.200 62.515 45.245 ;
        RECT 62.670 45.200 62.990 45.260 ;
        RECT 66.350 45.200 66.670 45.260 ;
        RECT 62.225 45.060 66.670 45.200 ;
        RECT 62.225 45.015 62.515 45.060 ;
        RECT 62.670 45.000 62.990 45.060 ;
        RECT 66.350 45.000 66.670 45.060 ;
        RECT 68.665 45.015 68.955 45.245 ;
        RECT 53.485 44.675 53.775 44.905 ;
        RECT 53.560 44.520 53.700 44.675 ;
        RECT 60.370 44.660 60.690 44.920 ;
        RECT 67.270 44.860 67.590 44.920 ;
        RECT 68.740 44.860 68.880 45.015 ;
        RECT 69.110 45.000 69.430 45.260 ;
        RECT 73.340 44.860 73.480 45.355 ;
        RECT 78.310 45.340 78.630 45.400 ;
        RECT 73.710 45.200 74.030 45.260 ;
        RECT 75.465 45.200 75.755 45.245 ;
        RECT 73.710 45.060 75.755 45.200 ;
        RECT 73.710 45.000 74.030 45.060 ;
        RECT 75.465 45.015 75.755 45.060 ;
        RECT 88.890 45.000 89.210 45.260 ;
        RECT 74.185 44.860 74.475 44.905 ;
        RECT 67.270 44.720 74.475 44.860 ;
        RECT 67.270 44.660 67.590 44.720 ;
        RECT 74.185 44.675 74.475 44.720 ;
        RECT 75.065 44.860 75.355 44.905 ;
        RECT 76.255 44.860 76.545 44.905 ;
        RECT 78.775 44.860 79.065 44.905 ;
        RECT 75.065 44.720 79.065 44.860 ;
        RECT 75.065 44.675 75.355 44.720 ;
        RECT 76.255 44.675 76.545 44.720 ;
        RECT 78.775 44.675 79.065 44.720 ;
        RECT 57.150 44.520 57.470 44.580 ;
        RECT 53.560 44.380 57.470 44.520 ;
        RECT 57.150 44.320 57.470 44.380 ;
        RECT 74.670 44.520 74.960 44.565 ;
        RECT 76.770 44.520 77.060 44.565 ;
        RECT 78.340 44.520 78.630 44.565 ;
        RECT 74.670 44.380 78.630 44.520 ;
        RECT 74.670 44.335 74.960 44.380 ;
        RECT 76.770 44.335 77.060 44.380 ;
        RECT 78.340 44.335 78.630 44.380 ;
        RECT 89.825 44.520 90.115 44.565 ;
        RECT 90.730 44.520 91.050 44.580 ;
        RECT 89.825 44.380 91.050 44.520 ;
        RECT 89.825 44.335 90.115 44.380 ;
        RECT 90.730 44.320 91.050 44.380 ;
        RECT 23.110 44.040 49.560 44.180 ;
        RECT 23.110 43.980 23.430 44.040 ;
        RECT 13.380 43.360 92.040 43.840 ;
        RECT 16.670 43.160 16.990 43.220 ;
        RECT 14.920 43.020 16.990 43.160 ;
        RECT 14.920 42.525 15.060 43.020 ;
        RECT 16.670 42.960 16.990 43.020 ;
        RECT 20.350 43.160 20.670 43.220 ;
        RECT 21.745 43.160 22.035 43.205 ;
        RECT 20.350 43.020 22.035 43.160 ;
        RECT 20.350 42.960 20.670 43.020 ;
        RECT 21.745 42.975 22.035 43.020 ;
        RECT 30.485 43.160 30.775 43.205 ;
        RECT 30.930 43.160 31.250 43.220 ;
        RECT 30.485 43.020 31.250 43.160 ;
        RECT 30.485 42.975 30.775 43.020 ;
        RECT 30.930 42.960 31.250 43.020 ;
        RECT 39.685 43.160 39.975 43.205 ;
        RECT 40.130 43.160 40.450 43.220 ;
        RECT 51.645 43.160 51.935 43.205 ;
        RECT 53.010 43.160 53.330 43.220 ;
        RECT 61.290 43.160 61.610 43.220 ;
        RECT 72.330 43.160 72.650 43.220 ;
        RECT 39.685 43.020 40.450 43.160 ;
        RECT 39.685 42.975 39.975 43.020 ;
        RECT 40.130 42.960 40.450 43.020 ;
        RECT 40.680 43.020 49.560 43.160 ;
        RECT 15.330 42.820 15.620 42.865 ;
        RECT 17.430 42.820 17.720 42.865 ;
        RECT 19.000 42.820 19.290 42.865 ;
        RECT 15.330 42.680 19.290 42.820 ;
        RECT 15.330 42.635 15.620 42.680 ;
        RECT 17.430 42.635 17.720 42.680 ;
        RECT 19.000 42.635 19.290 42.680 ;
        RECT 25.870 42.820 26.190 42.880 ;
        RECT 29.565 42.820 29.855 42.865 ;
        RECT 38.290 42.820 38.610 42.880 ;
        RECT 25.870 42.680 28.860 42.820 ;
        RECT 25.870 42.620 26.190 42.680 ;
        RECT 14.845 42.295 15.135 42.525 ;
        RECT 15.725 42.480 16.015 42.525 ;
        RECT 16.915 42.480 17.205 42.525 ;
        RECT 19.435 42.480 19.725 42.525 ;
        RECT 28.720 42.480 28.860 42.680 ;
        RECT 29.565 42.680 38.610 42.820 ;
        RECT 29.565 42.635 29.855 42.680 ;
        RECT 38.290 42.620 38.610 42.680 ;
        RECT 30.470 42.480 30.790 42.540 ;
        RECT 15.725 42.340 19.725 42.480 ;
        RECT 15.725 42.295 16.015 42.340 ;
        RECT 16.915 42.295 17.205 42.340 ;
        RECT 19.435 42.295 19.725 42.340 ;
        RECT 23.660 42.340 28.400 42.480 ;
        RECT 23.660 42.200 23.800 42.340 ;
        RECT 23.570 41.940 23.890 42.200 ;
        RECT 24.950 42.140 25.270 42.200 ;
        RECT 26.805 42.140 27.095 42.185 ;
        RECT 24.950 42.000 27.095 42.140 ;
        RECT 24.950 41.940 25.270 42.000 ;
        RECT 26.805 41.955 27.095 42.000 ;
        RECT 27.265 42.140 27.555 42.185 ;
        RECT 27.710 42.140 28.030 42.200 ;
        RECT 28.260 42.185 28.400 42.340 ;
        RECT 28.720 42.340 30.790 42.480 ;
        RECT 28.720 42.185 28.860 42.340 ;
        RECT 30.470 42.280 30.790 42.340 ;
        RECT 32.785 42.480 33.075 42.525 ;
        RECT 34.610 42.480 34.930 42.540 ;
        RECT 40.680 42.480 40.820 43.020 ;
        RECT 45.230 42.820 45.520 42.865 ;
        RECT 47.330 42.820 47.620 42.865 ;
        RECT 48.900 42.820 49.190 42.865 ;
        RECT 45.230 42.680 49.190 42.820 ;
        RECT 49.420 42.820 49.560 43.020 ;
        RECT 51.645 43.020 53.330 43.160 ;
        RECT 51.645 42.975 51.935 43.020 ;
        RECT 53.010 42.960 53.330 43.020 ;
        RECT 53.560 43.020 72.650 43.160 ;
        RECT 53.560 42.820 53.700 43.020 ;
        RECT 61.290 42.960 61.610 43.020 ;
        RECT 72.330 42.960 72.650 43.020 ;
        RECT 73.710 42.960 74.030 43.220 ;
        RECT 76.025 43.160 76.315 43.205 ;
        RECT 79.230 43.160 79.550 43.220 ;
        RECT 76.025 43.020 79.550 43.160 ;
        RECT 76.025 42.975 76.315 43.020 ;
        RECT 79.230 42.960 79.550 43.020 ;
        RECT 49.420 42.680 53.700 42.820 ;
        RECT 54.430 42.820 54.720 42.865 ;
        RECT 56.530 42.820 56.820 42.865 ;
        RECT 58.100 42.820 58.390 42.865 ;
        RECT 54.430 42.680 58.390 42.820 ;
        RECT 45.230 42.635 45.520 42.680 ;
        RECT 47.330 42.635 47.620 42.680 ;
        RECT 48.900 42.635 49.190 42.680 ;
        RECT 54.430 42.635 54.720 42.680 ;
        RECT 56.530 42.635 56.820 42.680 ;
        RECT 58.100 42.635 58.390 42.680 ;
        RECT 62.710 42.820 63.000 42.865 ;
        RECT 64.810 42.820 65.100 42.865 ;
        RECT 66.380 42.820 66.670 42.865 ;
        RECT 62.710 42.680 66.670 42.820 ;
        RECT 62.710 42.635 63.000 42.680 ;
        RECT 64.810 42.635 65.100 42.680 ;
        RECT 66.380 42.635 66.670 42.680 ;
        RECT 78.810 42.820 79.100 42.865 ;
        RECT 80.910 42.820 81.200 42.865 ;
        RECT 82.480 42.820 82.770 42.865 ;
        RECT 78.810 42.680 82.770 42.820 ;
        RECT 78.810 42.635 79.100 42.680 ;
        RECT 80.910 42.635 81.200 42.680 ;
        RECT 82.480 42.635 82.770 42.680 ;
        RECT 41.985 42.480 42.275 42.525 ;
        RECT 32.785 42.340 40.820 42.480 ;
        RECT 41.140 42.340 42.275 42.480 ;
        RECT 32.785 42.295 33.075 42.340 ;
        RECT 34.610 42.280 34.930 42.340 ;
        RECT 27.265 42.000 28.030 42.140 ;
        RECT 27.265 41.955 27.555 42.000 ;
        RECT 27.710 41.940 28.030 42.000 ;
        RECT 28.185 41.955 28.475 42.185 ;
        RECT 28.645 41.955 28.935 42.185 ;
        RECT 29.090 42.140 29.410 42.200 ;
        RECT 31.865 42.140 32.155 42.185 ;
        RECT 32.325 42.140 32.615 42.185 ;
        RECT 34.150 42.140 34.470 42.200 ;
        RECT 29.090 42.000 34.470 42.140 ;
        RECT 29.090 41.940 29.410 42.000 ;
        RECT 31.865 41.955 32.155 42.000 ;
        RECT 32.325 41.955 32.615 42.000 ;
        RECT 34.150 41.940 34.470 42.000 ;
        RECT 37.830 42.140 38.150 42.200 ;
        RECT 41.140 42.140 41.280 42.340 ;
        RECT 41.985 42.295 42.275 42.340 ;
        RECT 42.905 42.480 43.195 42.525 ;
        RECT 45.625 42.480 45.915 42.525 ;
        RECT 46.815 42.480 47.105 42.525 ;
        RECT 49.335 42.480 49.625 42.525 ;
        RECT 42.905 42.340 45.420 42.480 ;
        RECT 42.905 42.295 43.195 42.340 ;
        RECT 37.830 42.000 41.280 42.140 ;
        RECT 37.830 41.940 38.150 42.000 ;
        RECT 41.510 41.940 41.830 42.200 ;
        RECT 44.730 41.940 45.050 42.200 ;
        RECT 45.280 42.140 45.420 42.340 ;
        RECT 45.625 42.340 49.625 42.480 ;
        RECT 45.625 42.295 45.915 42.340 ;
        RECT 46.815 42.295 47.105 42.340 ;
        RECT 49.335 42.295 49.625 42.340 ;
        RECT 54.825 42.480 55.115 42.525 ;
        RECT 56.015 42.480 56.305 42.525 ;
        RECT 58.535 42.480 58.825 42.525 ;
        RECT 54.825 42.340 58.825 42.480 ;
        RECT 54.825 42.295 55.115 42.340 ;
        RECT 56.015 42.295 56.305 42.340 ;
        RECT 58.535 42.295 58.825 42.340 ;
        RECT 63.105 42.480 63.395 42.525 ;
        RECT 64.295 42.480 64.585 42.525 ;
        RECT 66.815 42.480 67.105 42.525 ;
        RECT 73.250 42.480 73.570 42.540 ;
        RECT 63.105 42.340 67.105 42.480 ;
        RECT 63.105 42.295 63.395 42.340 ;
        RECT 64.295 42.295 64.585 42.340 ;
        RECT 66.815 42.295 67.105 42.340 ;
        RECT 71.500 42.340 73.570 42.480 ;
        RECT 52.090 42.140 52.410 42.200 ;
        RECT 52.565 42.140 52.855 42.185 ;
        RECT 45.280 42.000 49.560 42.140 ;
        RECT 49.420 41.860 49.560 42.000 ;
        RECT 52.090 42.000 52.855 42.140 ;
        RECT 52.090 41.940 52.410 42.000 ;
        RECT 52.565 41.955 52.855 42.000 ;
        RECT 53.945 42.140 54.235 42.185 ;
        RECT 56.690 42.140 57.010 42.200 ;
        RECT 62.225 42.140 62.515 42.185 ;
        RECT 67.270 42.140 67.590 42.200 ;
        RECT 53.945 42.000 58.760 42.140 ;
        RECT 53.945 41.955 54.235 42.000 ;
        RECT 56.690 41.940 57.010 42.000 ;
        RECT 58.620 41.860 58.760 42.000 ;
        RECT 62.225 42.000 67.590 42.140 ;
        RECT 62.225 41.955 62.515 42.000 ;
        RECT 67.270 41.940 67.590 42.000 ;
        RECT 68.650 42.140 68.970 42.200 ;
        RECT 71.500 42.185 71.640 42.340 ;
        RECT 73.250 42.280 73.570 42.340 ;
        RECT 79.205 42.480 79.495 42.525 ;
        RECT 80.395 42.480 80.685 42.525 ;
        RECT 82.915 42.480 83.205 42.525 ;
        RECT 79.205 42.340 83.205 42.480 ;
        RECT 79.205 42.295 79.495 42.340 ;
        RECT 80.395 42.295 80.685 42.340 ;
        RECT 82.915 42.295 83.205 42.340 ;
        RECT 70.505 42.140 70.795 42.185 ;
        RECT 68.650 42.000 70.795 42.140 ;
        RECT 68.650 41.940 68.970 42.000 ;
        RECT 70.505 41.955 70.795 42.000 ;
        RECT 71.425 41.955 71.715 42.185 ;
        RECT 71.870 41.940 72.190 42.200 ;
        RECT 72.345 41.955 72.635 42.185 ;
        RECT 72.790 42.140 73.110 42.200 ;
        RECT 75.105 42.140 75.395 42.185 ;
        RECT 72.790 42.000 75.395 42.140 ;
        RECT 16.210 41.845 16.530 41.860 ;
        RECT 16.180 41.615 16.530 41.845 ;
        RECT 16.210 41.600 16.530 41.615 ;
        RECT 30.930 41.800 31.250 41.860 ;
        RECT 46.080 41.800 46.370 41.845 ;
        RECT 47.950 41.800 48.270 41.860 ;
        RECT 30.930 41.660 44.960 41.800 ;
        RECT 30.930 41.600 31.250 41.660 ;
        RECT 22.650 41.260 22.970 41.520 ;
        RECT 44.820 41.460 44.960 41.660 ;
        RECT 46.080 41.660 48.270 41.800 ;
        RECT 46.080 41.615 46.370 41.660 ;
        RECT 47.950 41.600 48.270 41.660 ;
        RECT 49.330 41.800 49.650 41.860 ;
        RECT 51.170 41.800 51.490 41.860 ;
        RECT 55.310 41.845 55.630 41.860 ;
        RECT 49.330 41.660 51.490 41.800 ;
        RECT 49.330 41.600 49.650 41.660 ;
        RECT 51.170 41.600 51.490 41.660 ;
        RECT 55.280 41.615 55.630 41.845 ;
        RECT 55.310 41.600 55.630 41.615 ;
        RECT 58.530 41.600 58.850 41.860 ;
        RECT 63.560 41.800 63.850 41.845 ;
        RECT 65.430 41.800 65.750 41.860 ;
        RECT 63.560 41.660 65.750 41.800 ;
        RECT 63.560 41.615 63.850 41.660 ;
        RECT 65.430 41.600 65.750 41.660 ;
        RECT 70.030 41.800 70.350 41.860 ;
        RECT 72.420 41.800 72.560 41.955 ;
        RECT 72.790 41.940 73.110 42.000 ;
        RECT 75.105 41.955 75.395 42.000 ;
        RECT 78.310 42.140 78.630 42.200 ;
        RECT 83.370 42.140 83.690 42.200 ;
        RECT 78.310 42.000 83.690 42.140 ;
        RECT 70.030 41.660 72.560 41.800 ;
        RECT 74.185 41.800 74.475 41.845 ;
        RECT 74.185 41.660 74.860 41.800 ;
        RECT 70.030 41.600 70.350 41.660 ;
        RECT 74.185 41.615 74.475 41.660 ;
        RECT 74.720 41.520 74.860 41.660 ;
        RECT 53.025 41.460 53.315 41.505 ;
        RECT 54.390 41.460 54.710 41.520 ;
        RECT 56.230 41.460 56.550 41.520 ;
        RECT 44.820 41.320 56.550 41.460 ;
        RECT 53.025 41.275 53.315 41.320 ;
        RECT 54.390 41.260 54.710 41.320 ;
        RECT 56.230 41.260 56.550 41.320 ;
        RECT 60.845 41.460 61.135 41.505 ;
        RECT 62.210 41.460 62.530 41.520 ;
        RECT 60.845 41.320 62.530 41.460 ;
        RECT 60.845 41.275 61.135 41.320 ;
        RECT 62.210 41.260 62.530 41.320 ;
        RECT 69.125 41.460 69.415 41.505 ;
        RECT 70.950 41.460 71.270 41.520 ;
        RECT 69.125 41.320 71.270 41.460 ;
        RECT 69.125 41.275 69.415 41.320 ;
        RECT 70.950 41.260 71.270 41.320 ;
        RECT 71.870 41.460 72.190 41.520 ;
        RECT 73.250 41.460 73.570 41.520 ;
        RECT 71.870 41.320 73.570 41.460 ;
        RECT 71.870 41.260 72.190 41.320 ;
        RECT 73.250 41.260 73.570 41.320 ;
        RECT 74.630 41.260 74.950 41.520 ;
        RECT 75.180 41.460 75.320 41.955 ;
        RECT 78.310 41.940 78.630 42.000 ;
        RECT 83.370 41.940 83.690 42.000 ;
        RECT 79.660 41.800 79.950 41.845 ;
        RECT 81.530 41.800 81.850 41.860 ;
        RECT 79.660 41.660 81.850 41.800 ;
        RECT 79.660 41.615 79.950 41.660 ;
        RECT 81.530 41.600 81.850 41.660 ;
        RECT 85.225 41.460 85.515 41.505 ;
        RECT 88.890 41.460 89.210 41.520 ;
        RECT 75.180 41.320 89.210 41.460 ;
        RECT 85.225 41.275 85.515 41.320 ;
        RECT 88.890 41.260 89.210 41.320 ;
        RECT 13.380 40.640 92.040 41.120 ;
        RECT 15.765 40.440 16.055 40.485 ;
        RECT 16.210 40.440 16.530 40.500 ;
        RECT 15.765 40.300 16.530 40.440 ;
        RECT 15.765 40.255 16.055 40.300 ;
        RECT 16.210 40.240 16.530 40.300 ;
        RECT 24.505 40.440 24.795 40.485 ;
        RECT 31.850 40.440 32.170 40.500 ;
        RECT 24.505 40.300 32.170 40.440 ;
        RECT 24.505 40.255 24.795 40.300 ;
        RECT 31.850 40.240 32.170 40.300 ;
        RECT 47.950 40.240 48.270 40.500 ;
        RECT 49.805 40.440 50.095 40.485 ;
        RECT 53.010 40.440 53.330 40.500 ;
        RECT 49.805 40.300 53.330 40.440 ;
        RECT 49.805 40.255 50.095 40.300 ;
        RECT 53.010 40.240 53.330 40.300 ;
        RECT 53.485 40.440 53.775 40.485 ;
        RECT 54.850 40.440 55.170 40.500 ;
        RECT 55.785 40.440 56.075 40.485 ;
        RECT 64.510 40.440 64.830 40.500 ;
        RECT 53.485 40.300 56.075 40.440 ;
        RECT 53.485 40.255 53.775 40.300 ;
        RECT 54.850 40.240 55.170 40.300 ;
        RECT 55.785 40.255 56.075 40.300 ;
        RECT 60.920 40.300 64.830 40.440 ;
        RECT 19.445 40.100 19.735 40.145 ;
        RECT 18.140 39.960 19.735 40.100 ;
        RECT 17.145 39.575 17.435 39.805 ;
        RECT 17.220 38.740 17.360 39.575 ;
        RECT 17.590 39.560 17.910 39.820 ;
        RECT 18.140 39.805 18.280 39.960 ;
        RECT 19.445 39.915 19.735 39.960 ;
        RECT 20.350 40.100 20.670 40.160 ;
        RECT 22.190 40.100 22.510 40.160 ;
        RECT 23.125 40.100 23.415 40.145 ;
        RECT 28.630 40.100 28.950 40.160 ;
        RECT 29.565 40.100 29.855 40.145 ;
        RECT 20.350 39.960 21.960 40.100 ;
        RECT 20.350 39.900 20.670 39.960 ;
        RECT 18.065 39.575 18.355 39.805 ;
        RECT 18.985 39.575 19.275 39.805 ;
        RECT 20.810 39.760 21.130 39.820 ;
        RECT 21.820 39.805 21.960 39.960 ;
        RECT 22.190 39.960 23.415 40.100 ;
        RECT 22.190 39.900 22.510 39.960 ;
        RECT 23.125 39.915 23.415 39.960 ;
        RECT 23.660 39.960 27.020 40.100 ;
        RECT 21.285 39.760 21.575 39.805 ;
        RECT 20.810 39.620 21.575 39.760 ;
        RECT 17.680 39.080 17.820 39.560 ;
        RECT 19.060 39.420 19.200 39.575 ;
        RECT 20.810 39.560 21.130 39.620 ;
        RECT 21.285 39.575 21.575 39.620 ;
        RECT 21.745 39.575 22.035 39.805 ;
        RECT 22.650 39.560 22.970 39.820 ;
        RECT 23.660 39.805 23.800 39.960 ;
        RECT 23.660 39.620 23.995 39.805 ;
        RECT 26.880 39.760 27.020 39.960 ;
        RECT 28.630 39.960 29.855 40.100 ;
        RECT 28.630 39.900 28.950 39.960 ;
        RECT 29.565 39.915 29.855 39.960 ;
        RECT 30.470 40.100 30.790 40.160 ;
        RECT 38.750 40.100 39.070 40.160 ;
        RECT 30.470 39.960 35.300 40.100 ;
        RECT 30.470 39.900 30.790 39.960 ;
        RECT 26.880 39.620 28.860 39.760 ;
        RECT 23.705 39.575 23.995 39.620 ;
        RECT 26.330 39.420 26.650 39.480 ;
        RECT 19.060 39.280 26.650 39.420 ;
        RECT 28.720 39.420 28.860 39.620 ;
        RECT 29.090 39.560 29.410 39.820 ;
        RECT 30.025 39.760 30.315 39.805 ;
        RECT 30.930 39.760 31.250 39.820 ;
        RECT 30.025 39.620 31.250 39.760 ;
        RECT 30.025 39.575 30.315 39.620 ;
        RECT 30.930 39.560 31.250 39.620 ;
        RECT 32.785 39.575 33.075 39.805 ;
        RECT 33.705 39.760 33.995 39.805 ;
        RECT 34.610 39.760 34.930 39.820 ;
        RECT 33.705 39.620 34.930 39.760 ;
        RECT 35.160 39.760 35.300 39.960 ;
        RECT 38.750 39.960 43.120 40.100 ;
        RECT 38.750 39.900 39.070 39.960 ;
        RECT 42.980 39.805 43.120 39.960 ;
        RECT 54.390 39.900 54.710 40.160 ;
        RECT 60.920 40.100 61.060 40.300 ;
        RECT 64.510 40.240 64.830 40.300 ;
        RECT 65.430 40.240 65.750 40.500 ;
        RECT 83.845 40.255 84.135 40.485 ;
        RECT 55.860 39.960 61.060 40.100 ;
        RECT 61.305 40.100 61.595 40.145 ;
        RECT 69.110 40.100 69.430 40.160 ;
        RECT 61.305 39.960 69.430 40.100 ;
        RECT 42.445 39.760 42.735 39.805 ;
        RECT 35.160 39.620 42.735 39.760 ;
        RECT 33.705 39.575 33.995 39.620 ;
        RECT 32.860 39.420 33.000 39.575 ;
        RECT 34.610 39.560 34.930 39.620 ;
        RECT 42.445 39.575 42.735 39.620 ;
        RECT 42.905 39.575 43.195 39.805 ;
        RECT 43.810 39.560 44.130 39.820 ;
        RECT 44.285 39.760 44.575 39.805 ;
        RECT 55.860 39.760 56.000 39.960 ;
        RECT 61.305 39.915 61.595 39.960 ;
        RECT 69.110 39.900 69.430 39.960 ;
        RECT 71.410 40.100 71.730 40.160 ;
        RECT 83.920 40.100 84.060 40.255 ;
        RECT 71.410 39.960 75.320 40.100 ;
        RECT 71.410 39.900 71.730 39.960 ;
        RECT 44.285 39.620 56.000 39.760 ;
        RECT 56.245 39.760 56.535 39.805 ;
        RECT 57.150 39.760 57.470 39.820 ;
        RECT 62.210 39.760 62.530 39.820 ;
        RECT 56.245 39.620 62.530 39.760 ;
        RECT 44.285 39.575 44.575 39.620 ;
        RECT 56.245 39.575 56.535 39.620 ;
        RECT 57.150 39.560 57.470 39.620 ;
        RECT 62.210 39.560 62.530 39.620 ;
        RECT 62.670 39.560 62.990 39.820 ;
        RECT 66.810 39.560 67.130 39.820 ;
        RECT 67.285 39.575 67.575 39.805 ;
        RECT 67.745 39.575 68.035 39.805 ;
        RECT 35.070 39.420 35.390 39.480 ;
        RECT 28.720 39.280 35.390 39.420 ;
        RECT 26.330 39.220 26.650 39.280 ;
        RECT 35.070 39.220 35.390 39.280 ;
        RECT 49.790 39.420 50.110 39.480 ;
        RECT 50.265 39.420 50.555 39.465 ;
        RECT 49.790 39.280 50.555 39.420 ;
        RECT 49.790 39.220 50.110 39.280 ;
        RECT 50.265 39.235 50.555 39.280 ;
        RECT 51.170 39.220 51.490 39.480 ;
        RECT 57.625 39.420 57.915 39.465 ;
        RECT 58.530 39.420 58.850 39.480 ;
        RECT 57.625 39.280 58.850 39.420 ;
        RECT 57.625 39.235 57.915 39.280 ;
        RECT 58.530 39.220 58.850 39.280 ;
        RECT 61.290 39.420 61.610 39.480 ;
        RECT 61.765 39.420 62.055 39.465 ;
        RECT 67.360 39.420 67.500 39.575 ;
        RECT 61.290 39.280 62.055 39.420 ;
        RECT 61.290 39.220 61.610 39.280 ;
        RECT 61.765 39.235 62.055 39.280 ;
        RECT 62.300 39.280 67.500 39.420 ;
        RECT 67.820 39.420 67.960 39.575 ;
        RECT 68.650 39.560 68.970 39.820 ;
        RECT 69.570 39.560 69.890 39.820 ;
        RECT 70.505 39.760 70.795 39.805 ;
        RECT 70.950 39.760 71.270 39.820 ;
        RECT 71.960 39.805 72.100 39.960 ;
        RECT 70.505 39.620 71.270 39.760 ;
        RECT 70.505 39.575 70.795 39.620 ;
        RECT 70.950 39.560 71.270 39.620 ;
        RECT 71.885 39.575 72.175 39.805 ;
        RECT 72.330 39.760 72.650 39.820 ;
        RECT 75.180 39.805 75.320 39.960 ;
        RECT 80.240 39.960 84.060 40.100 ;
        RECT 72.805 39.760 73.095 39.805 ;
        RECT 74.185 39.760 74.475 39.805 ;
        RECT 72.330 39.620 74.475 39.760 ;
        RECT 72.330 39.560 72.650 39.620 ;
        RECT 72.805 39.575 73.095 39.620 ;
        RECT 74.185 39.575 74.475 39.620 ;
        RECT 75.105 39.760 75.395 39.805 ;
        RECT 75.550 39.760 75.870 39.820 ;
        RECT 75.105 39.620 75.870 39.760 ;
        RECT 75.105 39.575 75.395 39.620 ;
        RECT 75.550 39.560 75.870 39.620 ;
        RECT 79.230 39.760 79.550 39.820 ;
        RECT 80.240 39.805 80.380 39.960 ;
        RECT 80.165 39.760 80.455 39.805 ;
        RECT 79.230 39.620 80.455 39.760 ;
        RECT 79.230 39.560 79.550 39.620 ;
        RECT 80.165 39.575 80.455 39.620 ;
        RECT 81.070 39.560 81.390 39.820 ;
        RECT 81.545 39.575 81.835 39.805 ;
        RECT 82.005 39.760 82.295 39.805 ;
        RECT 82.450 39.760 82.770 39.820 ;
        RECT 82.005 39.620 82.770 39.760 ;
        RECT 82.005 39.575 82.295 39.620 ;
        RECT 71.425 39.420 71.715 39.465 ;
        RECT 67.820 39.280 71.715 39.420 ;
        RECT 41.525 39.080 41.815 39.125 ;
        RECT 60.830 39.080 61.150 39.140 ;
        RECT 17.680 38.940 41.280 39.080 ;
        RECT 21.270 38.740 21.590 38.800 ;
        RECT 22.650 38.740 22.970 38.800 ;
        RECT 17.220 38.600 22.970 38.740 ;
        RECT 21.270 38.540 21.590 38.600 ;
        RECT 22.650 38.540 22.970 38.600 ;
        RECT 30.930 38.740 31.250 38.800 ;
        RECT 31.865 38.740 32.155 38.785 ;
        RECT 30.930 38.600 32.155 38.740 ;
        RECT 41.140 38.740 41.280 38.940 ;
        RECT 41.525 38.940 61.150 39.080 ;
        RECT 41.525 38.895 41.815 38.940 ;
        RECT 60.830 38.880 61.150 38.940 ;
        RECT 50.710 38.740 51.030 38.800 ;
        RECT 41.140 38.600 51.030 38.740 ;
        RECT 30.930 38.540 31.250 38.600 ;
        RECT 31.865 38.555 32.155 38.600 ;
        RECT 50.710 38.540 51.030 38.600 ;
        RECT 52.550 38.540 52.870 38.800 ;
        RECT 53.010 38.740 53.330 38.800 ;
        RECT 53.485 38.740 53.775 38.785 ;
        RECT 53.010 38.600 53.775 38.740 ;
        RECT 53.010 38.540 53.330 38.600 ;
        RECT 53.485 38.555 53.775 38.600 ;
        RECT 60.370 38.740 60.690 38.800 ;
        RECT 62.300 38.740 62.440 39.280 ;
        RECT 71.425 39.235 71.715 39.280 ;
        RECT 73.250 39.420 73.570 39.480 ;
        RECT 79.690 39.420 80.010 39.480 ;
        RECT 81.620 39.420 81.760 39.575 ;
        RECT 82.450 39.560 82.770 39.620 ;
        RECT 84.750 39.560 85.070 39.820 ;
        RECT 73.250 39.280 81.760 39.420 ;
        RECT 73.250 39.220 73.570 39.280 ;
        RECT 79.690 39.220 80.010 39.280 ;
        RECT 69.570 39.080 69.890 39.140 ;
        RECT 80.150 39.080 80.470 39.140 ;
        RECT 63.680 38.940 69.890 39.080 ;
        RECT 60.370 38.600 62.440 38.740 ;
        RECT 63.130 38.740 63.450 38.800 ;
        RECT 63.680 38.785 63.820 38.940 ;
        RECT 69.570 38.880 69.890 38.940 ;
        RECT 71.960 38.940 80.470 39.080 ;
        RECT 63.605 38.740 63.895 38.785 ;
        RECT 63.130 38.600 63.895 38.740 ;
        RECT 60.370 38.540 60.690 38.600 ;
        RECT 63.130 38.540 63.450 38.600 ;
        RECT 63.605 38.555 63.895 38.600 ;
        RECT 66.810 38.740 67.130 38.800 ;
        RECT 71.960 38.740 72.100 38.940 ;
        RECT 80.150 38.880 80.470 38.940 ;
        RECT 83.385 39.080 83.675 39.125 ;
        RECT 84.750 39.080 85.070 39.140 ;
        RECT 83.385 38.940 85.070 39.080 ;
        RECT 83.385 38.895 83.675 38.940 ;
        RECT 84.750 38.880 85.070 38.940 ;
        RECT 66.810 38.600 72.100 38.740 ;
        RECT 66.810 38.540 67.130 38.600 ;
        RECT 72.330 38.540 72.650 38.800 ;
        RECT 75.090 38.740 75.410 38.800 ;
        RECT 76.025 38.740 76.315 38.785 ;
        RECT 75.090 38.600 76.315 38.740 ;
        RECT 75.090 38.540 75.410 38.600 ;
        RECT 76.025 38.555 76.315 38.600 ;
        RECT 13.380 37.920 92.040 38.400 ;
        RECT 21.730 37.720 22.050 37.780 ;
        RECT 23.110 37.720 23.430 37.780 ;
        RECT 35.085 37.720 35.375 37.765 ;
        RECT 21.730 37.580 23.430 37.720 ;
        RECT 21.730 37.520 22.050 37.580 ;
        RECT 23.110 37.520 23.430 37.580 ;
        RECT 31.020 37.580 35.375 37.720 ;
        RECT 18.550 37.380 18.840 37.425 ;
        RECT 20.650 37.380 20.940 37.425 ;
        RECT 22.220 37.380 22.510 37.425 ;
        RECT 18.550 37.240 22.510 37.380 ;
        RECT 18.550 37.195 18.840 37.240 ;
        RECT 20.650 37.195 20.940 37.240 ;
        RECT 22.220 37.195 22.510 37.240 ;
        RECT 16.670 37.040 16.990 37.100 ;
        RECT 18.050 37.040 18.370 37.100 ;
        RECT 16.670 36.900 18.370 37.040 ;
        RECT 16.670 36.840 16.990 36.900 ;
        RECT 18.050 36.840 18.370 36.900 ;
        RECT 18.945 37.040 19.235 37.085 ;
        RECT 20.135 37.040 20.425 37.085 ;
        RECT 22.655 37.040 22.945 37.085 ;
        RECT 18.945 36.900 22.945 37.040 ;
        RECT 31.020 37.040 31.160 37.580 ;
        RECT 31.020 36.900 31.620 37.040 ;
        RECT 18.945 36.855 19.235 36.900 ;
        RECT 20.135 36.855 20.425 36.900 ;
        RECT 22.655 36.855 22.945 36.900 ;
        RECT 26.790 36.700 27.110 36.760 ;
        RECT 30.010 36.700 30.330 36.760 ;
        RECT 26.790 36.560 30.330 36.700 ;
        RECT 26.790 36.500 27.110 36.560 ;
        RECT 30.010 36.500 30.330 36.560 ;
        RECT 30.470 36.700 30.790 36.760 ;
        RECT 31.480 36.745 31.620 36.900 ;
        RECT 34.700 36.760 34.840 37.580 ;
        RECT 35.085 37.535 35.375 37.580 ;
        RECT 55.310 37.520 55.630 37.780 ;
        RECT 77.405 37.720 77.695 37.765 ;
        RECT 81.070 37.720 81.390 37.780 ;
        RECT 77.405 37.580 81.390 37.720 ;
        RECT 77.405 37.535 77.695 37.580 ;
        RECT 81.070 37.520 81.390 37.580 ;
        RECT 40.590 37.380 40.880 37.425 ;
        RECT 42.160 37.380 42.450 37.425 ;
        RECT 44.260 37.380 44.550 37.425 ;
        RECT 40.590 37.240 44.550 37.380 ;
        RECT 40.590 37.195 40.880 37.240 ;
        RECT 42.160 37.195 42.450 37.240 ;
        RECT 44.260 37.195 44.550 37.240 ;
        RECT 49.790 37.380 50.110 37.440 ;
        RECT 74.630 37.380 74.950 37.440 ;
        RECT 49.790 37.240 74.950 37.380 ;
        RECT 49.790 37.180 50.110 37.240 ;
        RECT 74.630 37.180 74.950 37.240 ;
        RECT 83.410 37.380 83.700 37.425 ;
        RECT 85.510 37.380 85.800 37.425 ;
        RECT 87.080 37.380 87.370 37.425 ;
        RECT 83.410 37.240 87.370 37.380 ;
        RECT 83.410 37.195 83.700 37.240 ;
        RECT 85.510 37.195 85.800 37.240 ;
        RECT 87.080 37.195 87.370 37.240 ;
        RECT 40.155 37.040 40.445 37.085 ;
        RECT 42.675 37.040 42.965 37.085 ;
        RECT 43.865 37.040 44.155 37.085 ;
        RECT 40.155 36.900 44.155 37.040 ;
        RECT 40.155 36.855 40.445 36.900 ;
        RECT 42.675 36.855 42.965 36.900 ;
        RECT 43.865 36.855 44.155 36.900 ;
        RECT 51.170 37.040 51.490 37.100 ;
        RECT 58.085 37.040 58.375 37.085 ;
        RECT 51.170 36.900 58.375 37.040 ;
        RECT 51.170 36.840 51.490 36.900 ;
        RECT 58.085 36.855 58.375 36.900 ;
        RECT 62.210 36.840 62.530 37.100 ;
        RECT 82.450 37.040 82.770 37.100 ;
        RECT 81.160 36.900 82.770 37.040 ;
        RECT 30.945 36.700 31.235 36.745 ;
        RECT 30.470 36.560 31.235 36.700 ;
        RECT 30.470 36.500 30.790 36.560 ;
        RECT 30.945 36.515 31.235 36.560 ;
        RECT 31.405 36.515 31.695 36.745 ;
        RECT 31.850 36.500 32.170 36.760 ;
        RECT 34.150 36.500 34.470 36.760 ;
        RECT 34.610 36.500 34.930 36.760 ;
        RECT 35.070 36.700 35.390 36.760 ;
        RECT 35.545 36.700 35.835 36.745 ;
        RECT 40.590 36.700 40.910 36.760 ;
        RECT 44.730 36.700 45.050 36.760 ;
        RECT 35.070 36.560 40.910 36.700 ;
        RECT 35.070 36.500 35.390 36.560 ;
        RECT 35.545 36.515 35.835 36.560 ;
        RECT 40.590 36.500 40.910 36.560 ;
        RECT 42.520 36.560 45.050 36.700 ;
        RECT 19.400 36.360 19.690 36.405 ;
        RECT 21.270 36.360 21.590 36.420 ;
        RECT 27.725 36.360 28.015 36.405 ;
        RECT 19.400 36.220 21.590 36.360 ;
        RECT 19.400 36.175 19.690 36.220 ;
        RECT 21.270 36.160 21.590 36.220 ;
        RECT 25.040 36.220 28.015 36.360 ;
        RECT 22.190 36.020 22.510 36.080 ;
        RECT 25.040 36.065 25.180 36.220 ;
        RECT 27.725 36.175 28.015 36.220 ;
        RECT 28.630 36.160 28.950 36.420 ;
        RECT 31.940 36.360 32.080 36.500 ;
        RECT 42.520 36.420 42.660 36.560 ;
        RECT 44.730 36.500 45.050 36.560 ;
        RECT 46.585 36.515 46.875 36.745 ;
        RECT 31.940 36.220 38.520 36.360 ;
        RECT 24.965 36.020 25.255 36.065 ;
        RECT 22.190 35.880 25.255 36.020 ;
        RECT 22.190 35.820 22.510 35.880 ;
        RECT 24.965 35.835 25.255 35.880 ;
        RECT 26.790 35.820 27.110 36.080 ;
        RECT 28.720 36.020 28.860 36.160 ;
        RECT 30.930 36.020 31.250 36.080 ;
        RECT 28.720 35.880 31.250 36.020 ;
        RECT 30.930 35.820 31.250 35.880 ;
        RECT 31.390 36.020 31.710 36.080 ;
        RECT 33.245 36.020 33.535 36.065 ;
        RECT 31.390 35.880 33.535 36.020 ;
        RECT 31.390 35.820 31.710 35.880 ;
        RECT 33.245 35.835 33.535 35.880 ;
        RECT 37.830 35.820 38.150 36.080 ;
        RECT 38.380 36.020 38.520 36.220 ;
        RECT 42.430 36.160 42.750 36.420 ;
        RECT 43.520 36.360 43.810 36.405 ;
        RECT 45.205 36.360 45.495 36.405 ;
        RECT 43.520 36.220 45.495 36.360 ;
        RECT 43.520 36.175 43.810 36.220 ;
        RECT 45.205 36.175 45.495 36.220 ;
        RECT 46.660 36.360 46.800 36.515 ;
        RECT 47.030 36.500 47.350 36.760 ;
        RECT 47.490 36.500 47.810 36.760 ;
        RECT 47.950 36.700 48.270 36.760 ;
        RECT 48.425 36.700 48.715 36.745 ;
        RECT 66.810 36.700 67.130 36.760 ;
        RECT 47.950 36.560 48.715 36.700 ;
        RECT 47.950 36.500 48.270 36.560 ;
        RECT 48.425 36.515 48.715 36.560 ;
        RECT 56.780 36.560 67.130 36.700 ;
        RECT 56.780 36.360 56.920 36.560 ;
        RECT 66.810 36.500 67.130 36.560 ;
        RECT 79.230 36.500 79.550 36.760 ;
        RECT 80.150 36.500 80.470 36.760 ;
        RECT 81.160 36.745 81.300 36.900 ;
        RECT 82.450 36.840 82.770 36.900 ;
        RECT 83.805 37.040 84.095 37.085 ;
        RECT 84.995 37.040 85.285 37.085 ;
        RECT 87.515 37.040 87.805 37.085 ;
        RECT 83.805 36.900 87.805 37.040 ;
        RECT 83.805 36.855 84.095 36.900 ;
        RECT 84.995 36.855 85.285 36.900 ;
        RECT 87.515 36.855 87.805 36.900 ;
        RECT 80.625 36.515 80.915 36.745 ;
        RECT 81.085 36.515 81.375 36.745 ;
        RECT 82.925 36.700 83.215 36.745 ;
        RECT 83.370 36.700 83.690 36.760 ;
        RECT 82.925 36.560 83.690 36.700 ;
        RECT 82.925 36.515 83.215 36.560 ;
        RECT 46.660 36.220 56.920 36.360 ;
        RECT 57.165 36.360 57.455 36.405 ;
        RECT 59.465 36.360 59.755 36.405 ;
        RECT 57.165 36.220 59.755 36.360 ;
        RECT 46.660 36.020 46.800 36.220 ;
        RECT 57.165 36.175 57.455 36.220 ;
        RECT 59.465 36.175 59.755 36.220 ;
        RECT 63.590 36.160 63.910 36.420 ;
        RECT 75.090 36.360 75.410 36.420 ;
        RECT 75.565 36.360 75.855 36.405 ;
        RECT 75.090 36.220 75.855 36.360 ;
        RECT 75.090 36.160 75.410 36.220 ;
        RECT 75.565 36.175 75.855 36.220 ;
        RECT 76.485 36.360 76.775 36.405 ;
        RECT 79.690 36.360 80.010 36.420 ;
        RECT 76.485 36.220 80.010 36.360 ;
        RECT 76.485 36.175 76.775 36.220 ;
        RECT 79.690 36.160 80.010 36.220 ;
        RECT 38.380 35.880 46.800 36.020 ;
        RECT 57.625 36.020 57.915 36.065 ;
        RECT 58.070 36.020 58.390 36.080 ;
        RECT 57.625 35.880 58.390 36.020 ;
        RECT 57.625 35.835 57.915 35.880 ;
        RECT 58.070 35.820 58.390 35.880 ;
        RECT 64.050 35.820 64.370 36.080 ;
        RECT 74.170 36.020 74.490 36.080 ;
        RECT 80.700 36.020 80.840 36.515 ;
        RECT 83.370 36.500 83.690 36.560 ;
        RECT 82.465 36.360 82.755 36.405 ;
        RECT 84.150 36.360 84.440 36.405 ;
        RECT 82.465 36.220 84.440 36.360 ;
        RECT 82.465 36.175 82.755 36.220 ;
        RECT 84.150 36.175 84.440 36.220 ;
        RECT 74.170 35.880 80.840 36.020 ;
        RECT 87.050 36.020 87.370 36.080 ;
        RECT 89.825 36.020 90.115 36.065 ;
        RECT 87.050 35.880 90.115 36.020 ;
        RECT 74.170 35.820 74.490 35.880 ;
        RECT 87.050 35.820 87.370 35.880 ;
        RECT 89.825 35.835 90.115 35.880 ;
        RECT 13.380 35.200 92.040 35.680 ;
        RECT 21.270 34.800 21.590 35.060 ;
        RECT 30.470 34.800 30.790 35.060 ;
        RECT 30.930 35.000 31.250 35.060 ;
        RECT 34.150 35.000 34.470 35.060 ;
        RECT 30.930 34.860 34.470 35.000 ;
        RECT 30.930 34.800 31.250 34.860 ;
        RECT 34.150 34.800 34.470 34.860 ;
        RECT 42.445 35.000 42.735 35.045 ;
        RECT 42.890 35.000 43.210 35.060 ;
        RECT 42.445 34.860 43.210 35.000 ;
        RECT 42.445 34.815 42.735 34.860 ;
        RECT 42.890 34.800 43.210 34.860 ;
        RECT 44.745 35.000 45.035 35.045 ;
        RECT 47.490 35.000 47.810 35.060 ;
        RECT 44.745 34.860 47.810 35.000 ;
        RECT 44.745 34.815 45.035 34.860 ;
        RECT 47.490 34.800 47.810 34.860 ;
        RECT 51.170 35.000 51.490 35.060 ;
        RECT 53.025 35.000 53.315 35.045 ;
        RECT 63.590 35.000 63.910 35.060 ;
        RECT 51.170 34.860 63.910 35.000 ;
        RECT 51.170 34.800 51.490 34.860 ;
        RECT 53.025 34.815 53.315 34.860 ;
        RECT 63.590 34.800 63.910 34.860 ;
        RECT 67.270 35.000 67.590 35.060 ;
        RECT 78.785 35.000 79.075 35.045 ;
        RECT 80.150 35.000 80.470 35.060 ;
        RECT 88.890 35.000 89.210 35.060 ;
        RECT 90.285 35.000 90.575 35.045 ;
        RECT 67.270 34.860 75.780 35.000 ;
        RECT 67.270 34.800 67.590 34.860 ;
        RECT 75.640 34.720 75.780 34.860 ;
        RECT 78.785 34.860 80.470 35.000 ;
        RECT 78.785 34.815 79.075 34.860 ;
        RECT 80.150 34.800 80.470 34.860 ;
        RECT 80.700 34.860 90.575 35.000 ;
        RECT 26.790 34.660 27.110 34.720 ;
        RECT 30.010 34.660 30.330 34.720 ;
        RECT 35.070 34.660 35.390 34.720 ;
        RECT 23.660 34.520 27.110 34.660 ;
        RECT 22.650 34.120 22.970 34.380 ;
        RECT 23.110 34.120 23.430 34.380 ;
        RECT 23.660 34.365 23.800 34.520 ;
        RECT 26.790 34.460 27.110 34.520 ;
        RECT 27.340 34.520 30.330 34.660 ;
        RECT 23.585 34.135 23.875 34.365 ;
        RECT 24.505 34.135 24.795 34.365 ;
        RECT 24.965 34.320 25.255 34.365 ;
        RECT 27.340 34.320 27.480 34.520 ;
        RECT 30.010 34.460 30.330 34.520 ;
        RECT 31.020 34.520 35.390 34.660 ;
        RECT 24.965 34.180 27.480 34.320 ;
        RECT 24.965 34.135 25.255 34.180 ;
        RECT 24.580 33.980 24.720 34.135 ;
        RECT 28.630 34.120 28.950 34.380 ;
        RECT 31.020 34.365 31.160 34.520 ;
        RECT 35.070 34.460 35.390 34.520 ;
        RECT 37.830 34.660 38.150 34.720 ;
        RECT 41.065 34.660 41.355 34.705 ;
        RECT 43.825 34.660 44.115 34.705 ;
        RECT 37.830 34.520 44.115 34.660 ;
        RECT 37.830 34.460 38.150 34.520 ;
        RECT 41.065 34.475 41.355 34.520 ;
        RECT 43.825 34.475 44.115 34.520 ;
        RECT 55.770 34.660 56.090 34.720 ;
        RECT 69.570 34.660 69.890 34.720 ;
        RECT 55.770 34.520 69.890 34.660 ;
        RECT 55.770 34.460 56.090 34.520 ;
        RECT 69.570 34.460 69.890 34.520 ;
        RECT 75.550 34.660 75.870 34.720 ;
        RECT 79.690 34.660 80.010 34.720 ;
        RECT 80.700 34.705 80.840 34.860 ;
        RECT 88.890 34.800 89.210 34.860 ;
        RECT 90.285 34.815 90.575 34.860 ;
        RECT 84.750 34.705 85.070 34.720 ;
        RECT 80.625 34.660 80.915 34.705 ;
        RECT 84.720 34.660 85.070 34.705 ;
        RECT 75.550 34.520 78.540 34.660 ;
        RECT 75.550 34.460 75.870 34.520 ;
        RECT 29.565 34.320 29.855 34.365 ;
        RECT 29.565 34.180 30.700 34.320 ;
        RECT 29.565 34.135 29.855 34.180 ;
        RECT 24.580 33.840 26.100 33.980 ;
        RECT 25.960 33.345 26.100 33.840 ;
        RECT 25.885 33.300 26.175 33.345 ;
        RECT 27.250 33.300 27.570 33.360 ;
        RECT 25.885 33.160 27.570 33.300 ;
        RECT 30.560 33.300 30.700 34.180 ;
        RECT 30.945 34.135 31.235 34.365 ;
        RECT 31.390 34.320 31.710 34.380 ;
        RECT 32.225 34.320 32.515 34.365 ;
        RECT 39.685 34.320 39.975 34.365 ;
        RECT 31.390 34.180 32.515 34.320 ;
        RECT 31.390 34.120 31.710 34.180 ;
        RECT 32.225 34.135 32.515 34.180 ;
        RECT 37.920 34.180 39.975 34.320 ;
        RECT 31.825 33.980 32.115 34.025 ;
        RECT 33.015 33.980 33.305 34.025 ;
        RECT 35.535 33.980 35.825 34.025 ;
        RECT 31.825 33.840 35.825 33.980 ;
        RECT 31.825 33.795 32.115 33.840 ;
        RECT 33.015 33.795 33.305 33.840 ;
        RECT 35.535 33.795 35.825 33.840 ;
        RECT 31.430 33.640 31.720 33.685 ;
        RECT 33.530 33.640 33.820 33.685 ;
        RECT 35.100 33.640 35.390 33.685 ;
        RECT 31.430 33.500 35.390 33.640 ;
        RECT 31.430 33.455 31.720 33.500 ;
        RECT 33.530 33.455 33.820 33.500 ;
        RECT 35.100 33.455 35.390 33.500 ;
        RECT 31.850 33.300 32.170 33.360 ;
        RECT 37.920 33.345 38.060 34.180 ;
        RECT 39.685 34.135 39.975 34.180 ;
        RECT 40.590 34.120 40.910 34.380 ;
        RECT 41.525 34.135 41.815 34.365 ;
        RECT 40.680 33.640 40.820 34.120 ;
        RECT 41.600 33.980 41.740 34.135 ;
        RECT 42.890 34.120 43.210 34.380 ;
        RECT 52.090 34.320 52.410 34.380 ;
        RECT 52.565 34.320 52.855 34.365 ;
        RECT 52.090 34.180 52.855 34.320 ;
        RECT 52.090 34.120 52.410 34.180 ;
        RECT 52.565 34.135 52.855 34.180 ;
        RECT 53.010 34.320 53.330 34.380 ;
        RECT 53.945 34.320 54.235 34.365 ;
        RECT 53.010 34.180 54.235 34.320 ;
        RECT 53.010 34.120 53.330 34.180 ;
        RECT 53.945 34.135 54.235 34.180 ;
        RECT 54.850 34.120 55.170 34.380 ;
        RECT 57.150 34.320 57.470 34.380 ;
        RECT 58.905 34.320 59.195 34.365 ;
        RECT 57.150 34.180 59.195 34.320 ;
        RECT 57.150 34.120 57.470 34.180 ;
        RECT 58.905 34.135 59.195 34.180 ;
        RECT 64.050 34.320 64.370 34.380 ;
        RECT 70.965 34.320 71.255 34.365 ;
        RECT 72.345 34.320 72.635 34.365 ;
        RECT 64.050 34.180 72.635 34.320 ;
        RECT 64.050 34.120 64.370 34.180 ;
        RECT 43.350 33.980 43.670 34.040 ;
        RECT 41.600 33.840 43.670 33.980 ;
        RECT 43.350 33.780 43.670 33.840 ;
        RECT 57.625 33.795 57.915 34.025 ;
        RECT 58.505 33.980 58.795 34.025 ;
        RECT 59.695 33.980 59.985 34.025 ;
        RECT 62.215 33.980 62.505 34.025 ;
        RECT 58.505 33.840 62.505 33.980 ;
        RECT 58.505 33.795 58.795 33.840 ;
        RECT 59.695 33.795 59.985 33.840 ;
        RECT 62.215 33.795 62.505 33.840 ;
        RECT 52.550 33.640 52.870 33.700 ;
        RECT 40.680 33.500 52.870 33.640 ;
        RECT 52.550 33.440 52.870 33.500 ;
        RECT 37.845 33.300 38.135 33.345 ;
        RECT 30.560 33.160 38.135 33.300 ;
        RECT 57.700 33.300 57.840 33.795 ;
        RECT 58.110 33.640 58.400 33.685 ;
        RECT 60.210 33.640 60.500 33.685 ;
        RECT 61.780 33.640 62.070 33.685 ;
        RECT 58.110 33.500 62.070 33.640 ;
        RECT 58.110 33.455 58.400 33.500 ;
        RECT 60.210 33.455 60.500 33.500 ;
        RECT 61.780 33.455 62.070 33.500 ;
        RECT 58.530 33.300 58.850 33.360 ;
        RECT 57.700 33.160 58.850 33.300 ;
        RECT 25.885 33.115 26.175 33.160 ;
        RECT 27.250 33.100 27.570 33.160 ;
        RECT 31.850 33.100 32.170 33.160 ;
        RECT 37.845 33.115 38.135 33.160 ;
        RECT 58.530 33.100 58.850 33.160 ;
        RECT 58.990 33.300 59.310 33.360 ;
        RECT 64.525 33.300 64.815 33.345 ;
        RECT 64.970 33.300 65.290 33.360 ;
        RECT 58.990 33.160 65.290 33.300 ;
        RECT 69.660 33.300 69.800 34.180 ;
        RECT 70.965 34.135 71.255 34.180 ;
        RECT 72.345 34.135 72.635 34.180 ;
        RECT 73.265 34.135 73.555 34.365 ;
        RECT 76.945 34.135 77.235 34.365 ;
        RECT 77.390 34.320 77.710 34.380 ;
        RECT 77.865 34.320 78.155 34.365 ;
        RECT 77.390 34.180 78.155 34.320 ;
        RECT 78.400 34.320 78.540 34.520 ;
        RECT 79.690 34.520 80.915 34.660 ;
        RECT 84.555 34.520 85.070 34.660 ;
        RECT 79.690 34.460 80.010 34.520 ;
        RECT 80.625 34.475 80.915 34.520 ;
        RECT 84.720 34.475 85.070 34.520 ;
        RECT 84.750 34.460 85.070 34.475 ;
        RECT 80.150 34.320 80.470 34.380 ;
        RECT 78.400 34.180 80.470 34.320 ;
        RECT 71.870 33.980 72.190 34.040 ;
        RECT 73.340 33.980 73.480 34.135 ;
        RECT 71.870 33.840 73.480 33.980 ;
        RECT 71.870 33.780 72.190 33.840 ;
        RECT 74.170 33.780 74.490 34.040 ;
        RECT 77.020 33.700 77.160 34.135 ;
        RECT 77.390 34.120 77.710 34.180 ;
        RECT 77.865 34.135 78.155 34.180 ;
        RECT 80.150 34.120 80.470 34.180 ;
        RECT 81.070 34.120 81.390 34.380 ;
        RECT 81.990 34.320 82.310 34.380 ;
        RECT 87.050 34.320 87.370 34.380 ;
        RECT 81.990 34.180 87.370 34.320 ;
        RECT 81.990 34.120 82.310 34.180 ;
        RECT 87.050 34.120 87.370 34.180 ;
        RECT 83.370 33.780 83.690 34.040 ;
        RECT 84.265 33.980 84.555 34.025 ;
        RECT 85.455 33.980 85.745 34.025 ;
        RECT 87.975 33.980 88.265 34.025 ;
        RECT 84.265 33.840 88.265 33.980 ;
        RECT 84.265 33.795 84.555 33.840 ;
        RECT 85.455 33.795 85.745 33.840 ;
        RECT 87.975 33.795 88.265 33.840 ;
        RECT 70.045 33.640 70.335 33.685 ;
        RECT 76.930 33.640 77.250 33.700 ;
        RECT 70.045 33.500 77.250 33.640 ;
        RECT 70.045 33.455 70.335 33.500 ;
        RECT 76.930 33.440 77.250 33.500 ;
        RECT 77.850 33.640 78.170 33.700 ;
        RECT 79.245 33.640 79.535 33.685 ;
        RECT 77.850 33.500 79.535 33.640 ;
        RECT 77.850 33.440 78.170 33.500 ;
        RECT 79.245 33.455 79.535 33.500 ;
        RECT 80.150 33.640 80.470 33.700 ;
        RECT 82.450 33.640 82.770 33.700 ;
        RECT 80.150 33.500 82.770 33.640 ;
        RECT 80.150 33.440 80.470 33.500 ;
        RECT 82.450 33.440 82.770 33.500 ;
        RECT 83.870 33.640 84.160 33.685 ;
        RECT 85.970 33.640 86.260 33.685 ;
        RECT 87.540 33.640 87.830 33.685 ;
        RECT 83.870 33.500 87.830 33.640 ;
        RECT 83.870 33.455 84.160 33.500 ;
        RECT 85.970 33.455 86.260 33.500 ;
        RECT 87.540 33.455 87.830 33.500 ;
        RECT 81.070 33.300 81.390 33.360 ;
        RECT 69.660 33.160 81.390 33.300 ;
        RECT 58.990 33.100 59.310 33.160 ;
        RECT 64.525 33.115 64.815 33.160 ;
        RECT 64.970 33.100 65.290 33.160 ;
        RECT 81.070 33.100 81.390 33.160 ;
        RECT 13.380 32.480 92.040 32.960 ;
        RECT 21.590 32.140 51.400 32.280 ;
        RECT 18.970 31.940 19.290 32.000 ;
        RECT 20.810 31.940 21.130 32.000 ;
        RECT 21.590 31.940 21.730 32.140 ;
        RECT 18.970 31.800 21.730 31.940 ;
        RECT 23.110 31.940 23.430 32.000 ;
        RECT 23.110 31.800 23.800 31.940 ;
        RECT 18.970 31.740 19.290 31.800 ;
        RECT 20.810 31.740 21.130 31.800 ;
        RECT 23.110 31.740 23.430 31.800 ;
        RECT 22.190 31.600 22.510 31.660 ;
        RECT 16.300 31.460 22.510 31.600 ;
        RECT 16.300 31.305 16.440 31.460 ;
        RECT 22.190 31.400 22.510 31.460 ;
        RECT 23.660 31.600 23.800 31.800 ;
        RECT 42.890 31.740 43.210 32.000 ;
        RECT 51.260 31.940 51.400 32.140 ;
        RECT 51.630 32.080 51.950 32.340 ;
        RECT 57.150 32.080 57.470 32.340 ;
        RECT 68.740 32.140 76.700 32.280 ;
        RECT 60.410 31.940 60.700 31.985 ;
        RECT 62.510 31.940 62.800 31.985 ;
        RECT 64.080 31.940 64.370 31.985 ;
        RECT 51.260 31.800 58.300 31.940 ;
        RECT 34.610 31.600 34.930 31.660 ;
        RECT 42.980 31.600 43.120 31.740 ;
        RECT 49.790 31.600 50.110 31.660 ;
        RECT 52.090 31.600 52.410 31.660 ;
        RECT 57.625 31.600 57.915 31.645 ;
        RECT 23.660 31.460 34.930 31.600 ;
        RECT 16.225 31.075 16.515 31.305 ;
        RECT 16.670 31.260 16.990 31.320 ;
        RECT 18.970 31.260 19.290 31.320 ;
        RECT 16.670 31.120 19.290 31.260 ;
        RECT 16.670 31.060 16.990 31.120 ;
        RECT 18.970 31.060 19.290 31.120 ;
        RECT 19.430 31.260 19.750 31.320 ;
        RECT 23.660 31.305 23.800 31.460 ;
        RECT 34.610 31.400 34.930 31.460 ;
        RECT 42.520 31.460 50.110 31.600 ;
        RECT 23.125 31.260 23.415 31.305 ;
        RECT 19.430 31.120 23.415 31.260 ;
        RECT 19.430 31.060 19.750 31.120 ;
        RECT 23.125 31.075 23.415 31.120 ;
        RECT 23.585 31.075 23.875 31.305 ;
        RECT 24.030 31.060 24.350 31.320 ;
        RECT 24.965 31.260 25.255 31.305 ;
        RECT 25.410 31.260 25.730 31.320 ;
        RECT 27.250 31.260 27.570 31.320 ;
        RECT 24.965 31.120 27.570 31.260 ;
        RECT 24.965 31.075 25.255 31.120 ;
        RECT 25.410 31.060 25.730 31.120 ;
        RECT 27.250 31.060 27.570 31.120 ;
        RECT 18.065 30.920 18.355 30.965 ;
        RECT 18.510 30.920 18.830 30.980 ;
        RECT 18.065 30.780 18.830 30.920 ;
        RECT 42.520 30.920 42.660 31.460 ;
        RECT 49.790 31.400 50.110 31.460 ;
        RECT 50.340 31.460 52.410 31.600 ;
        RECT 42.890 31.260 43.210 31.320 ;
        RECT 48.885 31.260 49.175 31.305 ;
        RECT 42.890 31.120 49.175 31.260 ;
        RECT 42.890 31.060 43.210 31.120 ;
        RECT 48.885 31.075 49.175 31.120 ;
        RECT 44.285 30.920 44.575 30.965 ;
        RECT 42.520 30.780 44.575 30.920 ;
        RECT 18.065 30.735 18.355 30.780 ;
        RECT 18.510 30.720 18.830 30.780 ;
        RECT 44.285 30.735 44.575 30.780 ;
        RECT 45.205 30.920 45.495 30.965 ;
        RECT 45.650 30.920 45.970 30.980 ;
        RECT 50.340 30.965 50.480 31.460 ;
        RECT 52.090 31.400 52.410 31.460 ;
        RECT 54.940 31.460 57.915 31.600 ;
        RECT 50.725 31.260 51.015 31.305 ;
        RECT 51.630 31.260 51.950 31.320 ;
        RECT 50.725 31.120 51.950 31.260 ;
        RECT 50.725 31.075 51.015 31.120 ;
        RECT 51.630 31.060 51.950 31.120 ;
        RECT 53.930 31.060 54.250 31.320 ;
        RECT 54.940 31.305 55.080 31.460 ;
        RECT 57.625 31.415 57.915 31.460 ;
        RECT 54.865 31.075 55.155 31.305 ;
        RECT 55.325 31.075 55.615 31.305 ;
        RECT 45.205 30.780 45.970 30.920 ;
        RECT 45.205 30.735 45.495 30.780 ;
        RECT 45.650 30.720 45.970 30.780 ;
        RECT 49.805 30.735 50.095 30.965 ;
        RECT 50.265 30.735 50.555 30.965 ;
        RECT 51.170 30.920 51.490 30.980 ;
        RECT 55.400 30.920 55.540 31.075 ;
        RECT 55.770 31.060 56.090 31.320 ;
        RECT 58.160 31.260 58.300 31.800 ;
        RECT 60.410 31.800 64.370 31.940 ;
        RECT 60.410 31.755 60.700 31.800 ;
        RECT 62.510 31.755 62.800 31.800 ;
        RECT 64.080 31.755 64.370 31.800 ;
        RECT 58.530 31.600 58.850 31.660 ;
        RECT 59.925 31.600 60.215 31.645 ;
        RECT 58.530 31.460 60.215 31.600 ;
        RECT 58.530 31.400 58.850 31.460 ;
        RECT 59.925 31.415 60.215 31.460 ;
        RECT 60.805 31.600 61.095 31.645 ;
        RECT 61.995 31.600 62.285 31.645 ;
        RECT 64.515 31.600 64.805 31.645 ;
        RECT 60.805 31.460 64.805 31.600 ;
        RECT 60.805 31.415 61.095 31.460 ;
        RECT 61.995 31.415 62.285 31.460 ;
        RECT 64.515 31.415 64.805 31.460 ;
        RECT 59.465 31.260 59.755 31.305 ;
        RECT 63.130 31.260 63.450 31.320 ;
        RECT 64.050 31.260 64.370 31.320 ;
        RECT 58.160 31.120 64.370 31.260 ;
        RECT 59.465 31.075 59.755 31.120 ;
        RECT 63.130 31.060 63.450 31.120 ;
        RECT 64.050 31.060 64.370 31.120 ;
        RECT 67.730 31.260 68.050 31.320 ;
        RECT 68.205 31.260 68.495 31.305 ;
        RECT 68.740 31.260 68.880 32.140 ;
        RECT 76.560 31.985 76.700 32.140 ;
        RECT 70.070 31.940 70.360 31.985 ;
        RECT 72.170 31.940 72.460 31.985 ;
        RECT 73.740 31.940 74.030 31.985 ;
        RECT 70.070 31.800 74.030 31.940 ;
        RECT 70.070 31.755 70.360 31.800 ;
        RECT 72.170 31.755 72.460 31.800 ;
        RECT 73.740 31.755 74.030 31.800 ;
        RECT 76.485 31.940 76.775 31.985 ;
        RECT 83.830 31.940 84.150 32.000 ;
        RECT 76.485 31.800 84.150 31.940 ;
        RECT 76.485 31.755 76.775 31.800 ;
        RECT 83.830 31.740 84.150 31.800 ;
        RECT 70.465 31.600 70.755 31.645 ;
        RECT 71.655 31.600 71.945 31.645 ;
        RECT 74.175 31.600 74.465 31.645 ;
        RECT 70.465 31.460 74.465 31.600 ;
        RECT 70.465 31.415 70.755 31.460 ;
        RECT 71.655 31.415 71.945 31.460 ;
        RECT 74.175 31.415 74.465 31.460 ;
        RECT 67.730 31.120 68.880 31.260 ;
        RECT 69.585 31.260 69.875 31.305 ;
        RECT 73.250 31.260 73.570 31.320 ;
        RECT 69.585 31.120 73.570 31.260 ;
        RECT 67.730 31.060 68.050 31.120 ;
        RECT 68.205 31.075 68.495 31.120 ;
        RECT 69.585 31.075 69.875 31.120 ;
        RECT 73.250 31.060 73.570 31.120 ;
        RECT 88.890 31.060 89.210 31.320 ;
        RECT 51.170 30.780 55.540 30.920 ;
        RECT 15.305 30.580 15.595 30.625 ;
        RECT 15.750 30.580 16.070 30.640 ;
        RECT 15.305 30.440 16.070 30.580 ;
        RECT 15.305 30.395 15.595 30.440 ;
        RECT 15.750 30.380 16.070 30.440 ;
        RECT 17.145 30.580 17.435 30.625 ;
        RECT 17.590 30.580 17.910 30.640 ;
        RECT 17.145 30.440 17.910 30.580 ;
        RECT 17.145 30.395 17.435 30.440 ;
        RECT 17.590 30.380 17.910 30.440 ;
        RECT 21.730 30.380 22.050 30.640 ;
        RECT 46.110 30.380 46.430 30.640 ;
        RECT 49.880 30.580 50.020 30.735 ;
        RECT 51.170 30.720 51.490 30.780 ;
        RECT 52.550 30.580 52.870 30.640 ;
        RECT 49.880 30.440 52.870 30.580 ;
        RECT 55.400 30.580 55.540 30.780 ;
        RECT 57.610 30.920 57.930 30.980 ;
        RECT 58.545 30.920 58.835 30.965 ;
        RECT 58.990 30.920 59.310 30.980 ;
        RECT 57.610 30.780 59.310 30.920 ;
        RECT 57.610 30.720 57.930 30.780 ;
        RECT 58.545 30.735 58.835 30.780 ;
        RECT 58.990 30.720 59.310 30.780 ;
        RECT 59.910 30.920 60.230 30.980 ;
        RECT 61.150 30.920 61.440 30.965 ;
        RECT 59.910 30.780 61.440 30.920 ;
        RECT 59.910 30.720 60.230 30.780 ;
        RECT 61.150 30.735 61.440 30.780 ;
        RECT 69.125 30.920 69.415 30.965 ;
        RECT 70.920 30.920 71.210 30.965 ;
        RECT 72.790 30.920 73.110 30.980 ;
        RECT 69.125 30.780 70.720 30.920 ;
        RECT 69.125 30.735 69.415 30.780 ;
        RECT 60.370 30.580 60.690 30.640 ;
        RECT 55.400 30.440 60.690 30.580 ;
        RECT 52.550 30.380 52.870 30.440 ;
        RECT 60.370 30.380 60.690 30.440 ;
        RECT 63.130 30.580 63.450 30.640 ;
        RECT 66.825 30.580 67.115 30.625 ;
        RECT 63.130 30.440 67.115 30.580 ;
        RECT 63.130 30.380 63.450 30.440 ;
        RECT 66.825 30.395 67.115 30.440 ;
        RECT 67.285 30.580 67.575 30.625 ;
        RECT 70.030 30.580 70.350 30.640 ;
        RECT 67.285 30.440 70.350 30.580 ;
        RECT 70.580 30.580 70.720 30.780 ;
        RECT 70.920 30.780 73.110 30.920 ;
        RECT 70.920 30.735 71.210 30.780 ;
        RECT 72.790 30.720 73.110 30.780 ;
        RECT 75.090 30.920 75.410 30.980 ;
        RECT 78.785 30.920 79.075 30.965 ;
        RECT 75.090 30.780 79.075 30.920 ;
        RECT 75.090 30.720 75.410 30.780 ;
        RECT 78.785 30.735 79.075 30.780 ;
        RECT 79.690 30.720 80.010 30.980 ;
        RECT 75.180 30.580 75.320 30.720 ;
        RECT 70.580 30.440 75.320 30.580 ;
        RECT 67.285 30.395 67.575 30.440 ;
        RECT 70.030 30.380 70.350 30.440 ;
        RECT 80.610 30.380 80.930 30.640 ;
        RECT 89.825 30.580 90.115 30.625 ;
        RECT 90.730 30.580 91.050 30.640 ;
        RECT 89.825 30.440 91.050 30.580 ;
        RECT 89.825 30.395 90.115 30.440 ;
        RECT 90.730 30.380 91.050 30.440 ;
        RECT 13.380 29.760 92.040 30.240 ;
        RECT 19.430 29.560 19.750 29.620 ;
        RECT 17.220 29.420 19.750 29.560 ;
        RECT 17.220 29.220 17.360 29.420 ;
        RECT 19.430 29.360 19.750 29.420 ;
        RECT 24.030 29.560 24.350 29.620 ;
        RECT 26.345 29.560 26.635 29.605 ;
        RECT 24.030 29.420 26.635 29.560 ;
        RECT 24.030 29.360 24.350 29.420 ;
        RECT 26.345 29.375 26.635 29.420 ;
        RECT 27.250 29.560 27.570 29.620 ;
        RECT 47.950 29.560 48.270 29.620 ;
        RECT 64.510 29.560 64.830 29.620 ;
        RECT 66.365 29.560 66.655 29.605 ;
        RECT 69.570 29.560 69.890 29.620 ;
        RECT 27.250 29.420 48.270 29.560 ;
        RECT 27.250 29.360 27.570 29.420 ;
        RECT 16.760 29.080 17.360 29.220 ;
        RECT 20.320 29.220 20.610 29.265 ;
        RECT 21.730 29.220 22.050 29.280 ;
        RECT 20.320 29.080 22.050 29.220 ;
        RECT 16.760 28.925 16.900 29.080 ;
        RECT 20.320 29.035 20.610 29.080 ;
        RECT 21.730 29.020 22.050 29.080 ;
        RECT 16.685 28.695 16.975 28.925 ;
        RECT 17.130 28.680 17.450 28.940 ;
        RECT 17.590 28.680 17.910 28.940 ;
        RECT 18.525 28.880 18.815 28.925 ;
        RECT 19.980 28.880 20.580 28.895 ;
        RECT 25.410 28.880 25.730 28.940 ;
        RECT 27.265 28.880 27.555 28.925 ;
        RECT 18.525 28.755 25.730 28.880 ;
        RECT 18.525 28.740 20.120 28.755 ;
        RECT 20.440 28.740 25.730 28.755 ;
        RECT 18.525 28.695 18.815 28.740 ;
        RECT 25.410 28.680 25.730 28.740 ;
        RECT 25.960 28.740 27.555 28.880 ;
        RECT 18.050 28.540 18.370 28.600 ;
        RECT 18.985 28.540 19.275 28.585 ;
        RECT 18.050 28.400 19.275 28.540 ;
        RECT 18.050 28.340 18.370 28.400 ;
        RECT 18.985 28.355 19.275 28.400 ;
        RECT 19.865 28.540 20.155 28.585 ;
        RECT 21.055 28.540 21.345 28.585 ;
        RECT 23.575 28.540 23.865 28.585 ;
        RECT 19.865 28.400 23.865 28.540 ;
        RECT 19.865 28.355 20.155 28.400 ;
        RECT 21.055 28.355 21.345 28.400 ;
        RECT 23.575 28.355 23.865 28.400 ;
        RECT 19.470 28.200 19.760 28.245 ;
        RECT 21.570 28.200 21.860 28.245 ;
        RECT 23.140 28.200 23.430 28.245 ;
        RECT 19.470 28.060 23.430 28.200 ;
        RECT 19.470 28.015 19.760 28.060 ;
        RECT 21.570 28.015 21.860 28.060 ;
        RECT 23.140 28.015 23.430 28.060 ;
        RECT 15.290 27.660 15.610 27.920 ;
        RECT 22.650 27.860 22.970 27.920 ;
        RECT 25.960 27.905 26.100 28.740 ;
        RECT 27.265 28.695 27.555 28.740 ;
        RECT 28.170 28.680 28.490 28.940 ;
        RECT 30.485 28.695 30.775 28.925 ;
        RECT 30.945 28.695 31.235 28.925 ;
        RECT 30.560 28.200 30.700 28.695 ;
        RECT 31.020 28.540 31.160 28.695 ;
        RECT 31.390 28.680 31.710 28.940 ;
        RECT 32.400 28.925 32.540 29.420 ;
        RECT 47.950 29.360 48.270 29.420 ;
        RECT 50.800 29.420 64.280 29.560 ;
        RECT 38.765 29.220 39.055 29.265 ;
        RECT 34.240 29.080 39.055 29.220 ;
        RECT 32.325 28.695 32.615 28.925 ;
        RECT 33.245 28.880 33.535 28.925 ;
        RECT 33.690 28.880 34.010 28.940 ;
        RECT 34.240 28.925 34.380 29.080 ;
        RECT 38.765 29.035 39.055 29.080 ;
        RECT 41.970 29.220 42.290 29.280 ;
        RECT 50.800 29.220 50.940 29.420 ;
        RECT 58.530 29.220 58.850 29.280 ;
        RECT 41.970 29.080 50.940 29.220 ;
        RECT 51.260 29.080 58.850 29.220 ;
        RECT 41.970 29.020 42.290 29.080 ;
        RECT 33.245 28.740 34.010 28.880 ;
        RECT 33.245 28.695 33.535 28.740 ;
        RECT 33.690 28.680 34.010 28.740 ;
        RECT 34.165 28.695 34.455 28.925 ;
        RECT 34.610 28.680 34.930 28.940 ;
        RECT 35.085 28.880 35.375 28.925 ;
        RECT 35.530 28.880 35.850 28.940 ;
        RECT 35.085 28.740 35.850 28.880 ;
        RECT 35.085 28.695 35.375 28.740 ;
        RECT 35.530 28.680 35.850 28.740 ;
        RECT 36.910 28.680 37.230 28.940 ;
        RECT 37.845 28.880 38.135 28.925 ;
        RECT 42.890 28.880 43.210 28.940 ;
        RECT 43.810 28.925 44.130 28.940 ;
        RECT 51.260 28.925 51.400 29.080 ;
        RECT 58.530 29.020 58.850 29.080 ;
        RECT 52.550 28.925 52.870 28.940 ;
        RECT 37.845 28.740 43.210 28.880 ;
        RECT 37.845 28.695 38.135 28.740 ;
        RECT 42.890 28.680 43.210 28.740 ;
        RECT 43.780 28.695 44.130 28.925 ;
        RECT 51.185 28.695 51.475 28.925 ;
        RECT 52.520 28.695 52.870 28.925 ;
        RECT 43.810 28.680 44.130 28.695 ;
        RECT 52.550 28.680 52.870 28.695 ;
        RECT 53.930 28.880 54.250 28.940 ;
        RECT 60.460 28.925 60.600 29.420 ;
        RECT 62.685 29.220 62.975 29.265 ;
        RECT 61.380 29.080 62.975 29.220 ;
        RECT 64.140 29.220 64.280 29.420 ;
        RECT 64.510 29.420 66.655 29.560 ;
        RECT 64.510 29.360 64.830 29.420 ;
        RECT 66.365 29.375 66.655 29.420 ;
        RECT 67.360 29.420 69.890 29.560 ;
        RECT 67.360 29.220 67.500 29.420 ;
        RECT 69.570 29.360 69.890 29.420 ;
        RECT 72.790 29.360 73.110 29.620 ;
        RECT 79.690 29.560 80.010 29.620 ;
        RECT 82.465 29.560 82.755 29.605 ;
        RECT 79.690 29.420 84.520 29.560 ;
        RECT 79.690 29.360 80.010 29.420 ;
        RECT 82.465 29.375 82.755 29.420 ;
        RECT 64.140 29.080 67.500 29.220 ;
        RECT 53.930 28.740 56.460 28.880 ;
        RECT 53.930 28.680 54.250 28.740 ;
        RECT 34.700 28.540 34.840 28.680 ;
        RECT 56.320 28.600 56.460 28.740 ;
        RECT 60.385 28.695 60.675 28.925 ;
        RECT 60.830 28.680 61.150 28.940 ;
        RECT 61.380 28.925 61.520 29.080 ;
        RECT 62.685 29.035 62.975 29.080 ;
        RECT 67.730 29.020 68.050 29.280 ;
        RECT 71.870 29.220 72.190 29.280 ;
        RECT 71.040 29.080 72.190 29.220 ;
        RECT 61.305 28.695 61.595 28.925 ;
        RECT 62.225 28.695 62.515 28.925 ;
        RECT 63.130 28.880 63.450 28.940 ;
        RECT 63.605 28.880 63.895 28.925 ;
        RECT 63.130 28.740 63.895 28.880 ;
        RECT 42.430 28.540 42.750 28.600 ;
        RECT 31.020 28.400 34.840 28.540 ;
        RECT 35.620 28.400 42.750 28.540 ;
        RECT 35.620 28.260 35.760 28.400 ;
        RECT 42.430 28.340 42.750 28.400 ;
        RECT 43.325 28.540 43.615 28.585 ;
        RECT 44.515 28.540 44.805 28.585 ;
        RECT 47.035 28.540 47.325 28.585 ;
        RECT 43.325 28.400 47.325 28.540 ;
        RECT 43.325 28.355 43.615 28.400 ;
        RECT 44.515 28.355 44.805 28.400 ;
        RECT 47.035 28.355 47.325 28.400 ;
        RECT 52.065 28.540 52.355 28.585 ;
        RECT 53.255 28.540 53.545 28.585 ;
        RECT 55.775 28.540 56.065 28.585 ;
        RECT 52.065 28.400 56.065 28.540 ;
        RECT 52.065 28.355 52.355 28.400 ;
        RECT 53.255 28.355 53.545 28.400 ;
        RECT 55.775 28.355 56.065 28.400 ;
        RECT 56.230 28.540 56.550 28.600 ;
        RECT 62.300 28.540 62.440 28.695 ;
        RECT 63.130 28.680 63.450 28.740 ;
        RECT 63.605 28.695 63.895 28.740 ;
        RECT 64.050 28.880 64.370 28.940 ;
        RECT 64.525 28.880 64.815 28.925 ;
        RECT 64.050 28.740 64.815 28.880 ;
        RECT 56.230 28.400 62.440 28.540 ;
        RECT 63.680 28.540 63.820 28.695 ;
        RECT 64.050 28.680 64.370 28.740 ;
        RECT 64.525 28.695 64.815 28.740 ;
        RECT 67.270 28.680 67.590 28.940 ;
        RECT 68.190 28.680 68.510 28.940 ;
        RECT 69.125 28.880 69.415 28.925 ;
        RECT 68.740 28.740 69.415 28.880 ;
        RECT 68.740 28.540 68.880 28.740 ;
        RECT 69.125 28.695 69.415 28.740 ;
        RECT 69.585 28.695 69.875 28.925 ;
        RECT 70.030 28.880 70.350 28.940 ;
        RECT 71.040 28.925 71.180 29.080 ;
        RECT 71.870 29.020 72.190 29.080 ;
        RECT 73.250 29.220 73.570 29.280 ;
        RECT 83.370 29.220 83.690 29.280 ;
        RECT 84.380 29.265 84.520 29.420 ;
        RECT 73.250 29.080 83.690 29.220 ;
        RECT 73.250 29.020 73.570 29.080 ;
        RECT 75.640 28.925 75.780 29.080 ;
        RECT 83.370 29.020 83.690 29.080 ;
        RECT 84.305 29.220 84.595 29.265 ;
        RECT 86.130 29.220 86.450 29.280 ;
        RECT 84.305 29.080 86.450 29.220 ;
        RECT 84.305 29.035 84.595 29.080 ;
        RECT 86.130 29.020 86.450 29.080 ;
        RECT 70.505 28.880 70.795 28.925 ;
        RECT 70.030 28.740 70.795 28.880 ;
        RECT 69.660 28.540 69.800 28.695 ;
        RECT 70.030 28.680 70.350 28.740 ;
        RECT 70.505 28.695 70.795 28.740 ;
        RECT 70.965 28.695 71.255 28.925 ;
        RECT 71.425 28.695 71.715 28.925 ;
        RECT 75.565 28.695 75.855 28.925 ;
        RECT 76.900 28.880 77.190 28.925 ;
        RECT 78.310 28.880 78.630 28.940 ;
        RECT 76.900 28.740 78.630 28.880 ;
        RECT 76.900 28.695 77.190 28.740 ;
        RECT 63.680 28.400 68.880 28.540 ;
        RECT 69.200 28.400 69.800 28.540 ;
        RECT 56.230 28.340 56.550 28.400 ;
        RECT 30.560 28.060 31.620 28.200 ;
        RECT 25.885 27.860 26.175 27.905 ;
        RECT 22.650 27.720 26.175 27.860 ;
        RECT 22.650 27.660 22.970 27.720 ;
        RECT 25.885 27.675 26.175 27.720 ;
        RECT 29.105 27.860 29.395 27.905 ;
        RECT 30.930 27.860 31.250 27.920 ;
        RECT 29.105 27.720 31.250 27.860 ;
        RECT 31.480 27.860 31.620 28.060 ;
        RECT 35.530 28.000 35.850 28.260 ;
        RECT 37.370 28.200 37.690 28.260 ;
        RECT 36.080 28.060 37.690 28.200 ;
        RECT 36.080 27.860 36.220 28.060 ;
        RECT 37.370 28.000 37.690 28.060 ;
        RECT 42.930 28.200 43.220 28.245 ;
        RECT 45.030 28.200 45.320 28.245 ;
        RECT 46.600 28.200 46.890 28.245 ;
        RECT 42.930 28.060 46.890 28.200 ;
        RECT 42.930 28.015 43.220 28.060 ;
        RECT 45.030 28.015 45.320 28.060 ;
        RECT 46.600 28.015 46.890 28.060 ;
        RECT 51.670 28.200 51.960 28.245 ;
        RECT 53.770 28.200 54.060 28.245 ;
        RECT 55.340 28.200 55.630 28.245 ;
        RECT 51.670 28.060 55.630 28.200 ;
        RECT 51.670 28.015 51.960 28.060 ;
        RECT 53.770 28.015 54.060 28.060 ;
        RECT 55.340 28.015 55.630 28.060 ;
        RECT 59.005 28.200 59.295 28.245 ;
        RECT 59.910 28.200 60.230 28.260 ;
        RECT 59.005 28.060 60.230 28.200 ;
        RECT 59.005 28.015 59.295 28.060 ;
        RECT 59.910 28.000 60.230 28.060 ;
        RECT 31.480 27.720 36.220 27.860 ;
        RECT 29.105 27.675 29.395 27.720 ;
        RECT 30.930 27.660 31.250 27.720 ;
        RECT 36.450 27.660 36.770 27.920 ;
        RECT 45.650 27.860 45.970 27.920 ;
        RECT 49.345 27.860 49.635 27.905 ;
        RECT 45.650 27.720 49.635 27.860 ;
        RECT 45.650 27.660 45.970 27.720 ;
        RECT 49.345 27.675 49.635 27.720 ;
        RECT 55.770 27.860 56.090 27.920 ;
        RECT 58.085 27.860 58.375 27.905 ;
        RECT 55.770 27.720 58.375 27.860 ;
        RECT 62.300 27.860 62.440 28.400 ;
        RECT 62.670 28.200 62.990 28.260 ;
        RECT 67.270 28.200 67.590 28.260 ;
        RECT 62.670 28.060 67.590 28.200 ;
        RECT 62.670 28.000 62.990 28.060 ;
        RECT 67.270 28.000 67.590 28.060 ;
        RECT 69.200 27.860 69.340 28.400 ;
        RECT 69.570 28.200 69.890 28.260 ;
        RECT 71.500 28.200 71.640 28.695 ;
        RECT 78.310 28.680 78.630 28.740 ;
        RECT 78.770 28.880 79.090 28.940 ;
        RECT 82.450 28.880 82.770 28.940 ;
        RECT 83.845 28.880 84.135 28.925 ;
        RECT 78.770 28.740 81.300 28.880 ;
        RECT 78.770 28.680 79.090 28.740 ;
        RECT 81.160 28.600 81.300 28.740 ;
        RECT 82.450 28.740 84.135 28.880 ;
        RECT 82.450 28.680 82.770 28.740 ;
        RECT 83.845 28.695 84.135 28.740 ;
        RECT 84.765 28.695 85.055 28.925 ;
        RECT 76.445 28.540 76.735 28.585 ;
        RECT 77.635 28.540 77.925 28.585 ;
        RECT 80.155 28.540 80.445 28.585 ;
        RECT 76.445 28.400 80.445 28.540 ;
        RECT 76.445 28.355 76.735 28.400 ;
        RECT 77.635 28.355 77.925 28.400 ;
        RECT 80.155 28.355 80.445 28.400 ;
        RECT 81.070 28.540 81.390 28.600 ;
        RECT 84.840 28.540 84.980 28.695 ;
        RECT 85.670 28.680 85.990 28.940 ;
        RECT 81.070 28.400 84.980 28.540 ;
        RECT 81.070 28.340 81.390 28.400 ;
        RECT 69.570 28.060 71.640 28.200 ;
        RECT 76.050 28.200 76.340 28.245 ;
        RECT 78.150 28.200 78.440 28.245 ;
        RECT 79.720 28.200 80.010 28.245 ;
        RECT 76.050 28.060 80.010 28.200 ;
        RECT 69.570 28.000 69.890 28.060 ;
        RECT 76.050 28.015 76.340 28.060 ;
        RECT 78.150 28.015 78.440 28.060 ;
        RECT 79.720 28.015 80.010 28.060 ;
        RECT 81.530 27.860 81.850 27.920 ;
        RECT 62.300 27.720 81.850 27.860 ;
        RECT 55.770 27.660 56.090 27.720 ;
        RECT 58.085 27.675 58.375 27.720 ;
        RECT 81.530 27.660 81.850 27.720 ;
        RECT 82.910 27.660 83.230 27.920 ;
        RECT 13.380 27.040 92.040 27.520 ;
        RECT 18.510 26.840 18.830 26.900 ;
        RECT 21.745 26.840 22.035 26.885 ;
        RECT 18.510 26.700 22.035 26.840 ;
        RECT 18.510 26.640 18.830 26.700 ;
        RECT 21.745 26.655 22.035 26.700 ;
        RECT 15.330 26.500 15.620 26.545 ;
        RECT 17.430 26.500 17.720 26.545 ;
        RECT 19.000 26.500 19.290 26.545 ;
        RECT 15.330 26.360 19.290 26.500 ;
        RECT 15.330 26.315 15.620 26.360 ;
        RECT 17.430 26.315 17.720 26.360 ;
        RECT 19.000 26.315 19.290 26.360 ;
        RECT 15.725 26.160 16.015 26.205 ;
        RECT 16.915 26.160 17.205 26.205 ;
        RECT 19.435 26.160 19.725 26.205 ;
        RECT 15.725 26.020 19.725 26.160 ;
        RECT 15.725 25.975 16.015 26.020 ;
        RECT 16.915 25.975 17.205 26.020 ;
        RECT 19.435 25.975 19.725 26.020 ;
        RECT 14.845 25.820 15.135 25.865 ;
        RECT 18.050 25.820 18.370 25.880 ;
        RECT 14.845 25.680 18.370 25.820 ;
        RECT 21.820 25.820 21.960 26.655 ;
        RECT 24.950 26.640 25.270 26.900 ;
        RECT 27.710 26.840 28.030 26.900 ;
        RECT 42.445 26.840 42.735 26.885 ;
        RECT 42.890 26.840 43.210 26.900 ;
        RECT 27.710 26.700 42.200 26.840 ;
        RECT 27.710 26.640 28.030 26.700 ;
        RECT 28.670 26.500 28.960 26.545 ;
        RECT 30.770 26.500 31.060 26.545 ;
        RECT 32.340 26.500 32.630 26.545 ;
        RECT 28.670 26.360 32.630 26.500 ;
        RECT 28.670 26.315 28.960 26.360 ;
        RECT 30.770 26.315 31.060 26.360 ;
        RECT 32.340 26.315 32.630 26.360 ;
        RECT 36.030 26.500 36.320 26.545 ;
        RECT 38.130 26.500 38.420 26.545 ;
        RECT 39.700 26.500 39.990 26.545 ;
        RECT 36.030 26.360 39.990 26.500 ;
        RECT 42.060 26.500 42.200 26.700 ;
        RECT 42.445 26.700 43.210 26.840 ;
        RECT 42.445 26.655 42.735 26.700 ;
        RECT 42.890 26.640 43.210 26.700 ;
        RECT 43.810 26.640 44.130 26.900 ;
        RECT 46.660 26.700 70.030 26.840 ;
        RECT 46.660 26.500 46.800 26.700 ;
        RECT 42.060 26.360 46.800 26.500 ;
        RECT 36.030 26.315 36.320 26.360 ;
        RECT 38.130 26.315 38.420 26.360 ;
        RECT 39.700 26.315 39.990 26.360 ;
        RECT 47.030 26.300 47.350 26.560 ;
        RECT 52.550 26.300 52.870 26.560 ;
        RECT 69.890 26.500 70.030 26.700 ;
        RECT 78.310 26.640 78.630 26.900 ;
        RECT 82.910 26.500 83.230 26.560 ;
        RECT 69.890 26.360 83.230 26.500 ;
        RECT 82.910 26.300 83.230 26.360 ;
        RECT 83.870 26.500 84.160 26.545 ;
        RECT 85.970 26.500 86.260 26.545 ;
        RECT 87.540 26.500 87.830 26.545 ;
        RECT 83.870 26.360 87.830 26.500 ;
        RECT 83.870 26.315 84.160 26.360 ;
        RECT 85.970 26.315 86.260 26.360 ;
        RECT 87.540 26.315 87.830 26.360 ;
        RECT 29.065 26.160 29.355 26.205 ;
        RECT 30.255 26.160 30.545 26.205 ;
        RECT 32.775 26.160 33.065 26.205 ;
        RECT 29.065 26.020 33.065 26.160 ;
        RECT 29.065 25.975 29.355 26.020 ;
        RECT 30.255 25.975 30.545 26.020 ;
        RECT 32.775 25.975 33.065 26.020 ;
        RECT 36.425 26.160 36.715 26.205 ;
        RECT 37.615 26.160 37.905 26.205 ;
        RECT 40.135 26.160 40.425 26.205 ;
        RECT 47.120 26.160 47.260 26.300 ;
        RECT 48.870 26.160 49.190 26.220 ;
        RECT 74.170 26.160 74.490 26.220 ;
        RECT 78.310 26.160 78.630 26.220 ;
        RECT 81.070 26.160 81.390 26.220 ;
        RECT 83.370 26.160 83.690 26.220 ;
        RECT 36.425 26.020 40.425 26.160 ;
        RECT 36.425 25.975 36.715 26.020 ;
        RECT 37.615 25.975 37.905 26.020 ;
        RECT 40.135 25.975 40.425 26.020 ;
        RECT 45.740 26.020 78.080 26.160 ;
        RECT 22.205 25.820 22.495 25.865 ;
        RECT 21.820 25.680 22.495 25.820 ;
        RECT 14.845 25.635 15.135 25.680 ;
        RECT 18.050 25.620 18.370 25.680 ;
        RECT 22.205 25.635 22.495 25.680 ;
        RECT 22.650 25.820 22.970 25.880 ;
        RECT 23.585 25.820 23.875 25.865 ;
        RECT 22.650 25.680 23.875 25.820 ;
        RECT 22.650 25.620 22.970 25.680 ;
        RECT 23.585 25.635 23.875 25.680 ;
        RECT 24.045 25.820 24.335 25.865 ;
        RECT 25.410 25.820 25.730 25.880 ;
        RECT 24.045 25.680 25.730 25.820 ;
        RECT 24.045 25.635 24.335 25.680 ;
        RECT 25.410 25.620 25.730 25.680 ;
        RECT 28.170 25.620 28.490 25.880 ;
        RECT 29.520 25.820 29.810 25.865 ;
        RECT 30.930 25.820 31.250 25.880 ;
        RECT 29.520 25.680 31.250 25.820 ;
        RECT 29.520 25.635 29.810 25.680 ;
        RECT 30.930 25.620 31.250 25.680 ;
        RECT 35.530 25.620 35.850 25.880 ;
        RECT 45.740 25.865 45.880 26.020 ;
        RECT 48.870 25.960 49.190 26.020 ;
        RECT 36.880 25.635 37.170 25.865 ;
        RECT 45.205 25.635 45.495 25.865 ;
        RECT 45.665 25.635 45.955 25.865 ;
        RECT 15.290 25.480 15.610 25.540 ;
        RECT 16.070 25.480 16.360 25.525 ;
        RECT 23.125 25.480 23.415 25.525 ;
        RECT 15.290 25.340 16.360 25.480 ;
        RECT 15.290 25.280 15.610 25.340 ;
        RECT 16.070 25.295 16.360 25.340 ;
        RECT 22.280 25.340 23.415 25.480 ;
        RECT 22.280 25.200 22.420 25.340 ;
        RECT 23.125 25.295 23.415 25.340 ;
        RECT 36.450 25.480 36.770 25.540 ;
        RECT 37.000 25.480 37.140 25.635 ;
        RECT 36.450 25.340 37.140 25.480 ;
        RECT 37.370 25.480 37.690 25.540 ;
        RECT 41.970 25.480 42.290 25.540 ;
        RECT 45.280 25.480 45.420 25.635 ;
        RECT 46.110 25.620 46.430 25.880 ;
        RECT 47.045 25.820 47.335 25.865 ;
        RECT 47.950 25.820 48.270 25.880 ;
        RECT 53.930 25.820 54.250 25.880 ;
        RECT 54.480 25.865 54.620 26.020 ;
        RECT 74.170 25.960 74.490 26.020 ;
        RECT 47.045 25.680 48.270 25.820 ;
        RECT 47.045 25.635 47.335 25.680 ;
        RECT 47.950 25.620 48.270 25.680 ;
        RECT 50.340 25.680 54.250 25.820 ;
        RECT 37.370 25.340 45.420 25.480 ;
        RECT 36.450 25.280 36.770 25.340 ;
        RECT 37.370 25.280 37.690 25.340 ;
        RECT 41.970 25.280 42.290 25.340 ;
        RECT 49.790 25.280 50.110 25.540 ;
        RECT 22.190 24.940 22.510 25.200 ;
        RECT 30.930 25.140 31.250 25.200 ;
        RECT 35.085 25.140 35.375 25.185 ;
        RECT 30.930 25.000 35.375 25.140 ;
        RECT 30.930 24.940 31.250 25.000 ;
        RECT 35.085 24.955 35.375 25.000 ;
        RECT 35.990 25.140 36.310 25.200 ;
        RECT 50.340 25.140 50.480 25.680 ;
        RECT 53.930 25.620 54.250 25.680 ;
        RECT 54.405 25.635 54.695 25.865 ;
        RECT 54.865 25.635 55.155 25.865 ;
        RECT 55.785 25.635 56.075 25.865 ;
        RECT 59.465 25.820 59.755 25.865 ;
        RECT 68.650 25.820 68.970 25.880 ;
        RECT 75.565 25.820 75.855 25.865 ;
        RECT 77.390 25.820 77.710 25.880 ;
        RECT 59.465 25.680 68.970 25.820 ;
        RECT 59.465 25.635 59.755 25.680 ;
        RECT 50.725 25.295 51.015 25.525 ;
        RECT 51.645 25.480 51.935 25.525 ;
        RECT 54.940 25.480 55.080 25.635 ;
        RECT 51.645 25.340 55.080 25.480 ;
        RECT 51.645 25.295 51.935 25.340 ;
        RECT 35.990 25.000 50.480 25.140 ;
        RECT 50.800 25.140 50.940 25.295 ;
        RECT 55.860 25.200 56.000 25.635 ;
        RECT 68.650 25.620 68.970 25.680 ;
        RECT 69.890 25.680 77.710 25.820 ;
        RECT 77.940 25.820 78.080 26.020 ;
        RECT 78.310 26.020 80.380 26.160 ;
        RECT 78.310 25.960 78.630 26.020 ;
        RECT 79.230 25.820 79.550 25.880 ;
        RECT 77.940 25.680 79.550 25.820 ;
        RECT 56.230 25.480 56.550 25.540 ;
        RECT 69.890 25.480 70.030 25.680 ;
        RECT 75.565 25.635 75.855 25.680 ;
        RECT 77.390 25.620 77.710 25.680 ;
        RECT 79.230 25.620 79.550 25.680 ;
        RECT 79.690 25.620 80.010 25.880 ;
        RECT 80.240 25.865 80.380 26.020 ;
        RECT 81.070 26.020 83.690 26.160 ;
        RECT 81.070 25.960 81.390 26.020 ;
        RECT 83.370 25.960 83.690 26.020 ;
        RECT 84.265 26.160 84.555 26.205 ;
        RECT 85.455 26.160 85.745 26.205 ;
        RECT 87.975 26.160 88.265 26.205 ;
        RECT 84.265 26.020 88.265 26.160 ;
        RECT 84.265 25.975 84.555 26.020 ;
        RECT 85.455 25.975 85.745 26.020 ;
        RECT 87.975 25.975 88.265 26.020 ;
        RECT 80.165 25.635 80.455 25.865 ;
        RECT 80.610 25.620 80.930 25.880 ;
        RECT 81.530 25.620 81.850 25.880 ;
        RECT 56.230 25.340 70.030 25.480 ;
        RECT 76.485 25.480 76.775 25.525 ;
        RECT 83.370 25.480 83.690 25.540 ;
        RECT 84.610 25.480 84.900 25.525 ;
        RECT 76.485 25.340 83.140 25.480 ;
        RECT 56.230 25.280 56.550 25.340 ;
        RECT 76.485 25.295 76.775 25.340 ;
        RECT 52.090 25.140 52.410 25.200 ;
        RECT 55.310 25.140 55.630 25.200 ;
        RECT 50.800 25.000 55.630 25.140 ;
        RECT 35.990 24.940 36.310 25.000 ;
        RECT 52.090 24.940 52.410 25.000 ;
        RECT 55.310 24.940 55.630 25.000 ;
        RECT 55.770 25.140 56.090 25.200 ;
        RECT 58.545 25.140 58.835 25.185 ;
        RECT 55.770 25.000 58.835 25.140 ;
        RECT 55.770 24.940 56.090 25.000 ;
        RECT 58.545 24.955 58.835 25.000 ;
        RECT 77.405 25.140 77.695 25.185 ;
        RECT 80.610 25.140 80.930 25.200 ;
        RECT 77.405 25.000 80.930 25.140 ;
        RECT 83.000 25.140 83.140 25.340 ;
        RECT 83.370 25.340 84.900 25.480 ;
        RECT 83.370 25.280 83.690 25.340 ;
        RECT 84.610 25.295 84.900 25.340 ;
        RECT 85.670 25.140 85.990 25.200 ;
        RECT 90.270 25.140 90.590 25.200 ;
        RECT 83.000 25.000 90.590 25.140 ;
        RECT 77.405 24.955 77.695 25.000 ;
        RECT 80.610 24.940 80.930 25.000 ;
        RECT 85.670 24.940 85.990 25.000 ;
        RECT 90.270 24.940 90.590 25.000 ;
        RECT 13.380 24.320 92.040 24.800 ;
        RECT 30.485 24.120 30.775 24.165 ;
        RECT 31.390 24.120 31.710 24.180 ;
        RECT 30.485 23.980 31.710 24.120 ;
        RECT 30.485 23.935 30.775 23.980 ;
        RECT 31.390 23.920 31.710 23.980 ;
        RECT 43.810 24.120 44.130 24.180 ;
        RECT 49.790 24.120 50.110 24.180 ;
        RECT 56.230 24.120 56.550 24.180 ;
        RECT 43.810 23.980 47.720 24.120 ;
        RECT 43.810 23.920 44.130 23.980 ;
        RECT 22.190 23.780 22.510 23.840 ;
        RECT 23.585 23.780 23.875 23.825 ;
        RECT 22.190 23.640 23.875 23.780 ;
        RECT 22.190 23.580 22.510 23.640 ;
        RECT 23.585 23.595 23.875 23.640 ;
        RECT 27.710 23.780 28.030 23.840 ;
        RECT 28.645 23.780 28.935 23.825 ;
        RECT 27.710 23.640 28.935 23.780 ;
        RECT 27.710 23.580 28.030 23.640 ;
        RECT 28.645 23.595 28.935 23.640 ;
        RECT 29.565 23.780 29.855 23.825 ;
        RECT 30.930 23.780 31.250 23.840 ;
        RECT 29.565 23.640 31.250 23.780 ;
        RECT 29.565 23.595 29.855 23.640 ;
        RECT 30.930 23.580 31.250 23.640 ;
        RECT 40.590 23.780 40.910 23.840 ;
        RECT 42.445 23.780 42.735 23.825 ;
        RECT 45.650 23.780 45.970 23.840 ;
        RECT 40.590 23.640 42.735 23.780 ;
        RECT 40.590 23.580 40.910 23.640 ;
        RECT 42.445 23.595 42.735 23.640 ;
        RECT 42.980 23.640 45.970 23.780 ;
        RECT 16.225 23.255 16.515 23.485 ;
        RECT 18.510 23.440 18.830 23.500 ;
        RECT 19.445 23.440 19.735 23.485 ;
        RECT 18.510 23.300 19.735 23.440 ;
        RECT 16.300 22.760 16.440 23.255 ;
        RECT 18.510 23.240 18.830 23.300 ;
        RECT 19.445 23.255 19.735 23.300 ;
        RECT 21.285 23.440 21.575 23.485 ;
        RECT 21.730 23.440 22.050 23.500 ;
        RECT 22.665 23.440 22.955 23.485 ;
        RECT 21.285 23.300 22.955 23.440 ;
        RECT 21.285 23.255 21.575 23.300 ;
        RECT 21.730 23.240 22.050 23.300 ;
        RECT 22.665 23.255 22.955 23.300 ;
        RECT 24.045 23.255 24.335 23.485 ;
        RECT 24.505 23.440 24.795 23.485 ;
        RECT 25.410 23.440 25.730 23.500 ;
        RECT 24.505 23.300 25.730 23.440 ;
        RECT 24.505 23.255 24.795 23.300 ;
        RECT 24.120 23.100 24.260 23.255 ;
        RECT 25.410 23.240 25.730 23.300 ;
        RECT 25.885 23.440 26.175 23.485 ;
        RECT 26.330 23.440 26.650 23.500 ;
        RECT 25.885 23.300 26.650 23.440 ;
        RECT 31.020 23.440 31.160 23.580 ;
        RECT 42.980 23.485 43.120 23.640 ;
        RECT 45.650 23.580 45.970 23.640 ;
        RECT 47.030 23.580 47.350 23.840 ;
        RECT 47.580 23.780 47.720 23.980 ;
        RECT 49.790 23.980 56.550 24.120 ;
        RECT 49.790 23.920 50.110 23.980 ;
        RECT 56.230 23.920 56.550 23.980 ;
        RECT 65.890 24.120 66.210 24.180 ;
        RECT 71.870 24.120 72.190 24.180 ;
        RECT 78.310 24.120 78.630 24.180 ;
        RECT 65.890 23.980 68.420 24.120 ;
        RECT 65.890 23.920 66.210 23.980 ;
        RECT 51.630 23.780 51.950 23.840 ;
        RECT 47.580 23.640 51.950 23.780 ;
        RECT 41.525 23.440 41.815 23.485 ;
        RECT 31.020 23.300 41.815 23.440 ;
        RECT 25.885 23.255 26.175 23.300 ;
        RECT 25.960 23.100 26.100 23.255 ;
        RECT 26.330 23.240 26.650 23.300 ;
        RECT 41.525 23.255 41.815 23.300 ;
        RECT 42.905 23.255 43.195 23.485 ;
        RECT 43.365 23.440 43.655 23.485 ;
        RECT 43.810 23.440 44.130 23.500 ;
        RECT 48.040 23.485 48.180 23.640 ;
        RECT 51.630 23.580 51.950 23.640 ;
        RECT 55.770 23.780 56.090 23.840 ;
        RECT 63.605 23.780 63.895 23.825 ;
        RECT 68.280 23.780 68.420 23.980 ;
        RECT 70.580 23.980 78.630 24.120 ;
        RECT 55.770 23.640 62.440 23.780 ;
        RECT 55.770 23.580 56.090 23.640 ;
        RECT 43.365 23.300 44.130 23.440 ;
        RECT 43.365 23.255 43.655 23.300 ;
        RECT 43.810 23.240 44.130 23.300 ;
        RECT 46.125 23.255 46.415 23.485 ;
        RECT 47.505 23.255 47.795 23.485 ;
        RECT 47.965 23.255 48.255 23.485 ;
        RECT 58.070 23.440 58.390 23.500 ;
        RECT 60.385 23.440 60.675 23.485 ;
        RECT 58.070 23.300 60.675 23.440 ;
        RECT 24.120 22.960 26.100 23.100 ;
        RECT 41.970 23.100 42.290 23.160 ;
        RECT 46.200 23.100 46.340 23.255 ;
        RECT 41.970 22.960 46.340 23.100 ;
        RECT 47.580 23.100 47.720 23.255 ;
        RECT 58.070 23.240 58.390 23.300 ;
        RECT 60.385 23.255 60.675 23.300 ;
        RECT 60.830 23.240 61.150 23.500 ;
        RECT 62.300 23.485 62.440 23.640 ;
        RECT 63.605 23.640 67.960 23.780 ;
        RECT 68.280 23.640 68.880 23.780 ;
        RECT 63.605 23.595 63.895 23.640 ;
        RECT 67.820 23.500 67.960 23.640 ;
        RECT 61.305 23.255 61.595 23.485 ;
        RECT 62.225 23.255 62.515 23.485 ;
        RECT 64.050 23.440 64.370 23.500 ;
        RECT 64.525 23.440 64.815 23.485 ;
        RECT 64.050 23.300 64.815 23.440 ;
        RECT 49.330 23.100 49.650 23.160 ;
        RECT 47.580 22.960 49.650 23.100 ;
        RECT 41.970 22.900 42.290 22.960 ;
        RECT 49.330 22.900 49.650 22.960 ;
        RECT 56.690 23.100 57.010 23.160 ;
        RECT 60.920 23.100 61.060 23.240 ;
        RECT 56.690 22.960 61.060 23.100 ;
        RECT 61.380 23.100 61.520 23.255 ;
        RECT 64.050 23.240 64.370 23.300 ;
        RECT 64.525 23.255 64.815 23.300 ;
        RECT 66.350 23.240 66.670 23.500 ;
        RECT 66.825 23.255 67.115 23.485 ;
        RECT 62.685 23.100 62.975 23.145 ;
        RECT 65.890 23.100 66.210 23.160 ;
        RECT 61.380 22.960 62.975 23.100 ;
        RECT 56.690 22.900 57.010 22.960 ;
        RECT 62.685 22.915 62.975 22.960 ;
        RECT 63.220 22.960 66.210 23.100 ;
        RECT 66.900 23.100 67.040 23.255 ;
        RECT 67.270 23.240 67.590 23.500 ;
        RECT 67.730 23.440 68.050 23.500 ;
        RECT 68.205 23.440 68.495 23.485 ;
        RECT 67.730 23.300 68.495 23.440 ;
        RECT 68.740 23.440 68.880 23.640 ;
        RECT 70.580 23.485 70.720 23.980 ;
        RECT 71.870 23.920 72.190 23.980 ;
        RECT 78.310 23.920 78.630 23.980 ;
        RECT 79.230 23.920 79.550 24.180 ;
        RECT 79.690 24.120 80.010 24.180 ;
        RECT 79.690 23.980 82.220 24.120 ;
        RECT 79.690 23.920 80.010 23.980 ;
        RECT 74.185 23.780 74.475 23.825 ;
        RECT 75.090 23.780 75.410 23.840 ;
        RECT 74.185 23.640 75.410 23.780 ;
        RECT 74.185 23.595 74.475 23.640 ;
        RECT 75.090 23.580 75.410 23.640 ;
        RECT 75.550 23.780 75.870 23.840 ;
        RECT 79.320 23.780 79.460 23.920 ;
        RECT 82.080 23.780 82.220 23.980 ;
        RECT 82.450 23.780 82.770 23.840 ;
        RECT 75.550 23.640 78.080 23.780 ;
        RECT 79.320 23.640 81.760 23.780 ;
        RECT 75.550 23.580 75.870 23.640 ;
        RECT 70.045 23.440 70.335 23.485 ;
        RECT 68.740 23.300 70.335 23.440 ;
        RECT 67.730 23.240 68.050 23.300 ;
        RECT 68.205 23.255 68.495 23.300 ;
        RECT 70.045 23.255 70.335 23.300 ;
        RECT 70.505 23.255 70.795 23.485 ;
        RECT 70.965 23.255 71.255 23.485 ;
        RECT 71.885 23.440 72.175 23.485 ;
        RECT 71.885 23.300 73.020 23.440 ;
        RECT 71.885 23.255 72.175 23.300 ;
        RECT 69.110 23.100 69.430 23.160 ;
        RECT 66.900 22.960 69.430 23.100 ;
        RECT 71.040 23.100 71.180 23.255 ;
        RECT 72.345 23.100 72.635 23.145 ;
        RECT 71.040 22.960 72.635 23.100 ;
        RECT 72.880 23.100 73.020 23.300 ;
        RECT 73.250 23.240 73.570 23.500 ;
        RECT 76.930 23.440 77.250 23.500 ;
        RECT 77.940 23.485 78.080 23.640 ;
        RECT 73.800 23.300 77.250 23.440 ;
        RECT 73.800 23.100 73.940 23.300 ;
        RECT 76.930 23.240 77.250 23.300 ;
        RECT 77.865 23.255 78.155 23.485 ;
        RECT 78.325 23.255 78.615 23.485 ;
        RECT 72.880 22.960 73.940 23.100 ;
        RECT 78.400 23.100 78.540 23.255 ;
        RECT 78.770 23.240 79.090 23.500 ;
        RECT 79.230 23.440 79.550 23.500 ;
        RECT 79.705 23.440 79.995 23.485 ;
        RECT 79.230 23.300 79.995 23.440 ;
        RECT 79.230 23.240 79.550 23.300 ;
        RECT 79.705 23.255 79.995 23.300 ;
        RECT 80.150 23.240 80.470 23.500 ;
        RECT 80.610 23.440 80.930 23.500 ;
        RECT 81.620 23.485 81.760 23.640 ;
        RECT 82.080 23.640 82.770 23.780 ;
        RECT 82.080 23.485 82.220 23.640 ;
        RECT 82.450 23.580 82.770 23.640 ;
        RECT 81.085 23.440 81.375 23.485 ;
        RECT 80.610 23.300 81.375 23.440 ;
        RECT 80.610 23.240 80.930 23.300 ;
        RECT 81.085 23.255 81.375 23.300 ;
        RECT 81.545 23.255 81.835 23.485 ;
        RECT 82.005 23.255 82.295 23.485 ;
        RECT 85.225 23.440 85.515 23.485 ;
        RECT 85.670 23.440 85.990 23.500 ;
        RECT 82.495 23.300 85.990 23.440 ;
        RECT 82.495 23.100 82.635 23.300 ;
        RECT 85.225 23.255 85.515 23.300 ;
        RECT 85.670 23.240 85.990 23.300 ;
        RECT 87.050 23.240 87.370 23.500 ;
        RECT 90.270 23.240 90.590 23.500 ;
        RECT 78.400 22.960 82.635 23.100 ;
        RECT 23.570 22.760 23.890 22.820 ;
        RECT 16.300 22.620 23.890 22.760 ;
        RECT 23.570 22.560 23.890 22.620 ;
        RECT 24.490 22.760 24.810 22.820 ;
        RECT 26.805 22.760 27.095 22.805 ;
        RECT 24.490 22.620 27.095 22.760 ;
        RECT 24.490 22.560 24.810 22.620 ;
        RECT 26.805 22.575 27.095 22.620 ;
        RECT 44.270 22.560 44.590 22.820 ;
        RECT 48.885 22.760 49.175 22.805 ;
        RECT 50.250 22.760 50.570 22.820 ;
        RECT 48.885 22.620 50.570 22.760 ;
        RECT 48.885 22.575 49.175 22.620 ;
        RECT 50.250 22.560 50.570 22.620 ;
        RECT 56.230 22.760 56.550 22.820 ;
        RECT 63.220 22.760 63.360 22.960 ;
        RECT 65.890 22.900 66.210 22.960 ;
        RECT 69.110 22.900 69.430 22.960 ;
        RECT 72.345 22.915 72.635 22.960 ;
        RECT 83.370 22.900 83.690 23.160 ;
        RECT 94.870 23.100 95.190 23.160 ;
        RECT 86.220 22.960 95.190 23.100 ;
        RECT 56.230 22.620 63.360 22.760 ;
        RECT 56.230 22.560 56.550 22.620 ;
        RECT 65.430 22.560 65.750 22.820 ;
        RECT 70.490 22.760 70.810 22.820 ;
        RECT 86.220 22.805 86.360 22.960 ;
        RECT 94.870 22.900 95.190 22.960 ;
        RECT 76.945 22.760 77.235 22.805 ;
        RECT 70.490 22.620 77.235 22.760 ;
        RECT 70.490 22.560 70.810 22.620 ;
        RECT 76.945 22.575 77.235 22.620 ;
        RECT 86.145 22.575 86.435 22.805 ;
        RECT 87.985 22.760 88.275 22.805 ;
        RECT 91.650 22.760 91.970 22.820 ;
        RECT 87.985 22.620 91.970 22.760 ;
        RECT 87.985 22.575 88.275 22.620 ;
        RECT 91.650 22.560 91.970 22.620 ;
        RECT 14.830 22.420 15.150 22.480 ;
        RECT 15.305 22.420 15.595 22.465 ;
        RECT 14.830 22.280 15.595 22.420 ;
        RECT 14.830 22.220 15.150 22.280 ;
        RECT 15.305 22.235 15.595 22.280 ;
        RECT 18.510 22.220 18.830 22.480 ;
        RECT 19.430 22.420 19.750 22.480 ;
        RECT 20.365 22.420 20.655 22.465 ;
        RECT 19.430 22.280 20.655 22.420 ;
        RECT 19.430 22.220 19.750 22.280 ;
        RECT 20.365 22.235 20.655 22.280 ;
        RECT 24.950 22.420 25.270 22.480 ;
        RECT 25.425 22.420 25.715 22.465 ;
        RECT 24.950 22.280 25.715 22.420 ;
        RECT 24.950 22.220 25.270 22.280 ;
        RECT 25.425 22.235 25.715 22.280 ;
        RECT 58.990 22.220 59.310 22.480 ;
        RECT 67.270 22.420 67.590 22.480 ;
        RECT 68.665 22.420 68.955 22.465 ;
        RECT 67.270 22.280 68.955 22.420 ;
        RECT 67.270 22.220 67.590 22.280 ;
        RECT 68.665 22.235 68.955 22.280 ;
        RECT 78.310 22.420 78.630 22.480 ;
        RECT 80.150 22.420 80.470 22.480 ;
        RECT 78.310 22.280 80.470 22.420 ;
        RECT 78.310 22.220 78.630 22.280 ;
        RECT 80.150 22.220 80.470 22.280 ;
        RECT 88.430 22.420 88.750 22.480 ;
        RECT 89.365 22.420 89.655 22.465 ;
        RECT 88.430 22.280 89.655 22.420 ;
        RECT 88.430 22.220 88.750 22.280 ;
        RECT 89.365 22.235 89.655 22.280 ;
        RECT 13.380 21.600 92.040 22.080 ;
        RECT 25.870 21.400 26.190 21.460 ;
        RECT 41.525 21.400 41.815 21.445 ;
        RECT 41.970 21.400 42.290 21.460 ;
        RECT 25.870 21.260 41.280 21.400 ;
        RECT 25.870 21.200 26.190 21.260 ;
        RECT 23.110 21.060 23.430 21.120 ;
        RECT 35.110 21.060 35.400 21.105 ;
        RECT 37.210 21.060 37.500 21.105 ;
        RECT 38.780 21.060 39.070 21.105 ;
        RECT 23.110 20.920 23.800 21.060 ;
        RECT 23.110 20.860 23.430 20.920 ;
        RECT 19.890 20.720 20.210 20.780 ;
        RECT 23.660 20.720 23.800 20.920 ;
        RECT 35.110 20.920 39.070 21.060 ;
        RECT 35.110 20.875 35.400 20.920 ;
        RECT 37.210 20.875 37.500 20.920 ;
        RECT 38.780 20.875 39.070 20.920 ;
        RECT 35.505 20.720 35.795 20.765 ;
        RECT 36.695 20.720 36.985 20.765 ;
        RECT 39.215 20.720 39.505 20.765 ;
        RECT 16.760 20.580 23.340 20.720 ;
        RECT 16.760 20.425 16.900 20.580 ;
        RECT 19.890 20.520 20.210 20.580 ;
        RECT 16.685 20.195 16.975 20.425 ;
        RECT 17.130 20.180 17.450 20.440 ;
        RECT 17.590 20.180 17.910 20.440 ;
        RECT 18.525 20.195 18.815 20.425 ;
        RECT 21.285 20.380 21.575 20.425 ;
        RECT 22.650 20.380 22.970 20.440 ;
        RECT 23.200 20.425 23.340 20.580 ;
        RECT 23.660 20.580 32.540 20.720 ;
        RECT 23.660 20.425 23.800 20.580 ;
        RECT 21.285 20.240 22.970 20.380 ;
        RECT 21.285 20.195 21.575 20.240 ;
        RECT 18.600 20.040 18.740 20.195 ;
        RECT 22.650 20.180 22.970 20.240 ;
        RECT 23.125 20.195 23.415 20.425 ;
        RECT 23.585 20.195 23.875 20.425 ;
        RECT 24.030 20.180 24.350 20.440 ;
        RECT 24.965 20.380 25.255 20.425 ;
        RECT 27.250 20.380 27.570 20.440 ;
        RECT 28.720 20.425 28.860 20.580 ;
        RECT 24.965 20.240 27.570 20.380 ;
        RECT 24.965 20.195 25.255 20.240 ;
        RECT 25.040 20.040 25.180 20.195 ;
        RECT 27.250 20.180 27.570 20.240 ;
        RECT 28.185 20.195 28.475 20.425 ;
        RECT 28.645 20.195 28.935 20.425 ;
        RECT 18.600 19.900 25.180 20.040 ;
        RECT 15.290 19.500 15.610 19.760 ;
        RECT 20.350 19.500 20.670 19.760 ;
        RECT 20.810 19.700 21.130 19.760 ;
        RECT 21.745 19.700 22.035 19.745 ;
        RECT 20.810 19.560 22.035 19.700 ;
        RECT 28.260 19.700 28.400 20.195 ;
        RECT 29.090 20.180 29.410 20.440 ;
        RECT 30.945 20.195 31.235 20.425 ;
        RECT 31.020 20.040 31.160 20.195 ;
        RECT 31.850 20.180 32.170 20.440 ;
        RECT 32.400 20.425 32.540 20.580 ;
        RECT 35.505 20.580 39.505 20.720 ;
        RECT 41.140 20.720 41.280 21.260 ;
        RECT 41.525 21.260 42.290 21.400 ;
        RECT 41.525 21.215 41.815 21.260 ;
        RECT 41.970 21.200 42.290 21.260 ;
        RECT 44.270 21.400 44.590 21.460 ;
        RECT 58.070 21.400 58.390 21.460 ;
        RECT 69.570 21.400 69.890 21.460 ;
        RECT 44.270 21.260 58.390 21.400 ;
        RECT 44.270 21.200 44.590 21.260 ;
        RECT 58.070 21.200 58.390 21.260 ;
        RECT 58.620 21.260 69.890 21.400 ;
        RECT 58.620 21.060 58.760 21.260 ;
        RECT 69.570 21.200 69.890 21.260 ;
        RECT 72.805 21.400 73.095 21.445 ;
        RECT 73.250 21.400 73.570 21.460 ;
        RECT 72.805 21.260 73.570 21.400 ;
        RECT 72.805 21.215 73.095 21.260 ;
        RECT 73.250 21.200 73.570 21.260 ;
        RECT 74.630 21.400 74.950 21.460 ;
        RECT 74.630 21.260 84.060 21.400 ;
        RECT 74.630 21.200 74.950 21.260 ;
        RECT 44.360 20.920 58.760 21.060 ;
        RECT 59.030 21.060 59.320 21.105 ;
        RECT 61.130 21.060 61.420 21.105 ;
        RECT 62.700 21.060 62.990 21.105 ;
        RECT 59.030 20.920 62.990 21.060 ;
        RECT 44.360 20.720 44.500 20.920 ;
        RECT 59.030 20.875 59.320 20.920 ;
        RECT 61.130 20.875 61.420 20.920 ;
        RECT 62.700 20.875 62.990 20.920 ;
        RECT 66.390 21.060 66.680 21.105 ;
        RECT 68.490 21.060 68.780 21.105 ;
        RECT 70.060 21.060 70.350 21.105 ;
        RECT 66.390 20.920 70.350 21.060 ;
        RECT 66.390 20.875 66.680 20.920 ;
        RECT 68.490 20.875 68.780 20.920 ;
        RECT 70.060 20.875 70.350 20.920 ;
        RECT 79.690 20.860 80.010 21.120 ;
        RECT 83.920 21.060 84.060 21.260 ;
        RECT 85.210 21.060 85.530 21.120 ;
        RECT 88.905 21.060 89.195 21.105 ;
        RECT 83.920 20.920 84.520 21.060 ;
        RECT 48.870 20.720 49.190 20.780 ;
        RECT 59.425 20.720 59.715 20.765 ;
        RECT 60.615 20.720 60.905 20.765 ;
        RECT 63.135 20.720 63.425 20.765 ;
        RECT 41.140 20.580 44.500 20.720 ;
        RECT 44.820 20.580 50.480 20.720 ;
        RECT 35.505 20.535 35.795 20.580 ;
        RECT 36.695 20.535 36.985 20.580 ;
        RECT 39.215 20.535 39.505 20.580 ;
        RECT 32.325 20.195 32.615 20.425 ;
        RECT 32.770 20.180 33.090 20.440 ;
        RECT 34.625 20.380 34.915 20.425 ;
        RECT 35.070 20.380 35.390 20.440 ;
        RECT 34.625 20.240 35.390 20.380 ;
        RECT 34.625 20.195 34.915 20.240 ;
        RECT 35.070 20.180 35.390 20.240 ;
        RECT 44.270 20.180 44.590 20.440 ;
        RECT 44.820 20.425 44.960 20.580 ;
        RECT 48.870 20.520 49.190 20.580 ;
        RECT 44.745 20.195 45.035 20.425 ;
        RECT 45.190 20.180 45.510 20.440 ;
        RECT 46.125 20.380 46.415 20.425 ;
        RECT 47.950 20.380 48.270 20.440 ;
        RECT 50.340 20.425 50.480 20.580 ;
        RECT 51.260 20.580 56.460 20.720 ;
        RECT 46.125 20.240 48.270 20.380 ;
        RECT 46.125 20.195 46.415 20.240 ;
        RECT 47.950 20.180 48.270 20.240 ;
        RECT 49.805 20.195 50.095 20.425 ;
        RECT 50.265 20.195 50.555 20.425 ;
        RECT 33.690 20.040 34.010 20.100 ;
        RECT 31.020 19.900 34.010 20.040 ;
        RECT 33.690 19.840 34.010 19.900 ;
        RECT 34.165 20.040 34.455 20.085 ;
        RECT 35.850 20.040 36.140 20.085 ;
        RECT 49.880 20.040 50.020 20.195 ;
        RECT 50.710 20.180 51.030 20.440 ;
        RECT 51.260 20.040 51.400 20.580 ;
        RECT 56.320 20.440 56.460 20.580 ;
        RECT 59.425 20.580 63.425 20.720 ;
        RECT 59.425 20.535 59.715 20.580 ;
        RECT 60.615 20.535 60.905 20.580 ;
        RECT 63.135 20.535 63.425 20.580 ;
        RECT 66.785 20.720 67.075 20.765 ;
        RECT 67.975 20.720 68.265 20.765 ;
        RECT 70.495 20.720 70.785 20.765 ;
        RECT 66.785 20.580 70.785 20.720 ;
        RECT 66.785 20.535 67.075 20.580 ;
        RECT 67.975 20.535 68.265 20.580 ;
        RECT 70.495 20.535 70.785 20.580 ;
        RECT 74.170 20.720 74.490 20.780 ;
        RECT 76.930 20.720 77.250 20.780 ;
        RECT 79.780 20.720 79.920 20.860 ;
        RECT 74.170 20.580 75.320 20.720 ;
        RECT 74.170 20.520 74.490 20.580 ;
        RECT 51.645 20.195 51.935 20.425 ;
        RECT 34.165 19.900 36.140 20.040 ;
        RECT 34.165 19.855 34.455 19.900 ;
        RECT 35.850 19.855 36.140 19.900 ;
        RECT 36.540 19.900 51.400 20.040 ;
        RECT 51.720 20.040 51.860 20.195 ;
        RECT 55.770 20.180 56.090 20.440 ;
        RECT 56.230 20.180 56.550 20.440 ;
        RECT 56.690 20.180 57.010 20.440 ;
        RECT 57.150 20.180 57.470 20.440 ;
        RECT 58.085 20.195 58.375 20.425 ;
        RECT 55.860 20.040 56.000 20.180 ;
        RECT 58.160 20.040 58.300 20.195 ;
        RECT 58.530 20.180 58.850 20.440 ;
        RECT 58.990 20.380 59.310 20.440 ;
        RECT 59.825 20.380 60.115 20.425 ;
        RECT 58.990 20.240 60.115 20.380 ;
        RECT 58.990 20.180 59.310 20.240 ;
        RECT 59.825 20.195 60.115 20.240 ;
        RECT 65.905 20.380 66.195 20.425 ;
        RECT 70.030 20.380 70.350 20.440 ;
        RECT 65.905 20.240 70.350 20.380 ;
        RECT 65.905 20.195 66.195 20.240 ;
        RECT 70.030 20.180 70.350 20.240 ;
        RECT 74.630 20.180 74.950 20.440 ;
        RECT 75.180 20.425 75.320 20.580 ;
        RECT 76.560 20.580 79.920 20.720 ;
        RECT 80.255 20.580 84.060 20.720 ;
        RECT 75.105 20.195 75.395 20.425 ;
        RECT 75.550 20.180 75.870 20.440 ;
        RECT 76.560 20.425 76.700 20.580 ;
        RECT 76.930 20.520 77.250 20.580 ;
        RECT 80.255 20.440 80.395 20.580 ;
        RECT 76.485 20.195 76.775 20.425 ;
        RECT 78.770 20.180 79.090 20.440 ;
        RECT 79.690 20.180 80.010 20.440 ;
        RECT 80.150 20.180 80.470 20.440 ;
        RECT 80.610 20.180 80.930 20.440 ;
        RECT 81.530 20.380 81.850 20.440 ;
        RECT 83.920 20.425 84.060 20.580 ;
        RECT 84.380 20.425 84.520 20.920 ;
        RECT 85.210 20.920 89.195 21.060 ;
        RECT 85.210 20.860 85.530 20.920 ;
        RECT 88.905 20.875 89.195 20.920 ;
        RECT 82.465 20.380 82.755 20.425 ;
        RECT 81.530 20.240 82.755 20.380 ;
        RECT 81.530 20.180 81.850 20.240 ;
        RECT 82.465 20.195 82.755 20.240 ;
        RECT 83.385 20.180 83.675 20.410 ;
        RECT 83.845 20.195 84.135 20.425 ;
        RECT 84.305 20.195 84.595 20.425 ;
        RECT 86.130 20.180 86.450 20.440 ;
        RECT 87.970 20.180 88.290 20.440 ;
        RECT 67.270 20.085 67.590 20.100 ;
        RECT 67.240 20.040 67.590 20.085 ;
        RECT 51.720 19.900 58.300 20.040 ;
        RECT 67.075 19.900 67.590 20.040 ;
        RECT 28.630 19.700 28.950 19.760 ;
        RECT 28.260 19.560 28.950 19.700 ;
        RECT 20.810 19.500 21.130 19.560 ;
        RECT 21.745 19.515 22.035 19.560 ;
        RECT 28.630 19.500 28.950 19.560 ;
        RECT 30.470 19.500 30.790 19.760 ;
        RECT 32.770 19.700 33.090 19.760 ;
        RECT 36.540 19.700 36.680 19.900 ;
        RECT 67.240 19.855 67.590 19.900 ;
        RECT 67.270 19.840 67.590 19.855 ;
        RECT 83.460 19.760 83.600 20.180 ;
        RECT 32.770 19.560 36.680 19.700 ;
        RECT 32.770 19.500 33.090 19.560 ;
        RECT 42.890 19.500 43.210 19.760 ;
        RECT 48.410 19.500 48.730 19.760 ;
        RECT 54.865 19.700 55.155 19.745 ;
        RECT 55.770 19.700 56.090 19.760 ;
        RECT 54.865 19.560 56.090 19.700 ;
        RECT 54.865 19.515 55.155 19.560 ;
        RECT 55.770 19.500 56.090 19.560 ;
        RECT 58.070 19.700 58.390 19.760 ;
        RECT 62.670 19.700 62.990 19.760 ;
        RECT 58.070 19.560 62.990 19.700 ;
        RECT 58.070 19.500 58.390 19.560 ;
        RECT 62.670 19.500 62.990 19.560 ;
        RECT 65.445 19.700 65.735 19.745 ;
        RECT 67.730 19.700 68.050 19.760 ;
        RECT 65.445 19.560 68.050 19.700 ;
        RECT 65.445 19.515 65.735 19.560 ;
        RECT 67.730 19.500 68.050 19.560 ;
        RECT 73.250 19.500 73.570 19.760 ;
        RECT 78.770 19.700 79.090 19.760 ;
        RECT 81.530 19.700 81.850 19.760 ;
        RECT 78.770 19.560 81.850 19.700 ;
        RECT 78.770 19.500 79.090 19.560 ;
        RECT 81.530 19.500 81.850 19.560 ;
        RECT 82.005 19.700 82.295 19.745 ;
        RECT 82.450 19.700 82.770 19.760 ;
        RECT 82.005 19.560 82.770 19.700 ;
        RECT 82.005 19.515 82.295 19.560 ;
        RECT 82.450 19.500 82.770 19.560 ;
        RECT 83.370 19.500 83.690 19.760 ;
        RECT 84.750 19.700 85.070 19.760 ;
        RECT 85.685 19.700 85.975 19.745 ;
        RECT 84.750 19.560 85.975 19.700 ;
        RECT 84.750 19.500 85.070 19.560 ;
        RECT 85.685 19.515 85.975 19.560 ;
        RECT 87.050 19.500 87.370 19.760 ;
        RECT 13.380 18.880 92.040 19.360 ;
        RECT 17.590 18.480 17.910 18.740 ;
        RECT 21.730 18.680 22.050 18.740 ;
        RECT 18.140 18.540 22.050 18.680 ;
        RECT 15.765 18.340 16.055 18.385 ;
        RECT 16.210 18.340 16.530 18.400 ;
        RECT 15.765 18.200 16.530 18.340 ;
        RECT 15.765 18.155 16.055 18.200 ;
        RECT 16.210 18.140 16.530 18.200 ;
        RECT 16.685 18.340 16.975 18.385 ;
        RECT 18.140 18.340 18.280 18.540 ;
        RECT 21.730 18.480 22.050 18.540 ;
        RECT 28.630 18.480 28.950 18.740 ;
        RECT 31.850 18.680 32.170 18.740 ;
        RECT 36.465 18.680 36.755 18.725 ;
        RECT 31.850 18.540 36.755 18.680 ;
        RECT 31.850 18.480 32.170 18.540 ;
        RECT 36.465 18.495 36.755 18.540 ;
        RECT 49.330 18.680 49.650 18.740 ;
        RECT 54.865 18.680 55.155 18.725 ;
        RECT 49.330 18.540 55.155 18.680 ;
        RECT 49.330 18.480 49.650 18.540 ;
        RECT 54.865 18.495 55.155 18.540 ;
        RECT 57.150 18.680 57.470 18.740 ;
        RECT 62.685 18.680 62.975 18.725 ;
        RECT 72.790 18.680 73.110 18.740 ;
        RECT 57.150 18.540 62.975 18.680 ;
        RECT 57.150 18.480 57.470 18.540 ;
        RECT 62.685 18.495 62.975 18.540 ;
        RECT 66.900 18.540 73.110 18.680 ;
        RECT 30.470 18.385 30.790 18.400 ;
        RECT 30.440 18.340 30.790 18.385 ;
        RECT 16.685 18.200 18.280 18.340 ;
        RECT 18.600 18.200 28.400 18.340 ;
        RECT 30.275 18.200 30.790 18.340 ;
        RECT 16.685 18.155 16.975 18.200 ;
        RECT 18.050 18.000 18.370 18.060 ;
        RECT 18.600 18.000 18.740 18.200 ;
        RECT 28.260 18.060 28.400 18.200 ;
        RECT 30.440 18.155 30.790 18.200 ;
        RECT 30.470 18.140 30.790 18.155 ;
        RECT 35.070 18.340 35.390 18.400 ;
        RECT 37.385 18.340 37.675 18.385 ;
        RECT 41.970 18.340 42.290 18.400 ;
        RECT 35.070 18.200 42.290 18.340 ;
        RECT 35.070 18.140 35.390 18.200 ;
        RECT 37.385 18.155 37.675 18.200 ;
        RECT 41.970 18.140 42.290 18.200 ;
        RECT 42.890 18.340 43.210 18.400 ;
        RECT 45.710 18.340 46.000 18.385 ;
        RECT 58.530 18.340 58.850 18.400 ;
        RECT 42.890 18.200 46.000 18.340 ;
        RECT 42.890 18.140 43.210 18.200 ;
        RECT 45.710 18.155 46.000 18.200 ;
        RECT 48.040 18.200 58.850 18.340 ;
        RECT 18.970 18.000 19.290 18.060 ;
        RECT 20.810 18.045 21.130 18.060 ;
        RECT 19.445 18.000 19.735 18.045 ;
        RECT 20.780 18.000 21.130 18.045 ;
        RECT 18.050 17.860 19.735 18.000 ;
        RECT 20.615 17.860 21.130 18.000 ;
        RECT 18.050 17.800 18.370 17.860 ;
        RECT 18.970 17.800 19.290 17.860 ;
        RECT 19.445 17.815 19.735 17.860 ;
        RECT 20.780 17.815 21.130 17.860 ;
        RECT 20.810 17.800 21.130 17.815 ;
        RECT 23.570 18.000 23.890 18.060 ;
        RECT 26.805 18.000 27.095 18.045 ;
        RECT 27.250 18.000 27.570 18.060 ;
        RECT 23.570 17.860 26.560 18.000 ;
        RECT 23.570 17.800 23.890 17.860 ;
        RECT 20.325 17.660 20.615 17.705 ;
        RECT 21.515 17.660 21.805 17.705 ;
        RECT 24.035 17.660 24.325 17.705 ;
        RECT 20.325 17.520 24.325 17.660 ;
        RECT 26.420 17.660 26.560 17.860 ;
        RECT 26.805 17.860 27.570 18.000 ;
        RECT 26.805 17.815 27.095 17.860 ;
        RECT 27.250 17.800 27.570 17.860 ;
        RECT 27.725 17.815 28.015 18.045 ;
        RECT 28.170 18.000 28.490 18.060 ;
        RECT 48.040 18.045 48.180 18.200 ;
        RECT 29.105 18.000 29.395 18.045 ;
        RECT 28.170 17.860 29.395 18.000 ;
        RECT 27.800 17.660 27.940 17.815 ;
        RECT 28.170 17.800 28.490 17.860 ;
        RECT 29.105 17.815 29.395 17.860 ;
        RECT 29.640 17.860 35.760 18.000 ;
        RECT 29.640 17.660 29.780 17.860 ;
        RECT 26.420 17.520 27.940 17.660 ;
        RECT 20.325 17.475 20.615 17.520 ;
        RECT 21.515 17.475 21.805 17.520 ;
        RECT 24.035 17.475 24.325 17.520 ;
        RECT 19.930 17.320 20.220 17.365 ;
        RECT 22.030 17.320 22.320 17.365 ;
        RECT 23.600 17.320 23.890 17.365 ;
        RECT 19.930 17.180 23.890 17.320 ;
        RECT 19.930 17.135 20.220 17.180 ;
        RECT 22.030 17.135 22.320 17.180 ;
        RECT 23.600 17.135 23.890 17.180 ;
        RECT 26.330 16.780 26.650 17.040 ;
        RECT 27.800 16.980 27.940 17.520 ;
        RECT 28.260 17.520 29.780 17.660 ;
        RECT 29.985 17.660 30.275 17.705 ;
        RECT 31.175 17.660 31.465 17.705 ;
        RECT 33.695 17.660 33.985 17.705 ;
        RECT 29.985 17.520 33.985 17.660 ;
        RECT 35.620 17.660 35.760 17.860 ;
        RECT 38.305 17.815 38.595 18.045 ;
        RECT 47.045 18.000 47.335 18.045 ;
        RECT 47.965 18.000 48.255 18.045 ;
        RECT 47.045 17.860 48.255 18.000 ;
        RECT 47.045 17.815 47.335 17.860 ;
        RECT 47.965 17.815 48.255 17.860 ;
        RECT 48.410 18.000 48.730 18.060 ;
        RECT 55.400 18.045 55.540 18.200 ;
        RECT 58.530 18.140 58.850 18.200 ;
        RECT 64.050 18.340 64.370 18.400 ;
        RECT 66.900 18.385 67.040 18.540 ;
        RECT 72.790 18.480 73.110 18.540 ;
        RECT 75.550 18.680 75.870 18.740 ;
        RECT 79.245 18.680 79.535 18.725 ;
        RECT 75.550 18.540 79.535 18.680 ;
        RECT 75.550 18.480 75.870 18.540 ;
        RECT 79.245 18.495 79.535 18.540 ;
        RECT 80.150 18.680 80.470 18.740 ;
        RECT 87.970 18.680 88.290 18.740 ;
        RECT 80.150 18.540 88.290 18.680 ;
        RECT 80.150 18.480 80.470 18.540 ;
        RECT 87.970 18.480 88.290 18.540 ;
        RECT 64.525 18.340 64.815 18.385 ;
        RECT 64.050 18.200 64.815 18.340 ;
        RECT 64.050 18.140 64.370 18.200 ;
        RECT 64.525 18.155 64.815 18.200 ;
        RECT 66.825 18.155 67.115 18.385 ;
        RECT 67.270 18.140 67.590 18.400 ;
        RECT 81.070 18.340 81.390 18.400 ;
        RECT 71.040 18.200 81.390 18.340 ;
        RECT 49.245 18.000 49.535 18.045 ;
        RECT 48.410 17.860 49.535 18.000 ;
        RECT 36.910 17.660 37.230 17.720 ;
        RECT 38.380 17.660 38.520 17.815 ;
        RECT 48.410 17.800 48.730 17.860 ;
        RECT 49.245 17.815 49.535 17.860 ;
        RECT 55.325 17.815 55.615 18.045 ;
        RECT 55.770 18.000 56.090 18.060 ;
        RECT 56.605 18.000 56.895 18.045 ;
        RECT 55.770 17.860 56.895 18.000 ;
        RECT 55.770 17.800 56.090 17.860 ;
        RECT 56.605 17.815 56.895 17.860 ;
        RECT 63.605 17.815 63.895 18.045 ;
        RECT 35.620 17.520 38.520 17.660 ;
        RECT 42.455 17.660 42.745 17.705 ;
        RECT 44.975 17.660 45.265 17.705 ;
        RECT 46.165 17.660 46.455 17.705 ;
        RECT 42.455 17.520 46.455 17.660 ;
        RECT 28.260 17.380 28.400 17.520 ;
        RECT 29.985 17.475 30.275 17.520 ;
        RECT 31.175 17.475 31.465 17.520 ;
        RECT 33.695 17.475 33.985 17.520 ;
        RECT 36.910 17.460 37.230 17.520 ;
        RECT 42.455 17.475 42.745 17.520 ;
        RECT 44.975 17.475 45.265 17.520 ;
        RECT 46.165 17.475 46.455 17.520 ;
        RECT 48.845 17.660 49.135 17.705 ;
        RECT 50.035 17.660 50.325 17.705 ;
        RECT 52.555 17.660 52.845 17.705 ;
        RECT 48.845 17.520 52.845 17.660 ;
        RECT 48.845 17.475 49.135 17.520 ;
        RECT 50.035 17.475 50.325 17.520 ;
        RECT 52.555 17.475 52.845 17.520 ;
        RECT 56.205 17.660 56.495 17.705 ;
        RECT 57.395 17.660 57.685 17.705 ;
        RECT 59.915 17.660 60.205 17.705 ;
        RECT 63.680 17.660 63.820 17.815 ;
        RECT 66.350 17.800 66.670 18.060 ;
        RECT 68.205 17.815 68.495 18.045 ;
        RECT 71.040 18.000 71.180 18.200 ;
        RECT 81.070 18.140 81.390 18.200 ;
        RECT 70.580 17.860 71.180 18.000 ;
        RECT 71.380 18.000 71.670 18.045 ;
        RECT 73.250 18.000 73.570 18.060 ;
        RECT 71.380 17.860 73.570 18.000 ;
        RECT 64.970 17.660 65.290 17.720 ;
        RECT 68.280 17.660 68.420 17.815 ;
        RECT 56.205 17.520 60.205 17.660 ;
        RECT 56.205 17.475 56.495 17.520 ;
        RECT 57.395 17.475 57.685 17.520 ;
        RECT 59.915 17.475 60.205 17.520 ;
        RECT 62.300 17.520 68.420 17.660 ;
        RECT 70.030 17.660 70.350 17.720 ;
        RECT 70.580 17.660 70.720 17.860 ;
        RECT 71.380 17.815 71.670 17.860 ;
        RECT 73.250 17.800 73.570 17.860 ;
        RECT 77.390 17.800 77.710 18.060 ;
        RECT 78.325 18.000 78.615 18.045 ;
        RECT 79.230 18.000 79.550 18.060 ;
        RECT 82.450 18.045 82.770 18.060 ;
        RECT 82.420 18.000 82.770 18.045 ;
        RECT 78.325 17.860 79.550 18.000 ;
        RECT 82.255 17.860 82.770 18.000 ;
        RECT 78.325 17.815 78.615 17.860 ;
        RECT 70.030 17.520 70.720 17.660 ;
        RECT 70.925 17.660 71.215 17.705 ;
        RECT 72.115 17.660 72.405 17.705 ;
        RECT 74.635 17.660 74.925 17.705 ;
        RECT 70.925 17.520 74.925 17.660 ;
        RECT 28.170 17.120 28.490 17.380 ;
        RECT 29.590 17.320 29.880 17.365 ;
        RECT 31.690 17.320 31.980 17.365 ;
        RECT 33.260 17.320 33.550 17.365 ;
        RECT 40.590 17.320 40.910 17.380 ;
        RECT 62.300 17.365 62.440 17.520 ;
        RECT 64.970 17.460 65.290 17.520 ;
        RECT 70.030 17.460 70.350 17.520 ;
        RECT 70.925 17.475 71.215 17.520 ;
        RECT 72.115 17.475 72.405 17.520 ;
        RECT 74.635 17.475 74.925 17.520 ;
        RECT 29.590 17.180 33.550 17.320 ;
        RECT 29.590 17.135 29.880 17.180 ;
        RECT 31.690 17.135 31.980 17.180 ;
        RECT 33.260 17.135 33.550 17.180 ;
        RECT 36.080 17.180 40.910 17.320 ;
        RECT 36.080 17.025 36.220 17.180 ;
        RECT 40.590 17.120 40.910 17.180 ;
        RECT 42.890 17.320 43.180 17.365 ;
        RECT 44.460 17.320 44.750 17.365 ;
        RECT 46.560 17.320 46.850 17.365 ;
        RECT 42.890 17.180 46.850 17.320 ;
        RECT 42.890 17.135 43.180 17.180 ;
        RECT 44.460 17.135 44.750 17.180 ;
        RECT 46.560 17.135 46.850 17.180 ;
        RECT 48.450 17.320 48.740 17.365 ;
        RECT 50.550 17.320 50.840 17.365 ;
        RECT 52.120 17.320 52.410 17.365 ;
        RECT 48.450 17.180 52.410 17.320 ;
        RECT 48.450 17.135 48.740 17.180 ;
        RECT 50.550 17.135 50.840 17.180 ;
        RECT 52.120 17.135 52.410 17.180 ;
        RECT 55.810 17.320 56.100 17.365 ;
        RECT 57.910 17.320 58.200 17.365 ;
        RECT 59.480 17.320 59.770 17.365 ;
        RECT 55.810 17.180 59.770 17.320 ;
        RECT 55.810 17.135 56.100 17.180 ;
        RECT 57.910 17.135 58.200 17.180 ;
        RECT 59.480 17.135 59.770 17.180 ;
        RECT 62.225 17.135 62.515 17.365 ;
        RECT 62.670 17.320 62.990 17.380 ;
        RECT 70.530 17.320 70.820 17.365 ;
        RECT 72.630 17.320 72.920 17.365 ;
        RECT 74.200 17.320 74.490 17.365 ;
        RECT 62.670 17.180 70.030 17.320 ;
        RECT 62.670 17.120 62.990 17.180 ;
        RECT 36.005 16.980 36.295 17.025 ;
        RECT 27.800 16.840 36.295 16.980 ;
        RECT 36.005 16.795 36.295 16.840 ;
        RECT 38.750 16.980 39.070 17.040 ;
        RECT 40.145 16.980 40.435 17.025 ;
        RECT 38.750 16.840 40.435 16.980 ;
        RECT 38.750 16.780 39.070 16.840 ;
        RECT 40.145 16.795 40.435 16.840 ;
        RECT 53.470 16.980 53.790 17.040 ;
        RECT 65.445 16.980 65.735 17.025 ;
        RECT 53.470 16.840 65.735 16.980 ;
        RECT 69.890 16.980 70.030 17.180 ;
        RECT 70.530 17.180 74.490 17.320 ;
        RECT 70.530 17.135 70.820 17.180 ;
        RECT 72.630 17.135 72.920 17.180 ;
        RECT 74.200 17.135 74.490 17.180 ;
        RECT 76.945 17.320 77.235 17.365 ;
        RECT 77.390 17.320 77.710 17.380 ;
        RECT 78.400 17.320 78.540 17.815 ;
        RECT 79.230 17.800 79.550 17.860 ;
        RECT 82.420 17.815 82.770 17.860 ;
        RECT 82.450 17.800 82.770 17.815 ;
        RECT 83.830 18.000 84.150 18.060 ;
        RECT 88.445 18.000 88.735 18.045 ;
        RECT 83.830 17.860 88.735 18.000 ;
        RECT 83.830 17.800 84.150 17.860 ;
        RECT 88.445 17.815 88.735 17.860 ;
        RECT 81.070 17.460 81.390 17.720 ;
        RECT 81.965 17.660 82.255 17.705 ;
        RECT 83.155 17.660 83.445 17.705 ;
        RECT 85.675 17.660 85.965 17.705 ;
        RECT 81.965 17.520 85.965 17.660 ;
        RECT 81.965 17.475 82.255 17.520 ;
        RECT 83.155 17.475 83.445 17.520 ;
        RECT 85.675 17.475 85.965 17.520 ;
        RECT 76.945 17.180 78.540 17.320 ;
        RECT 81.570 17.320 81.860 17.365 ;
        RECT 83.670 17.320 83.960 17.365 ;
        RECT 85.240 17.320 85.530 17.365 ;
        RECT 81.570 17.180 85.530 17.320 ;
        RECT 76.945 17.135 77.235 17.180 ;
        RECT 77.390 17.120 77.710 17.180 ;
        RECT 81.570 17.135 81.860 17.180 ;
        RECT 83.670 17.135 83.960 17.180 ;
        RECT 85.240 17.135 85.530 17.180 ;
        RECT 80.610 16.980 80.930 17.040 ;
        RECT 69.890 16.840 80.930 16.980 ;
        RECT 53.470 16.780 53.790 16.840 ;
        RECT 65.445 16.795 65.735 16.840 ;
        RECT 80.610 16.780 80.930 16.840 ;
        RECT 89.350 16.780 89.670 17.040 ;
        RECT 13.380 16.160 92.040 16.640 ;
        RECT 21.730 15.760 22.050 16.020 ;
        RECT 23.125 15.960 23.415 16.005 ;
        RECT 24.030 15.960 24.350 16.020 ;
        RECT 42.430 15.960 42.750 16.020 ;
        RECT 23.125 15.820 24.350 15.960 ;
        RECT 23.125 15.775 23.415 15.820 ;
        RECT 24.030 15.760 24.350 15.820 ;
        RECT 33.320 15.820 42.750 15.960 ;
        RECT 15.330 15.620 15.620 15.665 ;
        RECT 17.430 15.620 17.720 15.665 ;
        RECT 19.000 15.620 19.290 15.665 ;
        RECT 15.330 15.480 19.290 15.620 ;
        RECT 15.330 15.435 15.620 15.480 ;
        RECT 17.430 15.435 17.720 15.480 ;
        RECT 19.000 15.435 19.290 15.480 ;
        RECT 15.725 15.280 16.015 15.325 ;
        RECT 16.915 15.280 17.205 15.325 ;
        RECT 19.435 15.280 19.725 15.325 ;
        RECT 15.725 15.140 19.725 15.280 ;
        RECT 15.725 15.095 16.015 15.140 ;
        RECT 16.915 15.095 17.205 15.140 ;
        RECT 19.435 15.095 19.725 15.140 ;
        RECT 14.845 14.940 15.135 14.985 ;
        RECT 18.970 14.940 19.290 15.000 ;
        RECT 14.845 14.800 19.290 14.940 ;
        RECT 14.845 14.755 15.135 14.800 ;
        RECT 18.970 14.740 19.290 14.800 ;
        RECT 24.045 14.940 24.335 14.985 ;
        RECT 26.330 14.940 26.650 15.000 ;
        RECT 24.045 14.800 26.650 14.940 ;
        RECT 24.045 14.755 24.335 14.800 ;
        RECT 26.330 14.740 26.650 14.800 ;
        RECT 29.105 14.940 29.395 14.985 ;
        RECT 30.930 14.940 31.250 15.000 ;
        RECT 29.105 14.800 31.250 14.940 ;
        RECT 29.105 14.755 29.395 14.800 ;
        RECT 30.930 14.740 31.250 14.800 ;
        RECT 31.390 14.740 31.710 15.000 ;
        RECT 33.320 14.985 33.460 15.820 ;
        RECT 42.430 15.760 42.750 15.820 ;
        RECT 45.190 15.960 45.510 16.020 ;
        RECT 45.665 15.960 45.955 16.005 ;
        RECT 45.190 15.820 45.955 15.960 ;
        RECT 45.190 15.760 45.510 15.820 ;
        RECT 45.665 15.775 45.955 15.820 ;
        RECT 50.710 15.960 51.030 16.020 ;
        RECT 51.645 15.960 51.935 16.005 ;
        RECT 50.710 15.820 51.935 15.960 ;
        RECT 50.710 15.760 51.030 15.820 ;
        RECT 51.645 15.775 51.935 15.820 ;
        RECT 79.690 15.960 80.010 16.020 ;
        RECT 80.165 15.960 80.455 16.005 ;
        RECT 79.690 15.820 80.455 15.960 ;
        RECT 79.690 15.760 80.010 15.820 ;
        RECT 80.165 15.775 80.455 15.820 ;
        RECT 82.465 15.960 82.755 16.005 ;
        RECT 83.370 15.960 83.690 16.020 ;
        RECT 82.465 15.820 83.690 15.960 ;
        RECT 82.465 15.775 82.755 15.820 ;
        RECT 83.370 15.760 83.690 15.820 ;
        RECT 34.165 15.620 34.455 15.665 ;
        RECT 36.910 15.620 37.230 15.680 ;
        RECT 34.165 15.480 37.230 15.620 ;
        RECT 34.165 15.435 34.455 15.480 ;
        RECT 36.910 15.420 37.230 15.480 ;
        RECT 43.365 15.620 43.655 15.665 ;
        RECT 47.950 15.620 48.270 15.680 ;
        RECT 43.365 15.480 48.270 15.620 ;
        RECT 43.365 15.435 43.655 15.480 ;
        RECT 47.950 15.420 48.270 15.480 ;
        RECT 83.870 15.620 84.160 15.665 ;
        RECT 85.970 15.620 86.260 15.665 ;
        RECT 87.540 15.620 87.830 15.665 ;
        RECT 83.870 15.480 87.830 15.620 ;
        RECT 83.870 15.435 84.160 15.480 ;
        RECT 85.970 15.435 86.260 15.480 ;
        RECT 87.540 15.435 87.830 15.480 ;
        RECT 55.310 15.280 55.630 15.340 ;
        RECT 69.110 15.280 69.430 15.340 ;
        RECT 80.150 15.280 80.470 15.340 ;
        RECT 38.840 15.140 44.960 15.280 ;
        RECT 38.840 15.000 38.980 15.140 ;
        RECT 33.245 14.755 33.535 14.985 ;
        RECT 35.070 14.740 35.390 15.000 ;
        RECT 36.925 14.940 37.215 14.985 ;
        RECT 37.830 14.940 38.150 15.000 ;
        RECT 36.925 14.800 38.150 14.940 ;
        RECT 36.925 14.755 37.215 14.800 ;
        RECT 37.830 14.740 38.150 14.800 ;
        RECT 38.750 14.740 39.070 15.000 ;
        RECT 40.590 14.740 40.910 15.000 ;
        RECT 41.050 14.940 41.370 15.000 ;
        RECT 42.060 14.985 42.200 15.140 ;
        RECT 41.525 14.940 41.815 14.985 ;
        RECT 41.050 14.800 41.815 14.940 ;
        RECT 41.050 14.740 41.370 14.800 ;
        RECT 41.525 14.755 41.815 14.800 ;
        RECT 41.985 14.755 42.275 14.985 ;
        RECT 42.445 14.940 42.735 14.985 ;
        RECT 44.270 14.940 44.590 15.000 ;
        RECT 44.820 14.985 44.960 15.140 ;
        RECT 55.310 15.140 60.140 15.280 ;
        RECT 55.310 15.080 55.630 15.140 ;
        RECT 42.445 14.800 44.590 14.940 ;
        RECT 42.445 14.755 42.735 14.800 ;
        RECT 44.270 14.740 44.590 14.800 ;
        RECT 44.745 14.755 45.035 14.985 ;
        RECT 45.650 14.940 45.970 15.000 ;
        RECT 47.505 14.940 47.795 14.985 ;
        RECT 45.650 14.800 47.795 14.940 ;
        RECT 45.650 14.740 45.970 14.800 ;
        RECT 47.505 14.755 47.795 14.800 ;
        RECT 47.965 14.940 48.255 14.985 ;
        RECT 49.330 14.940 49.650 15.000 ;
        RECT 50.725 14.940 51.015 14.985 ;
        RECT 47.965 14.800 51.015 14.940 ;
        RECT 47.965 14.755 48.255 14.800 ;
        RECT 49.330 14.740 49.650 14.800 ;
        RECT 50.725 14.755 51.015 14.800 ;
        RECT 54.865 14.940 55.155 14.985 ;
        RECT 57.610 14.940 57.930 15.000 ;
        RECT 60.000 14.985 60.140 15.140 ;
        RECT 69.110 15.140 80.470 15.280 ;
        RECT 69.110 15.080 69.430 15.140 ;
        RECT 54.865 14.800 57.930 14.940 ;
        RECT 54.865 14.755 55.155 14.800 ;
        RECT 57.610 14.740 57.930 14.800 ;
        RECT 58.085 14.755 58.375 14.985 ;
        RECT 59.925 14.755 60.215 14.985 ;
        RECT 64.525 14.940 64.815 14.985 ;
        RECT 64.970 14.940 65.290 15.000 ;
        RECT 64.525 14.800 65.290 14.940 ;
        RECT 64.525 14.755 64.815 14.800 ;
        RECT 15.290 14.600 15.610 14.660 ;
        RECT 16.070 14.600 16.360 14.645 ;
        RECT 15.290 14.460 16.360 14.600 ;
        RECT 15.290 14.400 15.610 14.460 ;
        RECT 16.070 14.415 16.360 14.460 ;
        RECT 24.965 14.600 25.255 14.645 ;
        RECT 26.790 14.600 27.110 14.660 ;
        RECT 40.130 14.600 40.450 14.660 ;
        RECT 24.965 14.460 27.110 14.600 ;
        RECT 24.965 14.415 25.255 14.460 ;
        RECT 26.790 14.400 27.110 14.460 ;
        RECT 36.080 14.460 40.450 14.600 ;
        RECT 27.250 14.260 27.570 14.320 ;
        RECT 28.185 14.260 28.475 14.305 ;
        RECT 27.250 14.120 28.475 14.260 ;
        RECT 27.250 14.060 27.570 14.120 ;
        RECT 28.185 14.075 28.475 14.120 ;
        RECT 30.470 14.060 30.790 14.320 ;
        RECT 32.325 14.260 32.615 14.305 ;
        RECT 33.690 14.260 34.010 14.320 ;
        RECT 36.080 14.305 36.220 14.460 ;
        RECT 40.130 14.400 40.450 14.460 ;
        RECT 43.825 14.600 44.115 14.645 ;
        RECT 49.790 14.600 50.110 14.660 ;
        RECT 43.825 14.460 50.110 14.600 ;
        RECT 58.160 14.600 58.300 14.755 ;
        RECT 64.970 14.740 65.290 14.800 ;
        RECT 67.730 14.740 68.050 15.000 ;
        RECT 70.950 14.740 71.270 15.000 ;
        RECT 72.790 14.740 73.110 15.000 ;
        RECT 77.390 14.740 77.710 15.000 ;
        RECT 79.320 14.985 79.460 15.140 ;
        RECT 80.150 15.080 80.470 15.140 ;
        RECT 81.070 15.280 81.390 15.340 ;
        RECT 83.385 15.280 83.675 15.325 ;
        RECT 81.070 15.140 83.675 15.280 ;
        RECT 81.070 15.080 81.390 15.140 ;
        RECT 83.385 15.095 83.675 15.140 ;
        RECT 84.265 15.280 84.555 15.325 ;
        RECT 85.455 15.280 85.745 15.325 ;
        RECT 87.975 15.280 88.265 15.325 ;
        RECT 84.265 15.140 88.265 15.280 ;
        RECT 84.265 15.095 84.555 15.140 ;
        RECT 85.455 15.095 85.745 15.140 ;
        RECT 87.975 15.095 88.265 15.140 ;
        RECT 84.750 14.985 85.070 15.000 ;
        RECT 79.245 14.755 79.535 14.985 ;
        RECT 84.720 14.940 85.070 14.985 ;
        RECT 84.555 14.800 85.070 14.940 ;
        RECT 84.720 14.755 85.070 14.800 ;
        RECT 84.750 14.740 85.070 14.755 ;
        RECT 63.130 14.600 63.450 14.660 ;
        RECT 58.160 14.460 63.450 14.600 ;
        RECT 43.825 14.415 44.115 14.460 ;
        RECT 49.790 14.400 50.110 14.460 ;
        RECT 63.130 14.400 63.450 14.460 ;
        RECT 74.170 14.600 74.490 14.660 ;
        RECT 78.325 14.600 78.615 14.645 ;
        RECT 80.625 14.600 80.915 14.645 ;
        RECT 74.170 14.460 80.915 14.600 ;
        RECT 74.170 14.400 74.490 14.460 ;
        RECT 78.325 14.415 78.615 14.460 ;
        RECT 80.625 14.415 80.915 14.460 ;
        RECT 81.545 14.600 81.835 14.645 ;
        RECT 85.670 14.600 85.990 14.660 ;
        RECT 81.545 14.460 90.500 14.600 ;
        RECT 81.545 14.415 81.835 14.460 ;
        RECT 85.670 14.400 85.990 14.460 ;
        RECT 32.325 14.120 34.010 14.260 ;
        RECT 32.325 14.075 32.615 14.120 ;
        RECT 33.690 14.060 34.010 14.120 ;
        RECT 36.005 14.075 36.295 14.305 ;
        RECT 37.845 14.260 38.135 14.305 ;
        RECT 42.890 14.260 43.210 14.320 ;
        RECT 37.845 14.120 43.210 14.260 ;
        RECT 37.845 14.075 38.135 14.120 ;
        RECT 42.890 14.060 43.210 14.120 ;
        RECT 46.570 14.060 46.890 14.320 ;
        RECT 48.885 14.260 49.175 14.305 ;
        RECT 49.330 14.260 49.650 14.320 ;
        RECT 48.885 14.120 49.650 14.260 ;
        RECT 48.885 14.075 49.175 14.120 ;
        RECT 49.330 14.060 49.650 14.120 ;
        RECT 53.010 14.260 53.330 14.320 ;
        RECT 53.945 14.260 54.235 14.305 ;
        RECT 53.010 14.120 54.235 14.260 ;
        RECT 53.010 14.060 53.330 14.120 ;
        RECT 53.945 14.075 54.235 14.120 ;
        RECT 56.230 14.260 56.550 14.320 ;
        RECT 57.165 14.260 57.455 14.305 ;
        RECT 56.230 14.120 57.455 14.260 ;
        RECT 56.230 14.060 56.550 14.120 ;
        RECT 57.165 14.075 57.455 14.120 ;
        RECT 59.450 14.260 59.770 14.320 ;
        RECT 60.845 14.260 61.135 14.305 ;
        RECT 59.450 14.120 61.135 14.260 ;
        RECT 59.450 14.060 59.770 14.120 ;
        RECT 60.845 14.075 61.135 14.120 ;
        RECT 62.670 14.260 62.990 14.320 ;
        RECT 63.605 14.260 63.895 14.305 ;
        RECT 62.670 14.120 63.895 14.260 ;
        RECT 62.670 14.060 62.990 14.120 ;
        RECT 63.605 14.075 63.895 14.120 ;
        RECT 65.890 14.260 66.210 14.320 ;
        RECT 66.825 14.260 67.115 14.305 ;
        RECT 65.890 14.120 67.115 14.260 ;
        RECT 65.890 14.060 66.210 14.120 ;
        RECT 66.825 14.075 67.115 14.120 ;
        RECT 69.110 14.260 69.430 14.320 ;
        RECT 70.045 14.260 70.335 14.305 ;
        RECT 69.110 14.120 70.335 14.260 ;
        RECT 69.110 14.060 69.430 14.120 ;
        RECT 70.045 14.075 70.335 14.120 ;
        RECT 72.330 14.260 72.650 14.320 ;
        RECT 73.725 14.260 74.015 14.305 ;
        RECT 72.330 14.120 74.015 14.260 ;
        RECT 72.330 14.060 72.650 14.120 ;
        RECT 73.725 14.075 74.015 14.120 ;
        RECT 75.550 14.260 75.870 14.320 ;
        RECT 90.360 14.305 90.500 14.460 ;
        RECT 76.485 14.260 76.775 14.305 ;
        RECT 75.550 14.120 76.775 14.260 ;
        RECT 75.550 14.060 75.870 14.120 ;
        RECT 76.485 14.075 76.775 14.120 ;
        RECT 90.285 14.075 90.575 14.305 ;
        RECT 13.380 13.440 92.040 13.920 ;
        RECT 7.930 9.500 8.250 9.560 ;
        RECT 15.750 9.500 16.070 9.560 ;
        RECT 7.930 9.360 16.070 9.500 ;
        RECT 7.930 9.300 8.250 9.360 ;
        RECT 15.750 9.300 16.070 9.360 ;
        RECT 78.770 9.500 79.090 9.560 ;
        RECT 89.350 9.500 89.670 9.560 ;
        RECT 78.770 9.360 89.670 9.500 ;
        RECT 78.770 9.300 79.090 9.360 ;
        RECT 89.350 9.300 89.670 9.360 ;
        RECT 11.150 9.160 11.470 9.220 ;
        RECT 19.430 9.160 19.750 9.220 ;
        RECT 11.150 9.020 19.750 9.160 ;
        RECT 11.150 8.960 11.470 9.020 ;
        RECT 19.430 8.960 19.750 9.020 ;
        RECT 81.990 8.480 82.310 8.540 ;
        RECT 87.050 8.480 87.370 8.540 ;
        RECT 81.990 8.340 87.370 8.480 ;
        RECT 81.990 8.280 82.310 8.340 ;
        RECT 87.050 8.280 87.370 8.340 ;
      LAYER met2 ;
        RECT 69.205 222.560 69.595 222.640 ;
        RECT 69.205 222.420 127.660 222.560 ;
        RECT 69.205 222.340 69.595 222.420 ;
        RECT 72.120 222.090 72.420 222.215 ;
        RECT 72.120 221.950 126.920 222.090 ;
        RECT 72.120 221.825 72.420 221.950 ;
        RECT 74.770 221.725 75.160 221.785 ;
        RECT 125.240 221.770 125.770 221.780 ;
        RECT 125.240 221.725 125.805 221.770 ;
        RECT 74.770 221.540 125.805 221.725 ;
        RECT 74.770 221.485 75.160 221.540 ;
        RECT 125.240 221.490 125.805 221.540 ;
        RECT 126.780 221.620 126.920 221.950 ;
        RECT 127.520 222.060 127.660 222.420 ;
        RECT 149.680 222.060 150.000 222.120 ;
        RECT 127.520 221.920 150.000 222.060 ;
        RECT 149.680 221.860 150.000 221.920 ;
        RECT 125.240 221.480 125.770 221.490 ;
        RECT 126.780 221.480 140.200 221.620 ;
        RECT 138.880 221.310 139.370 221.320 ;
        RECT 80.275 221.240 80.665 221.305 ;
        RECT 82.770 221.240 83.840 221.280 ;
        RECT 80.275 221.160 117.550 221.240 ;
        RECT 138.880 221.160 139.405 221.310 ;
        RECT 80.275 221.120 139.405 221.160 ;
        RECT 80.275 221.070 82.940 221.120 ;
        RECT 83.620 221.070 139.405 221.120 ;
        RECT 80.275 221.005 80.665 221.070 ;
        RECT 117.055 221.030 139.405 221.070 ;
        RECT 117.055 221.020 139.370 221.030 ;
        RECT 83.085 220.900 83.475 220.980 ;
        RECT 117.055 220.965 139.130 221.020 ;
        RECT 140.060 221.000 140.200 221.480 ;
        RECT 149.120 221.000 149.440 221.060 ;
        RECT 83.085 220.800 116.760 220.900 ;
        RECT 140.060 220.860 149.440 221.000 ;
        RECT 149.120 220.800 149.440 220.860 ;
        RECT 83.085 220.760 133.370 220.800 ;
        RECT 83.085 220.680 83.475 220.760 ;
        RECT 116.620 220.660 133.370 220.760 ;
        RECT 85.785 220.525 86.175 220.595 ;
        RECT 115.915 220.580 116.285 220.585 ;
        RECT 115.570 220.525 116.285 220.580 ;
        RECT 85.785 220.365 116.285 220.525 ;
        RECT 85.785 220.295 86.175 220.365 ;
        RECT 115.570 220.310 116.285 220.365 ;
        RECT 115.915 220.305 116.285 220.310 ;
        RECT 91.280 220.140 91.670 220.220 ;
        RECT 132.220 220.210 132.610 220.480 ;
        RECT 93.670 220.140 94.650 220.160 ;
        RECT 116.845 220.140 132.610 220.210 ;
        RECT 91.280 220.040 132.610 220.140 ;
        RECT 133.230 220.250 133.370 220.660 ;
        RECT 148.660 220.250 148.920 220.340 ;
        RECT 133.230 220.110 148.920 220.250 ;
        RECT 91.280 220.035 132.510 220.040 ;
        RECT 91.280 220.020 117.005 220.035 ;
        RECT 148.660 220.020 148.920 220.110 ;
        RECT 91.280 219.995 93.810 220.020 ;
        RECT 94.490 220.000 117.005 220.020 ;
        RECT 94.490 219.995 116.860 220.000 ;
        RECT 91.280 219.920 91.670 219.995 ;
        RECT 93.955 219.800 94.345 219.880 ;
        RECT 148.110 219.800 148.430 219.860 ;
        RECT 93.955 219.660 148.430 219.800 ;
        RECT 88.600 219.490 88.900 219.615 ;
        RECT 93.955 219.580 94.345 219.660 ;
        RECT 148.110 219.600 148.430 219.660 ;
        RECT 88.600 219.440 93.810 219.490 ;
        RECT 94.490 219.440 111.950 219.490 ;
        RECT 88.600 219.350 111.950 219.440 ;
        RECT 88.600 219.225 88.900 219.350 ;
        RECT 93.560 219.310 94.730 219.350 ;
        RECT 93.670 219.290 94.610 219.310 ;
        RECT 77.535 219.090 77.925 219.170 ;
        RECT 96.090 219.090 111.560 219.180 ;
        RECT 77.535 219.080 88.440 219.090 ;
        RECT 89.070 219.080 111.560 219.090 ;
        RECT 77.535 219.040 111.560 219.080 ;
        RECT 77.535 218.950 96.230 219.040 ;
        RECT 77.535 218.870 77.925 218.950 ;
        RECT 88.330 218.940 89.190 218.950 ;
        RECT 66.485 218.730 66.875 218.810 ;
        RECT 96.750 218.730 111.150 218.830 ;
        RECT 66.485 218.690 111.150 218.730 ;
        RECT 66.485 218.590 96.890 218.690 ;
        RECT 66.485 218.510 66.875 218.590 ;
        RECT 63.655 218.200 64.045 218.280 ;
        RECT 63.655 218.060 110.150 218.200 ;
        RECT 63.655 217.980 64.045 218.060 ;
        RECT 62.690 208.800 62.970 212.800 ;
        RECT 72.350 208.800 72.630 212.800 ;
        RECT 28.930 201.175 30.470 201.545 ;
        RECT 51.200 200.690 51.460 201.010 ;
        RECT 48.900 199.330 49.160 199.650 ;
        RECT 8.410 198.115 8.690 198.485 ;
        RECT 32.230 198.455 33.770 198.825 ;
        RECT 8.480 112.610 8.620 198.115 ;
        RECT 42.920 197.630 43.180 197.950 ;
        RECT 44.760 197.630 45.020 197.950 ;
        RECT 42.460 197.290 42.720 197.610 ;
        RECT 38.320 196.950 38.580 197.270 ;
        RECT 28.930 195.735 30.470 196.105 ;
        RECT 38.380 194.890 38.520 196.950 ;
        RECT 38.320 194.570 38.580 194.890 ;
        RECT 32.230 193.015 33.770 193.385 ;
        RECT 28.930 190.295 30.470 190.665 ;
        RECT 32.230 187.575 33.770 187.945 ;
        RECT 22.680 186.750 22.940 187.070 ;
        RECT 18.080 186.070 18.340 186.390 ;
        RECT 18.140 184.690 18.280 186.070 ;
        RECT 21.760 185.390 22.020 185.710 ;
        RECT 18.080 184.370 18.340 184.690 ;
        RECT 21.820 183.670 21.960 185.390 ;
        RECT 18.540 183.350 18.800 183.670 ;
        RECT 21.760 183.350 22.020 183.670 ;
        RECT 18.600 181.290 18.740 183.350 ;
        RECT 22.740 181.970 22.880 186.750 ;
        RECT 38.380 186.730 38.520 194.570 ;
        RECT 41.080 193.890 41.340 194.210 ;
        RECT 41.140 192.850 41.280 193.890 ;
        RECT 41.080 192.530 41.340 192.850 ;
        RECT 42.520 191.150 42.660 197.290 ;
        RECT 42.980 192.510 43.120 197.630 ;
        RECT 43.380 197.520 43.640 197.610 ;
        RECT 43.380 197.380 44.040 197.520 ;
        RECT 43.380 197.290 43.640 197.380 ;
        RECT 43.380 196.270 43.640 196.590 ;
        RECT 43.440 192.850 43.580 196.270 ;
        RECT 43.900 192.850 44.040 197.380 ;
        RECT 44.820 195.230 44.960 197.630 ;
        RECT 48.960 197.610 49.100 199.330 ;
        RECT 48.900 197.290 49.160 197.610 ;
        RECT 47.520 196.270 47.780 196.590 ;
        RECT 47.580 195.570 47.720 196.270 ;
        RECT 46.600 195.250 46.860 195.570 ;
        RECT 47.520 195.250 47.780 195.570 ;
        RECT 44.760 194.910 45.020 195.230 ;
        RECT 45.680 193.550 45.940 193.870 ;
        RECT 46.140 193.550 46.400 193.870 ;
        RECT 43.380 192.530 43.640 192.850 ;
        RECT 43.840 192.530 44.100 192.850 ;
        RECT 42.920 192.190 43.180 192.510 ;
        RECT 42.000 190.830 42.260 191.150 ;
        RECT 42.460 190.830 42.720 191.150 ;
        RECT 42.060 190.130 42.200 190.830 ;
        RECT 42.000 189.810 42.260 190.130 ;
        RECT 41.540 188.110 41.800 188.430 ;
        RECT 41.600 187.070 41.740 188.110 ;
        RECT 41.540 186.750 41.800 187.070 ;
        RECT 28.200 186.410 28.460 186.730 ;
        RECT 38.320 186.410 38.580 186.730 ;
        RECT 25.900 186.070 26.160 186.390 ;
        RECT 25.960 183.670 26.100 186.070 ;
        RECT 27.740 185.390 28.000 185.710 ;
        RECT 27.800 184.090 27.940 185.390 ;
        RECT 28.260 184.690 28.400 186.410 ;
        RECT 34.640 185.390 34.900 185.710 ;
        RECT 28.930 184.855 30.470 185.225 ;
        RECT 28.200 184.370 28.460 184.690 ;
        RECT 28.660 184.370 28.920 184.690 ;
        RECT 28.720 184.090 28.860 184.370 ;
        RECT 27.800 183.950 28.860 184.090 ;
        RECT 25.900 183.350 26.160 183.670 ;
        RECT 24.060 182.670 24.320 182.990 ;
        RECT 22.680 181.650 22.940 181.970 ;
        RECT 24.120 181.630 24.260 182.670 ;
        RECT 24.060 181.310 24.320 181.630 ;
        RECT 18.540 180.970 18.800 181.290 ;
        RECT 18.600 179.250 18.740 180.970 ;
        RECT 18.540 178.930 18.800 179.250 ;
        RECT 18.600 176.190 18.740 178.930 ;
        RECT 25.960 178.230 26.100 183.350 ;
        RECT 28.720 180.690 28.860 183.950 ;
        RECT 31.420 183.690 31.680 184.010 ;
        RECT 31.940 183.950 33.000 184.090 ;
        RECT 30.500 183.350 30.760 183.670 ;
        RECT 30.560 181.630 30.700 183.350 ;
        RECT 30.960 182.670 31.220 182.990 ;
        RECT 30.500 181.310 30.760 181.630 ;
        RECT 27.800 180.550 28.860 180.690 ;
        RECT 25.900 177.910 26.160 178.230 ;
        RECT 27.800 177.970 27.940 180.550 ;
        RECT 28.660 180.180 28.920 180.270 ;
        RECT 28.260 180.040 28.920 180.180 ;
        RECT 28.260 178.910 28.400 180.040 ;
        RECT 28.660 179.950 28.920 180.040 ;
        RECT 28.930 179.415 30.470 179.785 ;
        RECT 31.020 179.250 31.160 182.670 ;
        RECT 31.480 181.200 31.620 183.690 ;
        RECT 31.940 183.670 32.080 183.950 ;
        RECT 31.880 183.350 32.140 183.670 ;
        RECT 32.340 183.350 32.600 183.670 ;
        RECT 32.400 182.900 32.540 183.350 ;
        RECT 32.860 182.990 33.000 183.950 ;
        RECT 34.700 183.670 34.840 185.390 ;
        RECT 34.640 183.350 34.900 183.670 ;
        RECT 36.020 183.350 36.280 183.670 ;
        RECT 37.400 183.350 37.660 183.670 ;
        RECT 33.720 183.240 33.980 183.330 ;
        RECT 33.720 183.100 34.380 183.240 ;
        RECT 33.720 183.010 33.980 183.100 ;
        RECT 31.940 182.760 32.540 182.900 ;
        RECT 31.940 181.970 32.080 182.760 ;
        RECT 32.800 182.670 33.060 182.990 ;
        RECT 32.230 182.135 33.770 182.505 ;
        RECT 34.240 181.970 34.380 183.100 ;
        RECT 34.640 182.670 34.900 182.990 ;
        RECT 31.880 181.650 32.140 181.970 ;
        RECT 34.180 181.650 34.440 181.970 ;
        RECT 31.880 181.200 32.140 181.290 ;
        RECT 31.480 181.060 32.140 181.200 ;
        RECT 31.880 180.970 32.140 181.060 ;
        RECT 34.700 180.950 34.840 182.670 ;
        RECT 35.560 181.650 35.820 181.970 ;
        RECT 35.620 181.290 35.760 181.650 ;
        RECT 36.080 181.290 36.220 183.350 ;
        RECT 35.560 180.970 35.820 181.290 ;
        RECT 36.020 180.970 36.280 181.290 ;
        RECT 36.480 180.970 36.740 181.290 ;
        RECT 34.640 180.630 34.900 180.950 ;
        RECT 31.420 179.950 31.680 180.270 ;
        RECT 34.640 179.950 34.900 180.270 ;
        RECT 30.960 178.930 31.220 179.250 ;
        RECT 28.200 178.590 28.460 178.910 ;
        RECT 23.140 177.570 23.400 177.890 ;
        RECT 23.200 176.530 23.340 177.570 ;
        RECT 23.140 176.210 23.400 176.530 ;
        RECT 18.540 175.870 18.800 176.190 ;
        RECT 22.220 174.850 22.480 175.170 ;
        RECT 22.280 161.820 22.420 174.850 ;
        RECT 25.960 170.750 26.100 177.910 ;
        RECT 27.800 177.830 28.860 177.970 ;
        RECT 28.720 177.550 28.860 177.830 ;
        RECT 28.660 177.230 28.920 177.550 ;
        RECT 28.720 175.170 28.860 177.230 ;
        RECT 28.660 174.850 28.920 175.170 ;
        RECT 28.930 173.975 30.470 174.345 ;
        RECT 30.500 173.490 30.760 173.810 ;
        RECT 28.660 173.150 28.920 173.470 ;
        RECT 27.740 172.130 28.000 172.450 ;
        RECT 25.900 170.430 26.160 170.750 ;
        RECT 22.680 170.090 22.940 170.410 ;
        RECT 22.740 168.370 22.880 170.090 ;
        RECT 27.280 169.070 27.540 169.390 ;
        RECT 22.680 168.050 22.940 168.370 ;
        RECT 27.340 167.350 27.480 169.070 ;
        RECT 27.280 167.030 27.540 167.350 ;
        RECT 27.800 166.670 27.940 172.130 ;
        RECT 28.720 169.300 28.860 173.150 ;
        RECT 30.040 172.810 30.300 173.130 ;
        RECT 29.580 172.470 29.840 172.790 ;
        RECT 29.640 170.410 29.780 172.470 ;
        RECT 30.100 170.410 30.240 172.810 ;
        RECT 30.560 171.090 30.700 173.490 ;
        RECT 31.480 172.790 31.620 179.950 ;
        RECT 32.230 176.695 33.770 177.065 ;
        RECT 31.420 172.470 31.680 172.790 ;
        RECT 30.960 171.790 31.220 172.110 ;
        RECT 31.880 171.790 32.140 172.110 ;
        RECT 31.020 171.170 31.160 171.790 ;
        RECT 30.500 170.770 30.760 171.090 ;
        RECT 31.020 171.030 31.620 171.170 ;
        RECT 30.960 170.430 31.220 170.750 ;
        RECT 29.580 170.090 29.840 170.410 ;
        RECT 30.040 170.090 30.300 170.410 ;
        RECT 29.640 169.390 29.780 170.090 ;
        RECT 28.260 169.160 28.860 169.300 ;
        RECT 28.260 168.030 28.400 169.160 ;
        RECT 29.580 169.070 29.840 169.390 ;
        RECT 28.930 168.535 30.470 168.905 ;
        RECT 28.200 167.770 28.460 168.030 ;
        RECT 28.200 167.710 28.860 167.770 ;
        RECT 28.260 167.630 28.860 167.710 ;
        RECT 25.440 166.350 25.700 166.670 ;
        RECT 27.740 166.350 28.000 166.670 ;
        RECT 28.200 166.350 28.460 166.670 ;
        RECT 22.680 161.820 22.940 161.910 ;
        RECT 22.280 161.680 22.940 161.820 ;
        RECT 22.680 161.590 22.940 161.680 ;
        RECT 22.740 154.430 22.880 161.590 ;
        RECT 23.600 155.470 23.860 155.790 ;
        RECT 22.680 154.110 22.940 154.430 ;
        RECT 19.000 150.710 19.260 151.030 ;
        RECT 19.060 140.490 19.200 150.710 ;
        RECT 20.380 150.370 20.640 150.690 ;
        RECT 20.440 149.330 20.580 150.370 ;
        RECT 22.740 149.330 22.880 154.110 ;
        RECT 23.660 153.070 23.800 155.470 ;
        RECT 23.600 152.750 23.860 153.070 ;
        RECT 20.380 149.010 20.640 149.330 ;
        RECT 22.680 149.010 22.940 149.330 ;
        RECT 19.000 140.170 19.260 140.490 ;
        RECT 21.300 139.490 21.560 139.810 ;
        RECT 21.360 138.450 21.500 139.490 ;
        RECT 22.740 139.470 22.880 149.010 ;
        RECT 24.060 147.650 24.320 147.970 ;
        RECT 24.120 143.210 24.260 147.650 ;
        RECT 24.060 142.890 24.320 143.210 ;
        RECT 23.140 139.830 23.400 140.150 ;
        RECT 22.680 139.150 22.940 139.470 ;
        RECT 22.740 138.450 22.880 139.150 ;
        RECT 21.300 138.130 21.560 138.450 ;
        RECT 22.680 138.130 22.940 138.450 ;
        RECT 12.100 136.605 12.360 136.750 ;
        RECT 12.090 136.235 12.370 136.605 ;
        RECT 23.200 121.450 23.340 139.830 ;
        RECT 25.500 139.810 25.640 166.350 ;
        RECT 28.260 165.050 28.400 166.350 ;
        RECT 28.720 165.310 28.860 167.630 ;
        RECT 31.020 167.350 31.160 170.430 ;
        RECT 29.120 167.030 29.380 167.350 ;
        RECT 30.960 167.030 31.220 167.350 ;
        RECT 29.180 165.650 29.320 167.030 ;
        RECT 29.580 166.690 29.840 167.010 ;
        RECT 29.120 165.330 29.380 165.650 ;
        RECT 27.800 164.970 28.400 165.050 ;
        RECT 28.660 164.990 28.920 165.310 ;
        RECT 29.640 164.970 29.780 166.690 ;
        RECT 27.740 164.910 28.400 164.970 ;
        RECT 27.740 164.650 28.000 164.910 ;
        RECT 29.580 164.650 29.840 164.970 ;
        RECT 31.020 164.630 31.160 167.030 ;
        RECT 30.960 164.310 31.220 164.630 ;
        RECT 25.900 163.630 26.160 163.950 ;
        RECT 26.360 163.630 26.620 163.950 ;
        RECT 25.960 162.930 26.100 163.630 ;
        RECT 25.900 162.610 26.160 162.930 ;
        RECT 26.420 162.590 26.560 163.630 ;
        RECT 28.930 163.095 30.470 163.465 ;
        RECT 26.360 162.270 26.620 162.590 ;
        RECT 26.420 156.810 26.560 162.270 ;
        RECT 29.580 160.910 29.840 161.230 ;
        RECT 29.640 159.870 29.780 160.910 ;
        RECT 29.580 159.550 29.840 159.870 ;
        RECT 31.020 159.610 31.160 164.310 ;
        RECT 31.480 162.930 31.620 171.030 ;
        RECT 31.940 170.320 32.080 171.790 ;
        RECT 32.230 171.255 33.770 171.625 ;
        RECT 32.340 170.320 32.600 170.410 ;
        RECT 31.940 170.180 32.600 170.320 ;
        RECT 32.340 170.090 32.600 170.180 ;
        RECT 31.880 169.070 32.140 169.390 ;
        RECT 31.940 167.690 32.080 169.070 ;
        RECT 31.880 167.370 32.140 167.690 ;
        RECT 31.940 165.050 32.080 167.370 ;
        RECT 32.230 165.815 33.770 166.185 ;
        RECT 33.720 165.330 33.980 165.650 ;
        RECT 31.940 164.910 32.540 165.050 ;
        RECT 31.880 163.970 32.140 164.290 ;
        RECT 31.420 162.610 31.680 162.930 ;
        RECT 31.940 162.330 32.080 163.970 ;
        RECT 31.480 162.190 32.080 162.330 ;
        RECT 31.480 160.210 31.620 162.190 ;
        RECT 32.400 161.910 32.540 164.910 ;
        RECT 32.800 163.630 33.060 163.950 ;
        RECT 32.860 161.910 33.000 163.630 ;
        RECT 33.780 162.590 33.920 165.330 ;
        RECT 34.180 164.650 34.440 164.970 ;
        RECT 33.720 162.270 33.980 162.590 ;
        RECT 32.340 161.590 32.600 161.910 ;
        RECT 32.800 161.590 33.060 161.910 ;
        RECT 31.880 161.250 32.140 161.570 ;
        RECT 31.940 160.210 32.080 161.250 ;
        RECT 32.230 160.375 33.770 160.745 ;
        RECT 31.420 159.890 31.680 160.210 ;
        RECT 31.880 159.890 32.140 160.210 ;
        RECT 31.020 159.470 31.620 159.610 ;
        RECT 31.480 159.190 31.620 159.470 ;
        RECT 33.720 159.210 33.980 159.530 ;
        RECT 31.420 158.870 31.680 159.190 ;
        RECT 28.930 157.655 30.470 158.025 ;
        RECT 26.360 156.490 26.620 156.810 ;
        RECT 26.420 154.430 26.560 156.490 ;
        RECT 27.280 156.150 27.540 156.470 ;
        RECT 27.340 154.770 27.480 156.150 ;
        RECT 27.280 154.450 27.540 154.770 ;
        RECT 26.360 154.110 26.620 154.430 ;
        RECT 26.420 151.370 26.560 154.110 ;
        RECT 26.360 151.050 26.620 151.370 ;
        RECT 25.900 150.030 26.160 150.350 ;
        RECT 25.960 148.990 26.100 150.030 ;
        RECT 26.420 149.330 26.560 151.050 ;
        RECT 27.340 150.350 27.480 154.450 ;
        RECT 31.480 154.430 31.620 158.870 ;
        RECT 33.780 156.810 33.920 159.210 ;
        RECT 33.720 156.490 33.980 156.810 ;
        RECT 31.880 155.470 32.140 155.790 ;
        RECT 31.420 154.110 31.680 154.430 ;
        RECT 28.930 152.215 30.470 152.585 ;
        RECT 31.420 151.050 31.680 151.370 ;
        RECT 26.820 150.030 27.080 150.350 ;
        RECT 27.280 150.030 27.540 150.350 ;
        RECT 26.360 149.010 26.620 149.330 ;
        RECT 25.900 148.670 26.160 148.990 ;
        RECT 26.880 147.970 27.020 150.030 ;
        RECT 26.820 147.650 27.080 147.970 ;
        RECT 27.340 147.630 27.480 150.030 ;
        RECT 31.480 149.330 31.620 151.050 ;
        RECT 31.420 149.010 31.680 149.330 ;
        RECT 31.940 149.240 32.080 155.470 ;
        RECT 32.230 154.935 33.770 155.305 ;
        RECT 32.230 149.495 33.770 149.865 ;
        RECT 31.940 149.100 32.540 149.240 ;
        RECT 27.280 147.310 27.540 147.630 ;
        RECT 28.930 146.775 30.470 147.145 ;
        RECT 29.120 145.950 29.380 146.270 ;
        RECT 27.740 145.610 28.000 145.930 ;
        RECT 26.360 144.590 26.620 144.910 ;
        RECT 25.900 143.570 26.160 143.890 ;
        RECT 25.440 139.490 25.700 139.810 ;
        RECT 25.500 133.010 25.640 139.490 ;
        RECT 25.960 138.110 26.100 143.570 ;
        RECT 26.420 142.530 26.560 144.590 ;
        RECT 27.800 143.290 27.940 145.610 ;
        RECT 29.180 145.590 29.320 145.950 ;
        RECT 31.480 145.590 31.620 149.010 ;
        RECT 32.400 148.650 32.540 149.100 ;
        RECT 31.880 148.330 32.140 148.650 ;
        RECT 32.340 148.330 32.600 148.650 ;
        RECT 31.940 146.610 32.080 148.330 ;
        RECT 31.880 146.290 32.140 146.610 ;
        RECT 28.200 145.270 28.460 145.590 ;
        RECT 29.120 145.270 29.380 145.590 ;
        RECT 29.580 145.270 29.840 145.590 ;
        RECT 31.420 145.270 31.680 145.590 ;
        RECT 28.260 143.890 28.400 145.270 ;
        RECT 28.200 143.570 28.460 143.890 ;
        RECT 29.180 143.550 29.320 145.270 ;
        RECT 27.340 143.210 27.940 143.290 ;
        RECT 29.120 143.230 29.380 143.550 ;
        RECT 29.640 143.210 29.780 145.270 ;
        RECT 31.880 144.590 32.140 144.910 ;
        RECT 27.280 143.150 27.940 143.210 ;
        RECT 27.280 142.890 27.540 143.150 ;
        RECT 26.820 142.550 27.080 142.870 ;
        RECT 26.360 142.210 26.620 142.530 ;
        RECT 25.900 137.790 26.160 138.110 ;
        RECT 26.420 137.090 26.560 142.210 ;
        RECT 26.880 137.770 27.020 142.550 ;
        RECT 27.800 142.190 27.940 143.150 ;
        RECT 29.580 142.890 29.840 143.210 ;
        RECT 30.960 142.550 31.220 142.870 ;
        RECT 27.280 141.870 27.540 142.190 ;
        RECT 27.740 141.870 28.000 142.190 ;
        RECT 26.820 137.450 27.080 137.770 ;
        RECT 26.360 136.770 26.620 137.090 ;
        RECT 27.340 136.750 27.480 141.870 ;
        RECT 27.800 141.170 27.940 141.870 ;
        RECT 28.930 141.335 30.470 141.705 ;
        RECT 27.740 140.850 28.000 141.170 ;
        RECT 28.200 140.510 28.460 140.830 ;
        RECT 28.260 139.470 28.400 140.510 ;
        RECT 31.020 140.150 31.160 142.550 ;
        RECT 31.420 141.870 31.680 142.190 ;
        RECT 30.960 139.830 31.220 140.150 ;
        RECT 28.200 139.150 28.460 139.470 ;
        RECT 28.260 138.110 28.400 139.150 ;
        RECT 28.200 137.790 28.460 138.110 ;
        RECT 31.020 137.770 31.160 139.830 ;
        RECT 30.960 137.450 31.220 137.770 ;
        RECT 28.200 137.110 28.460 137.430 ;
        RECT 27.280 136.430 27.540 136.750 ;
        RECT 28.260 135.130 28.400 137.110 ;
        RECT 28.930 135.895 30.470 136.265 ;
        RECT 28.260 134.990 28.860 135.130 ;
        RECT 25.440 132.690 25.700 133.010 ;
        RECT 28.720 131.730 28.860 134.990 ;
        RECT 31.020 134.710 31.160 137.450 ;
        RECT 30.960 134.390 31.220 134.710 ;
        RECT 31.480 134.450 31.620 141.870 ;
        RECT 31.940 139.470 32.080 144.590 ;
        RECT 32.230 144.055 33.770 144.425 ;
        RECT 34.240 143.550 34.380 164.650 ;
        RECT 34.700 162.250 34.840 179.950 ;
        RECT 36.540 179.250 36.680 180.970 ;
        RECT 36.480 178.930 36.740 179.250 ;
        RECT 37.460 178.910 37.600 183.350 ;
        RECT 37.860 180.630 38.120 180.950 ;
        RECT 37.920 179.250 38.060 180.630 ;
        RECT 37.860 178.930 38.120 179.250 ;
        RECT 37.400 178.590 37.660 178.910 ;
        RECT 38.380 178.230 38.520 186.410 ;
        RECT 42.520 184.010 42.660 190.830 ;
        RECT 42.980 189.110 43.120 192.190 ;
        RECT 45.740 192.170 45.880 193.550 ;
        RECT 46.200 192.850 46.340 193.550 ;
        RECT 46.140 192.530 46.400 192.850 ;
        RECT 46.130 192.250 46.410 192.365 ;
        RECT 46.660 192.250 46.800 195.250 ;
        RECT 48.440 194.230 48.700 194.550 ;
        RECT 47.060 193.550 47.320 193.870 ;
        RECT 47.120 192.510 47.260 193.550 ;
        RECT 48.500 192.850 48.640 194.230 ;
        RECT 48.960 194.210 49.100 197.290 ;
        RECT 49.360 196.270 49.620 196.590 ;
        RECT 48.900 193.890 49.160 194.210 ;
        RECT 48.440 192.530 48.700 192.850 ;
        RECT 45.680 191.850 45.940 192.170 ;
        RECT 46.130 192.110 46.800 192.250 ;
        RECT 47.060 192.190 47.320 192.510 ;
        RECT 46.130 191.995 46.410 192.110 ;
        RECT 46.140 191.850 46.400 191.995 ;
        RECT 42.920 188.790 43.180 189.110 ;
        RECT 42.920 188.110 43.180 188.430 ;
        RECT 42.980 184.690 43.120 188.110 ;
        RECT 44.300 185.450 44.560 185.710 ;
        RECT 43.900 185.390 44.560 185.450 ;
        RECT 43.900 185.310 44.500 185.390 ;
        RECT 42.920 184.370 43.180 184.690 ;
        RECT 42.460 183.690 42.720 184.010 ;
        RECT 41.540 180.970 41.800 181.290 ;
        RECT 38.320 177.910 38.580 178.230 ;
        RECT 35.560 177.570 35.820 177.890 ;
        RECT 35.100 172.130 35.360 172.450 ;
        RECT 35.160 164.630 35.300 172.130 ;
        RECT 35.620 167.350 35.760 177.570 ;
        RECT 37.400 173.490 37.660 173.810 ;
        RECT 37.460 169.390 37.600 173.490 ;
        RECT 38.380 173.130 38.520 177.910 ;
        RECT 41.600 177.890 41.740 180.970 ;
        RECT 42.000 178.590 42.260 178.910 ;
        RECT 41.540 177.570 41.800 177.890 ;
        RECT 38.320 172.810 38.580 173.130 ;
        RECT 38.380 170.750 38.520 172.810 ;
        RECT 38.320 170.430 38.580 170.750 ;
        RECT 37.400 169.070 37.660 169.390 ;
        RECT 35.560 167.030 35.820 167.350 ;
        RECT 35.100 164.310 35.360 164.630 ;
        RECT 35.100 162.270 35.360 162.590 ;
        RECT 34.640 161.930 34.900 162.250 ;
        RECT 34.640 161.250 34.900 161.570 ;
        RECT 34.700 156.470 34.840 161.250 ;
        RECT 34.640 156.150 34.900 156.470 ;
        RECT 34.640 154.450 34.900 154.770 ;
        RECT 34.700 150.350 34.840 154.450 ;
        RECT 34.640 150.030 34.900 150.350 ;
        RECT 34.640 148.330 34.900 148.650 ;
        RECT 34.700 146.270 34.840 148.330 ;
        RECT 35.160 148.310 35.300 162.270 ;
        RECT 35.620 161.570 35.760 167.030 ;
        RECT 36.940 166.410 37.200 166.670 ;
        RECT 37.460 166.410 37.600 169.070 ;
        RECT 38.380 167.350 38.520 170.430 ;
        RECT 42.060 170.410 42.200 178.590 ;
        RECT 42.520 172.700 42.660 183.690 ;
        RECT 43.900 183.670 44.040 185.310 ;
        RECT 43.840 183.350 44.100 183.670 ;
        RECT 43.380 183.010 43.640 183.330 ;
        RECT 42.920 172.700 43.180 172.790 ;
        RECT 42.520 172.560 43.180 172.700 ;
        RECT 42.920 172.470 43.180 172.560 ;
        RECT 42.460 171.790 42.720 172.110 ;
        RECT 43.440 171.850 43.580 183.010 ;
        RECT 43.900 181.290 44.040 183.350 ;
        RECT 45.220 182.670 45.480 182.990 ;
        RECT 45.280 181.290 45.420 182.670 ;
        RECT 43.840 180.970 44.100 181.290 ;
        RECT 45.220 180.970 45.480 181.290 ;
        RECT 45.740 178.230 45.880 191.850 ;
        RECT 48.960 186.050 49.100 193.890 ;
        RECT 49.420 193.870 49.560 196.270 ;
        RECT 51.260 195.570 51.400 200.690 ;
        RECT 62.760 199.990 62.900 208.800 ;
        RECT 72.420 199.990 72.560 208.800 ;
        RECT 110.010 206.150 110.150 218.060 ;
        RECT 111.010 206.600 111.150 218.690 ;
        RECT 110.920 206.340 111.240 206.600 ;
        RECT 109.920 205.890 110.240 206.150 ;
        RECT 111.420 206.120 111.560 219.040 ;
        RECT 111.330 205.860 111.650 206.120 ;
        RECT 101.480 205.335 105.480 205.405 ;
        RECT 111.810 205.335 111.950 219.350 ;
        RECT 121.210 218.215 121.530 218.275 ;
        RECT 125.435 218.215 125.805 218.285 ;
        RECT 121.210 218.075 125.805 218.215 ;
        RECT 121.210 218.015 121.530 218.075 ;
        RECT 125.435 218.005 125.805 218.075 ;
        RECT 128.010 218.215 128.330 218.275 ;
        RECT 132.235 218.215 132.605 218.285 ;
        RECT 139.035 218.275 139.405 218.285 ;
        RECT 128.010 218.075 132.605 218.215 ;
        RECT 128.010 218.015 128.330 218.075 ;
        RECT 132.235 218.005 132.605 218.075 ;
        RECT 138.890 218.015 139.405 218.275 ;
        RECT 139.035 218.005 139.405 218.015 ;
        RECT 116.450 217.755 116.770 217.815 ;
        RECT 119.850 217.755 120.170 217.815 ;
        RECT 121.550 217.755 121.870 217.815 ;
        RECT 116.450 217.615 121.870 217.755 ;
        RECT 116.450 217.555 116.770 217.615 ;
        RECT 119.850 217.555 120.170 217.615 ;
        RECT 121.550 217.555 121.870 217.615 ;
        RECT 124.610 217.755 124.930 217.815 ;
        RECT 126.650 217.755 126.970 217.815 ;
        RECT 124.610 217.615 126.970 217.755 ;
        RECT 124.610 217.555 124.930 217.615 ;
        RECT 126.650 217.555 126.970 217.615 ;
        RECT 127.330 217.755 127.650 217.815 ;
        RECT 130.050 217.755 130.370 217.815 ;
        RECT 131.750 217.755 132.070 217.815 ;
        RECT 127.330 217.615 132.070 217.755 ;
        RECT 127.330 217.555 127.650 217.615 ;
        RECT 130.050 217.555 130.370 217.615 ;
        RECT 131.750 217.555 132.070 217.615 ;
        RECT 133.110 217.755 133.430 217.815 ;
        RECT 134.470 217.755 134.790 217.815 ;
        RECT 133.110 217.615 134.790 217.755 ;
        RECT 133.110 217.555 133.430 217.615 ;
        RECT 134.470 217.555 134.790 217.615 ;
        RECT 138.890 215.915 139.210 215.975 ;
        RECT 140.250 215.915 140.570 215.975 ;
        RECT 138.890 215.775 140.570 215.915 ;
        RECT 138.890 215.715 139.210 215.775 ;
        RECT 140.250 215.715 140.570 215.775 ;
        RECT 123.930 215.455 124.250 215.515 ;
        RECT 126.310 215.455 126.630 215.515 ;
        RECT 123.930 215.315 126.630 215.455 ;
        RECT 123.930 215.255 124.250 215.315 ;
        RECT 126.310 215.255 126.630 215.315 ;
        RECT 135.490 215.455 135.810 215.515 ;
        RECT 137.530 215.455 137.850 215.515 ;
        RECT 135.490 215.315 137.850 215.455 ;
        RECT 135.490 215.255 135.810 215.315 ;
        RECT 137.530 215.255 137.850 215.315 ;
        RECT 117.130 214.995 117.450 215.055 ;
        RECT 118.490 214.995 118.810 215.055 ;
        RECT 117.130 214.855 118.810 214.995 ;
        RECT 117.130 214.795 117.450 214.855 ;
        RECT 118.490 214.795 118.810 214.855 ;
        RECT 144.330 213.615 144.650 213.675 ;
        RECT 146.030 213.615 146.350 213.675 ;
        RECT 144.330 213.475 146.350 213.615 ;
        RECT 144.330 213.415 144.650 213.475 ;
        RECT 146.030 213.415 146.350 213.475 ;
        RECT 117.130 213.155 117.450 213.215 ;
        RECT 120.870 213.155 121.190 213.215 ;
        RECT 117.130 213.015 121.190 213.155 ;
        RECT 117.130 212.955 117.450 213.015 ;
        RECT 120.870 212.955 121.190 213.015 ;
        RECT 130.730 213.155 131.050 213.215 ;
        RECT 134.470 213.155 134.790 213.215 ;
        RECT 130.730 213.015 134.790 213.155 ;
        RECT 130.730 212.955 131.050 213.015 ;
        RECT 134.470 212.955 134.790 213.015 ;
        RECT 117.130 212.695 117.450 212.755 ;
        RECT 121.210 212.695 121.530 212.755 ;
        RECT 126.990 212.695 127.310 212.755 ;
        RECT 117.130 212.555 127.310 212.695 ;
        RECT 117.130 212.495 117.450 212.555 ;
        RECT 121.210 212.495 121.530 212.555 ;
        RECT 126.990 212.495 127.310 212.555 ;
        RECT 128.010 212.695 128.330 212.755 ;
        RECT 129.030 212.695 129.350 212.755 ;
        RECT 128.010 212.555 129.350 212.695 ;
        RECT 128.010 212.495 128.330 212.555 ;
        RECT 129.030 212.495 129.350 212.555 ;
        RECT 126.990 212.235 127.310 212.295 ;
        RECT 134.810 212.235 135.130 212.295 ;
        RECT 137.870 212.235 138.190 212.295 ;
        RECT 126.990 212.095 138.190 212.235 ;
        RECT 126.990 212.035 127.310 212.095 ;
        RECT 134.810 212.035 135.130 212.095 ;
        RECT 137.870 212.035 138.190 212.095 ;
        RECT 119.170 210.855 119.490 210.915 ;
        RECT 124.270 210.855 124.590 210.915 ;
        RECT 119.170 210.715 124.590 210.855 ;
        RECT 119.170 210.655 119.490 210.715 ;
        RECT 124.270 210.655 124.590 210.715 ;
        RECT 132.770 210.855 133.090 210.915 ;
        RECT 135.150 210.855 135.470 210.915 ;
        RECT 132.770 210.715 135.470 210.855 ;
        RECT 132.770 210.655 133.090 210.715 ;
        RECT 135.150 210.655 135.470 210.715 ;
        RECT 138.210 210.855 138.530 210.915 ;
        RECT 139.910 210.855 140.230 210.915 ;
        RECT 138.210 210.715 140.230 210.855 ;
        RECT 138.210 210.655 138.530 210.715 ;
        RECT 139.910 210.655 140.230 210.715 ;
        RECT 117.130 210.395 117.450 210.455 ;
        RECT 121.550 210.395 121.870 210.455 ;
        RECT 117.130 210.255 121.870 210.395 ;
        RECT 117.130 210.195 117.450 210.255 ;
        RECT 121.550 210.195 121.870 210.255 ;
        RECT 138.890 210.395 139.210 210.455 ;
        RECT 139.910 210.395 140.230 210.455 ;
        RECT 138.890 210.255 140.230 210.395 ;
        RECT 138.890 210.195 139.210 210.255 ;
        RECT 139.910 210.195 140.230 210.255 ;
        RECT 121.890 209.935 122.210 209.995 ;
        RECT 125.290 209.935 125.610 209.995 ;
        RECT 129.710 209.935 130.030 209.995 ;
        RECT 121.890 209.795 130.030 209.935 ;
        RECT 121.890 209.735 122.210 209.795 ;
        RECT 125.290 209.735 125.610 209.795 ;
        RECT 129.710 209.735 130.030 209.795 ;
        RECT 144.330 209.015 144.650 209.075 ;
        RECT 146.030 209.015 146.350 209.075 ;
        RECT 144.330 208.875 146.350 209.015 ;
        RECT 144.330 208.815 144.650 208.875 ;
        RECT 146.030 208.815 146.350 208.875 ;
        RECT 143.795 208.555 144.165 208.625 ;
        RECT 146.030 208.555 146.350 208.615 ;
        RECT 143.795 208.415 146.350 208.555 ;
        RECT 143.795 208.345 144.165 208.415 ;
        RECT 146.030 208.355 146.350 208.415 ;
        RECT 113.390 208.095 113.710 208.155 ;
        RECT 117.130 208.095 117.450 208.155 ;
        RECT 113.390 207.955 117.450 208.095 ;
        RECT 113.390 207.895 113.710 207.955 ;
        RECT 117.130 207.895 117.450 207.955 ;
        RECT 135.150 208.095 135.470 208.155 ;
        RECT 138.890 208.095 139.210 208.155 ;
        RECT 140.590 208.095 140.910 208.155 ;
        RECT 142.630 208.095 142.950 208.155 ;
        RECT 135.150 207.955 142.950 208.095 ;
        RECT 135.150 207.895 135.470 207.955 ;
        RECT 138.890 207.895 139.210 207.955 ;
        RECT 140.590 207.895 140.910 207.955 ;
        RECT 142.630 207.895 142.950 207.955 ;
        RECT 133.110 207.175 133.430 207.235 ;
        RECT 142.435 207.175 142.805 207.245 ;
        RECT 133.110 207.035 142.805 207.175 ;
        RECT 133.110 206.975 133.430 207.035 ;
        RECT 142.435 206.965 142.805 207.035 ;
        RECT 143.990 206.715 144.310 206.775 ;
        RECT 145.350 206.715 145.670 206.775 ;
        RECT 143.990 206.575 145.670 206.715 ;
        RECT 143.990 206.515 144.310 206.575 ;
        RECT 145.350 206.515 145.670 206.575 ;
        RECT 116.110 206.255 116.430 206.315 ;
        RECT 121.550 206.255 121.870 206.315 ;
        RECT 127.670 206.255 127.990 206.315 ;
        RECT 116.110 206.115 127.990 206.255 ;
        RECT 116.110 206.055 116.430 206.115 ;
        RECT 121.550 206.055 121.870 206.115 ;
        RECT 127.670 206.055 127.990 206.115 ;
        RECT 135.490 205.795 135.810 205.855 ;
        RECT 138.890 205.795 139.210 205.855 ;
        RECT 135.490 205.655 139.210 205.795 ;
        RECT 135.490 205.595 135.810 205.655 ;
        RECT 138.890 205.595 139.210 205.655 ;
        RECT 141.610 205.795 141.930 205.855 ;
        RECT 143.650 205.795 143.970 205.855 ;
        RECT 141.610 205.655 143.970 205.795 ;
        RECT 141.610 205.595 141.930 205.655 ;
        RECT 143.650 205.595 143.970 205.655 ;
        RECT 112.710 205.335 113.030 205.395 ;
        RECT 101.480 205.195 113.030 205.335 ;
        RECT 101.480 205.125 105.480 205.195 ;
        RECT 112.710 205.135 113.030 205.195 ;
        RECT 147.050 205.335 147.370 205.395 ;
        RECT 149.680 205.335 150.000 205.430 ;
        RECT 155.245 205.335 159.245 205.405 ;
        RECT 147.050 205.195 159.245 205.335 ;
        RECT 147.050 205.135 147.370 205.195 ;
        RECT 149.680 205.100 150.000 205.195 ;
        RECT 155.245 205.125 159.245 205.195 ;
        RECT 123.930 204.875 124.250 204.935 ;
        RECT 126.650 204.875 126.970 204.935 ;
        RECT 123.930 204.735 126.970 204.875 ;
        RECT 123.930 204.675 124.250 204.735 ;
        RECT 126.650 204.675 126.970 204.735 ;
        RECT 127.670 204.875 127.990 204.935 ;
        RECT 130.730 204.875 131.050 204.935 ;
        RECT 136.170 204.875 136.490 204.935 ;
        RECT 138.890 204.875 139.210 204.935 ;
        RECT 127.670 204.735 139.210 204.875 ;
        RECT 127.670 204.675 127.990 204.735 ;
        RECT 130.730 204.675 131.050 204.735 ;
        RECT 136.170 204.675 136.490 204.735 ;
        RECT 138.890 204.675 139.210 204.735 ;
        RECT 128.010 204.415 128.330 204.475 ;
        RECT 129.710 204.415 130.030 204.475 ;
        RECT 128.010 204.275 130.030 204.415 ;
        RECT 128.010 204.215 128.330 204.275 ;
        RECT 129.710 204.215 130.030 204.275 ;
        RECT 130.730 204.415 131.050 204.475 ;
        RECT 143.795 204.415 144.165 204.485 ;
        RECT 130.730 204.275 144.165 204.415 ;
        RECT 130.730 204.215 131.050 204.275 ;
        RECT 143.795 204.205 144.165 204.275 ;
        RECT 113.390 202.835 113.710 203.095 ;
        RECT 111.360 202.575 111.620 202.665 ;
        RECT 112.710 202.575 113.030 202.635 ;
        RECT 107.190 202.435 113.030 202.575 ;
        RECT 101.480 202.115 105.480 202.185 ;
        RECT 107.190 202.115 107.330 202.435 ;
        RECT 111.360 202.345 111.620 202.435 ;
        RECT 112.710 202.375 113.030 202.435 ;
        RECT 101.480 201.975 107.330 202.115 ;
        RECT 101.480 201.905 105.480 201.975 ;
        RECT 113.480 201.655 113.620 202.835 ;
        RECT 114.895 202.205 115.265 203.745 ;
        RECT 120.335 202.205 120.705 203.745 ;
        RECT 125.775 202.205 126.145 203.745 ;
        RECT 131.215 202.205 131.585 203.745 ;
        RECT 136.655 202.205 137.025 203.745 ;
        RECT 142.095 202.205 142.465 203.745 ;
        RECT 147.535 202.205 147.905 203.745 ;
        RECT 155.245 202.115 159.245 202.185 ;
        RECT 148.670 201.975 159.245 202.115 ;
        RECT 117.130 201.655 117.450 201.715 ;
        RECT 120.870 201.655 121.190 201.715 ;
        RECT 113.480 201.515 116.850 201.655 ;
        RECT 116.710 200.795 116.850 201.515 ;
        RECT 117.130 201.515 121.190 201.655 ;
        RECT 117.130 201.455 117.450 201.515 ;
        RECT 120.870 201.455 121.190 201.515 ;
        RECT 129.710 201.655 130.030 201.715 ;
        RECT 139.910 201.655 140.230 201.715 ;
        RECT 129.710 201.515 140.230 201.655 ;
        RECT 129.710 201.455 130.030 201.515 ;
        RECT 139.910 201.455 140.230 201.515 ;
        RECT 140.590 201.655 140.910 201.715 ;
        RECT 145.350 201.655 145.670 201.715 ;
        RECT 140.590 201.515 145.670 201.655 ;
        RECT 140.590 201.455 140.910 201.515 ;
        RECT 145.350 201.455 145.670 201.515 ;
        RECT 118.830 201.195 119.150 201.255 ;
        RECT 131.750 201.195 132.070 201.255 ;
        RECT 138.210 201.195 138.530 201.255 ;
        RECT 118.830 201.055 138.530 201.195 ;
        RECT 118.830 200.995 119.150 201.055 ;
        RECT 131.750 200.995 132.070 201.055 ;
        RECT 138.210 200.995 138.530 201.055 ;
        RECT 138.890 201.195 139.210 201.255 ;
        RECT 140.590 201.195 140.910 201.255 ;
        RECT 138.890 201.055 140.910 201.195 ;
        RECT 138.890 200.995 139.210 201.055 ;
        RECT 140.590 200.995 140.910 201.055 ;
        RECT 142.970 201.195 143.290 201.255 ;
        RECT 148.110 201.195 148.440 201.290 ;
        RECT 148.670 201.195 148.810 201.975 ;
        RECT 155.245 201.905 159.245 201.975 ;
        RECT 142.970 201.055 148.810 201.195 ;
        RECT 142.970 200.995 143.290 201.055 ;
        RECT 148.110 200.960 148.440 201.055 ;
        RECT 113.050 200.735 113.370 200.795 ;
        RECT 115.430 200.735 115.750 200.795 ;
        RECT 113.050 200.595 115.750 200.735 ;
        RECT 116.710 200.735 117.110 200.795 ;
        RECT 119.850 200.735 120.170 200.795 ;
        RECT 121.890 200.735 122.210 200.795 ;
        RECT 123.590 200.735 123.910 200.795 ;
        RECT 116.710 200.595 123.910 200.735 ;
        RECT 113.050 200.535 113.370 200.595 ;
        RECT 115.430 200.535 115.750 200.595 ;
        RECT 116.790 200.535 117.110 200.595 ;
        RECT 119.850 200.535 120.170 200.595 ;
        RECT 121.890 200.535 122.210 200.595 ;
        RECT 123.590 200.535 123.910 200.595 ;
        RECT 129.710 200.735 130.030 200.795 ;
        RECT 132.430 200.735 132.750 200.795 ;
        RECT 137.190 200.735 137.510 200.795 ;
        RECT 129.710 200.595 132.750 200.735 ;
        RECT 129.710 200.535 130.030 200.595 ;
        RECT 132.430 200.535 132.750 200.595 ;
        RECT 133.030 200.595 137.510 200.735 ;
        RECT 62.700 199.670 62.960 199.990 ;
        RECT 72.360 199.670 72.620 199.990 ;
        RECT 58.100 198.990 58.360 199.310 ;
        RECT 61.780 198.990 62.040 199.310 ;
        RECT 64.540 198.990 64.800 199.310 ;
        RECT 70.980 198.990 71.240 199.310 ;
        RECT 58.160 198.290 58.300 198.990 ;
        RECT 58.100 197.970 58.360 198.290 ;
        RECT 56.720 196.950 56.980 197.270 ;
        RECT 51.200 195.250 51.460 195.570 ;
        RECT 50.280 194.230 50.540 194.550 ;
        RECT 49.360 193.550 49.620 193.870 ;
        RECT 49.420 191.490 49.560 193.550 ;
        RECT 49.360 191.170 49.620 191.490 ;
        RECT 47.520 185.730 47.780 186.050 ;
        RECT 48.900 185.730 49.160 186.050 ;
        RECT 47.060 180.290 47.320 180.610 ;
        RECT 47.120 178.230 47.260 180.290 ;
        RECT 45.680 177.910 45.940 178.230 ;
        RECT 47.060 177.910 47.320 178.230 ;
        RECT 45.220 175.530 45.480 175.850 ;
        RECT 44.300 174.850 44.560 175.170 ;
        RECT 43.840 174.510 44.100 174.830 ;
        RECT 43.900 172.450 44.040 174.510 ;
        RECT 44.360 173.810 44.500 174.850 ;
        RECT 44.300 173.490 44.560 173.810 ;
        RECT 44.760 173.150 45.020 173.470 ;
        RECT 44.820 172.450 44.960 173.150 ;
        RECT 43.840 172.130 44.100 172.450 ;
        RECT 44.760 172.130 45.020 172.450 ;
        RECT 42.000 170.090 42.260 170.410 ;
        RECT 42.060 168.370 42.200 170.090 ;
        RECT 42.000 168.050 42.260 168.370 ;
        RECT 42.520 167.350 42.660 171.790 ;
        RECT 42.980 171.710 43.580 171.850 ;
        RECT 38.320 167.030 38.580 167.350 ;
        RECT 40.160 167.030 40.420 167.350 ;
        RECT 42.460 167.030 42.720 167.350 ;
        RECT 36.940 166.350 37.600 166.410 ;
        RECT 39.240 166.350 39.500 166.670 ;
        RECT 37.000 166.270 37.600 166.350 ;
        RECT 37.460 164.970 37.600 166.270 ;
        RECT 39.300 165.310 39.440 166.350 ;
        RECT 39.240 164.990 39.500 165.310 ;
        RECT 37.400 164.650 37.660 164.970 ;
        RECT 37.460 162.930 37.600 164.650 ;
        RECT 37.860 164.310 38.120 164.630 ;
        RECT 37.400 162.610 37.660 162.930 ;
        RECT 37.460 162.250 37.600 162.610 ;
        RECT 37.400 161.930 37.660 162.250 ;
        RECT 37.920 161.910 38.060 164.310 ;
        RECT 38.780 162.270 39.040 162.590 ;
        RECT 37.860 161.590 38.120 161.910 ;
        RECT 35.620 161.430 36.220 161.570 ;
        RECT 36.080 159.190 36.220 161.430 ;
        RECT 38.840 159.530 38.980 162.270 ;
        RECT 39.300 161.910 39.440 164.990 ;
        RECT 39.240 161.590 39.500 161.910 ;
        RECT 38.780 159.210 39.040 159.530 ;
        RECT 36.020 158.870 36.280 159.190 ;
        RECT 35.560 158.190 35.820 158.510 ;
        RECT 35.620 154.770 35.760 158.190 ;
        RECT 35.560 154.450 35.820 154.770 ;
        RECT 36.080 153.410 36.220 158.870 ;
        RECT 39.300 156.210 39.440 161.590 ;
        RECT 40.220 159.530 40.360 167.030 ;
        RECT 42.980 167.010 43.120 171.710 ;
        RECT 44.820 167.350 44.960 172.130 ;
        RECT 45.280 172.110 45.420 175.530 ;
        RECT 47.120 173.810 47.260 177.910 ;
        RECT 47.060 173.490 47.320 173.810 ;
        RECT 47.120 172.700 47.260 173.490 ;
        RECT 47.580 173.470 47.720 185.730 ;
        RECT 48.900 182.670 49.160 182.990 ;
        RECT 47.980 180.630 48.240 180.950 ;
        RECT 48.040 179.250 48.180 180.630 ;
        RECT 48.960 180.270 49.100 182.670 ;
        RECT 48.440 179.950 48.700 180.270 ;
        RECT 48.900 179.950 49.160 180.270 ;
        RECT 47.980 178.930 48.240 179.250 ;
        RECT 48.500 178.570 48.640 179.950 ;
        RECT 48.440 178.250 48.700 178.570 ;
        RECT 47.520 173.150 47.780 173.470 ;
        RECT 47.980 172.700 48.240 172.790 ;
        RECT 47.120 172.560 48.240 172.700 ;
        RECT 47.980 172.470 48.240 172.560 ;
        RECT 45.220 171.790 45.480 172.110 ;
        RECT 44.760 167.030 45.020 167.350 ;
        RECT 45.280 167.010 45.420 171.790 ;
        RECT 46.140 169.410 46.400 169.730 ;
        RECT 42.920 166.690 43.180 167.010 ;
        RECT 45.220 166.690 45.480 167.010 ;
        RECT 42.980 162.930 43.120 166.690 ;
        RECT 46.200 165.650 46.340 169.410 ;
        RECT 48.040 168.370 48.180 172.470 ;
        RECT 48.500 172.110 48.640 178.250 ;
        RECT 49.420 177.890 49.560 191.170 ;
        RECT 49.820 178.930 50.080 179.250 ;
        RECT 49.360 177.570 49.620 177.890 ;
        RECT 49.880 176.530 50.020 178.930 ;
        RECT 49.820 176.210 50.080 176.530 ;
        RECT 48.900 175.530 49.160 175.850 ;
        RECT 48.960 173.810 49.100 175.530 ;
        RECT 48.900 173.490 49.160 173.810 ;
        RECT 48.440 171.790 48.700 172.110 ;
        RECT 50.340 170.410 50.480 194.230 ;
        RECT 50.740 193.550 51.000 193.870 ;
        RECT 50.800 191.830 50.940 193.550 ;
        RECT 50.740 191.510 51.000 191.830 ;
        RECT 51.260 190.130 51.400 195.250 ;
        RECT 56.780 194.550 56.920 196.950 ;
        RECT 61.840 195.570 61.980 198.990 ;
        RECT 63.160 196.270 63.420 196.590 ;
        RECT 61.780 195.250 62.040 195.570 ;
        RECT 63.220 194.550 63.360 196.270 ;
        RECT 56.720 194.230 56.980 194.550 ;
        RECT 60.860 194.230 61.120 194.550 ;
        RECT 63.160 194.230 63.420 194.550 ;
        RECT 59.480 193.550 59.740 193.870 ;
        RECT 59.540 192.850 59.680 193.550 ;
        RECT 60.920 192.850 61.060 194.230 ;
        RECT 51.660 192.530 51.920 192.850 ;
        RECT 57.640 192.530 57.900 192.850 ;
        RECT 59.480 192.530 59.740 192.850 ;
        RECT 60.860 192.530 61.120 192.850 ;
        RECT 51.720 192.365 51.860 192.530 ;
        RECT 51.650 191.995 51.930 192.365 ;
        RECT 51.660 191.850 51.920 191.995 ;
        RECT 51.200 189.810 51.460 190.130 ;
        RECT 50.740 183.010 51.000 183.330 ;
        RECT 50.800 181.970 50.940 183.010 ;
        RECT 50.740 181.650 51.000 181.970 ;
        RECT 51.260 175.170 51.400 189.810 ;
        RECT 57.700 189.110 57.840 192.530 ;
        RECT 63.220 192.170 63.360 194.230 ;
        RECT 63.160 191.850 63.420 192.170 ;
        RECT 62.240 190.830 62.500 191.150 ;
        RECT 62.300 189.790 62.440 190.830 ;
        RECT 60.860 189.470 61.120 189.790 ;
        RECT 62.240 189.470 62.500 189.790 ;
        RECT 57.180 188.790 57.440 189.110 ;
        RECT 57.640 188.790 57.900 189.110 ;
        RECT 53.040 186.750 53.300 187.070 ;
        RECT 53.100 182.990 53.240 186.750 ;
        RECT 57.240 186.390 57.380 188.790 ;
        RECT 57.700 187.410 57.840 188.790 ;
        RECT 58.100 188.110 58.360 188.430 ;
        RECT 57.640 187.090 57.900 187.410 ;
        RECT 58.160 186.730 58.300 188.110 ;
        RECT 58.100 186.410 58.360 186.730 ;
        RECT 59.940 186.410 60.200 186.730 ;
        RECT 57.180 186.070 57.440 186.390 ;
        RECT 58.160 184.690 58.300 186.410 ;
        RECT 59.020 186.070 59.280 186.390 ;
        RECT 58.100 184.370 58.360 184.690 ;
        RECT 53.500 183.350 53.760 183.670 ;
        RECT 57.640 183.350 57.900 183.670 ;
        RECT 53.040 182.670 53.300 182.990 ;
        RECT 52.580 180.630 52.840 180.950 ;
        RECT 52.640 179.250 52.780 180.630 ;
        RECT 52.580 178.930 52.840 179.250 ;
        RECT 51.200 174.850 51.460 175.170 ;
        RECT 53.100 174.830 53.240 182.670 ;
        RECT 53.560 181.970 53.700 183.350 ;
        RECT 57.700 181.970 57.840 183.350 ;
        RECT 59.080 181.970 59.220 186.070 ;
        RECT 53.500 181.650 53.760 181.970 ;
        RECT 57.640 181.650 57.900 181.970 ;
        RECT 59.020 181.650 59.280 181.970 ;
        RECT 59.480 181.310 59.740 181.630 ;
        RECT 55.340 180.970 55.600 181.290 ;
        RECT 57.640 180.970 57.900 181.290 ;
        RECT 59.020 180.970 59.280 181.290 ;
        RECT 54.420 178.590 54.680 178.910 ;
        RECT 53.960 174.850 54.220 175.170 ;
        RECT 53.040 174.510 53.300 174.830 ;
        RECT 53.100 172.790 53.240 174.510 ;
        RECT 53.040 172.470 53.300 172.790 ;
        RECT 54.020 172.450 54.160 174.850 ;
        RECT 53.960 172.130 54.220 172.450 ;
        RECT 49.360 170.090 49.620 170.410 ;
        RECT 50.280 170.090 50.540 170.410 ;
        RECT 51.200 170.090 51.460 170.410 ;
        RECT 47.980 168.050 48.240 168.370 ;
        RECT 49.420 168.030 49.560 170.090 ;
        RECT 51.260 168.370 51.400 170.090 ;
        RECT 51.660 169.070 51.920 169.390 ;
        RECT 51.200 168.050 51.460 168.370 ;
        RECT 49.360 167.710 49.620 168.030 ;
        RECT 51.720 167.350 51.860 169.070 ;
        RECT 49.360 167.090 49.620 167.350 ;
        RECT 49.360 167.030 50.940 167.090 ;
        RECT 51.660 167.030 51.920 167.350 ;
        RECT 53.040 167.090 53.300 167.350 ;
        RECT 54.020 167.090 54.160 172.130 ;
        RECT 54.480 168.370 54.620 178.590 ;
        RECT 55.400 178.230 55.540 180.970 ;
        RECT 56.260 180.630 56.520 180.950 ;
        RECT 56.720 180.630 56.980 180.950 ;
        RECT 56.320 178.230 56.460 180.630 ;
        RECT 56.780 179.250 56.920 180.630 ;
        RECT 57.180 179.950 57.440 180.270 ;
        RECT 56.720 178.930 56.980 179.250 ;
        RECT 57.240 178.650 57.380 179.950 ;
        RECT 57.700 179.250 57.840 180.970 ;
        RECT 59.080 179.250 59.220 180.970 ;
        RECT 57.640 178.930 57.900 179.250 ;
        RECT 59.020 178.930 59.280 179.250 ;
        RECT 57.240 178.570 57.840 178.650 ;
        RECT 57.240 178.510 57.900 178.570 ;
        RECT 55.340 177.910 55.600 178.230 ;
        RECT 56.260 177.910 56.520 178.230 ;
        RECT 55.400 169.390 55.540 177.910 ;
        RECT 57.240 172.790 57.380 178.510 ;
        RECT 57.640 178.250 57.900 178.510 ;
        RECT 59.540 177.890 59.680 181.310 ;
        RECT 60.000 178.910 60.140 186.410 ;
        RECT 60.400 185.390 60.660 185.710 ;
        RECT 60.460 181.290 60.600 185.390 ;
        RECT 60.920 183.670 61.060 189.470 ;
        RECT 61.780 189.020 62.040 189.110 ;
        RECT 62.300 189.020 62.440 189.470 ;
        RECT 63.220 189.110 63.360 191.850 ;
        RECT 64.080 191.510 64.340 191.830 ;
        RECT 63.620 190.830 63.880 191.150 ;
        RECT 61.780 188.880 62.440 189.020 ;
        RECT 61.780 188.790 62.040 188.880 ;
        RECT 61.780 185.390 62.040 185.710 ;
        RECT 61.840 184.350 61.980 185.390 ;
        RECT 61.780 184.030 62.040 184.350 ;
        RECT 60.860 183.525 61.120 183.670 ;
        RECT 60.850 183.155 61.130 183.525 ;
        RECT 60.860 182.670 61.120 182.990 ;
        RECT 60.920 181.290 61.060 182.670 ;
        RECT 60.400 180.970 60.660 181.290 ;
        RECT 60.860 180.970 61.120 181.290 ;
        RECT 61.840 178.910 61.980 184.030 ;
        RECT 62.300 180.610 62.440 188.880 ;
        RECT 63.160 188.790 63.420 189.110 ;
        RECT 63.680 187.070 63.820 190.830 ;
        RECT 64.140 189.110 64.280 191.510 ;
        RECT 64.080 188.790 64.340 189.110 ;
        RECT 64.140 188.430 64.280 188.790 ;
        RECT 64.080 188.110 64.340 188.430 ;
        RECT 63.620 186.750 63.880 187.070 ;
        RECT 64.140 186.730 64.280 188.110 ;
        RECT 64.080 186.410 64.340 186.730 ;
        RECT 64.600 184.090 64.740 198.990 ;
        RECT 68.220 196.270 68.480 196.590 ;
        RECT 65.460 194.230 65.720 194.550 ;
        RECT 65.520 190.130 65.660 194.230 ;
        RECT 67.300 193.890 67.560 194.210 ;
        RECT 66.380 191.170 66.640 191.490 ;
        RECT 66.440 190.130 66.580 191.170 ;
        RECT 67.360 191.150 67.500 193.890 ;
        RECT 68.280 192.170 68.420 196.270 ;
        RECT 68.680 195.480 68.940 195.570 ;
        RECT 68.680 195.340 69.340 195.480 ;
        RECT 68.680 195.250 68.940 195.340 ;
        RECT 68.680 194.230 68.940 194.550 ;
        RECT 68.220 191.850 68.480 192.170 ;
        RECT 67.300 190.830 67.560 191.150 ;
        RECT 65.460 189.810 65.720 190.130 ;
        RECT 66.380 189.810 66.640 190.130 ;
        RECT 66.440 189.450 66.580 189.810 ;
        RECT 66.380 189.130 66.640 189.450 ;
        RECT 66.440 186.390 66.580 189.130 ;
        RECT 68.280 188.770 68.420 191.850 ;
        RECT 68.740 191.490 68.880 194.230 ;
        RECT 69.200 192.850 69.340 195.340 ;
        RECT 69.600 193.550 69.860 193.870 ;
        RECT 69.140 192.530 69.400 192.850 ;
        RECT 68.680 191.170 68.940 191.490 ;
        RECT 68.220 188.450 68.480 188.770 ;
        RECT 66.380 186.070 66.640 186.390 ;
        RECT 68.680 185.730 68.940 186.050 ;
        RECT 68.740 184.690 68.880 185.730 ;
        RECT 65.000 184.370 65.260 184.690 ;
        RECT 68.680 184.370 68.940 184.690 ;
        RECT 64.140 183.950 64.740 184.090 ;
        RECT 65.060 184.010 65.200 184.370 ;
        RECT 68.220 184.030 68.480 184.350 ;
        RECT 63.620 183.525 63.880 183.670 ;
        RECT 63.610 183.155 63.890 183.525 ;
        RECT 63.160 182.670 63.420 182.990 ;
        RECT 63.220 181.630 63.360 182.670 ;
        RECT 63.160 181.310 63.420 181.630 ;
        RECT 62.700 180.860 62.960 180.950 ;
        RECT 64.140 180.860 64.280 183.950 ;
        RECT 65.000 183.690 65.260 184.010 ;
        RECT 65.460 183.350 65.720 183.670 ;
        RECT 64.540 183.010 64.800 183.330 ;
        RECT 62.700 180.720 64.280 180.860 ;
        RECT 62.700 180.630 62.960 180.720 ;
        RECT 62.240 180.290 62.500 180.610 ;
        RECT 59.940 178.590 60.200 178.910 ;
        RECT 61.780 178.590 62.040 178.910 ;
        RECT 60.400 177.910 60.660 178.230 ;
        RECT 62.300 177.970 62.440 180.290 ;
        RECT 59.020 177.570 59.280 177.890 ;
        RECT 59.480 177.570 59.740 177.890 ;
        RECT 59.940 177.570 60.200 177.890 ;
        RECT 58.100 172.810 58.360 173.130 ;
        RECT 57.180 172.470 57.440 172.790 ;
        RECT 57.640 172.470 57.900 172.790 ;
        RECT 57.700 171.090 57.840 172.470 ;
        RECT 57.640 170.770 57.900 171.090 ;
        RECT 57.640 170.090 57.900 170.410 ;
        RECT 55.340 169.070 55.600 169.390 ;
        RECT 54.420 168.050 54.680 168.370 ;
        RECT 57.180 168.050 57.440 168.370 ;
        RECT 54.880 167.710 55.140 168.030 ;
        RECT 53.040 167.030 54.160 167.090 ;
        RECT 49.420 167.010 50.940 167.030 ;
        RECT 49.420 166.950 51.000 167.010 ;
        RECT 53.100 166.950 54.160 167.030 ;
        RECT 50.740 166.690 51.000 166.950 ;
        RECT 54.020 166.670 54.160 166.950 ;
        RECT 53.500 166.350 53.760 166.670 ;
        RECT 53.960 166.350 54.220 166.670 ;
        RECT 46.140 165.330 46.400 165.650 ;
        RECT 42.920 162.610 43.180 162.930 ;
        RECT 42.920 161.930 43.180 162.250 ;
        RECT 42.460 161.590 42.720 161.910 ;
        RECT 42.000 161.250 42.260 161.570 ;
        RECT 40.620 160.910 40.880 161.230 ;
        RECT 39.700 159.210 39.960 159.530 ;
        RECT 40.160 159.210 40.420 159.530 ;
        RECT 38.840 156.070 39.440 156.210 ;
        RECT 36.020 153.090 36.280 153.410 ;
        RECT 36.940 151.050 37.200 151.370 ;
        RECT 35.560 150.030 35.820 150.350 ;
        RECT 35.620 148.990 35.760 150.030 ;
        RECT 35.560 148.670 35.820 148.990 ;
        RECT 35.100 147.990 35.360 148.310 ;
        RECT 37.000 146.610 37.140 151.050 ;
        RECT 38.840 151.030 38.980 156.070 ;
        RECT 39.760 154.430 39.900 159.210 ;
        RECT 40.680 156.810 40.820 160.910 ;
        RECT 42.060 159.870 42.200 161.250 ;
        RECT 42.520 159.870 42.660 161.590 ;
        RECT 42.980 160.210 43.120 161.930 ;
        RECT 50.280 161.590 50.540 161.910 ;
        RECT 47.520 160.910 47.780 161.230 ;
        RECT 48.440 160.910 48.700 161.230 ;
        RECT 42.920 159.890 43.180 160.210 ;
        RECT 42.000 159.550 42.260 159.870 ;
        RECT 42.460 159.550 42.720 159.870 ;
        RECT 41.540 159.210 41.800 159.530 ;
        RECT 41.600 157.490 41.740 159.210 ;
        RECT 41.540 157.170 41.800 157.490 ;
        RECT 40.620 156.490 40.880 156.810 ;
        RECT 39.700 154.110 39.960 154.430 ;
        RECT 39.240 153.090 39.500 153.410 ;
        RECT 39.300 151.030 39.440 153.090 ;
        RECT 39.760 151.030 39.900 154.110 ;
        RECT 42.060 151.030 42.200 159.550 ;
        RECT 47.580 155.790 47.720 160.910 ;
        RECT 47.980 156.380 48.240 156.470 ;
        RECT 48.500 156.380 48.640 160.910 ;
        RECT 50.340 160.210 50.480 161.590 ;
        RECT 53.560 161.570 53.700 166.350 ;
        RECT 54.420 161.590 54.680 161.910 ;
        RECT 53.560 161.430 54.160 161.570 ;
        RECT 53.500 160.910 53.760 161.230 ;
        RECT 50.280 159.890 50.540 160.210 ;
        RECT 48.900 159.210 49.160 159.530 ;
        RECT 48.960 157.490 49.100 159.210 ;
        RECT 48.900 157.170 49.160 157.490 ;
        RECT 47.980 156.240 48.640 156.380 ;
        RECT 47.980 156.150 48.240 156.240 ;
        RECT 49.820 155.810 50.080 156.130 ;
        RECT 42.920 155.470 43.180 155.790 ;
        RECT 47.520 155.470 47.780 155.790 ;
        RECT 42.980 152.130 43.120 155.470 ;
        RECT 49.360 153.770 49.620 154.090 ;
        RECT 42.520 151.990 43.120 152.130 ;
        RECT 38.780 150.710 39.040 151.030 ;
        RECT 39.240 150.710 39.500 151.030 ;
        RECT 39.700 150.710 39.960 151.030 ;
        RECT 42.000 150.710 42.260 151.030 ;
        RECT 39.760 149.330 39.900 150.710 ;
        RECT 39.700 149.010 39.960 149.330 ;
        RECT 41.540 147.650 41.800 147.970 ;
        RECT 36.940 146.290 37.200 146.610 ;
        RECT 34.640 145.950 34.900 146.270 ;
        RECT 39.240 144.590 39.500 144.910 ;
        RECT 39.300 143.550 39.440 144.590 ;
        RECT 34.180 143.290 34.440 143.550 ;
        RECT 34.180 143.230 35.760 143.290 ;
        RECT 39.240 143.230 39.500 143.550 ;
        RECT 34.240 143.150 35.760 143.230 ;
        RECT 41.600 143.210 41.740 147.650 ;
        RECT 42.520 145.930 42.660 151.990 ;
        RECT 42.920 151.050 43.180 151.370 ;
        RECT 42.980 145.930 43.120 151.050 ;
        RECT 44.760 150.710 45.020 151.030 ;
        RECT 43.840 148.330 44.100 148.650 ;
        RECT 43.900 146.610 44.040 148.330 ;
        RECT 43.840 146.290 44.100 146.610 ;
        RECT 42.460 145.610 42.720 145.930 ;
        RECT 42.920 145.610 43.180 145.930 ;
        RECT 44.820 143.210 44.960 150.710 ;
        RECT 49.420 148.650 49.560 153.770 ;
        RECT 49.360 148.330 49.620 148.650 ;
        RECT 46.600 147.990 46.860 148.310 ;
        RECT 46.660 143.550 46.800 147.990 ;
        RECT 47.060 145.950 47.320 146.270 ;
        RECT 46.600 143.230 46.860 143.550 ;
        RECT 31.880 139.150 32.140 139.470 ;
        RECT 32.230 138.615 33.770 138.985 ;
        RECT 35.620 138.110 35.760 143.150 ;
        RECT 39.700 142.890 39.960 143.210 ;
        RECT 41.540 142.890 41.800 143.210 ;
        RECT 44.760 142.890 45.020 143.210 ;
        RECT 36.480 142.550 36.740 142.870 ;
        RECT 36.540 141.170 36.680 142.550 ;
        RECT 39.240 141.870 39.500 142.190 ;
        RECT 36.480 140.850 36.740 141.170 ;
        RECT 39.300 140.150 39.440 141.870 ;
        RECT 39.760 140.490 39.900 142.890 ;
        RECT 42.460 141.870 42.720 142.190 ;
        RECT 45.680 141.870 45.940 142.190 ;
        RECT 39.700 140.170 39.960 140.490 ;
        RECT 36.940 139.830 37.200 140.150 ;
        RECT 39.240 139.830 39.500 140.150 ;
        RECT 35.560 137.790 35.820 138.110 ;
        RECT 37.000 137.430 37.140 139.830 ;
        RECT 36.940 137.110 37.200 137.430 ;
        RECT 34.180 135.070 34.440 135.390 ;
        RECT 31.880 134.450 32.140 134.710 ;
        RECT 31.480 134.390 32.140 134.450 ;
        RECT 31.480 134.310 32.080 134.390 ;
        RECT 29.120 133.710 29.380 134.030 ;
        RECT 28.260 131.590 28.860 131.730 ;
        RECT 28.260 129.860 28.400 131.590 ;
        RECT 29.180 131.310 29.320 133.710 ;
        RECT 31.480 133.010 31.620 134.310 ;
        RECT 32.230 133.175 33.770 133.545 ;
        RECT 31.420 132.690 31.680 133.010 ;
        RECT 30.960 131.670 31.220 131.990 ;
        RECT 29.120 130.990 29.380 131.310 ;
        RECT 28.930 130.455 30.470 130.825 ;
        RECT 28.260 129.720 28.860 129.860 ;
        RECT 28.720 128.930 28.860 129.720 ;
        RECT 28.660 128.610 28.920 128.930 ;
        RECT 26.820 128.270 27.080 128.590 ;
        RECT 26.880 124.170 27.020 128.270 ;
        RECT 28.720 127.570 28.860 128.610 ;
        RECT 28.660 127.250 28.920 127.570 ;
        RECT 28.930 125.015 30.470 125.385 ;
        RECT 26.820 123.850 27.080 124.170 ;
        RECT 31.020 122.130 31.160 131.670 ;
        RECT 31.420 130.990 31.680 131.310 ;
        RECT 30.960 121.810 31.220 122.130 ;
        RECT 23.140 121.130 23.400 121.450 ;
        RECT 23.600 121.130 23.860 121.450 ;
        RECT 23.200 118.730 23.340 121.130 ;
        RECT 23.660 119.410 23.800 121.130 ;
        RECT 28.930 119.575 30.470 119.945 ;
        RECT 31.480 119.410 31.620 130.990 ;
        RECT 34.240 129.610 34.380 135.070 ;
        RECT 37.000 134.710 37.140 137.110 ;
        RECT 42.520 134.710 42.660 141.870 ;
        RECT 45.220 139.490 45.480 139.810 ;
        RECT 45.280 138.450 45.420 139.490 ;
        RECT 45.220 138.130 45.480 138.450 ;
        RECT 45.740 137.770 45.880 141.870 ;
        RECT 47.120 138.450 47.260 145.950 ;
        RECT 48.900 145.270 49.160 145.590 ;
        RECT 47.520 144.930 47.780 145.250 ;
        RECT 47.580 142.190 47.720 144.930 ;
        RECT 47.520 141.870 47.780 142.190 ;
        RECT 47.580 138.450 47.720 141.870 ;
        RECT 48.960 139.470 49.100 145.270 ;
        RECT 49.880 145.250 50.020 155.810 ;
        RECT 50.340 154.770 50.480 159.890 ;
        RECT 53.560 159.530 53.700 160.910 ;
        RECT 53.500 159.210 53.760 159.530 ;
        RECT 52.580 158.530 52.840 158.850 ;
        RECT 52.640 157.150 52.780 158.530 ;
        RECT 52.580 156.830 52.840 157.150 ;
        RECT 50.280 154.680 50.540 154.770 ;
        RECT 50.280 154.540 50.940 154.680 ;
        RECT 50.280 154.450 50.540 154.540 ;
        RECT 50.280 152.750 50.540 153.070 ;
        RECT 50.340 152.050 50.480 152.750 ;
        RECT 50.280 151.730 50.540 152.050 ;
        RECT 50.800 151.030 50.940 154.540 ;
        RECT 53.560 154.090 53.700 159.210 ;
        RECT 53.500 153.770 53.760 154.090 ;
        RECT 51.660 152.750 51.920 153.070 ;
        RECT 51.720 151.370 51.860 152.750 ;
        RECT 51.660 151.050 51.920 151.370 ;
        RECT 50.740 150.710 51.000 151.030 ;
        RECT 51.200 150.370 51.460 150.690 ;
        RECT 50.280 148.330 50.540 148.650 ;
        RECT 49.820 144.930 50.080 145.250 ;
        RECT 50.340 143.550 50.480 148.330 ;
        RECT 51.260 143.890 51.400 150.370 ;
        RECT 51.200 143.570 51.460 143.890 ;
        RECT 50.280 143.230 50.540 143.550 ;
        RECT 49.360 142.890 49.620 143.210 ;
        RECT 49.420 140.830 49.560 142.890 ;
        RECT 49.820 142.210 50.080 142.530 ;
        RECT 49.360 140.510 49.620 140.830 ;
        RECT 48.900 139.150 49.160 139.470 ;
        RECT 47.060 138.130 47.320 138.450 ;
        RECT 47.520 138.130 47.780 138.450 ;
        RECT 45.680 137.450 45.940 137.770 ;
        RECT 47.120 135.730 47.260 138.130 ;
        RECT 48.960 137.430 49.100 139.150 ;
        RECT 49.880 138.450 50.020 142.210 ;
        RECT 50.340 141.170 50.480 143.230 ;
        RECT 50.280 140.850 50.540 141.170 ;
        RECT 50.340 138.450 50.480 140.850 ;
        RECT 51.260 140.490 51.400 143.570 ;
        RECT 53.500 141.870 53.760 142.190 ;
        RECT 52.580 140.510 52.840 140.830 ;
        RECT 51.200 140.170 51.460 140.490 ;
        RECT 50.740 139.490 51.000 139.810 ;
        RECT 49.820 138.130 50.080 138.450 ;
        RECT 50.280 138.130 50.540 138.450 ;
        RECT 50.800 137.850 50.940 139.490 ;
        RECT 50.340 137.770 50.940 137.850 ;
        RECT 51.260 137.770 51.400 140.170 ;
        RECT 52.640 137.770 52.780 140.510 ;
        RECT 53.560 140.150 53.700 141.870 ;
        RECT 53.500 139.830 53.760 140.150 ;
        RECT 53.040 139.490 53.300 139.810 ;
        RECT 53.100 138.450 53.240 139.490 ;
        RECT 53.040 138.130 53.300 138.450 ;
        RECT 53.560 137.850 53.700 139.830 ;
        RECT 50.280 137.710 50.940 137.770 ;
        RECT 50.280 137.450 50.540 137.710 ;
        RECT 51.200 137.450 51.460 137.770 ;
        RECT 52.580 137.450 52.840 137.770 ;
        RECT 53.100 137.710 53.700 137.850 ;
        RECT 48.900 137.110 49.160 137.430 ;
        RECT 42.920 135.410 43.180 135.730 ;
        RECT 47.060 135.410 47.320 135.730 ;
        RECT 36.940 134.390 37.200 134.710 ;
        RECT 42.460 134.390 42.720 134.710 ;
        RECT 34.640 134.050 34.900 134.370 ;
        RECT 34.700 131.310 34.840 134.050 ;
        RECT 36.020 131.670 36.280 131.990 ;
        RECT 34.640 130.990 34.900 131.310 ;
        RECT 34.180 129.290 34.440 129.610 ;
        RECT 32.230 127.735 33.770 128.105 ;
        RECT 36.080 127.570 36.220 131.670 ;
        RECT 37.000 129.270 37.140 134.390 ;
        RECT 39.700 134.050 39.960 134.370 ;
        RECT 39.760 131.650 39.900 134.050 ;
        RECT 42.980 132.330 43.120 135.410 ;
        RECT 48.960 135.050 49.100 137.110 ;
        RECT 49.820 136.430 50.080 136.750 ;
        RECT 48.900 134.730 49.160 135.050 ;
        RECT 47.520 133.710 47.780 134.030 ;
        RECT 47.580 132.330 47.720 133.710 ;
        RECT 48.960 132.670 49.100 134.730 ;
        RECT 48.900 132.350 49.160 132.670 ;
        RECT 42.920 132.010 43.180 132.330 ;
        RECT 47.060 132.010 47.320 132.330 ;
        RECT 47.520 132.010 47.780 132.330 ;
        RECT 39.700 131.330 39.960 131.650 ;
        RECT 37.860 130.990 38.120 131.310 ;
        RECT 42.920 130.990 43.180 131.310 ;
        RECT 45.680 130.990 45.940 131.310 ;
        RECT 37.920 129.270 38.060 130.990 ;
        RECT 42.460 129.630 42.720 129.950 ;
        RECT 36.940 128.950 37.200 129.270 ;
        RECT 37.860 128.950 38.120 129.270 ;
        RECT 40.620 129.010 40.880 129.270 ;
        RECT 40.620 128.950 41.280 129.010 ;
        RECT 36.020 127.250 36.280 127.570 ;
        RECT 35.100 126.570 35.360 126.890 ;
        RECT 35.160 124.850 35.300 126.570 ;
        RECT 37.000 126.210 37.140 128.950 ;
        RECT 40.680 128.870 41.280 128.950 ;
        RECT 40.620 128.270 40.880 128.590 ;
        RECT 37.400 126.230 37.660 126.550 ;
        RECT 40.160 126.230 40.420 126.550 ;
        RECT 36.940 125.890 37.200 126.210 ;
        RECT 37.460 124.930 37.600 126.230 ;
        RECT 39.700 125.550 39.960 125.870 ;
        RECT 35.100 124.530 35.360 124.850 ;
        RECT 37.000 124.790 37.600 124.930 ;
        RECT 37.000 124.170 37.140 124.790 ;
        RECT 37.400 124.190 37.660 124.510 ;
        RECT 39.760 124.250 39.900 125.550 ;
        RECT 40.220 124.850 40.360 126.230 ;
        RECT 40.160 124.530 40.420 124.850 ;
        RECT 36.940 123.850 37.200 124.170 ;
        RECT 31.880 122.830 32.140 123.150 ;
        RECT 23.600 119.090 23.860 119.410 ;
        RECT 24.520 119.090 24.780 119.410 ;
        RECT 31.420 119.090 31.680 119.410 ;
        RECT 23.140 118.410 23.400 118.730 ;
        RECT 18.080 117.390 18.340 117.710 ;
        RECT 12.090 115.835 12.370 116.205 ;
        RECT 12.100 115.690 12.360 115.835 ;
        RECT 16.700 115.010 16.960 115.330 ;
        RECT 12.100 112.805 12.360 112.950 ;
        RECT 8.420 112.290 8.680 112.610 ;
        RECT 12.090 112.435 12.370 112.805 ;
        RECT 16.760 110.570 16.900 115.010 ;
        RECT 17.160 112.630 17.420 112.950 ;
        RECT 16.700 110.250 16.960 110.570 ;
        RECT 14.390 108.355 14.670 108.725 ;
        RECT 14.460 104.450 14.600 108.355 ;
        RECT 16.760 107.170 16.900 110.250 ;
        RECT 15.320 106.850 15.580 107.170 ;
        RECT 16.700 106.850 16.960 107.170 ;
        RECT 15.380 105.810 15.520 106.850 ;
        RECT 15.320 105.490 15.580 105.810 ;
        RECT 16.760 105.470 16.900 106.850 ;
        RECT 17.220 105.470 17.360 112.630 ;
        RECT 18.140 110.570 18.280 117.390 ;
        RECT 23.200 112.950 23.340 118.410 ;
        RECT 24.580 118.390 24.720 119.090 ;
        RECT 24.520 118.070 24.780 118.390 ;
        RECT 24.980 118.070 25.240 118.390 ;
        RECT 24.060 117.730 24.320 118.050 ;
        RECT 24.120 116.350 24.260 117.730 ;
        RECT 24.520 117.390 24.780 117.710 ;
        RECT 24.060 116.030 24.320 116.350 ;
        RECT 21.760 112.630 22.020 112.950 ;
        RECT 23.140 112.630 23.400 112.950 ;
        RECT 19.460 111.950 19.720 112.270 ;
        RECT 18.080 110.250 18.340 110.570 ;
        RECT 17.620 109.910 17.880 110.230 ;
        RECT 16.700 105.150 16.960 105.470 ;
        RECT 17.160 105.150 17.420 105.470 ;
        RECT 17.680 104.790 17.820 109.910 ;
        RECT 17.620 104.470 17.880 104.790 ;
        RECT 14.400 104.130 14.660 104.450 ;
        RECT 12.090 102.235 12.370 102.605 ;
        RECT 12.160 102.070 12.300 102.235 ;
        RECT 18.140 102.070 18.280 110.250 ;
        RECT 18.540 109.230 18.800 109.550 ;
        RECT 18.600 105.130 18.740 109.230 ;
        RECT 19.520 105.470 19.660 111.950 ;
        RECT 21.820 111.160 21.960 112.630 ;
        RECT 23.200 111.250 23.340 112.630 ;
        RECT 21.360 111.020 21.960 111.160 ;
        RECT 21.360 108.530 21.500 111.020 ;
        RECT 22.220 110.930 22.480 111.250 ;
        RECT 23.140 110.930 23.400 111.250 ;
        RECT 21.760 110.250 22.020 110.570 ;
        RECT 21.300 108.210 21.560 108.530 ;
        RECT 19.460 105.150 19.720 105.470 ;
        RECT 21.360 105.130 21.500 108.210 ;
        RECT 21.820 107.510 21.960 110.250 ;
        RECT 21.760 107.190 22.020 107.510 ;
        RECT 22.280 105.470 22.420 110.930 ;
        RECT 23.140 110.250 23.400 110.570 ;
        RECT 23.200 108.530 23.340 110.250 ;
        RECT 23.140 108.210 23.400 108.530 ;
        RECT 23.600 107.530 23.860 107.850 ;
        RECT 22.680 107.190 22.940 107.510 ;
        RECT 22.220 105.150 22.480 105.470 ;
        RECT 18.540 104.810 18.800 105.130 ;
        RECT 21.300 104.810 21.560 105.130 ;
        RECT 22.740 103.090 22.880 107.190 ;
        RECT 23.660 105.810 23.800 107.530 ;
        RECT 24.580 107.510 24.720 117.390 ;
        RECT 25.040 116.010 25.180 118.070 ;
        RECT 26.360 117.730 26.620 118.050 ;
        RECT 24.980 115.690 25.240 116.010 ;
        RECT 26.420 115.330 26.560 117.730 ;
        RECT 30.960 117.390 31.220 117.710 ;
        RECT 27.280 116.030 27.540 116.350 ;
        RECT 27.340 115.670 27.480 116.030 ;
        RECT 27.280 115.350 27.540 115.670 ;
        RECT 26.360 115.010 26.620 115.330 ;
        RECT 26.820 112.290 27.080 112.610 ;
        RECT 26.360 107.870 26.620 108.190 ;
        RECT 24.520 107.190 24.780 107.510 ;
        RECT 25.900 107.190 26.160 107.510 ;
        RECT 25.960 105.890 26.100 107.190 ;
        RECT 23.600 105.490 23.860 105.810 ;
        RECT 24.120 105.750 26.100 105.890 ;
        RECT 23.130 104.955 23.410 105.325 ;
        RECT 23.140 104.810 23.400 104.955 ;
        RECT 23.600 104.470 23.860 104.790 ;
        RECT 21.760 102.770 22.020 103.090 ;
        RECT 22.680 102.770 22.940 103.090 ;
        RECT 12.100 101.750 12.360 102.070 ;
        RECT 18.080 101.750 18.340 102.070 ;
        RECT 19.460 101.750 19.720 102.070 ;
        RECT 18.540 101.070 18.800 101.390 ;
        RECT 14.860 99.370 15.120 99.690 ;
        RECT 14.920 91.530 15.060 99.370 ;
        RECT 18.600 97.650 18.740 101.070 ;
        RECT 19.520 97.650 19.660 101.750 ;
        RECT 21.820 99.090 21.960 102.770 ;
        RECT 23.660 102.410 23.800 104.470 ;
        RECT 24.120 102.750 24.260 105.750 ;
        RECT 25.440 105.150 25.700 105.470 ;
        RECT 24.520 104.130 24.780 104.450 ;
        RECT 24.060 102.430 24.320 102.750 ;
        RECT 23.600 102.090 23.860 102.410 ;
        RECT 23.600 101.410 23.860 101.730 ;
        RECT 22.220 101.070 22.480 101.390 ;
        RECT 22.280 99.690 22.420 101.070 ;
        RECT 23.660 100.370 23.800 101.410 ;
        RECT 24.120 100.370 24.260 102.430 ;
        RECT 23.600 100.050 23.860 100.370 ;
        RECT 24.060 100.050 24.320 100.370 ;
        RECT 22.220 99.370 22.480 99.690 ;
        RECT 24.580 99.470 24.720 104.130 ;
        RECT 21.360 98.950 21.960 99.090 ;
        RECT 24.120 99.330 24.720 99.470 ;
        RECT 25.500 99.350 25.640 105.150 ;
        RECT 25.960 104.790 26.100 105.750 ;
        RECT 26.420 105.130 26.560 107.870 ;
        RECT 26.880 107.170 27.020 112.290 ;
        RECT 27.340 110.570 27.480 115.350 ;
        RECT 31.020 115.330 31.160 117.390 ;
        RECT 31.940 116.010 32.080 122.830 ;
        RECT 32.230 122.295 33.770 122.665 ;
        RECT 34.180 117.390 34.440 117.710 ;
        RECT 32.230 116.855 33.770 117.225 ;
        RECT 34.240 116.350 34.380 117.390 ;
        RECT 34.180 116.030 34.440 116.350 ;
        RECT 31.880 115.690 32.140 116.010 ;
        RECT 30.960 115.010 31.220 115.330 ;
        RECT 28.930 114.135 30.470 114.505 ;
        RECT 31.020 110.570 31.160 115.010 ;
        RECT 31.940 114.990 32.080 115.690 ;
        RECT 36.940 115.350 37.200 115.670 ;
        RECT 37.460 115.410 37.600 124.190 ;
        RECT 38.380 124.110 39.900 124.250 ;
        RECT 37.860 123.740 38.120 123.830 ;
        RECT 38.380 123.740 38.520 124.110 ;
        RECT 39.760 123.830 39.900 124.110 ;
        RECT 37.860 123.600 38.520 123.740 ;
        RECT 37.860 123.510 38.120 123.600 ;
        RECT 37.860 117.390 38.120 117.710 ;
        RECT 37.920 116.010 38.060 117.390 ;
        RECT 37.860 115.690 38.120 116.010 ;
        RECT 31.880 114.670 32.140 114.990 ;
        RECT 36.020 114.670 36.280 114.990 ;
        RECT 31.420 112.630 31.680 112.950 ;
        RECT 31.480 110.570 31.620 112.630 ;
        RECT 32.230 111.415 33.770 111.785 ;
        RECT 36.080 110.910 36.220 114.670 ;
        RECT 37.000 112.690 37.140 115.350 ;
        RECT 37.460 115.270 38.060 115.410 ;
        RECT 37.400 114.670 37.660 114.990 ;
        RECT 36.540 112.550 37.140 112.690 ;
        RECT 36.020 110.590 36.280 110.910 ;
        RECT 36.540 110.570 36.680 112.550 ;
        RECT 36.940 111.950 37.200 112.270 ;
        RECT 27.280 110.250 27.540 110.570 ;
        RECT 30.960 110.250 31.220 110.570 ;
        RECT 31.420 110.250 31.680 110.570 ;
        RECT 36.480 110.250 36.740 110.570 ;
        RECT 27.340 108.530 27.480 110.250 ;
        RECT 27.740 109.230 28.000 109.550 ;
        RECT 28.200 109.230 28.460 109.550 ;
        RECT 27.800 108.530 27.940 109.230 ;
        RECT 27.280 108.210 27.540 108.530 ;
        RECT 27.740 108.210 28.000 108.530 ;
        RECT 28.260 108.190 28.400 109.230 ;
        RECT 28.930 108.695 30.470 109.065 ;
        RECT 28.200 107.870 28.460 108.190 ;
        RECT 31.020 107.510 31.160 110.250 ;
        RECT 36.540 108.530 36.680 110.250 ;
        RECT 36.480 108.210 36.740 108.530 ;
        RECT 37.000 107.850 37.140 111.950 ;
        RECT 36.940 107.530 37.200 107.850 ;
        RECT 37.460 107.510 37.600 114.670 ;
        RECT 30.960 107.190 31.220 107.510 ;
        RECT 37.400 107.190 37.660 107.510 ;
        RECT 26.820 106.850 27.080 107.170 ;
        RECT 31.420 106.850 31.680 107.170 ;
        RECT 26.360 104.810 26.620 105.130 ;
        RECT 26.820 104.810 27.080 105.130 ;
        RECT 25.900 104.470 26.160 104.790 ;
        RECT 25.900 103.790 26.160 104.110 ;
        RECT 26.360 103.790 26.620 104.110 ;
        RECT 18.540 97.330 18.800 97.650 ;
        RECT 19.460 97.330 19.720 97.650 ;
        RECT 18.600 94.590 18.740 97.330 ;
        RECT 18.540 94.270 18.800 94.590 ;
        RECT 21.360 93.910 21.500 98.950 ;
        RECT 21.760 98.350 22.020 98.670 ;
        RECT 22.220 98.350 22.480 98.670 ;
        RECT 21.820 96.630 21.960 98.350 ;
        RECT 21.760 96.310 22.020 96.630 ;
        RECT 19.000 93.590 19.260 93.910 ;
        RECT 21.300 93.590 21.560 93.910 ;
        RECT 16.240 92.910 16.500 93.230 ;
        RECT 14.860 91.210 15.120 91.530 ;
        RECT 16.300 90.850 16.440 92.910 ;
        RECT 19.060 91.610 19.200 93.590 ;
        RECT 21.820 93.230 21.960 96.310 ;
        RECT 21.760 92.910 22.020 93.230 ;
        RECT 18.600 91.470 19.200 91.610 ;
        RECT 16.240 90.530 16.500 90.850 ;
        RECT 18.600 89.490 18.740 91.470 ;
        RECT 21.760 90.870 22.020 91.190 ;
        RECT 19.000 90.530 19.260 90.850 ;
        RECT 18.540 89.170 18.800 89.490 ;
        RECT 19.060 88.810 19.200 90.530 ;
        RECT 21.820 89.150 21.960 90.870 ;
        RECT 22.280 90.510 22.420 98.350 ;
        RECT 22.680 95.970 22.940 96.290 ;
        RECT 22.740 94.250 22.880 95.970 ;
        RECT 23.140 94.610 23.400 94.930 ;
        RECT 22.680 93.930 22.940 94.250 ;
        RECT 22.680 93.250 22.940 93.570 ;
        RECT 22.740 92.210 22.880 93.250 ;
        RECT 22.680 91.890 22.940 92.210 ;
        RECT 23.200 91.610 23.340 94.610 ;
        RECT 23.200 91.530 23.800 91.610 ;
        RECT 23.140 91.470 23.800 91.530 ;
        RECT 23.140 91.210 23.400 91.470 ;
        RECT 23.140 90.530 23.400 90.850 ;
        RECT 22.220 90.420 22.480 90.510 ;
        RECT 22.220 90.280 22.880 90.420 ;
        RECT 22.220 90.190 22.480 90.280 ;
        RECT 21.760 88.830 22.020 89.150 ;
        RECT 19.000 88.490 19.260 88.810 ;
        RECT 20.380 84.750 20.640 85.070 ;
        RECT 20.440 80.310 20.580 84.750 ;
        RECT 20.380 80.220 20.640 80.310 ;
        RECT 20.380 80.080 21.040 80.220 ;
        RECT 20.380 79.990 20.640 80.080 ;
        RECT 20.900 79.630 21.040 80.080 ;
        RECT 21.300 79.650 21.560 79.970 ;
        RECT 18.540 79.310 18.800 79.630 ;
        RECT 20.840 79.310 21.100 79.630 ;
        RECT 17.160 77.610 17.420 77.930 ;
        RECT 17.220 75.890 17.360 77.610 ;
        RECT 17.160 75.570 17.420 75.890 ;
        RECT 18.080 74.890 18.340 75.210 ;
        RECT 18.140 72.150 18.280 74.890 ;
        RECT 18.600 74.870 18.740 79.310 ;
        RECT 18.540 74.550 18.800 74.870 ;
        RECT 20.900 74.530 21.040 79.310 ;
        RECT 21.360 75.210 21.500 79.650 ;
        RECT 21.820 78.270 21.960 88.830 ;
        RECT 22.220 88.490 22.480 88.810 ;
        RECT 22.280 86.770 22.420 88.490 ;
        RECT 22.220 86.450 22.480 86.770 ;
        RECT 22.220 85.090 22.480 85.410 ;
        RECT 22.280 84.130 22.420 85.090 ;
        RECT 22.740 85.070 22.880 90.280 ;
        RECT 23.200 87.790 23.340 90.530 ;
        RECT 23.140 87.470 23.400 87.790 ;
        RECT 22.680 84.750 22.940 85.070 ;
        RECT 23.200 84.130 23.340 87.470 ;
        RECT 23.660 86.430 23.800 91.470 ;
        RECT 23.600 86.110 23.860 86.430 ;
        RECT 23.600 85.430 23.860 85.750 ;
        RECT 22.280 83.990 23.340 84.130 ;
        RECT 22.280 80.990 22.420 83.990 ;
        RECT 22.680 81.010 22.940 81.330 ;
        RECT 22.220 80.670 22.480 80.990 ;
        RECT 22.740 80.310 22.880 81.010 ;
        RECT 23.660 80.650 23.800 85.430 ;
        RECT 23.600 80.330 23.860 80.650 ;
        RECT 22.680 79.990 22.940 80.310 ;
        RECT 22.740 78.610 22.880 79.990 ;
        RECT 23.600 79.650 23.860 79.970 ;
        RECT 22.680 78.290 22.940 78.610 ;
        RECT 21.760 77.950 22.020 78.270 ;
        RECT 21.300 74.890 21.560 75.210 ;
        RECT 20.840 74.210 21.100 74.530 ;
        RECT 21.820 72.830 21.960 77.950 ;
        RECT 22.740 75.890 22.880 78.290 ;
        RECT 23.660 77.930 23.800 79.650 ;
        RECT 23.600 77.610 23.860 77.930 ;
        RECT 23.660 75.890 23.800 77.610 ;
        RECT 22.680 75.570 22.940 75.890 ;
        RECT 23.600 75.570 23.860 75.890 ;
        RECT 22.740 74.870 22.880 75.570 ;
        RECT 22.680 74.550 22.940 74.870 ;
        RECT 22.220 73.870 22.480 74.190 ;
        RECT 21.760 72.510 22.020 72.830 ;
        RECT 21.300 72.170 21.560 72.490 ;
        RECT 18.080 71.830 18.340 72.150 ;
        RECT 20.840 71.490 21.100 71.810 ;
        RECT 15.320 71.150 15.580 71.470 ;
        RECT 19.000 71.150 19.260 71.470 ;
        RECT 15.380 69.090 15.520 71.150 ;
        RECT 15.320 68.770 15.580 69.090 ;
        RECT 14.390 67.555 14.670 67.925 ;
        RECT 14.400 67.410 14.660 67.555 ;
        RECT 19.060 67.050 19.200 71.150 ;
        RECT 20.900 70.450 21.040 71.490 ;
        RECT 19.460 70.130 19.720 70.450 ;
        RECT 20.840 70.130 21.100 70.450 ;
        RECT 19.000 66.730 19.260 67.050 ;
        RECT 19.520 66.030 19.660 70.130 ;
        RECT 21.360 70.110 21.500 72.170 ;
        RECT 21.300 69.790 21.560 70.110 ;
        RECT 21.360 66.450 21.500 69.790 ;
        RECT 21.820 69.430 21.960 72.510 ;
        RECT 22.280 72.150 22.420 73.870 ;
        RECT 22.680 72.850 22.940 73.170 ;
        RECT 22.740 72.490 22.880 72.850 ;
        RECT 22.680 72.170 22.940 72.490 ;
        RECT 22.220 71.830 22.480 72.150 ;
        RECT 21.760 69.110 22.020 69.430 ;
        RECT 21.820 67.390 21.960 69.110 ;
        RECT 21.760 67.070 22.020 67.390 ;
        RECT 20.900 66.310 21.500 66.450 ;
        RECT 19.460 65.710 19.720 66.030 ;
        RECT 12.090 63.475 12.370 63.845 ;
        RECT 16.240 63.670 16.500 63.990 ;
        RECT 12.160 63.310 12.300 63.475 ;
        RECT 12.100 62.990 12.360 63.310 ;
        RECT 13.470 60.755 13.750 61.125 ;
        RECT 16.300 60.930 16.440 63.670 ;
        RECT 17.160 62.990 17.420 63.310 ;
        RECT 13.540 59.570 13.680 60.755 ;
        RECT 16.240 60.610 16.500 60.930 ;
        RECT 13.480 59.250 13.740 59.570 ;
        RECT 16.700 58.230 16.960 58.550 ;
        RECT 14.390 53.955 14.670 54.325 ;
        RECT 13.010 50.555 13.290 50.925 ;
        RECT 13.080 50.050 13.220 50.555 ;
        RECT 13.020 49.730 13.280 50.050 ;
        RECT 14.460 49.710 14.600 53.955 ;
        RECT 16.760 53.450 16.900 58.230 ;
        RECT 17.220 57.725 17.360 62.990 ;
        RECT 18.540 60.270 18.800 60.590 ;
        RECT 18.080 57.890 18.340 58.210 ;
        RECT 17.150 57.355 17.430 57.725 ;
        RECT 18.140 56.850 18.280 57.890 ;
        RECT 18.080 56.530 18.340 56.850 ;
        RECT 18.600 56.170 18.740 60.270 ;
        RECT 19.000 57.890 19.260 58.210 ;
        RECT 19.060 56.170 19.200 57.890 ;
        RECT 19.460 57.550 19.720 57.870 ;
        RECT 18.540 55.850 18.800 56.170 ;
        RECT 19.000 55.850 19.260 56.170 ;
        RECT 16.700 53.130 16.960 53.450 ;
        RECT 14.860 52.450 15.120 52.770 ;
        RECT 14.400 49.390 14.660 49.710 ;
        RECT 12.100 48.205 12.360 48.350 ;
        RECT 12.090 47.835 12.370 48.205 ;
        RECT 14.920 45.630 15.060 52.450 ;
        RECT 16.240 52.110 16.500 52.430 ;
        RECT 16.300 50.730 16.440 52.110 ;
        RECT 16.240 50.410 16.500 50.730 ;
        RECT 16.240 49.390 16.500 49.710 ;
        RECT 16.300 47.670 16.440 49.390 ;
        RECT 16.240 47.350 16.500 47.670 ;
        RECT 14.860 45.310 15.120 45.630 ;
        RECT 16.760 44.950 16.900 53.130 ;
        RECT 19.520 47.670 19.660 57.550 ;
        RECT 20.900 56.930 21.040 66.310 ;
        RECT 21.300 65.710 21.560 66.030 ;
        RECT 21.360 57.870 21.500 65.710 ;
        RECT 21.820 61.610 21.960 67.070 ;
        RECT 22.680 63.670 22.940 63.990 ;
        RECT 22.220 61.630 22.480 61.950 ;
        RECT 21.760 61.290 22.020 61.610 ;
        RECT 22.280 59.230 22.420 61.630 ;
        RECT 22.740 61.270 22.880 63.670 ;
        RECT 23.140 62.990 23.400 63.310 ;
        RECT 22.680 60.950 22.940 61.270 ;
        RECT 22.740 59.570 22.880 60.950 ;
        RECT 22.680 59.250 22.940 59.570 ;
        RECT 22.220 58.910 22.480 59.230 ;
        RECT 22.280 58.550 22.420 58.910 ;
        RECT 22.220 58.230 22.480 58.550 ;
        RECT 23.200 58.210 23.340 62.990 ;
        RECT 24.120 61.270 24.260 99.330 ;
        RECT 25.440 99.030 25.700 99.350 ;
        RECT 25.500 96.290 25.640 99.030 ;
        RECT 25.440 95.970 25.700 96.290 ;
        RECT 25.440 93.590 25.700 93.910 ;
        RECT 24.980 93.250 25.240 93.570 ;
        RECT 24.520 91.890 24.780 92.210 ;
        RECT 24.580 89.490 24.720 91.890 ;
        RECT 24.520 89.170 24.780 89.490 ;
        RECT 24.580 88.130 24.720 89.170 ;
        RECT 24.520 87.810 24.780 88.130 ;
        RECT 24.580 81.330 24.720 87.810 ;
        RECT 24.520 81.010 24.780 81.330 ;
        RECT 25.040 77.840 25.180 93.250 ;
        RECT 25.500 91.190 25.640 93.590 ;
        RECT 25.960 92.210 26.100 103.790 ;
        RECT 26.420 102.070 26.560 103.790 ;
        RECT 26.880 102.410 27.020 104.810 ;
        RECT 28.930 103.255 30.470 103.625 ;
        RECT 26.820 102.090 27.080 102.410 ;
        RECT 26.360 101.750 26.620 102.070 ;
        RECT 26.360 99.030 26.620 99.350 ;
        RECT 26.420 94.930 26.560 99.030 ;
        RECT 26.880 96.970 27.020 102.090 ;
        RECT 28.930 97.815 30.470 98.185 ;
        RECT 26.820 96.650 27.080 96.970 ;
        RECT 26.360 94.610 26.620 94.930 ;
        RECT 26.880 94.250 27.020 96.650 ;
        RECT 26.820 93.930 27.080 94.250 ;
        RECT 27.740 93.930 28.000 94.250 ;
        RECT 25.900 91.890 26.160 92.210 ;
        RECT 25.440 90.870 25.700 91.190 ;
        RECT 26.360 89.170 26.620 89.490 ;
        RECT 26.420 87.790 26.560 89.170 ;
        RECT 26.880 88.470 27.020 93.930 ;
        RECT 27.800 92.210 27.940 93.930 ;
        RECT 28.930 92.375 30.470 92.745 ;
        RECT 27.740 91.890 28.000 92.210 ;
        RECT 27.740 90.870 28.000 91.190 ;
        RECT 27.280 88.830 27.540 89.150 ;
        RECT 26.820 88.150 27.080 88.470 ;
        RECT 26.360 87.470 26.620 87.790 ;
        RECT 26.880 86.090 27.020 88.150 ;
        RECT 27.340 86.770 27.480 88.830 ;
        RECT 27.280 86.450 27.540 86.770 ;
        RECT 25.440 85.770 25.700 86.090 ;
        RECT 26.820 85.770 27.080 86.090 ;
        RECT 24.580 77.700 25.180 77.840 ;
        RECT 24.060 60.950 24.320 61.270 ;
        RECT 23.140 57.890 23.400 58.210 ;
        RECT 21.300 57.550 21.560 57.870 ;
        RECT 19.980 56.790 21.500 56.930 ;
        RECT 19.980 56.170 20.120 56.790 ;
        RECT 20.840 56.365 21.100 56.510 ;
        RECT 19.920 55.850 20.180 56.170 ;
        RECT 20.830 55.995 21.110 56.365 ;
        RECT 19.920 54.830 20.180 55.150 ;
        RECT 20.380 54.830 20.640 55.150 ;
        RECT 19.980 52.770 20.120 54.830 ;
        RECT 19.920 52.450 20.180 52.770 ;
        RECT 20.440 52.170 20.580 54.830 ;
        RECT 19.980 52.030 20.580 52.170 ;
        RECT 18.080 47.350 18.340 47.670 ;
        RECT 19.460 47.350 19.720 47.670 ;
        RECT 18.140 45.970 18.280 47.350 ;
        RECT 18.080 45.650 18.340 45.970 ;
        RECT 16.700 44.630 16.960 44.950 ;
        RECT 16.760 43.250 16.900 44.630 ;
        RECT 16.700 42.930 16.960 43.250 ;
        RECT 16.240 41.570 16.500 41.890 ;
        RECT 16.300 40.530 16.440 41.570 ;
        RECT 16.240 40.210 16.500 40.530 ;
        RECT 16.760 37.130 16.900 42.930 ;
        RECT 17.620 39.760 17.880 39.850 ;
        RECT 17.220 39.620 17.880 39.760 ;
        RECT 16.700 36.810 16.960 37.130 ;
        RECT 16.700 31.090 16.960 31.350 ;
        RECT 16.300 31.030 16.960 31.090 ;
        RECT 16.300 30.950 16.900 31.030 ;
        RECT 15.780 30.350 16.040 30.670 ;
        RECT 15.320 27.630 15.580 27.950 ;
        RECT 15.380 25.570 15.520 27.630 ;
        RECT 15.320 25.250 15.580 25.570 ;
        RECT 14.860 22.190 15.120 22.510 ;
        RECT 7.960 9.270 8.220 9.590 ;
        RECT 14.920 9.330 15.060 22.190 ;
        RECT 15.320 19.470 15.580 19.790 ;
        RECT 15.380 14.690 15.520 19.470 ;
        RECT 15.320 14.370 15.580 14.690 ;
        RECT 15.840 9.590 15.980 30.350 ;
        RECT 16.300 18.430 16.440 30.950 ;
        RECT 17.220 28.970 17.360 39.620 ;
        RECT 17.620 39.530 17.880 39.620 ;
        RECT 18.080 36.810 18.340 37.130 ;
        RECT 17.620 30.350 17.880 30.670 ;
        RECT 17.680 28.970 17.820 30.350 ;
        RECT 17.160 28.650 17.420 28.970 ;
        RECT 17.620 28.650 17.880 28.970 ;
        RECT 17.220 20.470 17.360 28.650 ;
        RECT 18.140 28.630 18.280 36.810 ;
        RECT 19.000 31.710 19.260 32.030 ;
        RECT 19.060 31.350 19.200 31.710 ;
        RECT 19.520 31.350 19.660 47.350 ;
        RECT 19.980 39.365 20.120 52.030 ;
        RECT 20.380 50.410 20.640 50.730 ;
        RECT 20.440 43.250 20.580 50.410 ;
        RECT 20.900 48.010 21.040 55.995 ;
        RECT 20.840 47.690 21.100 48.010 ;
        RECT 20.840 46.670 21.100 46.990 ;
        RECT 20.900 45.630 21.040 46.670 ;
        RECT 20.840 45.310 21.100 45.630 ;
        RECT 20.380 42.930 20.640 43.250 ;
        RECT 20.440 40.190 20.580 42.930 ;
        RECT 20.380 39.870 20.640 40.190 ;
        RECT 20.840 39.530 21.100 39.850 ;
        RECT 19.910 38.995 20.190 39.365 ;
        RECT 19.000 31.030 19.260 31.350 ;
        RECT 19.460 31.030 19.720 31.350 ;
        RECT 18.540 30.690 18.800 31.010 ;
        RECT 18.080 28.310 18.340 28.630 ;
        RECT 18.140 25.910 18.280 28.310 ;
        RECT 18.600 26.930 18.740 30.690 ;
        RECT 19.520 29.650 19.660 31.030 ;
        RECT 19.460 29.330 19.720 29.650 ;
        RECT 18.540 26.610 18.800 26.930 ;
        RECT 18.080 25.590 18.340 25.910 ;
        RECT 17.160 20.150 17.420 20.470 ;
        RECT 17.620 20.150 17.880 20.470 ;
        RECT 17.680 18.770 17.820 20.150 ;
        RECT 17.620 18.450 17.880 18.770 ;
        RECT 16.240 18.110 16.500 18.430 ;
        RECT 18.140 18.090 18.280 25.590 ;
        RECT 18.600 23.530 18.740 26.610 ;
        RECT 18.540 23.210 18.800 23.530 ;
        RECT 18.540 22.190 18.800 22.510 ;
        RECT 19.460 22.190 19.720 22.510 ;
        RECT 18.080 17.770 18.340 18.090 ;
        RECT 18.600 16.670 18.740 22.190 ;
        RECT 19.000 17.770 19.260 18.090 ;
        RECT 18.140 16.530 18.740 16.670 ;
        RECT 18.140 12.730 18.280 16.530 ;
        RECT 19.060 15.030 19.200 17.770 ;
        RECT 19.000 14.710 19.260 15.030 ;
        RECT 17.680 12.590 18.280 12.730 ;
        RECT 8.020 6.800 8.160 9.270 ;
        RECT 11.180 8.930 11.440 9.250 ;
        RECT 14.460 9.190 15.060 9.330 ;
        RECT 15.780 9.270 16.040 9.590 ;
        RECT 11.240 6.800 11.380 8.930 ;
        RECT 14.460 6.800 14.600 9.190 ;
        RECT 17.680 6.800 17.820 12.590 ;
        RECT 19.520 9.250 19.660 22.190 ;
        RECT 19.980 20.810 20.120 38.995 ;
        RECT 20.900 32.030 21.040 39.530 ;
        RECT 21.360 38.830 21.500 56.790 ;
        RECT 21.760 56.530 22.020 56.850 ;
        RECT 21.820 56.365 21.960 56.530 ;
        RECT 21.750 56.170 22.030 56.365 ;
        RECT 23.200 56.170 23.340 57.890 ;
        RECT 24.580 56.930 24.720 77.700 ;
        RECT 24.980 76.930 25.240 77.250 ;
        RECT 25.040 72.150 25.180 76.930 ;
        RECT 25.500 76.910 25.640 85.770 ;
        RECT 27.800 83.710 27.940 90.870 ;
        RECT 30.960 87.470 31.220 87.790 ;
        RECT 28.930 86.935 30.470 87.305 ;
        RECT 28.200 85.090 28.460 85.410 ;
        RECT 28.260 84.050 28.400 85.090 ;
        RECT 28.200 83.730 28.460 84.050 ;
        RECT 27.740 83.390 28.000 83.710 ;
        RECT 27.800 80.310 27.940 83.390 ;
        RECT 31.020 83.030 31.160 87.470 ;
        RECT 31.480 86.170 31.620 106.850 ;
        RECT 36.480 106.510 36.740 106.830 ;
        RECT 32.230 105.975 33.770 106.345 ;
        RECT 36.540 105.470 36.680 106.510 ;
        RECT 36.480 105.150 36.740 105.470 ;
        RECT 32.230 100.535 33.770 100.905 ;
        RECT 34.180 98.350 34.440 98.670 ;
        RECT 32.230 95.095 33.770 95.465 ;
        RECT 34.240 94.930 34.380 98.350 ;
        RECT 37.920 97.650 38.060 115.270 ;
        RECT 37.860 97.330 38.120 97.650 ;
        RECT 35.560 95.970 35.820 96.290 ;
        RECT 35.620 94.930 35.760 95.970 ;
        RECT 34.180 94.610 34.440 94.930 ;
        RECT 35.560 94.610 35.820 94.930 ;
        RECT 34.240 90.850 34.380 94.610 ;
        RECT 37.920 94.590 38.060 97.330 ;
        RECT 37.860 94.270 38.120 94.590 ;
        RECT 38.380 93.910 38.520 123.600 ;
        RECT 39.240 123.510 39.500 123.830 ;
        RECT 39.700 123.510 39.960 123.830 ;
        RECT 39.300 116.690 39.440 123.510 ;
        RECT 40.680 123.490 40.820 128.270 ;
        RECT 40.620 123.170 40.880 123.490 ;
        RECT 41.140 120.770 41.280 128.870 ;
        RECT 42.000 126.230 42.260 126.550 ;
        RECT 42.060 125.870 42.200 126.230 ;
        RECT 42.000 125.550 42.260 125.870 ;
        RECT 41.540 124.250 41.800 124.510 ;
        RECT 42.520 124.250 42.660 129.630 ;
        RECT 42.980 124.850 43.120 130.990 ;
        RECT 45.740 129.270 45.880 130.990 ;
        RECT 43.380 128.950 43.640 129.270 ;
        RECT 45.680 128.950 45.940 129.270 ;
        RECT 42.920 124.530 43.180 124.850 ;
        RECT 41.540 124.190 42.660 124.250 ;
        RECT 41.600 124.110 42.660 124.190 ;
        RECT 41.080 120.450 41.340 120.770 ;
        RECT 41.140 118.810 41.280 120.450 ;
        RECT 40.680 118.670 41.280 118.810 ;
        RECT 39.240 116.370 39.500 116.690 ;
        RECT 40.680 116.010 40.820 118.670 ;
        RECT 41.080 118.070 41.340 118.390 ;
        RECT 40.620 115.690 40.880 116.010 ;
        RECT 40.620 111.950 40.880 112.270 ;
        RECT 40.680 109.550 40.820 111.950 ;
        RECT 41.140 110.570 41.280 118.070 ;
        RECT 42.000 115.690 42.260 116.010 ;
        RECT 41.540 115.350 41.800 115.670 ;
        RECT 41.600 112.270 41.740 115.350 ;
        RECT 41.540 111.950 41.800 112.270 ;
        RECT 41.600 110.910 41.740 111.950 ;
        RECT 41.540 110.590 41.800 110.910 ;
        RECT 41.080 110.250 41.340 110.570 ;
        RECT 40.160 109.230 40.420 109.550 ;
        RECT 40.620 109.230 40.880 109.550 ;
        RECT 39.700 107.870 39.960 108.190 ;
        RECT 40.220 108.100 40.360 109.230 ;
        RECT 40.620 108.100 40.880 108.190 ;
        RECT 40.220 107.960 40.880 108.100 ;
        RECT 40.620 107.870 40.880 107.960 ;
        RECT 42.060 107.930 42.200 115.690 ;
        RECT 42.920 115.010 43.180 115.330 ;
        RECT 42.980 112.950 43.120 115.010 ;
        RECT 42.920 112.630 43.180 112.950 ;
        RECT 42.980 111.250 43.120 112.630 ;
        RECT 42.920 110.930 43.180 111.250 ;
        RECT 42.460 110.250 42.720 110.570 ;
        RECT 42.520 108.530 42.660 110.250 ;
        RECT 42.460 108.210 42.720 108.530 ;
        RECT 38.780 106.850 39.040 107.170 ;
        RECT 38.840 105.810 38.980 106.850 ;
        RECT 39.760 105.810 39.900 107.870 ;
        RECT 41.600 107.790 42.200 107.930 ;
        RECT 38.780 105.490 39.040 105.810 ;
        RECT 39.700 105.490 39.960 105.810 ;
        RECT 39.700 104.810 39.960 105.130 ;
        RECT 39.760 103.090 39.900 104.810 ;
        RECT 39.700 102.770 39.960 103.090 ;
        RECT 41.080 101.750 41.340 102.070 ;
        RECT 41.140 100.370 41.280 101.750 ;
        RECT 41.600 101.390 41.740 107.790 ;
        RECT 42.000 107.190 42.260 107.510 ;
        RECT 42.060 105.810 42.200 107.190 ;
        RECT 42.000 105.490 42.260 105.810 ;
        RECT 42.060 102.070 42.200 105.490 ;
        RECT 42.920 104.810 43.180 105.130 ;
        RECT 42.980 102.490 43.120 104.810 ;
        RECT 43.440 103.090 43.580 128.950 ;
        RECT 45.220 128.610 45.480 128.930 ;
        RECT 45.280 126.890 45.420 128.610 ;
        RECT 45.740 127.230 45.880 128.950 ;
        RECT 46.140 128.270 46.400 128.590 ;
        RECT 45.680 126.910 45.940 127.230 ;
        RECT 46.200 126.890 46.340 128.270 ;
        RECT 45.220 126.570 45.480 126.890 ;
        RECT 46.140 126.570 46.400 126.890 ;
        RECT 44.300 126.290 44.560 126.550 ;
        RECT 44.300 126.230 45.420 126.290 ;
        RECT 45.680 126.230 45.940 126.550 ;
        RECT 46.600 126.230 46.860 126.550 ;
        RECT 44.360 126.150 45.420 126.230 ;
        RECT 43.840 125.550 44.100 125.870 ;
        RECT 44.760 125.550 45.020 125.870 ;
        RECT 43.900 123.490 44.040 125.550 ;
        RECT 44.820 123.830 44.960 125.550 ;
        RECT 45.280 124.850 45.420 126.150 ;
        RECT 45.740 125.870 45.880 126.230 ;
        RECT 45.680 125.550 45.940 125.870 ;
        RECT 45.220 124.530 45.480 124.850 ;
        RECT 44.760 123.510 45.020 123.830 ;
        RECT 43.840 123.170 44.100 123.490 ;
        RECT 44.300 115.690 44.560 116.010 ;
        RECT 43.840 114.670 44.100 114.990 ;
        RECT 43.900 112.950 44.040 114.670 ;
        RECT 44.360 112.950 44.500 115.690 ;
        RECT 44.820 113.290 44.960 123.510 ;
        RECT 46.660 123.150 46.800 126.230 ;
        RECT 47.120 124.850 47.260 132.010 ;
        RECT 47.580 129.610 47.720 132.010 ;
        RECT 48.960 131.650 49.100 132.350 ;
        RECT 49.880 132.330 50.020 136.430 ;
        RECT 49.820 132.010 50.080 132.330 ;
        RECT 50.340 131.990 50.480 137.450 ;
        RECT 53.100 132.670 53.240 137.710 ;
        RECT 53.500 136.770 53.760 137.090 ;
        RECT 53.560 134.710 53.700 136.770 ;
        RECT 53.500 134.390 53.760 134.710 ;
        RECT 53.040 132.350 53.300 132.670 ;
        RECT 50.280 131.670 50.540 131.990 ;
        RECT 48.900 131.330 49.160 131.650 ;
        RECT 47.520 129.290 47.780 129.610 ;
        RECT 48.960 125.870 49.100 131.330 ;
        RECT 49.360 128.950 49.620 129.270 ;
        RECT 48.900 125.550 49.160 125.870 ;
        RECT 47.060 124.530 47.320 124.850 ;
        RECT 48.440 124.530 48.700 124.850 ;
        RECT 46.600 122.830 46.860 123.150 ;
        RECT 46.660 122.130 46.800 122.830 ;
        RECT 46.600 121.810 46.860 122.130 ;
        RECT 48.500 121.450 48.640 124.530 ;
        RECT 49.420 124.170 49.560 128.950 ;
        RECT 49.820 128.270 50.080 128.590 ;
        RECT 49.360 123.850 49.620 124.170 ;
        RECT 48.900 123.510 49.160 123.830 ;
        RECT 48.960 122.130 49.100 123.510 ;
        RECT 48.900 121.810 49.160 122.130 ;
        RECT 49.880 121.450 50.020 128.270 ;
        RECT 53.560 126.210 53.700 134.390 ;
        RECT 53.500 125.890 53.760 126.210 ;
        RECT 51.200 122.830 51.460 123.150 ;
        RECT 48.440 121.130 48.700 121.450 ;
        RECT 49.820 121.130 50.080 121.450 ;
        RECT 45.220 120.110 45.480 120.430 ;
        RECT 45.280 116.010 45.420 120.110 ;
        RECT 50.280 118.070 50.540 118.390 ;
        RECT 50.340 116.010 50.480 118.070 ;
        RECT 45.220 115.690 45.480 116.010 ;
        RECT 50.280 115.690 50.540 116.010 ;
        RECT 49.820 115.350 50.080 115.670 ;
        RECT 45.220 115.010 45.480 115.330 ;
        RECT 44.760 112.970 45.020 113.290 ;
        RECT 43.840 112.630 44.100 112.950 ;
        RECT 44.300 112.630 44.560 112.950 ;
        RECT 44.360 110.570 44.500 112.630 ;
        RECT 44.760 112.290 45.020 112.610 ;
        RECT 44.300 110.250 44.560 110.570 ;
        RECT 44.820 109.970 44.960 112.290 ;
        RECT 45.280 110.570 45.420 115.010 ;
        RECT 45.680 114.670 45.940 114.990 ;
        RECT 45.220 110.250 45.480 110.570 ;
        RECT 45.740 110.230 45.880 114.670 ;
        RECT 49.880 113.630 50.020 115.350 ;
        RECT 49.820 113.310 50.080 113.630 ;
        RECT 46.140 112.290 46.400 112.610 ;
        RECT 46.200 111.250 46.340 112.290 ;
        RECT 46.140 110.930 46.400 111.250 ;
        RECT 44.360 109.830 44.960 109.970 ;
        RECT 45.680 109.910 45.940 110.230 ;
        RECT 44.360 107.510 44.500 109.830 ;
        RECT 44.760 109.230 45.020 109.550 ;
        RECT 44.300 107.190 44.560 107.510 ;
        RECT 43.840 104.470 44.100 104.790 ;
        RECT 43.380 102.770 43.640 103.090 ;
        RECT 42.980 102.350 43.580 102.490 ;
        RECT 42.000 101.750 42.260 102.070 ;
        RECT 42.920 101.750 43.180 102.070 ;
        RECT 41.540 101.070 41.800 101.390 ;
        RECT 41.080 100.050 41.340 100.370 ;
        RECT 42.000 93.930 42.260 94.250 ;
        RECT 38.320 93.590 38.580 93.910 ;
        RECT 34.180 90.530 34.440 90.850 ;
        RECT 32.230 89.655 33.770 90.025 ;
        RECT 31.480 86.030 32.080 86.170 ;
        RECT 31.420 83.050 31.680 83.370 ;
        RECT 30.960 82.710 31.220 83.030 ;
        RECT 28.930 81.495 30.470 81.865 ;
        RECT 27.740 79.990 28.000 80.310 ;
        RECT 25.440 76.590 25.700 76.910 ;
        RECT 25.500 74.870 25.640 76.590 ;
        RECT 25.440 74.550 25.700 74.870 ;
        RECT 25.900 73.870 26.160 74.190 ;
        RECT 24.980 71.830 25.240 72.150 ;
        RECT 24.980 69.790 25.240 70.110 ;
        RECT 25.040 67.390 25.180 69.790 ;
        RECT 24.980 67.070 25.240 67.390 ;
        RECT 25.960 66.710 26.100 73.870 ;
        RECT 27.800 73.170 27.940 79.990 ;
        RECT 29.120 79.310 29.380 79.630 ;
        RECT 29.180 77.930 29.320 79.310 ;
        RECT 29.120 77.610 29.380 77.930 ;
        RECT 28.930 76.055 30.470 76.425 ;
        RECT 28.200 74.210 28.460 74.530 ;
        RECT 28.260 73.170 28.400 74.210 ;
        RECT 27.740 72.850 28.000 73.170 ;
        RECT 28.200 72.850 28.460 73.170 ;
        RECT 26.820 72.510 27.080 72.830 ;
        RECT 26.880 69.770 27.020 72.510 ;
        RECT 26.820 69.450 27.080 69.770 ;
        RECT 27.800 67.730 27.940 72.850 ;
        RECT 28.930 70.615 30.470 70.985 ;
        RECT 29.120 68.770 29.380 69.090 ;
        RECT 29.180 67.730 29.320 68.770 ;
        RECT 27.740 67.410 28.000 67.730 ;
        RECT 29.120 67.410 29.380 67.730 ;
        RECT 31.480 67.130 31.620 83.050 ;
        RECT 31.020 66.990 31.620 67.130 ;
        RECT 25.900 66.390 26.160 66.710 ;
        RECT 28.200 66.390 28.460 66.710 ;
        RECT 28.260 65.010 28.400 66.390 ;
        RECT 28.930 65.175 30.470 65.545 ;
        RECT 28.200 64.970 28.460 65.010 ;
        RECT 27.340 64.830 28.460 64.970 ;
        RECT 27.340 64.330 27.480 64.830 ;
        RECT 28.200 64.690 28.460 64.830 ;
        RECT 27.280 64.010 27.540 64.330 ;
        RECT 30.040 63.670 30.300 63.990 ;
        RECT 27.280 63.330 27.540 63.650 ;
        RECT 25.900 62.990 26.160 63.310 ;
        RECT 25.960 61.610 26.100 62.990 ;
        RECT 26.820 61.970 27.080 62.290 ;
        RECT 25.900 61.290 26.160 61.610 ;
        RECT 26.360 59.250 26.620 59.570 ;
        RECT 24.980 58.910 25.240 59.230 ;
        RECT 24.120 56.790 24.720 56.930 ;
        RECT 21.745 55.995 22.030 56.170 ;
        RECT 21.745 55.850 22.005 55.995 ;
        RECT 23.140 55.850 23.400 56.170 ;
        RECT 22.680 55.170 22.940 55.490 ;
        RECT 22.740 54.130 22.880 55.170 ;
        RECT 22.680 53.810 22.940 54.130 ;
        RECT 23.200 51.170 23.340 55.850 ;
        RECT 24.120 55.150 24.260 56.790 ;
        RECT 25.040 56.170 25.180 58.910 ;
        RECT 26.420 56.170 26.560 59.250 ;
        RECT 26.880 58.550 27.020 61.970 ;
        RECT 26.820 58.230 27.080 58.550 ;
        RECT 24.520 55.850 24.780 56.170 ;
        RECT 24.980 55.850 25.240 56.170 ;
        RECT 25.440 55.850 25.700 56.170 ;
        RECT 26.360 55.850 26.620 56.170 ;
        RECT 24.060 54.830 24.320 55.150 ;
        RECT 21.820 51.030 23.340 51.170 ;
        RECT 21.820 48.350 21.960 51.030 ;
        RECT 21.760 48.030 22.020 48.350 ;
        RECT 22.680 47.350 22.940 47.670 ;
        RECT 21.760 46.670 22.020 46.990 ;
        RECT 21.820 44.125 21.960 46.670 ;
        RECT 22.740 45.630 22.880 47.350 ;
        RECT 23.600 45.650 23.860 45.970 ;
        RECT 22.680 45.310 22.940 45.630 ;
        RECT 21.750 43.755 22.030 44.125 ;
        RECT 23.140 43.950 23.400 44.270 ;
        RECT 22.680 41.230 22.940 41.550 ;
        RECT 22.740 40.725 22.880 41.230 ;
        RECT 22.670 40.355 22.950 40.725 ;
        RECT 22.220 39.870 22.480 40.190 ;
        RECT 21.300 38.510 21.560 38.830 ;
        RECT 21.760 37.490 22.020 37.810 ;
        RECT 21.300 36.130 21.560 36.450 ;
        RECT 21.360 35.090 21.500 36.130 ;
        RECT 21.300 34.770 21.560 35.090 ;
        RECT 20.840 31.710 21.100 32.030 ;
        RECT 21.820 31.090 21.960 37.490 ;
        RECT 22.280 36.110 22.420 39.870 ;
        RECT 22.680 39.760 22.940 39.850 ;
        RECT 23.200 39.760 23.340 43.950 ;
        RECT 23.660 42.230 23.800 45.650 ;
        RECT 23.600 41.910 23.860 42.230 ;
        RECT 22.680 39.620 23.340 39.760 ;
        RECT 22.680 39.530 22.940 39.620 ;
        RECT 22.680 38.510 22.940 38.830 ;
        RECT 22.220 35.790 22.480 36.110 ;
        RECT 22.280 31.690 22.420 35.790 ;
        RECT 22.740 34.410 22.880 38.510 ;
        RECT 23.200 37.810 23.340 39.620 ;
        RECT 23.140 37.490 23.400 37.810 ;
        RECT 22.680 34.090 22.940 34.410 ;
        RECT 23.140 34.090 23.400 34.410 ;
        RECT 23.200 32.030 23.340 34.090 ;
        RECT 23.140 31.710 23.400 32.030 ;
        RECT 22.220 31.370 22.480 31.690 ;
        RECT 21.820 30.950 22.420 31.090 ;
        RECT 21.760 30.350 22.020 30.670 ;
        RECT 21.820 29.310 21.960 30.350 ;
        RECT 21.760 28.990 22.020 29.310 ;
        RECT 22.280 25.230 22.420 30.950 ;
        RECT 22.680 27.630 22.940 27.950 ;
        RECT 22.740 25.910 22.880 27.630 ;
        RECT 22.680 25.590 22.940 25.910 ;
        RECT 22.220 24.910 22.480 25.230 ;
        RECT 22.280 23.870 22.420 24.910 ;
        RECT 22.220 23.550 22.480 23.870 ;
        RECT 21.760 23.210 22.020 23.530 ;
        RECT 19.920 20.490 20.180 20.810 ;
        RECT 20.380 19.470 20.640 19.790 ;
        RECT 20.840 19.470 21.100 19.790 ;
        RECT 20.440 11.370 20.580 19.470 ;
        RECT 20.900 18.090 21.040 19.470 ;
        RECT 21.820 18.770 21.960 23.210 ;
        RECT 22.740 20.470 22.880 25.590 ;
        RECT 23.200 21.150 23.340 31.710 ;
        RECT 24.060 31.030 24.320 31.350 ;
        RECT 24.120 29.650 24.260 31.030 ;
        RECT 24.060 29.330 24.320 29.650 ;
        RECT 24.580 23.610 24.720 55.850 ;
        RECT 24.980 55.170 25.240 55.490 ;
        RECT 25.040 42.650 25.180 55.170 ;
        RECT 25.500 53.110 25.640 55.850 ;
        RECT 25.440 52.790 25.700 53.110 ;
        RECT 25.500 51.170 25.640 52.790 ;
        RECT 25.500 51.030 26.100 51.170 ;
        RECT 25.440 48.030 25.700 48.350 ;
        RECT 25.500 44.950 25.640 48.030 ;
        RECT 25.440 44.630 25.700 44.950 ;
        RECT 25.960 42.910 26.100 51.030 ;
        RECT 26.420 47.670 26.560 55.850 ;
        RECT 26.880 51.070 27.020 58.230 ;
        RECT 27.340 56.510 27.480 63.330 ;
        RECT 28.200 62.990 28.460 63.310 ;
        RECT 29.580 62.990 29.840 63.310 ;
        RECT 27.740 60.270 28.000 60.590 ;
        RECT 27.800 58.550 27.940 60.270 ;
        RECT 28.260 59.570 28.400 62.990 ;
        RECT 29.640 62.290 29.780 62.990 ;
        RECT 29.580 61.970 29.840 62.290 ;
        RECT 30.100 60.500 30.240 63.670 ;
        RECT 31.020 60.840 31.160 66.990 ;
        RECT 31.420 66.390 31.680 66.710 ;
        RECT 31.480 63.990 31.620 66.390 ;
        RECT 31.940 64.970 32.080 86.030 ;
        RECT 32.230 84.215 33.770 84.585 ;
        RECT 34.240 81.410 34.380 90.530 ;
        RECT 36.940 88.150 37.200 88.470 ;
        RECT 34.640 84.750 34.900 85.070 ;
        RECT 34.700 83.370 34.840 84.750 ;
        RECT 34.640 83.050 34.900 83.370 ;
        RECT 34.700 82.350 34.840 83.050 ;
        RECT 34.640 82.030 34.900 82.350 ;
        RECT 34.240 81.270 34.840 81.410 ;
        RECT 32.230 78.775 33.770 79.145 ;
        RECT 32.230 73.335 33.770 73.705 ;
        RECT 34.180 68.430 34.440 68.750 ;
        RECT 32.230 67.895 33.770 68.265 ;
        RECT 34.240 65.010 34.380 68.430 ;
        RECT 31.940 64.830 33.920 64.970 ;
        RECT 31.420 63.670 31.680 63.990 ;
        RECT 31.480 62.290 31.620 63.670 ;
        RECT 33.780 63.560 33.920 64.830 ;
        RECT 34.180 64.690 34.440 65.010 ;
        RECT 34.700 64.970 34.840 81.270 ;
        RECT 35.560 80.670 35.820 80.990 ;
        RECT 35.620 79.630 35.760 80.670 ;
        RECT 35.560 79.310 35.820 79.630 ;
        RECT 35.620 78.610 35.760 79.310 ;
        RECT 35.560 78.290 35.820 78.610 ;
        RECT 34.700 64.830 35.300 64.970 ;
        RECT 34.640 64.350 34.900 64.670 ;
        RECT 33.780 63.420 34.380 63.560 ;
        RECT 31.880 62.990 32.140 63.310 ;
        RECT 31.420 61.970 31.680 62.290 ;
        RECT 31.020 60.700 31.620 60.840 ;
        RECT 30.100 60.360 31.160 60.500 ;
        RECT 28.930 59.735 30.470 60.105 ;
        RECT 28.200 59.250 28.460 59.570 ;
        RECT 31.020 59.230 31.160 60.360 ;
        RECT 30.960 58.910 31.220 59.230 ;
        RECT 27.740 58.230 28.000 58.550 ;
        RECT 29.120 57.890 29.380 58.210 ;
        RECT 28.660 57.550 28.920 57.870 ;
        RECT 27.280 56.190 27.540 56.510 ;
        RECT 28.720 56.170 28.860 57.550 ;
        RECT 29.180 56.510 29.320 57.890 ;
        RECT 31.480 57.870 31.620 60.700 ;
        RECT 31.940 58.890 32.080 62.990 ;
        RECT 32.230 62.455 33.770 62.825 ;
        RECT 32.340 61.630 32.600 61.950 ;
        RECT 31.880 58.570 32.140 58.890 ;
        RECT 32.400 58.550 32.540 61.630 ;
        RECT 33.260 61.290 33.520 61.610 ;
        RECT 33.320 59.570 33.460 61.290 ;
        RECT 33.260 59.250 33.520 59.570 ;
        RECT 32.340 58.230 32.600 58.550 ;
        RECT 31.420 57.550 31.680 57.870 ;
        RECT 32.230 57.015 33.770 57.385 ;
        RECT 29.120 56.190 29.380 56.510 ;
        RECT 28.660 56.080 28.920 56.170 ;
        RECT 28.260 55.940 28.920 56.080 ;
        RECT 28.260 51.410 28.400 55.940 ;
        RECT 28.660 55.850 28.920 55.940 ;
        RECT 30.960 55.850 31.220 56.170 ;
        RECT 28.930 54.295 30.470 54.665 ;
        RECT 28.660 52.450 28.920 52.770 ;
        RECT 28.200 51.090 28.460 51.410 ;
        RECT 26.820 50.750 27.080 51.070 ;
        RECT 26.880 48.090 27.020 50.750 ;
        RECT 28.720 50.390 28.860 52.450 ;
        RECT 31.020 50.390 31.160 55.850 ;
        RECT 31.420 54.830 31.680 55.150 ;
        RECT 31.480 50.390 31.620 54.830 ;
        RECT 32.340 52.850 32.600 53.110 ;
        RECT 31.940 52.790 32.600 52.850 ;
        RECT 31.940 52.710 32.540 52.790 ;
        RECT 28.660 50.070 28.920 50.390 ;
        RECT 30.960 50.070 31.220 50.390 ;
        RECT 31.420 50.070 31.680 50.390 ;
        RECT 28.200 49.390 28.460 49.710 ;
        RECT 26.880 47.950 27.480 48.090 ;
        RECT 26.360 47.350 26.620 47.670 ;
        RECT 25.040 42.510 25.640 42.650 ;
        RECT 25.900 42.590 26.160 42.910 ;
        RECT 24.980 41.910 25.240 42.230 ;
        RECT 25.040 26.930 25.180 41.910 ;
        RECT 25.500 31.770 25.640 42.510 ;
        RECT 26.420 39.510 26.560 47.350 ;
        RECT 27.340 45.290 27.480 47.950 ;
        RECT 28.260 47.670 28.400 49.390 ;
        RECT 28.930 48.855 30.470 49.225 ;
        RECT 30.040 48.370 30.300 48.690 ;
        RECT 29.580 47.690 29.840 48.010 ;
        RECT 28.200 47.350 28.460 47.670 ;
        RECT 29.640 45.290 29.780 47.690 ;
        RECT 30.100 45.290 30.240 48.370 ;
        RECT 31.020 48.010 31.160 50.070 ;
        RECT 30.960 47.690 31.220 48.010 ;
        RECT 31.420 47.350 31.680 47.670 ;
        RECT 27.280 44.970 27.540 45.290 ;
        RECT 29.580 44.970 29.840 45.290 ;
        RECT 30.040 44.970 30.300 45.290 ;
        RECT 26.820 44.630 27.080 44.950 ;
        RECT 26.360 39.190 26.620 39.510 ;
        RECT 26.880 36.790 27.020 44.630 ;
        RECT 27.340 43.160 27.480 44.970 ;
        RECT 30.960 44.630 31.220 44.950 ;
        RECT 28.930 43.415 30.470 43.785 ;
        RECT 31.020 43.250 31.160 44.630 ;
        RECT 27.340 43.020 28.860 43.160 ;
        RECT 27.740 41.910 28.000 42.230 ;
        RECT 26.820 36.470 27.080 36.790 ;
        RECT 26.820 35.790 27.080 36.110 ;
        RECT 26.880 34.750 27.020 35.790 ;
        RECT 26.820 34.430 27.080 34.750 ;
        RECT 27.280 33.070 27.540 33.390 ;
        RECT 25.500 31.630 26.100 31.770 ;
        RECT 25.440 31.030 25.700 31.350 ;
        RECT 25.500 28.970 25.640 31.030 ;
        RECT 25.440 28.650 25.700 28.970 ;
        RECT 24.980 26.610 25.240 26.930 ;
        RECT 25.440 25.590 25.700 25.910 ;
        RECT 25.500 23.725 25.640 25.590 ;
        RECT 24.580 23.470 25.180 23.610 ;
        RECT 23.600 22.530 23.860 22.850 ;
        RECT 24.520 22.530 24.780 22.850 ;
        RECT 23.140 20.830 23.400 21.150 ;
        RECT 22.680 20.150 22.940 20.470 ;
        RECT 21.760 18.450 22.020 18.770 ;
        RECT 20.840 17.770 21.100 18.090 ;
        RECT 21.820 16.050 21.960 18.450 ;
        RECT 23.660 18.090 23.800 22.530 ;
        RECT 24.060 20.150 24.320 20.470 ;
        RECT 23.600 17.770 23.860 18.090 ;
        RECT 24.120 16.050 24.260 20.150 ;
        RECT 21.760 15.730 22.020 16.050 ;
        RECT 24.060 15.730 24.320 16.050 ;
        RECT 24.580 12.730 24.720 22.530 ;
        RECT 25.040 22.510 25.180 23.470 ;
        RECT 25.430 23.355 25.710 23.725 ;
        RECT 25.440 23.210 25.700 23.355 ;
        RECT 24.980 22.190 25.240 22.510 ;
        RECT 25.960 21.490 26.100 31.630 ;
        RECT 27.340 31.350 27.480 33.070 ;
        RECT 27.280 31.030 27.540 31.350 ;
        RECT 27.340 29.650 27.480 31.030 ;
        RECT 27.280 29.330 27.540 29.650 ;
        RECT 26.360 23.210 26.620 23.530 ;
        RECT 25.900 21.170 26.160 21.490 ;
        RECT 26.420 17.070 26.560 23.210 ;
        RECT 27.340 20.470 27.480 29.330 ;
        RECT 27.800 26.930 27.940 41.910 ;
        RECT 28.720 40.190 28.860 43.020 ;
        RECT 30.960 42.930 31.220 43.250 ;
        RECT 30.500 42.250 30.760 42.570 ;
        RECT 29.120 41.910 29.380 42.230 ;
        RECT 28.660 39.870 28.920 40.190 ;
        RECT 29.180 39.850 29.320 41.910 ;
        RECT 30.560 40.190 30.700 42.250 ;
        RECT 30.960 41.570 31.220 41.890 ;
        RECT 30.500 39.870 30.760 40.190 ;
        RECT 31.020 39.850 31.160 41.570 ;
        RECT 29.120 39.530 29.380 39.850 ;
        RECT 30.960 39.530 31.220 39.850 ;
        RECT 30.960 38.510 31.220 38.830 ;
        RECT 28.930 37.975 30.470 38.345 ;
        RECT 30.040 36.470 30.300 36.790 ;
        RECT 30.500 36.470 30.760 36.790 ;
        RECT 28.660 36.130 28.920 36.450 ;
        RECT 28.720 34.410 28.860 36.130 ;
        RECT 30.100 34.750 30.240 36.470 ;
        RECT 30.560 35.090 30.700 36.470 ;
        RECT 31.020 36.110 31.160 38.510 ;
        RECT 31.480 36.700 31.620 47.350 ;
        RECT 31.940 40.530 32.080 52.710 ;
        RECT 32.230 51.575 33.770 51.945 ;
        RECT 33.260 51.090 33.520 51.410 ;
        RECT 33.720 51.090 33.980 51.410 ;
        RECT 33.320 47.330 33.460 51.090 ;
        RECT 33.780 47.525 33.920 51.090 ;
        RECT 33.260 47.010 33.520 47.330 ;
        RECT 33.710 47.155 33.990 47.525 ;
        RECT 32.230 46.135 33.770 46.505 ;
        RECT 34.240 42.230 34.380 63.420 ;
        RECT 34.700 55.060 34.840 64.350 ;
        RECT 35.160 55.570 35.300 64.830 ;
        RECT 35.620 61.950 35.760 78.290 ;
        RECT 36.480 68.430 36.740 68.750 ;
        RECT 36.540 63.650 36.680 68.430 ;
        RECT 36.480 63.330 36.740 63.650 ;
        RECT 35.560 61.860 35.820 61.950 ;
        RECT 35.560 61.720 36.220 61.860 ;
        RECT 35.560 61.630 35.820 61.720 ;
        RECT 35.560 60.270 35.820 60.590 ;
        RECT 35.620 56.510 35.760 60.270 ;
        RECT 35.560 56.190 35.820 56.510 ;
        RECT 35.160 55.430 35.760 55.570 ;
        RECT 35.100 55.060 35.360 55.150 ;
        RECT 34.700 54.920 35.360 55.060 ;
        RECT 34.700 52.770 34.840 54.920 ;
        RECT 35.100 54.830 35.360 54.920 ;
        RECT 35.620 54.210 35.760 55.430 ;
        RECT 35.160 54.070 35.760 54.210 ;
        RECT 34.640 52.450 34.900 52.770 ;
        RECT 34.700 50.730 34.840 52.450 ;
        RECT 34.640 50.410 34.900 50.730 ;
        RECT 35.160 47.670 35.300 54.070 ;
        RECT 36.080 51.410 36.220 61.720 ;
        RECT 37.000 56.850 37.140 88.150 ;
        RECT 38.380 80.650 38.520 93.590 ;
        RECT 42.060 91.530 42.200 93.930 ;
        RECT 38.780 91.210 39.040 91.530 ;
        RECT 42.000 91.210 42.260 91.530 ;
        RECT 38.840 89.490 38.980 91.210 ;
        RECT 41.540 90.190 41.800 90.510 ;
        RECT 41.600 89.490 41.740 90.190 ;
        RECT 42.980 89.490 43.120 101.750 ;
        RECT 43.440 99.470 43.580 102.350 ;
        RECT 43.900 100.030 44.040 104.470 ;
        RECT 43.840 99.710 44.100 100.030 ;
        RECT 44.360 99.470 44.500 107.190 ;
        RECT 44.820 102.410 44.960 109.230 ;
        RECT 45.220 107.190 45.480 107.510 ;
        RECT 45.680 107.190 45.940 107.510 ;
        RECT 45.280 105.810 45.420 107.190 ;
        RECT 45.220 105.490 45.480 105.810 ;
        RECT 44.760 102.090 45.020 102.410 ;
        RECT 45.280 102.070 45.420 105.490 ;
        RECT 45.740 102.070 45.880 107.190 ;
        RECT 47.060 106.850 47.320 107.170 ;
        RECT 49.820 106.850 50.080 107.170 ;
        RECT 46.600 104.810 46.860 105.130 ;
        RECT 46.660 103.090 46.800 104.810 ;
        RECT 46.600 102.770 46.860 103.090 ;
        RECT 45.220 101.750 45.480 102.070 ;
        RECT 45.680 101.750 45.940 102.070 ;
        RECT 45.280 99.470 45.420 101.750 ;
        RECT 43.440 99.330 44.500 99.470 ;
        RECT 44.360 94.590 44.500 99.330 ;
        RECT 44.820 99.330 45.420 99.470 ;
        RECT 46.140 99.370 46.400 99.690 ;
        RECT 44.300 94.270 44.560 94.590 ;
        RECT 38.780 89.170 39.040 89.490 ;
        RECT 41.540 89.170 41.800 89.490 ;
        RECT 42.920 89.170 43.180 89.490 ;
        RECT 44.360 88.810 44.500 94.270 ;
        RECT 44.820 93.140 44.960 99.330 ;
        RECT 45.220 96.650 45.480 96.970 ;
        RECT 45.280 94.930 45.420 96.650 ;
        RECT 45.220 94.610 45.480 94.930 ;
        RECT 45.220 93.140 45.480 93.230 ;
        RECT 44.820 93.000 45.480 93.140 ;
        RECT 45.220 92.910 45.480 93.000 ;
        RECT 44.300 88.490 44.560 88.810 ;
        RECT 44.360 86.430 44.500 88.490 ;
        RECT 45.280 86.770 45.420 92.910 ;
        RECT 45.220 86.450 45.480 86.770 ;
        RECT 44.300 86.110 44.560 86.430 ;
        RECT 45.680 85.090 45.940 85.410 ;
        RECT 40.160 84.750 40.420 85.070 ;
        RECT 40.220 80.650 40.360 84.750 ;
        RECT 45.740 84.050 45.880 85.090 ;
        RECT 45.680 83.730 45.940 84.050 ;
        RECT 42.460 83.390 42.720 83.710 ;
        RECT 41.080 83.050 41.340 83.370 ;
        RECT 41.140 81.330 41.280 83.050 ;
        RECT 41.080 81.010 41.340 81.330 ;
        RECT 38.320 80.330 38.580 80.650 ;
        RECT 40.160 80.330 40.420 80.650 ;
        RECT 42.000 79.990 42.260 80.310 ;
        RECT 41.080 77.610 41.340 77.930 ;
        RECT 41.140 75.890 41.280 77.610 ;
        RECT 41.080 75.570 41.340 75.890 ;
        RECT 42.060 75.550 42.200 79.990 ;
        RECT 42.520 78.270 42.660 83.390 ;
        RECT 46.200 80.650 46.340 99.370 ;
        RECT 47.120 99.010 47.260 106.850 ;
        RECT 49.880 104.110 50.020 106.850 ;
        RECT 50.740 106.510 51.000 106.830 ;
        RECT 49.820 103.790 50.080 104.110 ;
        RECT 50.800 103.090 50.940 106.510 ;
        RECT 50.740 102.770 51.000 103.090 ;
        RECT 48.900 99.710 49.160 100.030 ;
        RECT 48.440 99.370 48.700 99.690 ;
        RECT 47.060 98.690 47.320 99.010 ;
        RECT 47.120 90.850 47.260 98.690 ;
        RECT 48.500 97.650 48.640 99.370 ;
        RECT 48.440 97.330 48.700 97.650 ;
        RECT 48.440 92.910 48.700 93.230 ;
        RECT 48.500 91.190 48.640 92.910 ;
        RECT 48.440 90.870 48.700 91.190 ;
        RECT 47.060 90.530 47.320 90.850 ;
        RECT 46.600 84.750 46.860 85.070 ;
        RECT 46.660 83.030 46.800 84.750 ;
        RECT 47.120 83.370 47.260 90.530 ;
        RECT 47.980 88.490 48.240 88.810 ;
        RECT 48.040 84.050 48.180 88.490 ;
        RECT 48.440 86.110 48.700 86.430 ;
        RECT 47.980 83.730 48.240 84.050 ;
        RECT 47.060 83.050 47.320 83.370 ;
        RECT 46.600 82.710 46.860 83.030 ;
        RECT 48.500 80.650 48.640 86.110 ;
        RECT 48.960 83.710 49.100 99.710 ;
        RECT 50.740 96.990 51.000 97.310 ;
        RECT 49.360 91.890 49.620 92.210 ;
        RECT 49.420 89.490 49.560 91.890 ;
        RECT 49.820 90.190 50.080 90.510 ;
        RECT 49.360 89.170 49.620 89.490 ;
        RECT 49.880 88.810 50.020 90.190 ;
        RECT 49.820 88.490 50.080 88.810 ;
        RECT 49.360 87.810 49.620 88.130 ;
        RECT 49.420 86.430 49.560 87.810 ;
        RECT 50.280 87.470 50.540 87.790 ;
        RECT 50.340 86.770 50.480 87.470 ;
        RECT 50.280 86.450 50.540 86.770 ;
        RECT 49.360 86.110 49.620 86.430 ;
        RECT 50.340 85.410 50.480 86.450 ;
        RECT 50.280 85.090 50.540 85.410 ;
        RECT 49.360 84.750 49.620 85.070 ;
        RECT 49.420 83.710 49.560 84.750 ;
        RECT 48.900 83.390 49.160 83.710 ;
        RECT 49.360 83.390 49.620 83.710 ;
        RECT 48.960 83.030 49.100 83.390 ;
        RECT 48.900 82.710 49.160 83.030 ;
        RECT 49.360 82.030 49.620 82.350 ;
        RECT 49.420 81.330 49.560 82.030 ;
        RECT 49.360 81.010 49.620 81.330 ;
        RECT 46.140 80.330 46.400 80.650 ;
        RECT 48.440 80.330 48.700 80.650 ;
        RECT 42.920 79.310 43.180 79.630 ;
        RECT 44.760 79.310 45.020 79.630 ;
        RECT 42.460 77.950 42.720 78.270 ;
        RECT 42.000 75.230 42.260 75.550 ;
        RECT 42.520 74.870 42.660 77.950 ;
        RECT 42.460 74.550 42.720 74.870 ;
        RECT 37.860 74.210 38.120 74.530 ;
        RECT 37.920 72.150 38.060 74.210 ;
        RECT 42.520 72.830 42.660 74.550 ;
        RECT 39.700 72.510 39.960 72.830 ;
        RECT 41.080 72.510 41.340 72.830 ;
        RECT 42.460 72.510 42.720 72.830 ;
        RECT 37.860 71.830 38.120 72.150 ;
        RECT 36.940 56.530 37.200 56.850 ;
        RECT 36.020 51.090 36.280 51.410 ;
        RECT 37.400 48.600 37.660 48.690 ;
        RECT 37.920 48.600 38.060 71.830 ;
        RECT 38.320 68.430 38.580 68.750 ;
        RECT 38.780 68.430 39.040 68.750 ;
        RECT 38.380 67.730 38.520 68.430 ;
        RECT 38.320 67.410 38.580 67.730 ;
        RECT 38.840 64.970 38.980 68.430 ;
        RECT 37.400 48.460 38.060 48.600 ;
        RECT 37.400 48.370 37.660 48.460 ;
        RECT 35.100 47.350 35.360 47.670 ;
        RECT 34.640 47.010 34.900 47.330 ;
        RECT 34.700 43.160 34.840 47.010 ;
        RECT 34.700 43.020 35.300 43.160 ;
        RECT 34.640 42.250 34.900 42.570 ;
        RECT 34.180 41.910 34.440 42.230 ;
        RECT 32.230 40.695 33.770 41.065 ;
        RECT 31.880 40.210 32.140 40.530 ;
        RECT 34.700 39.850 34.840 42.250 ;
        RECT 35.160 39.930 35.300 43.020 ;
        RECT 37.920 42.230 38.060 48.460 ;
        RECT 38.380 64.830 38.980 64.970 ;
        RECT 38.380 42.910 38.520 64.830 ;
        RECT 39.240 57.890 39.500 58.210 ;
        RECT 39.300 56.850 39.440 57.890 ;
        RECT 39.240 56.530 39.500 56.850 ;
        RECT 39.760 51.070 39.900 72.510 ;
        RECT 41.140 69.430 41.280 72.510 ;
        RECT 41.080 69.110 41.340 69.430 ;
        RECT 40.620 64.690 40.880 65.010 ;
        RECT 40.680 59.230 40.820 64.690 ;
        RECT 41.140 63.990 41.280 69.110 ;
        RECT 41.080 63.670 41.340 63.990 ;
        RECT 41.140 61.610 41.280 63.670 ;
        RECT 41.080 61.290 41.340 61.610 ;
        RECT 40.620 58.910 40.880 59.230 ;
        RECT 41.140 58.550 41.280 61.290 ;
        RECT 42.980 59.570 43.120 79.310 ;
        RECT 44.820 75.210 44.960 79.310 ;
        RECT 46.200 78.610 46.340 80.330 ;
        RECT 48.500 78.610 48.640 80.330 ;
        RECT 46.140 78.290 46.400 78.610 ;
        RECT 48.440 78.290 48.700 78.610 ;
        RECT 44.760 74.890 45.020 75.210 ;
        RECT 47.520 74.550 47.780 74.870 ;
        RECT 43.380 67.410 43.640 67.730 ;
        RECT 43.440 67.050 43.580 67.410 ;
        RECT 43.380 66.730 43.640 67.050 ;
        RECT 43.840 66.730 44.100 67.050 ;
        RECT 44.760 66.730 45.020 67.050 ;
        RECT 43.440 65.010 43.580 66.730 ;
        RECT 43.900 65.885 44.040 66.730 ;
        RECT 43.830 65.515 44.110 65.885 ;
        RECT 43.380 64.690 43.640 65.010 ;
        RECT 44.820 64.970 44.960 66.730 ;
        RECT 47.580 66.030 47.720 74.550 ;
        RECT 48.440 73.870 48.700 74.190 ;
        RECT 48.500 67.730 48.640 73.870 ;
        RECT 48.900 69.110 49.160 69.430 ;
        RECT 48.440 67.410 48.700 67.730 ;
        RECT 48.440 66.390 48.700 66.710 ;
        RECT 47.520 65.710 47.780 66.030 ;
        RECT 44.820 64.830 46.800 64.970 ;
        RECT 44.760 62.990 45.020 63.310 ;
        RECT 44.820 61.950 44.960 62.990 ;
        RECT 44.760 61.630 45.020 61.950 ;
        RECT 42.920 59.250 43.180 59.570 ;
        RECT 41.080 58.230 41.340 58.550 ;
        RECT 44.300 57.550 44.560 57.870 ;
        RECT 44.360 56.170 44.500 57.550 ;
        RECT 44.300 55.850 44.560 56.170 ;
        RECT 42.000 55.510 42.260 55.830 ;
        RECT 42.060 54.130 42.200 55.510 ;
        RECT 42.000 53.810 42.260 54.130 ;
        RECT 39.700 50.750 39.960 51.070 ;
        RECT 38.780 45.650 39.040 45.970 ;
        RECT 38.840 44.610 38.980 45.650 ;
        RECT 39.760 45.630 39.900 50.750 ;
        RECT 41.080 50.410 41.340 50.730 ;
        RECT 41.540 50.410 41.800 50.730 ;
        RECT 42.460 50.640 42.720 50.730 ;
        RECT 42.460 50.500 43.120 50.640 ;
        RECT 42.460 50.410 42.720 50.500 ;
        RECT 40.160 47.010 40.420 47.330 ;
        RECT 39.700 45.310 39.960 45.630 ;
        RECT 38.780 44.290 39.040 44.610 ;
        RECT 38.320 42.590 38.580 42.910 ;
        RECT 37.860 42.140 38.120 42.230 ;
        RECT 37.460 42.000 38.120 42.140 ;
        RECT 34.640 39.530 34.900 39.850 ;
        RECT 35.160 39.790 35.760 39.930 ;
        RECT 34.700 37.210 34.840 39.530 ;
        RECT 35.100 39.190 35.360 39.510 ;
        RECT 34.240 37.070 34.840 37.210 ;
        RECT 34.240 36.790 34.380 37.070 ;
        RECT 35.160 36.790 35.300 39.190 ;
        RECT 31.880 36.700 32.140 36.790 ;
        RECT 31.480 36.560 32.140 36.700 ;
        RECT 31.880 36.470 32.140 36.560 ;
        RECT 34.180 36.470 34.440 36.790 ;
        RECT 34.640 36.470 34.900 36.790 ;
        RECT 35.100 36.470 35.360 36.790 ;
        RECT 30.960 35.790 31.220 36.110 ;
        RECT 31.420 35.790 31.680 36.110 ;
        RECT 30.500 34.770 30.760 35.090 ;
        RECT 30.960 34.770 31.220 35.090 ;
        RECT 30.040 34.490 30.300 34.750 ;
        RECT 31.020 34.490 31.160 34.770 ;
        RECT 30.040 34.430 31.160 34.490 ;
        RECT 28.660 34.090 28.920 34.410 ;
        RECT 30.100 34.350 31.160 34.430 ;
        RECT 31.480 34.410 31.620 35.790 ;
        RECT 32.230 35.255 33.770 35.625 ;
        RECT 34.180 34.770 34.440 35.090 ;
        RECT 31.420 34.090 31.680 34.410 ;
        RECT 28.720 33.810 28.860 34.090 ;
        RECT 28.260 33.670 28.860 33.810 ;
        RECT 28.260 28.970 28.400 33.670 ;
        RECT 31.880 33.070 32.140 33.390 ;
        RECT 28.930 32.535 30.470 32.905 ;
        RECT 28.200 28.650 28.460 28.970 ;
        RECT 31.420 28.650 31.680 28.970 ;
        RECT 27.740 26.610 28.000 26.930 ;
        RECT 28.260 26.330 28.400 28.650 ;
        RECT 30.960 27.630 31.220 27.950 ;
        RECT 28.930 27.095 30.470 27.465 ;
        RECT 27.800 26.190 28.400 26.330 ;
        RECT 27.800 23.870 27.940 26.190 ;
        RECT 31.020 25.910 31.160 27.630 ;
        RECT 28.200 25.590 28.460 25.910 ;
        RECT 30.960 25.590 31.220 25.910 ;
        RECT 27.740 23.550 28.000 23.870 ;
        RECT 27.280 20.150 27.540 20.470 ;
        RECT 27.280 17.770 27.540 18.090 ;
        RECT 27.340 17.490 27.480 17.770 ;
        RECT 27.800 17.490 27.940 23.550 ;
        RECT 28.260 18.090 28.400 25.590 ;
        RECT 30.960 24.910 31.220 25.230 ;
        RECT 31.020 23.870 31.160 24.910 ;
        RECT 31.480 24.210 31.620 28.650 ;
        RECT 31.420 23.890 31.680 24.210 ;
        RECT 30.960 23.550 31.220 23.870 ;
        RECT 31.940 23.610 32.080 33.070 ;
        RECT 32.230 29.815 33.770 30.185 ;
        RECT 33.720 28.880 33.980 28.970 ;
        RECT 34.240 28.880 34.380 34.770 ;
        RECT 34.700 31.690 34.840 36.470 ;
        RECT 35.100 34.430 35.360 34.750 ;
        RECT 34.640 31.370 34.900 31.690 ;
        RECT 34.700 28.970 34.840 31.370 ;
        RECT 33.720 28.740 34.380 28.880 ;
        RECT 33.720 28.650 33.980 28.740 ;
        RECT 32.230 24.375 33.770 24.745 ;
        RECT 28.930 21.655 30.470 22.025 ;
        RECT 29.110 20.635 29.390 21.005 ;
        RECT 29.180 20.470 29.320 20.635 ;
        RECT 29.120 20.150 29.380 20.470 ;
        RECT 28.660 19.470 28.920 19.790 ;
        RECT 30.500 19.470 30.760 19.790 ;
        RECT 28.720 18.770 28.860 19.470 ;
        RECT 28.660 18.450 28.920 18.770 ;
        RECT 30.560 18.430 30.700 19.470 ;
        RECT 30.500 18.110 30.760 18.430 ;
        RECT 28.200 17.770 28.460 18.090 ;
        RECT 27.340 17.410 28.400 17.490 ;
        RECT 27.340 17.350 28.460 17.410 ;
        RECT 26.360 16.750 26.620 17.070 ;
        RECT 26.420 15.030 26.560 16.750 ;
        RECT 27.340 16.670 27.480 17.350 ;
        RECT 28.200 17.090 28.460 17.350 ;
        RECT 26.880 16.530 27.480 16.670 ;
        RECT 26.360 14.710 26.620 15.030 ;
        RECT 26.880 14.690 27.020 16.530 ;
        RECT 28.930 16.215 30.470 16.585 ;
        RECT 31.020 15.030 31.160 23.550 ;
        RECT 31.480 23.470 32.080 23.610 ;
        RECT 31.480 15.030 31.620 23.470 ;
        RECT 31.880 20.150 32.140 20.470 ;
        RECT 32.800 20.150 33.060 20.470 ;
        RECT 31.940 18.770 32.080 20.150 ;
        RECT 32.860 19.790 33.000 20.150 ;
        RECT 33.720 20.040 33.980 20.130 ;
        RECT 34.240 20.040 34.380 28.740 ;
        RECT 34.640 28.650 34.900 28.970 ;
        RECT 35.160 27.690 35.300 34.430 ;
        RECT 35.620 28.970 35.760 39.790 ;
        RECT 35.560 28.880 35.820 28.970 ;
        RECT 35.560 28.740 36.220 28.880 ;
        RECT 35.560 28.650 35.820 28.740 ;
        RECT 35.560 27.970 35.820 28.290 ;
        RECT 35.620 27.690 35.760 27.970 ;
        RECT 35.160 27.550 35.760 27.690 ;
        RECT 35.160 25.650 35.300 27.550 ;
        RECT 35.560 25.650 35.820 25.910 ;
        RECT 35.160 25.590 35.820 25.650 ;
        RECT 35.160 25.510 35.760 25.590 ;
        RECT 35.160 20.470 35.300 25.510 ;
        RECT 36.080 25.230 36.220 28.740 ;
        RECT 36.940 28.650 37.200 28.970 ;
        RECT 36.480 27.630 36.740 27.950 ;
        RECT 36.540 25.570 36.680 27.630 ;
        RECT 36.480 25.250 36.740 25.570 ;
        RECT 36.020 24.910 36.280 25.230 ;
        RECT 35.100 20.150 35.360 20.470 ;
        RECT 33.720 19.900 34.380 20.040 ;
        RECT 33.720 19.810 33.980 19.900 ;
        RECT 32.800 19.470 33.060 19.790 ;
        RECT 32.230 18.935 33.770 19.305 ;
        RECT 31.880 18.450 32.140 18.770 ;
        RECT 35.100 18.110 35.360 18.430 ;
        RECT 35.160 15.030 35.300 18.110 ;
        RECT 37.000 17.750 37.140 28.650 ;
        RECT 37.460 28.290 37.600 42.000 ;
        RECT 37.860 41.910 38.120 42.000 ;
        RECT 38.840 40.190 38.980 44.290 ;
        RECT 40.220 43.250 40.360 47.010 ;
        RECT 41.140 46.990 41.280 50.410 ;
        RECT 41.600 50.050 41.740 50.410 ;
        RECT 41.540 49.730 41.800 50.050 ;
        RECT 42.460 49.730 42.720 50.050 ;
        RECT 41.600 48.690 41.740 49.730 ;
        RECT 41.540 48.370 41.800 48.690 ;
        RECT 42.520 47.670 42.660 49.730 ;
        RECT 42.460 47.350 42.720 47.670 ;
        RECT 41.080 46.670 41.340 46.990 ;
        RECT 41.540 45.310 41.800 45.630 ;
        RECT 40.160 42.930 40.420 43.250 ;
        RECT 41.600 42.230 41.740 45.310 ;
        RECT 42.520 45.290 42.660 47.350 ;
        RECT 42.460 44.970 42.720 45.290 ;
        RECT 41.540 41.910 41.800 42.230 ;
        RECT 38.780 39.870 39.040 40.190 ;
        RECT 40.620 36.470 40.880 36.790 ;
        RECT 37.860 35.790 38.120 36.110 ;
        RECT 37.920 34.750 38.060 35.790 ;
        RECT 37.860 34.430 38.120 34.750 ;
        RECT 37.400 27.970 37.660 28.290 ;
        RECT 37.460 25.570 37.600 27.970 ;
        RECT 37.400 25.250 37.660 25.570 ;
        RECT 36.940 17.430 37.200 17.750 ;
        RECT 36.940 15.390 37.200 15.710 ;
        RECT 30.960 14.710 31.220 15.030 ;
        RECT 31.420 14.710 31.680 15.030 ;
        RECT 35.100 14.710 35.360 15.030 ;
        RECT 26.820 14.370 27.080 14.690 ;
        RECT 27.280 14.030 27.540 14.350 ;
        RECT 30.500 14.030 30.760 14.350 ;
        RECT 33.720 14.260 33.980 14.350 ;
        RECT 33.720 14.120 34.380 14.260 ;
        RECT 33.720 14.030 33.980 14.120 ;
        RECT 24.120 12.590 24.720 12.730 ;
        RECT 20.440 11.230 21.040 11.370 ;
        RECT 19.460 8.930 19.720 9.250 ;
        RECT 20.900 6.800 21.040 11.230 ;
        RECT 24.120 6.800 24.260 12.590 ;
        RECT 27.340 6.800 27.480 14.030 ;
        RECT 30.560 6.800 30.700 14.030 ;
        RECT 32.230 13.495 33.770 13.865 ;
        RECT 34.240 8.650 34.380 14.120 ;
        RECT 33.780 8.510 34.380 8.650 ;
        RECT 33.780 6.800 33.920 8.510 ;
        RECT 37.000 6.800 37.140 15.390 ;
        RECT 37.920 15.030 38.060 34.430 ;
        RECT 40.680 34.410 40.820 36.470 ;
        RECT 42.460 36.130 42.720 36.450 ;
        RECT 40.620 34.090 40.880 34.410 ;
        RECT 40.680 23.870 40.820 34.090 ;
        RECT 42.000 28.990 42.260 29.310 ;
        RECT 42.060 25.570 42.200 28.990 ;
        RECT 42.520 28.630 42.660 36.130 ;
        RECT 42.980 35.090 43.120 50.500 ;
        RECT 44.300 50.410 44.560 50.730 ;
        RECT 45.220 50.410 45.480 50.730 ;
        RECT 44.360 48.350 44.500 50.410 ;
        RECT 45.280 48.690 45.420 50.410 ;
        RECT 45.220 48.370 45.480 48.690 ;
        RECT 44.300 48.030 44.560 48.350 ;
        RECT 45.220 46.670 45.480 46.990 ;
        RECT 45.280 45.290 45.420 46.670 ;
        RECT 45.220 44.970 45.480 45.290 ;
        RECT 44.760 44.630 45.020 44.950 ;
        RECT 44.820 42.230 44.960 44.630 ;
        RECT 44.760 41.910 45.020 42.230 ;
        RECT 43.840 39.760 44.100 39.850 ;
        RECT 43.840 39.620 44.500 39.760 ;
        RECT 43.840 39.530 44.100 39.620 ;
        RECT 42.920 34.770 43.180 35.090 ;
        RECT 42.920 34.090 43.180 34.410 ;
        RECT 42.980 32.030 43.120 34.090 ;
        RECT 43.380 33.750 43.640 34.070 ;
        RECT 42.920 31.710 43.180 32.030 ;
        RECT 42.920 31.030 43.180 31.350 ;
        RECT 42.980 28.970 43.120 31.030 ;
        RECT 42.920 28.650 43.180 28.970 ;
        RECT 42.460 28.310 42.720 28.630 ;
        RECT 42.980 26.930 43.120 28.650 ;
        RECT 42.920 26.610 43.180 26.930 ;
        RECT 42.000 25.250 42.260 25.570 ;
        RECT 40.620 23.725 40.880 23.870 ;
        RECT 40.610 23.610 40.890 23.725 ;
        RECT 40.610 23.470 41.280 23.610 ;
        RECT 40.610 23.355 40.890 23.470 ;
        RECT 40.620 17.090 40.880 17.410 ;
        RECT 38.780 16.750 39.040 17.070 ;
        RECT 38.840 15.030 38.980 16.750 ;
        RECT 40.680 15.030 40.820 17.090 ;
        RECT 41.140 15.030 41.280 23.470 ;
        RECT 42.000 22.870 42.260 23.190 ;
        RECT 42.060 21.490 42.200 22.870 ;
        RECT 42.000 21.170 42.260 21.490 ;
        RECT 42.060 18.430 42.200 21.170 ;
        RECT 42.980 20.720 43.120 26.610 ;
        RECT 43.440 24.120 43.580 33.750 ;
        RECT 43.840 28.650 44.100 28.970 ;
        RECT 43.900 26.930 44.040 28.650 ;
        RECT 43.840 26.610 44.100 26.930 ;
        RECT 43.840 24.120 44.100 24.210 ;
        RECT 43.440 23.980 44.100 24.120 ;
        RECT 43.840 23.890 44.100 23.980 ;
        RECT 43.900 23.530 44.040 23.890 ;
        RECT 43.840 23.210 44.100 23.530 ;
        RECT 42.520 20.580 43.120 20.720 ;
        RECT 42.000 18.110 42.260 18.430 ;
        RECT 42.520 16.050 42.660 20.580 ;
        RECT 42.920 19.470 43.180 19.790 ;
        RECT 42.980 18.430 43.120 19.470 ;
        RECT 42.920 18.110 43.180 18.430 ;
        RECT 42.460 15.730 42.720 16.050 ;
        RECT 37.860 14.710 38.120 15.030 ;
        RECT 38.780 14.710 39.040 15.030 ;
        RECT 40.620 14.710 40.880 15.030 ;
        RECT 41.080 14.710 41.340 15.030 ;
        RECT 43.900 14.940 44.040 23.210 ;
        RECT 44.360 22.850 44.500 39.620 ;
        RECT 44.820 36.790 44.960 41.910 ;
        RECT 44.760 36.470 45.020 36.790 ;
        RECT 45.680 30.690 45.940 31.010 ;
        RECT 45.740 27.950 45.880 30.690 ;
        RECT 46.140 30.350 46.400 30.670 ;
        RECT 45.680 27.630 45.940 27.950 ;
        RECT 45.740 23.870 45.880 27.630 ;
        RECT 46.200 25.910 46.340 30.350 ;
        RECT 46.140 25.590 46.400 25.910 ;
        RECT 45.680 23.550 45.940 23.870 ;
        RECT 44.300 22.530 44.560 22.850 ;
        RECT 44.300 21.170 44.560 21.490 ;
        RECT 44.360 21.005 44.500 21.170 ;
        RECT 44.290 20.635 44.570 21.005 ;
        RECT 44.360 20.470 44.500 20.635 ;
        RECT 44.300 20.150 44.560 20.470 ;
        RECT 45.220 20.150 45.480 20.470 ;
        RECT 45.280 16.050 45.420 20.150 ;
        RECT 45.220 15.730 45.480 16.050 ;
        RECT 45.740 15.030 45.880 23.550 ;
        RECT 46.660 16.670 46.800 64.830 ;
        RECT 47.060 62.990 47.320 63.310 ;
        RECT 47.120 56.850 47.260 62.990 ;
        RECT 47.580 58.890 47.720 65.710 ;
        RECT 48.500 63.990 48.640 66.390 ;
        RECT 48.960 64.410 49.100 69.110 ;
        RECT 49.820 68.430 50.080 68.750 ;
        RECT 49.360 66.730 49.620 67.050 ;
        RECT 49.420 65.010 49.560 66.730 ;
        RECT 49.360 64.690 49.620 65.010 ;
        RECT 48.960 64.330 49.560 64.410 ;
        RECT 48.900 64.270 49.560 64.330 ;
        RECT 48.900 64.010 49.160 64.270 ;
        RECT 48.440 63.670 48.700 63.990 ;
        RECT 49.420 63.310 49.560 64.270 ;
        RECT 49.360 62.990 49.620 63.310 ;
        RECT 49.880 59.570 50.020 68.430 ;
        RECT 50.280 64.690 50.540 65.010 ;
        RECT 49.820 59.250 50.080 59.570 ;
        RECT 50.340 58.970 50.480 64.690 ;
        RECT 47.520 58.570 47.780 58.890 ;
        RECT 49.880 58.830 50.480 58.970 ;
        RECT 47.060 56.530 47.320 56.850 ;
        RECT 48.440 55.850 48.700 56.170 ;
        RECT 48.500 53.110 48.640 55.850 ;
        RECT 49.360 55.510 49.620 55.830 ;
        RECT 48.440 52.790 48.700 53.110 ;
        RECT 49.420 49.710 49.560 55.510 ;
        RECT 49.880 53.110 50.020 58.830 ;
        RECT 50.280 55.850 50.540 56.170 ;
        RECT 49.820 52.790 50.080 53.110 ;
        RECT 47.520 49.390 47.780 49.710 ;
        RECT 49.360 49.390 49.620 49.710 ;
        RECT 47.580 48.010 47.720 49.390 ;
        RECT 49.420 48.010 49.560 49.390 ;
        RECT 47.520 47.690 47.780 48.010 ;
        RECT 49.360 47.690 49.620 48.010 ;
        RECT 49.420 41.890 49.560 47.690 ;
        RECT 49.880 45.290 50.020 52.790 ;
        RECT 49.820 44.970 50.080 45.290 ;
        RECT 47.980 41.570 48.240 41.890 ;
        RECT 49.360 41.570 49.620 41.890 ;
        RECT 48.040 40.530 48.180 41.570 ;
        RECT 47.980 40.210 48.240 40.530 ;
        RECT 49.820 39.365 50.080 39.510 ;
        RECT 49.810 38.995 50.090 39.365 ;
        RECT 49.880 37.470 50.020 38.995 ;
        RECT 49.820 37.150 50.080 37.470 ;
        RECT 47.060 36.470 47.320 36.790 ;
        RECT 47.520 36.470 47.780 36.790 ;
        RECT 47.980 36.470 48.240 36.790 ;
        RECT 47.120 26.590 47.260 36.470 ;
        RECT 47.580 35.090 47.720 36.470 ;
        RECT 47.520 34.770 47.780 35.090 ;
        RECT 48.040 29.650 48.180 36.470 ;
        RECT 49.820 31.370 50.080 31.690 ;
        RECT 47.980 29.330 48.240 29.650 ;
        RECT 47.060 26.270 47.320 26.590 ;
        RECT 48.040 25.910 48.180 29.330 ;
        RECT 48.900 25.930 49.160 26.250 ;
        RECT 47.980 25.590 48.240 25.910 ;
        RECT 47.060 23.725 47.320 23.870 ;
        RECT 47.050 23.355 47.330 23.725 ;
        RECT 48.040 20.470 48.180 25.590 ;
        RECT 48.960 20.810 49.100 25.930 ;
        RECT 49.880 25.570 50.020 31.370 ;
        RECT 49.820 25.250 50.080 25.570 ;
        RECT 49.880 24.210 50.020 25.250 ;
        RECT 49.820 23.890 50.080 24.210 ;
        RECT 49.360 22.870 49.620 23.190 ;
        RECT 48.900 20.490 49.160 20.810 ;
        RECT 47.980 20.150 48.240 20.470 ;
        RECT 48.440 19.470 48.700 19.790 ;
        RECT 48.500 18.090 48.640 19.470 ;
        RECT 49.420 18.770 49.560 22.870 ;
        RECT 49.360 18.450 49.620 18.770 ;
        RECT 48.440 17.770 48.700 18.090 ;
        RECT 46.660 16.530 48.180 16.670 ;
        RECT 48.040 15.710 48.180 16.530 ;
        RECT 47.980 15.390 48.240 15.710 ;
        RECT 49.420 15.030 49.560 18.450 ;
        RECT 44.300 14.940 44.560 15.030 ;
        RECT 43.900 14.800 44.560 14.940 ;
        RECT 44.300 14.710 44.560 14.800 ;
        RECT 45.680 14.710 45.940 15.030 ;
        RECT 49.360 14.710 49.620 15.030 ;
        RECT 49.880 14.690 50.020 23.890 ;
        RECT 50.340 22.850 50.480 55.850 ;
        RECT 50.800 50.050 50.940 96.990 ;
        RECT 51.260 96.970 51.400 122.830 ;
        RECT 54.020 118.050 54.160 161.430 ;
        RECT 54.480 160.210 54.620 161.590 ;
        RECT 54.940 161.570 55.080 167.710 ;
        RECT 54.940 161.430 56.000 161.570 ;
        RECT 54.880 160.910 55.140 161.230 ;
        RECT 55.340 160.910 55.600 161.230 ;
        RECT 54.420 159.890 54.680 160.210 ;
        RECT 54.480 156.470 54.620 159.890 ;
        RECT 54.940 159.190 55.080 160.910 ;
        RECT 54.880 158.870 55.140 159.190 ;
        RECT 54.940 157.490 55.080 158.870 ;
        RECT 54.880 157.170 55.140 157.490 ;
        RECT 54.420 156.150 54.680 156.470 ;
        RECT 55.400 155.790 55.540 160.910 ;
        RECT 54.420 155.470 54.680 155.790 ;
        RECT 55.340 155.470 55.600 155.790 ;
        RECT 54.480 153.410 54.620 155.470 ;
        RECT 54.880 153.770 55.140 154.090 ;
        RECT 54.420 153.090 54.680 153.410 ;
        RECT 54.940 151.710 55.080 153.770 ;
        RECT 55.860 153.410 56.000 161.430 ;
        RECT 57.240 154.090 57.380 168.050 ;
        RECT 57.700 167.690 57.840 170.090 ;
        RECT 57.640 167.370 57.900 167.690 ;
        RECT 57.700 159.530 57.840 167.370 ;
        RECT 58.160 167.350 58.300 172.810 ;
        RECT 59.080 172.700 59.220 177.570 ;
        RECT 60.000 173.810 60.140 177.570 ;
        RECT 59.940 173.490 60.200 173.810 ;
        RECT 59.940 172.700 60.200 172.790 ;
        RECT 59.080 172.560 60.200 172.700 ;
        RECT 59.940 172.470 60.200 172.560 ;
        RECT 58.560 170.430 58.820 170.750 ;
        RECT 58.620 167.690 58.760 170.430 ;
        RECT 60.000 169.730 60.140 172.470 ;
        RECT 59.940 169.410 60.200 169.730 ;
        RECT 60.460 169.390 60.600 177.910 ;
        RECT 61.840 177.830 62.440 177.970 ;
        RECT 61.320 175.870 61.580 176.190 ;
        RECT 60.400 169.070 60.660 169.390 ;
        RECT 60.860 169.070 61.120 169.390 ;
        RECT 58.560 167.370 58.820 167.690 ;
        RECT 58.100 167.030 58.360 167.350 ;
        RECT 58.160 165.310 58.300 167.030 ;
        RECT 58.100 164.990 58.360 165.310 ;
        RECT 58.620 164.970 58.760 167.370 ;
        RECT 60.920 167.350 61.060 169.070 ;
        RECT 60.860 167.030 61.120 167.350 ;
        RECT 59.020 166.690 59.280 167.010 ;
        RECT 59.080 164.970 59.220 166.690 ;
        RECT 61.380 166.410 61.520 175.870 ;
        RECT 61.840 171.090 61.980 177.830 ;
        RECT 63.680 176.530 63.820 180.720 ;
        RECT 64.600 180.610 64.740 183.010 ;
        RECT 65.520 181.970 65.660 183.350 ;
        RECT 65.460 181.650 65.720 181.970 ;
        RECT 65.000 181.310 65.260 181.630 ;
        RECT 64.540 180.290 64.800 180.610 ;
        RECT 65.060 180.010 65.200 181.310 ;
        RECT 64.600 179.870 65.200 180.010 ;
        RECT 64.600 178.230 64.740 179.870 ;
        RECT 65.520 178.230 65.660 181.650 ;
        RECT 68.280 181.290 68.420 184.030 ;
        RECT 68.740 181.630 68.880 184.370 ;
        RECT 69.200 182.990 69.340 192.530 ;
        RECT 69.660 192.170 69.800 193.550 ;
        RECT 71.040 192.510 71.180 198.990 ;
        RECT 101.480 198.895 105.480 198.965 ;
        RECT 112.175 198.905 112.545 200.445 ;
        RECT 117.615 198.905 117.985 200.445 ;
        RECT 123.055 198.905 123.425 200.445 ;
        RECT 128.495 198.905 128.865 200.445 ;
        RECT 130.390 200.275 130.710 200.335 ;
        RECT 133.030 200.275 133.170 200.595 ;
        RECT 137.190 200.535 137.510 200.595 ;
        RECT 141.610 200.735 141.930 200.795 ;
        RECT 146.710 200.735 147.030 200.795 ;
        RECT 141.610 200.595 147.030 200.735 ;
        RECT 141.610 200.535 141.930 200.595 ;
        RECT 146.710 200.535 147.030 200.595 ;
        RECT 130.390 200.135 133.170 200.275 ;
        RECT 130.390 200.075 130.710 200.135 ;
        RECT 133.935 198.905 134.305 200.445 ;
        RECT 139.375 198.905 139.745 200.445 ;
        RECT 140.590 200.275 140.910 200.335 ;
        RECT 143.310 200.275 143.630 200.335 ;
        RECT 140.590 200.135 143.630 200.275 ;
        RECT 140.590 200.075 140.910 200.135 ;
        RECT 143.310 200.075 143.630 200.135 ;
        RECT 144.815 198.905 145.185 200.445 ;
        RECT 147.050 198.895 147.370 198.955 ;
        RECT 148.660 198.895 148.920 198.985 ;
        RECT 155.245 198.895 159.245 198.965 ;
        RECT 101.480 198.755 107.330 198.895 ;
        RECT 101.480 198.685 105.480 198.755 ;
        RECT 107.190 198.435 107.330 198.755 ;
        RECT 147.050 198.755 159.245 198.895 ;
        RECT 147.050 198.695 147.370 198.755 ;
        RECT 148.660 198.665 148.920 198.755 ;
        RECT 155.245 198.685 159.245 198.755 ;
        RECT 111.410 198.435 111.740 198.530 ;
        RECT 112.710 198.435 113.030 198.495 ;
        RECT 107.190 198.295 113.030 198.435 ;
        RECT 111.410 198.200 111.740 198.295 ;
        RECT 112.710 198.235 113.030 198.295 ;
        RECT 126.990 198.435 127.310 198.495 ;
        RECT 134.470 198.435 134.790 198.495 ;
        RECT 136.170 198.435 136.490 198.495 ;
        RECT 140.590 198.435 140.910 198.495 ;
        RECT 126.990 198.295 135.890 198.435 ;
        RECT 126.990 198.235 127.310 198.295 ;
        RECT 134.470 198.235 134.790 198.295 ;
        RECT 114.410 197.975 114.730 198.035 ;
        RECT 123.590 197.975 123.910 198.035 ;
        RECT 126.990 197.975 127.310 198.035 ;
        RECT 114.410 197.835 127.310 197.975 ;
        RECT 114.410 197.775 114.730 197.835 ;
        RECT 123.590 197.775 123.910 197.835 ;
        RECT 126.990 197.775 127.310 197.835 ;
        RECT 133.450 197.975 133.770 198.035 ;
        RECT 134.810 197.975 135.130 198.035 ;
        RECT 133.450 197.835 135.130 197.975 ;
        RECT 135.750 197.975 135.890 198.295 ;
        RECT 136.170 198.295 140.910 198.435 ;
        RECT 136.170 198.235 136.490 198.295 ;
        RECT 140.590 198.235 140.910 198.295 ;
        RECT 144.330 198.435 144.650 198.495 ;
        RECT 146.030 198.435 146.350 198.495 ;
        RECT 144.330 198.295 146.350 198.435 ;
        RECT 144.330 198.235 144.650 198.295 ;
        RECT 146.030 198.235 146.350 198.295 ;
        RECT 140.590 197.975 140.910 198.035 ;
        RECT 135.750 197.835 140.910 197.975 ;
        RECT 133.450 197.775 133.770 197.835 ;
        RECT 134.810 197.775 135.130 197.835 ;
        RECT 140.590 197.775 140.910 197.835 ;
        RECT 143.990 197.975 144.310 198.035 ;
        RECT 145.350 197.975 145.670 198.035 ;
        RECT 143.990 197.835 145.670 197.975 ;
        RECT 143.990 197.775 144.310 197.835 ;
        RECT 145.350 197.775 145.670 197.835 ;
        RECT 71.440 197.290 71.700 197.610 ;
        RECT 124.610 197.515 124.930 197.575 ;
        RECT 124.610 197.315 125.010 197.515 ;
        RECT 128.010 197.315 128.330 197.575 ;
        RECT 135.150 197.515 135.470 197.575 ;
        RECT 137.870 197.515 138.190 197.575 ;
        RECT 135.150 197.375 138.190 197.515 ;
        RECT 135.150 197.315 135.470 197.375 ;
        RECT 137.870 197.315 138.190 197.375 ;
        RECT 140.930 197.515 141.250 197.575 ;
        RECT 142.630 197.515 142.950 197.575 ;
        RECT 140.930 197.375 142.950 197.515 ;
        RECT 140.930 197.315 141.250 197.375 ;
        RECT 142.630 197.315 142.950 197.375 ;
        RECT 71.500 195.570 71.640 197.290 ;
        RECT 77.420 196.950 77.680 197.270 ;
        RECT 124.870 197.055 125.010 197.315 ;
        RECT 128.100 197.055 128.240 197.315 ;
        RECT 130.050 197.055 130.370 197.115 ;
        RECT 135.830 197.055 136.150 197.115 ;
        RECT 71.440 195.250 71.700 195.570 ;
        RECT 77.480 194.890 77.620 196.950 ;
        RECT 124.870 196.915 136.150 197.055 ;
        RECT 130.050 196.855 130.370 196.915 ;
        RECT 135.830 196.855 136.150 196.915 ;
        RECT 140.590 197.055 140.910 197.115 ;
        RECT 143.650 197.055 143.970 197.115 ;
        RECT 140.590 196.915 143.970 197.055 ;
        RECT 140.590 196.855 140.910 196.915 ;
        RECT 143.650 196.855 143.970 196.915 ;
        RECT 124.950 196.595 125.270 196.655 ;
        RECT 134.810 196.595 135.130 196.655 ;
        RECT 124.950 196.455 135.130 196.595 ;
        RECT 124.950 196.395 125.270 196.455 ;
        RECT 134.810 196.395 135.130 196.455 ;
        RECT 117.130 196.135 117.450 196.195 ;
        RECT 122.230 196.135 122.550 196.195 ;
        RECT 126.650 196.135 126.970 196.195 ;
        RECT 117.130 195.995 126.970 196.135 ;
        RECT 117.130 195.935 117.450 195.995 ;
        RECT 122.230 195.935 122.550 195.995 ;
        RECT 126.650 195.935 126.970 195.995 ;
        RECT 130.390 196.135 130.710 196.195 ;
        RECT 131.750 196.135 132.070 196.195 ;
        RECT 138.550 196.135 138.870 196.195 ;
        RECT 143.310 196.135 143.630 196.195 ;
        RECT 130.390 195.995 143.630 196.135 ;
        RECT 130.390 195.935 130.710 195.995 ;
        RECT 131.750 195.935 132.070 195.995 ;
        RECT 138.550 195.935 138.870 195.995 ;
        RECT 143.310 195.935 143.630 195.995 ;
        RECT 133.450 195.675 133.770 195.735 ;
        RECT 137.530 195.675 137.850 195.735 ;
        RECT 140.250 195.675 140.570 195.735 ;
        RECT 141.610 195.675 141.930 195.735 ;
        RECT 143.650 195.675 143.970 195.735 ;
        RECT 133.450 195.535 140.570 195.675 ;
        RECT 133.450 195.475 133.770 195.535 ;
        RECT 137.530 195.475 137.850 195.535 ;
        RECT 140.250 195.475 140.570 195.535 ;
        RECT 141.190 195.535 143.970 195.675 ;
        RECT 116.110 195.215 116.430 195.275 ;
        RECT 121.890 195.215 122.210 195.275 ;
        RECT 125.290 195.215 125.610 195.275 ;
        RECT 141.190 195.215 141.330 195.535 ;
        RECT 141.610 195.475 141.930 195.535 ;
        RECT 143.650 195.475 143.970 195.535 ;
        RECT 146.030 195.675 146.350 195.735 ;
        RECT 148.050 195.675 148.470 195.800 ;
        RECT 155.245 195.675 159.245 195.745 ;
        RECT 146.030 195.535 159.245 195.675 ;
        RECT 146.030 195.475 146.350 195.535 ;
        RECT 148.050 195.410 148.470 195.535 ;
        RECT 155.245 195.465 159.245 195.535 ;
        RECT 116.110 195.075 141.330 195.215 ;
        RECT 116.110 195.015 116.430 195.075 ;
        RECT 121.890 195.015 122.210 195.075 ;
        RECT 125.290 195.015 125.610 195.075 ;
        RECT 77.420 194.570 77.680 194.890 ;
        RECT 113.390 194.755 113.710 194.815 ;
        RECT 114.070 194.755 114.390 194.815 ;
        RECT 116.110 194.755 116.430 194.815 ;
        RECT 113.390 194.615 116.430 194.755 ;
        RECT 73.280 193.890 73.540 194.210 ;
        RECT 73.340 192.850 73.480 193.890 ;
        RECT 73.280 192.530 73.540 192.850 ;
        RECT 70.980 192.190 71.240 192.510 ;
        RECT 69.600 191.850 69.860 192.170 ;
        RECT 71.900 191.850 72.160 192.170 ;
        RECT 74.660 191.850 74.920 192.170 ;
        RECT 69.660 189.450 69.800 191.850 ;
        RECT 70.980 191.510 71.240 191.830 ;
        RECT 69.600 189.130 69.860 189.450 ;
        RECT 71.040 189.110 71.180 191.510 ;
        RECT 71.960 190.130 72.100 191.850 ;
        RECT 71.900 189.810 72.160 190.130 ;
        RECT 74.720 189.110 74.860 191.850 ;
        RECT 70.980 188.790 71.240 189.110 ;
        RECT 74.660 188.790 74.920 189.110 ;
        RECT 72.820 188.450 73.080 188.770 ;
        RECT 71.900 183.010 72.160 183.330 ;
        RECT 69.140 182.670 69.400 182.990 ;
        RECT 70.060 182.670 70.320 182.990 ;
        RECT 68.680 181.310 68.940 181.630 ;
        RECT 68.220 180.970 68.480 181.290 ;
        RECT 64.540 177.910 64.800 178.230 ;
        RECT 65.460 177.910 65.720 178.230 ;
        RECT 65.920 177.910 66.180 178.230 ;
        RECT 63.620 176.210 63.880 176.530 ;
        RECT 63.680 172.790 63.820 176.210 ;
        RECT 64.600 176.190 64.740 177.910 ;
        RECT 64.540 175.870 64.800 176.190 ;
        RECT 63.620 172.470 63.880 172.790 ;
        RECT 64.080 172.470 64.340 172.790 ;
        RECT 61.780 170.770 62.040 171.090 ;
        RECT 61.840 170.410 61.980 170.770 ;
        RECT 61.780 170.090 62.040 170.410 ;
        RECT 61.840 169.390 61.980 170.090 ;
        RECT 61.780 169.070 62.040 169.390 ;
        RECT 63.680 168.280 63.820 172.470 ;
        RECT 64.140 170.070 64.280 172.470 ;
        RECT 65.980 171.090 66.120 177.910 ;
        RECT 68.280 177.890 68.420 180.970 ;
        RECT 69.200 180.270 69.340 182.670 ;
        RECT 69.600 181.310 69.860 181.630 ;
        RECT 70.120 181.540 70.260 182.670 ;
        RECT 70.520 181.540 70.780 181.630 ;
        RECT 70.120 181.400 70.780 181.540 ;
        RECT 70.520 181.310 70.780 181.400 ;
        RECT 69.140 179.950 69.400 180.270 ;
        RECT 69.200 178.570 69.340 179.950 ;
        RECT 69.660 179.250 69.800 181.310 ;
        RECT 70.060 180.630 70.320 180.950 ;
        RECT 70.980 180.630 71.240 180.950 ;
        RECT 69.600 178.930 69.860 179.250 ;
        RECT 69.140 178.250 69.400 178.570 ;
        RECT 68.220 177.570 68.480 177.890 ;
        RECT 68.280 172.110 68.420 177.570 ;
        RECT 70.120 177.550 70.260 180.630 ;
        RECT 70.060 177.230 70.320 177.550 ;
        RECT 69.140 175.530 69.400 175.850 ;
        RECT 69.200 172.790 69.340 175.530 ;
        RECT 70.120 175.510 70.260 177.230 ;
        RECT 70.520 175.530 70.780 175.850 ;
        RECT 70.060 175.190 70.320 175.510 ;
        RECT 69.600 174.510 69.860 174.830 ;
        RECT 69.140 172.470 69.400 172.790 ;
        RECT 68.220 171.790 68.480 172.110 ;
        RECT 65.920 170.770 66.180 171.090 ;
        RECT 66.380 170.770 66.640 171.090 ;
        RECT 64.080 169.750 64.340 170.070 ;
        RECT 63.680 168.140 64.280 168.280 ;
        RECT 62.240 167.370 62.500 167.690 ;
        RECT 63.620 167.370 63.880 167.690 ;
        RECT 60.460 166.270 61.520 166.410 ;
        RECT 60.460 165.650 60.600 166.270 ;
        RECT 60.400 165.330 60.660 165.650 ;
        RECT 58.560 164.650 58.820 164.970 ;
        RECT 59.020 164.650 59.280 164.970 ;
        RECT 59.080 161.910 59.220 164.650 ;
        RECT 59.020 161.590 59.280 161.910 ;
        RECT 57.640 159.210 57.900 159.530 ;
        RECT 59.080 156.890 59.220 161.590 ;
        RECT 59.080 156.750 59.680 156.890 ;
        RECT 57.640 156.150 57.900 156.470 ;
        RECT 59.020 156.150 59.280 156.470 ;
        RECT 57.700 154.770 57.840 156.150 ;
        RECT 57.640 154.450 57.900 154.770 ;
        RECT 57.180 153.770 57.440 154.090 ;
        RECT 55.800 153.090 56.060 153.410 ;
        RECT 55.340 152.750 55.600 153.070 ;
        RECT 54.880 151.390 55.140 151.710 ;
        RECT 54.940 149.330 55.080 151.390 ;
        RECT 55.400 151.030 55.540 152.750 ;
        RECT 55.340 150.710 55.600 151.030 ;
        RECT 59.080 150.690 59.220 156.150 ;
        RECT 59.020 150.370 59.280 150.690 ;
        RECT 54.880 149.010 55.140 149.330 ;
        RECT 59.020 148.330 59.280 148.650 ;
        RECT 59.080 146.610 59.220 148.330 ;
        RECT 59.020 146.290 59.280 146.610 ;
        RECT 59.540 143.550 59.680 156.750 ;
        RECT 59.940 151.730 60.200 152.050 ;
        RECT 60.000 151.370 60.140 151.730 ;
        RECT 59.940 151.050 60.200 151.370 ;
        RECT 59.480 143.230 59.740 143.550 ;
        RECT 60.000 143.210 60.140 151.050 ;
        RECT 60.460 145.590 60.600 165.330 ;
        RECT 62.300 159.870 62.440 167.370 ;
        RECT 63.680 164.970 63.820 167.370 ;
        RECT 64.140 164.970 64.280 168.140 ;
        RECT 66.440 165.650 66.580 170.770 ;
        RECT 67.760 170.320 68.020 170.410 ;
        RECT 68.280 170.320 68.420 171.790 ;
        RECT 69.200 170.410 69.340 172.470 ;
        RECT 69.660 172.450 69.800 174.510 ;
        RECT 70.580 173.810 70.720 175.530 ;
        RECT 70.520 173.490 70.780 173.810 ;
        RECT 70.050 172.955 70.330 173.325 ;
        RECT 70.060 172.810 70.320 172.955 ;
        RECT 69.600 172.130 69.860 172.450 ;
        RECT 71.040 170.750 71.180 180.630 ;
        RECT 71.960 180.270 72.100 183.010 ;
        RECT 71.900 179.950 72.160 180.270 ;
        RECT 72.880 178.230 73.020 188.450 ;
        RECT 77.480 184.010 77.620 194.570 ;
        RECT 113.390 194.555 113.710 194.615 ;
        RECT 114.070 194.555 114.390 194.615 ;
        RECT 116.110 194.555 116.430 194.615 ;
        RECT 140.590 194.755 140.910 194.815 ;
        RECT 142.630 194.755 142.950 194.815 ;
        RECT 140.590 194.615 142.950 194.755 ;
        RECT 140.590 194.555 140.910 194.615 ;
        RECT 142.630 194.555 142.950 194.615 ;
        RECT 120.870 194.295 121.190 194.355 ;
        RECT 121.550 194.295 121.870 194.355 ;
        RECT 129.030 194.295 129.350 194.355 ;
        RECT 120.870 194.155 129.350 194.295 ;
        RECT 120.870 194.095 121.190 194.155 ;
        RECT 121.550 194.095 121.870 194.155 ;
        RECT 129.030 194.095 129.350 194.155 ;
        RECT 115.235 193.835 115.605 193.905 ;
        RECT 118.830 193.835 119.150 193.895 ;
        RECT 115.235 193.695 119.150 193.835 ;
        RECT 115.235 193.625 115.605 193.695 ;
        RECT 118.830 193.635 119.150 193.695 ;
        RECT 127.330 193.835 127.650 193.895 ;
        RECT 130.730 193.835 131.050 193.895 ;
        RECT 137.190 193.835 137.510 193.895 ;
        RECT 127.330 193.695 137.510 193.835 ;
        RECT 127.330 193.635 127.650 193.695 ;
        RECT 130.730 193.635 131.050 193.695 ;
        RECT 137.190 193.635 137.510 193.695 ;
        RECT 143.650 193.835 143.970 193.895 ;
        RECT 146.710 193.835 147.030 193.895 ;
        RECT 143.650 193.695 147.030 193.835 ;
        RECT 143.650 193.635 143.970 193.695 ;
        RECT 146.710 193.635 147.030 193.695 ;
        RECT 132.770 192.915 133.090 192.975 ;
        RECT 134.470 192.915 134.790 192.975 ;
        RECT 132.770 192.775 134.790 192.915 ;
        RECT 132.770 192.715 133.090 192.775 ;
        RECT 134.470 192.715 134.790 192.775 ;
        RECT 101.480 192.455 105.480 192.525 ;
        RECT 109.920 192.455 110.240 192.515 ;
        RECT 112.710 192.455 113.030 192.515 ;
        RECT 101.480 192.315 113.030 192.455 ;
        RECT 101.480 192.245 105.480 192.315 ;
        RECT 109.920 192.255 110.240 192.315 ;
        RECT 112.710 192.255 113.030 192.315 ;
        RECT 118.830 192.455 119.150 192.515 ;
        RECT 125.435 192.455 125.805 192.525 ;
        RECT 118.830 192.315 125.805 192.455 ;
        RECT 118.830 192.255 119.150 192.315 ;
        RECT 125.435 192.245 125.805 192.315 ;
        RECT 147.050 192.455 147.370 192.515 ;
        RECT 148.570 192.455 148.900 192.550 ;
        RECT 155.245 192.455 159.245 192.525 ;
        RECT 147.050 192.315 159.245 192.455 ;
        RECT 147.050 192.255 147.370 192.315 ;
        RECT 148.570 192.220 148.900 192.315 ;
        RECT 155.245 192.245 159.245 192.315 ;
        RECT 113.390 191.995 113.710 192.055 ;
        RECT 120.870 191.995 121.190 192.055 ;
        RECT 124.270 191.995 124.590 192.055 ;
        RECT 113.390 191.855 124.590 191.995 ;
        RECT 113.390 191.795 113.710 191.855 ;
        RECT 120.870 191.795 121.190 191.855 ;
        RECT 124.270 191.795 124.590 191.855 ;
        RECT 132.770 191.995 133.090 192.055 ;
        RECT 138.210 191.995 138.530 192.055 ;
        RECT 145.350 191.995 145.670 192.055 ;
        RECT 132.770 191.855 145.670 191.995 ;
        RECT 132.770 191.795 133.090 191.855 ;
        RECT 138.210 191.795 138.530 191.855 ;
        RECT 145.350 191.795 145.670 191.855 ;
        RECT 127.330 191.535 127.650 191.595 ;
        RECT 129.030 191.535 129.350 191.595 ;
        RECT 127.330 191.395 129.350 191.535 ;
        RECT 127.330 191.335 127.650 191.395 ;
        RECT 129.030 191.335 129.350 191.395 ;
        RECT 138.550 191.535 138.870 191.595 ;
        RECT 138.550 191.395 143.880 191.535 ;
        RECT 138.550 191.335 138.870 191.395 ;
        RECT 143.740 191.145 143.880 191.395 ;
        RECT 118.635 191.135 119.005 191.145 ;
        RECT 143.740 191.135 144.165 191.145 ;
        RECT 118.635 190.875 119.150 191.135 ;
        RECT 122.570 191.075 122.890 191.135 ;
        RECT 123.590 191.075 123.910 191.135 ;
        RECT 122.570 190.935 123.910 191.075 ;
        RECT 122.570 190.875 122.890 190.935 ;
        RECT 123.590 190.875 123.910 190.935 ;
        RECT 129.710 191.075 130.030 191.135 ;
        RECT 135.150 191.075 135.470 191.135 ;
        RECT 137.530 191.075 137.850 191.135 ;
        RECT 138.550 191.075 138.870 191.135 ;
        RECT 129.710 190.935 130.450 191.075 ;
        RECT 129.710 190.875 130.030 190.935 ;
        RECT 118.635 190.865 119.005 190.875 ;
        RECT 128.835 190.155 129.205 190.225 ;
        RECT 129.710 190.155 130.030 190.215 ;
        RECT 128.835 190.015 130.030 190.155 ;
        RECT 130.310 190.155 130.450 190.935 ;
        RECT 135.150 190.935 138.870 191.075 ;
        RECT 135.150 190.875 135.470 190.935 ;
        RECT 137.530 190.875 137.850 190.935 ;
        RECT 138.550 190.875 138.870 190.935 ;
        RECT 143.650 190.875 144.165 191.135 ;
        RECT 143.795 190.865 144.165 190.875 ;
        RECT 141.610 190.615 141.930 190.675 ;
        RECT 142.970 190.615 143.290 190.675 ;
        RECT 146.030 190.615 146.350 190.675 ;
        RECT 141.610 190.475 146.350 190.615 ;
        RECT 141.610 190.415 141.930 190.475 ;
        RECT 142.970 190.415 143.290 190.475 ;
        RECT 146.030 190.415 146.350 190.475 ;
        RECT 135.830 190.155 136.150 190.215 ;
        RECT 130.310 190.015 136.150 190.155 ;
        RECT 128.835 189.945 129.205 190.015 ;
        RECT 129.710 189.955 130.030 190.015 ;
        RECT 135.830 189.955 136.150 190.015 ;
        RECT 113.730 189.695 114.050 189.755 ;
        RECT 116.110 189.695 116.430 189.755 ;
        RECT 118.150 189.695 118.470 189.755 ;
        RECT 113.730 189.555 118.470 189.695 ;
        RECT 113.730 189.495 114.050 189.555 ;
        RECT 116.110 189.495 116.430 189.555 ;
        RECT 118.150 189.495 118.470 189.555 ;
        RECT 124.610 189.695 124.930 189.755 ;
        RECT 127.670 189.695 127.990 189.755 ;
        RECT 129.370 189.695 129.690 189.755 ;
        RECT 131.750 189.695 132.070 189.755 ;
        RECT 124.610 189.555 132.070 189.695 ;
        RECT 124.610 189.495 124.930 189.555 ;
        RECT 127.670 189.495 127.990 189.555 ;
        RECT 129.370 189.495 129.690 189.555 ;
        RECT 131.750 189.495 132.070 189.555 ;
        RECT 111.835 189.235 112.205 189.305 ;
        RECT 113.390 189.235 113.710 189.295 ;
        RECT 111.835 189.095 113.710 189.235 ;
        RECT 111.835 189.025 112.205 189.095 ;
        RECT 113.390 189.035 113.710 189.095 ;
        RECT 116.450 189.235 116.770 189.295 ;
        RECT 118.150 189.235 118.470 189.295 ;
        RECT 116.450 189.095 118.470 189.235 ;
        RECT 116.450 189.035 116.770 189.095 ;
        RECT 118.150 189.035 118.470 189.095 ;
        RECT 119.850 189.235 120.170 189.295 ;
        RECT 121.550 189.235 121.870 189.295 ;
        RECT 124.270 189.235 124.590 189.295 ;
        RECT 119.850 189.095 124.590 189.235 ;
        RECT 119.850 189.035 120.170 189.095 ;
        RECT 121.550 189.035 121.870 189.095 ;
        RECT 124.270 189.035 124.590 189.095 ;
        RECT 125.290 189.235 125.610 189.295 ;
        RECT 135.490 189.235 135.810 189.295 ;
        RECT 125.290 189.095 135.810 189.235 ;
        RECT 125.290 189.035 125.610 189.095 ;
        RECT 135.490 189.035 135.810 189.095 ;
        RECT 122.035 188.835 122.405 188.845 ;
        RECT 114.070 188.775 114.390 188.835 ;
        RECT 119.510 188.775 119.830 188.835 ;
        RECT 114.070 188.635 119.830 188.775 ;
        RECT 114.070 188.575 114.390 188.635 ;
        RECT 119.510 188.575 119.830 188.635 ;
        RECT 121.890 188.575 122.405 188.835 ;
        RECT 140.590 188.775 140.910 188.835 ;
        RECT 142.630 188.775 142.950 188.835 ;
        RECT 140.590 188.635 142.950 188.775 ;
        RECT 140.590 188.575 140.910 188.635 ;
        RECT 142.630 188.575 142.950 188.635 ;
        RECT 122.035 188.565 122.405 188.575 ;
        RECT 114.410 188.315 114.730 188.375 ;
        RECT 118.830 188.315 119.150 188.375 ;
        RECT 120.870 188.315 121.190 188.375 ;
        RECT 127.330 188.315 127.650 188.375 ;
        RECT 114.410 188.175 127.650 188.315 ;
        RECT 114.410 188.115 114.730 188.175 ;
        RECT 118.830 188.115 119.150 188.175 ;
        RECT 120.870 188.115 121.190 188.175 ;
        RECT 127.330 188.115 127.650 188.175 ;
        RECT 135.150 188.315 135.470 188.375 ;
        RECT 138.210 188.315 138.530 188.375 ;
        RECT 138.890 188.315 139.210 188.375 ;
        RECT 145.350 188.315 145.670 188.375 ;
        RECT 135.150 188.175 145.670 188.315 ;
        RECT 135.150 188.115 135.470 188.175 ;
        RECT 138.210 188.115 138.530 188.175 ;
        RECT 138.890 188.115 139.210 188.175 ;
        RECT 145.350 188.115 145.670 188.175 ;
        RECT 119.850 187.855 120.170 187.915 ;
        RECT 127.330 187.855 127.650 187.915 ;
        RECT 119.850 187.715 127.650 187.855 ;
        RECT 119.850 187.655 120.170 187.715 ;
        RECT 127.330 187.655 127.650 187.715 ;
        RECT 128.010 187.855 128.330 187.915 ;
        RECT 129.710 187.855 130.030 187.915 ;
        RECT 128.010 187.715 130.030 187.855 ;
        RECT 128.010 187.655 128.330 187.715 ;
        RECT 129.710 187.655 130.030 187.715 ;
        RECT 130.390 187.855 130.710 187.915 ;
        RECT 135.150 187.855 135.470 187.915 ;
        RECT 141.610 187.855 141.930 187.915 ;
        RECT 143.650 187.855 143.970 187.915 ;
        RECT 130.390 187.715 141.330 187.855 ;
        RECT 130.390 187.655 130.710 187.715 ;
        RECT 135.150 187.655 135.470 187.715 ;
        RECT 118.830 187.395 119.150 187.455 ;
        RECT 121.890 187.395 122.210 187.455 ;
        RECT 118.830 187.255 122.210 187.395 ;
        RECT 118.830 187.195 119.150 187.255 ;
        RECT 121.890 187.195 122.210 187.255 ;
        RECT 122.570 187.395 122.890 187.455 ;
        RECT 126.990 187.395 127.310 187.455 ;
        RECT 122.570 187.255 127.310 187.395 ;
        RECT 122.570 187.195 122.890 187.255 ;
        RECT 126.990 187.195 127.310 187.255 ;
        RECT 129.710 187.395 130.030 187.455 ;
        RECT 132.770 187.395 133.090 187.455 ;
        RECT 129.710 187.255 133.090 187.395 ;
        RECT 129.710 187.195 130.030 187.255 ;
        RECT 132.770 187.195 133.090 187.255 ;
        RECT 135.635 187.395 136.005 187.465 ;
        RECT 140.590 187.395 140.910 187.455 ;
        RECT 135.635 187.255 140.910 187.395 ;
        RECT 141.190 187.395 141.330 187.715 ;
        RECT 141.610 187.715 143.970 187.855 ;
        RECT 141.610 187.655 141.930 187.715 ;
        RECT 143.650 187.655 143.970 187.715 ;
        RECT 146.030 187.855 146.350 187.915 ;
        RECT 149.235 187.855 149.605 187.925 ;
        RECT 146.030 187.715 149.605 187.855 ;
        RECT 146.030 187.655 146.350 187.715 ;
        RECT 149.235 187.645 149.605 187.715 ;
        RECT 142.970 187.395 143.290 187.455 ;
        RECT 141.190 187.255 143.290 187.395 ;
        RECT 135.635 187.185 136.005 187.255 ;
        RECT 140.590 187.195 140.910 187.255 ;
        RECT 142.970 187.195 143.290 187.255 ;
        RECT 122.230 186.935 122.550 186.995 ;
        RECT 124.270 186.935 124.590 186.995 ;
        RECT 129.370 186.935 129.690 186.995 ;
        RECT 122.230 186.795 129.690 186.935 ;
        RECT 122.230 186.735 122.550 186.795 ;
        RECT 124.270 186.735 124.590 186.795 ;
        RECT 129.370 186.735 129.690 186.795 ;
        RECT 136.170 186.935 136.490 186.995 ;
        RECT 138.210 186.935 138.530 186.995 ;
        RECT 136.170 186.795 138.530 186.935 ;
        RECT 136.170 186.735 136.490 186.795 ;
        RECT 138.210 186.735 138.530 186.795 ;
        RECT 145.835 186.535 146.205 186.545 ;
        RECT 117.130 186.475 117.450 186.535 ;
        RECT 124.270 186.475 124.590 186.535 ;
        RECT 117.130 186.335 124.590 186.475 ;
        RECT 117.130 186.275 117.450 186.335 ;
        RECT 124.270 186.275 124.590 186.335 ;
        RECT 130.730 186.475 131.050 186.535 ;
        RECT 135.150 186.475 135.470 186.535 ;
        RECT 139.910 186.475 140.230 186.535 ;
        RECT 130.730 186.335 135.470 186.475 ;
        RECT 130.730 186.275 131.050 186.335 ;
        RECT 135.150 186.275 135.470 186.335 ;
        RECT 135.750 186.335 140.230 186.475 ;
        RECT 114.410 186.015 114.730 186.075 ;
        RECT 118.830 186.015 119.150 186.075 ;
        RECT 114.410 185.875 119.150 186.015 ;
        RECT 114.410 185.815 114.730 185.875 ;
        RECT 118.830 185.815 119.150 185.875 ;
        RECT 121.550 186.015 121.870 186.075 ;
        RECT 127.330 186.015 127.650 186.075 ;
        RECT 121.550 185.875 127.650 186.015 ;
        RECT 121.550 185.815 121.870 185.875 ;
        RECT 127.330 185.815 127.650 185.875 ;
        RECT 132.770 186.015 133.090 186.075 ;
        RECT 135.150 186.015 135.470 186.075 ;
        RECT 135.750 186.015 135.890 186.335 ;
        RECT 139.910 186.275 140.230 186.335 ;
        RECT 145.835 186.275 146.350 186.535 ;
        RECT 145.835 186.265 146.205 186.275 ;
        RECT 132.770 185.875 135.890 186.015 ;
        RECT 138.890 186.015 139.210 186.075 ;
        RECT 139.910 186.015 140.230 186.075 ;
        RECT 138.890 185.875 140.230 186.015 ;
        RECT 132.770 185.815 133.090 185.875 ;
        RECT 135.150 185.815 135.470 185.875 ;
        RECT 138.890 185.815 139.210 185.875 ;
        RECT 139.910 185.815 140.230 185.875 ;
        RECT 108.435 185.555 108.805 185.625 ;
        RECT 119.170 185.555 119.490 185.615 ;
        RECT 108.435 185.415 119.490 185.555 ;
        RECT 108.435 185.345 108.805 185.415 ;
        RECT 119.170 185.355 119.490 185.415 ;
        RECT 135.830 185.555 136.150 185.615 ;
        RECT 138.210 185.555 138.530 185.615 ;
        RECT 145.350 185.555 145.670 185.615 ;
        RECT 135.830 185.415 145.670 185.555 ;
        RECT 135.830 185.355 136.150 185.415 ;
        RECT 138.210 185.355 138.530 185.415 ;
        RECT 145.350 185.355 145.670 185.415 ;
        RECT 116.110 185.095 116.430 185.155 ;
        RECT 118.830 185.095 119.150 185.155 ;
        RECT 121.210 185.095 121.530 185.155 ;
        RECT 116.110 184.955 121.530 185.095 ;
        RECT 116.110 184.895 116.430 184.955 ;
        RECT 118.830 184.895 119.150 184.955 ;
        RECT 121.210 184.895 121.530 184.955 ;
        RECT 132.235 185.095 132.605 185.165 ;
        RECT 132.770 185.095 133.090 185.155 ;
        RECT 132.235 184.955 133.090 185.095 ;
        RECT 132.235 184.885 132.605 184.955 ;
        RECT 132.770 184.895 133.090 184.955 ;
        RECT 139.035 185.095 139.405 185.165 ;
        RECT 140.590 185.095 140.910 185.155 ;
        RECT 139.035 184.955 140.910 185.095 ;
        RECT 139.035 184.885 139.405 184.955 ;
        RECT 140.590 184.895 140.910 184.955 ;
        RECT 142.435 185.095 142.805 185.165 ;
        RECT 143.650 185.095 143.970 185.155 ;
        RECT 142.435 184.955 143.970 185.095 ;
        RECT 142.435 184.885 142.805 184.955 ;
        RECT 143.650 184.895 143.970 184.955 ;
        RECT 146.030 185.095 146.350 185.155 ;
        RECT 152.635 185.095 153.005 185.165 ;
        RECT 146.030 184.955 153.005 185.095 ;
        RECT 146.030 184.895 146.350 184.955 ;
        RECT 152.635 184.885 153.005 184.955 ;
        RECT 77.420 183.690 77.680 184.010 ;
        RECT 73.280 183.350 73.540 183.670 ;
        RECT 73.340 181.970 73.480 183.350 ;
        RECT 73.280 181.650 73.540 181.970 ;
        RECT 72.820 177.910 73.080 178.230 ;
        RECT 71.440 177.230 71.700 177.550 ;
        RECT 71.500 175.850 71.640 177.230 ;
        RECT 71.440 175.530 71.700 175.850 ;
        RECT 71.900 175.530 72.160 175.850 ;
        RECT 71.960 175.170 72.100 175.530 ;
        RECT 72.360 175.190 72.620 175.510 ;
        RECT 71.900 174.850 72.160 175.170 ;
        RECT 71.440 174.510 71.700 174.830 ;
        RECT 71.500 173.470 71.640 174.510 ;
        RECT 71.440 173.150 71.700 173.470 ;
        RECT 71.960 172.790 72.100 174.850 ;
        RECT 71.900 172.470 72.160 172.790 ;
        RECT 70.980 170.430 71.240 170.750 ;
        RECT 67.760 170.180 68.420 170.320 ;
        RECT 67.760 170.090 68.020 170.180 ;
        RECT 69.140 170.090 69.400 170.410 ;
        RECT 71.900 170.090 72.160 170.410 ;
        RECT 68.680 169.750 68.940 170.070 ;
        RECT 68.740 167.690 68.880 169.750 ;
        RECT 71.440 169.070 71.700 169.390 ;
        RECT 68.680 167.370 68.940 167.690 ;
        RECT 66.380 165.330 66.640 165.650 ;
        RECT 63.620 164.650 63.880 164.970 ;
        RECT 64.080 164.650 64.340 164.970 ;
        RECT 65.000 163.630 65.260 163.950 ;
        RECT 65.060 161.910 65.200 163.630 ;
        RECT 65.000 161.590 65.260 161.910 ;
        RECT 65.460 161.590 65.720 161.910 ;
        RECT 63.160 160.910 63.420 161.230 ;
        RECT 62.240 159.550 62.500 159.870 ;
        RECT 61.320 158.190 61.580 158.510 ;
        RECT 61.780 158.190 62.040 158.510 ;
        RECT 61.380 156.470 61.520 158.190 ;
        RECT 61.840 157.150 61.980 158.190 ;
        RECT 63.220 157.490 63.360 160.910 ;
        RECT 65.520 159.530 65.660 161.590 ;
        RECT 65.460 159.210 65.720 159.530 ;
        RECT 63.160 157.170 63.420 157.490 ;
        RECT 61.780 156.830 62.040 157.150 ;
        RECT 61.320 156.150 61.580 156.470 ;
        RECT 62.700 156.380 62.960 156.470 ;
        RECT 63.220 156.380 63.360 157.170 ;
        RECT 66.440 156.810 66.580 165.330 ;
        RECT 67.300 164.990 67.560 165.310 ;
        RECT 63.620 156.490 63.880 156.810 ;
        RECT 66.380 156.490 66.640 156.810 ;
        RECT 62.700 156.240 63.360 156.380 ;
        RECT 62.700 156.150 62.960 156.240 ;
        RECT 61.780 155.470 62.040 155.790 ;
        RECT 61.840 151.030 61.980 155.470 ;
        RECT 63.160 153.770 63.420 154.090 ;
        RECT 61.320 150.710 61.580 151.030 ;
        RECT 61.780 150.710 62.040 151.030 ;
        RECT 60.860 150.030 61.120 150.350 ;
        RECT 60.920 149.330 61.060 150.030 ;
        RECT 61.380 149.330 61.520 150.710 ;
        RECT 62.240 150.600 62.500 150.690 ;
        RECT 63.220 150.600 63.360 153.770 ;
        RECT 63.680 152.130 63.820 156.490 ;
        RECT 64.540 156.150 64.800 156.470 ;
        RECT 64.080 155.470 64.340 155.790 ;
        RECT 64.140 153.070 64.280 155.470 ;
        RECT 64.600 154.090 64.740 156.150 ;
        RECT 64.540 153.770 64.800 154.090 ;
        RECT 64.080 152.750 64.340 153.070 ;
        RECT 65.000 152.750 65.260 153.070 ;
        RECT 63.680 152.050 64.280 152.130 ;
        RECT 63.680 151.990 64.340 152.050 ;
        RECT 64.080 151.730 64.340 151.990 ;
        RECT 62.240 150.460 63.360 150.600 ;
        RECT 62.240 150.370 62.500 150.460 ;
        RECT 60.860 149.010 61.120 149.330 ;
        RECT 61.320 149.010 61.580 149.330 ;
        RECT 60.860 148.330 61.120 148.650 ;
        RECT 60.920 145.590 61.060 148.330 ;
        RECT 63.220 146.610 63.360 150.460 ;
        RECT 65.060 148.990 65.200 152.750 ;
        RECT 65.920 150.370 66.180 150.690 ;
        RECT 65.000 148.670 65.260 148.990 ;
        RECT 63.160 146.290 63.420 146.610 ;
        RECT 60.400 145.270 60.660 145.590 ;
        RECT 60.860 145.270 61.120 145.590 ;
        RECT 65.460 145.270 65.720 145.590 ;
        RECT 60.460 143.210 60.600 145.270 ;
        RECT 60.920 143.890 61.060 145.270 ;
        RECT 61.320 144.930 61.580 145.250 ;
        RECT 65.000 144.930 65.260 145.250 ;
        RECT 60.860 143.570 61.120 143.890 ;
        RECT 61.380 143.210 61.520 144.930 ;
        RECT 57.180 142.890 57.440 143.210 ;
        RECT 59.940 142.890 60.200 143.210 ;
        RECT 60.400 142.890 60.660 143.210 ;
        RECT 61.320 142.890 61.580 143.210 ;
        RECT 55.400 141.170 56.920 141.250 ;
        RECT 57.240 141.170 57.380 142.890 ;
        RECT 58.560 142.550 58.820 142.870 ;
        RECT 55.340 141.110 56.920 141.170 ;
        RECT 55.340 140.850 55.600 141.110 ;
        RECT 56.260 140.510 56.520 140.830 ;
        RECT 54.420 140.005 54.680 140.150 ;
        RECT 54.410 139.635 54.690 140.005 ;
        RECT 55.800 139.490 56.060 139.810 ;
        RECT 54.420 139.150 54.680 139.470 ;
        RECT 54.480 135.730 54.620 139.150 ;
        RECT 55.860 137.430 56.000 139.490 ;
        RECT 56.320 137.770 56.460 140.510 ;
        RECT 56.780 139.470 56.920 141.110 ;
        RECT 57.180 140.850 57.440 141.170 ;
        RECT 58.620 140.490 58.760 142.550 ;
        RECT 60.000 141.930 60.140 142.890 ;
        RECT 59.540 141.790 60.140 141.930 ;
        RECT 58.560 140.170 58.820 140.490 ;
        RECT 56.720 139.150 56.980 139.470 ;
        RECT 56.260 137.450 56.520 137.770 ;
        RECT 55.800 137.110 56.060 137.430 ;
        RECT 56.780 136.750 56.920 139.150 ;
        RECT 58.620 137.770 58.760 140.170 ;
        RECT 59.020 139.490 59.280 139.810 ;
        RECT 59.080 138.110 59.220 139.490 ;
        RECT 59.020 137.790 59.280 138.110 ;
        RECT 58.560 137.450 58.820 137.770 ;
        RECT 56.720 136.430 56.980 136.750 ;
        RECT 54.420 135.410 54.680 135.730 ;
        RECT 54.480 133.010 54.620 135.410 ;
        RECT 54.420 132.690 54.680 133.010 ;
        RECT 54.480 128.590 54.620 132.690 ;
        RECT 58.620 132.410 58.760 137.450 ;
        RECT 58.160 132.330 58.760 132.410 ;
        RECT 58.100 132.270 58.760 132.330 ;
        RECT 58.100 132.010 58.360 132.270 ;
        RECT 55.340 130.990 55.600 131.310 ;
        RECT 55.400 128.930 55.540 130.990 ;
        RECT 58.160 129.270 58.300 132.010 ;
        RECT 58.100 128.950 58.360 129.270 ;
        RECT 55.340 128.610 55.600 128.930 ;
        RECT 54.420 128.270 54.680 128.590 ;
        RECT 56.720 122.830 56.980 123.150 ;
        RECT 56.780 121.450 56.920 122.830 ;
        RECT 58.160 121.790 58.300 128.950 ;
        RECT 58.100 121.470 58.360 121.790 ;
        RECT 56.720 121.130 56.980 121.450 ;
        RECT 58.160 118.390 58.300 121.470 ;
        RECT 58.100 118.070 58.360 118.390 ;
        RECT 53.960 117.730 54.220 118.050 ;
        RECT 57.180 117.390 57.440 117.710 ;
        RECT 51.660 115.690 51.920 116.010 ;
        RECT 51.720 106.830 51.860 115.690 ;
        RECT 57.240 112.610 57.380 117.390 ;
        RECT 57.640 113.650 57.900 113.970 ;
        RECT 57.180 112.290 57.440 112.610 ;
        RECT 56.260 111.950 56.520 112.270 ;
        RECT 56.320 110.570 56.460 111.950 ;
        RECT 57.240 110.570 57.380 112.290 ;
        RECT 57.700 110.570 57.840 113.650 ;
        RECT 58.160 113.290 58.300 118.070 ;
        RECT 58.100 112.970 58.360 113.290 ;
        RECT 56.260 110.250 56.520 110.570 ;
        RECT 57.180 110.250 57.440 110.570 ;
        RECT 57.640 110.250 57.900 110.570 ;
        RECT 51.660 106.510 51.920 106.830 ;
        RECT 51.200 96.650 51.460 96.970 ;
        RECT 51.720 93.140 51.860 106.510 ;
        RECT 56.320 105.470 56.460 110.250 ;
        RECT 56.720 109.910 56.980 110.230 ;
        RECT 56.780 107.170 56.920 109.910 ;
        RECT 59.080 108.530 59.220 137.790 ;
        RECT 59.540 135.050 59.680 141.790 ;
        RECT 60.860 139.210 61.120 139.470 ;
        RECT 61.380 139.210 61.520 142.890 ;
        RECT 61.780 140.170 62.040 140.490 ;
        RECT 60.860 139.150 61.520 139.210 ;
        RECT 60.920 139.070 61.520 139.150 ;
        RECT 59.940 138.130 60.200 138.450 ;
        RECT 60.000 135.050 60.140 138.130 ;
        RECT 59.480 134.730 59.740 135.050 ;
        RECT 59.940 134.730 60.200 135.050 ;
        RECT 60.920 130.290 61.060 139.070 ;
        RECT 61.320 137.790 61.580 138.110 ;
        RECT 61.380 134.710 61.520 137.790 ;
        RECT 61.840 134.710 61.980 140.170 ;
        RECT 63.620 139.830 63.880 140.150 ;
        RECT 63.680 134.710 63.820 139.830 ;
        RECT 65.060 139.810 65.200 144.930 ;
        RECT 65.520 143.890 65.660 145.270 ;
        RECT 65.460 143.570 65.720 143.890 ;
        RECT 65.000 139.490 65.260 139.810 ;
        RECT 65.980 139.470 66.120 150.370 ;
        RECT 66.440 148.990 66.580 156.490 ;
        RECT 66.840 156.150 67.100 156.470 ;
        RECT 66.900 154.090 67.040 156.150 ;
        RECT 66.840 153.770 67.100 154.090 ;
        RECT 66.380 148.670 66.640 148.990 ;
        RECT 66.900 148.650 67.040 153.770 ;
        RECT 66.840 148.330 67.100 148.650 ;
        RECT 67.360 145.250 67.500 164.990 ;
        RECT 68.740 156.810 68.880 167.370 ;
        RECT 70.060 161.590 70.320 161.910 ;
        RECT 70.980 161.590 71.240 161.910 ;
        RECT 70.120 156.890 70.260 161.590 ;
        RECT 71.040 158.850 71.180 161.590 ;
        RECT 70.980 158.530 71.240 158.850 ;
        RECT 68.680 156.490 68.940 156.810 ;
        RECT 70.120 156.750 71.180 156.890 ;
        RECT 68.740 154.090 68.880 156.490 ;
        RECT 70.060 156.150 70.320 156.470 ;
        RECT 70.120 154.090 70.260 156.150 ;
        RECT 71.040 154.430 71.180 156.750 ;
        RECT 70.980 154.110 71.240 154.430 ;
        RECT 68.680 153.770 68.940 154.090 ;
        RECT 70.060 153.770 70.320 154.090 ;
        RECT 70.120 153.410 70.260 153.770 ;
        RECT 70.060 153.090 70.320 153.410 ;
        RECT 71.040 153.070 71.180 154.110 ;
        RECT 69.600 152.750 69.860 153.070 ;
        RECT 70.980 152.750 71.240 153.070 ;
        RECT 69.660 151.030 69.800 152.750 ;
        RECT 67.760 150.710 68.020 151.030 ;
        RECT 69.600 150.710 69.860 151.030 ;
        RECT 67.820 148.650 67.960 150.710 ;
        RECT 68.680 150.370 68.940 150.690 ;
        RECT 68.740 148.650 68.880 150.370 ;
        RECT 67.760 148.330 68.020 148.650 ;
        RECT 68.680 148.330 68.940 148.650 ;
        RECT 68.220 147.990 68.480 148.310 ;
        RECT 67.300 144.930 67.560 145.250 ;
        RECT 68.280 143.210 68.420 147.990 ;
        RECT 69.660 146.010 69.800 150.710 ;
        RECT 71.500 148.990 71.640 169.070 ;
        RECT 71.960 168.370 72.100 170.090 ;
        RECT 71.900 168.050 72.160 168.370 ;
        RECT 72.420 167.010 72.560 175.190 ;
        RECT 72.880 174.830 73.020 177.910 ;
        RECT 73.340 175.850 73.480 181.650 ;
        RECT 73.740 175.870 74.000 176.190 ;
        RECT 73.280 175.530 73.540 175.850 ;
        RECT 72.820 174.510 73.080 174.830 ;
        RECT 73.340 173.810 73.480 175.530 ;
        RECT 73.280 173.490 73.540 173.810 ;
        RECT 72.820 173.150 73.080 173.470 ;
        RECT 73.340 173.325 73.480 173.490 ;
        RECT 72.880 172.110 73.020 173.150 ;
        RECT 73.270 172.955 73.550 173.325 ;
        RECT 73.800 172.790 73.940 175.870 ;
        RECT 74.660 175.530 74.920 175.850 ;
        RECT 74.720 173.470 74.860 175.530 ;
        RECT 76.500 173.490 76.760 173.810 ;
        RECT 74.660 173.150 74.920 173.470 ;
        RECT 73.740 172.470 74.000 172.790 ;
        RECT 74.720 172.110 74.860 173.150 ;
        RECT 76.560 172.450 76.700 173.490 ;
        RECT 77.480 173.130 77.620 183.690 ;
        RECT 100.970 182.410 102.630 184.070 ;
        RECT 123.240 180.480 125.770 180.490 ;
        RECT 100.360 180.380 108.770 180.390 ;
        RECT 100.360 180.100 108.805 180.380 ;
        RECT 123.240 180.200 125.805 180.480 ;
        RECT 123.240 180.190 125.770 180.200 ;
        RECT 100.360 180.090 108.770 180.100 ;
        RECT 77.420 172.810 77.680 173.130 ;
        RECT 76.500 172.130 76.760 172.450 ;
        RECT 72.820 171.790 73.080 172.110 ;
        RECT 73.280 171.790 73.540 172.110 ;
        RECT 73.740 171.790 74.000 172.110 ;
        RECT 74.660 171.790 74.920 172.110 ;
        RECT 73.340 168.370 73.480 171.790 ;
        RECT 73.280 168.050 73.540 168.370 ;
        RECT 73.800 167.010 73.940 171.790 ;
        RECT 77.480 170.410 77.620 172.810 ;
        RECT 77.420 170.090 77.680 170.410 ;
        RECT 77.480 167.350 77.620 170.090 ;
        RECT 77.420 167.030 77.680 167.350 ;
        RECT 72.360 166.690 72.620 167.010 ;
        RECT 73.740 166.690 74.000 167.010 ;
        RECT 77.480 165.310 77.620 167.030 ;
        RECT 77.420 164.990 77.680 165.310 ;
        RECT 72.360 161.590 72.620 161.910 ;
        RECT 72.820 161.590 73.080 161.910 ;
        RECT 71.900 158.530 72.160 158.850 ;
        RECT 71.960 157.490 72.100 158.530 ;
        RECT 71.900 157.170 72.160 157.490 ;
        RECT 71.900 156.150 72.160 156.470 ;
        RECT 71.960 154.770 72.100 156.150 ;
        RECT 71.900 154.450 72.160 154.770 ;
        RECT 72.420 151.710 72.560 161.590 ;
        RECT 72.880 159.190 73.020 161.590 ;
        RECT 77.480 161.570 77.620 164.990 ;
        RECT 77.480 161.430 78.540 161.570 ;
        RECT 74.660 160.910 74.920 161.230 ;
        RECT 74.720 159.870 74.860 160.910 ;
        RECT 73.740 159.550 74.000 159.870 ;
        RECT 74.660 159.550 74.920 159.870 ;
        RECT 75.580 159.550 75.840 159.870 ;
        RECT 72.820 158.870 73.080 159.190 ;
        RECT 72.820 158.190 73.080 158.510 ;
        RECT 72.880 157.150 73.020 158.190 ;
        RECT 72.820 156.830 73.080 157.150 ;
        RECT 72.360 151.390 72.620 151.710 ;
        RECT 72.360 150.030 72.620 150.350 ;
        RECT 71.440 148.670 71.700 148.990 ;
        RECT 71.900 148.330 72.160 148.650 ;
        RECT 71.440 147.990 71.700 148.310 ;
        RECT 69.200 145.870 69.800 146.010 ;
        RECT 66.380 142.890 66.640 143.210 ;
        RECT 68.220 142.890 68.480 143.210 ;
        RECT 66.440 140.150 66.580 142.890 ;
        RECT 66.380 139.830 66.640 140.150 ;
        RECT 66.840 139.490 67.100 139.810 ;
        RECT 65.920 139.150 66.180 139.470 ;
        RECT 65.980 138.360 66.120 139.150 ;
        RECT 65.980 138.220 66.580 138.360 ;
        RECT 65.920 137.450 66.180 137.770 ;
        RECT 65.980 135.730 66.120 137.450 ;
        RECT 66.440 137.090 66.580 138.220 ;
        RECT 66.380 136.770 66.640 137.090 ;
        RECT 66.440 135.730 66.580 136.770 ;
        RECT 65.920 135.410 66.180 135.730 ;
        RECT 66.380 135.410 66.640 135.730 ;
        RECT 65.000 135.070 65.260 135.390 ;
        RECT 61.320 134.390 61.580 134.710 ;
        RECT 61.780 134.390 62.040 134.710 ;
        RECT 63.620 134.390 63.880 134.710 ;
        RECT 61.320 133.710 61.580 134.030 ;
        RECT 61.380 132.670 61.520 133.710 ;
        RECT 63.680 133.010 63.820 134.390 ;
        RECT 63.620 132.690 63.880 133.010 ;
        RECT 61.320 132.350 61.580 132.670 ;
        RECT 60.860 129.970 61.120 130.290 ;
        RECT 65.060 129.270 65.200 135.070 ;
        RECT 66.900 134.370 67.040 139.490 ;
        RECT 68.280 139.470 68.420 142.890 ;
        RECT 69.200 139.810 69.340 145.870 ;
        RECT 69.600 144.930 69.860 145.250 ;
        RECT 70.980 144.930 71.240 145.250 ;
        RECT 69.660 142.870 69.800 144.930 ;
        RECT 69.600 142.550 69.860 142.870 ;
        RECT 69.140 139.490 69.400 139.810 ;
        RECT 68.220 139.380 68.480 139.470 ;
        RECT 67.820 139.240 68.480 139.380 ;
        RECT 67.820 134.370 67.960 139.240 ;
        RECT 68.220 139.150 68.480 139.240 ;
        RECT 68.220 137.450 68.480 137.770 ;
        RECT 68.280 135.730 68.420 137.450 ;
        RECT 68.680 136.430 68.940 136.750 ;
        RECT 68.220 135.410 68.480 135.730 ;
        RECT 66.840 134.050 67.100 134.370 ;
        RECT 67.760 134.050 68.020 134.370 ;
        RECT 67.820 133.010 67.960 134.050 ;
        RECT 67.760 132.690 68.020 133.010 ;
        RECT 67.760 132.010 68.020 132.330 ;
        RECT 67.820 130.290 67.960 132.010 ;
        RECT 67.760 129.970 68.020 130.290 ;
        RECT 68.740 129.610 68.880 136.430 ;
        RECT 69.200 135.730 69.340 139.490 ;
        RECT 69.140 135.410 69.400 135.730 ;
        RECT 69.660 132.670 69.800 142.550 ;
        RECT 71.040 138.450 71.180 144.930 ;
        RECT 70.980 138.130 71.240 138.450 ;
        RECT 71.500 138.110 71.640 147.990 ;
        RECT 71.960 140.005 72.100 148.330 ;
        RECT 72.420 148.310 72.560 150.030 ;
        RECT 72.880 149.330 73.020 156.830 ;
        RECT 73.280 155.470 73.540 155.790 ;
        RECT 72.820 149.010 73.080 149.330 ;
        RECT 73.340 148.650 73.480 155.470 ;
        RECT 73.800 154.430 73.940 159.550 ;
        RECT 74.200 157.170 74.460 157.490 ;
        RECT 74.260 156.470 74.400 157.170 ;
        RECT 75.120 156.830 75.380 157.150 ;
        RECT 75.180 156.470 75.320 156.830 ;
        RECT 74.200 156.150 74.460 156.470 ;
        RECT 75.120 156.150 75.380 156.470 ;
        RECT 73.740 154.110 74.000 154.430 ;
        RECT 73.800 153.750 73.940 154.110 ;
        RECT 73.740 153.430 74.000 153.750 ;
        RECT 73.740 151.390 74.000 151.710 ;
        RECT 73.280 148.330 73.540 148.650 ;
        RECT 72.360 147.990 72.620 148.310 ;
        RECT 73.800 145.590 73.940 151.390 ;
        RECT 74.260 150.770 74.400 156.150 ;
        RECT 74.660 154.450 74.920 154.770 ;
        RECT 74.720 153.490 74.860 154.450 ;
        RECT 74.720 153.350 75.320 153.490 ;
        RECT 75.180 151.030 75.320 153.350 ;
        RECT 74.260 150.630 74.860 150.770 ;
        RECT 75.120 150.710 75.380 151.030 ;
        RECT 74.720 146.270 74.860 150.630 ;
        RECT 75.120 147.990 75.380 148.310 ;
        RECT 74.660 145.950 74.920 146.270 ;
        RECT 75.180 145.930 75.320 147.990 ;
        RECT 75.120 145.610 75.380 145.930 ;
        RECT 73.740 145.270 74.000 145.590 ;
        RECT 75.640 145.250 75.780 159.550 ;
        RECT 78.400 158.510 78.540 161.430 ;
        RECT 78.340 158.190 78.600 158.510 ;
        RECT 80.180 158.190 80.440 158.510 ;
        RECT 78.400 156.810 78.540 158.190 ;
        RECT 77.880 156.490 78.140 156.810 ;
        RECT 78.340 156.490 78.600 156.810 ;
        RECT 76.500 153.430 76.760 153.750 ;
        RECT 76.040 153.090 76.300 153.410 ;
        RECT 76.100 151.030 76.240 153.090 ;
        RECT 76.040 150.710 76.300 151.030 ;
        RECT 76.560 145.250 76.700 153.430 ;
        RECT 77.940 153.410 78.080 156.490 ;
        RECT 78.340 155.470 78.600 155.790 ;
        RECT 78.400 154.430 78.540 155.470 ;
        RECT 78.340 154.110 78.600 154.430 ;
        RECT 80.240 154.090 80.380 158.190 ;
        RECT 80.180 153.770 80.440 154.090 ;
        RECT 77.880 153.090 78.140 153.410 ;
        RECT 82.020 150.710 82.280 151.030 ;
        RECT 82.080 149.330 82.220 150.710 ;
        RECT 82.020 149.010 82.280 149.330 ;
        RECT 76.960 145.270 77.220 145.590 ;
        RECT 75.580 144.930 75.840 145.250 ;
        RECT 76.500 144.930 76.760 145.250 ;
        RECT 72.360 144.590 72.620 144.910 ;
        RECT 72.420 143.550 72.560 144.590 ;
        RECT 76.560 143.890 76.700 144.930 ;
        RECT 76.500 143.570 76.760 143.890 ;
        RECT 72.360 143.230 72.620 143.550 ;
        RECT 71.890 139.635 72.170 140.005 ;
        RECT 70.060 137.790 70.320 138.110 ;
        RECT 71.440 137.790 71.700 138.110 ;
        RECT 70.120 137.430 70.260 137.790 ;
        RECT 70.060 137.110 70.320 137.430 ;
        RECT 71.440 137.170 71.700 137.430 ;
        RECT 71.960 137.170 72.100 139.635 ;
        RECT 77.020 137.770 77.160 145.270 ;
        RECT 76.960 137.450 77.220 137.770 ;
        RECT 77.420 137.450 77.680 137.770 ;
        RECT 71.440 137.110 72.100 137.170 ;
        RECT 73.280 137.110 73.540 137.430 ;
        RECT 69.600 132.350 69.860 132.670 ;
        RECT 70.120 129.950 70.260 137.110 ;
        RECT 71.500 137.030 72.100 137.110 ;
        RECT 73.340 135.730 73.480 137.110 ;
        RECT 73.280 135.410 73.540 135.730 ;
        RECT 77.480 134.280 77.620 137.450 ;
        RECT 76.560 134.140 77.620 134.280 ;
        RECT 76.560 132.670 76.700 134.140 ;
        RECT 74.200 132.350 74.460 132.670 ;
        RECT 76.500 132.350 76.760 132.670 ;
        RECT 70.060 129.630 70.320 129.950 ;
        RECT 68.680 129.290 68.940 129.610 ;
        RECT 65.000 128.950 65.260 129.270 ;
        RECT 59.940 123.510 60.200 123.830 ;
        RECT 67.760 123.510 68.020 123.830 ;
        RECT 68.220 123.510 68.480 123.830 ;
        RECT 69.140 123.740 69.400 123.830 ;
        RECT 68.740 123.600 69.400 123.740 ;
        RECT 60.000 116.690 60.140 123.510 ;
        RECT 65.920 123.170 66.180 123.490 ;
        RECT 61.780 122.830 62.040 123.150 ;
        RECT 61.840 118.390 61.980 122.830 ;
        RECT 61.780 118.070 62.040 118.390 ;
        RECT 59.940 116.370 60.200 116.690 ;
        RECT 65.980 116.010 66.120 123.170 ;
        RECT 67.300 121.130 67.560 121.450 ;
        RECT 67.360 119.410 67.500 121.130 ;
        RECT 67.820 119.410 67.960 123.510 ;
        RECT 67.300 119.090 67.560 119.410 ;
        RECT 67.760 119.090 68.020 119.410 ;
        RECT 66.380 117.730 66.640 118.050 ;
        RECT 66.440 116.690 66.580 117.730 ;
        RECT 68.280 116.690 68.420 123.510 ;
        RECT 68.740 120.430 68.880 123.600 ;
        RECT 69.140 123.510 69.400 123.600 ;
        RECT 74.260 121.450 74.400 132.350 ;
        RECT 73.740 121.130 74.000 121.450 ;
        RECT 74.200 121.130 74.460 121.450 ;
        RECT 76.960 121.130 77.220 121.450 ;
        RECT 68.680 120.110 68.940 120.430 ;
        RECT 68.740 118.390 68.880 120.110 ;
        RECT 73.800 119.410 73.940 121.130 ;
        RECT 73.740 119.090 74.000 119.410 ;
        RECT 68.680 118.070 68.940 118.390 ;
        RECT 71.900 118.070 72.160 118.390 ;
        RECT 73.280 118.070 73.540 118.390 ;
        RECT 66.380 116.370 66.640 116.690 ;
        RECT 68.220 116.370 68.480 116.690 ;
        RECT 65.920 115.690 66.180 116.010 ;
        RECT 68.680 115.690 68.940 116.010 ;
        RECT 70.060 115.690 70.320 116.010 ;
        RECT 65.980 113.270 66.120 115.690 ;
        RECT 65.060 113.130 66.120 113.270 ;
        RECT 64.540 112.630 64.800 112.950 ;
        RECT 64.600 111.250 64.740 112.630 ;
        RECT 65.060 112.270 65.200 113.130 ;
        RECT 68.740 112.270 68.880 115.690 ;
        RECT 70.120 113.630 70.260 115.690 ;
        RECT 71.960 115.670 72.100 118.070 ;
        RECT 72.820 117.730 73.080 118.050 ;
        RECT 71.900 115.350 72.160 115.670 ;
        RECT 70.060 113.310 70.320 113.630 ;
        RECT 65.000 111.950 65.260 112.270 ;
        RECT 66.840 111.950 67.100 112.270 ;
        RECT 68.680 111.950 68.940 112.270 ;
        RECT 69.140 111.950 69.400 112.270 ;
        RECT 65.060 111.250 65.200 111.950 ;
        RECT 64.540 110.930 64.800 111.250 ;
        RECT 65.000 110.930 65.260 111.250 ;
        RECT 63.620 110.250 63.880 110.570 ;
        RECT 63.680 108.530 63.820 110.250 ;
        RECT 66.900 110.230 67.040 111.950 ;
        RECT 66.840 109.910 67.100 110.230 ;
        RECT 67.760 109.910 68.020 110.230 ;
        RECT 64.080 109.570 64.340 109.890 ;
        RECT 59.020 108.210 59.280 108.530 ;
        RECT 63.620 108.210 63.880 108.530 ;
        RECT 57.180 107.870 57.440 108.190 ;
        RECT 56.720 106.850 56.980 107.170 ;
        RECT 56.260 105.150 56.520 105.470 ;
        RECT 53.960 104.470 54.220 104.790 ;
        RECT 55.340 104.470 55.600 104.790 ;
        RECT 52.120 103.790 52.380 104.110 ;
        RECT 52.180 96.630 52.320 103.790 ;
        RECT 54.020 100.370 54.160 104.470 ;
        RECT 55.400 103.090 55.540 104.470 ;
        RECT 55.340 102.770 55.600 103.090 ;
        RECT 53.960 100.050 54.220 100.370 ;
        RECT 52.120 96.310 52.380 96.630 ;
        RECT 55.400 96.290 55.540 102.770 ;
        RECT 55.800 101.410 56.060 101.730 ;
        RECT 55.860 98.670 56.000 101.410 ;
        RECT 56.320 99.690 56.460 105.150 ;
        RECT 56.780 104.110 56.920 106.850 ;
        RECT 57.240 105.810 57.380 107.870 ;
        RECT 57.180 105.490 57.440 105.810 ;
        RECT 56.720 103.790 56.980 104.110 ;
        RECT 56.780 100.030 56.920 103.790 ;
        RECT 57.180 101.750 57.440 102.070 ;
        RECT 56.720 99.710 56.980 100.030 ;
        RECT 56.260 99.370 56.520 99.690 ;
        RECT 57.240 99.010 57.380 101.750 ;
        RECT 57.180 98.690 57.440 99.010 ;
        RECT 55.800 98.350 56.060 98.670 ;
        RECT 55.860 96.970 56.000 98.350 ;
        RECT 55.800 96.650 56.060 96.970 ;
        RECT 55.340 95.970 55.600 96.290 ;
        RECT 55.860 93.910 56.000 96.650 ;
        RECT 55.800 93.590 56.060 93.910 ;
        RECT 57.240 93.230 57.380 98.690 ;
        RECT 58.560 96.650 58.820 96.970 ;
        RECT 51.260 93.000 51.860 93.140 ;
        RECT 51.260 86.430 51.400 93.000 ;
        RECT 57.180 92.910 57.440 93.230 ;
        RECT 52.580 90.530 52.840 90.850 ;
        RECT 52.640 89.490 52.780 90.530 ;
        RECT 52.120 89.170 52.380 89.490 ;
        RECT 52.580 89.170 52.840 89.490 ;
        RECT 52.180 88.810 52.320 89.170 ;
        RECT 56.720 88.830 56.980 89.150 ;
        RECT 52.120 88.490 52.380 88.810 ;
        RECT 51.200 86.110 51.460 86.430 ;
        RECT 51.260 74.610 51.400 86.110 ;
        RECT 52.180 79.970 52.320 88.490 ;
        RECT 53.500 87.810 53.760 88.130 ;
        RECT 53.040 85.090 53.300 85.410 ;
        RECT 52.580 84.750 52.840 85.070 ;
        RECT 52.640 83.710 52.780 84.750 ;
        RECT 52.580 83.390 52.840 83.710 ;
        RECT 53.100 81.330 53.240 85.090 ;
        RECT 53.040 81.010 53.300 81.330 ;
        RECT 52.120 79.650 52.380 79.970 ;
        RECT 51.660 79.310 51.920 79.630 ;
        RECT 51.720 75.210 51.860 79.310 ;
        RECT 52.120 77.950 52.380 78.270 ;
        RECT 52.180 75.890 52.320 77.950 ;
        RECT 53.040 77.610 53.300 77.930 ;
        RECT 52.580 76.590 52.840 76.910 ;
        RECT 52.120 75.570 52.380 75.890 ;
        RECT 51.660 74.890 51.920 75.210 ;
        RECT 51.260 74.470 51.860 74.610 ;
        RECT 51.200 66.390 51.460 66.710 ;
        RECT 51.260 62.290 51.400 66.390 ;
        RECT 51.720 63.990 51.860 74.470 ;
        RECT 52.180 69.770 52.320 75.570 ;
        RECT 52.640 74.870 52.780 76.590 ;
        RECT 53.100 75.890 53.240 77.610 ;
        RECT 53.040 75.570 53.300 75.890 ;
        RECT 52.580 74.550 52.840 74.870 ;
        RECT 52.120 69.450 52.380 69.770 ;
        RECT 52.640 64.330 52.780 74.550 ;
        RECT 53.560 72.830 53.700 87.810 ;
        RECT 55.800 85.770 56.060 86.090 ;
        RECT 54.420 84.750 54.680 85.070 ;
        RECT 54.480 81.330 54.620 84.750 ;
        RECT 54.420 81.010 54.680 81.330 ;
        RECT 55.340 79.310 55.600 79.630 ;
        RECT 54.420 73.870 54.680 74.190 ;
        RECT 53.500 72.510 53.760 72.830 ;
        RECT 53.560 72.150 53.700 72.510 ;
        RECT 53.500 71.830 53.760 72.150 ;
        RECT 54.480 67.730 54.620 73.870 ;
        RECT 55.400 69.770 55.540 79.310 ;
        RECT 55.860 78.270 56.000 85.770 ;
        RECT 56.780 84.050 56.920 88.830 ;
        RECT 57.240 88.470 57.380 92.910 ;
        RECT 57.180 88.150 57.440 88.470 ;
        RECT 57.240 86.090 57.380 88.150 ;
        RECT 57.180 85.770 57.440 86.090 ;
        RECT 56.720 83.730 56.980 84.050 ;
        RECT 55.800 77.950 56.060 78.270 ;
        RECT 55.860 75.210 56.000 77.950 ;
        RECT 55.800 74.890 56.060 75.210 ;
        RECT 55.860 71.720 56.000 74.890 ;
        RECT 57.240 74.870 57.380 85.770 ;
        RECT 57.640 84.750 57.900 85.070 ;
        RECT 57.700 84.050 57.840 84.750 ;
        RECT 57.640 83.730 57.900 84.050 ;
        RECT 58.620 80.650 58.760 96.650 ;
        RECT 58.560 80.330 58.820 80.650 ;
        RECT 58.100 79.990 58.360 80.310 ;
        RECT 58.160 78.610 58.300 79.990 ;
        RECT 58.100 78.290 58.360 78.610 ;
        RECT 57.180 74.550 57.440 74.870 ;
        RECT 57.640 72.170 57.900 72.490 ;
        RECT 56.260 71.720 56.520 71.810 ;
        RECT 55.860 71.580 56.520 71.720 ;
        RECT 56.260 71.490 56.520 71.580 ;
        RECT 55.340 69.450 55.600 69.770 ;
        RECT 57.180 68.770 57.440 69.090 ;
        RECT 57.240 67.730 57.380 68.770 ;
        RECT 54.420 67.410 54.680 67.730 ;
        RECT 57.180 67.410 57.440 67.730 ;
        RECT 53.040 66.050 53.300 66.370 ;
        RECT 52.580 64.010 52.840 64.330 ;
        RECT 51.660 63.670 51.920 63.990 ;
        RECT 52.580 62.990 52.840 63.310 ;
        RECT 51.200 61.970 51.460 62.290 ;
        RECT 51.260 58.550 51.400 61.970 ;
        RECT 52.640 61.270 52.780 62.990 ;
        RECT 53.100 62.290 53.240 66.050 ;
        RECT 55.340 63.330 55.600 63.650 ;
        RECT 55.400 62.290 55.540 63.330 ;
        RECT 53.040 61.970 53.300 62.290 ;
        RECT 55.340 61.970 55.600 62.290 ;
        RECT 52.580 60.950 52.840 61.270 ;
        RECT 55.800 60.950 56.060 61.270 ;
        RECT 51.200 58.230 51.460 58.550 ;
        RECT 55.340 57.890 55.600 58.210 ;
        RECT 55.400 56.510 55.540 57.890 ;
        RECT 55.340 56.190 55.600 56.510 ;
        RECT 53.500 55.510 53.760 55.830 ;
        RECT 54.880 55.510 55.140 55.830 ;
        RECT 52.580 54.830 52.840 55.150 ;
        RECT 51.660 52.790 51.920 53.110 ;
        RECT 50.740 49.730 51.000 50.050 ;
        RECT 50.800 48.010 50.940 49.730 ;
        RECT 50.740 47.690 51.000 48.010 ;
        RECT 51.200 41.570 51.460 41.890 ;
        RECT 51.260 39.510 51.400 41.570 ;
        RECT 51.200 39.190 51.460 39.510 ;
        RECT 50.740 38.510 51.000 38.830 ;
        RECT 50.800 31.090 50.940 38.510 ;
        RECT 51.260 37.130 51.400 39.190 ;
        RECT 51.200 36.810 51.460 37.130 ;
        RECT 51.200 34.770 51.460 35.090 ;
        RECT 51.260 31.770 51.400 34.770 ;
        RECT 51.720 32.370 51.860 52.790 ;
        RECT 52.640 51.070 52.780 54.830 ;
        RECT 52.580 50.750 52.840 51.070 ;
        RECT 53.040 48.370 53.300 48.690 ;
        RECT 53.100 45.290 53.240 48.370 ;
        RECT 52.120 44.970 52.380 45.290 ;
        RECT 53.040 44.970 53.300 45.290 ;
        RECT 52.180 42.230 52.320 44.970 ;
        RECT 53.100 43.250 53.240 44.970 ;
        RECT 53.040 42.930 53.300 43.250 ;
        RECT 52.120 41.910 52.380 42.230 ;
        RECT 52.180 34.410 52.320 41.910 ;
        RECT 53.100 40.530 53.240 42.930 ;
        RECT 53.040 40.210 53.300 40.530 ;
        RECT 53.100 38.830 53.240 40.210 ;
        RECT 52.580 38.510 52.840 38.830 ;
        RECT 53.040 38.510 53.300 38.830 ;
        RECT 52.120 34.090 52.380 34.410 ;
        RECT 52.640 33.730 52.780 38.510 ;
        RECT 53.100 34.410 53.240 38.510 ;
        RECT 53.040 34.090 53.300 34.410 ;
        RECT 52.580 33.410 52.840 33.730 ;
        RECT 51.660 32.050 51.920 32.370 ;
        RECT 51.260 31.630 51.860 31.770 ;
        RECT 51.720 31.350 51.860 31.630 ;
        RECT 52.120 31.370 52.380 31.690 ;
        RECT 50.800 31.010 51.400 31.090 ;
        RECT 51.660 31.030 51.920 31.350 ;
        RECT 50.800 30.950 51.460 31.010 ;
        RECT 51.200 30.690 51.460 30.950 ;
        RECT 51.720 23.870 51.860 31.030 ;
        RECT 52.180 25.230 52.320 31.370 ;
        RECT 52.640 30.670 52.780 33.410 ;
        RECT 52.580 30.350 52.840 30.670 ;
        RECT 52.580 28.650 52.840 28.970 ;
        RECT 52.640 26.590 52.780 28.650 ;
        RECT 52.580 26.270 52.840 26.590 ;
        RECT 52.120 24.910 52.380 25.230 ;
        RECT 51.660 23.550 51.920 23.870 ;
        RECT 50.280 22.530 50.540 22.850 ;
        RECT 50.740 20.150 51.000 20.470 ;
        RECT 50.800 16.050 50.940 20.150 ;
        RECT 53.560 17.070 53.700 55.510 ;
        RECT 54.940 54.130 55.080 55.510 ;
        RECT 55.400 54.130 55.540 56.190 ;
        RECT 55.860 55.830 56.000 60.950 ;
        RECT 57.700 59.570 57.840 72.170 ;
        RECT 58.620 66.030 58.760 80.330 ;
        RECT 59.080 73.170 59.220 108.210 ;
        RECT 64.140 105.810 64.280 109.570 ;
        RECT 65.920 109.230 66.180 109.550 ;
        RECT 65.460 108.210 65.720 108.530 ;
        RECT 64.080 105.490 64.340 105.810 ;
        RECT 65.520 105.130 65.660 108.210 ;
        RECT 65.460 104.810 65.720 105.130 ;
        RECT 65.980 104.530 66.120 109.230 ;
        RECT 66.900 107.510 67.040 109.910 ;
        RECT 66.840 107.190 67.100 107.510 ;
        RECT 67.300 105.490 67.560 105.810 ;
        RECT 66.840 105.150 67.100 105.470 ;
        RECT 65.520 104.390 66.120 104.530 ;
        RECT 65.520 104.110 65.660 104.390 ;
        RECT 61.780 103.790 62.040 104.110 ;
        RECT 65.460 103.790 65.720 104.110 ;
        RECT 61.840 102.410 61.980 103.790 ;
        RECT 61.780 102.090 62.040 102.410 ;
        RECT 65.000 101.750 65.260 102.070 ;
        RECT 65.060 100.370 65.200 101.750 ;
        RECT 65.000 100.050 65.260 100.370 ;
        RECT 61.780 96.310 62.040 96.630 ;
        RECT 61.840 94.930 61.980 96.310 ;
        RECT 61.780 94.610 62.040 94.930 ;
        RECT 65.060 87.790 65.200 100.050 ;
        RECT 65.520 96.970 65.660 103.790 ;
        RECT 66.900 102.070 67.040 105.150 ;
        RECT 67.360 102.070 67.500 105.490 ;
        RECT 67.820 105.470 67.960 109.910 ;
        RECT 68.680 109.570 68.940 109.890 ;
        RECT 68.740 108.190 68.880 109.570 ;
        RECT 69.200 108.530 69.340 111.950 ;
        RECT 69.600 110.250 69.860 110.570 ;
        RECT 69.140 108.210 69.400 108.530 ;
        RECT 68.680 107.870 68.940 108.190 ;
        RECT 68.680 107.190 68.940 107.510 ;
        RECT 69.660 107.250 69.800 110.250 ;
        RECT 70.120 109.970 70.260 113.310 ;
        RECT 70.520 112.630 70.780 112.950 ;
        RECT 70.580 111.250 70.720 112.630 ;
        RECT 70.980 112.290 71.240 112.610 ;
        RECT 70.520 110.930 70.780 111.250 ;
        RECT 71.040 110.910 71.180 112.290 ;
        RECT 70.980 110.590 71.240 110.910 ;
        RECT 70.120 109.890 70.720 109.970 ;
        RECT 70.120 109.830 70.780 109.890 ;
        RECT 70.520 109.570 70.780 109.830 ;
        RECT 71.960 108.190 72.100 115.350 ;
        RECT 72.880 112.950 73.020 117.730 ;
        RECT 72.820 112.630 73.080 112.950 ;
        RECT 73.340 110.910 73.480 118.070 ;
        RECT 77.020 112.950 77.160 121.130 ;
        RECT 88.460 115.690 88.720 116.010 ;
        RECT 79.260 114.670 79.520 114.990 ;
        RECT 76.960 112.630 77.220 112.950 ;
        RECT 74.660 112.290 74.920 112.610 ;
        RECT 74.200 111.950 74.460 112.270 ;
        RECT 73.280 110.590 73.540 110.910 ;
        RECT 74.260 110.230 74.400 111.950 ;
        RECT 74.200 109.910 74.460 110.230 ;
        RECT 72.360 109.570 72.620 109.890 ;
        RECT 72.420 108.530 72.560 109.570 ;
        RECT 74.720 109.550 74.860 112.290 ;
        RECT 75.120 110.250 75.380 110.570 ;
        RECT 74.660 109.230 74.920 109.550 ;
        RECT 75.180 108.530 75.320 110.250 ;
        RECT 78.800 109.570 79.060 109.890 ;
        RECT 72.360 108.210 72.620 108.530 ;
        RECT 73.280 108.210 73.540 108.530 ;
        RECT 75.120 108.210 75.380 108.530 ;
        RECT 71.900 107.870 72.160 108.190 ;
        RECT 67.760 105.150 68.020 105.470 ;
        RECT 67.760 103.790 68.020 104.110 ;
        RECT 66.840 101.750 67.100 102.070 ;
        RECT 67.300 101.750 67.560 102.070 ;
        RECT 66.380 101.070 66.640 101.390 ;
        RECT 65.920 100.050 66.180 100.370 ;
        RECT 65.460 96.650 65.720 96.970 ;
        RECT 65.980 88.470 66.120 100.050 ;
        RECT 66.440 99.690 66.580 101.070 ;
        RECT 67.820 100.370 67.960 103.790 ;
        RECT 68.220 102.430 68.480 102.750 ;
        RECT 67.760 100.050 68.020 100.370 ;
        RECT 66.380 99.370 66.640 99.690 ;
        RECT 66.440 88.810 66.580 99.370 ;
        RECT 68.280 99.350 68.420 102.430 ;
        RECT 68.220 99.030 68.480 99.350 ;
        RECT 68.220 96.310 68.480 96.630 ;
        RECT 67.300 95.860 67.560 95.950 ;
        RECT 67.300 95.720 67.960 95.860 ;
        RECT 67.300 95.630 67.560 95.720 ;
        RECT 66.830 94.755 67.110 95.125 ;
        RECT 66.900 94.590 67.040 94.755 ;
        RECT 66.840 94.270 67.100 94.590 ;
        RECT 67.300 92.910 67.560 93.230 ;
        RECT 67.360 90.850 67.500 92.910 ;
        RECT 67.300 90.530 67.560 90.850 ;
        RECT 66.380 88.490 66.640 88.810 ;
        RECT 66.840 88.490 67.100 88.810 ;
        RECT 65.920 88.150 66.180 88.470 ;
        RECT 65.000 87.470 65.260 87.790 ;
        RECT 65.980 86.170 66.120 88.150 ;
        RECT 65.520 86.030 66.120 86.170 ;
        RECT 65.520 85.750 65.660 86.030 ;
        RECT 65.460 85.430 65.720 85.750 ;
        RECT 66.380 85.430 66.640 85.750 ;
        RECT 65.920 84.750 66.180 85.070 ;
        RECT 59.480 79.310 59.740 79.630 ;
        RECT 59.020 72.850 59.280 73.170 ;
        RECT 59.080 69.430 59.220 72.850 ;
        RECT 59.020 69.110 59.280 69.430 ;
        RECT 59.020 66.730 59.280 67.050 ;
        RECT 58.560 65.710 58.820 66.030 ;
        RECT 58.100 63.670 58.360 63.990 ;
        RECT 58.160 62.290 58.300 63.670 ;
        RECT 58.100 61.970 58.360 62.290 ;
        RECT 57.640 59.250 57.900 59.570 ;
        RECT 58.160 58.890 58.300 61.970 ;
        RECT 58.100 58.570 58.360 58.890 ;
        RECT 59.080 55.830 59.220 66.730 ;
        RECT 59.540 65.010 59.680 79.310 ;
        RECT 64.080 77.610 64.340 77.930 ;
        RECT 64.140 74.870 64.280 77.610 ;
        RECT 65.980 74.870 66.120 84.750 ;
        RECT 66.440 83.370 66.580 85.430 ;
        RECT 66.900 84.050 67.040 88.490 ;
        RECT 66.840 83.730 67.100 84.050 ;
        RECT 66.380 83.050 66.640 83.370 ;
        RECT 66.440 79.970 66.580 83.050 ;
        RECT 66.380 79.650 66.640 79.970 ;
        RECT 67.360 77.930 67.500 90.530 ;
        RECT 67.820 85.750 67.960 95.720 ;
        RECT 68.280 94.250 68.420 96.310 ;
        RECT 68.740 96.290 68.880 107.190 ;
        RECT 69.660 107.110 70.260 107.250 ;
        RECT 70.120 106.830 70.260 107.110 ;
        RECT 69.140 106.510 69.400 106.830 ;
        RECT 70.060 106.510 70.320 106.830 ;
        RECT 69.200 105.130 69.340 106.510 ;
        RECT 69.140 104.810 69.400 105.130 ;
        RECT 69.200 99.690 69.340 104.810 ;
        RECT 69.140 99.370 69.400 99.690 ;
        RECT 69.200 97.650 69.340 99.370 ;
        RECT 70.520 99.030 70.780 99.350 ;
        RECT 73.340 99.205 73.480 108.210 ;
        RECT 75.580 107.870 75.840 108.190 ;
        RECT 75.120 104.810 75.380 105.130 ;
        RECT 73.740 104.470 74.000 104.790 ;
        RECT 73.800 104.110 73.940 104.470 ;
        RECT 75.180 104.110 75.320 104.810 ;
        RECT 73.740 103.790 74.000 104.110 ;
        RECT 75.120 103.790 75.380 104.110 ;
        RECT 69.140 97.330 69.400 97.650 ;
        RECT 69.200 96.910 70.260 97.050 ;
        RECT 68.680 95.970 68.940 96.290 ;
        RECT 68.220 93.930 68.480 94.250 ;
        RECT 69.200 93.910 69.340 96.910 ;
        RECT 69.600 96.310 69.860 96.630 ;
        RECT 69.140 93.590 69.400 93.910 ;
        RECT 69.660 93.230 69.800 96.310 ;
        RECT 70.120 95.950 70.260 96.910 ;
        RECT 70.580 96.630 70.720 99.030 ;
        RECT 72.820 98.690 73.080 99.010 ;
        RECT 73.270 98.835 73.550 99.205 ;
        RECT 72.880 96.630 73.020 98.690 ;
        RECT 70.520 96.310 70.780 96.630 ;
        RECT 72.820 96.310 73.080 96.630 ;
        RECT 70.060 95.630 70.320 95.950 ;
        RECT 70.580 94.250 70.720 96.310 ;
        RECT 72.360 95.970 72.620 96.290 ;
        RECT 70.060 93.930 70.320 94.250 ;
        RECT 70.520 93.930 70.780 94.250 ;
        RECT 71.900 93.930 72.160 94.250 ;
        RECT 69.600 92.910 69.860 93.230 ;
        RECT 68.680 91.210 68.940 91.530 ;
        RECT 68.740 89.490 68.880 91.210 ;
        RECT 70.120 90.510 70.260 93.930 ;
        RECT 70.580 90.850 70.720 93.930 ;
        RECT 71.960 93.230 72.100 93.930 ;
        RECT 71.900 92.910 72.160 93.230 ;
        RECT 70.520 90.760 70.780 90.850 ;
        RECT 70.520 90.620 71.180 90.760 ;
        RECT 70.520 90.530 70.780 90.620 ;
        RECT 70.060 90.190 70.320 90.510 ;
        RECT 68.680 89.170 68.940 89.490 ;
        RECT 68.740 88.810 68.880 89.170 ;
        RECT 69.600 88.830 69.860 89.150 ;
        RECT 68.680 88.490 68.940 88.810 ;
        RECT 68.680 87.470 68.940 87.790 ;
        RECT 68.220 86.450 68.480 86.770 ;
        RECT 67.760 85.430 68.020 85.750 ;
        RECT 67.300 77.610 67.560 77.930 ;
        RECT 67.300 76.930 67.560 77.250 ;
        RECT 67.360 75.550 67.500 76.930 ;
        RECT 67.300 75.230 67.560 75.550 ;
        RECT 64.080 74.550 64.340 74.870 ;
        RECT 65.920 74.550 66.180 74.870 ;
        RECT 64.140 72.490 64.280 74.550 ;
        RECT 67.360 73.170 67.500 75.230 ;
        RECT 67.300 72.850 67.560 73.170 ;
        RECT 66.380 72.510 66.640 72.830 ;
        RECT 64.080 72.170 64.340 72.490 ;
        RECT 64.140 69.770 64.280 72.170 ;
        RECT 64.080 69.450 64.340 69.770 ;
        RECT 65.460 69.110 65.720 69.430 ;
        RECT 64.540 66.390 64.800 66.710 ;
        RECT 60.400 65.710 60.660 66.030 ;
        RECT 59.480 64.690 59.740 65.010 ;
        RECT 59.940 62.990 60.200 63.310 ;
        RECT 60.000 61.950 60.140 62.990 ;
        RECT 59.940 61.630 60.200 61.950 ;
        RECT 60.460 58.890 60.600 65.710 ;
        RECT 64.600 61.610 64.740 66.390 ;
        RECT 65.520 63.650 65.660 69.110 ;
        RECT 65.920 63.670 66.180 63.990 ;
        RECT 65.460 63.330 65.720 63.650 ;
        RECT 65.980 61.610 66.120 63.670 ;
        RECT 64.540 61.290 64.800 61.610 ;
        RECT 65.920 61.290 66.180 61.610 ;
        RECT 66.440 61.520 66.580 72.510 ;
        RECT 66.840 71.150 67.100 71.470 ;
        RECT 66.900 69.090 67.040 71.150 ;
        RECT 66.840 68.770 67.100 69.090 ;
        RECT 67.300 68.430 67.560 68.750 ;
        RECT 67.360 67.730 67.500 68.430 ;
        RECT 67.300 67.410 67.560 67.730 ;
        RECT 67.820 64.330 67.960 85.430 ;
        RECT 68.280 82.350 68.420 86.450 ;
        RECT 68.740 85.750 68.880 87.470 ;
        RECT 69.660 86.770 69.800 88.830 ;
        RECT 70.520 88.490 70.780 88.810 ;
        RECT 69.600 86.450 69.860 86.770 ;
        RECT 70.580 85.750 70.720 88.490 ;
        RECT 68.680 85.430 68.940 85.750 ;
        RECT 70.520 85.660 70.780 85.750 ;
        RECT 70.120 85.520 70.780 85.660 ;
        RECT 69.140 83.730 69.400 84.050 ;
        RECT 68.220 82.030 68.480 82.350 ;
        RECT 68.280 81.330 68.420 82.030 ;
        RECT 68.220 81.010 68.480 81.330 ;
        RECT 69.200 79.970 69.340 83.730 ;
        RECT 70.120 82.690 70.260 85.520 ;
        RECT 70.520 85.430 70.780 85.520 ;
        RECT 70.520 84.750 70.780 85.070 ;
        RECT 70.580 84.050 70.720 84.750 ;
        RECT 70.520 83.730 70.780 84.050 ;
        RECT 70.060 82.370 70.320 82.690 ;
        RECT 70.050 82.090 70.330 82.205 ;
        RECT 69.660 81.950 70.330 82.090 ;
        RECT 69.140 79.650 69.400 79.970 ;
        RECT 69.140 74.550 69.400 74.870 ;
        RECT 68.670 72.315 68.950 72.685 ;
        RECT 68.680 72.170 68.940 72.315 ;
        RECT 69.200 72.005 69.340 74.550 ;
        RECT 69.130 71.635 69.410 72.005 ;
        RECT 68.220 69.450 68.480 69.770 ;
        RECT 67.760 64.010 68.020 64.330 ;
        RECT 68.280 63.990 68.420 69.450 ;
        RECT 68.680 66.730 68.940 67.050 ;
        RECT 68.220 63.670 68.480 63.990 ;
        RECT 67.760 63.330 68.020 63.650 ;
        RECT 66.840 62.990 67.100 63.310 ;
        RECT 67.300 62.990 67.560 63.310 ;
        RECT 66.900 62.290 67.040 62.990 ;
        RECT 66.840 61.970 67.100 62.290 ;
        RECT 67.360 61.950 67.500 62.990 ;
        RECT 67.300 61.630 67.560 61.950 ;
        RECT 66.840 61.520 67.100 61.610 ;
        RECT 66.440 61.380 67.100 61.520 ;
        RECT 66.840 61.290 67.100 61.380 ;
        RECT 65.460 58.910 65.720 59.230 ;
        RECT 60.400 58.570 60.660 58.890 ;
        RECT 64.540 58.230 64.800 58.550 ;
        RECT 60.400 57.550 60.660 57.870 ;
        RECT 60.460 55.830 60.600 57.550 ;
        RECT 55.800 55.510 56.060 55.830 ;
        RECT 59.020 55.510 59.280 55.830 ;
        RECT 60.400 55.510 60.660 55.830 ;
        RECT 54.880 53.810 55.140 54.130 ;
        RECT 55.340 53.810 55.600 54.130 ;
        RECT 53.960 52.450 54.220 52.770 ;
        RECT 54.020 50.730 54.160 52.450 ;
        RECT 53.960 50.410 54.220 50.730 ;
        RECT 54.020 45.290 54.160 50.410 ;
        RECT 55.860 49.710 56.000 55.510 ;
        RECT 58.560 52.450 58.820 52.770 ;
        RECT 58.620 51.410 58.760 52.450 ;
        RECT 58.560 51.090 58.820 51.410 ;
        RECT 59.080 50.050 59.220 55.510 ;
        RECT 60.460 54.130 60.600 55.510 ;
        RECT 60.860 54.830 61.120 55.150 ;
        RECT 60.400 53.810 60.660 54.130 ;
        RECT 60.920 51.410 61.060 54.830 ;
        RECT 64.600 54.130 64.740 58.230 ;
        RECT 64.540 53.810 64.800 54.130 ;
        RECT 61.320 52.790 61.580 53.110 ;
        RECT 61.380 51.410 61.520 52.790 ;
        RECT 62.240 52.110 62.500 52.430 ;
        RECT 60.860 51.090 61.120 51.410 ;
        RECT 61.320 51.090 61.580 51.410 ;
        RECT 60.860 50.070 61.120 50.390 ;
        RECT 59.020 49.730 59.280 50.050 ;
        RECT 55.800 49.390 56.060 49.710 ;
        RECT 55.800 47.690 56.060 48.010 ;
        RECT 55.860 45.630 56.000 47.690 ;
        RECT 56.260 47.010 56.520 47.330 ;
        RECT 55.800 45.310 56.060 45.630 ;
        RECT 53.960 44.970 54.220 45.290 ;
        RECT 55.340 41.570 55.600 41.890 ;
        RECT 54.420 41.230 54.680 41.550 ;
        RECT 54.480 40.190 54.620 41.230 ;
        RECT 54.880 40.210 55.140 40.530 ;
        RECT 54.420 39.870 54.680 40.190 ;
        RECT 54.940 34.410 55.080 40.210 ;
        RECT 55.400 37.810 55.540 41.570 ;
        RECT 56.320 41.550 56.460 47.010 ;
        RECT 57.180 46.670 57.440 46.990 ;
        RECT 56.720 44.970 56.980 45.290 ;
        RECT 56.780 42.230 56.920 44.970 ;
        RECT 57.240 44.610 57.380 46.670 ;
        RECT 60.400 44.630 60.660 44.950 ;
        RECT 57.180 44.290 57.440 44.610 ;
        RECT 56.720 41.910 56.980 42.230 ;
        RECT 56.260 41.230 56.520 41.550 ;
        RECT 57.240 39.850 57.380 44.290 ;
        RECT 58.560 41.570 58.820 41.890 ;
        RECT 57.180 39.530 57.440 39.850 ;
        RECT 58.620 39.510 58.760 41.570 ;
        RECT 58.560 39.190 58.820 39.510 ;
        RECT 55.340 37.490 55.600 37.810 ;
        RECT 58.100 35.790 58.360 36.110 ;
        RECT 55.800 34.430 56.060 34.750 ;
        RECT 54.880 34.090 55.140 34.410 ;
        RECT 55.860 31.350 56.000 34.430 ;
        RECT 57.180 34.090 57.440 34.410 ;
        RECT 57.240 32.370 57.380 34.090 ;
        RECT 57.180 32.050 57.440 32.370 ;
        RECT 53.960 31.030 54.220 31.350 ;
        RECT 55.800 31.030 56.060 31.350 ;
        RECT 54.020 28.970 54.160 31.030 ;
        RECT 53.960 28.650 54.220 28.970 ;
        RECT 55.860 28.370 56.000 31.030 ;
        RECT 57.640 30.690 57.900 31.010 ;
        RECT 54.020 28.230 56.000 28.370 ;
        RECT 56.260 28.310 56.520 28.630 ;
        RECT 54.020 25.910 54.160 28.230 ;
        RECT 55.800 27.690 56.060 27.950 ;
        RECT 55.400 27.630 56.060 27.690 ;
        RECT 55.400 27.550 56.000 27.630 ;
        RECT 53.960 25.590 54.220 25.910 ;
        RECT 55.400 25.230 55.540 27.550 ;
        RECT 56.320 27.010 56.460 28.310 ;
        RECT 55.860 26.870 56.460 27.010 ;
        RECT 55.860 25.230 56.000 26.870 ;
        RECT 56.260 25.250 56.520 25.570 ;
        RECT 55.340 24.910 55.600 25.230 ;
        RECT 55.800 24.910 56.060 25.230 ;
        RECT 53.500 16.750 53.760 17.070 ;
        RECT 50.740 15.730 51.000 16.050 ;
        RECT 55.400 15.370 55.540 24.910 ;
        RECT 55.860 23.870 56.000 24.910 ;
        RECT 56.320 24.210 56.460 25.250 ;
        RECT 56.260 23.890 56.520 24.210 ;
        RECT 55.800 23.550 56.060 23.870 ;
        RECT 55.860 20.470 56.000 23.550 ;
        RECT 56.720 22.870 56.980 23.190 ;
        RECT 56.260 22.530 56.520 22.850 ;
        RECT 56.320 20.470 56.460 22.530 ;
        RECT 56.780 20.470 56.920 22.870 ;
        RECT 55.800 20.150 56.060 20.470 ;
        RECT 56.260 20.150 56.520 20.470 ;
        RECT 56.720 20.150 56.980 20.470 ;
        RECT 57.180 20.150 57.440 20.470 ;
        RECT 55.800 19.470 56.060 19.790 ;
        RECT 55.860 18.090 56.000 19.470 ;
        RECT 57.240 18.770 57.380 20.150 ;
        RECT 57.180 18.450 57.440 18.770 ;
        RECT 55.800 17.770 56.060 18.090 ;
        RECT 55.340 15.050 55.600 15.370 ;
        RECT 57.700 15.030 57.840 30.690 ;
        RECT 58.160 23.530 58.300 35.790 ;
        RECT 58.620 33.390 58.760 39.190 ;
        RECT 60.460 38.830 60.600 44.630 ;
        RECT 60.920 39.170 61.060 50.070 ;
        RECT 62.300 48.690 62.440 52.110 ;
        RECT 62.240 48.370 62.500 48.690 ;
        RECT 63.160 48.370 63.420 48.690 ;
        RECT 63.220 47.670 63.360 48.370 ;
        RECT 63.160 47.350 63.420 47.670 ;
        RECT 65.000 47.350 65.260 47.670 ;
        RECT 62.700 47.010 62.960 47.330 ;
        RECT 62.760 45.290 62.900 47.010 ;
        RECT 61.320 44.970 61.580 45.290 ;
        RECT 62.700 44.970 62.960 45.290 ;
        RECT 61.380 43.250 61.520 44.970 ;
        RECT 61.320 42.930 61.580 43.250 ;
        RECT 61.380 39.510 61.520 42.930 ;
        RECT 62.240 41.230 62.500 41.550 ;
        RECT 62.300 39.850 62.440 41.230 ;
        RECT 62.760 39.850 62.900 44.970 ;
        RECT 64.540 40.210 64.800 40.530 ;
        RECT 62.240 39.530 62.500 39.850 ;
        RECT 62.700 39.530 62.960 39.850 ;
        RECT 61.320 39.190 61.580 39.510 ;
        RECT 60.860 38.850 61.120 39.170 ;
        RECT 60.400 38.510 60.660 38.830 ;
        RECT 58.560 33.070 58.820 33.390 ;
        RECT 59.020 33.070 59.280 33.390 ;
        RECT 58.620 31.690 58.760 33.070 ;
        RECT 58.560 31.370 58.820 31.690 ;
        RECT 58.620 29.310 58.760 31.370 ;
        RECT 59.080 31.010 59.220 33.070 ;
        RECT 59.020 30.690 59.280 31.010 ;
        RECT 59.940 30.690 60.200 31.010 ;
        RECT 58.560 28.990 58.820 29.310 ;
        RECT 58.100 23.210 58.360 23.530 ;
        RECT 58.160 21.490 58.300 23.210 ;
        RECT 58.100 21.170 58.360 21.490 ;
        RECT 58.160 19.790 58.300 21.170 ;
        RECT 58.620 20.470 58.760 28.990 ;
        RECT 60.000 28.290 60.140 30.690 ;
        RECT 60.460 30.670 60.600 38.510 ;
        RECT 62.300 37.130 62.440 39.530 ;
        RECT 62.240 36.810 62.500 37.130 ;
        RECT 60.400 30.350 60.660 30.670 ;
        RECT 60.460 28.880 60.600 30.350 ;
        RECT 60.860 28.880 61.120 28.970 ;
        RECT 60.460 28.740 61.120 28.880 ;
        RECT 60.860 28.650 61.120 28.740 ;
        RECT 59.940 27.970 60.200 28.290 ;
        RECT 60.920 23.530 61.060 28.650 ;
        RECT 62.760 28.290 62.900 39.530 ;
        RECT 63.160 38.510 63.420 38.830 ;
        RECT 63.220 31.350 63.360 38.510 ;
        RECT 63.620 36.130 63.880 36.450 ;
        RECT 63.680 35.090 63.820 36.130 ;
        RECT 64.080 35.790 64.340 36.110 ;
        RECT 63.620 34.770 63.880 35.090 ;
        RECT 64.140 34.410 64.280 35.790 ;
        RECT 64.080 34.090 64.340 34.410 ;
        RECT 63.160 31.030 63.420 31.350 ;
        RECT 64.080 31.030 64.340 31.350 ;
        RECT 63.160 30.350 63.420 30.670 ;
        RECT 63.220 28.970 63.360 30.350 ;
        RECT 64.140 28.970 64.280 31.030 ;
        RECT 64.600 29.650 64.740 40.210 ;
        RECT 65.060 33.390 65.200 47.350 ;
        RECT 65.520 42.650 65.660 58.910 ;
        RECT 65.980 55.830 66.120 61.290 ;
        RECT 66.900 59.570 67.040 61.290 ;
        RECT 67.820 61.010 67.960 63.330 ;
        RECT 68.740 61.610 68.880 66.730 ;
        RECT 69.660 66.710 69.800 81.950 ;
        RECT 70.050 81.835 70.330 81.950 ;
        RECT 71.040 80.730 71.180 90.620 ;
        RECT 72.420 89.490 72.560 95.970 ;
        RECT 72.880 94.250 73.020 96.310 ;
        RECT 72.820 93.930 73.080 94.250 ;
        RECT 72.880 92.210 73.020 93.930 ;
        RECT 73.340 93.910 73.480 98.835 ;
        RECT 73.280 93.590 73.540 93.910 ;
        RECT 72.820 91.890 73.080 92.210 ;
        RECT 72.820 90.870 73.080 91.190 ;
        RECT 72.360 89.400 72.620 89.490 ;
        RECT 71.960 89.260 72.620 89.400 ;
        RECT 71.440 83.730 71.700 84.050 ;
        RECT 70.580 80.590 71.180 80.730 ;
        RECT 70.060 79.310 70.320 79.630 ;
        RECT 70.120 78.270 70.260 79.310 ;
        RECT 70.580 78.610 70.720 80.590 ;
        RECT 70.980 79.990 71.240 80.310 ;
        RECT 70.520 78.290 70.780 78.610 ;
        RECT 70.060 77.950 70.320 78.270 ;
        RECT 71.040 77.930 71.180 79.990 ;
        RECT 70.980 77.610 71.240 77.930 ;
        RECT 71.500 77.590 71.640 83.730 ;
        RECT 71.960 77.930 72.100 89.260 ;
        RECT 72.360 89.170 72.620 89.260 ;
        RECT 72.880 88.810 73.020 90.870 ;
        RECT 72.820 88.490 73.080 88.810 ;
        RECT 72.880 85.750 73.020 88.490 ;
        RECT 73.340 86.090 73.480 93.590 ;
        RECT 73.280 85.770 73.540 86.090 ;
        RECT 72.820 85.430 73.080 85.750 ;
        RECT 72.880 83.710 73.020 85.430 ;
        RECT 72.820 83.390 73.080 83.710 ;
        RECT 72.360 82.710 72.620 83.030 ;
        RECT 71.900 77.610 72.160 77.930 ;
        RECT 70.520 77.500 70.780 77.590 ;
        RECT 70.120 77.360 70.780 77.500 ;
        RECT 70.120 73.170 70.260 77.360 ;
        RECT 70.520 77.270 70.780 77.360 ;
        RECT 71.440 77.270 71.700 77.590 ;
        RECT 71.960 76.820 72.100 77.610 ;
        RECT 71.040 76.680 72.100 76.820 ;
        RECT 70.520 74.890 70.780 75.210 ;
        RECT 70.580 74.530 70.720 74.890 ;
        RECT 70.520 74.210 70.780 74.530 ;
        RECT 70.580 73.170 70.720 74.210 ;
        RECT 71.040 73.170 71.180 76.680 ;
        RECT 71.440 74.890 71.700 75.210 ;
        RECT 70.060 72.850 70.320 73.170 ;
        RECT 70.520 72.850 70.780 73.170 ;
        RECT 70.980 72.850 71.240 73.170 ;
        RECT 70.060 72.400 70.320 72.490 ;
        RECT 70.060 72.260 71.180 72.400 ;
        RECT 70.060 72.170 70.320 72.260 ;
        RECT 70.520 71.490 70.780 71.810 ;
        RECT 70.580 69.430 70.720 71.490 ;
        RECT 71.040 69.430 71.180 72.260 ;
        RECT 70.520 69.110 70.780 69.430 ;
        RECT 70.980 69.110 71.240 69.430 ;
        RECT 71.040 67.050 71.180 69.110 ;
        RECT 71.500 69.090 71.640 74.890 ;
        RECT 72.420 74.870 72.560 82.710 ;
        RECT 72.820 82.205 73.080 82.350 ;
        RECT 72.810 81.835 73.090 82.205 ;
        RECT 73.800 80.990 73.940 103.790 ;
        RECT 75.120 102.090 75.380 102.410 ;
        RECT 74.660 101.410 74.920 101.730 ;
        RECT 74.720 100.370 74.860 101.410 ;
        RECT 75.180 101.390 75.320 102.090 ;
        RECT 75.120 101.070 75.380 101.390 ;
        RECT 74.660 100.050 74.920 100.370 ;
        RECT 74.200 99.370 74.460 99.690 ;
        RECT 74.260 97.310 74.400 99.370 ;
        RECT 74.660 99.030 74.920 99.350 ;
        RECT 74.720 97.650 74.860 99.030 ;
        RECT 75.180 97.650 75.320 101.070 ;
        RECT 75.640 99.690 75.780 107.870 ;
        RECT 78.860 107.510 79.000 109.570 ;
        RECT 78.800 107.190 79.060 107.510 ;
        RECT 76.960 106.510 77.220 106.830 ;
        RECT 76.040 105.490 76.300 105.810 ;
        RECT 76.100 99.690 76.240 105.490 ;
        RECT 77.020 105.130 77.160 106.510 ;
        RECT 76.500 104.810 76.760 105.130 ;
        RECT 76.960 104.810 77.220 105.130 ;
        RECT 76.560 100.370 76.700 104.810 ;
        RECT 76.960 103.790 77.220 104.110 ;
        RECT 77.020 102.410 77.160 103.790 ;
        RECT 77.420 102.430 77.680 102.750 ;
        RECT 76.960 102.090 77.220 102.410 ;
        RECT 76.500 100.050 76.760 100.370 ;
        RECT 75.580 99.370 75.840 99.690 ;
        RECT 76.040 99.370 76.300 99.690 ;
        RECT 75.580 98.690 75.840 99.010 ;
        RECT 76.500 98.690 76.760 99.010 ;
        RECT 74.660 97.330 74.920 97.650 ;
        RECT 75.120 97.330 75.380 97.650 ;
        RECT 74.200 96.990 74.460 97.310 ;
        RECT 74.260 88.470 74.400 96.990 ;
        RECT 74.660 96.310 74.920 96.630 ;
        RECT 74.720 89.490 74.860 96.310 ;
        RECT 75.640 95.125 75.780 98.690 ;
        RECT 76.560 95.950 76.700 98.690 ;
        RECT 76.500 95.630 76.760 95.950 ;
        RECT 75.570 94.755 75.850 95.125 ;
        RECT 74.660 89.170 74.920 89.490 ;
        RECT 74.200 88.150 74.460 88.470 ;
        RECT 74.200 87.470 74.460 87.790 ;
        RECT 74.260 84.050 74.400 87.470 ;
        RECT 74.720 85.750 74.860 89.170 ;
        RECT 75.120 88.150 75.380 88.470 ;
        RECT 74.660 85.430 74.920 85.750 ;
        RECT 74.200 83.730 74.460 84.050 ;
        RECT 74.660 82.370 74.920 82.690 ;
        RECT 73.740 80.670 74.000 80.990 ;
        RECT 73.800 80.310 73.940 80.670 ;
        RECT 73.740 79.990 74.000 80.310 ;
        RECT 73.280 78.290 73.540 78.610 ;
        RECT 73.730 78.435 74.010 78.805 ;
        RECT 72.820 75.570 73.080 75.890 ;
        RECT 72.360 74.780 72.620 74.870 ;
        RECT 71.960 74.640 72.620 74.780 ;
        RECT 71.440 68.770 71.700 69.090 ;
        RECT 70.980 66.730 71.240 67.050 ;
        RECT 69.600 66.390 69.860 66.710 ;
        RECT 71.960 66.370 72.100 74.640 ;
        RECT 72.360 74.550 72.620 74.640 ;
        RECT 72.350 71.635 72.630 72.005 ;
        RECT 72.420 71.470 72.560 71.635 ;
        RECT 72.360 71.150 72.620 71.470 ;
        RECT 72.360 69.790 72.620 70.110 ;
        RECT 72.420 67.050 72.560 69.790 ;
        RECT 72.360 66.730 72.620 67.050 ;
        RECT 71.900 66.050 72.160 66.370 ;
        RECT 70.520 64.010 70.780 64.330 ;
        RECT 68.680 61.290 68.940 61.610 ;
        RECT 67.360 60.870 67.960 61.010 ;
        RECT 66.840 59.250 67.100 59.570 ;
        RECT 66.900 58.550 67.040 59.250 ;
        RECT 66.840 58.230 67.100 58.550 ;
        RECT 66.380 57.550 66.640 57.870 ;
        RECT 65.920 55.510 66.180 55.830 ;
        RECT 66.440 53.110 66.580 57.550 ;
        RECT 66.380 52.790 66.640 53.110 ;
        RECT 66.380 47.010 66.640 47.330 ;
        RECT 66.440 45.290 66.580 47.010 ;
        RECT 67.360 45.630 67.500 60.870 ;
        RECT 67.750 60.075 68.030 60.445 ;
        RECT 70.060 60.270 70.320 60.590 ;
        RECT 67.820 58.890 67.960 60.075 ;
        RECT 67.760 58.570 68.020 58.890 ;
        RECT 68.680 58.230 68.940 58.550 ;
        RECT 69.140 58.290 69.400 58.550 ;
        RECT 70.120 58.290 70.260 60.270 ;
        RECT 70.580 58.550 70.720 64.010 ;
        RECT 70.980 61.970 71.240 62.290 ;
        RECT 71.040 58.550 71.180 61.970 ;
        RECT 69.140 58.230 70.260 58.290 ;
        RECT 70.520 58.230 70.780 58.550 ;
        RECT 70.980 58.230 71.240 58.550 ;
        RECT 71.440 58.230 71.700 58.550 ;
        RECT 67.760 57.890 68.020 58.210 ;
        RECT 67.820 55.490 67.960 57.890 ;
        RECT 68.740 56.850 68.880 58.230 ;
        RECT 69.200 58.150 70.260 58.230 ;
        RECT 69.140 57.550 69.400 57.870 ;
        RECT 68.680 56.530 68.940 56.850 ;
        RECT 69.200 56.170 69.340 57.550 ;
        RECT 69.140 55.850 69.400 56.170 ;
        RECT 67.760 55.170 68.020 55.490 ;
        RECT 70.120 55.150 70.260 58.150 ;
        RECT 71.500 57.870 71.640 58.230 ;
        RECT 70.980 57.550 71.240 57.870 ;
        RECT 71.440 57.550 71.700 57.870 ;
        RECT 71.040 55.830 71.180 57.550 ;
        RECT 71.440 56.190 71.700 56.510 ;
        RECT 70.980 55.510 71.240 55.830 ;
        RECT 70.060 54.830 70.320 55.150 ;
        RECT 71.500 52.770 71.640 56.190 ;
        RECT 71.960 56.170 72.100 66.050 ;
        RECT 72.880 66.030 73.020 75.570 ;
        RECT 73.340 75.210 73.480 78.290 ;
        RECT 73.800 78.270 73.940 78.435 ;
        RECT 73.740 77.950 74.000 78.270 ;
        RECT 74.200 77.610 74.460 77.930 ;
        RECT 74.260 77.250 74.400 77.610 ;
        RECT 74.200 76.930 74.460 77.250 ;
        RECT 73.280 74.890 73.540 75.210 ;
        RECT 74.720 74.870 74.860 82.370 ;
        RECT 75.180 74.870 75.320 88.150 ;
        RECT 75.640 87.790 75.780 94.755 ;
        RECT 76.560 94.250 76.700 95.630 ;
        RECT 76.500 93.930 76.760 94.250 ;
        RECT 77.020 93.910 77.160 102.090 ;
        RECT 77.480 99.010 77.620 102.430 ;
        RECT 79.320 99.600 79.460 114.670 ;
        RECT 88.520 113.970 88.660 115.690 ;
        RECT 89.830 115.155 90.110 115.525 ;
        RECT 89.840 115.010 90.100 115.155 ;
        RECT 88.460 113.650 88.720 113.970 ;
        RECT 79.720 112.630 79.980 112.950 ;
        RECT 87.540 112.630 87.800 112.950 ;
        RECT 88.460 112.630 88.720 112.950 ;
        RECT 79.780 110.570 79.920 112.630 ;
        RECT 79.720 110.250 79.980 110.570 ;
        RECT 81.100 110.250 81.360 110.570 ;
        RECT 81.160 108.530 81.300 110.250 ;
        RECT 87.600 110.230 87.740 112.630 ;
        RECT 87.540 109.910 87.800 110.230 ;
        RECT 87.080 109.230 87.340 109.550 ;
        RECT 81.100 108.210 81.360 108.530 ;
        RECT 84.780 107.530 85.040 107.850 ;
        RECT 82.940 106.510 83.200 106.830 ;
        RECT 80.180 104.130 80.440 104.450 ;
        RECT 79.720 99.600 79.980 99.690 ;
        RECT 78.860 99.460 79.980 99.600 ;
        RECT 78.340 99.030 78.600 99.350 ;
        RECT 77.420 98.690 77.680 99.010 ;
        RECT 77.880 98.350 78.140 98.670 ;
        RECT 77.940 97.310 78.080 98.350 ;
        RECT 78.400 97.650 78.540 99.030 ;
        RECT 78.340 97.330 78.600 97.650 ;
        RECT 77.880 96.990 78.140 97.310 ;
        RECT 77.880 93.930 78.140 94.250 ;
        RECT 76.960 93.590 77.220 93.910 ;
        RECT 77.940 93.570 78.080 93.930 ;
        RECT 77.880 93.250 78.140 93.570 ;
        RECT 77.940 90.510 78.080 93.250 ;
        RECT 78.860 93.230 79.000 99.460 ;
        RECT 79.720 99.370 79.980 99.460 ;
        RECT 79.250 98.835 79.530 99.205 ;
        RECT 79.320 98.670 79.460 98.835 ;
        RECT 79.260 98.350 79.520 98.670 ;
        RECT 80.240 96.970 80.380 104.130 ;
        RECT 80.640 101.750 80.900 102.070 ;
        RECT 80.180 96.650 80.440 96.970 ;
        RECT 80.180 93.930 80.440 94.250 ;
        RECT 79.260 93.590 79.520 93.910 ;
        RECT 78.800 92.910 79.060 93.230 ;
        RECT 78.860 91.190 79.000 92.910 ;
        RECT 79.320 91.190 79.460 93.590 ;
        RECT 80.240 91.530 80.380 93.930 ;
        RECT 80.180 91.210 80.440 91.530 ;
        RECT 78.800 90.870 79.060 91.190 ;
        RECT 79.260 90.870 79.520 91.190 ;
        RECT 77.880 90.190 78.140 90.510 ;
        RECT 75.580 87.470 75.840 87.790 ;
        RECT 75.580 86.450 75.840 86.770 ;
        RECT 75.640 80.730 75.780 86.450 ;
        RECT 77.940 86.430 78.080 90.190 ;
        RECT 79.320 89.400 79.460 90.870 ;
        RECT 79.320 89.260 79.920 89.400 ;
        RECT 78.800 88.830 79.060 89.150 ;
        RECT 77.880 86.110 78.140 86.430 ;
        RECT 76.960 85.770 77.220 86.090 ;
        RECT 76.500 85.090 76.760 85.410 ;
        RECT 76.040 84.750 76.300 85.070 ;
        RECT 76.100 82.350 76.240 84.750 ;
        RECT 76.040 82.030 76.300 82.350 ;
        RECT 75.640 80.590 76.240 80.730 ;
        RECT 76.100 80.310 76.240 80.590 ;
        RECT 75.580 79.990 75.840 80.310 ;
        RECT 76.040 79.990 76.300 80.310 ;
        RECT 75.640 78.805 75.780 79.990 ;
        RECT 75.570 78.435 75.850 78.805 ;
        RECT 75.580 76.930 75.840 77.250 ;
        RECT 74.660 74.550 74.920 74.870 ;
        RECT 75.120 74.550 75.380 74.870 ;
        RECT 73.280 74.210 73.540 74.530 ;
        RECT 73.340 69.430 73.480 74.210 ;
        RECT 73.740 73.870 74.000 74.190 ;
        RECT 74.200 73.870 74.460 74.190 ;
        RECT 73.800 73.170 73.940 73.870 ;
        RECT 73.740 72.850 74.000 73.170 ;
        RECT 73.740 72.170 74.000 72.490 ;
        RECT 73.800 70.450 73.940 72.170 ;
        RECT 74.260 72.150 74.400 73.870 ;
        RECT 74.200 71.830 74.460 72.150 ;
        RECT 73.740 70.130 74.000 70.450 ;
        RECT 74.200 69.790 74.460 70.110 ;
        RECT 73.280 69.110 73.540 69.430 ;
        RECT 73.740 68.770 74.000 69.090 ;
        RECT 73.800 67.050 73.940 68.770 ;
        RECT 73.740 66.730 74.000 67.050 ;
        RECT 72.820 65.710 73.080 66.030 ;
        RECT 72.880 63.990 73.020 65.710 ;
        RECT 73.800 64.330 73.940 66.730 ;
        RECT 73.740 64.010 74.000 64.330 ;
        RECT 72.820 63.670 73.080 63.990 ;
        RECT 72.880 60.445 73.020 63.670 ;
        RECT 73.800 61.270 73.940 64.010 ;
        RECT 73.740 60.950 74.000 61.270 ;
        RECT 72.810 60.075 73.090 60.445 ;
        RECT 73.740 60.270 74.000 60.590 ;
        RECT 72.360 59.250 72.620 59.570 ;
        RECT 72.820 59.250 73.080 59.570 ;
        RECT 72.420 58.550 72.560 59.250 ;
        RECT 72.880 58.550 73.020 59.250 ;
        RECT 73.280 58.910 73.540 59.230 ;
        RECT 72.360 58.230 72.620 58.550 ;
        RECT 72.820 58.230 73.080 58.550 ;
        RECT 72.420 56.850 72.560 58.230 ;
        RECT 73.340 58.210 73.480 58.910 ;
        RECT 73.800 58.550 73.940 60.270 ;
        RECT 74.260 58.890 74.400 69.790 ;
        RECT 74.720 61.950 74.860 74.550 ;
        RECT 75.640 74.190 75.780 76.930 ;
        RECT 75.580 74.100 75.840 74.190 ;
        RECT 75.180 73.960 75.840 74.100 ;
        RECT 75.180 72.685 75.320 73.960 ;
        RECT 75.580 73.870 75.840 73.960 ;
        RECT 76.100 73.250 76.240 79.990 ;
        RECT 76.560 75.890 76.700 85.090 ;
        RECT 77.020 83.710 77.160 85.770 ;
        RECT 77.420 85.090 77.680 85.410 ;
        RECT 76.960 83.390 77.220 83.710 ;
        RECT 76.960 80.730 77.220 80.990 ;
        RECT 77.480 80.730 77.620 85.090 ;
        RECT 76.960 80.670 77.620 80.730 ;
        RECT 77.020 80.590 77.620 80.670 ;
        RECT 76.500 75.570 76.760 75.890 ;
        RECT 76.960 74.890 77.220 75.210 ;
        RECT 77.020 73.930 77.160 74.890 ;
        RECT 75.640 73.110 76.240 73.250 ;
        RECT 76.560 73.790 77.160 73.930 ;
        RECT 75.110 72.315 75.390 72.685 ;
        RECT 75.180 69.770 75.320 72.315 ;
        RECT 75.640 71.470 75.780 73.110 ;
        RECT 76.040 72.570 76.300 72.830 ;
        RECT 76.560 72.570 76.700 73.790 ;
        RECT 76.960 72.850 77.220 73.170 ;
        RECT 76.040 72.510 76.700 72.570 ;
        RECT 76.100 72.430 76.700 72.510 ;
        RECT 76.040 72.060 76.300 72.150 ;
        RECT 77.020 72.060 77.160 72.850 ;
        RECT 77.480 72.490 77.620 80.590 ;
        RECT 77.940 78.010 78.080 86.110 ;
        RECT 78.860 80.310 79.000 88.830 ;
        RECT 79.780 88.810 79.920 89.260 ;
        RECT 80.240 89.150 80.380 91.210 ;
        RECT 80.180 88.830 80.440 89.150 ;
        RECT 80.700 88.810 80.840 101.750 ;
        RECT 82.480 101.410 82.740 101.730 ;
        RECT 82.540 100.370 82.680 101.410 ;
        RECT 82.480 100.050 82.740 100.370 ;
        RECT 81.560 98.690 81.820 99.010 ;
        RECT 81.100 95.630 81.360 95.950 ;
        RECT 81.160 94.930 81.300 95.630 ;
        RECT 81.100 94.610 81.360 94.930 ;
        RECT 79.260 88.490 79.520 88.810 ;
        RECT 79.720 88.490 79.980 88.810 ;
        RECT 80.640 88.490 80.900 88.810 ;
        RECT 79.320 83.370 79.460 88.490 ;
        RECT 79.780 85.320 79.920 88.490 ;
        RECT 79.780 85.180 80.380 85.320 ;
        RECT 79.260 83.050 79.520 83.370 ;
        RECT 80.240 80.310 80.380 85.180 ;
        RECT 80.700 80.650 80.840 88.490 ;
        RECT 81.620 85.750 81.760 98.690 ;
        RECT 83.000 94.930 83.140 106.510 ;
        RECT 84.840 105.810 84.980 107.530 ;
        RECT 87.140 107.510 87.280 109.230 ;
        RECT 88.520 108.530 88.660 112.630 ;
        RECT 89.840 112.125 90.100 112.270 ;
        RECT 89.830 111.755 90.110 112.125 ;
        RECT 88.460 108.210 88.720 108.530 ;
        RECT 87.080 107.190 87.340 107.510 ;
        RECT 87.540 107.190 87.800 107.510 ;
        RECT 84.780 105.490 85.040 105.810 ;
        RECT 87.600 104.790 87.740 107.190 ;
        RECT 100.360 105.820 100.660 180.090 ;
        RECT 100.860 179.630 118.970 179.640 ;
        RECT 100.860 179.350 119.005 179.630 ;
        RECT 100.860 179.340 118.970 179.350 ;
        RECT 100.860 120.760 101.160 179.340 ;
        RECT 101.580 178.940 122.370 178.950 ;
        RECT 101.580 178.660 122.405 178.940 ;
        RECT 101.580 178.650 122.370 178.660 ;
        RECT 101.580 135.760 101.880 178.650 ;
        RECT 102.210 178.350 115.570 178.360 ;
        RECT 102.210 178.070 115.605 178.350 ;
        RECT 102.210 178.060 115.570 178.070 ;
        RECT 102.210 150.840 102.510 178.060 ;
        RECT 102.770 177.660 112.170 177.670 ;
        RECT 102.770 177.380 112.205 177.660 ;
        RECT 102.770 177.370 112.170 177.380 ;
        RECT 102.790 165.570 103.090 177.370 ;
        RECT 106.840 176.770 107.540 176.780 ;
        RECT 106.500 176.030 107.850 176.770 ;
        RECT 106.840 166.600 107.540 176.030 ;
        RECT 117.980 174.620 118.880 176.640 ;
        RECT 116.255 172.705 116.575 172.760 ;
        RECT 116.255 172.550 118.860 172.705 ;
        RECT 116.255 172.500 116.575 172.550 ;
        RECT 108.890 171.080 116.880 171.470 ;
        RECT 108.820 168.770 109.400 169.400 ;
        RECT 111.430 168.020 114.090 171.080 ;
        RECT 108.930 167.570 116.870 168.020 ;
        RECT 106.750 165.810 107.610 166.600 ;
        RECT 106.840 161.770 107.540 161.780 ;
        RECT 106.500 161.030 107.850 161.770 ;
        RECT 106.840 151.600 107.540 161.030 ;
        RECT 116.160 157.690 116.480 157.750 ;
        RECT 116.160 157.550 118.510 157.690 ;
        RECT 116.160 157.490 116.480 157.550 ;
        RECT 108.890 156.080 116.880 156.470 ;
        RECT 108.790 153.690 109.370 154.320 ;
        RECT 111.430 153.020 114.090 156.080 ;
        RECT 108.930 152.570 116.870 153.020 ;
        RECT 102.210 150.540 103.050 150.840 ;
        RECT 106.750 150.810 107.610 151.600 ;
        RECT 106.840 146.720 107.540 146.730 ;
        RECT 106.500 145.980 107.850 146.720 ;
        RECT 106.840 136.550 107.540 145.980 ;
        RECT 116.400 142.635 116.720 142.690 ;
        RECT 116.400 142.485 118.115 142.635 ;
        RECT 116.400 142.430 116.720 142.485 ;
        RECT 108.890 141.030 116.880 141.420 ;
        RECT 108.790 138.740 109.370 139.370 ;
        RECT 111.430 137.970 114.090 141.030 ;
        RECT 108.930 137.520 116.870 137.970 ;
        RECT 106.750 135.760 107.610 136.550 ;
        RECT 101.580 135.460 103.130 135.760 ;
        RECT 106.840 131.720 107.540 131.730 ;
        RECT 106.500 130.980 107.850 131.720 ;
        RECT 106.840 121.550 107.540 130.980 ;
        RECT 116.290 127.640 116.610 127.680 ;
        RECT 116.290 127.460 117.690 127.640 ;
        RECT 116.290 127.420 116.610 127.460 ;
        RECT 108.890 126.030 116.880 126.420 ;
        RECT 108.790 123.740 109.370 124.370 ;
        RECT 111.430 122.970 114.090 126.030 ;
        RECT 108.930 122.520 116.870 122.970 ;
        RECT 106.750 120.760 107.610 121.550 ;
        RECT 100.860 120.460 103.170 120.760 ;
        RECT 106.790 116.780 107.490 116.790 ;
        RECT 106.450 116.040 107.800 116.780 ;
        RECT 106.790 106.610 107.490 116.040 ;
        RECT 116.510 112.675 116.830 112.720 ;
        RECT 116.510 112.505 117.195 112.675 ;
        RECT 116.510 112.460 116.830 112.505 ;
        RECT 108.840 111.090 116.830 111.480 ;
        RECT 108.750 108.700 109.330 109.330 ;
        RECT 111.380 108.030 114.040 111.090 ;
        RECT 108.880 107.580 116.820 108.030 ;
        RECT 106.700 105.820 107.560 106.610 ;
        RECT 100.360 105.520 103.080 105.820 ;
        RECT 87.540 104.470 87.800 104.790 ;
        RECT 84.320 103.790 84.580 104.110 ;
        RECT 84.380 100.370 84.520 103.790 ;
        RECT 87.600 103.090 87.740 104.470 ;
        RECT 100.180 103.665 112.290 103.900 ;
        RECT 100.180 103.175 110.620 103.390 ;
        RECT 87.540 102.770 87.800 103.090 ;
        RECT 100.180 102.760 109.045 102.970 ;
        RECT 100.180 102.210 107.455 102.480 ;
        RECT 100.180 101.665 105.905 101.930 ;
        RECT 85.240 101.070 85.500 101.390 ;
        RECT 100.180 101.075 104.305 101.360 ;
        RECT 84.320 100.050 84.580 100.370 ;
        RECT 85.300 99.350 85.440 101.070 ;
        RECT 100.180 100.400 102.800 100.700 ;
        RECT 100.180 99.790 101.275 100.035 ;
        RECT 84.780 99.030 85.040 99.350 ;
        RECT 85.240 99.030 85.500 99.350 ;
        RECT 84.840 97.650 84.980 99.030 ;
        RECT 84.780 97.330 85.040 97.650 ;
        RECT 82.940 94.610 83.200 94.930 ;
        RECT 101.030 92.875 101.275 99.790 ;
        RECT 102.500 92.925 102.800 100.400 ;
        RECT 104.020 92.925 104.305 101.075 ;
        RECT 105.640 92.955 105.905 101.665 ;
        RECT 100.620 92.615 101.680 92.875 ;
        RECT 102.120 92.625 103.180 92.925 ;
        RECT 103.630 92.640 104.690 92.925 ;
        RECT 105.240 92.690 106.300 92.955 ;
        RECT 107.185 92.925 107.455 102.210 ;
        RECT 108.835 92.955 109.045 102.760 ;
        RECT 106.790 92.655 107.850 92.925 ;
        RECT 108.410 92.695 109.470 92.955 ;
        RECT 110.405 92.925 110.620 103.175 ;
        RECT 112.055 92.945 112.290 103.665 ;
        RECT 117.025 101.605 117.195 112.505 ;
        RECT 117.510 102.010 117.690 127.460 ;
        RECT 117.965 102.335 118.115 142.485 ;
        RECT 118.370 102.640 118.510 157.550 ;
        RECT 118.705 102.965 118.860 172.550 ;
        RECT 123.240 169.890 123.540 180.190 ;
        RECT 120.480 169.590 123.540 169.890 ;
        RECT 123.830 179.710 129.170 179.720 ;
        RECT 123.830 179.430 129.205 179.710 ;
        RECT 152.680 179.480 152.960 179.515 ;
        RECT 123.830 179.420 129.170 179.430 ;
        RECT 120.480 105.740 120.780 169.590 ;
        RECT 123.830 168.770 124.130 179.420 ;
        RECT 143.320 179.180 152.970 179.480 ;
        RECT 121.150 168.470 124.130 168.770 ;
        RECT 124.430 179.000 132.570 179.010 ;
        RECT 124.430 178.720 132.605 179.000 ;
        RECT 124.430 178.710 132.570 178.720 ;
        RECT 121.150 120.900 121.450 168.470 ;
        RECT 124.430 167.820 124.730 178.710 ;
        RECT 121.750 167.520 124.730 167.820 ;
        RECT 124.920 178.280 135.970 178.290 ;
        RECT 124.920 178.000 136.005 178.280 ;
        RECT 124.920 177.990 135.970 178.000 ;
        RECT 121.750 135.710 122.050 167.520 ;
        RECT 124.920 166.810 125.220 177.990 ;
        RECT 122.310 166.510 125.220 166.810 ;
        RECT 125.540 177.560 142.770 177.570 ;
        RECT 125.540 177.280 142.805 177.560 ;
        RECT 125.540 177.270 142.770 177.280 ;
        RECT 122.310 150.820 122.610 166.510 ;
        RECT 125.540 166.000 125.840 177.270 ;
        RECT 126.720 176.720 127.420 176.730 ;
        RECT 126.380 175.980 127.730 176.720 ;
        RECT 126.720 166.550 127.420 175.980 ;
        RECT 137.800 174.600 138.700 176.620 ;
        RECT 136.460 172.635 136.780 172.690 ;
        RECT 136.460 172.485 138.465 172.635 ;
        RECT 136.460 172.430 136.780 172.485 ;
        RECT 128.770 171.030 136.760 171.420 ;
        RECT 128.680 168.760 129.260 169.390 ;
        RECT 131.310 167.970 133.970 171.030 ;
        RECT 128.810 167.520 136.750 167.970 ;
        RECT 122.900 165.700 125.840 166.000 ;
        RECT 126.630 165.760 127.490 166.550 ;
        RECT 126.720 161.770 127.420 161.780 ;
        RECT 126.380 161.030 127.730 161.770 ;
        RECT 126.720 151.600 127.420 161.030 ;
        RECT 136.270 157.695 136.590 157.720 ;
        RECT 136.270 157.485 138.095 157.695 ;
        RECT 136.270 157.460 136.590 157.485 ;
        RECT 128.770 156.080 136.760 156.470 ;
        RECT 128.680 153.800 129.260 154.430 ;
        RECT 131.310 153.020 133.970 156.080 ;
        RECT 128.810 152.570 136.750 153.020 ;
        RECT 122.310 150.520 122.980 150.820 ;
        RECT 126.630 150.810 127.490 151.600 ;
        RECT 126.720 146.720 127.420 146.730 ;
        RECT 126.380 145.980 127.730 146.720 ;
        RECT 126.720 136.550 127.420 145.980 ;
        RECT 136.150 142.705 136.470 142.750 ;
        RECT 136.150 142.535 137.715 142.705 ;
        RECT 136.150 142.490 136.470 142.535 ;
        RECT 128.770 141.030 136.760 141.420 ;
        RECT 128.680 138.730 129.260 139.360 ;
        RECT 131.310 137.970 133.970 141.030 ;
        RECT 128.810 137.520 136.750 137.970 ;
        RECT 126.630 135.760 127.490 136.550 ;
        RECT 121.750 135.410 122.980 135.710 ;
        RECT 126.720 131.780 127.420 131.790 ;
        RECT 126.380 131.040 127.730 131.780 ;
        RECT 126.720 121.610 127.420 131.040 ;
        RECT 136.335 127.700 136.655 127.760 ;
        RECT 136.335 127.555 137.375 127.700 ;
        RECT 136.335 127.500 136.655 127.555 ;
        RECT 128.770 126.090 136.760 126.480 ;
        RECT 128.610 123.790 129.190 124.420 ;
        RECT 131.310 123.030 133.970 126.090 ;
        RECT 128.810 122.580 136.750 123.030 ;
        RECT 121.150 120.600 123.010 120.900 ;
        RECT 126.630 120.820 127.490 121.610 ;
        RECT 126.720 116.780 127.420 116.790 ;
        RECT 126.380 116.040 127.730 116.780 ;
        RECT 126.720 106.610 127.420 116.040 ;
        RECT 136.160 112.690 136.480 112.750 ;
        RECT 136.160 112.550 137.090 112.690 ;
        RECT 136.160 112.490 136.480 112.550 ;
        RECT 128.770 111.090 136.760 111.480 ;
        RECT 128.730 108.760 129.310 109.390 ;
        RECT 131.310 108.030 133.970 111.090 ;
        RECT 128.810 107.580 136.750 108.030 ;
        RECT 126.630 105.820 127.490 106.610 ;
        RECT 120.480 105.440 123.040 105.740 ;
        RECT 136.950 103.450 137.090 112.550 ;
        RECT 137.230 103.740 137.375 127.555 ;
        RECT 137.545 104.065 137.715 142.535 ;
        RECT 137.885 104.455 138.095 157.485 ;
        RECT 138.315 104.825 138.465 172.485 ;
        RECT 143.320 169.390 143.620 179.180 ;
        RECT 152.680 179.145 152.960 179.180 ;
        RECT 140.280 169.090 143.620 169.390 ;
        RECT 144.050 178.740 146.170 178.750 ;
        RECT 144.050 178.460 146.205 178.740 ;
        RECT 144.050 178.450 146.170 178.460 ;
        RECT 140.280 105.820 140.580 169.090 ;
        RECT 144.050 168.490 144.350 178.450 ;
        RECT 145.290 178.030 149.570 178.040 ;
        RECT 145.290 177.750 149.605 178.030 ;
        RECT 145.290 177.740 149.570 177.750 ;
        RECT 144.680 176.850 144.960 176.885 ;
        RECT 140.940 168.190 144.350 168.490 ;
        RECT 140.940 120.830 141.240 168.190 ;
        RECT 144.670 167.700 144.970 176.850 ;
        RECT 141.710 167.400 144.970 167.700 ;
        RECT 141.710 135.850 142.010 167.400 ;
        RECT 145.290 166.930 145.590 177.740 ;
        RECT 142.350 166.630 145.590 166.930 ;
        RECT 145.960 177.370 148.420 177.380 ;
        RECT 145.960 177.090 148.455 177.370 ;
        RECT 145.960 177.080 148.420 177.090 ;
        RECT 142.350 150.730 142.650 166.630 ;
        RECT 145.960 166.020 146.260 177.080 ;
        RECT 146.750 176.770 147.450 176.780 ;
        RECT 146.410 176.030 147.760 176.770 ;
        RECT 146.750 166.600 147.450 176.030 ;
        RECT 157.570 174.580 158.470 176.600 ;
        RECT 156.415 172.650 156.735 172.710 ;
        RECT 156.415 172.505 158.350 172.650 ;
        RECT 156.415 172.450 156.735 172.505 ;
        RECT 148.800 171.080 156.790 171.470 ;
        RECT 148.880 168.740 149.460 169.370 ;
        RECT 151.340 168.020 154.000 171.080 ;
        RECT 148.840 167.570 156.780 168.020 ;
        RECT 142.960 165.720 146.260 166.020 ;
        RECT 146.660 165.810 147.520 166.600 ;
        RECT 146.800 161.720 147.500 161.730 ;
        RECT 146.460 160.980 147.810 161.720 ;
        RECT 146.800 151.550 147.500 160.980 ;
        RECT 156.500 157.640 156.820 157.700 ;
        RECT 156.500 157.500 158.030 157.640 ;
        RECT 156.500 157.440 156.820 157.500 ;
        RECT 148.850 156.030 156.840 156.420 ;
        RECT 148.920 153.710 149.500 154.340 ;
        RECT 151.390 152.970 154.050 156.030 ;
        RECT 148.890 152.520 156.830 152.970 ;
        RECT 146.710 150.760 147.570 151.550 ;
        RECT 142.350 150.430 142.970 150.730 ;
        RECT 146.750 146.720 147.450 146.730 ;
        RECT 146.410 145.980 147.760 146.720 ;
        RECT 146.750 136.550 147.450 145.980 ;
        RECT 156.330 142.625 156.590 142.710 ;
        RECT 156.330 142.475 157.705 142.625 ;
        RECT 156.330 142.390 156.590 142.475 ;
        RECT 148.800 141.030 156.790 141.420 ;
        RECT 148.830 138.670 149.410 139.300 ;
        RECT 151.340 137.970 154.000 141.030 ;
        RECT 148.840 137.520 156.780 137.970 ;
        RECT 141.710 135.550 143.010 135.850 ;
        RECT 146.660 135.760 147.520 136.550 ;
        RECT 146.750 131.780 147.450 131.790 ;
        RECT 146.410 131.040 147.760 131.780 ;
        RECT 146.750 121.610 147.450 131.040 ;
        RECT 156.410 127.660 156.730 127.720 ;
        RECT 156.410 127.520 157.410 127.660 ;
        RECT 156.410 127.460 156.730 127.520 ;
        RECT 148.800 126.090 156.790 126.480 ;
        RECT 148.950 123.750 149.530 124.380 ;
        RECT 151.340 123.030 154.000 126.090 ;
        RECT 148.840 122.580 156.780 123.030 ;
        RECT 140.940 120.530 142.990 120.830 ;
        RECT 146.660 120.820 147.520 121.610 ;
        RECT 146.750 116.780 147.450 116.790 ;
        RECT 146.410 116.040 147.760 116.780 ;
        RECT 146.750 106.610 147.450 116.040 ;
        RECT 156.000 112.715 156.320 112.770 ;
        RECT 156.000 112.565 157.115 112.715 ;
        RECT 156.000 112.510 156.320 112.565 ;
        RECT 148.800 111.090 156.790 111.480 ;
        RECT 148.910 108.790 149.490 109.420 ;
        RECT 151.340 108.030 154.000 111.090 ;
        RECT 148.840 107.580 156.780 108.030 ;
        RECT 146.660 105.820 147.520 106.610 ;
        RECT 140.280 105.520 143.020 105.820 ;
        RECT 138.315 104.675 149.650 104.825 ;
        RECT 137.885 104.245 147.750 104.455 ;
        RECT 137.545 103.895 146.220 104.065 ;
        RECT 137.230 103.595 144.785 103.740 ;
        RECT 136.950 103.310 143.320 103.450 ;
        RECT 118.705 102.810 141.785 102.965 ;
        RECT 118.370 102.500 140.290 102.640 ;
        RECT 117.965 102.185 138.860 102.335 ;
        RECT 117.510 101.970 137.340 102.010 ;
        RECT 117.510 101.830 137.730 101.970 ;
        RECT 137.160 101.620 137.730 101.830 ;
        RECT 117.025 101.435 135.840 101.605 ;
        RECT 137.210 101.500 137.730 101.620 ;
        RECT 135.670 99.200 135.840 101.435 ;
        RECT 138.710 99.390 138.860 102.185 ;
        RECT 140.150 101.990 140.290 102.500 ;
        RECT 140.150 101.620 140.700 101.990 ;
        RECT 140.180 101.520 140.700 101.620 ;
        RECT 135.670 98.995 136.300 99.200 ;
        RECT 138.710 99.015 139.270 99.390 ;
        RECT 135.690 98.720 136.300 98.995 ;
        RECT 138.750 98.920 139.270 99.015 ;
        RECT 141.630 99.310 141.785 102.810 ;
        RECT 143.180 102.050 143.320 103.310 ;
        RECT 143.180 101.580 143.700 102.050 ;
        RECT 144.640 99.340 144.785 103.595 ;
        RECT 146.050 102.080 146.220 103.895 ;
        RECT 146.050 101.950 146.610 102.080 ;
        RECT 146.090 101.610 146.610 101.950 ;
        RECT 147.540 99.390 147.750 104.245 ;
        RECT 149.500 101.940 149.650 104.675 ;
        RECT 156.965 103.015 157.115 112.565 ;
        RECT 149.120 101.705 149.650 101.940 ;
        RECT 150.960 102.865 157.115 103.015 ;
        RECT 149.120 101.470 149.640 101.705 ;
        RECT 141.630 98.955 142.180 99.310 ;
        RECT 141.660 98.840 142.180 98.955 ;
        RECT 144.640 98.870 145.160 99.340 ;
        RECT 147.540 99.075 148.230 99.390 ;
        RECT 150.960 99.310 151.110 102.865 ;
        RECT 157.270 102.720 157.410 127.520 ;
        RECT 152.470 102.580 157.410 102.720 ;
        RECT 152.470 102.060 152.610 102.580 ;
        RECT 157.555 102.375 157.705 142.475 ;
        RECT 152.090 101.590 152.610 102.060 ;
        RECT 153.960 102.225 157.705 102.375 ;
        RECT 147.560 98.860 148.230 99.075 ;
        RECT 150.570 99.055 151.110 99.310 ;
        RECT 153.960 99.280 154.110 102.225 ;
        RECT 155.040 101.990 155.560 102.050 ;
        RECT 157.890 101.990 158.030 157.500 ;
        RECT 155.040 101.850 158.030 101.990 ;
        RECT 155.040 101.580 155.560 101.850 ;
        RECT 158.205 99.285 158.350 172.505 ;
        RECT 153.580 99.115 154.110 99.280 ;
        RECT 156.480 99.140 158.350 99.285 ;
        RECT 150.570 98.840 151.090 99.055 ;
        RECT 153.580 98.810 154.100 99.115 ;
        RECT 156.510 98.780 157.030 99.140 ;
        RECT 109.980 92.665 111.040 92.925 ;
        RECT 111.640 92.685 112.700 92.945 ;
        RECT 82.020 90.870 82.280 91.190 ;
        RECT 89.840 90.870 90.100 91.190 ;
        RECT 81.560 85.430 81.820 85.750 ;
        RECT 80.640 80.330 80.900 80.650 ;
        RECT 78.340 79.990 78.600 80.310 ;
        RECT 78.800 79.990 79.060 80.310 ;
        RECT 80.180 79.990 80.440 80.310 ;
        RECT 78.400 78.610 78.540 79.990 ;
        RECT 78.340 78.290 78.600 78.610 ;
        RECT 77.940 77.930 78.540 78.010 ;
        RECT 77.940 77.870 78.600 77.930 ;
        RECT 78.340 77.610 78.600 77.870 ;
        RECT 77.420 72.170 77.680 72.490 ;
        RECT 77.880 72.170 78.140 72.490 ;
        RECT 76.040 71.920 77.160 72.060 ;
        RECT 76.040 71.830 76.300 71.920 ;
        RECT 75.580 71.150 75.840 71.470 ;
        RECT 75.640 70.450 75.780 71.150 ;
        RECT 75.580 70.130 75.840 70.450 ;
        RECT 76.960 69.790 77.220 70.110 ;
        RECT 75.120 69.450 75.380 69.770 ;
        RECT 77.020 67.050 77.160 69.790 ;
        RECT 77.480 67.390 77.620 72.170 ;
        RECT 77.940 70.450 78.080 72.170 ;
        RECT 77.880 70.130 78.140 70.450 ;
        RECT 78.400 69.850 78.540 77.610 ;
        RECT 78.860 75.210 79.000 79.990 ;
        RECT 79.260 79.310 79.520 79.630 ;
        RECT 78.800 74.890 79.060 75.210 ;
        RECT 77.940 69.710 78.540 69.850 ;
        RECT 77.420 67.070 77.680 67.390 ;
        RECT 76.500 66.730 76.760 67.050 ;
        RECT 76.960 66.730 77.220 67.050 ;
        RECT 76.560 66.370 76.700 66.730 ;
        RECT 76.500 66.050 76.760 66.370 ;
        RECT 77.020 64.970 77.160 66.730 ;
        RECT 77.480 66.370 77.620 67.070 ;
        RECT 77.420 66.050 77.680 66.370 ;
        RECT 76.560 64.830 77.160 64.970 ;
        RECT 74.660 61.630 74.920 61.950 ;
        RECT 74.200 58.570 74.460 58.890 ;
        RECT 74.720 58.800 74.860 61.630 ;
        RECT 75.580 58.800 75.840 58.890 ;
        RECT 74.720 58.660 75.840 58.800 ;
        RECT 75.580 58.570 75.840 58.660 ;
        RECT 73.740 58.230 74.000 58.550 ;
        RECT 73.280 57.890 73.540 58.210 ;
        RECT 72.360 56.530 72.620 56.850 ;
        RECT 71.900 55.850 72.160 56.170 ;
        RECT 72.420 56.080 72.560 56.530 ;
        RECT 74.260 56.510 74.400 58.570 ;
        RECT 76.560 58.550 76.700 64.830 ;
        RECT 76.960 64.010 77.220 64.330 ;
        RECT 77.020 61.610 77.160 64.010 ;
        RECT 77.940 63.990 78.080 69.710 ;
        RECT 78.860 69.090 79.000 74.890 ;
        RECT 79.320 72.490 79.460 79.310 ;
        RECT 79.720 77.270 79.980 77.590 ;
        RECT 79.260 72.170 79.520 72.490 ;
        RECT 79.320 70.110 79.460 72.170 ;
        RECT 79.780 72.150 79.920 77.270 ;
        RECT 80.240 73.170 80.380 79.990 ;
        RECT 80.700 75.210 80.840 80.330 ;
        RECT 81.620 79.970 81.760 85.430 ;
        RECT 81.560 79.650 81.820 79.970 ;
        RECT 80.640 74.890 80.900 75.210 ;
        RECT 81.560 74.890 81.820 75.210 ;
        RECT 81.100 74.210 81.360 74.530 ;
        RECT 80.180 72.850 80.440 73.170 ;
        RECT 79.720 71.830 79.980 72.150 ;
        RECT 79.260 69.790 79.520 70.110 ;
        RECT 80.240 69.770 80.380 72.850 ;
        RECT 80.180 69.450 80.440 69.770 ;
        RECT 79.260 69.110 79.520 69.430 ;
        RECT 78.800 68.770 79.060 69.090 ;
        RECT 78.860 68.490 79.000 68.770 ;
        RECT 78.400 68.350 79.000 68.490 ;
        RECT 77.880 63.670 78.140 63.990 ;
        RECT 76.960 61.290 77.220 61.610 ;
        RECT 77.880 61.290 78.140 61.610 ;
        RECT 77.420 60.610 77.680 60.930 ;
        RECT 77.480 59.570 77.620 60.610 ;
        RECT 76.960 59.250 77.220 59.570 ;
        RECT 77.420 59.250 77.680 59.570 ;
        RECT 76.040 58.230 76.300 58.550 ;
        RECT 76.500 58.230 76.760 58.550 ;
        RECT 76.100 57.870 76.240 58.230 ;
        RECT 76.040 57.550 76.300 57.870 ;
        RECT 74.200 56.190 74.460 56.510 ;
        RECT 72.820 56.080 73.080 56.170 ;
        RECT 72.420 55.940 73.080 56.080 ;
        RECT 72.820 55.850 73.080 55.940 ;
        RECT 75.580 54.830 75.840 55.150 ;
        RECT 75.640 53.110 75.780 54.830 ;
        RECT 76.100 53.790 76.240 57.550 ;
        RECT 76.560 56.170 76.700 58.230 ;
        RECT 77.020 56.930 77.160 59.250 ;
        RECT 77.020 56.790 77.620 56.930 ;
        RECT 77.940 56.850 78.080 61.290 ;
        RECT 78.400 58.460 78.540 68.350 ;
        RECT 78.800 66.730 79.060 67.050 ;
        RECT 78.860 65.010 79.000 66.730 ;
        RECT 78.800 64.690 79.060 65.010 ;
        RECT 79.320 62.290 79.460 69.110 ;
        RECT 79.720 68.770 79.980 69.090 ;
        RECT 79.780 67.390 79.920 68.770 ;
        RECT 79.720 67.070 79.980 67.390 ;
        RECT 80.240 66.960 80.380 69.450 ;
        RECT 80.640 66.960 80.900 67.050 ;
        RECT 80.240 66.820 80.900 66.960 ;
        RECT 79.720 63.670 79.980 63.990 ;
        RECT 79.260 61.970 79.520 62.290 ;
        RECT 78.800 58.460 79.060 58.550 ;
        RECT 78.400 58.320 79.060 58.460 ;
        RECT 78.800 58.230 79.060 58.320 ;
        RECT 76.960 56.190 77.220 56.510 ;
        RECT 76.500 55.850 76.760 56.170 ;
        RECT 76.040 53.470 76.300 53.790 ;
        RECT 77.020 53.110 77.160 56.190 ;
        RECT 75.580 52.790 75.840 53.110 ;
        RECT 76.960 52.790 77.220 53.110 ;
        RECT 71.440 52.450 71.700 52.770 ;
        RECT 77.480 51.070 77.620 56.790 ;
        RECT 77.880 56.530 78.140 56.850 ;
        RECT 79.780 56.510 79.920 63.670 ;
        RECT 80.240 58.550 80.380 66.820 ;
        RECT 80.640 66.730 80.900 66.820 ;
        RECT 80.640 66.050 80.900 66.370 ;
        RECT 80.700 60.590 80.840 66.050 ;
        RECT 81.160 61.610 81.300 74.210 ;
        RECT 81.620 67.050 81.760 74.890 ;
        RECT 82.080 74.190 82.220 90.870 ;
        RECT 87.080 90.190 87.340 90.510 ;
        RECT 82.940 88.490 83.200 88.810 ;
        RECT 83.000 86.770 83.140 88.490 ;
        RECT 84.780 87.470 85.040 87.790 ;
        RECT 82.940 86.450 83.200 86.770 ;
        RECT 84.840 85.410 84.980 87.470 ;
        RECT 87.140 85.750 87.280 90.190 ;
        RECT 89.900 89.490 90.040 90.870 ;
        RECT 100.150 90.045 100.470 90.915 ;
        RECT 87.540 89.170 87.800 89.490 ;
        RECT 89.840 89.170 90.100 89.490 ;
        RECT 87.600 85.750 87.740 89.170 ;
        RECT 100.140 89.015 100.470 90.045 ;
        RECT 101.820 90.025 102.140 90.905 ;
        RECT 88.920 88.490 89.180 88.810 ;
        RECT 88.980 86.770 89.120 88.490 ;
        RECT 89.830 87.955 90.110 88.325 ;
        RECT 89.840 87.810 90.100 87.955 ;
        RECT 100.140 87.255 100.450 89.015 ;
        RECT 101.800 89.005 102.140 90.025 ;
        RECT 103.380 89.005 103.700 90.905 ;
        RECT 104.920 90.015 105.240 90.915 ;
        RECT 104.900 89.015 105.240 90.015 ;
        RECT 106.510 89.825 106.830 90.935 ;
        RECT 101.800 87.365 102.110 89.005 ;
        RECT 100.140 87.095 100.360 87.255 ;
        RECT 100.610 87.095 101.150 87.235 ;
        RECT 88.920 86.450 89.180 86.770 ;
        RECT 87.080 85.430 87.340 85.750 ;
        RECT 87.540 85.430 87.800 85.750 ;
        RECT 84.780 85.090 85.040 85.410 ;
        RECT 100.140 85.005 101.150 87.095 ;
        RECT 100.180 84.985 101.150 85.005 ;
        RECT 101.800 87.045 102.610 87.365 ;
        RECT 103.380 87.235 103.690 89.005 ;
        RECT 101.800 84.985 102.530 87.045 ;
        RECT 100.540 84.895 101.150 84.985 ;
        RECT 102.080 84.955 102.530 84.985 ;
        RECT 102.110 84.925 102.480 84.955 ;
        RECT 103.380 84.945 104.050 87.235 ;
        RECT 104.900 87.215 105.210 89.015 ;
        RECT 106.470 87.245 106.840 89.825 ;
        RECT 108.070 89.815 108.390 90.905 ;
        RECT 109.660 89.855 109.980 90.925 ;
        RECT 111.260 90.165 111.540 90.915 ;
        RECT 108.050 87.275 108.420 89.815 ;
        RECT 104.900 84.975 105.560 87.215 ;
        RECT 103.500 84.885 104.050 84.945 ;
        RECT 105.010 84.865 105.560 84.975 ;
        RECT 106.470 84.895 107.020 87.245 ;
        RECT 107.950 84.925 108.500 87.275 ;
        RECT 109.660 87.265 110.010 89.855 ;
        RECT 111.240 87.275 111.540 90.165 ;
        RECT 109.400 85.015 110.010 87.265 ;
        RECT 109.400 84.915 109.950 85.015 ;
        RECT 110.900 84.985 111.540 87.275 ;
        RECT 122.930 88.730 123.320 91.520 ;
        RECT 126.380 88.730 126.830 91.510 ;
        RECT 122.930 86.070 126.830 88.730 ;
        RECT 110.900 84.925 111.450 84.985 ;
        RECT 121.560 83.790 122.110 84.300 ;
        RECT 122.930 83.530 123.320 86.070 ;
        RECT 125.240 84.070 125.500 84.390 ;
        RECT 88.460 83.050 88.720 83.370 ;
        RECT 86.620 82.030 86.880 82.350 ;
        RECT 87.080 82.030 87.340 82.350 ;
        RECT 86.160 81.010 86.420 81.330 ;
        RECT 83.400 79.650 83.660 79.970 ;
        RECT 83.460 78.610 83.600 79.650 ;
        RECT 85.700 79.310 85.960 79.630 ;
        RECT 83.400 78.290 83.660 78.610 ;
        RECT 85.760 78.270 85.900 79.310 ;
        RECT 85.700 77.950 85.960 78.270 ;
        RECT 86.220 77.590 86.360 81.010 ;
        RECT 86.680 80.310 86.820 82.030 ;
        RECT 86.620 79.990 86.880 80.310 ;
        RECT 87.140 78.610 87.280 82.030 ;
        RECT 88.520 81.330 88.660 83.050 ;
        RECT 125.245 82.985 125.495 84.070 ;
        RECT 126.380 83.570 126.830 86.070 ;
        RECT 135.870 84.040 138.500 84.390 ;
        RECT 135.870 83.840 136.140 84.040 ;
        RECT 133.725 82.985 134.115 83.010 ;
        RECT 100.740 82.395 101.000 82.810 ;
        RECT 112.835 82.735 134.115 82.985 ;
        RECT 112.835 82.395 113.085 82.735 ;
        RECT 133.725 82.710 134.115 82.735 ;
        RECT 100.740 82.145 113.085 82.395 ;
        RECT 117.630 82.180 118.370 82.490 ;
        RECT 127.800 82.180 128.590 82.250 ;
        RECT 100.740 81.730 101.000 82.145 ;
        RECT 88.460 81.010 88.720 81.330 ;
        RECT 89.830 81.155 90.110 81.525 ;
        RECT 117.620 81.480 128.590 82.180 ;
        RECT 89.840 81.010 90.100 81.155 ;
        RECT 117.630 81.140 118.370 81.480 ;
        RECT 127.800 81.390 128.590 81.480 ;
        RECT 135.460 79.960 136.140 83.840 ;
        RECT 135.850 79.740 136.130 79.960 ;
        RECT 135.850 79.420 138.990 79.740 ;
        RECT 136.730 79.410 137.060 79.420 ;
        RECT 137.690 79.410 138.020 79.420 ;
        RECT 138.650 79.410 138.980 79.420 ;
        RECT 87.080 78.290 87.340 78.610 ;
        RECT 134.410 78.430 135.590 79.090 ;
        RECT 136.950 78.440 137.470 78.900 ;
        RECT 134.410 78.090 136.250 78.430 ;
        RECT 139.240 78.300 139.890 78.860 ;
        RECT 134.410 78.080 135.590 78.090 ;
        RECT 88.460 77.610 88.720 77.930 ;
        RECT 135.980 77.880 136.210 78.090 ;
        RECT 86.160 77.270 86.420 77.590 ;
        RECT 88.520 75.890 88.660 77.610 ;
        RECT 135.980 77.560 138.490 77.880 ;
        RECT 88.920 76.590 89.180 76.910 ;
        RECT 88.460 75.570 88.720 75.890 ;
        RECT 88.000 74.550 88.260 74.870 ;
        RECT 82.940 74.210 83.200 74.530 ;
        RECT 82.020 73.870 82.280 74.190 ;
        RECT 83.000 73.170 83.140 74.210 ;
        RECT 82.940 72.850 83.200 73.170 ;
        RECT 87.540 69.110 87.800 69.430 ;
        RECT 82.940 68.770 83.200 69.090 ;
        RECT 81.560 66.730 81.820 67.050 ;
        RECT 82.480 66.730 82.740 67.050 ;
        RECT 81.620 64.330 81.760 66.730 ;
        RECT 81.560 64.010 81.820 64.330 ;
        RECT 81.100 61.290 81.360 61.610 ;
        RECT 80.640 60.270 80.900 60.590 ;
        RECT 80.180 58.230 80.440 58.550 ;
        RECT 79.720 56.190 79.980 56.510 ;
        RECT 80.180 55.740 80.440 55.830 ;
        RECT 80.700 55.740 80.840 60.270 ;
        RECT 81.620 58.890 81.760 64.010 ;
        RECT 81.560 58.800 81.820 58.890 ;
        RECT 81.160 58.660 81.820 58.800 ;
        RECT 81.160 56.170 81.300 58.660 ;
        RECT 81.560 58.570 81.820 58.660 ;
        RECT 81.100 55.850 81.360 56.170 ;
        RECT 82.020 55.850 82.280 56.170 ;
        RECT 80.180 55.600 80.840 55.740 ;
        RECT 80.180 55.510 80.440 55.600 ;
        RECT 81.160 53.790 81.300 55.850 ;
        RECT 82.080 54.130 82.220 55.850 ;
        RECT 82.020 53.810 82.280 54.130 ;
        RECT 81.100 53.470 81.360 53.790 ;
        RECT 78.340 52.110 78.600 52.430 ;
        RECT 77.880 51.090 78.140 51.410 ;
        RECT 77.420 50.750 77.680 51.070 ;
        RECT 71.900 48.370 72.160 48.690 ;
        RECT 71.960 47.670 72.100 48.370 ;
        RECT 74.200 47.690 74.460 48.010 ;
        RECT 68.680 47.350 68.940 47.670 ;
        RECT 70.520 47.580 70.780 47.670 ;
        RECT 71.900 47.580 72.160 47.670 ;
        RECT 70.520 47.440 71.180 47.580 ;
        RECT 70.520 47.350 70.780 47.440 ;
        RECT 68.740 46.990 68.880 47.350 ;
        RECT 68.680 46.670 68.940 46.990 ;
        RECT 67.300 45.310 67.560 45.630 ;
        RECT 66.380 44.970 66.640 45.290 ;
        RECT 67.300 44.630 67.560 44.950 ;
        RECT 65.520 42.510 66.120 42.650 ;
        RECT 65.460 41.570 65.720 41.890 ;
        RECT 65.520 40.530 65.660 41.570 ;
        RECT 65.460 40.210 65.720 40.530 ;
        RECT 65.000 33.070 65.260 33.390 ;
        RECT 64.540 29.330 64.800 29.650 ;
        RECT 63.160 28.650 63.420 28.970 ;
        RECT 64.080 28.650 64.340 28.970 ;
        RECT 62.700 27.970 62.960 28.290 ;
        RECT 60.860 23.210 61.120 23.530 ;
        RECT 59.020 22.190 59.280 22.510 ;
        RECT 59.080 20.470 59.220 22.190 ;
        RECT 58.560 20.150 58.820 20.470 ;
        RECT 59.020 20.150 59.280 20.470 ;
        RECT 58.100 19.470 58.360 19.790 ;
        RECT 58.620 18.430 58.760 20.150 ;
        RECT 62.700 19.470 62.960 19.790 ;
        RECT 58.560 18.110 58.820 18.430 ;
        RECT 62.760 17.410 62.900 19.470 ;
        RECT 62.700 17.090 62.960 17.410 ;
        RECT 57.640 14.710 57.900 15.030 ;
        RECT 63.220 14.690 63.360 28.650 ;
        RECT 64.140 23.530 64.280 28.650 ;
        RECT 65.980 24.210 66.120 42.510 ;
        RECT 67.360 42.230 67.500 44.630 ;
        RECT 68.740 42.230 68.880 46.670 ;
        RECT 69.140 44.970 69.400 45.290 ;
        RECT 67.300 41.910 67.560 42.230 ;
        RECT 68.680 41.910 68.940 42.230 ;
        RECT 68.740 39.850 68.880 41.910 ;
        RECT 69.200 40.190 69.340 44.970 ;
        RECT 70.060 41.570 70.320 41.890 ;
        RECT 69.140 39.870 69.400 40.190 ;
        RECT 66.840 39.530 67.100 39.850 ;
        RECT 68.680 39.530 68.940 39.850 ;
        RECT 69.600 39.530 69.860 39.850 ;
        RECT 66.900 38.830 67.040 39.530 ;
        RECT 66.840 38.510 67.100 38.830 ;
        RECT 66.900 36.790 67.040 38.510 ;
        RECT 66.840 36.470 67.100 36.790 ;
        RECT 67.300 34.770 67.560 35.090 ;
        RECT 67.360 28.970 67.500 34.770 ;
        RECT 67.760 31.030 68.020 31.350 ;
        RECT 67.820 29.310 67.960 31.030 ;
        RECT 67.760 28.990 68.020 29.310 ;
        RECT 67.300 28.880 67.560 28.970 ;
        RECT 66.440 28.740 67.560 28.880 ;
        RECT 65.920 23.890 66.180 24.210 ;
        RECT 64.080 23.210 64.340 23.530 ;
        RECT 64.140 18.430 64.280 23.210 ;
        RECT 65.980 23.190 66.120 23.890 ;
        RECT 66.440 23.530 66.580 28.740 ;
        RECT 67.300 28.650 67.560 28.740 ;
        RECT 68.220 28.650 68.480 28.970 ;
        RECT 68.280 28.370 68.420 28.650 ;
        RECT 67.360 28.290 68.420 28.370 ;
        RECT 67.300 28.230 68.420 28.290 ;
        RECT 67.300 27.970 67.560 28.230 ;
        RECT 67.360 23.530 67.500 27.970 ;
        RECT 68.740 25.910 68.880 39.530 ;
        RECT 69.660 39.170 69.800 39.530 ;
        RECT 69.600 38.850 69.860 39.170 ;
        RECT 69.600 34.430 69.860 34.750 ;
        RECT 69.660 32.450 69.800 34.430 ;
        RECT 70.120 32.450 70.260 41.570 ;
        RECT 71.040 41.550 71.180 47.440 ;
        RECT 71.500 47.440 72.160 47.580 ;
        RECT 70.980 41.230 71.240 41.550 ;
        RECT 71.040 39.850 71.180 41.230 ;
        RECT 71.500 40.190 71.640 47.440 ;
        RECT 71.900 47.350 72.160 47.440 ;
        RECT 74.260 47.330 74.400 47.690 ;
        RECT 72.360 47.010 72.620 47.330 ;
        RECT 74.200 47.010 74.460 47.330 ;
        RECT 75.120 47.010 75.380 47.330 ;
        RECT 72.420 44.010 72.560 47.010 ;
        RECT 73.280 46.670 73.540 46.990 ;
        RECT 72.420 43.870 73.020 44.010 ;
        RECT 72.360 42.930 72.620 43.250 ;
        RECT 71.900 41.910 72.160 42.230 ;
        RECT 71.960 41.550 72.100 41.910 ;
        RECT 71.900 41.230 72.160 41.550 ;
        RECT 71.440 39.870 71.700 40.190 ;
        RECT 72.420 39.850 72.560 42.930 ;
        RECT 72.880 42.230 73.020 43.870 ;
        RECT 73.340 42.570 73.480 46.670 ;
        RECT 74.260 45.970 74.400 47.010 ;
        RECT 74.200 45.650 74.460 45.970 ;
        RECT 73.740 44.970 74.000 45.290 ;
        RECT 73.800 43.250 73.940 44.970 ;
        RECT 73.740 42.930 74.000 43.250 ;
        RECT 73.280 42.250 73.540 42.570 ;
        RECT 72.820 41.910 73.080 42.230 ;
        RECT 73.280 41.230 73.540 41.550 ;
        RECT 74.660 41.460 74.920 41.550 ;
        RECT 75.180 41.460 75.320 47.010 ;
        RECT 74.660 41.320 75.320 41.460 ;
        RECT 74.660 41.230 74.920 41.320 ;
        RECT 70.980 39.530 71.240 39.850 ;
        RECT 72.360 39.760 72.620 39.850 ;
        RECT 71.960 39.620 72.620 39.760 ;
        RECT 69.660 32.310 70.260 32.450 ;
        RECT 70.060 30.350 70.320 30.670 ;
        RECT 69.600 29.330 69.860 29.650 ;
        RECT 69.660 28.290 69.800 29.330 ;
        RECT 70.120 28.970 70.260 30.350 ;
        RECT 70.060 28.650 70.320 28.970 ;
        RECT 69.600 27.970 69.860 28.290 ;
        RECT 68.680 25.590 68.940 25.910 ;
        RECT 66.380 23.210 66.640 23.530 ;
        RECT 67.300 23.440 67.560 23.530 ;
        RECT 66.900 23.300 67.560 23.440 ;
        RECT 65.450 22.675 65.730 23.045 ;
        RECT 65.920 22.870 66.180 23.190 ;
        RECT 65.460 22.530 65.720 22.675 ;
        RECT 64.080 18.110 64.340 18.430 ;
        RECT 66.440 18.090 66.580 23.210 ;
        RECT 66.900 18.340 67.040 23.300 ;
        RECT 67.300 23.210 67.560 23.300 ;
        RECT 67.760 23.210 68.020 23.530 ;
        RECT 67.300 22.190 67.560 22.510 ;
        RECT 67.360 20.130 67.500 22.190 ;
        RECT 67.300 19.810 67.560 20.130 ;
        RECT 67.820 19.790 67.960 23.210 ;
        RECT 69.140 22.870 69.400 23.190 ;
        RECT 67.760 19.470 68.020 19.790 ;
        RECT 67.300 18.340 67.560 18.430 ;
        RECT 66.900 18.200 67.560 18.340 ;
        RECT 67.300 18.110 67.560 18.200 ;
        RECT 66.380 17.770 66.640 18.090 ;
        RECT 65.000 17.430 65.260 17.750 ;
        RECT 65.060 15.030 65.200 17.430 ;
        RECT 67.820 15.030 67.960 19.470 ;
        RECT 69.200 15.370 69.340 22.870 ;
        RECT 70.520 22.760 70.780 22.850 ;
        RECT 69.660 22.620 70.780 22.760 ;
        RECT 69.660 21.490 69.800 22.620 ;
        RECT 70.520 22.530 70.780 22.620 ;
        RECT 69.600 21.170 69.860 21.490 ;
        RECT 70.060 20.150 70.320 20.470 ;
        RECT 70.120 17.750 70.260 20.150 ;
        RECT 70.060 17.430 70.320 17.750 ;
        RECT 69.140 15.050 69.400 15.370 ;
        RECT 71.040 15.030 71.180 39.530 ;
        RECT 71.960 34.070 72.100 39.620 ;
        RECT 72.360 39.530 72.620 39.620 ;
        RECT 73.340 39.510 73.480 41.230 ;
        RECT 73.280 39.190 73.540 39.510 ;
        RECT 72.360 38.740 72.620 38.830 ;
        RECT 73.340 38.740 73.480 39.190 ;
        RECT 75.180 38.830 75.320 41.320 ;
        RECT 75.580 39.530 75.840 39.850 ;
        RECT 72.360 38.600 73.480 38.740 ;
        RECT 72.360 38.510 72.620 38.600 ;
        RECT 75.120 38.510 75.380 38.830 ;
        RECT 71.900 33.750 72.160 34.070 ;
        RECT 71.900 29.220 72.160 29.310 ;
        RECT 72.420 29.220 72.560 38.510 ;
        RECT 74.660 37.150 74.920 37.470 ;
        RECT 74.200 35.790 74.460 36.110 ;
        RECT 74.260 34.070 74.400 35.790 ;
        RECT 74.200 33.750 74.460 34.070 ;
        RECT 73.280 31.030 73.540 31.350 ;
        RECT 72.820 30.690 73.080 31.010 ;
        RECT 72.880 29.650 73.020 30.690 ;
        RECT 72.820 29.330 73.080 29.650 ;
        RECT 73.340 29.310 73.480 31.030 ;
        RECT 71.900 29.080 72.560 29.220 ;
        RECT 71.900 28.990 72.160 29.080 ;
        RECT 73.280 28.990 73.540 29.310 ;
        RECT 71.960 24.210 72.100 28.990 ;
        RECT 74.260 26.250 74.400 33.750 ;
        RECT 74.200 25.930 74.460 26.250 ;
        RECT 71.900 23.890 72.160 24.210 ;
        RECT 73.280 23.210 73.540 23.530 ;
        RECT 73.340 21.490 73.480 23.210 ;
        RECT 73.280 21.400 73.540 21.490 ;
        RECT 72.880 21.260 73.540 21.400 ;
        RECT 72.880 18.770 73.020 21.260 ;
        RECT 73.280 21.170 73.540 21.260 ;
        RECT 74.260 20.810 74.400 25.930 ;
        RECT 74.720 21.490 74.860 37.150 ;
        RECT 75.180 36.450 75.320 38.510 ;
        RECT 75.120 36.130 75.380 36.450 ;
        RECT 75.180 31.010 75.320 36.130 ;
        RECT 75.640 34.750 75.780 39.530 ;
        RECT 75.580 34.430 75.840 34.750 ;
        RECT 75.120 30.690 75.380 31.010 ;
        RECT 75.180 23.870 75.320 30.690 ;
        RECT 75.640 23.870 75.780 34.430 ;
        RECT 77.410 34.235 77.690 34.605 ;
        RECT 77.420 34.090 77.680 34.235 ;
        RECT 77.940 33.730 78.080 51.090 ;
        RECT 78.400 50.730 78.540 52.110 ;
        RECT 78.340 50.410 78.600 50.730 ;
        RECT 79.260 47.350 79.520 47.670 ;
        RECT 79.720 47.350 79.980 47.670 ;
        RECT 80.180 47.350 80.440 47.670 ;
        RECT 78.340 45.310 78.600 45.630 ;
        RECT 78.400 42.230 78.540 45.310 ;
        RECT 79.320 43.250 79.460 47.350 ;
        RECT 79.260 42.930 79.520 43.250 ;
        RECT 78.340 41.910 78.600 42.230 ;
        RECT 79.260 39.530 79.520 39.850 ;
        RECT 79.320 36.790 79.460 39.530 ;
        RECT 79.780 39.510 79.920 47.350 ;
        RECT 79.720 39.190 79.980 39.510 ;
        RECT 80.240 39.170 80.380 47.350 ;
        RECT 81.560 46.670 81.820 46.990 ;
        RECT 81.620 41.890 81.760 46.670 ;
        RECT 81.560 41.570 81.820 41.890 ;
        RECT 82.540 39.850 82.680 66.730 ;
        RECT 81.100 39.530 81.360 39.850 ;
        RECT 82.480 39.530 82.740 39.850 ;
        RECT 80.180 38.850 80.440 39.170 ;
        RECT 81.160 37.810 81.300 39.530 ;
        RECT 81.100 37.490 81.360 37.810 ;
        RECT 82.540 37.130 82.680 39.530 ;
        RECT 82.480 36.810 82.740 37.130 ;
        RECT 79.260 36.470 79.520 36.790 ;
        RECT 80.180 36.470 80.440 36.790 ;
        RECT 76.960 33.410 77.220 33.730 ;
        RECT 77.880 33.410 78.140 33.730 ;
        RECT 77.020 25.820 77.160 33.410 ;
        RECT 79.320 29.050 79.460 36.470 ;
        RECT 79.720 36.130 79.980 36.450 ;
        RECT 79.780 34.750 79.920 36.130 ;
        RECT 80.240 35.090 80.380 36.470 ;
        RECT 80.180 34.770 80.440 35.090 ;
        RECT 79.720 34.430 79.980 34.750 ;
        RECT 80.180 34.090 80.440 34.410 ;
        RECT 81.100 34.090 81.360 34.410 ;
        RECT 82.010 34.235 82.290 34.605 ;
        RECT 82.020 34.090 82.280 34.235 ;
        RECT 80.240 33.730 80.380 34.090 ;
        RECT 80.180 33.410 80.440 33.730 ;
        RECT 81.160 33.390 81.300 34.090 ;
        RECT 82.480 33.410 82.740 33.730 ;
        RECT 81.100 33.070 81.360 33.390 ;
        RECT 79.720 30.690 79.980 31.010 ;
        RECT 79.780 29.650 79.920 30.690 ;
        RECT 80.640 30.350 80.900 30.670 ;
        RECT 79.720 29.330 79.980 29.650 ;
        RECT 78.340 28.650 78.600 28.970 ;
        RECT 78.800 28.650 79.060 28.970 ;
        RECT 79.320 28.910 80.380 29.050 ;
        RECT 78.400 26.930 78.540 28.650 ;
        RECT 78.340 26.610 78.600 26.930 ;
        RECT 78.340 25.930 78.600 26.250 ;
        RECT 77.420 25.820 77.680 25.910 ;
        RECT 77.020 25.680 77.680 25.820 ;
        RECT 77.420 25.590 77.680 25.680 ;
        RECT 75.120 23.550 75.380 23.870 ;
        RECT 75.580 23.550 75.840 23.870 ;
        RECT 74.660 21.170 74.920 21.490 ;
        RECT 74.200 20.490 74.460 20.810 ;
        RECT 74.720 20.470 74.860 21.170 ;
        RECT 74.660 20.150 74.920 20.470 ;
        RECT 73.280 19.470 73.540 19.790 ;
        RECT 72.820 18.450 73.080 18.770 ;
        RECT 72.880 15.030 73.020 18.450 ;
        RECT 73.340 18.090 73.480 19.470 ;
        RECT 73.280 17.770 73.540 18.090 ;
        RECT 75.180 16.670 75.320 23.550 ;
        RECT 76.960 23.210 77.220 23.530 ;
        RECT 77.020 20.810 77.160 23.210 ;
        RECT 76.960 20.490 77.220 20.810 ;
        RECT 75.580 20.150 75.840 20.470 ;
        RECT 75.640 18.770 75.780 20.150 ;
        RECT 75.580 18.450 75.840 18.770 ;
        RECT 77.480 18.090 77.620 25.590 ;
        RECT 78.400 24.210 78.540 25.930 ;
        RECT 78.340 23.890 78.600 24.210 ;
        RECT 78.400 22.510 78.540 23.890 ;
        RECT 78.860 23.530 79.000 28.650 ;
        RECT 79.260 25.590 79.520 25.910 ;
        RECT 79.720 25.590 79.980 25.910 ;
        RECT 79.320 24.210 79.460 25.590 ;
        RECT 79.780 24.210 79.920 25.590 ;
        RECT 79.260 23.890 79.520 24.210 ;
        RECT 79.720 23.890 79.980 24.210 ;
        RECT 80.240 23.530 80.380 28.910 ;
        RECT 80.700 25.910 80.840 30.350 ;
        RECT 81.160 28.630 81.300 33.070 ;
        RECT 82.540 28.970 82.680 33.410 ;
        RECT 82.480 28.650 82.740 28.970 ;
        RECT 81.100 28.310 81.360 28.630 ;
        RECT 83.000 28.370 83.140 68.770 ;
        RECT 84.780 68.430 85.040 68.750 ;
        RECT 85.700 68.430 85.960 68.750 ;
        RECT 87.080 68.430 87.340 68.750 ;
        RECT 83.860 67.070 84.120 67.390 ;
        RECT 83.920 65.010 84.060 67.070 ;
        RECT 83.860 64.690 84.120 65.010 ;
        RECT 83.400 60.270 83.660 60.590 ;
        RECT 83.460 58.550 83.600 60.270 ;
        RECT 83.400 58.230 83.660 58.550 ;
        RECT 83.860 55.850 84.120 56.170 ;
        RECT 83.920 45.970 84.060 55.850 ;
        RECT 84.840 53.450 84.980 68.430 ;
        RECT 85.760 67.925 85.900 68.430 ;
        RECT 85.690 67.555 85.970 67.925 ;
        RECT 86.620 67.410 86.880 67.730 ;
        RECT 85.700 65.710 85.960 66.030 ;
        RECT 85.760 64.330 85.900 65.710 ;
        RECT 86.680 64.330 86.820 67.410 ;
        RECT 85.700 64.010 85.960 64.330 ;
        RECT 86.620 64.010 86.880 64.330 ;
        RECT 87.140 63.650 87.280 68.430 ;
        RECT 87.080 63.330 87.340 63.650 ;
        RECT 85.240 62.990 85.500 63.310 ;
        RECT 85.300 62.290 85.440 62.990 ;
        RECT 87.600 62.290 87.740 69.110 ;
        RECT 88.060 66.370 88.200 74.550 ;
        RECT 88.520 72.490 88.660 75.570 ;
        RECT 88.980 74.870 89.120 76.590 ;
        RECT 135.980 76.240 136.210 77.560 ;
        RECT 137.200 77.550 137.530 77.560 ;
        RECT 138.160 77.550 138.490 77.560 ;
        RECT 135.980 75.900 138.980 76.240 ;
        RECT 88.920 74.550 89.180 74.870 ;
        RECT 89.830 74.355 90.110 74.725 ;
        RECT 89.900 74.190 90.040 74.355 ;
        RECT 89.840 73.870 90.100 74.190 ;
        RECT 88.460 72.170 88.720 72.490 ;
        RECT 90.290 70.955 90.570 71.325 ;
        RECT 89.840 69.110 90.100 69.430 ;
        RECT 89.900 67.730 90.040 69.110 ;
        RECT 88.460 67.410 88.720 67.730 ;
        RECT 89.840 67.410 90.100 67.730 ;
        RECT 88.000 66.050 88.260 66.370 ;
        RECT 88.000 63.670 88.260 63.990 ;
        RECT 85.240 61.970 85.500 62.290 ;
        RECT 87.540 61.970 87.800 62.290 ;
        RECT 85.700 60.950 85.960 61.270 ;
        RECT 85.760 59.570 85.900 60.950 ;
        RECT 88.060 59.570 88.200 63.670 ;
        RECT 88.520 61.610 88.660 67.410 ;
        RECT 90.360 67.050 90.500 70.955 ;
        RECT 90.300 66.730 90.560 67.050 ;
        RECT 89.840 64.525 90.100 64.670 ;
        RECT 89.830 64.155 90.110 64.525 ;
        RECT 89.380 63.670 89.640 63.990 ;
        RECT 88.460 61.290 88.720 61.610 ;
        RECT 88.920 61.290 89.180 61.610 ;
        RECT 85.700 59.250 85.960 59.570 ;
        RECT 88.000 59.250 88.260 59.570 ;
        RECT 85.240 54.830 85.500 55.150 ;
        RECT 87.540 54.830 87.800 55.150 ;
        RECT 85.300 53.450 85.440 54.830 ;
        RECT 87.600 53.450 87.740 54.830 ;
        RECT 84.780 53.130 85.040 53.450 ;
        RECT 85.240 53.130 85.500 53.450 ;
        RECT 87.540 53.130 87.800 53.450 ;
        RECT 88.980 50.050 89.120 61.290 ;
        RECT 89.440 59.570 89.580 63.670 ;
        RECT 89.830 60.755 90.110 61.125 ;
        RECT 89.840 60.610 90.100 60.755 ;
        RECT 89.380 59.250 89.640 59.570 ;
        RECT 89.840 54.830 90.100 55.150 ;
        RECT 89.900 54.325 90.040 54.830 ;
        RECT 89.830 53.955 90.110 54.325 ;
        RECT 90.300 53.130 90.560 53.450 ;
        RECT 90.360 50.730 90.500 53.130 ;
        RECT 90.300 50.410 90.560 50.730 ;
        RECT 88.920 49.730 89.180 50.050 ;
        RECT 84.780 47.010 85.040 47.330 ;
        RECT 83.860 45.650 84.120 45.970 ;
        RECT 83.400 41.910 83.660 42.230 ;
        RECT 83.460 36.790 83.600 41.910 ;
        RECT 84.840 39.850 84.980 47.010 ;
        RECT 88.920 44.970 89.180 45.290 ;
        RECT 88.980 41.550 89.120 44.970 ;
        RECT 90.760 44.290 91.020 44.610 ;
        RECT 90.820 44.125 90.960 44.290 ;
        RECT 90.750 43.755 91.030 44.125 ;
        RECT 88.920 41.230 89.180 41.550 ;
        RECT 84.780 39.530 85.040 39.850 ;
        RECT 84.780 38.850 85.040 39.170 ;
        RECT 83.400 36.470 83.660 36.790 ;
        RECT 83.460 34.070 83.600 36.470 ;
        RECT 84.840 34.750 84.980 38.850 ;
        RECT 87.080 35.790 87.340 36.110 ;
        RECT 84.780 34.430 85.040 34.750 ;
        RECT 87.140 34.410 87.280 35.790 ;
        RECT 88.920 34.770 89.180 35.090 ;
        RECT 87.080 34.090 87.340 34.410 ;
        RECT 83.400 33.750 83.660 34.070 ;
        RECT 83.460 29.310 83.600 33.750 ;
        RECT 83.860 31.710 84.120 32.030 ;
        RECT 83.400 28.990 83.660 29.310 ;
        RECT 82.540 28.230 83.140 28.370 ;
        RECT 81.560 27.630 81.820 27.950 ;
        RECT 81.100 25.930 81.360 26.250 ;
        RECT 80.640 25.590 80.900 25.910 ;
        RECT 80.640 24.910 80.900 25.230 ;
        RECT 80.700 23.530 80.840 24.910 ;
        RECT 78.800 23.210 79.060 23.530 ;
        RECT 79.260 23.210 79.520 23.530 ;
        RECT 80.180 23.440 80.440 23.530 ;
        RECT 79.780 23.300 80.440 23.440 ;
        RECT 78.340 22.190 78.600 22.510 ;
        RECT 78.800 20.150 79.060 20.470 ;
        RECT 78.860 19.790 79.000 20.150 ;
        RECT 78.800 19.470 79.060 19.790 ;
        RECT 79.320 18.090 79.460 23.210 ;
        RECT 79.780 21.150 79.920 23.300 ;
        RECT 80.180 23.210 80.440 23.300 ;
        RECT 80.640 23.210 80.900 23.530 ;
        RECT 80.180 22.190 80.440 22.510 ;
        RECT 79.720 20.830 79.980 21.150 ;
        RECT 80.240 20.470 80.380 22.190 ;
        RECT 79.720 20.150 79.980 20.470 ;
        RECT 80.180 20.150 80.440 20.470 ;
        RECT 80.640 20.150 80.900 20.470 ;
        RECT 77.420 17.770 77.680 18.090 ;
        RECT 79.260 17.770 79.520 18.090 ;
        RECT 77.420 17.090 77.680 17.410 ;
        RECT 74.260 16.530 75.320 16.670 ;
        RECT 65.000 14.710 65.260 15.030 ;
        RECT 67.760 14.710 68.020 15.030 ;
        RECT 70.980 14.710 71.240 15.030 ;
        RECT 72.820 14.710 73.080 15.030 ;
        RECT 74.260 14.690 74.400 16.530 ;
        RECT 77.480 15.030 77.620 17.090 ;
        RECT 79.780 16.050 79.920 20.150 ;
        RECT 80.180 18.450 80.440 18.770 ;
        RECT 79.720 15.730 79.980 16.050 ;
        RECT 80.240 15.370 80.380 18.450 ;
        RECT 80.700 17.070 80.840 20.150 ;
        RECT 81.160 18.430 81.300 25.930 ;
        RECT 81.620 25.910 81.760 27.630 ;
        RECT 81.560 25.590 81.820 25.910 ;
        RECT 81.620 20.470 81.760 25.590 ;
        RECT 82.540 23.870 82.680 28.230 ;
        RECT 82.940 27.630 83.200 27.950 ;
        RECT 83.000 26.590 83.140 27.630 ;
        RECT 82.940 26.270 83.200 26.590 ;
        RECT 83.460 26.250 83.600 28.990 ;
        RECT 83.400 25.930 83.660 26.250 ;
        RECT 83.400 25.250 83.660 25.570 ;
        RECT 82.480 23.550 82.740 23.870 ;
        RECT 83.460 23.190 83.600 25.250 ;
        RECT 83.400 22.870 83.660 23.190 ;
        RECT 81.560 20.150 81.820 20.470 ;
        RECT 81.620 19.790 81.760 20.150 ;
        RECT 81.560 19.470 81.820 19.790 ;
        RECT 82.480 19.470 82.740 19.790 ;
        RECT 83.400 19.470 83.660 19.790 ;
        RECT 81.100 18.110 81.360 18.430 ;
        RECT 81.160 17.750 81.300 18.110 ;
        RECT 82.540 18.090 82.680 19.470 ;
        RECT 82.480 17.770 82.740 18.090 ;
        RECT 81.100 17.430 81.360 17.750 ;
        RECT 80.640 16.750 80.900 17.070 ;
        RECT 81.160 15.370 81.300 17.430 ;
        RECT 83.460 16.050 83.600 19.470 ;
        RECT 83.920 18.090 84.060 31.710 ;
        RECT 86.160 28.990 86.420 29.310 ;
        RECT 85.700 28.650 85.960 28.970 ;
        RECT 85.760 25.230 85.900 28.650 ;
        RECT 85.700 24.910 85.960 25.230 ;
        RECT 85.700 23.210 85.960 23.530 ;
        RECT 85.240 20.830 85.500 21.150 ;
        RECT 84.780 19.470 85.040 19.790 ;
        RECT 83.860 17.770 84.120 18.090 ;
        RECT 83.400 15.730 83.660 16.050 ;
        RECT 80.180 15.050 80.440 15.370 ;
        RECT 81.100 15.050 81.360 15.370 ;
        RECT 84.840 15.030 84.980 19.470 ;
        RECT 77.420 14.710 77.680 15.030 ;
        RECT 84.780 14.710 85.040 15.030 ;
        RECT 40.160 14.370 40.420 14.690 ;
        RECT 49.820 14.370 50.080 14.690 ;
        RECT 63.160 14.370 63.420 14.690 ;
        RECT 74.200 14.370 74.460 14.690 ;
        RECT 40.220 6.800 40.360 14.370 ;
        RECT 42.920 14.030 43.180 14.350 ;
        RECT 46.600 14.030 46.860 14.350 ;
        RECT 49.360 14.030 49.620 14.350 ;
        RECT 53.040 14.030 53.300 14.350 ;
        RECT 56.260 14.030 56.520 14.350 ;
        RECT 59.480 14.030 59.740 14.350 ;
        RECT 62.700 14.030 62.960 14.350 ;
        RECT 65.920 14.030 66.180 14.350 ;
        RECT 69.140 14.030 69.400 14.350 ;
        RECT 72.360 14.030 72.620 14.350 ;
        RECT 75.580 14.030 75.840 14.350 ;
        RECT 42.980 7.970 43.120 14.030 ;
        RECT 42.980 7.830 43.580 7.970 ;
        RECT 43.440 6.800 43.580 7.830 ;
        RECT 46.660 6.800 46.800 14.030 ;
        RECT 49.420 8.650 49.560 14.030 ;
        RECT 49.420 8.510 50.020 8.650 ;
        RECT 49.880 6.800 50.020 8.510 ;
        RECT 53.100 6.800 53.240 14.030 ;
        RECT 56.320 6.800 56.460 14.030 ;
        RECT 59.540 6.800 59.680 14.030 ;
        RECT 62.760 6.800 62.900 14.030 ;
        RECT 65.980 6.800 66.120 14.030 ;
        RECT 69.200 6.800 69.340 14.030 ;
        RECT 72.420 6.800 72.560 14.030 ;
        RECT 75.640 6.800 75.780 14.030 ;
        RECT 78.800 9.270 79.060 9.590 ;
        RECT 78.860 6.800 79.000 9.270 ;
        RECT 82.020 8.250 82.280 8.570 ;
        RECT 82.080 6.800 82.220 8.250 ;
        RECT 85.300 6.800 85.440 20.830 ;
        RECT 85.760 14.690 85.900 23.210 ;
        RECT 86.220 20.470 86.360 28.990 ;
        RECT 87.140 23.530 87.280 34.090 ;
        RECT 88.980 31.350 89.120 34.770 ;
        RECT 88.920 31.030 89.180 31.350 ;
        RECT 90.760 30.525 91.020 30.670 ;
        RECT 90.750 30.155 91.030 30.525 ;
        RECT 90.300 24.910 90.560 25.230 ;
        RECT 90.360 23.530 90.500 24.910 ;
        RECT 87.080 23.210 87.340 23.530 ;
        RECT 90.300 23.210 90.560 23.530 ;
        RECT 94.900 22.870 95.160 23.190 ;
        RECT 91.680 22.530 91.940 22.850 ;
        RECT 88.460 22.190 88.720 22.510 ;
        RECT 86.160 20.150 86.420 20.470 ;
        RECT 88.000 20.150 88.260 20.470 ;
        RECT 87.080 19.470 87.340 19.790 ;
        RECT 85.700 14.370 85.960 14.690 ;
        RECT 87.140 8.570 87.280 19.470 ;
        RECT 88.060 18.770 88.200 20.150 ;
        RECT 88.000 18.450 88.260 18.770 ;
        RECT 87.080 8.250 87.340 8.570 ;
        RECT 88.520 6.800 88.660 22.190 ;
        RECT 89.380 16.750 89.640 17.070 ;
        RECT 89.440 9.590 89.580 16.750 ;
        RECT 89.380 9.270 89.640 9.590 ;
        RECT 91.740 6.800 91.880 22.530 ;
        RECT 94.960 6.800 95.100 22.870 ;
        RECT 7.950 2.800 8.230 6.800 ;
        RECT 11.170 2.800 11.450 6.800 ;
        RECT 14.390 2.800 14.670 6.800 ;
        RECT 17.610 2.800 17.890 6.800 ;
        RECT 20.830 2.800 21.110 6.800 ;
        RECT 24.050 2.800 24.330 6.800 ;
        RECT 27.270 2.800 27.550 6.800 ;
        RECT 30.490 2.800 30.770 6.800 ;
        RECT 33.710 2.800 33.990 6.800 ;
        RECT 36.930 2.800 37.210 6.800 ;
        RECT 40.150 2.800 40.430 6.800 ;
        RECT 43.370 2.800 43.650 6.800 ;
        RECT 46.590 2.800 46.870 6.800 ;
        RECT 49.810 2.800 50.090 6.800 ;
        RECT 53.030 2.800 53.310 6.800 ;
        RECT 56.250 2.800 56.530 6.800 ;
        RECT 59.470 2.800 59.750 6.800 ;
        RECT 62.690 2.800 62.970 6.800 ;
        RECT 65.910 2.800 66.190 6.800 ;
        RECT 69.130 2.800 69.410 6.800 ;
        RECT 72.350 2.800 72.630 6.800 ;
        RECT 75.570 2.800 75.850 6.800 ;
        RECT 78.790 2.800 79.070 6.800 ;
        RECT 82.010 2.800 82.290 6.800 ;
        RECT 85.230 2.800 85.510 6.800 ;
        RECT 88.450 2.800 88.730 6.800 ;
        RECT 91.670 2.800 91.950 6.800 ;
        RECT 94.890 2.800 95.170 6.800 ;
      LAYER met3 ;
        RECT 63.690 224.960 64.010 225.340 ;
        RECT 63.700 218.305 64.000 224.960 ;
        RECT 66.520 224.940 66.840 225.320 ;
        RECT 69.240 224.980 69.560 225.360 ;
        RECT 72.110 225.020 72.430 225.400 ;
        RECT 66.530 218.835 66.830 224.940 ;
        RECT 69.250 222.665 69.550 224.980 ;
        RECT 69.225 222.315 69.575 222.665 ;
        RECT 72.120 222.195 72.420 225.020 ;
        RECT 74.805 224.950 75.125 225.330 ;
        RECT 77.570 224.970 77.890 225.350 ;
        RECT 72.095 221.845 72.445 222.195 ;
        RECT 74.815 221.810 75.115 224.950 ;
        RECT 74.790 221.460 75.140 221.810 ;
        RECT 77.580 219.195 77.880 224.970 ;
        RECT 80.310 224.890 80.630 225.270 ;
        RECT 83.120 224.920 83.440 225.300 ;
        RECT 85.820 225.000 86.140 225.380 ;
        RECT 80.320 221.330 80.620 224.890 ;
        RECT 80.295 220.980 80.645 221.330 ;
        RECT 83.130 221.005 83.430 224.920 ;
        RECT 83.105 220.655 83.455 221.005 ;
        RECT 85.830 220.620 86.130 225.000 ;
        RECT 88.590 224.930 88.910 225.310 ;
        RECT 91.315 224.960 91.635 225.340 ;
        RECT 93.990 224.990 94.310 225.370 ;
        RECT 142.460 225.130 142.780 225.440 ;
        RECT 85.805 220.270 86.155 220.620 ;
        RECT 88.600 219.595 88.900 224.930 ;
        RECT 91.325 220.245 91.625 224.960 ;
        RECT 91.300 219.895 91.650 220.245 ;
        RECT 94.000 219.905 94.300 224.990 ;
        RECT 142.400 224.815 142.840 225.130 ;
        RECT 115.120 220.825 115.720 224.815 ;
        RECT 115.120 220.815 116.250 220.825 ;
        RECT 125.320 220.815 125.920 224.815 ;
        RECT 132.120 220.815 132.720 224.815 ;
        RECT 138.920 220.815 139.520 224.815 ;
        RECT 142.320 220.815 142.920 224.815 ;
        RECT 115.270 220.610 116.250 220.815 ;
        RECT 115.270 220.525 116.265 220.610 ;
        RECT 115.935 220.280 116.265 220.525 ;
        RECT 88.575 219.245 88.925 219.595 ;
        RECT 93.975 219.555 94.325 219.905 ;
        RECT 77.555 218.845 77.905 219.195 ;
        RECT 66.505 218.485 66.855 218.835 ;
        RECT 125.470 218.310 125.770 220.815 ;
        RECT 132.270 220.455 132.570 220.815 ;
        RECT 132.255 220.125 132.585 220.455 ;
        RECT 132.270 218.310 132.570 220.125 ;
        RECT 139.070 218.310 139.370 220.815 ;
        RECT 63.675 217.955 64.025 218.305 ;
        RECT 125.455 217.980 125.785 218.310 ;
        RECT 132.255 217.980 132.585 218.310 ;
        RECT 139.055 217.980 139.385 218.310 ;
        RECT 142.470 207.270 142.770 220.815 ;
        RECT 143.815 208.320 144.145 208.650 ;
        RECT 142.455 206.940 142.785 207.270 ;
        RECT 143.830 204.510 144.130 208.320 ;
        RECT 143.815 204.180 144.145 204.510 ;
        RECT 103.875 203.765 105.465 203.770 ;
        RECT 103.850 202.185 105.490 203.765 ;
        RECT 114.915 202.185 115.245 203.765 ;
        RECT 120.355 202.185 120.685 203.765 ;
        RECT 125.795 202.185 126.125 203.765 ;
        RECT 131.235 202.185 131.565 203.765 ;
        RECT 136.675 202.185 137.005 203.765 ;
        RECT 142.115 202.185 142.445 203.765 ;
        RECT 28.910 201.195 30.490 201.525 ;
        RECT 100.980 199.740 102.620 200.510 ;
        RECT 32.210 198.475 33.790 198.805 ;
        RECT 8.385 198.450 8.715 198.465 ;
        RECT 8.385 198.150 13.070 198.450 ;
        RECT 8.385 198.135 8.715 198.150 ;
        RECT 7.860 197.090 11.860 197.240 ;
        RECT 12.770 197.090 13.070 198.150 ;
        RECT 7.860 196.790 13.070 197.090 ;
        RECT 7.860 196.640 11.860 196.790 ;
        RECT 28.910 195.755 30.490 196.085 ;
        RECT 32.210 193.035 33.790 193.365 ;
        RECT 46.105 192.330 46.435 192.345 ;
        RECT 51.625 192.330 51.955 192.345 ;
        RECT 46.105 192.030 51.955 192.330 ;
        RECT 46.105 192.015 46.435 192.030 ;
        RECT 51.625 192.015 51.955 192.030 ;
        RECT 28.910 190.315 30.490 190.645 ;
        RECT 32.210 187.595 33.790 187.925 ;
        RECT 28.910 184.875 30.490 185.205 ;
        RECT 101.005 184.070 102.595 199.740 ;
        RECT 60.825 183.490 61.155 183.505 ;
        RECT 63.585 183.490 63.915 183.505 ;
        RECT 60.825 183.190 63.915 183.490 ;
        RECT 60.825 183.175 61.155 183.190 ;
        RECT 63.585 183.175 63.915 183.190 ;
        RECT 32.210 182.155 33.790 182.485 ;
        RECT 100.970 182.410 102.630 184.070 ;
        RECT 28.910 179.435 30.490 179.765 ;
        RECT 32.210 176.715 33.790 177.045 ;
        RECT 103.875 176.485 105.465 202.185 ;
        RECT 109.840 198.890 113.500 200.480 ;
        RECT 112.195 198.885 112.525 198.890 ;
        RECT 117.635 198.885 117.965 200.465 ;
        RECT 123.075 198.885 123.405 200.465 ;
        RECT 128.515 198.885 128.845 200.465 ;
        RECT 133.955 198.885 134.285 200.465 ;
        RECT 139.395 198.885 139.725 200.465 ;
        RECT 115.255 193.600 115.585 193.930 ;
        RECT 111.855 189.000 112.185 189.330 ;
        RECT 108.455 185.320 108.785 185.650 ;
        RECT 108.470 181.770 108.770 185.320 ;
        RECT 111.870 181.770 112.170 189.000 ;
        RECT 115.270 181.770 115.570 193.600 ;
        RECT 125.455 192.220 125.785 192.550 ;
        RECT 118.655 190.840 118.985 191.170 ;
        RECT 118.670 181.770 118.970 190.840 ;
        RECT 122.055 188.540 122.385 188.870 ;
        RECT 122.070 181.770 122.370 188.540 ;
        RECT 125.470 181.770 125.770 192.220 ;
        RECT 143.830 191.170 144.130 204.180 ;
        RECT 147.555 202.185 147.885 203.765 ;
        RECT 144.835 198.885 145.165 200.465 ;
        RECT 148.095 195.430 148.445 195.780 ;
        RECT 143.815 190.840 144.145 191.170 ;
        RECT 128.855 189.920 129.185 190.250 ;
        RECT 128.870 181.770 129.170 189.920 ;
        RECT 135.655 187.160 135.985 187.490 ;
        RECT 132.255 184.860 132.585 185.190 ;
        RECT 132.270 181.770 132.570 184.860 ;
        RECT 135.670 181.770 135.970 187.160 ;
        RECT 145.855 186.240 146.185 186.570 ;
        RECT 139.055 184.860 139.385 185.190 ;
        RECT 142.455 184.860 142.785 185.190 ;
        RECT 139.070 181.770 139.370 184.860 ;
        RECT 142.470 181.770 142.770 184.860 ;
        RECT 145.870 181.770 146.170 186.240 ;
        RECT 108.320 177.770 108.920 181.770 ;
        RECT 111.720 177.770 112.320 181.770 ;
        RECT 115.120 177.770 115.720 181.770 ;
        RECT 118.520 177.770 119.120 181.770 ;
        RECT 121.920 177.770 122.520 181.770 ;
        RECT 125.320 177.770 125.920 181.770 ;
        RECT 128.720 177.770 129.320 181.770 ;
        RECT 132.120 177.770 132.720 181.770 ;
        RECT 135.520 177.770 136.120 181.770 ;
        RECT 138.920 177.770 139.520 181.770 ;
        RECT 142.320 177.770 142.920 181.770 ;
        RECT 145.720 177.770 146.320 181.770 ;
        RECT 111.850 177.430 112.190 177.770 ;
        RECT 111.855 177.355 112.185 177.430 ;
        RECT 139.070 176.850 139.370 177.770 ;
        RECT 142.450 177.440 142.790 177.770 ;
        RECT 142.455 177.255 142.785 177.440 ;
        RECT 148.120 177.395 148.420 195.430 ;
        RECT 149.255 187.620 149.585 187.950 ;
        RECT 149.270 181.770 149.570 187.620 ;
        RECT 152.655 184.860 152.985 185.190 ;
        RECT 152.670 181.770 152.970 184.860 ;
        RECT 149.120 177.770 149.720 181.770 ;
        RECT 152.520 177.770 153.120 181.770 ;
        RECT 149.255 177.725 149.585 177.770 ;
        RECT 148.105 177.065 148.435 177.395 ;
        RECT 144.655 176.850 144.985 176.865 ;
        RECT 117.980 176.485 118.880 176.640 ;
        RECT 137.800 176.485 138.700 176.620 ;
        RECT 139.070 176.550 144.985 176.850 ;
        RECT 144.655 176.535 144.985 176.550 ;
        RECT 103.865 176.250 138.700 176.485 ;
        RECT 157.570 176.250 158.470 176.600 ;
        RECT 103.865 176.230 144.350 176.250 ;
        RECT 145.300 176.230 158.470 176.250 ;
        RECT 103.865 175.110 158.470 176.230 ;
        RECT 103.865 174.875 138.700 175.110 ;
        RECT 117.980 174.620 118.880 174.875 ;
        RECT 137.800 174.600 138.700 174.875 ;
        RECT 157.570 174.580 158.470 175.110 ;
        RECT 28.910 173.995 30.490 174.325 ;
        RECT 70.025 173.290 70.355 173.305 ;
        RECT 73.245 173.290 73.575 173.305 ;
        RECT 70.025 172.990 73.575 173.290 ;
        RECT 70.025 172.975 70.355 172.990 ;
        RECT 73.245 172.975 73.575 172.990 ;
        RECT 32.210 171.275 33.790 171.605 ;
        RECT 108.820 169.350 109.400 169.400 ;
        RECT 128.680 169.350 129.260 169.390 ;
        RECT 148.880 169.350 149.460 169.370 ;
        RECT 28.910 168.555 30.490 168.885 ;
        RECT 108.800 168.720 149.480 169.350 ;
        RECT 32.210 165.835 33.790 166.165 ;
        RECT 28.910 163.115 30.490 163.445 ;
        RECT 32.210 160.395 33.790 160.725 ;
        RECT 28.910 157.675 30.490 158.005 ;
        RECT 32.210 154.955 33.790 155.285 ;
        RECT 128.680 154.340 129.260 154.430 ;
        RECT 139.065 154.340 139.695 168.720 ;
        RECT 108.740 153.710 149.500 154.340 ;
        RECT 108.790 153.690 109.370 153.710 ;
        RECT 28.910 152.235 30.490 152.565 ;
        RECT 32.210 149.515 33.790 149.845 ;
        RECT 28.910 146.795 30.490 147.125 ;
        RECT 32.210 144.075 33.790 144.405 ;
        RECT 28.910 141.355 30.490 141.685 ;
        RECT 54.385 139.970 54.715 139.985 ;
        RECT 71.865 139.970 72.195 139.985 ;
        RECT 54.385 139.670 72.195 139.970 ;
        RECT 54.385 139.655 54.715 139.670 ;
        RECT 71.865 139.655 72.195 139.670 ;
        RECT 108.790 139.340 109.370 139.370 ;
        RECT 128.680 139.340 129.260 139.360 ;
        RECT 139.065 139.340 139.695 153.710 ;
        RECT 32.210 138.635 33.790 138.965 ;
        RECT 108.790 138.740 149.490 139.340 ;
        RECT 108.810 138.710 149.490 138.740 ;
        RECT 12.065 136.570 12.395 136.585 ;
        RECT 11.850 136.255 12.395 136.570 ;
        RECT 11.850 136.040 12.150 136.255 ;
        RECT 7.860 135.590 12.150 136.040 ;
        RECT 28.910 135.915 30.490 136.245 ;
        RECT 7.860 135.440 11.860 135.590 ;
        RECT 32.210 133.195 33.790 133.525 ;
        RECT 28.910 130.475 30.490 130.805 ;
        RECT 32.210 127.755 33.790 128.085 ;
        RECT 28.910 125.035 30.490 125.365 ;
        RECT 128.610 124.380 129.190 124.420 ;
        RECT 139.065 124.380 139.695 138.710 ;
        RECT 148.830 138.670 149.410 138.710 ;
        RECT 108.800 124.370 149.530 124.380 ;
        RECT 108.790 123.750 149.530 124.370 ;
        RECT 108.790 123.740 109.370 123.750 ;
        RECT 32.210 122.315 33.790 122.645 ;
        RECT 28.910 119.595 30.490 119.925 ;
        RECT 32.210 116.875 33.790 117.205 ;
        RECT 12.065 116.170 12.395 116.185 ;
        RECT 11.850 115.855 12.395 116.170 ;
        RECT 11.850 115.640 12.150 115.855 ;
        RECT 7.860 115.190 12.150 115.640 ;
        RECT 89.805 115.490 90.135 115.505 ;
        RECT 93.860 115.490 97.860 115.640 ;
        RECT 89.805 115.190 97.860 115.490 ;
        RECT 7.860 115.040 11.860 115.190 ;
        RECT 89.805 115.175 90.135 115.190 ;
        RECT 93.860 115.040 97.860 115.190 ;
        RECT 28.910 114.155 30.490 114.485 ;
        RECT 12.065 112.770 12.395 112.785 ;
        RECT 11.850 112.455 12.395 112.770 ;
        RECT 11.850 112.240 12.150 112.455 ;
        RECT 7.860 111.790 12.150 112.240 ;
        RECT 89.805 112.090 90.135 112.105 ;
        RECT 93.860 112.090 97.860 112.240 ;
        RECT 89.805 111.790 97.860 112.090 ;
        RECT 7.860 111.640 11.860 111.790 ;
        RECT 89.805 111.775 90.135 111.790 ;
        RECT 32.210 111.435 33.790 111.765 ;
        RECT 93.860 111.640 97.860 111.790 ;
        RECT 128.730 109.330 129.310 109.390 ;
        RECT 139.065 109.330 139.695 123.750 ;
        RECT 148.910 109.330 149.490 109.420 ;
        RECT 7.860 108.690 11.860 108.840 ;
        RECT 28.910 108.715 30.490 109.045 ;
        RECT 108.740 108.790 149.490 109.330 ;
        RECT 14.365 108.690 14.695 108.705 ;
        RECT 108.740 108.700 149.420 108.790 ;
        RECT 7.860 108.390 14.695 108.690 ;
        RECT 7.860 108.240 11.860 108.390 ;
        RECT 14.365 108.375 14.695 108.390 ;
        RECT 32.210 105.995 33.790 106.325 ;
        RECT 7.860 105.290 11.860 105.440 ;
        RECT 23.105 105.290 23.435 105.305 ;
        RECT 7.860 104.990 23.435 105.290 ;
        RECT 7.860 104.840 11.860 104.990 ;
        RECT 23.105 104.975 23.435 104.990 ;
        RECT 28.910 103.275 30.490 103.605 ;
        RECT 12.065 102.570 12.395 102.585 ;
        RECT 11.850 102.255 12.395 102.570 ;
        RECT 139.065 102.305 139.695 108.700 ;
        RECT 11.850 102.040 12.150 102.255 ;
        RECT 7.860 101.590 12.150 102.040 ;
        RECT 139.065 101.675 158.365 102.305 ;
        RECT 7.860 101.440 11.860 101.590 ;
        RECT 32.210 100.555 33.790 100.885 ;
        RECT 73.245 99.170 73.575 99.185 ;
        RECT 79.225 99.170 79.555 99.185 ;
        RECT 73.245 98.870 79.555 99.170 ;
        RECT 73.245 98.855 73.575 98.870 ;
        RECT 79.225 98.855 79.555 98.870 ;
        RECT 28.910 97.835 30.490 98.165 ;
        RECT 157.735 96.565 158.365 101.675 ;
        RECT 32.210 95.115 33.790 95.445 ;
        RECT 66.805 95.090 67.135 95.105 ;
        RECT 75.545 95.090 75.875 95.105 ;
        RECT 66.805 94.790 75.875 95.090 ;
        RECT 66.805 94.775 67.135 94.790 ;
        RECT 75.545 94.775 75.875 94.790 ;
        RECT 28.910 92.395 30.490 92.725 ;
        RECT 32.210 89.675 33.790 90.005 ;
        RECT 89.805 88.290 90.135 88.305 ;
        RECT 93.860 88.290 97.860 88.440 ;
        RECT 89.805 87.990 97.860 88.290 ;
        RECT 89.805 87.975 90.135 87.990 ;
        RECT 93.860 87.840 97.860 87.990 ;
        RECT 28.910 86.955 30.490 87.285 ;
        RECT 32.210 84.235 33.790 84.565 ;
        RECT 121.560 83.790 122.110 84.300 ;
        RECT 133.745 83.010 134.095 83.035 ;
        RECT 133.745 82.710 137.340 83.010 ;
        RECT 133.745 82.685 134.095 82.710 ;
        RECT 70.025 82.170 70.355 82.185 ;
        RECT 72.785 82.170 73.115 82.185 ;
        RECT 70.025 81.870 73.115 82.170 ;
        RECT 70.025 81.855 70.355 81.870 ;
        RECT 72.785 81.855 73.115 81.870 ;
        RECT 28.910 81.515 30.490 81.845 ;
        RECT 89.805 81.490 90.135 81.505 ;
        RECT 93.860 81.490 97.860 81.640 ;
        RECT 89.805 81.190 97.860 81.490 ;
        RECT 89.805 81.175 90.135 81.190 ;
        RECT 93.860 81.040 97.860 81.190 ;
        RECT 32.210 78.795 33.790 79.125 ;
        RECT 137.040 78.825 137.340 82.710 ;
        RECT 73.705 78.770 74.035 78.785 ;
        RECT 75.545 78.770 75.875 78.785 ;
        RECT 73.705 78.470 75.875 78.770 ;
        RECT 137.025 78.495 137.355 78.825 ;
        RECT 73.705 78.455 74.035 78.470 ;
        RECT 75.545 78.455 75.875 78.470 ;
        RECT 139.240 78.300 139.890 78.860 ;
        RECT 28.910 76.075 30.490 76.405 ;
        RECT 89.805 74.690 90.135 74.705 ;
        RECT 93.860 74.690 97.860 74.840 ;
        RECT 89.805 74.390 97.860 74.690 ;
        RECT 89.805 74.375 90.135 74.390 ;
        RECT 93.860 74.240 97.860 74.390 ;
        RECT 32.210 73.355 33.790 73.685 ;
        RECT 68.645 72.650 68.975 72.665 ;
        RECT 75.085 72.650 75.415 72.665 ;
        RECT 68.645 72.350 75.415 72.650 ;
        RECT 68.645 72.335 68.975 72.350 ;
        RECT 75.085 72.335 75.415 72.350 ;
        RECT 69.105 71.970 69.435 71.985 ;
        RECT 72.325 71.970 72.655 71.985 ;
        RECT 69.105 71.670 72.655 71.970 ;
        RECT 69.105 71.655 69.435 71.670 ;
        RECT 72.325 71.655 72.655 71.670 ;
        RECT 90.265 71.290 90.595 71.305 ;
        RECT 93.860 71.290 97.860 71.440 ;
        RECT 90.265 70.990 97.860 71.290 ;
        RECT 90.265 70.975 90.595 70.990 ;
        RECT 28.910 70.635 30.490 70.965 ;
        RECT 93.860 70.840 97.860 70.990 ;
        RECT 7.860 67.890 11.860 68.040 ;
        RECT 32.210 67.915 33.790 68.245 ;
        RECT 14.365 67.890 14.695 67.905 ;
        RECT 7.860 67.590 14.695 67.890 ;
        RECT 7.860 67.440 11.860 67.590 ;
        RECT 14.365 67.575 14.695 67.590 ;
        RECT 85.665 67.890 85.995 67.905 ;
        RECT 93.860 67.890 97.860 68.040 ;
        RECT 85.665 67.590 97.860 67.890 ;
        RECT 85.665 67.575 85.995 67.590 ;
        RECT 93.860 67.440 97.860 67.590 ;
        RECT 43.805 65.860 44.135 65.865 ;
        RECT 43.805 65.850 44.390 65.860 ;
        RECT 43.805 65.550 44.590 65.850 ;
        RECT 43.805 65.540 44.390 65.550 ;
        RECT 43.805 65.535 44.135 65.540 ;
        RECT 28.910 65.195 30.490 65.525 ;
        RECT 7.860 64.490 11.860 64.640 ;
        RECT 89.805 64.490 90.135 64.505 ;
        RECT 93.860 64.490 97.860 64.640 ;
        RECT 7.860 64.040 12.150 64.490 ;
        RECT 89.805 64.190 97.860 64.490 ;
        RECT 89.805 64.175 90.135 64.190 ;
        RECT 93.860 64.040 97.860 64.190 ;
        RECT 11.850 63.825 12.150 64.040 ;
        RECT 11.850 63.510 12.395 63.825 ;
        RECT 12.065 63.495 12.395 63.510 ;
        RECT 32.210 62.475 33.790 62.805 ;
        RECT 7.860 61.090 11.860 61.240 ;
        RECT 13.445 61.090 13.775 61.105 ;
        RECT 7.860 60.790 13.775 61.090 ;
        RECT 7.860 60.640 11.860 60.790 ;
        RECT 13.445 60.775 13.775 60.790 ;
        RECT 89.805 61.090 90.135 61.105 ;
        RECT 93.860 61.090 97.860 61.240 ;
        RECT 89.805 60.790 97.860 61.090 ;
        RECT 89.805 60.775 90.135 60.790 ;
        RECT 93.860 60.640 97.860 60.790 ;
        RECT 67.725 60.410 68.055 60.425 ;
        RECT 72.785 60.410 73.115 60.425 ;
        RECT 67.725 60.110 73.115 60.410 ;
        RECT 67.725 60.095 68.055 60.110 ;
        RECT 72.785 60.095 73.115 60.110 ;
        RECT 28.910 59.755 30.490 60.085 ;
        RECT 7.860 57.690 11.860 57.840 ;
        RECT 17.125 57.690 17.455 57.705 ;
        RECT 7.860 57.390 17.455 57.690 ;
        RECT 7.860 57.240 11.860 57.390 ;
        RECT 17.125 57.375 17.455 57.390 ;
        RECT 32.210 57.035 33.790 57.365 ;
        RECT 20.805 56.330 21.135 56.345 ;
        RECT 21.725 56.330 22.055 56.345 ;
        RECT 20.805 56.030 22.055 56.330 ;
        RECT 20.805 56.015 21.135 56.030 ;
        RECT 21.725 56.015 22.055 56.030 ;
        RECT 7.860 54.290 11.860 54.440 ;
        RECT 28.910 54.315 30.490 54.645 ;
        RECT 14.365 54.290 14.695 54.305 ;
        RECT 7.860 53.990 14.695 54.290 ;
        RECT 7.860 53.840 11.860 53.990 ;
        RECT 14.365 53.975 14.695 53.990 ;
        RECT 89.805 54.290 90.135 54.305 ;
        RECT 93.860 54.290 97.860 54.440 ;
        RECT 89.805 53.990 97.860 54.290 ;
        RECT 89.805 53.975 90.135 53.990 ;
        RECT 93.860 53.840 97.860 53.990 ;
        RECT 32.210 51.595 33.790 51.925 ;
        RECT 7.860 50.890 11.860 51.040 ;
        RECT 12.985 50.890 13.315 50.905 ;
        RECT 7.860 50.590 13.315 50.890 ;
        RECT 7.860 50.440 11.860 50.590 ;
        RECT 12.985 50.575 13.315 50.590 ;
        RECT 28.910 48.875 30.490 49.205 ;
        RECT 12.065 48.170 12.395 48.185 ;
        RECT 11.850 47.855 12.395 48.170 ;
        RECT 11.850 47.640 12.150 47.855 ;
        RECT 7.860 47.190 12.150 47.640 ;
        RECT 31.130 47.490 31.510 47.500 ;
        RECT 33.685 47.490 34.015 47.505 ;
        RECT 31.130 47.190 34.015 47.490 ;
        RECT 7.860 47.040 11.860 47.190 ;
        RECT 31.130 47.180 31.510 47.190 ;
        RECT 33.685 47.175 34.015 47.190 ;
        RECT 32.210 46.155 33.790 46.485 ;
        RECT 7.860 44.090 11.860 44.240 ;
        RECT 21.725 44.090 22.055 44.105 ;
        RECT 7.860 43.790 22.055 44.090 ;
        RECT 7.860 43.640 11.860 43.790 ;
        RECT 21.725 43.775 22.055 43.790 ;
        RECT 90.725 44.090 91.055 44.105 ;
        RECT 93.860 44.090 97.860 44.240 ;
        RECT 90.725 43.790 97.860 44.090 ;
        RECT 90.725 43.775 91.055 43.790 ;
        RECT 28.910 43.435 30.490 43.765 ;
        RECT 93.860 43.640 97.860 43.790 ;
        RECT 7.860 40.690 11.860 40.840 ;
        RECT 32.210 40.715 33.790 41.045 ;
        RECT 22.645 40.690 22.975 40.705 ;
        RECT 7.860 40.390 22.975 40.690 ;
        RECT 7.860 40.240 11.860 40.390 ;
        RECT 22.645 40.375 22.975 40.390 ;
        RECT 19.885 39.330 20.215 39.345 ;
        RECT 49.785 39.330 50.115 39.345 ;
        RECT 19.885 39.030 50.115 39.330 ;
        RECT 19.885 39.015 20.215 39.030 ;
        RECT 49.785 39.015 50.115 39.030 ;
        RECT 28.910 37.995 30.490 38.325 ;
        RECT 32.210 35.275 33.790 35.605 ;
        RECT 77.385 34.570 77.715 34.585 ;
        RECT 81.985 34.570 82.315 34.585 ;
        RECT 77.385 34.270 82.315 34.570 ;
        RECT 77.385 34.255 77.715 34.270 ;
        RECT 81.985 34.255 82.315 34.270 ;
        RECT 28.910 32.555 30.490 32.885 ;
        RECT 90.725 30.490 91.055 30.505 ;
        RECT 93.860 30.490 97.860 30.640 ;
        RECT 90.725 30.190 97.860 30.490 ;
        RECT 90.725 30.175 91.055 30.190 ;
        RECT 32.210 29.835 33.790 30.165 ;
        RECT 93.860 30.040 97.860 30.190 ;
        RECT 28.910 27.115 30.490 27.445 ;
        RECT 32.210 24.395 33.790 24.725 ;
        RECT 25.405 23.690 25.735 23.705 ;
        RECT 40.585 23.690 40.915 23.705 ;
        RECT 47.025 23.690 47.355 23.705 ;
        RECT 25.405 23.390 47.355 23.690 ;
        RECT 25.405 23.375 25.735 23.390 ;
        RECT 40.585 23.375 40.915 23.390 ;
        RECT 47.025 23.375 47.355 23.390 ;
        RECT 44.010 23.010 44.390 23.020 ;
        RECT 65.425 23.010 65.755 23.025 ;
        RECT 44.010 22.710 65.755 23.010 ;
        RECT 44.010 22.700 44.390 22.710 ;
        RECT 65.425 22.695 65.755 22.710 ;
        RECT 28.910 21.675 30.490 22.005 ;
        RECT 29.085 20.970 29.415 20.985 ;
        RECT 31.130 20.970 31.510 20.980 ;
        RECT 44.265 20.970 44.595 20.985 ;
        RECT 29.085 20.670 44.595 20.970 ;
        RECT 29.085 20.655 29.415 20.670 ;
        RECT 31.130 20.660 31.510 20.670 ;
        RECT 44.265 20.655 44.595 20.670 ;
        RECT 32.210 18.955 33.790 19.285 ;
        RECT 28.910 16.235 30.490 16.565 ;
        RECT 32.210 13.515 33.790 13.845 ;
      LAYER met4 ;
        RECT 63.685 224.985 63.790 225.315 ;
        RECT 66.515 224.965 66.550 225.295 ;
        RECT 69.235 225.005 69.310 225.335 ;
        RECT 72.370 225.045 72.435 225.375 ;
        RECT 74.800 224.975 74.830 225.305 ;
        RECT 77.565 224.995 77.590 225.325 ;
        RECT 77.890 224.995 77.895 225.325 ;
        RECT 80.305 224.915 80.350 225.245 ;
        RECT 83.410 224.945 83.445 225.275 ;
        RECT 85.815 225.025 85.870 225.355 ;
        RECT 88.585 224.955 88.630 225.285 ;
        RECT 91.310 224.985 91.390 225.315 ;
        RECT 93.985 225.015 94.150 225.345 ;
        RECT 118.795 224.760 118.990 225.215 ;
        RECT 119.290 224.760 119.455 225.215 ;
        RECT 121.530 224.805 121.750 225.455 ;
        RECT 122.050 224.805 122.190 225.455 ;
        RECT 124.275 224.945 124.510 225.595 ;
        RECT 124.810 224.945 124.935 225.595 ;
        RECT 127.145 224.965 127.270 225.615 ;
        RECT 127.570 224.965 127.805 225.615 ;
        RECT 129.605 224.960 130.030 225.610 ;
        RECT 133.090 224.945 133.645 225.595 ;
        RECT 134.915 225.075 135.550 225.725 ;
        RECT 137.630 224.895 138.310 225.575 ;
        RECT 142.455 225.400 142.785 225.415 ;
        RECT 142.455 225.100 143.830 225.400 ;
        RECT 142.455 225.085 142.785 225.100 ;
        RECT 118.795 224.565 119.455 224.760 ;
        RECT 112.120 203.770 147.960 203.775 ;
        RECT 98.780 202.180 147.960 203.770 ;
        RECT 112.120 202.175 147.960 202.180 ;
        RECT 6.000 198.890 6.020 200.480 ;
        RECT 28.900 13.440 30.500 201.600 ;
        RECT 31.155 47.175 31.485 47.505 ;
        RECT 31.170 20.985 31.470 47.175 ;
        RECT 31.155 20.655 31.485 20.985 ;
        RECT 32.200 13.440 33.800 201.600 ;
        RECT 98.780 200.475 113.500 200.480 ;
        RECT 98.780 198.890 147.960 200.475 ;
        RECT 112.120 198.875 147.960 198.890 ;
        RECT 157.730 96.590 158.370 97.230 ;
        RECT 121.645 83.855 139.745 84.245 ;
        RECT 139.355 78.860 139.745 83.855 ;
        RECT 139.240 78.755 139.890 78.860 ;
        RECT 157.735 78.755 158.365 96.590 ;
        RECT 139.240 78.365 158.365 78.755 ;
        RECT 139.240 78.300 139.890 78.365 ;
        RECT 44.035 65.535 44.365 65.865 ;
        RECT 44.050 23.025 44.350 65.535 ;
        RECT 44.035 22.695 44.365 23.025 ;
        RECT 157.735 1.065 158.365 78.365 ;
        RECT 16.570 1.000 17.470 1.040 ;
        RECT 35.890 1.000 36.790 1.040 ;
        RECT 55.210 1.000 56.110 1.030 ;
        RECT 132.490 1.000 133.390 1.010 ;
        RECT 152.045 1.000 158.365 1.065 ;
        RECT 152.710 0.435 158.365 1.000 ;
  END
END tt_um_tim2305_adc_dac
END LIBRARY

