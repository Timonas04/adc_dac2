VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_tim2305_adc_dac
  CLASS BLOCK ;
  FOREIGN tt_um_tim2305_adc_dac ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER met1 ;
        RECT 147.680 220.250 147.940 220.570 ;
        RECT 147.240 219.710 147.500 220.030 ;
        RECT 146.840 219.250 147.160 219.510 ;
        RECT 146.310 218.730 146.570 219.050 ;
        RECT 146.370 214.650 146.510 218.730 ;
        RECT 146.930 214.650 147.070 219.250 ;
        RECT 147.300 214.650 147.440 219.710 ;
        RECT 147.740 214.650 147.880 220.250 ;
      LAYER met2 ;
        RECT 69.275 221.420 69.665 221.500 ;
        RECT 69.275 221.280 73.200 221.420 ;
        RECT 69.275 221.200 69.665 221.280 ;
        RECT 73.060 221.240 73.200 221.280 ;
        RECT 73.060 221.100 125.130 221.240 ;
        RECT 71.965 220.960 72.355 221.040 ;
        RECT 71.965 220.820 124.490 220.960 ;
        RECT 71.965 220.740 72.355 220.820 ;
        RECT 74.755 220.560 75.145 220.620 ;
        RECT 123.555 220.560 123.925 220.610 ;
        RECT 74.755 220.380 123.925 220.560 ;
        RECT 74.755 220.320 75.145 220.380 ;
        RECT 123.555 220.330 123.925 220.380 ;
        RECT 124.350 220.370 124.490 220.820 ;
        RECT 124.990 220.650 125.130 221.100 ;
        RECT 124.990 220.510 138.900 220.650 ;
        RECT 138.760 220.480 138.900 220.510 ;
        RECT 147.650 220.480 147.970 220.540 ;
        RECT 124.350 220.230 138.300 220.370 ;
        RECT 138.760 220.340 147.970 220.480 ;
        RECT 147.650 220.280 147.970 220.340 ;
        RECT 80.265 219.985 80.655 220.040 ;
        RECT 137.155 219.985 137.525 220.030 ;
        RECT 80.265 219.830 137.525 219.985 ;
        RECT 80.265 219.795 82.855 219.830 ;
        RECT 83.525 219.795 137.525 219.830 ;
        RECT 138.160 219.940 138.300 220.230 ;
        RECT 147.210 219.940 147.530 220.000 ;
        RECT 138.160 219.800 147.530 219.940 ;
        RECT 80.265 219.740 80.655 219.795 ;
        RECT 137.155 219.750 137.525 219.795 ;
        RECT 147.210 219.740 147.530 219.800 ;
        RECT 82.995 219.610 83.385 219.690 ;
        RECT 82.995 219.470 115.180 219.610 ;
        RECT 82.995 219.390 83.385 219.470 ;
        RECT 115.040 219.450 115.180 219.470 ;
        RECT 146.870 219.450 147.130 219.540 ;
        RECT 115.040 219.310 147.130 219.450 ;
        RECT 85.765 219.220 86.155 219.255 ;
        RECT 146.870 219.220 147.130 219.310 ;
        RECT 85.765 218.990 114.140 219.220 ;
        RECT 85.765 218.955 86.155 218.990 ;
        RECT 146.280 218.960 146.600 219.020 ;
        RECT 115.000 218.820 146.600 218.960 ;
        RECT 94.095 218.740 94.485 218.820 ;
        RECT 115.000 218.740 115.140 218.820 ;
        RECT 146.280 218.760 146.600 218.820 ;
        RECT 94.095 218.600 115.140 218.740 ;
        RECT 91.365 218.415 91.665 218.530 ;
        RECT 94.095 218.520 94.485 218.600 ;
        RECT 115.680 218.415 128.540 218.565 ;
        RECT 143.865 218.510 144.255 218.585 ;
        RECT 91.365 218.360 93.960 218.415 ;
        RECT 94.620 218.400 128.540 218.415 ;
        RECT 94.620 218.360 115.845 218.400 ;
        RECT 91.365 218.250 115.845 218.360 ;
        RECT 141.320 218.355 144.255 218.510 ;
        RECT 143.865 218.285 144.255 218.355 ;
        RECT 91.365 218.140 91.665 218.250 ;
        RECT 93.840 218.220 94.750 218.250 ;
        RECT 88.505 218.010 88.895 218.090 ;
        RECT 88.505 217.990 91.210 218.010 ;
        RECT 91.820 217.990 110.010 218.010 ;
        RECT 88.505 217.870 110.010 217.990 ;
        RECT 88.505 217.790 88.895 217.870 ;
        RECT 90.980 217.830 91.980 217.870 ;
        RECT 77.530 217.660 77.830 217.785 ;
        RECT 77.530 217.650 88.365 217.660 ;
        RECT 89.035 217.650 109.630 217.660 ;
        RECT 77.530 217.520 109.630 217.650 ;
        RECT 77.530 217.395 77.830 217.520 ;
        RECT 88.280 217.510 89.120 217.520 ;
        RECT 66.425 217.260 66.815 217.340 ;
        RECT 66.425 217.250 77.370 217.260 ;
        RECT 77.980 217.250 109.010 217.260 ;
        RECT 66.425 217.120 109.010 217.250 ;
        RECT 66.425 217.040 66.815 217.120 ;
        RECT 77.250 217.110 78.140 217.120 ;
        RECT 63.785 216.900 64.175 216.980 ;
        RECT 63.785 216.760 108.550 216.900 ;
        RECT 63.785 216.680 64.175 216.760 ;
        RECT 108.410 214.650 108.550 216.760 ;
        RECT 108.870 214.650 109.010 217.120 ;
        RECT 109.490 214.650 109.630 217.520 ;
        RECT 109.870 214.650 110.010 217.870 ;
      LAYER met3 ;
        RECT 63.820 225.030 64.140 225.410 ;
        RECT 63.830 217.005 64.130 225.030 ;
        RECT 66.460 224.940 66.780 225.320 ;
        RECT 69.310 225.110 69.630 225.490 ;
        RECT 66.470 217.365 66.770 224.940 ;
        RECT 69.320 221.525 69.620 225.110 ;
        RECT 72.000 224.870 72.320 225.250 ;
        RECT 74.790 224.920 75.110 225.300 ;
        RECT 69.295 221.175 69.645 221.525 ;
        RECT 72.010 221.065 72.310 224.870 ;
        RECT 71.985 220.715 72.335 221.065 ;
        RECT 74.800 220.645 75.100 224.920 ;
        RECT 77.520 224.730 77.840 225.110 ;
        RECT 80.300 224.900 80.620 225.280 ;
        RECT 74.775 220.295 75.125 220.645 ;
        RECT 77.530 217.765 77.830 224.730 ;
        RECT 80.310 220.065 80.610 224.900 ;
        RECT 83.030 224.730 83.350 225.110 ;
        RECT 85.800 224.890 86.120 225.270 ;
        RECT 88.540 224.890 88.860 225.270 ;
        RECT 80.285 219.715 80.635 220.065 ;
        RECT 83.040 219.715 83.340 224.730 ;
        RECT 83.015 219.365 83.365 219.715 ;
        RECT 85.810 219.280 86.110 224.890 ;
        RECT 85.785 218.930 86.135 219.280 ;
        RECT 88.550 218.115 88.850 224.890 ;
        RECT 91.355 224.810 91.675 225.190 ;
        RECT 91.365 218.510 91.665 224.810 ;
        RECT 94.130 224.790 94.450 225.170 ;
        RECT 143.900 225.090 144.220 225.470 ;
        RECT 94.140 218.845 94.440 224.790 ;
        RECT 123.575 220.305 123.905 220.635 ;
        RECT 91.340 218.160 91.690 218.510 ;
        RECT 94.115 218.495 94.465 218.845 ;
        RECT 123.590 218.540 123.890 220.305 ;
        RECT 137.175 219.725 137.505 220.055 ;
        RECT 137.190 218.280 137.490 219.725 ;
        RECT 143.910 218.610 144.210 225.090 ;
        RECT 143.885 218.260 144.235 218.610 ;
        RECT 88.525 217.765 88.875 218.115 ;
        RECT 77.505 217.415 77.855 217.765 ;
        RECT 66.445 217.015 66.795 217.365 ;
        RECT 63.805 216.655 64.155 217.005 ;
        RECT 8.565 202.460 10.155 202.485 ;
        RECT 1.070 200.860 10.160 202.460 ;
        RECT 8.565 200.835 10.155 200.860 ;
      LAYER met4 ;
        RECT 64.090 225.055 64.145 225.385 ;
        RECT 66.455 224.965 66.550 225.295 ;
        RECT 69.305 225.135 69.310 225.465 ;
        RECT 69.610 225.135 69.635 225.465 ;
        RECT 71.995 224.895 72.070 225.225 ;
        RECT 74.785 224.945 74.830 225.275 ;
        RECT 77.515 224.760 77.590 225.085 ;
        RECT 80.295 224.925 80.350 225.255 ;
        RECT 83.025 224.760 83.110 225.085 ;
        RECT 85.795 224.915 85.870 225.245 ;
        RECT 88.535 224.915 88.630 225.245 ;
        RECT 91.350 224.835 91.390 225.165 ;
        RECT 94.125 224.815 94.150 225.145 ;
        RECT 94.450 224.815 94.455 225.145 ;
        RECT 144.130 225.115 144.225 225.445 ;
        RECT 77.515 224.755 77.845 224.760 ;
        RECT 83.025 224.755 83.355 224.760 ;
        RECT 8.560 200.860 13.900 202.460 ;
        RECT 6.000 197.560 13.900 199.160 ;
        RECT 151.950 1.000 152.575 9.470 ;
  END
END tt_um_tim2305_adc_dac
END LIBRARY

