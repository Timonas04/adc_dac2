magic
tech sky130A
magscale 1 2
timestamp 1730882523
<< viali >>
rect 7941 33065 7975 33099
rect 11713 33065 11747 33099
rect 13737 33065 13771 33099
rect 11161 32997 11195 33031
rect 8125 32861 8159 32895
rect 10609 32861 10643 32895
rect 10977 32861 11011 32895
rect 11345 32861 11379 32895
rect 11529 32861 11563 32895
rect 12173 32861 12207 32895
rect 12725 32861 12759 32895
rect 13921 32861 13955 32895
rect 15025 32861 15059 32895
rect 15577 32861 15611 32895
rect 15945 32861 15979 32895
rect 12449 32793 12483 32827
rect 12633 32793 12667 32827
rect 12909 32793 12943 32827
rect 13093 32793 13127 32827
rect 13369 32793 13403 32827
rect 13553 32793 13587 32827
rect 14105 32793 14139 32827
rect 14289 32793 14323 32827
rect 14565 32793 14599 32827
rect 14749 32793 14783 32827
rect 15209 32793 15243 32827
rect 15761 32793 15795 32827
rect 15853 32793 15887 32827
rect 10425 32725 10459 32759
rect 10793 32725 10827 32759
rect 11989 32725 12023 32759
rect 12265 32725 12299 32759
rect 13185 32725 13219 32759
rect 14473 32725 14507 32759
rect 14933 32725 14967 32759
rect 15393 32725 15427 32759
rect 16129 32725 16163 32759
rect 12449 32521 12483 32555
rect 15853 32453 15887 32487
rect 6929 32385 6963 32419
rect 7205 32385 7239 32419
rect 7389 32385 7423 32419
rect 8953 32385 8987 32419
rect 9137 32385 9171 32419
rect 10609 32385 10643 32419
rect 13562 32385 13596 32419
rect 14381 32385 14415 32419
rect 14473 32385 14507 32419
rect 14565 32385 14599 32419
rect 14749 32385 14783 32419
rect 15117 32385 15151 32419
rect 15209 32385 15243 32419
rect 15301 32385 15335 32419
rect 15485 32385 15519 32419
rect 15761 32385 15795 32419
rect 15945 32385 15979 32419
rect 16129 32385 16163 32419
rect 10793 32317 10827 32351
rect 12081 32317 12115 32351
rect 13829 32317 13863 32351
rect 7021 32249 7055 32283
rect 7113 32249 7147 32283
rect 10425 32249 10459 32283
rect 11529 32249 11563 32283
rect 6745 32181 6779 32215
rect 9045 32181 9079 32215
rect 11345 32181 11379 32215
rect 14105 32181 14139 32215
rect 14841 32181 14875 32215
rect 15577 32181 15611 32215
rect 7849 31977 7883 32011
rect 8953 31977 8987 32011
rect 12173 31977 12207 32011
rect 13829 31977 13863 32011
rect 15485 31977 15519 32011
rect 11069 31909 11103 31943
rect 11161 31909 11195 31943
rect 16221 31909 16255 31943
rect 8401 31841 8435 31875
rect 11621 31841 11655 31875
rect 11713 31841 11747 31875
rect 6469 31773 6503 31807
rect 8125 31773 8159 31807
rect 8585 31773 8619 31807
rect 8677 31773 8711 31807
rect 9505 31773 9539 31807
rect 9689 31773 9723 31807
rect 9956 31773 9990 31807
rect 13553 31773 13587 31807
rect 13645 31773 13679 31807
rect 14105 31773 14139 31807
rect 15669 31773 15703 31807
rect 15853 31773 15887 31807
rect 16037 31773 16071 31807
rect 6736 31705 6770 31739
rect 8309 31705 8343 31739
rect 13286 31705 13320 31739
rect 14372 31705 14406 31739
rect 15945 31705 15979 31739
rect 7941 31637 7975 31671
rect 8401 31637 8435 31671
rect 11529 31637 11563 31671
rect 7481 31433 7515 31467
rect 11069 31433 11103 31467
rect 14933 31433 14967 31467
rect 8125 31365 8159 31399
rect 15025 31365 15059 31399
rect 7757 31297 7791 31331
rect 8484 31297 8518 31331
rect 9689 31297 9723 31331
rect 9956 31297 9990 31331
rect 12642 31297 12676 31331
rect 12909 31297 12943 31331
rect 13001 31297 13035 31331
rect 13369 31297 13403 31331
rect 13553 31297 13587 31331
rect 13820 31297 13854 31331
rect 15209 31297 15243 31331
rect 16313 31297 16347 31331
rect 7297 31229 7331 31263
rect 7665 31229 7699 31263
rect 8033 31229 8067 31263
rect 8217 31229 8251 31263
rect 16037 31229 16071 31263
rect 6745 31093 6779 31127
rect 9597 31093 9631 31127
rect 11529 31093 11563 31127
rect 15393 31093 15427 31127
rect 6101 30889 6135 30923
rect 8953 30889 8987 30923
rect 9873 30889 9907 30923
rect 10149 30889 10183 30923
rect 16313 30889 16347 30923
rect 12449 30821 12483 30855
rect 8309 30753 8343 30787
rect 9965 30753 9999 30787
rect 10701 30753 10735 30787
rect 10977 30753 11011 30787
rect 13001 30753 13035 30787
rect 13829 30753 13863 30787
rect 7481 30685 7515 30719
rect 7665 30685 7699 30719
rect 7757 30685 7791 30719
rect 7941 30685 7975 30719
rect 8217 30685 8251 30719
rect 8401 30685 8435 30719
rect 8493 30685 8527 30719
rect 8677 30685 8711 30719
rect 9137 30685 9171 30719
rect 9229 30685 9263 30719
rect 9413 30685 9447 30719
rect 9505 30685 9539 30719
rect 9781 30685 9815 30719
rect 10517 30685 10551 30719
rect 14381 30685 14415 30719
rect 14473 30685 14507 30719
rect 14565 30685 14599 30719
rect 14749 30685 14783 30719
rect 14933 30685 14967 30719
rect 7214 30617 7248 30651
rect 10057 30617 10091 30651
rect 10609 30617 10643 30651
rect 11244 30617 11278 30651
rect 12817 30617 12851 30651
rect 14105 30617 14139 30651
rect 15178 30617 15212 30651
rect 8033 30549 8067 30583
rect 9597 30549 9631 30583
rect 12357 30549 12391 30583
rect 12909 30549 12943 30583
rect 13277 30549 13311 30583
rect 6101 30345 6135 30379
rect 9321 30345 9355 30379
rect 11529 30345 11563 30379
rect 11897 30345 11931 30379
rect 12357 30345 12391 30379
rect 12725 30345 12759 30379
rect 16313 30345 16347 30379
rect 6644 30277 6678 30311
rect 8186 30277 8220 30311
rect 9413 30277 9447 30311
rect 10333 30277 10367 30311
rect 13921 30277 13955 30311
rect 5457 30209 5491 30243
rect 5641 30209 5675 30243
rect 5917 30209 5951 30243
rect 6193 30209 6227 30243
rect 6377 30209 6411 30243
rect 7941 30209 7975 30243
rect 9873 30209 9907 30243
rect 13737 30209 13771 30243
rect 14197 30209 14231 30243
rect 14289 30209 14323 30243
rect 14381 30209 14415 30243
rect 14565 30209 14599 30243
rect 14841 30209 14875 30243
rect 14933 30209 14967 30243
rect 15200 30209 15234 30243
rect 9781 30141 9815 30175
rect 10793 30141 10827 30175
rect 11253 30141 11287 30175
rect 11989 30141 12023 30175
rect 12081 30141 12115 30175
rect 12817 30141 12851 30175
rect 13001 30141 13035 30175
rect 10149 30073 10183 30107
rect 10701 30073 10735 30107
rect 10977 30073 11011 30107
rect 14657 30073 14691 30107
rect 5549 30005 5583 30039
rect 5733 30005 5767 30039
rect 7757 30005 7791 30039
rect 9781 30005 9815 30039
rect 10057 30005 10091 30039
rect 10333 30005 10367 30039
rect 13185 30005 13219 30039
rect 6101 29801 6135 29835
rect 7113 29801 7147 29835
rect 9229 29801 9263 29835
rect 9965 29801 9999 29835
rect 10149 29801 10183 29835
rect 10609 29801 10643 29835
rect 14841 29801 14875 29835
rect 15577 29801 15611 29835
rect 6653 29733 6687 29767
rect 10793 29733 10827 29767
rect 11805 29733 11839 29767
rect 6009 29665 6043 29699
rect 7849 29665 7883 29699
rect 8125 29665 8159 29699
rect 11069 29665 11103 29699
rect 12449 29665 12483 29699
rect 13185 29665 13219 29699
rect 6101 29597 6135 29631
rect 6193 29597 6227 29631
rect 6929 29597 6963 29631
rect 7205 29599 7239 29633
rect 8953 29597 8987 29631
rect 9137 29597 9171 29631
rect 9505 29597 9539 29631
rect 9597 29597 9631 29631
rect 9689 29597 9723 29631
rect 9873 29597 9907 29631
rect 10517 29597 10551 29631
rect 11345 29597 11379 29631
rect 11437 29597 11471 29631
rect 11621 29597 11655 29631
rect 11713 29597 11747 29631
rect 12173 29597 12207 29631
rect 13001 29597 13035 29631
rect 14105 29597 14139 29631
rect 14749 29597 14783 29631
rect 15117 29597 15151 29631
rect 15209 29597 15243 29631
rect 15301 29597 15335 29631
rect 15485 29597 15519 29631
rect 15853 29597 15887 29631
rect 15945 29597 15979 29631
rect 16037 29597 16071 29631
rect 16221 29597 16255 29631
rect 6377 29529 6411 29563
rect 11161 29529 11195 29563
rect 12265 29529 12299 29563
rect 13553 29529 13587 29563
rect 13737 29529 13771 29563
rect 5733 29461 5767 29495
rect 6561 29461 6595 29495
rect 7297 29461 7331 29495
rect 8677 29461 8711 29495
rect 9045 29461 9079 29495
rect 10149 29461 10183 29495
rect 12633 29461 12667 29495
rect 13093 29461 13127 29495
rect 13921 29461 13955 29495
rect 6561 29257 6595 29291
rect 9137 29257 9171 29291
rect 10977 29257 11011 29291
rect 11145 29257 11179 29291
rect 13645 29257 13679 29291
rect 16129 29257 16163 29291
rect 11345 29189 11379 29223
rect 12532 29189 12566 29223
rect 6929 29121 6963 29155
rect 7021 29121 7055 29155
rect 8421 29121 8455 29155
rect 8677 29121 8711 29155
rect 8953 29121 8987 29155
rect 9229 29121 9263 29155
rect 9505 29121 9539 29155
rect 9772 29121 9806 29155
rect 14381 29121 14415 29155
rect 14657 29121 14691 29155
rect 14749 29121 14783 29155
rect 14933 29121 14967 29155
rect 15025 29121 15059 29155
rect 15117 29121 15151 29155
rect 15669 29121 15703 29155
rect 15761 29121 15795 29155
rect 15945 29121 15979 29155
rect 16037 29121 16071 29155
rect 16313 29121 16347 29155
rect 6745 29053 6779 29087
rect 6837 29053 6871 29087
rect 8769 29053 8803 29087
rect 12081 29053 12115 29087
rect 12265 29053 12299 29087
rect 7297 28985 7331 29019
rect 10885 28985 10919 29019
rect 15301 28985 15335 29019
rect 11161 28917 11195 28951
rect 11529 28917 11563 28951
rect 13737 28917 13771 28951
rect 14473 28917 14507 28951
rect 15485 28917 15519 28951
rect 6837 28713 6871 28747
rect 7113 28713 7147 28747
rect 9137 28713 9171 28747
rect 9321 28713 9355 28747
rect 10149 28713 10183 28747
rect 13737 28713 13771 28747
rect 16313 28713 16347 28747
rect 8769 28645 8803 28679
rect 9873 28645 9907 28679
rect 8125 28577 8159 28611
rect 10701 28577 10735 28611
rect 14933 28577 14967 28611
rect 6745 28509 6779 28543
rect 7021 28509 7055 28543
rect 7205 28509 7239 28543
rect 8585 28509 8619 28543
rect 8769 28509 8803 28543
rect 10057 28509 10091 28543
rect 10609 28509 10643 28543
rect 11621 28509 11655 28543
rect 12357 28509 12391 28543
rect 14105 28509 14139 28543
rect 14289 28509 14323 28543
rect 14381 28509 14415 28543
rect 14473 28509 14507 28543
rect 3341 28441 3375 28475
rect 3525 28441 3559 28475
rect 8953 28441 8987 28475
rect 10977 28441 11011 28475
rect 12624 28441 12658 28475
rect 15200 28441 15234 28475
rect 7573 28373 7607 28407
rect 9153 28373 9187 28407
rect 10517 28373 10551 28407
rect 12265 28373 12299 28407
rect 14749 28373 14783 28407
rect 7757 28169 7791 28203
rect 8769 28169 8803 28203
rect 10609 28169 10643 28203
rect 10977 28169 11011 28203
rect 11529 28169 11563 28203
rect 13001 28169 13035 28203
rect 13369 28169 13403 28203
rect 15301 28169 15335 28203
rect 6837 28101 6871 28135
rect 8125 28101 8159 28135
rect 3045 28033 3079 28067
rect 4261 28033 4295 28067
rect 4445 28033 4479 28067
rect 6745 28033 6779 28067
rect 6929 28033 6963 28067
rect 7297 28033 7331 28067
rect 7573 28033 7607 28067
rect 7941 28033 7975 28067
rect 8401 28033 8435 28067
rect 9137 28033 9171 28067
rect 12642 28033 12676 28067
rect 12909 28033 12943 28067
rect 14381 28033 14415 28067
rect 15577 28033 15611 28067
rect 15669 28033 15703 28067
rect 15761 28033 15795 28067
rect 15945 28033 15979 28067
rect 16037 28033 16071 28067
rect 2789 27965 2823 27999
rect 7205 27965 7239 27999
rect 7665 27965 7699 27999
rect 9229 27965 9263 27999
rect 9413 27965 9447 27999
rect 11069 27965 11103 27999
rect 11161 27965 11195 27999
rect 13461 27965 13495 27999
rect 13553 27965 13587 27999
rect 15117 27965 15151 27999
rect 4261 27897 4295 27931
rect 8217 27897 8251 27931
rect 4169 27829 4203 27863
rect 7021 27829 7055 27863
rect 13829 27829 13863 27863
rect 14565 27829 14599 27863
rect 16221 27829 16255 27863
rect 10977 27625 11011 27659
rect 8953 27557 8987 27591
rect 12357 27557 12391 27591
rect 4077 27489 4111 27523
rect 11621 27489 11655 27523
rect 12817 27489 12851 27523
rect 12909 27489 12943 27523
rect 13737 27489 13771 27523
rect 2053 27421 2087 27455
rect 3801 27421 3835 27455
rect 3985 27421 4019 27455
rect 5549 27421 5583 27455
rect 7573 27421 7607 27455
rect 8769 27421 8803 27455
rect 8953 27421 8987 27455
rect 9137 27421 9171 27455
rect 9597 27421 9631 27455
rect 9864 27421 9898 27455
rect 11437 27421 11471 27455
rect 11805 27421 11839 27455
rect 13553 27421 13587 27455
rect 14105 27421 14139 27455
rect 15853 27421 15887 27455
rect 15945 27421 15979 27455
rect 16037 27421 16071 27455
rect 16221 27421 16255 27455
rect 2320 27353 2354 27387
rect 4344 27353 4378 27387
rect 5816 27353 5850 27387
rect 12725 27353 12759 27387
rect 14372 27353 14406 27387
rect 3433 27285 3467 27319
rect 3893 27285 3927 27319
rect 5457 27285 5491 27319
rect 6929 27285 6963 27319
rect 7021 27285 7055 27319
rect 8125 27285 8159 27319
rect 11253 27285 11287 27319
rect 11897 27285 11931 27319
rect 12265 27285 12299 27319
rect 13185 27285 13219 27319
rect 13645 27285 13679 27319
rect 15485 27285 15519 27319
rect 15577 27285 15611 27319
rect 2145 27081 2179 27115
rect 2881 27081 2915 27115
rect 4629 27081 4663 27115
rect 7757 27081 7791 27115
rect 9413 27081 9447 27115
rect 12541 27081 12575 27115
rect 12909 27081 12943 27115
rect 1593 27013 1627 27047
rect 2789 27013 2823 27047
rect 2998 27013 3032 27047
rect 11621 27013 11655 27047
rect 12449 27013 12483 27047
rect 15200 27013 15234 27047
rect 1501 26945 1535 26979
rect 1685 26945 1719 26979
rect 1777 26945 1811 26979
rect 3238 26945 3272 26979
rect 3516 26945 3550 26979
rect 4988 26945 5022 26979
rect 6377 26945 6411 26979
rect 6644 26945 6678 26979
rect 8033 26945 8067 26979
rect 8289 26945 8323 26979
rect 9965 26945 9999 26979
rect 10057 26945 10091 26979
rect 10425 26945 10459 26979
rect 13001 26945 13035 26979
rect 14585 26945 14619 26979
rect 14841 26945 14875 26979
rect 14933 26945 14967 26979
rect 2053 26877 2087 26911
rect 2262 26877 2296 26911
rect 2513 26877 2547 26911
rect 4721 26877 4755 26911
rect 10241 26877 10275 26911
rect 10977 26877 11011 26911
rect 13093 26877 13127 26911
rect 2421 26809 2455 26843
rect 3157 26809 3191 26843
rect 6101 26741 6135 26775
rect 9597 26741 9631 26775
rect 13461 26741 13495 26775
rect 16313 26741 16347 26775
rect 1961 26537 1995 26571
rect 2605 26537 2639 26571
rect 6377 26537 6411 26571
rect 8033 26537 8067 26571
rect 10333 26537 10367 26571
rect 14105 26537 14139 26571
rect 15577 26537 15611 26571
rect 3617 26469 3651 26503
rect 4629 26469 4663 26503
rect 5825 26469 5859 26503
rect 11897 26469 11931 26503
rect 2421 26401 2455 26435
rect 2764 26401 2798 26435
rect 2973 26401 3007 26435
rect 4721 26401 4755 26435
rect 4997 26401 5031 26435
rect 5089 26401 5123 26435
rect 5206 26401 5240 26435
rect 8493 26401 8527 26435
rect 8677 26401 8711 26435
rect 13921 26401 13955 26435
rect 2329 26333 2363 26367
rect 3249 26333 3283 26367
rect 3341 26333 3375 26367
rect 3617 26333 3651 26367
rect 3985 26333 4019 26367
rect 5457 26333 5491 26367
rect 5733 26333 5767 26367
rect 6101 26333 6135 26367
rect 6285 26333 6319 26367
rect 6469 26333 6503 26367
rect 6561 26333 6595 26367
rect 8953 26333 8987 26367
rect 9220 26333 9254 26367
rect 10425 26333 10459 26367
rect 13021 26333 13055 26367
rect 13277 26333 13311 26367
rect 14657 26333 14691 26367
rect 15393 26333 15427 26367
rect 15853 26333 15887 26367
rect 15945 26333 15979 26367
rect 16037 26333 16071 26367
rect 16221 26333 16255 26367
rect 4353 26265 4387 26299
rect 4470 26265 4504 26299
rect 5549 26265 5583 26299
rect 5825 26265 5859 26299
rect 6828 26265 6862 26299
rect 8401 26265 8435 26299
rect 10692 26265 10726 26299
rect 13553 26265 13587 26299
rect 13737 26265 13771 26299
rect 2881 26197 2915 26231
rect 3433 26197 3467 26231
rect 4261 26197 4295 26231
rect 5365 26197 5399 26231
rect 5634 26197 5668 26231
rect 6009 26197 6043 26231
rect 7941 26197 7975 26231
rect 11805 26197 11839 26231
rect 14841 26197 14875 26231
rect 3985 25993 4019 26027
rect 5386 25993 5420 26027
rect 5733 25993 5767 26027
rect 7113 25993 7147 26027
rect 9597 25993 9631 26027
rect 9689 25993 9723 26027
rect 10609 25993 10643 26027
rect 10977 25993 11011 26027
rect 14289 25993 14323 26027
rect 14657 25993 14691 26027
rect 15117 25993 15151 26027
rect 3309 25925 3343 25959
rect 3525 25925 3559 25959
rect 4169 25925 4203 25959
rect 5181 25925 5215 25959
rect 7205 25925 7239 25959
rect 10057 25925 10091 25959
rect 12940 25925 12974 25959
rect 14105 25925 14139 25959
rect 16129 25925 16163 25959
rect 3801 25857 3835 25891
rect 3893 25857 3927 25891
rect 4629 25857 4663 25891
rect 5641 25857 5675 25891
rect 5825 25857 5859 25891
rect 6193 25857 6227 25891
rect 7941 25857 7975 25891
rect 8484 25857 8518 25891
rect 10149 25857 10183 25891
rect 11069 25857 11103 25891
rect 13185 25857 13219 25891
rect 13277 25857 13311 25891
rect 15301 25857 15335 25891
rect 15393 25857 15427 25891
rect 15577 25857 15611 25891
rect 15669 25857 15703 25891
rect 15945 25857 15979 25891
rect 4261 25789 4295 25823
rect 4721 25789 4755 25823
rect 6561 25789 6595 25823
rect 8217 25789 8251 25823
rect 10241 25789 10275 25823
rect 11161 25789 11195 25823
rect 14749 25789 14783 25823
rect 14841 25789 14875 25823
rect 3157 25721 3191 25755
rect 3617 25721 3651 25755
rect 6101 25721 6135 25755
rect 15761 25721 15795 25755
rect 3341 25653 3375 25687
rect 5365 25653 5399 25687
rect 5549 25653 5583 25687
rect 11805 25653 11839 25687
rect 6653 25449 6687 25483
rect 7021 25449 7055 25483
rect 7665 25449 7699 25483
rect 7849 25449 7883 25483
rect 8125 25449 8159 25483
rect 9045 25449 9079 25483
rect 11069 25449 11103 25483
rect 6745 25313 6779 25347
rect 7941 25313 7975 25347
rect 8769 25313 8803 25347
rect 9597 25313 9631 25347
rect 11345 25313 11379 25347
rect 13185 25313 13219 25347
rect 14933 25313 14967 25347
rect 1409 25245 1443 25279
rect 6837 25245 6871 25279
rect 7113 25245 7147 25279
rect 7481 25245 7515 25279
rect 8033 25245 8067 25279
rect 10425 25245 10459 25279
rect 11253 25245 11287 25279
rect 12357 25245 12391 25279
rect 13001 25245 13035 25279
rect 14289 25245 14323 25279
rect 14381 25245 14415 25279
rect 14565 25245 14599 25279
rect 14657 25245 14691 25279
rect 5641 25177 5675 25211
rect 6469 25177 6503 25211
rect 9413 25177 9447 25211
rect 15200 25177 15234 25211
rect 1593 25109 1627 25143
rect 9505 25109 9539 25143
rect 9873 25109 9907 25143
rect 11989 25109 12023 25143
rect 12173 25109 12207 25143
rect 12449 25109 12483 25143
rect 13829 25109 13863 25143
rect 14105 25109 14139 25143
rect 16313 25109 16347 25143
rect 2053 24905 2087 24939
rect 8769 24905 8803 24939
rect 9321 24905 9355 24939
rect 11345 24905 11379 24939
rect 12909 24905 12943 24939
rect 13369 24905 13403 24939
rect 8677 24837 8711 24871
rect 1961 24769 1995 24803
rect 3525 24769 3559 24803
rect 3985 24769 4019 24803
rect 4169 24769 4203 24803
rect 4629 24769 4663 24803
rect 5273 24769 5307 24803
rect 5457 24769 5491 24803
rect 5641 24769 5675 24803
rect 6377 24769 6411 24803
rect 6561 24769 6595 24803
rect 6837 24769 6871 24803
rect 7104 24769 7138 24803
rect 9229 24769 9263 24803
rect 9965 24769 9999 24803
rect 10232 24769 10266 24803
rect 11785 24769 11819 24803
rect 13461 24769 13495 24803
rect 14105 24769 14139 24803
rect 14197 24769 14231 24803
rect 14381 24769 14415 24803
rect 14473 24769 14507 24803
rect 14565 24769 14599 24803
rect 14933 24769 14967 24803
rect 15200 24769 15234 24803
rect 1844 24701 1878 24735
rect 2329 24701 2363 24735
rect 3893 24701 3927 24735
rect 4813 24701 4847 24735
rect 6469 24701 6503 24735
rect 8953 24701 8987 24735
rect 11529 24701 11563 24735
rect 13553 24701 13587 24735
rect 4353 24633 4387 24667
rect 13921 24633 13955 24667
rect 1685 24565 1719 24599
rect 3709 24565 3743 24599
rect 4445 24565 4479 24599
rect 5457 24565 5491 24599
rect 8217 24565 8251 24599
rect 8309 24565 8343 24599
rect 13001 24565 13035 24599
rect 14841 24565 14875 24599
rect 16313 24565 16347 24599
rect 2973 24361 3007 24395
rect 6653 24361 6687 24395
rect 7205 24361 7239 24395
rect 7389 24361 7423 24395
rect 10149 24361 10183 24395
rect 15485 24361 15519 24395
rect 15577 24361 15611 24395
rect 3893 24293 3927 24327
rect 11989 24293 12023 24327
rect 4629 24225 4663 24259
rect 4997 24225 5031 24259
rect 5114 24225 5148 24259
rect 5641 24225 5675 24259
rect 7021 24225 7055 24259
rect 10609 24225 10643 24259
rect 10701 24225 10735 24259
rect 13369 24225 13403 24259
rect 1501 24157 1535 24191
rect 1768 24157 1802 24191
rect 2973 24157 3007 24191
rect 3157 24157 3191 24191
rect 3463 24157 3497 24191
rect 3617 24157 3651 24191
rect 3801 24157 3835 24191
rect 3985 24157 4019 24191
rect 4169 24157 4203 24191
rect 5365 24157 5399 24191
rect 6377 24157 6411 24191
rect 6469 24157 6503 24191
rect 6929 24157 6963 24191
rect 8502 24157 8536 24191
rect 8769 24157 8803 24191
rect 9781 24157 9815 24191
rect 9873 24157 9907 24191
rect 10057 24157 10091 24191
rect 11253 24157 11287 24191
rect 11345 24157 11379 24191
rect 11529 24157 11563 24191
rect 11621 24157 11655 24191
rect 11805 24157 11839 24191
rect 13553 24157 13587 24191
rect 13737 24157 13771 24191
rect 14381 24157 14415 24191
rect 14473 24157 14507 24191
rect 14565 24154 14599 24188
rect 14749 24157 14783 24191
rect 14841 24157 14875 24191
rect 15025 24157 15059 24191
rect 15117 24157 15151 24191
rect 15209 24157 15243 24191
rect 15761 24157 15795 24191
rect 16129 24157 16163 24191
rect 3249 24089 3283 24123
rect 4905 24089 4939 24123
rect 5850 24089 5884 24123
rect 6101 24089 6135 24123
rect 9965 24089 9999 24123
rect 13102 24089 13136 24123
rect 13921 24089 13955 24123
rect 15853 24089 15887 24123
rect 15945 24089 15979 24123
rect 2881 24021 2915 24055
rect 4261 24021 4295 24055
rect 5273 24021 5307 24055
rect 5733 24021 5767 24055
rect 6009 24021 6043 24055
rect 6285 24021 6319 24055
rect 9689 24021 9723 24055
rect 10517 24021 10551 24055
rect 11069 24021 11103 24055
rect 11437 24021 11471 24055
rect 11713 24021 11747 24055
rect 14105 24021 14139 24055
rect 2973 23817 3007 23851
rect 10609 23817 10643 23851
rect 13093 23817 13127 23851
rect 14565 23817 14599 23851
rect 15025 23817 15059 23851
rect 11805 23749 11839 23783
rect 13452 23749 13486 23783
rect 14841 23749 14875 23783
rect 15945 23749 15979 23783
rect 16129 23749 16163 23783
rect 1409 23681 1443 23715
rect 1676 23681 1710 23715
rect 2881 23681 2915 23715
rect 3065 23681 3099 23715
rect 3157 23681 3191 23715
rect 3341 23681 3375 23715
rect 3433 23681 3467 23715
rect 3525 23681 3559 23715
rect 4169 23681 4203 23715
rect 4261 23681 4295 23715
rect 4537 23681 4571 23715
rect 4813 23681 4847 23715
rect 5080 23681 5114 23715
rect 9496 23681 9530 23715
rect 10701 23681 10735 23715
rect 11713 23681 11747 23715
rect 11897 23681 11931 23715
rect 12081 23681 12115 23715
rect 12449 23681 12483 23715
rect 12541 23681 12575 23715
rect 12725 23681 12759 23715
rect 12817 23681 12851 23715
rect 12909 23681 12943 23715
rect 14657 23681 14691 23715
rect 15117 23681 15151 23715
rect 15301 23681 15335 23715
rect 15393 23681 15427 23715
rect 15485 23681 15519 23715
rect 9229 23613 9263 23647
rect 11345 23613 11379 23647
rect 13185 23613 13219 23647
rect 4445 23545 4479 23579
rect 11529 23545 11563 23579
rect 15761 23545 15795 23579
rect 2789 23477 2823 23511
rect 3801 23477 3835 23511
rect 3985 23477 4019 23511
rect 6193 23477 6227 23511
rect 12265 23477 12299 23511
rect 15669 23477 15703 23511
rect 1593 23273 1627 23307
rect 2605 23273 2639 23307
rect 3249 23273 3283 23307
rect 8033 23273 8067 23307
rect 9137 23273 9171 23307
rect 10701 23273 10735 23307
rect 11161 23273 11195 23307
rect 11437 23273 11471 23307
rect 11529 23273 11563 23307
rect 11805 23273 11839 23307
rect 3157 23205 3191 23239
rect 1961 23137 1995 23171
rect 2237 23137 2271 23171
rect 3341 23137 3375 23171
rect 7941 23137 7975 23171
rect 9689 23137 9723 23171
rect 11621 23145 11655 23179
rect 11713 23137 11747 23171
rect 11897 23137 11931 23171
rect 12725 23137 12759 23171
rect 1869 23069 1903 23103
rect 2329 23069 2363 23103
rect 2513 23069 2547 23103
rect 2973 23069 3007 23103
rect 3249 23069 3283 23103
rect 3801 23069 3835 23103
rect 3985 23069 4019 23103
rect 4077 23069 4111 23103
rect 4169 23069 4203 23103
rect 4721 23069 4755 23103
rect 6202 23069 6236 23103
rect 6469 23069 6503 23103
rect 8033 23069 8067 23103
rect 8217 23069 8251 23103
rect 9597 23069 9631 23103
rect 9965 23069 9999 23103
rect 10885 23069 10919 23103
rect 10977 23069 11011 23103
rect 11253 23069 11287 23103
rect 11345 23069 11379 23103
rect 11989 23069 12023 23103
rect 12265 23069 12299 23103
rect 12357 23069 12391 23103
rect 12633 23069 12667 23103
rect 14105 23069 14139 23103
rect 14289 23069 14323 23103
rect 14381 23069 14415 23103
rect 14473 23069 14507 23103
rect 14841 23069 14875 23103
rect 1752 23001 1786 23035
rect 2421 23001 2455 23035
rect 4537 23001 4571 23035
rect 7696 23001 7730 23035
rect 12449 23001 12483 23035
rect 13461 23001 13495 23035
rect 14749 23001 14783 23035
rect 15086 23001 15120 23035
rect 2789 22933 2823 22967
rect 2881 22933 2915 22967
rect 3617 22933 3651 22967
rect 4445 22933 4479 22967
rect 4905 22933 4939 22967
rect 5089 22933 5123 22967
rect 6561 22933 6595 22967
rect 9505 22933 9539 22967
rect 10609 22933 10643 22967
rect 12081 22933 12115 22967
rect 13369 22933 13403 22967
rect 16221 22933 16255 22967
rect 2529 22729 2563 22763
rect 2697 22729 2731 22763
rect 9781 22729 9815 22763
rect 11161 22729 11195 22763
rect 15301 22729 15335 22763
rect 16221 22729 16255 22763
rect 2329 22661 2363 22695
rect 6377 22661 6411 22695
rect 6561 22661 6595 22695
rect 8668 22661 8702 22695
rect 13737 22661 13771 22695
rect 15577 22661 15611 22695
rect 15761 22661 15795 22695
rect 15853 22661 15887 22695
rect 1961 22593 1995 22627
rect 2053 22593 2087 22627
rect 2237 22593 2271 22627
rect 3065 22593 3099 22627
rect 3893 22593 3927 22627
rect 4261 22593 4295 22627
rect 4537 22593 4571 22627
rect 4721 22593 4755 22627
rect 5181 22593 5215 22627
rect 5825 22593 5859 22627
rect 5917 22593 5951 22627
rect 6929 22593 6963 22627
rect 7196 22593 7230 22627
rect 10425 22593 10459 22627
rect 10609 22593 10643 22627
rect 10793 22593 10827 22627
rect 10885 22593 10919 22627
rect 10977 22593 11011 22627
rect 11529 22593 11563 22627
rect 13286 22593 13320 22627
rect 13553 22593 13587 22627
rect 13645 22593 13679 22627
rect 13829 22593 13863 22627
rect 14188 22593 14222 22627
rect 16037 22593 16071 22627
rect 3157 22525 3191 22559
rect 5273 22525 5307 22559
rect 5549 22525 5583 22559
rect 6009 22525 6043 22559
rect 6101 22525 6135 22559
rect 8401 22525 8435 22559
rect 13921 22525 13955 22559
rect 2237 22457 2271 22491
rect 3433 22457 3467 22491
rect 4445 22457 4479 22491
rect 12173 22457 12207 22491
rect 15393 22457 15427 22491
rect 2513 22389 2547 22423
rect 4077 22389 4111 22423
rect 4629 22389 4663 22423
rect 4905 22389 4939 22423
rect 5641 22389 5675 22423
rect 8309 22389 8343 22423
rect 9873 22389 9907 22423
rect 8309 22185 8343 22219
rect 8953 22185 8987 22219
rect 10333 22185 10367 22219
rect 11989 22185 12023 22219
rect 13553 22185 13587 22219
rect 3617 22117 3651 22151
rect 3341 22049 3375 22083
rect 6929 22049 6963 22083
rect 9505 22049 9539 22083
rect 10517 22049 10551 22083
rect 12357 22049 12391 22083
rect 12449 22049 12483 22083
rect 12909 22049 12943 22083
rect 13093 22049 13127 22083
rect 3249 21981 3283 22015
rect 3985 21981 4019 22015
rect 4133 21981 4167 22015
rect 4491 21981 4525 22015
rect 5457 21981 5491 22015
rect 6377 21981 6411 22015
rect 6653 21981 6687 22015
rect 6837 21981 6871 22015
rect 9781 21981 9815 22015
rect 9873 21981 9907 22015
rect 10057 21981 10091 22015
rect 10149 21981 10183 22015
rect 10701 21981 10735 22015
rect 12173 21981 12207 22015
rect 12265 21981 12299 22015
rect 13185 21981 13219 22015
rect 13921 21981 13955 22015
rect 15393 21981 15427 22015
rect 15669 21981 15703 22015
rect 16037 21981 16071 22015
rect 4261 21913 4295 21947
rect 4353 21913 4387 21947
rect 5641 21913 5675 21947
rect 7196 21913 7230 21947
rect 10977 21913 11011 21947
rect 11805 21913 11839 21947
rect 14105 21913 14139 21947
rect 14841 21913 14875 21947
rect 4629 21845 4663 21879
rect 6745 21845 6779 21879
rect 9321 21845 9355 21879
rect 9413 21845 9447 21879
rect 10885 21845 10919 21879
rect 13737 21845 13771 21879
rect 15209 21845 15243 21879
rect 15853 21845 15887 21879
rect 16221 21845 16255 21879
rect 3893 21641 3927 21675
rect 5273 21641 5307 21675
rect 5365 21641 5399 21675
rect 7573 21641 7607 21675
rect 10885 21641 10919 21675
rect 14565 21641 14599 21675
rect 15485 21641 15519 21675
rect 3525 21573 3559 21607
rect 4721 21573 4755 21607
rect 5482 21573 5516 21607
rect 6101 21573 6135 21607
rect 8217 21573 8251 21607
rect 1409 21505 1443 21539
rect 2881 21505 2915 21539
rect 3065 21505 3099 21539
rect 3249 21505 3283 21539
rect 3433 21505 3467 21539
rect 3617 21505 3651 21539
rect 4077 21505 4111 21539
rect 4169 21505 4203 21539
rect 4353 21505 4387 21539
rect 4445 21505 4479 21539
rect 4905 21505 4939 21539
rect 5917 21505 5951 21539
rect 6190 21495 6224 21529
rect 6561 21505 6595 21539
rect 6929 21505 6963 21539
rect 7665 21505 7699 21539
rect 7849 21505 7883 21539
rect 9505 21505 9539 21539
rect 9772 21505 9806 21539
rect 10977 21505 11011 21539
rect 11529 21505 11563 21539
rect 11713 21505 11747 21539
rect 12081 21505 12115 21539
rect 12624 21505 12658 21539
rect 14841 21505 14875 21539
rect 14933 21505 14967 21539
rect 15025 21505 15059 21539
rect 15209 21505 15243 21539
rect 15301 21505 15335 21539
rect 15761 21505 15795 21539
rect 15945 21505 15979 21539
rect 16037 21505 16071 21539
rect 2973 21437 3007 21471
rect 4997 21437 5031 21471
rect 8953 21437 8987 21471
rect 11069 21437 11103 21471
rect 11805 21437 11839 21471
rect 11897 21437 11931 21471
rect 12357 21437 12391 21471
rect 14381 21437 14415 21471
rect 6377 21369 6411 21403
rect 13737 21369 13771 21403
rect 15577 21369 15611 21403
rect 1593 21301 1627 21335
rect 3801 21301 3835 21335
rect 4537 21301 4571 21335
rect 5641 21301 5675 21335
rect 5733 21301 5767 21335
rect 7665 21301 7699 21335
rect 10977 21301 11011 21335
rect 11345 21301 11379 21335
rect 12265 21301 12299 21335
rect 13829 21301 13863 21335
rect 16221 21301 16255 21335
rect 3341 21097 3375 21131
rect 3801 21097 3835 21131
rect 6193 21097 6227 21131
rect 8309 21097 8343 21131
rect 9781 21097 9815 21131
rect 10793 21097 10827 21131
rect 12357 21097 12391 21131
rect 12725 21097 12759 21131
rect 2237 21029 2271 21063
rect 10149 21029 10183 21063
rect 12541 21029 12575 21063
rect 1685 20961 1719 20995
rect 2697 20961 2731 20995
rect 2789 20961 2823 20995
rect 3065 20961 3099 20995
rect 4445 20961 4479 20995
rect 5549 20961 5583 20995
rect 6745 20961 6779 20995
rect 6929 20961 6963 20995
rect 10057 20961 10091 20995
rect 10977 20961 11011 20995
rect 13185 20961 13219 20995
rect 13277 20961 13311 20995
rect 1777 20893 1811 20927
rect 2580 20893 2614 20927
rect 3157 20893 3191 20927
rect 3311 20893 3345 20927
rect 3982 20893 4016 20927
rect 4353 20893 4387 20927
rect 4537 20893 4571 20927
rect 4813 20893 4847 20927
rect 5825 20893 5859 20927
rect 6653 20893 6687 20927
rect 8953 20893 8987 20927
rect 9965 20893 9999 20927
rect 10241 20893 10275 20927
rect 10425 20893 10459 20927
rect 10609 20893 10643 20927
rect 10701 20893 10735 20927
rect 10885 20893 10919 20927
rect 11713 20893 11747 20927
rect 11897 20893 11931 20927
rect 11989 20893 12023 20927
rect 12081 20893 12115 20927
rect 12449 20893 12483 20927
rect 12633 20893 12667 20927
rect 13093 20893 13127 20927
rect 14933 20893 14967 20927
rect 2237 20825 2271 20859
rect 5917 20825 5951 20859
rect 6034 20825 6068 20859
rect 7196 20825 7230 20859
rect 10517 20825 10551 20859
rect 14381 20825 14415 20859
rect 14565 20825 14599 20859
rect 15178 20825 15212 20859
rect 1501 20757 1535 20791
rect 2421 20757 2455 20791
rect 3985 20757 4019 20791
rect 6285 20757 6319 20791
rect 11621 20757 11655 20791
rect 14197 20757 14231 20791
rect 16313 20757 16347 20791
rect 2881 20553 2915 20587
rect 4445 20553 4479 20587
rect 6377 20553 6411 20587
rect 8861 20553 8895 20587
rect 10609 20553 10643 20587
rect 11621 20553 11655 20587
rect 14841 20553 14875 20587
rect 14933 20553 14967 20587
rect 15669 20553 15703 20587
rect 1768 20485 1802 20519
rect 7490 20485 7524 20519
rect 13369 20485 13403 20519
rect 13706 20485 13740 20519
rect 3341 20417 3375 20451
rect 3801 20417 3835 20451
rect 4169 20417 4203 20451
rect 4261 20417 4295 20451
rect 4997 20417 5031 20451
rect 5641 20417 5675 20451
rect 8677 20417 8711 20451
rect 11069 20417 11103 20451
rect 11529 20417 11563 20451
rect 12725 20417 12759 20451
rect 12909 20417 12943 20451
rect 13001 20417 13035 20451
rect 13093 20417 13127 20451
rect 15209 20417 15243 20451
rect 15301 20417 15335 20451
rect 15393 20417 15427 20451
rect 15577 20417 15611 20451
rect 15853 20417 15887 20451
rect 15945 20417 15979 20451
rect 16129 20417 16163 20451
rect 16221 20417 16255 20451
rect 1501 20349 1535 20383
rect 2973 20349 3007 20383
rect 3249 20349 3283 20383
rect 5273 20349 5307 20383
rect 5549 20349 5583 20383
rect 7757 20349 7791 20383
rect 9413 20349 9447 20383
rect 10793 20349 10827 20383
rect 10885 20349 10919 20383
rect 10977 20349 11011 20383
rect 13461 20349 13495 20383
rect 5457 20281 5491 20315
rect 3893 20213 3927 20247
rect 8125 20213 8159 20247
rect 3617 20009 3651 20043
rect 4169 20009 4203 20043
rect 4353 20009 4387 20043
rect 6745 20009 6779 20043
rect 8493 20009 8527 20043
rect 15485 20009 15519 20043
rect 16221 20009 16255 20043
rect 2789 19941 2823 19975
rect 9045 19941 9079 19975
rect 11713 19941 11747 19975
rect 1409 19873 1443 19907
rect 3157 19873 3191 19907
rect 4997 19873 5031 19907
rect 8217 19873 8251 19907
rect 8493 19873 8527 19907
rect 8585 19873 8619 19907
rect 9229 19873 9263 19907
rect 11161 19873 11195 19907
rect 11529 19873 11563 19907
rect 1665 19805 1699 19839
rect 3249 19805 3283 19839
rect 3433 19805 3467 19839
rect 4353 19805 4387 19839
rect 4445 19805 4479 19839
rect 4905 19805 4939 19839
rect 5365 19805 5399 19839
rect 5632 19805 5666 19839
rect 7573 19805 7607 19839
rect 7757 19805 7791 19839
rect 7849 19805 7883 19839
rect 7941 19805 7975 19839
rect 8677 19805 8711 19839
rect 8953 19805 8987 19839
rect 9689 19805 9723 19839
rect 9781 19805 9815 19839
rect 9965 19805 9999 19839
rect 10057 19805 10091 19839
rect 11069 19805 11103 19839
rect 11437 19805 11471 19839
rect 11805 19805 11839 19839
rect 12265 19805 12299 19839
rect 13921 19805 13955 19839
rect 14105 19805 14139 19839
rect 15669 19805 15703 19839
rect 15945 19805 15979 19839
rect 16037 19805 16071 19839
rect 4629 19737 4663 19771
rect 8309 19737 8343 19771
rect 9229 19737 9263 19771
rect 14372 19737 14406 19771
rect 15853 19737 15887 19771
rect 5273 19669 5307 19703
rect 9505 19669 9539 19703
rect 11897 19669 11931 19703
rect 11989 19669 12023 19703
rect 13737 19669 13771 19703
rect 4077 19465 4111 19499
rect 5365 19465 5399 19499
rect 5457 19465 5491 19499
rect 8309 19465 8343 19499
rect 10701 19465 10735 19499
rect 10885 19465 10919 19499
rect 11253 19465 11287 19499
rect 11621 19465 11655 19499
rect 12449 19465 12483 19499
rect 13001 19465 13035 19499
rect 14105 19465 14139 19499
rect 2513 19397 2547 19431
rect 3617 19397 3651 19431
rect 5917 19397 5951 19431
rect 8769 19397 8803 19431
rect 9312 19397 9346 19431
rect 12081 19397 12115 19431
rect 1961 19329 1995 19363
rect 2881 19329 2915 19363
rect 3340 19329 3374 19363
rect 3433 19329 3467 19363
rect 4169 19329 4203 19363
rect 4261 19329 4295 19363
rect 4905 19329 4939 19363
rect 5181 19329 5215 19363
rect 5641 19329 5675 19363
rect 5733 19329 5767 19363
rect 7196 19329 7230 19363
rect 8401 19329 8435 19363
rect 10609 19329 10643 19363
rect 10793 19329 10827 19363
rect 11069 19329 11103 19363
rect 11345 19329 11379 19363
rect 11529 19329 11563 19363
rect 11713 19329 11747 19363
rect 11897 19329 11931 19363
rect 12173 19329 12207 19363
rect 12265 19329 12299 19363
rect 12909 19329 12943 19363
rect 13369 19329 13403 19363
rect 14381 19329 14415 19363
rect 14473 19329 14507 19363
rect 14565 19329 14599 19363
rect 14749 19329 14783 19363
rect 15189 19329 15223 19363
rect 2053 19261 2087 19295
rect 5089 19261 5123 19295
rect 6929 19261 6963 19295
rect 9045 19261 9079 19295
rect 13093 19261 13127 19295
rect 13921 19261 13955 19295
rect 14933 19261 14967 19295
rect 3985 19193 4019 19227
rect 4997 19193 5031 19227
rect 2329 19125 2363 19159
rect 3249 19125 3283 19159
rect 5917 19125 5951 19159
rect 8769 19125 8803 19159
rect 8953 19125 8987 19159
rect 10425 19125 10459 19159
rect 12541 19125 12575 19159
rect 16313 19125 16347 19159
rect 8953 18921 8987 18955
rect 10149 18921 10183 18955
rect 10701 18921 10735 18955
rect 11897 18921 11931 18955
rect 14289 18921 14323 18955
rect 14933 18921 14967 18955
rect 8677 18853 8711 18887
rect 9965 18853 9999 18887
rect 10517 18853 10551 18887
rect 13645 18853 13679 18887
rect 9321 18785 9355 18819
rect 9689 18785 9723 18819
rect 11345 18785 11379 18819
rect 5917 18717 5951 18751
rect 6101 18717 6135 18751
rect 6285 18717 6319 18751
rect 8309 18717 8343 18751
rect 8493 18717 8527 18751
rect 8769 18717 8803 18751
rect 9597 18717 9631 18751
rect 10977 18717 11011 18751
rect 11161 18717 11195 18751
rect 11253 18717 11287 18751
rect 11529 18717 11563 18751
rect 11805 18717 11839 18751
rect 11989 18717 12023 18751
rect 12265 18717 12299 18751
rect 12532 18717 12566 18751
rect 13921 18717 13955 18751
rect 14473 18717 14507 18751
rect 14565 18717 14599 18751
rect 14749 18717 14783 18751
rect 14841 18717 14875 18751
rect 15209 18717 15243 18751
rect 15301 18717 15335 18751
rect 15393 18717 15427 18751
rect 15577 18717 15611 18751
rect 15853 18717 15887 18751
rect 16221 18717 16255 18751
rect 6837 18649 6871 18683
rect 8064 18649 8098 18683
rect 9112 18649 9146 18683
rect 10241 18649 10275 18683
rect 15945 18649 15979 18683
rect 16037 18649 16071 18683
rect 6009 18581 6043 18615
rect 6929 18581 6963 18615
rect 9229 18581 9263 18615
rect 11713 18581 11747 18615
rect 13737 18581 13771 18615
rect 15669 18581 15703 18615
rect 6561 18377 6595 18411
rect 8493 18377 8527 18411
rect 10149 18377 10183 18411
rect 10977 18377 11011 18411
rect 11345 18377 11379 18411
rect 14197 18377 14231 18411
rect 16313 18377 16347 18411
rect 3893 18309 3927 18343
rect 7380 18309 7414 18343
rect 8585 18309 8619 18343
rect 9781 18309 9815 18343
rect 9997 18309 10031 18343
rect 16129 18309 16163 18343
rect 2329 18241 2363 18275
rect 2513 18241 2547 18275
rect 4813 18241 4847 18275
rect 5549 18241 5583 18275
rect 6377 18241 6411 18275
rect 6561 18241 6595 18275
rect 6837 18241 6871 18275
rect 7113 18241 7147 18275
rect 9413 18241 9447 18275
rect 9505 18241 9539 18275
rect 10241 18241 10275 18275
rect 10425 18241 10459 18275
rect 10609 18241 10643 18275
rect 10885 18241 10919 18275
rect 11161 18241 11195 18275
rect 11897 18241 11931 18275
rect 12164 18241 12198 18275
rect 14381 18241 14415 18275
rect 14729 18241 14763 18275
rect 15945 18241 15979 18275
rect 13921 18173 13955 18207
rect 14473 18173 14507 18207
rect 8861 18105 8895 18139
rect 9045 18105 9079 18139
rect 13277 18105 13311 18139
rect 2329 18037 2363 18071
rect 6745 18037 6779 18071
rect 9413 18037 9447 18071
rect 9965 18037 9999 18071
rect 13369 18037 13403 18071
rect 15853 18037 15887 18071
rect 1593 17833 1627 17867
rect 2053 17833 2087 17867
rect 3525 17833 3559 17867
rect 4537 17833 4571 17867
rect 5365 17833 5399 17867
rect 7297 17833 7331 17867
rect 7573 17833 7607 17867
rect 10241 17833 10275 17867
rect 12265 17833 12299 17867
rect 14381 17833 14415 17867
rect 2789 17765 2823 17799
rect 8585 17765 8619 17799
rect 12817 17697 12851 17731
rect 15117 17697 15151 17731
rect 2421 17629 2455 17663
rect 2605 17629 2639 17663
rect 2697 17629 2731 17663
rect 3160 17629 3194 17663
rect 3433 17629 3467 17663
rect 3617 17629 3651 17663
rect 3801 17629 3835 17663
rect 3893 17629 3927 17663
rect 4721 17629 4755 17663
rect 5181 17629 5215 17663
rect 5274 17629 5308 17663
rect 7297 17629 7331 17663
rect 7481 17629 7515 17663
rect 7757 17629 7791 17663
rect 7849 17629 7883 17663
rect 7941 17629 7975 17663
rect 8125 17629 8159 17663
rect 8401 17629 8435 17663
rect 8677 17629 8711 17663
rect 8953 17629 8987 17663
rect 12633 17629 12667 17663
rect 13553 17629 13587 17663
rect 13645 17629 13679 17663
rect 13737 17629 13771 17663
rect 13921 17629 13955 17663
rect 14105 17629 14139 17663
rect 14657 17629 14691 17663
rect 14749 17629 14783 17663
rect 14841 17629 14875 17663
rect 15025 17629 15059 17663
rect 15485 17629 15519 17663
rect 16313 17629 16347 17663
rect 1777 17561 1811 17595
rect 2237 17561 2271 17595
rect 4905 17561 4939 17595
rect 15301 17561 15335 17595
rect 15577 17561 15611 17595
rect 15761 17561 15795 17595
rect 1409 17493 1443 17527
rect 1577 17493 1611 17527
rect 1869 17493 1903 17527
rect 2037 17493 2071 17527
rect 2513 17493 2547 17527
rect 3157 17493 3191 17527
rect 3341 17493 3375 17527
rect 8217 17493 8251 17527
rect 12725 17493 12759 17527
rect 13369 17493 13403 17527
rect 14289 17493 14323 17527
rect 15945 17493 15979 17527
rect 16129 17493 16163 17527
rect 2973 17289 3007 17323
rect 9045 17289 9079 17323
rect 9229 17289 9263 17323
rect 10701 17289 10735 17323
rect 13093 17289 13127 17323
rect 13829 17289 13863 17323
rect 14473 17289 14507 17323
rect 15485 17289 15519 17323
rect 5181 17221 5215 17255
rect 5381 17221 5415 17255
rect 5733 17221 5767 17255
rect 9965 17221 9999 17255
rect 1593 17153 1627 17187
rect 1860 17153 1894 17187
rect 3157 17153 3191 17187
rect 3341 17153 3375 17187
rect 3433 17153 3467 17187
rect 3700 17153 3734 17187
rect 5641 17153 5675 17187
rect 5917 17153 5951 17187
rect 8493 17153 8527 17187
rect 9137 17153 9171 17187
rect 9443 17153 9477 17187
rect 9597 17153 9631 17187
rect 10149 17153 10183 17187
rect 10425 17153 10459 17187
rect 10609 17153 10643 17187
rect 10885 17153 10919 17187
rect 11161 17153 11195 17187
rect 13277 17153 13311 17187
rect 13645 17153 13679 17187
rect 14013 17153 14047 17187
rect 14105 17153 14139 17187
rect 14289 17153 14323 17187
rect 14657 17153 14691 17187
rect 14841 17153 14875 17187
rect 15025 17153 15059 17187
rect 15669 17153 15703 17187
rect 15761 17153 15795 17187
rect 15853 17153 15887 17187
rect 16037 17153 16071 17187
rect 8585 17085 8619 17119
rect 11253 17085 11287 17119
rect 8861 17017 8895 17051
rect 10333 17017 10367 17051
rect 13461 17017 13495 17051
rect 15209 17017 15243 17051
rect 3341 16949 3375 16983
rect 4813 16949 4847 16983
rect 5365 16949 5399 16983
rect 5549 16949 5583 16983
rect 6101 16949 6135 16983
rect 8493 16949 8527 16983
rect 14841 16949 14875 16983
rect 3617 16745 3651 16779
rect 5089 16745 5123 16779
rect 6745 16745 6779 16779
rect 9781 16745 9815 16779
rect 10425 16745 10459 16779
rect 3065 16677 3099 16711
rect 10793 16677 10827 16711
rect 1409 16609 1443 16643
rect 5273 16609 5307 16643
rect 10885 16609 10919 16643
rect 1665 16541 1699 16575
rect 3801 16541 3835 16575
rect 4077 16541 4111 16575
rect 4169 16541 4203 16575
rect 4813 16541 4847 16575
rect 4997 16541 5031 16575
rect 5181 16541 5215 16575
rect 5540 16541 5574 16575
rect 8125 16541 8159 16575
rect 9321 16541 9355 16575
rect 9505 16541 9539 16575
rect 10425 16541 10459 16575
rect 10517 16541 10551 16575
rect 10609 16541 10643 16575
rect 10701 16541 10735 16575
rect 13185 16541 13219 16575
rect 13277 16541 13311 16575
rect 13461 16541 13495 16575
rect 13553 16541 13587 16575
rect 13645 16541 13679 16575
rect 14105 16541 14139 16575
rect 15853 16541 15887 16575
rect 15945 16541 15979 16575
rect 16037 16541 16071 16575
rect 16221 16541 16255 16575
rect 3249 16473 3283 16507
rect 3985 16473 4019 16507
rect 7858 16473 7892 16507
rect 9597 16473 9631 16507
rect 9813 16473 9847 16507
rect 10977 16473 11011 16507
rect 11161 16473 11195 16507
rect 13921 16473 13955 16507
rect 14350 16473 14384 16507
rect 2789 16405 2823 16439
rect 3341 16405 3375 16439
rect 3433 16405 3467 16439
rect 4353 16405 4387 16439
rect 4537 16405 4571 16439
rect 6653 16405 6687 16439
rect 9413 16405 9447 16439
rect 9965 16405 9999 16439
rect 10149 16405 10183 16439
rect 11345 16405 11379 16439
rect 13093 16405 13127 16439
rect 15485 16405 15519 16439
rect 15577 16405 15611 16439
rect 3157 16201 3191 16235
rect 3525 16201 3559 16235
rect 3985 16201 4019 16235
rect 4445 16201 4479 16235
rect 6009 16201 6043 16235
rect 9137 16201 9171 16235
rect 9413 16201 9447 16235
rect 10885 16201 10919 16235
rect 11345 16201 11379 16235
rect 11529 16201 11563 16235
rect 12633 16201 12667 16235
rect 4997 16133 5031 16167
rect 5197 16133 5231 16167
rect 5825 16133 5859 16167
rect 7021 16133 7055 16167
rect 10977 16133 11011 16167
rect 11681 16133 11715 16167
rect 11897 16133 11931 16167
rect 12357 16133 12391 16167
rect 13093 16133 13127 16167
rect 14013 16133 14047 16167
rect 14381 16133 14415 16167
rect 15200 16133 15234 16167
rect 11207 16099 11241 16133
rect 1409 16065 1443 16099
rect 1676 16065 1710 16099
rect 2881 16065 2915 16099
rect 3065 16065 3099 16099
rect 3249 16065 3283 16099
rect 3433 16065 3467 16099
rect 3709 16065 3743 16099
rect 3893 16065 3927 16099
rect 4260 16065 4294 16099
rect 4353 16065 4387 16099
rect 4629 16065 4663 16099
rect 5457 16065 5491 16099
rect 7297 16065 7331 16099
rect 7481 16065 7515 16099
rect 8769 16065 8803 16099
rect 8953 16065 8987 16099
rect 9321 16065 9355 16099
rect 9597 16065 9631 16099
rect 9689 16065 9723 16099
rect 9873 16065 9907 16099
rect 10425 16065 10459 16099
rect 10517 16065 10551 16099
rect 12265 16065 12299 16099
rect 12817 16065 12851 16099
rect 12909 16065 12943 16099
rect 13369 16065 13403 16099
rect 13553 16065 13587 16099
rect 14197 16065 14231 16099
rect 14657 16065 14691 16099
rect 14749 16065 14783 16099
rect 4813 15997 4847 16031
rect 9781 15997 9815 16031
rect 10333 15997 10367 16031
rect 10609 15997 10643 16031
rect 14473 15997 14507 16031
rect 14933 15997 14967 16031
rect 2789 15929 2823 15963
rect 5365 15929 5399 15963
rect 6653 15929 6687 15963
rect 7665 15929 7699 15963
rect 13645 15929 13679 15963
rect 5181 15861 5215 15895
rect 5825 15861 5859 15895
rect 7021 15861 7055 15895
rect 7205 15861 7239 15895
rect 8953 15861 8987 15895
rect 10057 15861 10091 15895
rect 10333 15861 10367 15895
rect 10517 15861 10551 15895
rect 11161 15861 11195 15895
rect 11713 15861 11747 15895
rect 13185 15861 13219 15895
rect 16313 15861 16347 15895
rect 1593 15657 1627 15691
rect 1777 15657 1811 15691
rect 2789 15657 2823 15691
rect 3433 15657 3467 15691
rect 4721 15657 4755 15691
rect 5457 15657 5491 15691
rect 6653 15657 6687 15691
rect 8125 15657 8159 15691
rect 8309 15657 8343 15691
rect 9781 15657 9815 15691
rect 13001 15657 13035 15691
rect 13461 15657 13495 15691
rect 14289 15657 14323 15691
rect 14473 15657 14507 15691
rect 14749 15657 14783 15691
rect 2973 15589 3007 15623
rect 3065 15589 3099 15623
rect 4537 15589 4571 15623
rect 9137 15589 9171 15623
rect 15117 15589 15151 15623
rect 15761 15589 15795 15623
rect 2145 15521 2179 15555
rect 4721 15521 4755 15555
rect 4813 15521 4847 15555
rect 8033 15521 8067 15555
rect 9229 15521 9263 15555
rect 11529 15521 11563 15555
rect 2421 15453 2455 15487
rect 2697 15453 2731 15487
rect 3801 15453 3835 15487
rect 3985 15453 4019 15487
rect 4077 15453 4111 15487
rect 4169 15453 4203 15487
rect 4905 15453 4939 15487
rect 4997 15453 5031 15487
rect 5181 15453 5215 15487
rect 5641 15453 5675 15487
rect 5917 15453 5951 15487
rect 6010 15453 6044 15487
rect 6285 15453 6319 15487
rect 6382 15453 6416 15487
rect 7766 15453 7800 15487
rect 8677 15453 8711 15487
rect 8953 15453 8987 15487
rect 9045 15453 9079 15487
rect 9506 15453 9540 15487
rect 9643 15453 9677 15487
rect 9873 15453 9907 15487
rect 9965 15453 9999 15487
rect 10057 15453 10091 15487
rect 10241 15453 10275 15487
rect 10425 15453 10459 15487
rect 10517 15453 10551 15487
rect 10609 15453 10643 15487
rect 11161 15453 11195 15487
rect 11345 15453 11379 15487
rect 11437 15453 11471 15487
rect 11713 15453 11747 15487
rect 11989 15453 12023 15487
rect 12357 15453 12391 15487
rect 12633 15453 12667 15487
rect 14657 15453 14691 15487
rect 14933 15453 14967 15487
rect 15301 15453 15335 15487
rect 15393 15453 15427 15487
rect 15577 15453 15611 15487
rect 15669 15453 15703 15487
rect 15945 15453 15979 15487
rect 16037 15453 16071 15487
rect 16129 15453 16163 15487
rect 16313 15453 16347 15487
rect 1777 15385 1811 15419
rect 5825 15385 5859 15419
rect 6193 15385 6227 15419
rect 12173 15385 12207 15419
rect 12265 15385 12299 15419
rect 12817 15385 12851 15419
rect 13277 15385 13311 15419
rect 13461 15385 13495 15419
rect 14105 15385 14139 15419
rect 3433 15317 3467 15351
rect 3617 15317 3651 15351
rect 4445 15317 4479 15351
rect 5181 15317 5215 15351
rect 6561 15317 6595 15351
rect 8309 15317 8343 15351
rect 9321 15317 9355 15351
rect 10885 15317 10919 15351
rect 11897 15317 11931 15351
rect 12541 15317 12575 15351
rect 13645 15317 13679 15351
rect 14289 15317 14323 15351
rect 2053 15113 2087 15147
rect 2605 15113 2639 15147
rect 5733 15113 5767 15147
rect 6193 15113 6227 15147
rect 7849 15113 7883 15147
rect 9597 15113 9631 15147
rect 10609 15113 10643 15147
rect 12081 15113 12115 15147
rect 12633 15113 12667 15147
rect 14197 15113 14231 15147
rect 5089 15045 5123 15079
rect 5825 15045 5859 15079
rect 9965 15045 9999 15079
rect 10057 15045 10091 15079
rect 16221 15045 16255 15079
rect 1961 14977 1995 15011
rect 2145 14977 2179 15011
rect 2513 14977 2547 15011
rect 2697 14977 2731 15011
rect 5273 14977 5307 15011
rect 5549 14977 5583 15011
rect 6009 14977 6043 15011
rect 6469 14977 6503 15011
rect 6725 14977 6759 15011
rect 8217 14977 8251 15011
rect 8484 14977 8518 15011
rect 9689 14977 9723 15011
rect 9873 14977 9907 15011
rect 10175 14977 10209 15011
rect 10425 14977 10459 15011
rect 10609 14977 10643 15011
rect 10701 14977 10735 15011
rect 10885 14977 10919 15011
rect 10977 14977 11011 15011
rect 11069 14977 11103 15011
rect 11529 14977 11563 15011
rect 11713 14977 11747 15011
rect 11805 14977 11839 15011
rect 11897 14977 11931 15011
rect 12541 14977 12575 15011
rect 13001 14977 13035 15011
rect 14013 14977 14047 15011
rect 14657 14977 14691 15011
rect 14749 14977 14783 15011
rect 14841 14977 14875 15011
rect 15025 14977 15059 15011
rect 15393 14977 15427 15011
rect 15485 14977 15519 15011
rect 15577 14977 15611 15011
rect 15761 14977 15795 15011
rect 16037 14977 16071 15011
rect 5365 14909 5399 14943
rect 10333 14909 10367 14943
rect 12725 14909 12759 14943
rect 13553 14909 13587 14943
rect 13829 14909 13863 14943
rect 15853 14909 15887 14943
rect 11345 14841 11379 14875
rect 4905 14773 4939 14807
rect 12173 14773 12207 14807
rect 14381 14773 14415 14807
rect 15117 14773 15151 14807
rect 5641 14569 5675 14603
rect 10425 14569 10459 14603
rect 10701 14569 10735 14603
rect 11069 14569 11103 14603
rect 13645 14569 13679 14603
rect 14289 14569 14323 14603
rect 16313 14569 16347 14603
rect 8769 14501 8803 14535
rect 10057 14501 10091 14535
rect 10609 14501 10643 14535
rect 14197 14501 14231 14535
rect 4261 14433 4295 14467
rect 5733 14433 5767 14467
rect 9413 14433 9447 14467
rect 9597 14433 9631 14467
rect 10793 14433 10827 14467
rect 3341 14365 3375 14399
rect 4445 14365 4479 14399
rect 4537 14365 4571 14399
rect 5089 14365 5123 14399
rect 5457 14365 5491 14399
rect 6009 14365 6043 14399
rect 6193 14365 6227 14399
rect 6285 14365 6319 14399
rect 6469 14365 6503 14399
rect 6745 14365 6779 14399
rect 7849 14365 7883 14399
rect 8125 14365 8159 14399
rect 8309 14365 8343 14399
rect 8585 14365 8619 14399
rect 9321 14365 9355 14399
rect 10701 14365 10735 14399
rect 11161 14365 11195 14399
rect 11345 14365 11379 14399
rect 11437 14365 11471 14399
rect 11529 14365 11563 14399
rect 11805 14365 11839 14399
rect 13277 14365 13311 14399
rect 13737 14365 13771 14399
rect 14094 14359 14128 14393
rect 14473 14365 14507 14399
rect 14740 14365 14774 14399
rect 16129 14365 16163 14399
rect 12072 14297 12106 14331
rect 13461 14297 13495 14331
rect 14381 14297 14415 14331
rect 15945 14297 15979 14331
rect 3433 14229 3467 14263
rect 4537 14229 4571 14263
rect 5273 14229 5307 14263
rect 5825 14229 5859 14263
rect 6561 14229 6595 14263
rect 6929 14229 6963 14263
rect 8953 14229 8987 14263
rect 10425 14229 10459 14263
rect 11713 14229 11747 14263
rect 13185 14229 13219 14263
rect 13829 14229 13863 14263
rect 15853 14229 15887 14263
rect 4629 14025 4663 14059
rect 6929 14025 6963 14059
rect 9413 14025 9447 14059
rect 9781 14025 9815 14059
rect 10793 14025 10827 14059
rect 12817 14025 12851 14059
rect 14197 14025 14231 14059
rect 14473 14025 14507 14059
rect 16221 14025 16255 14059
rect 3709 13957 3743 13991
rect 14832 13957 14866 13991
rect 3939 13923 3973 13957
rect 1869 13889 1903 13923
rect 2053 13889 2087 13923
rect 3433 13889 3467 13923
rect 3617 13889 3651 13923
rect 4353 13889 4387 13923
rect 4537 13889 4571 13923
rect 5742 13889 5776 13923
rect 6009 13889 6043 13923
rect 6377 13889 6411 13923
rect 6929 13889 6963 13923
rect 7021 13889 7055 13923
rect 7849 13889 7883 13923
rect 8033 13889 8067 13923
rect 8300 13889 8334 13923
rect 9965 13889 9999 13923
rect 10149 13889 10183 13923
rect 10609 13889 10643 13923
rect 10977 13889 11011 13923
rect 11345 13889 11379 13923
rect 12725 13889 12759 13923
rect 13185 13889 13219 13923
rect 13921 13889 13955 13923
rect 14197 13889 14231 13923
rect 14289 13889 14323 13923
rect 16037 13889 16071 13923
rect 4169 13821 4203 13855
rect 10425 13821 10459 13855
rect 11529 13821 11563 13855
rect 12909 13821 12943 13855
rect 13829 13821 13863 13855
rect 14565 13821 14599 13855
rect 6653 13753 6687 13787
rect 6745 13753 6779 13787
rect 14105 13753 14139 13787
rect 1961 13685 1995 13719
rect 3525 13685 3559 13719
rect 3893 13685 3927 13719
rect 4077 13685 4111 13719
rect 6515 13685 6549 13719
rect 12173 13685 12207 13719
rect 12357 13685 12391 13719
rect 15945 13685 15979 13719
rect 7205 13481 7239 13515
rect 15393 13481 15427 13515
rect 15577 13481 15611 13515
rect 2789 13413 2823 13447
rect 3249 13413 3283 13447
rect 4169 13413 4203 13447
rect 13369 13413 13403 13447
rect 1409 13345 1443 13379
rect 3341 13345 3375 13379
rect 4077 13345 4111 13379
rect 5365 13345 5399 13379
rect 6101 13345 6135 13379
rect 7205 13345 7239 13379
rect 14657 13345 14691 13379
rect 2973 13277 3007 13311
rect 3525 13277 3559 13311
rect 3617 13277 3651 13311
rect 3801 13277 3835 13311
rect 3985 13277 4019 13311
rect 4261 13277 4295 13311
rect 4629 13277 4663 13311
rect 7297 13277 7331 13311
rect 8401 13277 8435 13311
rect 9873 13277 9907 13311
rect 10241 13277 10275 13311
rect 10333 13277 10367 13311
rect 10701 13277 10735 13311
rect 11253 13277 11287 13311
rect 11345 13277 11379 13311
rect 11621 13277 11655 13311
rect 11713 13277 11747 13311
rect 11989 13277 12023 13311
rect 12256 13277 12290 13311
rect 13921 13277 13955 13311
rect 15025 13277 15059 13311
rect 15209 13277 15243 13311
rect 15761 13277 15795 13311
rect 16129 13277 16163 13311
rect 1676 13209 1710 13243
rect 3249 13209 3283 13243
rect 3341 13209 3375 13243
rect 6837 13209 6871 13243
rect 10517 13209 10551 13243
rect 11529 13209 11563 13243
rect 14841 13209 14875 13243
rect 15853 13209 15887 13243
rect 15945 13209 15979 13243
rect 3065 13141 3099 13175
rect 4445 13141 4479 13175
rect 6745 13141 6779 13175
rect 7481 13141 7515 13175
rect 7849 13141 7883 13175
rect 10057 13141 10091 13175
rect 10425 13141 10459 13175
rect 11897 13141 11931 13175
rect 13737 13141 13771 13175
rect 14105 13141 14139 13175
rect 1593 12937 1627 12971
rect 1869 12937 1903 12971
rect 3433 12937 3467 12971
rect 4997 12937 5031 12971
rect 5825 12937 5859 12971
rect 6469 12937 6503 12971
rect 8217 12937 8251 12971
rect 8309 12937 8343 12971
rect 10425 12937 10459 12971
rect 10885 12937 10919 12971
rect 11897 12937 11931 12971
rect 12817 12937 12851 12971
rect 13645 12937 13679 12971
rect 15485 12937 15519 12971
rect 1777 12869 1811 12903
rect 2237 12869 2271 12903
rect 2421 12869 2455 12903
rect 2789 12869 2823 12903
rect 3893 12869 3927 12903
rect 4813 12869 4847 12903
rect 10793 12869 10827 12903
rect 1961 12801 1995 12835
rect 2605 12801 2639 12835
rect 2697 12801 2731 12835
rect 2973 12801 3007 12835
rect 3249 12801 3283 12835
rect 3709 12801 3743 12835
rect 3801 12801 3835 12835
rect 4077 12801 4111 12835
rect 4169 12801 4203 12835
rect 5089 12801 5123 12835
rect 5273 12801 5307 12835
rect 5641 12801 5675 12835
rect 6009 12801 6043 12835
rect 6193 12801 6227 12835
rect 6561 12801 6595 12835
rect 7766 12801 7800 12835
rect 8033 12801 8067 12835
rect 8125 12801 8159 12835
rect 9045 12801 9079 12835
rect 9505 12801 9539 12835
rect 11989 12801 12023 12835
rect 14105 12801 14139 12835
rect 14841 12801 14875 12835
rect 14933 12801 14967 12835
rect 15117 12801 15151 12835
rect 15301 12801 15335 12835
rect 15577 12801 15611 12835
rect 15761 12801 15795 12835
rect 15853 12801 15887 12835
rect 15945 12801 15979 12835
rect 2145 12733 2179 12767
rect 3065 12733 3099 12767
rect 5365 12733 5399 12767
rect 5457 12733 5491 12767
rect 6101 12733 6135 12767
rect 8585 12733 8619 12767
rect 9137 12733 9171 12767
rect 9321 12733 9355 12767
rect 10057 12733 10091 12767
rect 10977 12733 11011 12767
rect 12081 12733 12115 12767
rect 12909 12733 12943 12767
rect 13093 12733 13127 12767
rect 13737 12733 13771 12767
rect 13829 12733 13863 12767
rect 14657 12733 14691 12767
rect 2973 12665 3007 12699
rect 4445 12665 4479 12699
rect 6653 12665 6687 12699
rect 13277 12665 13311 12699
rect 16129 12665 16163 12699
rect 3525 12597 3559 12631
rect 4813 12597 4847 12631
rect 8677 12597 8711 12631
rect 11529 12597 11563 12631
rect 12449 12597 12483 12631
rect 2053 12393 2087 12427
rect 3157 12393 3191 12427
rect 6285 12393 6319 12427
rect 8217 12393 8251 12427
rect 9229 12393 9263 12427
rect 10057 12393 10091 12427
rect 11713 12393 11747 12427
rect 3525 12325 3559 12359
rect 4169 12325 4203 12359
rect 13369 12325 13403 12359
rect 3617 12257 3651 12291
rect 9781 12257 9815 12291
rect 11989 12257 12023 12291
rect 1685 12189 1719 12223
rect 1777 12189 1811 12223
rect 2513 12189 2547 12223
rect 2605 12189 2639 12223
rect 3341 12189 3375 12223
rect 4537 12189 4571 12223
rect 4813 12189 4847 12223
rect 6469 12189 6503 12223
rect 6745 12189 6779 12223
rect 6837 12189 6871 12223
rect 8493 12189 8527 12223
rect 9137 12189 9171 12223
rect 9597 12189 9631 12223
rect 11181 12189 11215 12223
rect 11437 12189 11471 12223
rect 11897 12189 11931 12223
rect 13461 12189 13495 12223
rect 14105 12189 14139 12223
rect 15393 12189 15427 12223
rect 15485 12189 15519 12223
rect 15577 12189 15611 12223
rect 15761 12189 15795 12223
rect 1501 12121 1535 12155
rect 1869 12121 1903 12155
rect 2069 12121 2103 12155
rect 2697 12121 2731 12155
rect 2881 12121 2915 12155
rect 4353 12121 4387 12155
rect 4721 12121 4755 12155
rect 5080 12121 5114 12155
rect 7104 12121 7138 12155
rect 8309 12121 8343 12155
rect 12256 12121 12290 12155
rect 14841 12121 14875 12155
rect 15853 12121 15887 12155
rect 16037 12121 16071 12155
rect 1599 12053 1633 12087
rect 2237 12053 2271 12087
rect 2329 12053 2363 12087
rect 4445 12053 4479 12087
rect 6193 12053 6227 12087
rect 6653 12053 6687 12087
rect 8677 12053 8711 12087
rect 9045 12053 9079 12087
rect 9689 12053 9723 12087
rect 15117 12053 15151 12087
rect 16221 12053 16255 12087
rect 1409 11849 1443 11883
rect 3525 11849 3559 11883
rect 4353 11849 4387 11883
rect 4997 11849 5031 11883
rect 6009 11849 6043 11883
rect 7139 11849 7173 11883
rect 9965 11849 9999 11883
rect 13645 11849 13679 11883
rect 3049 11781 3083 11815
rect 3249 11781 3283 11815
rect 5181 11781 5215 11815
rect 6929 11781 6963 11815
rect 8116 11781 8150 11815
rect 9873 11781 9907 11815
rect 11100 11781 11134 11815
rect 12348 11781 12382 11815
rect 2533 11713 2567 11747
rect 2789 11713 2823 11747
rect 3433 11713 3467 11747
rect 3801 11713 3835 11747
rect 4077 11713 4111 11747
rect 4169 11713 4203 11747
rect 4445 11713 4479 11747
rect 4629 11713 4663 11747
rect 5549 11713 5583 11747
rect 5825 11713 5859 11747
rect 6101 11713 6135 11747
rect 6653 11713 6687 11747
rect 7849 11713 7883 11747
rect 9321 11713 9355 11747
rect 9505 11713 9539 11747
rect 11345 11713 11379 11747
rect 12081 11713 12115 11747
rect 13829 11713 13863 11747
rect 14013 11713 14047 11747
rect 14105 11713 14139 11747
rect 14381 11713 14415 11747
rect 14565 11713 14599 11747
rect 14933 11713 14967 11747
rect 15189 11713 15223 11747
rect 2881 11577 2915 11611
rect 3893 11577 3927 11611
rect 6837 11577 6871 11611
rect 7297 11577 7331 11611
rect 13461 11577 13495 11611
rect 3065 11509 3099 11543
rect 4445 11509 4479 11543
rect 5181 11509 5215 11543
rect 5641 11509 5675 11543
rect 7113 11509 7147 11543
rect 9229 11509 9263 11543
rect 14289 11509 14323 11543
rect 14749 11509 14783 11543
rect 16313 11509 16347 11543
rect 2789 11305 2823 11339
rect 2881 11305 2915 11339
rect 5273 11305 5307 11339
rect 5457 11305 5491 11339
rect 8585 11305 8619 11339
rect 8953 11305 8987 11339
rect 9781 11305 9815 11339
rect 9965 11305 9999 11339
rect 13369 11305 13403 11339
rect 14841 11305 14875 11339
rect 4445 11237 4479 11271
rect 8769 11237 8803 11271
rect 16313 11237 16347 11271
rect 4721 11169 4755 11203
rect 9347 11169 9381 11203
rect 13921 11169 13955 11203
rect 14933 11169 14967 11203
rect 1409 11101 1443 11135
rect 2881 11101 2915 11135
rect 3065 11101 3099 11135
rect 4353 11101 4387 11135
rect 4537 11101 4571 11135
rect 4629 11101 4663 11135
rect 4813 11101 4847 11135
rect 9137 11101 9171 11135
rect 9505 11101 9539 11135
rect 11713 11101 11747 11135
rect 13277 11101 13311 11135
rect 13461 11101 13495 11135
rect 13737 11101 13771 11135
rect 14197 11101 14231 11135
rect 14381 11101 14415 11135
rect 14473 11101 14507 11135
rect 14565 11101 14599 11135
rect 15200 11101 15234 11135
rect 1676 11033 1710 11067
rect 5441 11033 5475 11067
rect 5641 11033 5675 11067
rect 8401 11033 8435 11067
rect 9597 11033 9631 11067
rect 12449 11033 12483 11067
rect 13553 11033 13587 11067
rect 8611 10965 8645 10999
rect 9797 10965 9831 10999
rect 1685 10761 1719 10795
rect 7481 10761 7515 10795
rect 13645 10761 13679 10795
rect 16313 10761 16347 10795
rect 1853 10693 1887 10727
rect 2053 10693 2087 10727
rect 2421 10693 2455 10727
rect 5733 10693 5767 10727
rect 7665 10693 7699 10727
rect 9137 10693 9171 10727
rect 14841 10693 14875 10727
rect 15178 10693 15212 10727
rect 2237 10625 2271 10659
rect 2513 10625 2547 10659
rect 2697 10625 2731 10659
rect 4077 10625 4111 10659
rect 4721 10625 4755 10659
rect 4997 10625 5031 10659
rect 5365 10625 5399 10659
rect 5549 10625 5583 10659
rect 7389 10625 7423 10659
rect 8309 10625 8343 10659
rect 8493 10625 8527 10659
rect 9321 10625 9355 10659
rect 9689 10625 9723 10659
rect 12081 10625 12115 10659
rect 13461 10625 13495 10659
rect 13829 10625 13863 10659
rect 14105 10625 14139 10659
rect 14197 10625 14231 10659
rect 14381 10625 14415 10659
rect 14473 10625 14507 10659
rect 14565 10625 14599 10659
rect 2605 10557 2639 10591
rect 9413 10557 9447 10591
rect 14933 10557 14967 10591
rect 4077 10489 4111 10523
rect 9505 10489 9539 10523
rect 13277 10489 13311 10523
rect 1869 10421 1903 10455
rect 5917 10421 5951 10455
rect 7665 10421 7699 10455
rect 8493 10421 8527 10455
rect 8953 10421 8987 10455
rect 9597 10421 9631 10455
rect 13921 10421 13955 10455
rect 3157 10217 3191 10251
rect 5273 10217 5307 10251
rect 7113 10217 7147 10251
rect 7297 10217 7331 10251
rect 8033 10217 8067 10251
rect 8769 10217 8803 10251
rect 13001 10217 13035 10251
rect 16221 10217 16255 10251
rect 8125 10149 8159 10183
rect 8953 10149 8987 10183
rect 4353 10081 4387 10115
rect 9505 10081 9539 10115
rect 3341 10013 3375 10047
rect 3617 10013 3651 10047
rect 5181 10013 5215 10047
rect 6653 10013 6687 10047
rect 6745 10013 6779 10047
rect 7389 10013 7423 10047
rect 8125 10013 8159 10047
rect 8401 10013 8435 10047
rect 8585 10013 8619 10047
rect 8769 10013 8803 10047
rect 10517 10013 10551 10047
rect 11161 10013 11195 10047
rect 13185 10013 13219 10047
rect 13553 10013 13587 10047
rect 13645 10013 13679 10047
rect 13737 10013 13771 10047
rect 13921 10013 13955 10047
rect 14105 10013 14139 10047
rect 15577 10013 15611 10047
rect 16037 10013 16071 10047
rect 3525 9945 3559 9979
rect 3985 9945 4019 9979
rect 6386 9945 6420 9979
rect 7113 9945 7147 9979
rect 11428 9945 11462 9979
rect 14350 9945 14384 9979
rect 15761 9945 15795 9979
rect 15945 9945 15979 9979
rect 4077 9877 4111 9911
rect 8309 9877 8343 9911
rect 9873 9877 9907 9911
rect 12541 9877 12575 9911
rect 13277 9877 13311 9911
rect 15485 9877 15519 9911
rect 3065 9673 3099 9707
rect 3709 9673 3743 9707
rect 4169 9673 4203 9707
rect 4445 9673 4479 9707
rect 6377 9673 6411 9707
rect 6929 9673 6963 9707
rect 9045 9673 9079 9707
rect 12909 9673 12943 9707
rect 4077 9605 4111 9639
rect 4286 9605 4320 9639
rect 6529 9605 6563 9639
rect 6745 9605 6779 9639
rect 14841 9605 14875 9639
rect 15393 9605 15427 9639
rect 15761 9605 15795 9639
rect 15853 9605 15887 9639
rect 2789 9537 2823 9571
rect 2881 9537 2915 9571
rect 3341 9537 3375 9571
rect 4813 9537 4847 9571
rect 6009 9537 6043 9571
rect 8053 9537 8087 9571
rect 8309 9537 8343 9571
rect 9321 9537 9355 9571
rect 9781 9537 9815 9571
rect 10048 9537 10082 9571
rect 11529 9537 11563 9571
rect 11796 9537 11830 9571
rect 13093 9537 13127 9571
rect 13360 9537 13394 9571
rect 14749 9537 14783 9571
rect 14933 9537 14967 9571
rect 15117 9537 15151 9571
rect 15577 9537 15611 9571
rect 16037 9537 16071 9571
rect 3065 9469 3099 9503
rect 3433 9469 3467 9503
rect 3801 9469 3835 9503
rect 5549 9469 5583 9503
rect 8401 9469 8435 9503
rect 9597 9469 9631 9503
rect 5733 9401 5767 9435
rect 9137 9401 9171 9435
rect 14565 9401 14599 9435
rect 6561 9333 6595 9367
rect 9505 9333 9539 9367
rect 11161 9333 11195 9367
rect 14473 9333 14507 9367
rect 16221 9333 16255 9367
rect 1961 9129 1995 9163
rect 3617 9129 3651 9163
rect 3985 9129 4019 9163
rect 4537 9129 4571 9163
rect 4997 9129 5031 9163
rect 8309 9129 8343 9163
rect 8585 9129 8619 9163
rect 11437 9129 11471 9163
rect 13461 9129 13495 9163
rect 16221 9129 16255 9163
rect 2513 9061 2547 9095
rect 8769 9061 8803 9095
rect 3985 8993 4019 9027
rect 11989 8993 12023 9027
rect 2237 8925 2271 8959
rect 3249 8925 3283 8959
rect 3801 8925 3835 8959
rect 4077 8925 4111 8959
rect 4721 8925 4755 8959
rect 4813 8925 4847 8959
rect 5089 8925 5123 8959
rect 5457 8925 5491 8959
rect 6837 8925 6871 8959
rect 6929 8925 6963 8959
rect 7196 8925 7230 8959
rect 8953 8925 8987 8959
rect 11345 8925 11379 8959
rect 13369 8925 13403 8959
rect 13461 8925 13495 8959
rect 13553 8925 13587 8959
rect 14289 8925 14323 8959
rect 15117 8925 15151 8959
rect 15209 8925 15243 8959
rect 15301 8925 15335 8959
rect 15485 8925 15519 8959
rect 15761 8925 15795 8959
rect 16037 8925 16071 8959
rect 1929 8857 1963 8891
rect 2145 8857 2179 8891
rect 2513 8857 2547 8891
rect 3433 8857 3467 8891
rect 6101 8857 6135 8891
rect 8401 8857 8435 8891
rect 9198 8857 9232 8891
rect 10517 8857 10551 8891
rect 11805 8857 11839 8891
rect 12541 8857 12575 8891
rect 14473 8857 14507 8891
rect 15577 8857 15611 8891
rect 15945 8857 15979 8891
rect 1777 8789 1811 8823
rect 2329 8789 2363 8823
rect 4261 8789 4295 8823
rect 8601 8789 8635 8823
rect 10333 8789 10367 8823
rect 11897 8789 11931 8823
rect 13829 8789 13863 8823
rect 14105 8789 14139 8823
rect 14841 8789 14875 8823
rect 1409 8585 1443 8619
rect 4353 8585 4387 8619
rect 5013 8585 5047 8619
rect 5273 8585 5307 8619
rect 8309 8585 8343 8619
rect 9781 8585 9815 8619
rect 10425 8585 10459 8619
rect 10793 8585 10827 8619
rect 12541 8585 12575 8619
rect 13001 8585 13035 8619
rect 13369 8585 13403 8619
rect 16313 8585 16347 8619
rect 2881 8517 2915 8551
rect 3081 8517 3115 8551
rect 4537 8517 4571 8551
rect 4813 8517 4847 8551
rect 6377 8517 6411 8551
rect 7196 8517 7230 8551
rect 12173 8517 12207 8551
rect 15178 8517 15212 8551
rect 2522 8449 2556 8483
rect 2789 8449 2823 8483
rect 3341 8449 3375 8483
rect 3525 8449 3559 8483
rect 4721 8449 4755 8483
rect 5457 8449 5491 8483
rect 5641 8449 5675 8483
rect 5733 8449 5767 8483
rect 6561 8449 6595 8483
rect 8401 8449 8435 8483
rect 8657 8449 8691 8483
rect 9873 8449 9907 8483
rect 10885 8449 10919 8483
rect 12081 8449 12115 8483
rect 12909 8449 12943 8483
rect 13645 8449 13679 8483
rect 13737 8449 13771 8483
rect 13829 8449 13863 8483
rect 14013 8449 14047 8483
rect 14197 8449 14231 8483
rect 14381 8449 14415 8483
rect 14473 8449 14507 8483
rect 14565 8449 14599 8483
rect 6745 8381 6779 8415
rect 6929 8381 6963 8415
rect 10977 8381 11011 8415
rect 12357 8381 12391 8415
rect 13093 8381 13127 8415
rect 14933 8381 14967 8415
rect 3249 8313 3283 8347
rect 3341 8313 3375 8347
rect 5181 8313 5215 8347
rect 5549 8313 5583 8347
rect 14841 8313 14875 8347
rect 3065 8245 3099 8279
rect 4997 8245 5031 8279
rect 11713 8245 11747 8279
rect 2973 8041 3007 8075
rect 5365 8041 5399 8075
rect 6469 8041 6503 8075
rect 8125 8041 8159 8075
rect 8953 8041 8987 8075
rect 9321 8041 9355 8075
rect 9505 8041 9539 8075
rect 11069 8041 11103 8075
rect 11345 8041 11379 8075
rect 13277 8041 13311 8075
rect 16313 8041 16347 8075
rect 3065 7973 3099 8007
rect 3617 7973 3651 8007
rect 4077 7973 4111 8007
rect 5733 7973 5767 8007
rect 5825 7973 5859 8007
rect 12909 7973 12943 8007
rect 1593 7905 1627 7939
rect 6929 7905 6963 7939
rect 8677 7905 8711 7939
rect 9229 7905 9263 7939
rect 11529 7905 11563 7939
rect 14933 7905 14967 7939
rect 1860 7837 1894 7871
rect 3433 7837 3467 7871
rect 3801 7837 3835 7871
rect 3893 7837 3927 7871
rect 4169 7837 4203 7871
rect 4353 7837 4387 7871
rect 6193 7837 6227 7871
rect 6653 7837 6687 7871
rect 6745 7837 6779 7871
rect 6837 7837 6871 7871
rect 7481 7837 7515 7871
rect 7849 7837 7883 7871
rect 8033 7837 8067 7871
rect 9321 7837 9355 7871
rect 10885 7837 10919 7871
rect 10977 7837 11011 7871
rect 11161 7837 11195 7871
rect 11796 7837 11830 7871
rect 13277 7837 13311 7871
rect 13645 7837 13679 7871
rect 14105 7837 14139 7871
rect 14289 7837 14323 7871
rect 14381 7837 14415 7871
rect 14473 7837 14507 7871
rect 15200 7837 15234 7871
rect 3249 7769 3283 7803
rect 4077 7769 4111 7803
rect 6377 7769 6411 7803
rect 7297 7769 7331 7803
rect 10618 7769 10652 7803
rect 3341 7701 3375 7735
rect 4261 7701 4295 7735
rect 5181 7701 5215 7735
rect 5365 7701 5399 7735
rect 6009 7701 6043 7735
rect 6101 7701 6135 7735
rect 7113 7701 7147 7735
rect 8033 7701 8067 7735
rect 13093 7701 13127 7735
rect 14749 7701 14783 7735
rect 3065 7497 3099 7531
rect 3157 7497 3191 7531
rect 3325 7497 3359 7531
rect 4721 7497 4755 7531
rect 6193 7497 6227 7531
rect 8125 7497 8159 7531
rect 16221 7497 16255 7531
rect 1501 7429 1535 7463
rect 1952 7429 1986 7463
rect 3525 7429 3559 7463
rect 4629 7429 4663 7463
rect 1409 7361 1443 7395
rect 1593 7361 1627 7395
rect 1685 7361 1719 7395
rect 3709 7361 3743 7395
rect 3893 7361 3927 7395
rect 3985 7361 4019 7395
rect 4077 7361 4111 7395
rect 4445 7361 4479 7395
rect 4721 7361 4755 7395
rect 4813 7361 4847 7395
rect 5080 7361 5114 7395
rect 6377 7361 6411 7395
rect 6644 7361 6678 7395
rect 7849 7361 7883 7395
rect 7941 7361 7975 7395
rect 8401 7361 8435 7395
rect 9045 7361 9079 7395
rect 9301 7361 9335 7395
rect 10517 7361 10551 7395
rect 11161 7361 11195 7395
rect 11529 7361 11563 7395
rect 11785 7361 11819 7395
rect 13093 7361 13127 7395
rect 13349 7361 13383 7395
rect 15678 7361 15712 7395
rect 15945 7361 15979 7395
rect 16037 7361 16071 7395
rect 8125 7293 8159 7327
rect 8493 7293 8527 7327
rect 4353 7225 4387 7259
rect 8769 7225 8803 7259
rect 12909 7225 12943 7259
rect 3341 7157 3375 7191
rect 7757 7157 7791 7191
rect 10425 7157 10459 7191
rect 14473 7157 14507 7191
rect 14565 7157 14599 7191
rect 2329 6953 2363 6987
rect 2973 6953 3007 6987
rect 3157 6953 3191 6987
rect 3433 6953 3467 6987
rect 5181 6953 5215 6987
rect 6929 6953 6963 6987
rect 7021 6953 7055 6987
rect 7205 6953 7239 6987
rect 11345 6953 11379 6987
rect 11529 6953 11563 6987
rect 13001 6953 13035 6987
rect 14657 6953 14691 6987
rect 1777 6817 1811 6851
rect 2053 6817 2087 6851
rect 3801 6817 3835 6851
rect 9229 6817 9263 6851
rect 10609 6817 10643 6851
rect 11186 6817 11220 6851
rect 12173 6817 12207 6851
rect 14933 6817 14967 6851
rect 1685 6749 1719 6783
rect 4068 6749 4102 6783
rect 5273 6749 5307 6783
rect 5457 6749 5491 6783
rect 5549 6749 5583 6783
rect 7849 6749 7883 6783
rect 8033 6749 8067 6783
rect 9873 6749 9907 6783
rect 10701 6749 10735 6783
rect 10977 6749 11011 6783
rect 12909 6749 12943 6783
rect 13277 6749 13311 6783
rect 13369 6749 13403 6783
rect 13461 6749 13495 6783
rect 13645 6749 13679 6783
rect 14105 6749 14139 6783
rect 14289 6749 14323 6783
rect 14473 6749 14507 6783
rect 2145 6681 2179 6715
rect 2345 6681 2379 6715
rect 2789 6681 2823 6715
rect 2989 6681 3023 6715
rect 3249 6681 3283 6715
rect 5365 6681 5399 6715
rect 5816 6681 5850 6715
rect 7173 6681 7207 6715
rect 7389 6681 7423 6715
rect 7941 6681 7975 6715
rect 11069 6681 11103 6715
rect 11989 6681 12023 6715
rect 14381 6681 14415 6715
rect 15200 6681 15234 6715
rect 2513 6613 2547 6647
rect 3449 6613 3483 6647
rect 3617 6613 3651 6647
rect 9965 6613 9999 6647
rect 11897 6613 11931 6647
rect 12725 6613 12759 6647
rect 16313 6613 16347 6647
rect 6377 6409 6411 6443
rect 6745 6409 6779 6443
rect 9505 6409 9539 6443
rect 10333 6409 10367 6443
rect 11161 6409 11195 6443
rect 11345 6409 11379 6443
rect 12081 6409 12115 6443
rect 13553 6409 13587 6443
rect 14105 6409 14139 6443
rect 14749 6409 14783 6443
rect 15577 6409 15611 6443
rect 15669 6409 15703 6443
rect 3494 6341 3528 6375
rect 4873 6341 4907 6375
rect 5089 6341 5123 6375
rect 5917 6341 5951 6375
rect 10501 6341 10535 6375
rect 10701 6341 10735 6375
rect 14473 6341 14507 6375
rect 15945 6341 15979 6375
rect 2789 6273 2823 6307
rect 3249 6273 3283 6307
rect 6561 6273 6595 6307
rect 6837 6273 6871 6307
rect 9505 6273 9539 6307
rect 9689 6273 9723 6307
rect 9781 6273 9815 6307
rect 9873 6273 9907 6307
rect 10793 6273 10827 6307
rect 11529 6273 11563 6307
rect 12633 6273 12667 6307
rect 13001 6273 13035 6307
rect 13277 6273 13311 6307
rect 13461 6273 13495 6307
rect 13737 6273 13771 6307
rect 13921 6273 13955 6307
rect 14289 6273 14323 6307
rect 14565 6273 14599 6307
rect 14933 6273 14967 6307
rect 15117 6276 15151 6310
rect 15212 6273 15246 6307
rect 15347 6273 15381 6307
rect 15853 6273 15887 6307
rect 16037 6273 16071 6307
rect 16221 6273 16255 6307
rect 2881 6205 2915 6239
rect 3157 6205 3191 6239
rect 10057 6205 10091 6239
rect 11805 6205 11839 6239
rect 5641 6137 5675 6171
rect 12449 6137 12483 6171
rect 4629 6069 4663 6103
rect 4721 6069 4755 6103
rect 4905 6069 4939 6103
rect 5457 6069 5491 6103
rect 9965 6069 9999 6103
rect 10517 6069 10551 6103
rect 11161 6069 11195 6103
rect 11713 6069 11747 6103
rect 12817 6069 12851 6103
rect 13093 6069 13127 6103
rect 3801 5865 3835 5899
rect 6653 5865 6687 5899
rect 10609 5865 10643 5899
rect 11989 5865 12023 5899
rect 12633 5865 12667 5899
rect 14749 5797 14783 5831
rect 5181 5661 5215 5695
rect 5273 5661 5307 5695
rect 5540 5661 5574 5695
rect 10517 5661 10551 5695
rect 10701 5661 10735 5695
rect 10793 5661 10827 5695
rect 10977 5661 11011 5695
rect 11345 5661 11379 5695
rect 12173 5661 12207 5695
rect 12541 5661 12575 5695
rect 12817 5661 12851 5695
rect 13277 5661 13311 5695
rect 14105 5661 14139 5695
rect 14289 5661 14323 5695
rect 14381 5661 14415 5695
rect 14473 5661 14507 5695
rect 14933 5661 14967 5695
rect 15117 5661 15151 5695
rect 15301 5661 15335 5695
rect 15761 5661 15795 5695
rect 15853 5661 15887 5695
rect 15945 5661 15979 5695
rect 16129 5661 16163 5695
rect 4914 5593 4948 5627
rect 13001 5593 13035 5627
rect 13093 5593 13127 5627
rect 13553 5593 13587 5627
rect 13737 5593 13771 5627
rect 13921 5593 13955 5627
rect 15025 5593 15059 5627
rect 10885 5525 10919 5559
rect 11437 5525 11471 5559
rect 12357 5525 12391 5559
rect 13461 5525 13495 5559
rect 14657 5525 14691 5559
rect 15485 5525 15519 5559
rect 10057 5321 10091 5355
rect 11989 5321 12023 5355
rect 12817 5321 12851 5355
rect 14013 5321 14047 5355
rect 10609 5253 10643 5287
rect 9965 5185 9999 5219
rect 10149 5185 10183 5219
rect 10425 5185 10459 5219
rect 10793 5185 10827 5219
rect 11161 5185 11195 5219
rect 12909 5185 12943 5219
rect 13553 5185 13587 5219
rect 13645 5185 13679 5219
rect 13737 5185 13771 5219
rect 13921 5185 13955 5219
rect 15025 5185 15059 5219
rect 15117 5185 15151 5219
rect 15209 5185 15243 5219
rect 15393 5185 15427 5219
rect 15761 5185 15795 5219
rect 15853 5185 15887 5219
rect 15945 5185 15979 5219
rect 16129 5185 16163 5219
rect 12081 5117 12115 5151
rect 12173 5117 12207 5151
rect 13001 5117 13035 5151
rect 14565 5117 14599 5151
rect 10241 5049 10275 5083
rect 11345 5049 11379 5083
rect 11161 4981 11195 5015
rect 11621 4981 11655 5015
rect 12449 4981 12483 5015
rect 13277 4981 13311 5015
rect 14749 4981 14783 5015
rect 15485 4981 15519 5015
rect 9045 4777 9079 4811
rect 11161 4777 11195 4811
rect 12817 4777 12851 4811
rect 14105 4777 14139 4811
rect 9229 4641 9263 4675
rect 13553 4641 13587 4675
rect 8953 4573 8987 4607
rect 9413 4573 9447 4607
rect 9505 4573 9539 4607
rect 9781 4573 9815 4607
rect 11437 4573 11471 4607
rect 11704 4573 11738 4607
rect 13461 4573 13495 4607
rect 15485 4573 15519 4607
rect 15853 4573 15887 4607
rect 15945 4573 15979 4607
rect 16037 4573 16071 4607
rect 16221 4573 16255 4607
rect 9689 4505 9723 4539
rect 10026 4505 10060 4539
rect 13369 4505 13403 4539
rect 15218 4505 15252 4539
rect 9229 4437 9263 4471
rect 13001 4437 13035 4471
rect 15577 4437 15611 4471
rect 11621 4233 11655 4267
rect 8217 4165 8251 4199
rect 9229 4165 9263 4199
rect 9321 4165 9355 4199
rect 9459 4165 9493 4199
rect 12756 4165 12790 4199
rect 8401 4097 8435 4131
rect 8493 4097 8527 4131
rect 8677 4097 8711 4131
rect 9137 4097 9171 4131
rect 9597 4097 9631 4131
rect 10140 4097 10174 4131
rect 13001 4097 13035 4131
rect 13093 4097 13127 4131
rect 13360 4097 13394 4131
rect 15770 4097 15804 4131
rect 16037 4097 16071 4131
rect 8861 4029 8895 4063
rect 9873 4029 9907 4063
rect 11253 3961 11287 3995
rect 14657 3961 14691 3995
rect 8033 3893 8067 3927
rect 8953 3893 8987 3927
rect 14473 3893 14507 3927
rect 9781 3689 9815 3723
rect 11253 3689 11287 3723
rect 11529 3689 11563 3723
rect 11713 3689 11747 3723
rect 13369 3689 13403 3723
rect 16313 3689 16347 3723
rect 9873 3553 9907 3587
rect 11989 3553 12023 3587
rect 13829 3553 13863 3587
rect 14933 3553 14967 3587
rect 8769 3485 8803 3519
rect 9229 3485 9263 3519
rect 10129 3485 10163 3519
rect 13461 3485 13495 3519
rect 14381 3485 14415 3519
rect 14473 3485 14507 3519
rect 14565 3485 14599 3519
rect 14749 3485 14783 3519
rect 15200 3485 15234 3519
rect 11345 3417 11379 3451
rect 11545 3417 11579 3451
rect 12256 3417 12290 3451
rect 13645 3417 13679 3451
rect 8585 3349 8619 3383
rect 14105 3349 14139 3383
rect 9413 3145 9447 3179
rect 10425 3145 10459 3179
rect 10793 3145 10827 3179
rect 14105 3145 14139 3179
rect 14841 3145 14875 3179
rect 8300 3077 8334 3111
rect 14657 3077 14691 3111
rect 15200 3077 15234 3111
rect 8033 3009 8067 3043
rect 12725 3009 12759 3043
rect 12992 3009 13026 3043
rect 14197 3009 14231 3043
rect 14473 3009 14507 3043
rect 14933 3009 14967 3043
rect 10885 2941 10919 2975
rect 10977 2941 11011 2975
rect 14381 2805 14415 2839
rect 16313 2805 16347 2839
rect 14841 2601 14875 2635
rect 15209 2601 15243 2635
rect 15761 2601 15795 2635
rect 16221 2601 16255 2635
rect 8401 2533 8435 2567
rect 10057 2533 10091 2567
rect 7481 2465 7515 2499
rect 7205 2397 7239 2431
rect 8769 2397 8803 2431
rect 9413 2397 9447 2431
rect 13277 2397 13311 2431
rect 13921 2397 13955 2431
rect 14565 2397 14599 2431
rect 14657 2397 14691 2431
rect 15025 2397 15059 2431
rect 15393 2397 15427 2431
rect 15577 2397 15611 2431
rect 16037 2397 16071 2431
rect 8217 2329 8251 2363
rect 9873 2329 9907 2363
rect 8585 2261 8619 2295
rect 9229 2261 9263 2295
rect 13093 2261 13127 2295
rect 13737 2261 13771 2295
rect 14381 2261 14415 2295
<< metal1 >>
rect 1104 33210 16652 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 16652 33210
rect 1104 33136 16652 33158
rect 7742 33056 7748 33108
rect 7800 33096 7806 33108
rect 7929 33099 7987 33105
rect 7929 33096 7941 33099
rect 7800 33068 7941 33096
rect 7800 33056 7806 33068
rect 7929 33065 7941 33068
rect 7975 33065 7987 33099
rect 7929 33059 7987 33065
rect 11701 33099 11759 33105
rect 11701 33065 11713 33099
rect 11747 33096 11759 33099
rect 12894 33096 12900 33108
rect 11747 33068 12900 33096
rect 11747 33065 11759 33068
rect 11701 33059 11759 33065
rect 12894 33056 12900 33068
rect 12952 33056 12958 33108
rect 12986 33056 12992 33108
rect 13044 33096 13050 33108
rect 13725 33099 13783 33105
rect 13044 33068 13676 33096
rect 13044 33056 13050 33068
rect 11149 33031 11207 33037
rect 11149 32997 11161 33031
rect 11195 33028 11207 33031
rect 13538 33028 13544 33040
rect 11195 33000 13544 33028
rect 11195 32997 11207 33000
rect 11149 32991 11207 32997
rect 13538 32988 13544 33000
rect 13596 32988 13602 33040
rect 13648 33028 13676 33068
rect 13725 33065 13737 33099
rect 13771 33096 13783 33099
rect 14826 33096 14832 33108
rect 13771 33068 14832 33096
rect 13771 33065 13783 33068
rect 13725 33059 13783 33065
rect 14826 33056 14832 33068
rect 14884 33056 14890 33108
rect 15286 33056 15292 33108
rect 15344 33096 15350 33108
rect 16482 33096 16488 33108
rect 15344 33068 16488 33096
rect 15344 33056 15350 33068
rect 16482 33056 16488 33068
rect 16540 33056 16546 33108
rect 13648 33000 15608 33028
rect 15470 32960 15476 32972
rect 12084 32932 15476 32960
rect 8110 32852 8116 32904
rect 8168 32852 8174 32904
rect 10594 32852 10600 32904
rect 10652 32852 10658 32904
rect 10870 32852 10876 32904
rect 10928 32892 10934 32904
rect 10965 32895 11023 32901
rect 10965 32892 10977 32895
rect 10928 32864 10977 32892
rect 10928 32852 10934 32864
rect 10965 32861 10977 32864
rect 11011 32861 11023 32895
rect 10965 32855 11023 32861
rect 11330 32852 11336 32904
rect 11388 32852 11394 32904
rect 11514 32852 11520 32904
rect 11572 32852 11578 32904
rect 10410 32716 10416 32768
rect 10468 32716 10474 32768
rect 10778 32716 10784 32768
rect 10836 32716 10842 32768
rect 11977 32759 12035 32765
rect 11977 32725 11989 32759
rect 12023 32756 12035 32759
rect 12084 32756 12112 32932
rect 15470 32920 15476 32932
rect 15528 32920 15534 32972
rect 12161 32895 12219 32901
rect 12161 32861 12173 32895
rect 12207 32861 12219 32895
rect 12161 32855 12219 32861
rect 12713 32895 12771 32901
rect 12713 32861 12725 32895
rect 12759 32892 12771 32895
rect 12759 32864 13860 32892
rect 12759 32861 12771 32864
rect 12713 32855 12771 32861
rect 12176 32824 12204 32855
rect 12437 32827 12495 32833
rect 12176 32796 12388 32824
rect 12023 32728 12112 32756
rect 12023 32725 12035 32728
rect 11977 32719 12035 32725
rect 12250 32716 12256 32768
rect 12308 32716 12314 32768
rect 12360 32756 12388 32796
rect 12437 32793 12449 32827
rect 12483 32824 12495 32827
rect 12526 32824 12532 32836
rect 12483 32796 12532 32824
rect 12483 32793 12495 32796
rect 12437 32787 12495 32793
rect 12526 32784 12532 32796
rect 12584 32784 12590 32836
rect 12621 32827 12679 32833
rect 12621 32793 12633 32827
rect 12667 32824 12679 32827
rect 12802 32824 12808 32836
rect 12667 32796 12808 32824
rect 12667 32793 12679 32796
rect 12621 32787 12679 32793
rect 12802 32784 12808 32796
rect 12860 32784 12866 32836
rect 12897 32827 12955 32833
rect 12897 32793 12909 32827
rect 12943 32824 12955 32827
rect 12986 32824 12992 32836
rect 12943 32796 12992 32824
rect 12943 32793 12955 32796
rect 12897 32787 12955 32793
rect 12912 32756 12940 32787
rect 12986 32784 12992 32796
rect 13044 32784 13050 32836
rect 13081 32827 13139 32833
rect 13081 32793 13093 32827
rect 13127 32824 13139 32827
rect 13127 32796 13308 32824
rect 13127 32793 13139 32796
rect 13081 32787 13139 32793
rect 12360 32728 12940 32756
rect 13170 32716 13176 32768
rect 13228 32716 13234 32768
rect 13280 32756 13308 32796
rect 13354 32784 13360 32836
rect 13412 32784 13418 32836
rect 13446 32784 13452 32836
rect 13504 32824 13510 32836
rect 13541 32827 13599 32833
rect 13541 32824 13553 32827
rect 13504 32796 13553 32824
rect 13504 32784 13510 32796
rect 13541 32793 13553 32796
rect 13587 32793 13599 32827
rect 13832 32824 13860 32864
rect 13906 32852 13912 32904
rect 13964 32852 13970 32904
rect 14918 32892 14924 32904
rect 14016 32864 14924 32892
rect 14016 32824 14044 32864
rect 14918 32852 14924 32864
rect 14976 32852 14982 32904
rect 15013 32895 15071 32901
rect 15013 32861 15025 32895
rect 15059 32892 15071 32895
rect 15286 32892 15292 32904
rect 15059 32864 15292 32892
rect 15059 32861 15071 32864
rect 15013 32855 15071 32861
rect 15286 32852 15292 32864
rect 15344 32852 15350 32904
rect 15378 32852 15384 32904
rect 15436 32892 15442 32904
rect 15580 32901 15608 33000
rect 15565 32895 15623 32901
rect 15565 32892 15577 32895
rect 15436 32864 15577 32892
rect 15436 32852 15442 32864
rect 15565 32861 15577 32864
rect 15611 32861 15623 32895
rect 15565 32855 15623 32861
rect 15933 32895 15991 32901
rect 15933 32861 15945 32895
rect 15979 32892 15991 32895
rect 16114 32892 16120 32904
rect 15979 32864 16120 32892
rect 15979 32861 15991 32864
rect 15933 32855 15991 32861
rect 16114 32852 16120 32864
rect 16172 32852 16178 32904
rect 13832 32796 14044 32824
rect 14093 32827 14151 32833
rect 13541 32787 13599 32793
rect 14093 32793 14105 32827
rect 14139 32824 14151 32827
rect 14182 32824 14188 32836
rect 14139 32796 14188 32824
rect 14139 32793 14151 32796
rect 14093 32787 14151 32793
rect 14108 32756 14136 32787
rect 14182 32784 14188 32796
rect 14240 32784 14246 32836
rect 14274 32784 14280 32836
rect 14332 32784 14338 32836
rect 14366 32784 14372 32836
rect 14424 32824 14430 32836
rect 14553 32827 14611 32833
rect 14553 32824 14565 32827
rect 14424 32796 14565 32824
rect 14424 32784 14430 32796
rect 14553 32793 14565 32796
rect 14599 32793 14611 32827
rect 14553 32787 14611 32793
rect 14642 32784 14648 32836
rect 14700 32824 14706 32836
rect 14737 32827 14795 32833
rect 14737 32824 14749 32827
rect 14700 32796 14749 32824
rect 14700 32784 14706 32796
rect 14737 32793 14749 32796
rect 14783 32793 14795 32827
rect 14737 32787 14795 32793
rect 15197 32827 15255 32833
rect 15197 32793 15209 32827
rect 15243 32824 15255 32827
rect 15654 32824 15660 32836
rect 15243 32796 15660 32824
rect 15243 32793 15255 32796
rect 15197 32787 15255 32793
rect 15654 32784 15660 32796
rect 15712 32784 15718 32836
rect 15746 32784 15752 32836
rect 15804 32784 15810 32836
rect 15838 32784 15844 32836
rect 15896 32824 15902 32836
rect 16206 32824 16212 32836
rect 15896 32796 16212 32824
rect 15896 32784 15902 32796
rect 16206 32784 16212 32796
rect 16264 32784 16270 32836
rect 13280 32728 14136 32756
rect 14458 32716 14464 32768
rect 14516 32716 14522 32768
rect 14826 32716 14832 32768
rect 14884 32756 14890 32768
rect 14921 32759 14979 32765
rect 14921 32756 14933 32759
rect 14884 32728 14933 32756
rect 14884 32716 14890 32728
rect 14921 32725 14933 32728
rect 14967 32725 14979 32759
rect 14921 32719 14979 32725
rect 15286 32716 15292 32768
rect 15344 32756 15350 32768
rect 15381 32759 15439 32765
rect 15381 32756 15393 32759
rect 15344 32728 15393 32756
rect 15344 32716 15350 32728
rect 15381 32725 15393 32728
rect 15427 32725 15439 32759
rect 15381 32719 15439 32725
rect 15470 32716 15476 32768
rect 15528 32756 15534 32768
rect 16117 32759 16175 32765
rect 16117 32756 16129 32759
rect 15528 32728 16129 32756
rect 15528 32716 15534 32728
rect 16117 32725 16129 32728
rect 16163 32725 16175 32759
rect 16117 32719 16175 32725
rect 1104 32666 16652 32688
rect 1104 32614 4874 32666
rect 4926 32614 4938 32666
rect 4990 32614 5002 32666
rect 5054 32614 5066 32666
rect 5118 32614 5130 32666
rect 5182 32614 16652 32666
rect 1104 32592 16652 32614
rect 11330 32512 11336 32564
rect 11388 32552 11394 32564
rect 12437 32555 12495 32561
rect 12437 32552 12449 32555
rect 11388 32524 12449 32552
rect 11388 32512 11394 32524
rect 12437 32521 12449 32524
rect 12483 32552 12495 32555
rect 13354 32552 13360 32564
rect 12483 32524 13360 32552
rect 12483 32521 12495 32524
rect 12437 32515 12495 32521
rect 13354 32512 13360 32524
rect 13412 32512 13418 32564
rect 13446 32512 13452 32564
rect 13504 32552 13510 32564
rect 14366 32552 14372 32564
rect 13504 32524 14372 32552
rect 13504 32512 13510 32524
rect 14366 32512 14372 32524
rect 14424 32512 14430 32564
rect 14458 32512 14464 32564
rect 14516 32512 14522 32564
rect 14752 32524 15516 32552
rect 10778 32444 10784 32496
rect 10836 32444 10842 32496
rect 13998 32444 14004 32496
rect 14056 32484 14062 32496
rect 14476 32484 14504 32512
rect 14056 32456 14412 32484
rect 14476 32456 14596 32484
rect 14056 32444 14062 32456
rect 6917 32419 6975 32425
rect 6917 32385 6929 32419
rect 6963 32385 6975 32419
rect 6917 32379 6975 32385
rect 6932 32348 6960 32379
rect 7190 32376 7196 32428
rect 7248 32376 7254 32428
rect 7374 32376 7380 32428
rect 7432 32376 7438 32428
rect 7466 32376 7472 32428
rect 7524 32416 7530 32428
rect 8941 32419 8999 32425
rect 8941 32416 8953 32419
rect 7524 32388 8953 32416
rect 7524 32376 7530 32388
rect 8941 32385 8953 32388
rect 8987 32385 8999 32419
rect 8941 32379 8999 32385
rect 9122 32376 9128 32428
rect 9180 32376 9186 32428
rect 10597 32419 10655 32425
rect 10597 32385 10609 32419
rect 10643 32416 10655 32419
rect 10796 32416 10824 32444
rect 10643 32388 12848 32416
rect 10643 32385 10655 32388
rect 10597 32379 10655 32385
rect 7650 32348 7656 32360
rect 6932 32320 7656 32348
rect 7650 32308 7656 32320
rect 7708 32308 7714 32360
rect 10778 32308 10784 32360
rect 10836 32308 10842 32360
rect 10980 32320 12020 32348
rect 7006 32240 7012 32292
rect 7064 32240 7070 32292
rect 7098 32240 7104 32292
rect 7156 32240 7162 32292
rect 10413 32283 10471 32289
rect 10413 32249 10425 32283
rect 10459 32280 10471 32283
rect 10980 32280 11008 32320
rect 10459 32252 11008 32280
rect 10459 32249 10471 32252
rect 10413 32243 10471 32249
rect 11054 32240 11060 32292
rect 11112 32280 11118 32292
rect 11517 32283 11575 32289
rect 11517 32280 11529 32283
rect 11112 32252 11529 32280
rect 11112 32240 11118 32252
rect 11517 32249 11529 32252
rect 11563 32249 11575 32283
rect 11992 32280 12020 32320
rect 12066 32308 12072 32360
rect 12124 32308 12130 32360
rect 12618 32280 12624 32292
rect 11992 32252 12624 32280
rect 11517 32243 11575 32249
rect 12618 32240 12624 32252
rect 12676 32240 12682 32292
rect 6730 32172 6736 32224
rect 6788 32172 6794 32224
rect 8386 32172 8392 32224
rect 8444 32212 8450 32224
rect 9033 32215 9091 32221
rect 9033 32212 9045 32215
rect 8444 32184 9045 32212
rect 8444 32172 8450 32184
rect 9033 32181 9045 32184
rect 9079 32181 9091 32215
rect 9033 32175 9091 32181
rect 11330 32172 11336 32224
rect 11388 32172 11394 32224
rect 12820 32212 12848 32388
rect 13538 32376 13544 32428
rect 13596 32425 13602 32428
rect 13596 32379 13608 32425
rect 13596 32376 13602 32379
rect 13722 32376 13728 32428
rect 13780 32416 13786 32428
rect 14384 32425 14412 32456
rect 14369 32419 14427 32425
rect 13780 32388 14044 32416
rect 13780 32376 13786 32388
rect 13817 32351 13875 32357
rect 13817 32317 13829 32351
rect 13863 32348 13875 32351
rect 13906 32348 13912 32360
rect 13863 32320 13912 32348
rect 13863 32317 13875 32320
rect 13817 32311 13875 32317
rect 13906 32308 13912 32320
rect 13964 32308 13970 32360
rect 14016 32348 14044 32388
rect 14369 32385 14381 32419
rect 14415 32385 14427 32419
rect 14369 32379 14427 32385
rect 14458 32376 14464 32428
rect 14516 32376 14522 32428
rect 14568 32425 14596 32456
rect 14752 32425 14780 32524
rect 14918 32444 14924 32496
rect 14976 32484 14982 32496
rect 14976 32456 15332 32484
rect 14976 32444 14982 32456
rect 14553 32419 14611 32425
rect 14553 32385 14565 32419
rect 14599 32385 14611 32419
rect 14553 32379 14611 32385
rect 14737 32419 14795 32425
rect 14737 32385 14749 32419
rect 14783 32385 14795 32419
rect 14737 32379 14795 32385
rect 14642 32348 14648 32360
rect 14016 32320 14648 32348
rect 14642 32308 14648 32320
rect 14700 32308 14706 32360
rect 14752 32348 14780 32379
rect 15010 32376 15016 32428
rect 15068 32416 15074 32428
rect 15304 32425 15332 32456
rect 15488 32425 15516 32524
rect 15654 32444 15660 32496
rect 15712 32484 15718 32496
rect 15841 32487 15899 32493
rect 15841 32484 15853 32487
rect 15712 32456 15853 32484
rect 15712 32444 15718 32456
rect 15841 32453 15853 32456
rect 15887 32453 15899 32487
rect 15841 32447 15899 32453
rect 15105 32419 15163 32425
rect 15105 32416 15117 32419
rect 15068 32388 15117 32416
rect 15068 32376 15074 32388
rect 15105 32385 15117 32388
rect 15151 32385 15163 32419
rect 15105 32379 15163 32385
rect 15197 32419 15255 32425
rect 15197 32385 15209 32419
rect 15243 32385 15255 32419
rect 15197 32379 15255 32385
rect 15289 32419 15347 32425
rect 15289 32385 15301 32419
rect 15335 32385 15347 32419
rect 15289 32379 15347 32385
rect 15473 32419 15531 32425
rect 15473 32385 15485 32419
rect 15519 32385 15531 32419
rect 15749 32419 15807 32425
rect 15749 32416 15761 32419
rect 15473 32379 15531 32385
rect 15672 32388 15761 32416
rect 14826 32348 14832 32360
rect 14752 32320 14832 32348
rect 14752 32280 14780 32320
rect 14826 32308 14832 32320
rect 14884 32308 14890 32360
rect 14016 32252 14780 32280
rect 14016 32212 14044 32252
rect 15102 32240 15108 32292
rect 15160 32280 15166 32292
rect 15212 32280 15240 32379
rect 15672 32360 15700 32388
rect 15749 32385 15761 32388
rect 15795 32385 15807 32419
rect 15749 32379 15807 32385
rect 15856 32360 15884 32447
rect 15930 32376 15936 32428
rect 15988 32376 15994 32428
rect 16117 32419 16175 32425
rect 16117 32385 16129 32419
rect 16163 32385 16175 32419
rect 16117 32379 16175 32385
rect 15654 32308 15660 32360
rect 15712 32308 15718 32360
rect 15838 32308 15844 32360
rect 15896 32308 15902 32360
rect 16132 32280 16160 32379
rect 15160 32252 15240 32280
rect 15304 32252 16160 32280
rect 15160 32240 15166 32252
rect 12820 32184 14044 32212
rect 14090 32172 14096 32224
rect 14148 32172 14154 32224
rect 14366 32172 14372 32224
rect 14424 32212 14430 32224
rect 14829 32215 14887 32221
rect 14829 32212 14841 32215
rect 14424 32184 14841 32212
rect 14424 32172 14430 32184
rect 14829 32181 14841 32184
rect 14875 32181 14887 32215
rect 14829 32175 14887 32181
rect 14918 32172 14924 32224
rect 14976 32212 14982 32224
rect 15304 32212 15332 32252
rect 14976 32184 15332 32212
rect 14976 32172 14982 32184
rect 15562 32172 15568 32224
rect 15620 32172 15626 32224
rect 1104 32122 16652 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 16652 32122
rect 1104 32048 16652 32070
rect 7837 32011 7895 32017
rect 7837 31977 7849 32011
rect 7883 32008 7895 32011
rect 8110 32008 8116 32020
rect 7883 31980 8116 32008
rect 7883 31977 7895 31980
rect 7837 31971 7895 31977
rect 8110 31968 8116 31980
rect 8168 31968 8174 32020
rect 8941 32011 8999 32017
rect 8941 31977 8953 32011
rect 8987 32008 8999 32011
rect 9122 32008 9128 32020
rect 8987 31980 9128 32008
rect 8987 31977 8999 31980
rect 8941 31971 8999 31977
rect 8386 31832 8392 31884
rect 8444 31832 8450 31884
rect 6457 31807 6515 31813
rect 6457 31773 6469 31807
rect 6503 31804 6515 31807
rect 6503 31776 6914 31804
rect 6503 31773 6515 31776
rect 6457 31767 6515 31773
rect 6886 31748 6914 31776
rect 8110 31764 8116 31816
rect 8168 31764 8174 31816
rect 8478 31764 8484 31816
rect 8536 31804 8542 31816
rect 8573 31807 8631 31813
rect 8573 31804 8585 31807
rect 8536 31776 8585 31804
rect 8536 31764 8542 31776
rect 8573 31773 8585 31776
rect 8619 31773 8631 31807
rect 8573 31767 8631 31773
rect 8665 31807 8723 31813
rect 8665 31773 8677 31807
rect 8711 31804 8723 31807
rect 8956 31804 8984 31971
rect 9122 31968 9128 31980
rect 9180 31968 9186 32020
rect 11514 31968 11520 32020
rect 11572 32008 11578 32020
rect 12161 32011 12219 32017
rect 12161 32008 12173 32011
rect 11572 31980 12173 32008
rect 11572 31968 11578 31980
rect 12161 31977 12173 31980
rect 12207 32008 12219 32011
rect 13722 32008 13728 32020
rect 12207 31980 13728 32008
rect 12207 31977 12219 31980
rect 12161 31971 12219 31977
rect 13722 31968 13728 31980
rect 13780 31968 13786 32020
rect 13814 31968 13820 32020
rect 13872 31968 13878 32020
rect 15378 31968 15384 32020
rect 15436 32008 15442 32020
rect 15473 32011 15531 32017
rect 15473 32008 15485 32011
rect 15436 31980 15485 32008
rect 15436 31968 15442 31980
rect 15473 31977 15485 31980
rect 15519 31977 15531 32011
rect 15473 31971 15531 31977
rect 10778 31900 10784 31952
rect 10836 31940 10842 31952
rect 10962 31940 10968 31952
rect 10836 31912 10968 31940
rect 10836 31900 10842 31912
rect 10962 31900 10968 31912
rect 11020 31940 11026 31952
rect 11057 31943 11115 31949
rect 11057 31940 11069 31943
rect 11020 31912 11069 31940
rect 11020 31900 11026 31912
rect 11057 31909 11069 31912
rect 11103 31909 11115 31943
rect 11057 31903 11115 31909
rect 11149 31943 11207 31949
rect 11149 31909 11161 31943
rect 11195 31909 11207 31943
rect 11149 31903 11207 31909
rect 8711 31776 8984 31804
rect 8711 31773 8723 31776
rect 8665 31767 8723 31773
rect 9398 31764 9404 31816
rect 9456 31804 9462 31816
rect 9493 31807 9551 31813
rect 9493 31804 9505 31807
rect 9456 31776 9505 31804
rect 9456 31764 9462 31776
rect 9493 31773 9505 31776
rect 9539 31773 9551 31807
rect 9493 31767 9551 31773
rect 9674 31764 9680 31816
rect 9732 31764 9738 31816
rect 9944 31807 10002 31813
rect 9944 31773 9956 31807
rect 9990 31804 10002 31807
rect 11164 31804 11192 31903
rect 16022 31900 16028 31952
rect 16080 31940 16086 31952
rect 16209 31943 16267 31949
rect 16209 31940 16221 31943
rect 16080 31912 16221 31940
rect 16080 31900 16086 31912
rect 16209 31909 16221 31912
rect 16255 31909 16267 31943
rect 16209 31903 16267 31909
rect 11330 31832 11336 31884
rect 11388 31872 11394 31884
rect 11609 31875 11667 31881
rect 11609 31872 11621 31875
rect 11388 31844 11621 31872
rect 11388 31832 11394 31844
rect 11609 31841 11621 31844
rect 11655 31841 11667 31875
rect 11609 31835 11667 31841
rect 11701 31875 11759 31881
rect 11701 31841 11713 31875
rect 11747 31841 11759 31875
rect 15930 31872 15936 31884
rect 11701 31835 11759 31841
rect 13565 31844 13768 31872
rect 11716 31804 11744 31835
rect 13565 31813 13593 31844
rect 13740 31816 13768 31844
rect 15856 31844 15936 31872
rect 9990 31776 11192 31804
rect 11256 31776 11744 31804
rect 13541 31807 13599 31813
rect 9990 31773 10002 31776
rect 9944 31767 10002 31773
rect 6730 31745 6736 31748
rect 6724 31699 6736 31745
rect 6730 31696 6736 31699
rect 6788 31696 6794 31748
rect 6886 31708 6920 31748
rect 6914 31696 6920 31708
rect 6972 31696 6978 31748
rect 8297 31739 8355 31745
rect 8297 31705 8309 31739
rect 8343 31736 8355 31739
rect 8846 31736 8852 31748
rect 8343 31708 8852 31736
rect 8343 31705 8355 31708
rect 8297 31699 8355 31705
rect 8846 31696 8852 31708
rect 8904 31696 8910 31748
rect 10686 31696 10692 31748
rect 10744 31736 10750 31748
rect 11256 31736 11284 31776
rect 13541 31773 13553 31807
rect 13587 31773 13599 31807
rect 13541 31767 13599 31773
rect 13633 31807 13691 31813
rect 13633 31773 13645 31807
rect 13679 31773 13691 31807
rect 13633 31767 13691 31773
rect 10744 31708 11284 31736
rect 10744 31696 10750 31708
rect 13078 31696 13084 31748
rect 13136 31736 13142 31748
rect 13274 31739 13332 31745
rect 13274 31736 13286 31739
rect 13136 31708 13286 31736
rect 13136 31696 13142 31708
rect 13274 31705 13286 31708
rect 13320 31705 13332 31739
rect 13274 31699 13332 31705
rect 13648 31680 13676 31767
rect 13722 31764 13728 31816
rect 13780 31804 13786 31816
rect 13906 31804 13912 31816
rect 13780 31776 13912 31804
rect 13780 31764 13786 31776
rect 13906 31764 13912 31776
rect 13964 31804 13970 31816
rect 14093 31807 14151 31813
rect 14093 31804 14105 31807
rect 13964 31776 14105 31804
rect 13964 31764 13970 31776
rect 14093 31773 14105 31776
rect 14139 31804 14151 31807
rect 14918 31804 14924 31816
rect 14139 31776 14924 31804
rect 14139 31773 14151 31776
rect 14093 31767 14151 31773
rect 14918 31764 14924 31776
rect 14976 31764 14982 31816
rect 15102 31804 15108 31816
rect 15028 31776 15108 31804
rect 14366 31745 14372 31748
rect 14360 31699 14372 31745
rect 14366 31696 14372 31699
rect 14424 31696 14430 31748
rect 14458 31696 14464 31748
rect 14516 31736 14522 31748
rect 15028 31736 15056 31776
rect 15102 31764 15108 31776
rect 15160 31764 15166 31816
rect 15194 31764 15200 31816
rect 15252 31804 15258 31816
rect 15856 31813 15884 31844
rect 15930 31832 15936 31844
rect 15988 31872 15994 31884
rect 16390 31872 16396 31884
rect 15988 31844 16396 31872
rect 15988 31832 15994 31844
rect 16390 31832 16396 31844
rect 16448 31832 16454 31884
rect 15657 31807 15715 31813
rect 15657 31804 15669 31807
rect 15252 31776 15669 31804
rect 15252 31764 15258 31776
rect 15657 31773 15669 31776
rect 15703 31773 15715 31807
rect 15657 31767 15715 31773
rect 15841 31807 15899 31813
rect 15841 31773 15853 31807
rect 15887 31773 15899 31807
rect 15841 31767 15899 31773
rect 16025 31807 16083 31813
rect 16025 31773 16037 31807
rect 16071 31804 16083 31807
rect 16114 31804 16120 31816
rect 16071 31776 16120 31804
rect 16071 31773 16083 31776
rect 16025 31767 16083 31773
rect 16114 31764 16120 31776
rect 16172 31764 16178 31816
rect 14516 31708 15056 31736
rect 15933 31739 15991 31745
rect 14516 31696 14522 31708
rect 15933 31705 15945 31739
rect 15979 31705 15991 31739
rect 15933 31699 15991 31705
rect 7926 31628 7932 31680
rect 7984 31628 7990 31680
rect 8389 31671 8447 31677
rect 8389 31637 8401 31671
rect 8435 31668 8447 31671
rect 8478 31668 8484 31680
rect 8435 31640 8484 31668
rect 8435 31637 8447 31640
rect 8389 31631 8447 31637
rect 8478 31628 8484 31640
rect 8536 31628 8542 31680
rect 11514 31628 11520 31680
rect 11572 31628 11578 31680
rect 13630 31628 13636 31680
rect 13688 31628 13694 31680
rect 15948 31668 15976 31699
rect 16114 31668 16120 31680
rect 15948 31640 16120 31668
rect 16114 31628 16120 31640
rect 16172 31628 16178 31680
rect 1104 31578 16652 31600
rect 1104 31526 4874 31578
rect 4926 31526 4938 31578
rect 4990 31526 5002 31578
rect 5054 31526 5066 31578
rect 5118 31526 5130 31578
rect 5182 31526 16652 31578
rect 1104 31504 16652 31526
rect 7374 31424 7380 31476
rect 7432 31464 7438 31476
rect 7469 31467 7527 31473
rect 7469 31464 7481 31467
rect 7432 31436 7481 31464
rect 7432 31424 7438 31436
rect 7469 31433 7481 31436
rect 7515 31433 7527 31467
rect 7469 31427 7527 31433
rect 11057 31467 11115 31473
rect 11057 31433 11069 31467
rect 11103 31464 11115 31467
rect 11238 31464 11244 31476
rect 11103 31436 11244 31464
rect 11103 31433 11115 31436
rect 11057 31427 11115 31433
rect 11238 31424 11244 31436
rect 11296 31464 11302 31476
rect 12066 31464 12072 31476
rect 11296 31436 12072 31464
rect 11296 31424 11302 31436
rect 12066 31424 12072 31436
rect 12124 31424 12130 31476
rect 14274 31424 14280 31476
rect 14332 31464 14338 31476
rect 14921 31467 14979 31473
rect 14921 31464 14933 31467
rect 14332 31436 14933 31464
rect 14332 31424 14338 31436
rect 14921 31433 14933 31436
rect 14967 31433 14979 31467
rect 14921 31427 14979 31433
rect 7926 31356 7932 31408
rect 7984 31396 7990 31408
rect 8113 31399 8171 31405
rect 8113 31396 8125 31399
rect 7984 31368 8125 31396
rect 7984 31356 7990 31368
rect 8113 31365 8125 31368
rect 8159 31365 8171 31399
rect 13722 31396 13728 31408
rect 8113 31359 8171 31365
rect 12912 31368 13728 31396
rect 7098 31288 7104 31340
rect 7156 31328 7162 31340
rect 7558 31328 7564 31340
rect 7156 31300 7564 31328
rect 7156 31288 7162 31300
rect 7558 31288 7564 31300
rect 7616 31328 7622 31340
rect 8478 31337 8484 31340
rect 7745 31331 7803 31337
rect 7745 31328 7757 31331
rect 7616 31300 7757 31328
rect 7616 31288 7622 31300
rect 7745 31297 7757 31300
rect 7791 31297 7803 31331
rect 8472 31328 8484 31337
rect 8439 31300 8484 31328
rect 7745 31291 7803 31297
rect 8472 31291 8484 31300
rect 8478 31288 8484 31291
rect 8536 31288 8542 31340
rect 9674 31288 9680 31340
rect 9732 31288 9738 31340
rect 9950 31337 9956 31340
rect 9944 31291 9956 31337
rect 9950 31288 9956 31291
rect 10008 31288 10014 31340
rect 12342 31288 12348 31340
rect 12400 31328 12406 31340
rect 12912 31337 12940 31368
rect 12630 31331 12688 31337
rect 12630 31328 12642 31331
rect 12400 31300 12642 31328
rect 12400 31288 12406 31300
rect 12630 31297 12642 31300
rect 12676 31297 12688 31331
rect 12630 31291 12688 31297
rect 12897 31331 12955 31337
rect 12897 31297 12909 31331
rect 12943 31297 12955 31331
rect 12897 31291 12955 31297
rect 12986 31288 12992 31340
rect 13044 31288 13050 31340
rect 13556 31337 13584 31368
rect 13722 31356 13728 31368
rect 13780 31356 13786 31408
rect 14182 31356 14188 31408
rect 14240 31396 14246 31408
rect 15013 31399 15071 31405
rect 15013 31396 15025 31399
rect 14240 31368 15025 31396
rect 14240 31356 14246 31368
rect 15013 31365 15025 31368
rect 15059 31365 15071 31399
rect 15013 31359 15071 31365
rect 13357 31331 13415 31337
rect 13357 31297 13369 31331
rect 13403 31297 13415 31331
rect 13357 31291 13415 31297
rect 13541 31331 13599 31337
rect 13541 31297 13553 31331
rect 13587 31297 13599 31331
rect 13541 31291 13599 31297
rect 6086 31220 6092 31272
rect 6144 31260 6150 31272
rect 7285 31263 7343 31269
rect 7285 31260 7297 31263
rect 6144 31232 7297 31260
rect 6144 31220 6150 31232
rect 7285 31229 7297 31232
rect 7331 31229 7343 31263
rect 7285 31223 7343 31229
rect 7650 31220 7656 31272
rect 7708 31220 7714 31272
rect 8018 31220 8024 31272
rect 8076 31220 8082 31272
rect 8205 31263 8263 31269
rect 8205 31229 8217 31263
rect 8251 31229 8263 31263
rect 13372 31260 13400 31291
rect 13630 31288 13636 31340
rect 13688 31288 13694 31340
rect 13808 31331 13866 31337
rect 13808 31297 13820 31331
rect 13854 31328 13866 31331
rect 14090 31328 14096 31340
rect 13854 31300 14096 31328
rect 13854 31297 13866 31300
rect 13808 31291 13866 31297
rect 14090 31288 14096 31300
rect 14148 31288 14154 31340
rect 15194 31288 15200 31340
rect 15252 31288 15258 31340
rect 16298 31288 16304 31340
rect 16356 31288 16362 31340
rect 13648 31260 13676 31288
rect 13372 31232 13676 31260
rect 8205 31223 8263 31229
rect 6914 31152 6920 31204
rect 6972 31192 6978 31204
rect 8220 31192 8248 31223
rect 15378 31220 15384 31272
rect 15436 31260 15442 31272
rect 16025 31263 16083 31269
rect 16025 31260 16037 31263
rect 15436 31232 16037 31260
rect 15436 31220 15442 31232
rect 16025 31229 16037 31232
rect 16071 31229 16083 31263
rect 16025 31223 16083 31229
rect 15838 31192 15844 31204
rect 6972 31164 8248 31192
rect 13004 31164 13584 31192
rect 6972 31152 6978 31164
rect 6730 31084 6736 31136
rect 6788 31084 6794 31136
rect 9398 31084 9404 31136
rect 9456 31124 9462 31136
rect 9585 31127 9643 31133
rect 9585 31124 9597 31127
rect 9456 31096 9597 31124
rect 9456 31084 9462 31096
rect 9585 31093 9597 31096
rect 9631 31093 9643 31127
rect 9585 31087 9643 31093
rect 11517 31127 11575 31133
rect 11517 31093 11529 31127
rect 11563 31124 11575 31127
rect 11882 31124 11888 31136
rect 11563 31096 11888 31124
rect 11563 31093 11575 31096
rect 11517 31087 11575 31093
rect 11882 31084 11888 31096
rect 11940 31084 11946 31136
rect 11974 31084 11980 31136
rect 12032 31124 12038 31136
rect 13004 31124 13032 31164
rect 12032 31096 13032 31124
rect 13556 31124 13584 31164
rect 15304 31164 15844 31192
rect 15304 31124 15332 31164
rect 15838 31152 15844 31164
rect 15896 31192 15902 31204
rect 16298 31192 16304 31204
rect 15896 31164 16304 31192
rect 15896 31152 15902 31164
rect 16298 31152 16304 31164
rect 16356 31152 16362 31204
rect 13556 31096 15332 31124
rect 15381 31127 15439 31133
rect 12032 31084 12038 31096
rect 15381 31093 15393 31127
rect 15427 31124 15439 31127
rect 15746 31124 15752 31136
rect 15427 31096 15752 31124
rect 15427 31093 15439 31096
rect 15381 31087 15439 31093
rect 15746 31084 15752 31096
rect 15804 31084 15810 31136
rect 1104 31034 16652 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 16652 31034
rect 1104 30960 16652 30982
rect 6086 30880 6092 30932
rect 6144 30880 6150 30932
rect 8018 30880 8024 30932
rect 8076 30920 8082 30932
rect 8941 30923 8999 30929
rect 8941 30920 8953 30923
rect 8076 30892 8953 30920
rect 8076 30880 8082 30892
rect 8941 30889 8953 30892
rect 8987 30889 8999 30923
rect 8941 30883 8999 30889
rect 9858 30880 9864 30932
rect 9916 30880 9922 30932
rect 9950 30880 9956 30932
rect 10008 30920 10014 30932
rect 10137 30923 10195 30929
rect 10137 30920 10149 30923
rect 10008 30892 10149 30920
rect 10008 30880 10014 30892
rect 10137 30889 10149 30892
rect 10183 30889 10195 30923
rect 10137 30883 10195 30889
rect 11882 30880 11888 30932
rect 11940 30920 11946 30932
rect 11940 30892 13860 30920
rect 11940 30880 11946 30892
rect 8478 30852 8484 30864
rect 7760 30824 8484 30852
rect 6454 30676 6460 30728
rect 6512 30716 6518 30728
rect 6914 30716 6920 30728
rect 6512 30688 6920 30716
rect 6512 30676 6518 30688
rect 6914 30676 6920 30688
rect 6972 30716 6978 30728
rect 7466 30716 7472 30728
rect 6972 30688 7472 30716
rect 6972 30676 6978 30688
rect 7466 30676 7472 30688
rect 7524 30676 7530 30728
rect 7760 30725 7788 30824
rect 8478 30812 8484 30824
rect 8536 30812 8542 30864
rect 9674 30812 9680 30864
rect 9732 30852 9738 30864
rect 12437 30855 12495 30861
rect 9732 30824 11008 30852
rect 9732 30812 9738 30824
rect 8297 30787 8355 30793
rect 8297 30753 8309 30787
rect 8343 30784 8355 30787
rect 8343 30756 9260 30784
rect 8343 30753 8355 30756
rect 8297 30747 8355 30753
rect 9232 30728 9260 30756
rect 9950 30744 9956 30796
rect 10008 30744 10014 30796
rect 10226 30744 10232 30796
rect 10284 30784 10290 30796
rect 10686 30784 10692 30796
rect 10284 30756 10692 30784
rect 10284 30744 10290 30756
rect 10686 30744 10692 30756
rect 10744 30744 10750 30796
rect 10980 30793 11008 30824
rect 12437 30821 12449 30855
rect 12483 30821 12495 30855
rect 12437 30815 12495 30821
rect 10965 30787 11023 30793
rect 10965 30753 10977 30787
rect 11011 30753 11023 30787
rect 10965 30747 11023 30753
rect 7653 30719 7711 30725
rect 7653 30685 7665 30719
rect 7699 30685 7711 30719
rect 7653 30679 7711 30685
rect 7745 30719 7803 30725
rect 7745 30685 7757 30719
rect 7791 30685 7803 30719
rect 7745 30679 7803 30685
rect 7929 30719 7987 30725
rect 7929 30685 7941 30719
rect 7975 30716 7987 30719
rect 8205 30719 8263 30725
rect 8205 30716 8217 30719
rect 7975 30688 8217 30716
rect 7975 30685 7987 30688
rect 7929 30679 7987 30685
rect 8205 30685 8217 30688
rect 8251 30685 8263 30719
rect 8205 30679 8263 30685
rect 7006 30608 7012 30660
rect 7064 30648 7070 30660
rect 7202 30651 7260 30657
rect 7202 30648 7214 30651
rect 7064 30620 7214 30648
rect 7064 30608 7070 30620
rect 7202 30617 7214 30620
rect 7248 30617 7260 30651
rect 7668 30648 7696 30679
rect 8386 30676 8392 30728
rect 8444 30676 8450 30728
rect 8478 30676 8484 30728
rect 8536 30676 8542 30728
rect 8665 30719 8723 30725
rect 8665 30685 8677 30719
rect 8711 30716 8723 30719
rect 8846 30716 8852 30728
rect 8711 30688 8852 30716
rect 8711 30685 8723 30688
rect 8665 30679 8723 30685
rect 8846 30676 8852 30688
rect 8904 30676 8910 30728
rect 9122 30676 9128 30728
rect 9180 30676 9186 30728
rect 9214 30676 9220 30728
rect 9272 30676 9278 30728
rect 9401 30719 9459 30725
rect 9401 30685 9413 30719
rect 9447 30685 9459 30719
rect 9401 30679 9459 30685
rect 8404 30648 8432 30676
rect 9416 30648 9444 30679
rect 9490 30676 9496 30728
rect 9548 30676 9554 30728
rect 9769 30719 9827 30725
rect 9769 30685 9781 30719
rect 9815 30716 9827 30719
rect 10134 30716 10140 30728
rect 9815 30688 10140 30716
rect 9815 30685 9827 30688
rect 9769 30679 9827 30685
rect 10134 30676 10140 30688
rect 10192 30676 10198 30728
rect 10505 30719 10563 30725
rect 10505 30685 10517 30719
rect 10551 30716 10563 30719
rect 12452 30716 12480 30815
rect 12710 30744 12716 30796
rect 12768 30784 12774 30796
rect 13832 30793 13860 30892
rect 16298 30880 16304 30932
rect 16356 30880 16362 30932
rect 14550 30812 14556 30864
rect 14608 30812 14614 30864
rect 12989 30787 13047 30793
rect 12989 30784 13001 30787
rect 12768 30756 13001 30784
rect 12768 30744 12774 30756
rect 12989 30753 13001 30756
rect 13035 30753 13047 30787
rect 12989 30747 13047 30753
rect 13817 30787 13875 30793
rect 13817 30753 13829 30787
rect 13863 30753 13875 30787
rect 14568 30784 14596 30812
rect 13817 30747 13875 30753
rect 13924 30756 14780 30784
rect 10551 30688 12480 30716
rect 10551 30685 10563 30688
rect 10505 30679 10563 30685
rect 12618 30676 12624 30728
rect 12676 30716 12682 30728
rect 13924 30716 13952 30756
rect 12676 30688 13952 30716
rect 12676 30676 12682 30688
rect 13998 30676 14004 30728
rect 14056 30716 14062 30728
rect 14366 30716 14372 30728
rect 14056 30688 14372 30716
rect 14056 30676 14062 30688
rect 14366 30676 14372 30688
rect 14424 30676 14430 30728
rect 14461 30719 14519 30725
rect 14461 30685 14473 30719
rect 14507 30685 14519 30719
rect 14461 30679 14519 30685
rect 14553 30719 14611 30725
rect 14553 30685 14565 30719
rect 14599 30716 14611 30719
rect 14642 30716 14648 30728
rect 14599 30688 14648 30716
rect 14599 30685 14611 30688
rect 14553 30679 14611 30685
rect 7668 30620 8340 30648
rect 8404 30620 9444 30648
rect 10045 30651 10103 30657
rect 7202 30611 7260 30617
rect 8018 30540 8024 30592
rect 8076 30540 8082 30592
rect 8312 30580 8340 30620
rect 10045 30617 10057 30651
rect 10091 30648 10103 30651
rect 10410 30648 10416 30660
rect 10091 30620 10416 30648
rect 10091 30617 10103 30620
rect 10045 30611 10103 30617
rect 10410 30608 10416 30620
rect 10468 30608 10474 30660
rect 10597 30651 10655 30657
rect 10597 30617 10609 30651
rect 10643 30648 10655 30651
rect 11054 30648 11060 30660
rect 10643 30620 11060 30648
rect 10643 30617 10655 30620
rect 10597 30611 10655 30617
rect 11054 30608 11060 30620
rect 11112 30608 11118 30660
rect 11232 30651 11290 30657
rect 11232 30617 11244 30651
rect 11278 30648 11290 30651
rect 11790 30648 11796 30660
rect 11278 30620 11796 30648
rect 11278 30617 11290 30620
rect 11232 30611 11290 30617
rect 11790 30608 11796 30620
rect 11848 30608 11854 30660
rect 12802 30648 12808 30660
rect 12360 30620 12808 30648
rect 9398 30580 9404 30592
rect 8312 30552 9404 30580
rect 9398 30540 9404 30552
rect 9456 30540 9462 30592
rect 9585 30583 9643 30589
rect 9585 30549 9597 30583
rect 9631 30580 9643 30583
rect 9766 30580 9772 30592
rect 9631 30552 9772 30580
rect 9631 30549 9643 30552
rect 9585 30543 9643 30549
rect 9766 30540 9772 30552
rect 9824 30540 9830 30592
rect 12360 30589 12388 30620
rect 12802 30608 12808 30620
rect 12860 30608 12866 30660
rect 13078 30608 13084 30660
rect 13136 30648 13142 30660
rect 14093 30651 14151 30657
rect 14093 30648 14105 30651
rect 13136 30620 14105 30648
rect 13136 30608 13142 30620
rect 14093 30617 14105 30620
rect 14139 30617 14151 30651
rect 14093 30611 14151 30617
rect 14274 30608 14280 30660
rect 14332 30648 14338 30660
rect 14476 30648 14504 30679
rect 14642 30676 14648 30688
rect 14700 30676 14706 30728
rect 14752 30725 14780 30756
rect 14737 30719 14795 30725
rect 14737 30685 14749 30719
rect 14783 30685 14795 30719
rect 14737 30679 14795 30685
rect 14918 30676 14924 30728
rect 14976 30676 14982 30728
rect 14332 30620 14504 30648
rect 14332 30608 14338 30620
rect 14826 30608 14832 30660
rect 14884 30648 14890 30660
rect 15166 30651 15224 30657
rect 15166 30648 15178 30651
rect 14884 30620 15178 30648
rect 14884 30608 14890 30620
rect 15166 30617 15178 30620
rect 15212 30617 15224 30651
rect 15166 30611 15224 30617
rect 12345 30583 12403 30589
rect 12345 30549 12357 30583
rect 12391 30549 12403 30583
rect 12345 30543 12403 30549
rect 12434 30540 12440 30592
rect 12492 30580 12498 30592
rect 12897 30583 12955 30589
rect 12897 30580 12909 30583
rect 12492 30552 12909 30580
rect 12492 30540 12498 30552
rect 12897 30549 12909 30552
rect 12943 30549 12955 30583
rect 12897 30543 12955 30549
rect 13262 30540 13268 30592
rect 13320 30540 13326 30592
rect 1104 30490 16652 30512
rect 1104 30438 4874 30490
rect 4926 30438 4938 30490
rect 4990 30438 5002 30490
rect 5054 30438 5066 30490
rect 5118 30438 5130 30490
rect 5182 30438 16652 30490
rect 1104 30416 16652 30438
rect 6089 30379 6147 30385
rect 6089 30345 6101 30379
rect 6135 30376 6147 30379
rect 6730 30376 6736 30388
rect 6135 30348 6736 30376
rect 6135 30345 6147 30348
rect 6089 30339 6147 30345
rect 6730 30336 6736 30348
rect 6788 30336 6794 30388
rect 6822 30336 6828 30388
rect 6880 30336 6886 30388
rect 8478 30336 8484 30388
rect 8536 30376 8542 30388
rect 9309 30379 9367 30385
rect 9309 30376 9321 30379
rect 8536 30348 9321 30376
rect 8536 30336 8542 30348
rect 9309 30345 9321 30348
rect 9355 30376 9367 30379
rect 9582 30376 9588 30388
rect 9355 30348 9588 30376
rect 9355 30345 9367 30348
rect 9309 30339 9367 30345
rect 9582 30336 9588 30348
rect 9640 30336 9646 30388
rect 9858 30336 9864 30388
rect 9916 30376 9922 30388
rect 10870 30376 10876 30388
rect 9916 30348 10876 30376
rect 9916 30336 9922 30348
rect 10870 30336 10876 30348
rect 10928 30336 10934 30388
rect 11514 30336 11520 30388
rect 11572 30336 11578 30388
rect 11882 30336 11888 30388
rect 11940 30336 11946 30388
rect 12342 30336 12348 30388
rect 12400 30336 12406 30388
rect 12713 30379 12771 30385
rect 12713 30345 12725 30379
rect 12759 30376 12771 30379
rect 13262 30376 13268 30388
rect 12759 30348 13268 30376
rect 12759 30345 12771 30348
rect 12713 30339 12771 30345
rect 13262 30336 13268 30348
rect 13320 30336 13326 30388
rect 16206 30336 16212 30388
rect 16264 30376 16270 30388
rect 16301 30379 16359 30385
rect 16301 30376 16313 30379
rect 16264 30348 16313 30376
rect 16264 30336 16270 30348
rect 16301 30345 16313 30348
rect 16347 30345 16359 30379
rect 16301 30339 16359 30345
rect 6454 30308 6460 30320
rect 5460 30280 6316 30308
rect 5460 30249 5488 30280
rect 5445 30243 5503 30249
rect 5445 30209 5457 30243
rect 5491 30209 5503 30243
rect 5445 30203 5503 30209
rect 5629 30243 5687 30249
rect 5629 30209 5641 30243
rect 5675 30209 5687 30243
rect 5629 30203 5687 30209
rect 5644 30172 5672 30203
rect 5902 30200 5908 30252
rect 5960 30200 5966 30252
rect 6178 30200 6184 30252
rect 6236 30200 6242 30252
rect 6086 30172 6092 30184
rect 5644 30144 6092 30172
rect 6086 30132 6092 30144
rect 6144 30132 6150 30184
rect 6288 30172 6316 30280
rect 6380 30280 6460 30308
rect 6380 30249 6408 30280
rect 6454 30268 6460 30280
rect 6512 30268 6518 30320
rect 6632 30311 6690 30317
rect 6632 30277 6644 30311
rect 6678 30308 6690 30311
rect 6840 30308 6868 30336
rect 6678 30280 6868 30308
rect 6678 30277 6690 30280
rect 6632 30271 6690 30277
rect 8018 30268 8024 30320
rect 8076 30308 8082 30320
rect 8174 30311 8232 30317
rect 8174 30308 8186 30311
rect 8076 30280 8186 30308
rect 8076 30268 8082 30280
rect 8174 30277 8186 30280
rect 8220 30277 8232 30311
rect 8174 30271 8232 30277
rect 9401 30311 9459 30317
rect 9401 30277 9413 30311
rect 9447 30308 9459 30311
rect 10134 30308 10140 30320
rect 9447 30280 10140 30308
rect 9447 30277 9459 30280
rect 9401 30271 9459 30277
rect 10134 30268 10140 30280
rect 10192 30268 10198 30320
rect 10321 30311 10379 30317
rect 10321 30277 10333 30311
rect 10367 30308 10379 30311
rect 10778 30308 10784 30320
rect 10367 30280 10784 30308
rect 10367 30277 10379 30280
rect 10321 30271 10379 30277
rect 10778 30268 10784 30280
rect 10836 30268 10842 30320
rect 12802 30268 12808 30320
rect 12860 30308 12866 30320
rect 12860 30280 13032 30308
rect 12860 30268 12866 30280
rect 6365 30243 6423 30249
rect 6365 30209 6377 30243
rect 6411 30209 6423 30243
rect 6365 30203 6423 30209
rect 6472 30212 7420 30240
rect 6472 30172 6500 30212
rect 6288 30144 6500 30172
rect 7392 30172 7420 30212
rect 7466 30200 7472 30252
rect 7524 30240 7530 30252
rect 7926 30240 7932 30252
rect 7524 30212 7932 30240
rect 7524 30200 7530 30212
rect 7926 30200 7932 30212
rect 7984 30200 7990 30252
rect 9861 30243 9919 30249
rect 9861 30209 9873 30243
rect 9907 30240 9919 30243
rect 10042 30240 10048 30252
rect 9907 30212 10048 30240
rect 9907 30209 9919 30212
rect 9861 30203 9919 30209
rect 10042 30200 10048 30212
rect 10100 30200 10106 30252
rect 10594 30200 10600 30252
rect 10652 30240 10658 30252
rect 13004 30240 13032 30280
rect 13538 30268 13544 30320
rect 13596 30308 13602 30320
rect 13909 30311 13967 30317
rect 13909 30308 13921 30311
rect 13596 30280 13921 30308
rect 13596 30268 13602 30280
rect 13909 30277 13921 30280
rect 13955 30277 13967 30311
rect 13909 30271 13967 30277
rect 13725 30243 13783 30249
rect 13725 30240 13737 30243
rect 10652 30212 12940 30240
rect 13004 30212 13737 30240
rect 10652 30200 10658 30212
rect 9769 30175 9827 30181
rect 7392 30144 7880 30172
rect 5534 29996 5540 30048
rect 5592 29996 5598 30048
rect 5721 30039 5779 30045
rect 5721 30005 5733 30039
rect 5767 30036 5779 30039
rect 7006 30036 7012 30048
rect 5767 30008 7012 30036
rect 5767 30005 5779 30008
rect 5721 29999 5779 30005
rect 7006 29996 7012 30008
rect 7064 29996 7070 30048
rect 7742 29996 7748 30048
rect 7800 29996 7806 30048
rect 7852 30036 7880 30144
rect 9769 30141 9781 30175
rect 9815 30172 9827 30175
rect 10781 30175 10839 30181
rect 10781 30172 10793 30175
rect 9815 30144 10793 30172
rect 9815 30141 9827 30144
rect 9769 30135 9827 30141
rect 10781 30141 10793 30144
rect 10827 30141 10839 30175
rect 11241 30175 11299 30181
rect 11241 30172 11253 30175
rect 10781 30135 10839 30141
rect 10888 30144 11253 30172
rect 10137 30107 10195 30113
rect 10137 30104 10149 30107
rect 9784 30076 10149 30104
rect 8846 30036 8852 30048
rect 7852 30008 8852 30036
rect 8846 29996 8852 30008
rect 8904 29996 8910 30048
rect 9784 30045 9812 30076
rect 10137 30073 10149 30076
rect 10183 30073 10195 30107
rect 10137 30067 10195 30073
rect 10686 30064 10692 30116
rect 10744 30064 10750 30116
rect 9769 30039 9827 30045
rect 9769 30005 9781 30039
rect 9815 30005 9827 30039
rect 9769 29999 9827 30005
rect 9858 29996 9864 30048
rect 9916 30036 9922 30048
rect 10045 30039 10103 30045
rect 10045 30036 10057 30039
rect 9916 30008 10057 30036
rect 9916 29996 9922 30008
rect 10045 30005 10057 30008
rect 10091 30005 10103 30039
rect 10045 29999 10103 30005
rect 10318 29996 10324 30048
rect 10376 30036 10382 30048
rect 10888 30036 10916 30144
rect 11241 30141 11253 30144
rect 11287 30141 11299 30175
rect 11241 30135 11299 30141
rect 11330 30132 11336 30184
rect 11388 30172 11394 30184
rect 11977 30175 12035 30181
rect 11977 30172 11989 30175
rect 11388 30144 11989 30172
rect 11388 30132 11394 30144
rect 11977 30141 11989 30144
rect 12023 30141 12035 30175
rect 11977 30135 12035 30141
rect 12069 30175 12127 30181
rect 12069 30141 12081 30175
rect 12115 30172 12127 30175
rect 12710 30172 12716 30184
rect 12115 30144 12716 30172
rect 12115 30141 12127 30144
rect 12069 30135 12127 30141
rect 10962 30064 10968 30116
rect 11020 30064 11026 30116
rect 11054 30064 11060 30116
rect 11112 30104 11118 30116
rect 12084 30104 12112 30135
rect 12710 30132 12716 30144
rect 12768 30132 12774 30184
rect 12805 30175 12863 30181
rect 12805 30141 12817 30175
rect 12851 30141 12863 30175
rect 12805 30135 12863 30141
rect 11112 30076 12112 30104
rect 11112 30064 11118 30076
rect 12342 30064 12348 30116
rect 12400 30104 12406 30116
rect 12820 30104 12848 30135
rect 12400 30076 12848 30104
rect 12912 30104 12940 30212
rect 13725 30209 13737 30212
rect 13771 30209 13783 30243
rect 13725 30203 13783 30209
rect 14090 30200 14096 30252
rect 14148 30240 14154 30252
rect 14185 30243 14243 30249
rect 14185 30240 14197 30243
rect 14148 30212 14197 30240
rect 14148 30200 14154 30212
rect 14185 30209 14197 30212
rect 14231 30209 14243 30243
rect 14185 30203 14243 30209
rect 14274 30200 14280 30252
rect 14332 30200 14338 30252
rect 14369 30243 14427 30249
rect 14369 30209 14381 30243
rect 14415 30209 14427 30243
rect 14369 30203 14427 30209
rect 12989 30175 13047 30181
rect 12989 30141 13001 30175
rect 13035 30172 13047 30175
rect 13078 30172 13084 30184
rect 13035 30144 13084 30172
rect 13035 30141 13047 30144
rect 12989 30135 13047 30141
rect 13078 30132 13084 30144
rect 13136 30132 13142 30184
rect 13170 30132 13176 30184
rect 13228 30172 13234 30184
rect 14384 30172 14412 30203
rect 14550 30200 14556 30252
rect 14608 30200 14614 30252
rect 14829 30243 14887 30249
rect 14829 30209 14841 30243
rect 14875 30209 14887 30243
rect 14829 30203 14887 30209
rect 13228 30144 14412 30172
rect 13228 30132 13234 30144
rect 14458 30132 14464 30184
rect 14516 30172 14522 30184
rect 14844 30172 14872 30203
rect 14918 30200 14924 30252
rect 14976 30200 14982 30252
rect 15010 30200 15016 30252
rect 15068 30200 15074 30252
rect 15188 30243 15246 30249
rect 15188 30209 15200 30243
rect 15234 30240 15246 30243
rect 15562 30240 15568 30252
rect 15234 30212 15568 30240
rect 15234 30209 15246 30212
rect 15188 30203 15246 30209
rect 15562 30200 15568 30212
rect 15620 30200 15626 30252
rect 15028 30172 15056 30200
rect 14516 30144 14872 30172
rect 14936 30144 15056 30172
rect 14516 30132 14522 30144
rect 14645 30107 14703 30113
rect 14645 30104 14657 30107
rect 12912 30076 14657 30104
rect 12400 30064 12406 30076
rect 14645 30073 14657 30076
rect 14691 30073 14703 30107
rect 14645 30067 14703 30073
rect 10376 30008 10916 30036
rect 10376 29996 10382 30008
rect 12158 29996 12164 30048
rect 12216 30036 12222 30048
rect 13173 30039 13231 30045
rect 13173 30036 13185 30039
rect 12216 30008 13185 30036
rect 12216 29996 12222 30008
rect 13173 30005 13185 30008
rect 13219 30005 13231 30039
rect 13173 29999 13231 30005
rect 14090 29996 14096 30048
rect 14148 30036 14154 30048
rect 14936 30036 14964 30144
rect 15838 30036 15844 30048
rect 14148 30008 15844 30036
rect 14148 29996 14154 30008
rect 15838 29996 15844 30008
rect 15896 29996 15902 30048
rect 1104 29946 16652 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 16652 29946
rect 1104 29872 16652 29894
rect 6086 29792 6092 29844
rect 6144 29792 6150 29844
rect 7098 29792 7104 29844
rect 7156 29832 7162 29844
rect 7374 29832 7380 29844
rect 7156 29804 7380 29832
rect 7156 29792 7162 29804
rect 7374 29792 7380 29804
rect 7432 29832 7438 29844
rect 7834 29832 7840 29844
rect 7432 29804 7840 29832
rect 7432 29792 7438 29804
rect 7834 29792 7840 29804
rect 7892 29792 7898 29844
rect 9217 29835 9275 29841
rect 9217 29801 9229 29835
rect 9263 29832 9275 29835
rect 9490 29832 9496 29844
rect 9263 29804 9496 29832
rect 9263 29801 9275 29804
rect 9217 29795 9275 29801
rect 9490 29792 9496 29804
rect 9548 29792 9554 29844
rect 9950 29792 9956 29844
rect 10008 29792 10014 29844
rect 10137 29835 10195 29841
rect 10137 29801 10149 29835
rect 10183 29832 10195 29835
rect 10318 29832 10324 29844
rect 10183 29804 10324 29832
rect 10183 29801 10195 29804
rect 10137 29795 10195 29801
rect 6641 29767 6699 29773
rect 6641 29764 6653 29767
rect 5920 29736 6653 29764
rect 5920 29628 5948 29736
rect 6641 29733 6653 29736
rect 6687 29764 6699 29767
rect 7190 29764 7196 29776
rect 6687 29736 7196 29764
rect 6687 29733 6699 29736
rect 6641 29727 6699 29733
rect 7190 29724 7196 29736
rect 7248 29724 7254 29776
rect 9582 29724 9588 29776
rect 9640 29764 9646 29776
rect 10152 29764 10180 29795
rect 10318 29792 10324 29804
rect 10376 29792 10382 29844
rect 10410 29792 10416 29844
rect 10468 29832 10474 29844
rect 10597 29835 10655 29841
rect 10597 29832 10609 29835
rect 10468 29804 10609 29832
rect 10468 29792 10474 29804
rect 10597 29801 10609 29804
rect 10643 29801 10655 29835
rect 12986 29832 12992 29844
rect 10597 29795 10655 29801
rect 11348 29804 12992 29832
rect 10781 29767 10839 29773
rect 9640 29736 10272 29764
rect 9640 29724 9646 29736
rect 5997 29699 6055 29705
rect 5997 29665 6009 29699
rect 6043 29696 6055 29699
rect 7742 29696 7748 29708
rect 6043 29668 7748 29696
rect 6043 29665 6055 29668
rect 5997 29659 6055 29665
rect 7742 29656 7748 29668
rect 7800 29696 7806 29708
rect 7837 29699 7895 29705
rect 7837 29696 7849 29699
rect 7800 29668 7849 29696
rect 7800 29656 7806 29668
rect 7837 29665 7849 29668
rect 7883 29665 7895 29699
rect 7837 29659 7895 29665
rect 8110 29656 8116 29708
rect 8168 29696 8174 29708
rect 9950 29696 9956 29708
rect 8168 29668 9956 29696
rect 8168 29656 8174 29668
rect 9950 29656 9956 29668
rect 10008 29696 10014 29708
rect 10134 29696 10140 29708
rect 10008 29668 10140 29696
rect 10008 29656 10014 29668
rect 10134 29656 10140 29668
rect 10192 29656 10198 29708
rect 10244 29696 10272 29736
rect 10781 29733 10793 29767
rect 10827 29764 10839 29767
rect 11238 29764 11244 29776
rect 10827 29736 11244 29764
rect 10827 29733 10839 29736
rect 10781 29727 10839 29733
rect 11238 29724 11244 29736
rect 11296 29724 11302 29776
rect 11057 29699 11115 29705
rect 11057 29696 11069 29699
rect 10244 29668 11069 29696
rect 11057 29665 11069 29668
rect 11103 29696 11115 29699
rect 11146 29696 11152 29708
rect 11103 29668 11152 29696
rect 11103 29665 11115 29668
rect 11057 29659 11115 29665
rect 11146 29656 11152 29668
rect 11204 29656 11210 29708
rect 6089 29631 6147 29637
rect 6089 29628 6101 29631
rect 5920 29600 6101 29628
rect 6089 29597 6101 29600
rect 6135 29597 6147 29631
rect 6089 29591 6147 29597
rect 6178 29588 6184 29640
rect 6236 29628 6242 29640
rect 6236 29600 6500 29628
rect 6236 29588 6242 29600
rect 6365 29563 6423 29569
rect 6365 29529 6377 29563
rect 6411 29529 6423 29563
rect 6472 29560 6500 29600
rect 6914 29588 6920 29640
rect 6972 29588 6978 29640
rect 7193 29638 7251 29639
rect 7193 29633 7420 29638
rect 7193 29599 7205 29633
rect 7239 29610 7420 29633
rect 7239 29599 7251 29610
rect 7193 29593 7251 29599
rect 7098 29560 7104 29572
rect 6472 29532 7104 29560
rect 6365 29523 6423 29529
rect 5718 29452 5724 29504
rect 5776 29452 5782 29504
rect 6086 29452 6092 29504
rect 6144 29492 6150 29504
rect 6380 29492 6408 29523
rect 7098 29520 7104 29532
rect 7156 29520 7162 29572
rect 7392 29560 7420 29610
rect 8846 29588 8852 29640
rect 8904 29628 8910 29640
rect 8941 29631 8999 29637
rect 8941 29628 8953 29631
rect 8904 29600 8953 29628
rect 8904 29588 8910 29600
rect 8941 29597 8953 29600
rect 8987 29597 8999 29631
rect 8941 29591 8999 29597
rect 9125 29631 9183 29637
rect 9125 29597 9137 29631
rect 9171 29628 9183 29631
rect 9214 29628 9220 29640
rect 9171 29600 9220 29628
rect 9171 29597 9183 29600
rect 9125 29591 9183 29597
rect 9140 29560 9168 29591
rect 9214 29588 9220 29600
rect 9272 29588 9278 29640
rect 9398 29588 9404 29640
rect 9456 29628 9462 29640
rect 9493 29631 9551 29637
rect 9493 29628 9505 29631
rect 9456 29600 9505 29628
rect 9456 29588 9462 29600
rect 9493 29597 9505 29600
rect 9539 29597 9551 29631
rect 9493 29591 9551 29597
rect 7392 29532 9168 29560
rect 9508 29560 9536 29591
rect 9582 29588 9588 29640
rect 9640 29588 9646 29640
rect 9677 29631 9735 29637
rect 9677 29597 9689 29631
rect 9723 29628 9735 29631
rect 9766 29628 9772 29640
rect 9723 29600 9772 29628
rect 9723 29597 9735 29600
rect 9677 29591 9735 29597
rect 9766 29588 9772 29600
rect 9824 29588 9830 29640
rect 9858 29588 9864 29640
rect 9916 29588 9922 29640
rect 10505 29631 10563 29637
rect 10505 29597 10517 29631
rect 10551 29628 10563 29631
rect 10686 29628 10692 29640
rect 10551 29600 10692 29628
rect 10551 29597 10563 29600
rect 10505 29591 10563 29597
rect 10520 29560 10548 29591
rect 10686 29588 10692 29600
rect 10744 29588 10750 29640
rect 11348 29637 11376 29804
rect 12986 29792 12992 29804
rect 13044 29832 13050 29844
rect 14090 29832 14096 29844
rect 13044 29804 14096 29832
rect 13044 29792 13050 29804
rect 14090 29792 14096 29804
rect 14148 29792 14154 29844
rect 14826 29792 14832 29844
rect 14884 29792 14890 29844
rect 15562 29792 15568 29844
rect 15620 29792 15626 29844
rect 11790 29724 11796 29776
rect 11848 29724 11854 29776
rect 12250 29724 12256 29776
rect 12308 29764 12314 29776
rect 12308 29736 16068 29764
rect 12308 29724 12314 29736
rect 12342 29696 12348 29708
rect 11808 29668 12348 29696
rect 11333 29631 11391 29637
rect 11333 29597 11345 29631
rect 11379 29597 11391 29631
rect 11333 29591 11391 29597
rect 11422 29588 11428 29640
rect 11480 29588 11486 29640
rect 11606 29588 11612 29640
rect 11664 29588 11670 29640
rect 11698 29588 11704 29640
rect 11756 29588 11762 29640
rect 9508 29532 10548 29560
rect 11149 29563 11207 29569
rect 11149 29529 11161 29563
rect 11195 29560 11207 29563
rect 11808 29560 11836 29668
rect 12342 29656 12348 29668
rect 12400 29656 12406 29708
rect 12437 29699 12495 29705
rect 12437 29665 12449 29699
rect 12483 29696 12495 29699
rect 12710 29696 12716 29708
rect 12483 29668 12716 29696
rect 12483 29665 12495 29668
rect 12437 29659 12495 29665
rect 12710 29656 12716 29668
rect 12768 29696 12774 29708
rect 13078 29696 13084 29708
rect 12768 29668 13084 29696
rect 12768 29656 12774 29668
rect 13078 29656 13084 29668
rect 13136 29696 13142 29708
rect 13173 29699 13231 29705
rect 13173 29696 13185 29699
rect 13136 29668 13185 29696
rect 13136 29656 13142 29668
rect 13173 29665 13185 29668
rect 13219 29665 13231 29699
rect 13173 29659 13231 29665
rect 13262 29656 13268 29708
rect 13320 29696 13326 29708
rect 14366 29696 14372 29708
rect 13320 29668 14372 29696
rect 13320 29656 13326 29668
rect 14366 29656 14372 29668
rect 14424 29696 14430 29708
rect 15654 29696 15660 29708
rect 14424 29668 15148 29696
rect 14424 29656 14430 29668
rect 12158 29588 12164 29640
rect 12216 29588 12222 29640
rect 12989 29631 13047 29637
rect 12989 29597 13001 29631
rect 13035 29628 13047 29631
rect 14093 29631 14151 29637
rect 14093 29628 14105 29631
rect 13035 29600 14105 29628
rect 13035 29597 13047 29600
rect 12989 29591 13047 29597
rect 14093 29597 14105 29600
rect 14139 29597 14151 29631
rect 14093 29591 14151 29597
rect 14737 29631 14795 29637
rect 14737 29597 14749 29631
rect 14783 29628 14795 29631
rect 14826 29628 14832 29640
rect 14783 29600 14832 29628
rect 14783 29597 14795 29600
rect 14737 29591 14795 29597
rect 11195 29532 11836 29560
rect 12253 29563 12311 29569
rect 11195 29529 11207 29532
rect 11149 29523 11207 29529
rect 12253 29529 12265 29563
rect 12299 29560 12311 29563
rect 13446 29560 13452 29572
rect 12299 29532 13452 29560
rect 12299 29529 12311 29532
rect 12253 29523 12311 29529
rect 13446 29520 13452 29532
rect 13504 29520 13510 29572
rect 13538 29520 13544 29572
rect 13596 29520 13602 29572
rect 13722 29520 13728 29572
rect 13780 29520 13786 29572
rect 14752 29560 14780 29591
rect 14826 29588 14832 29600
rect 14884 29588 14890 29640
rect 15120 29637 15148 29668
rect 15212 29668 15660 29696
rect 15212 29637 15240 29668
rect 15654 29656 15660 29668
rect 15712 29696 15718 29708
rect 15712 29668 15976 29696
rect 15712 29656 15718 29668
rect 15105 29631 15163 29637
rect 15105 29597 15117 29631
rect 15151 29597 15163 29631
rect 15105 29591 15163 29597
rect 15197 29631 15255 29637
rect 15197 29597 15209 29631
rect 15243 29597 15255 29631
rect 15197 29591 15255 29597
rect 15286 29588 15292 29640
rect 15344 29588 15350 29640
rect 15473 29631 15531 29637
rect 15473 29628 15485 29631
rect 15396 29600 15485 29628
rect 13832 29532 14780 29560
rect 15396 29560 15424 29600
rect 15473 29597 15485 29600
rect 15519 29597 15531 29631
rect 15473 29591 15531 29597
rect 15838 29588 15844 29640
rect 15896 29588 15902 29640
rect 15948 29637 15976 29668
rect 16040 29637 16068 29736
rect 15933 29631 15991 29637
rect 15933 29597 15945 29631
rect 15979 29597 15991 29631
rect 15933 29591 15991 29597
rect 16025 29631 16083 29637
rect 16025 29597 16037 29631
rect 16071 29597 16083 29631
rect 16025 29591 16083 29597
rect 16209 29631 16267 29637
rect 16209 29597 16221 29631
rect 16255 29597 16267 29631
rect 16209 29591 16267 29597
rect 16224 29560 16252 29591
rect 15396 29532 16252 29560
rect 6144 29464 6408 29492
rect 6549 29495 6607 29501
rect 6144 29452 6150 29464
rect 6549 29461 6561 29495
rect 6595 29492 6607 29495
rect 6730 29492 6736 29504
rect 6595 29464 6736 29492
rect 6595 29461 6607 29464
rect 6549 29455 6607 29461
rect 6730 29452 6736 29464
rect 6788 29452 6794 29504
rect 6914 29452 6920 29504
rect 6972 29492 6978 29504
rect 7285 29495 7343 29501
rect 7285 29492 7297 29495
rect 6972 29464 7297 29492
rect 6972 29452 6978 29464
rect 7285 29461 7297 29464
rect 7331 29461 7343 29495
rect 7285 29455 7343 29461
rect 8662 29452 8668 29504
rect 8720 29452 8726 29504
rect 9030 29452 9036 29504
rect 9088 29452 9094 29504
rect 10137 29495 10195 29501
rect 10137 29461 10149 29495
rect 10183 29492 10195 29495
rect 10318 29492 10324 29504
rect 10183 29464 10324 29492
rect 10183 29461 10195 29464
rect 10137 29455 10195 29461
rect 10318 29452 10324 29464
rect 10376 29452 10382 29504
rect 10502 29452 10508 29504
rect 10560 29492 10566 29504
rect 12526 29492 12532 29504
rect 10560 29464 12532 29492
rect 10560 29452 10566 29464
rect 12526 29452 12532 29464
rect 12584 29452 12590 29504
rect 12618 29452 12624 29504
rect 12676 29452 12682 29504
rect 12894 29452 12900 29504
rect 12952 29492 12958 29504
rect 13081 29495 13139 29501
rect 13081 29492 13093 29495
rect 12952 29464 13093 29492
rect 12952 29452 12958 29464
rect 13081 29461 13093 29464
rect 13127 29492 13139 29495
rect 13262 29492 13268 29504
rect 13127 29464 13268 29492
rect 13127 29461 13139 29464
rect 13081 29455 13139 29461
rect 13262 29452 13268 29464
rect 13320 29452 13326 29504
rect 13630 29452 13636 29504
rect 13688 29492 13694 29504
rect 13832 29492 13860 29532
rect 13688 29464 13860 29492
rect 13909 29495 13967 29501
rect 13688 29452 13694 29464
rect 13909 29461 13921 29495
rect 13955 29492 13967 29495
rect 14274 29492 14280 29504
rect 13955 29464 14280 29492
rect 13955 29461 13967 29464
rect 13909 29455 13967 29461
rect 14274 29452 14280 29464
rect 14332 29452 14338 29504
rect 14550 29452 14556 29504
rect 14608 29492 14614 29504
rect 15396 29492 15424 29532
rect 14608 29464 15424 29492
rect 14608 29452 14614 29464
rect 1104 29402 16652 29424
rect 1104 29350 4874 29402
rect 4926 29350 4938 29402
rect 4990 29350 5002 29402
rect 5054 29350 5066 29402
rect 5118 29350 5130 29402
rect 5182 29350 16652 29402
rect 1104 29328 16652 29350
rect 6549 29291 6607 29297
rect 6549 29257 6561 29291
rect 6595 29288 6607 29291
rect 6638 29288 6644 29300
rect 6595 29260 6644 29288
rect 6595 29257 6607 29260
rect 6549 29251 6607 29257
rect 6638 29248 6644 29260
rect 6696 29248 6702 29300
rect 6730 29248 6736 29300
rect 6788 29288 6794 29300
rect 8386 29288 8392 29300
rect 6788 29260 8392 29288
rect 6788 29248 6794 29260
rect 8386 29248 8392 29260
rect 8444 29248 8450 29300
rect 8662 29248 8668 29300
rect 8720 29288 8726 29300
rect 9125 29291 9183 29297
rect 9125 29288 9137 29291
rect 8720 29260 9137 29288
rect 8720 29248 8726 29260
rect 9125 29257 9137 29260
rect 9171 29257 9183 29291
rect 9125 29251 9183 29257
rect 10870 29248 10876 29300
rect 10928 29288 10934 29300
rect 10965 29291 11023 29297
rect 10965 29288 10977 29291
rect 10928 29260 10977 29288
rect 10928 29248 10934 29260
rect 10965 29257 10977 29260
rect 11011 29257 11023 29291
rect 10965 29251 11023 29257
rect 11133 29291 11191 29297
rect 11133 29257 11145 29291
rect 11179 29288 11191 29291
rect 11606 29288 11612 29300
rect 11179 29260 11612 29288
rect 11179 29257 11191 29260
rect 11133 29251 11191 29257
rect 11606 29248 11612 29260
rect 11664 29248 11670 29300
rect 13630 29248 13636 29300
rect 13688 29248 13694 29300
rect 14090 29248 14096 29300
rect 14148 29288 14154 29300
rect 14642 29288 14648 29300
rect 14148 29260 14648 29288
rect 14148 29248 14154 29260
rect 14642 29248 14648 29260
rect 14700 29288 14706 29300
rect 14700 29260 15700 29288
rect 14700 29248 14706 29260
rect 5902 29180 5908 29232
rect 5960 29220 5966 29232
rect 6822 29220 6828 29232
rect 5960 29192 6828 29220
rect 5960 29180 5966 29192
rect 6822 29180 6828 29192
rect 6880 29220 6886 29232
rect 6880 29192 7052 29220
rect 6880 29180 6886 29192
rect 5534 29112 5540 29164
rect 5592 29152 5598 29164
rect 6638 29152 6644 29164
rect 5592 29124 6644 29152
rect 5592 29112 5598 29124
rect 6638 29112 6644 29124
rect 6696 29152 6702 29164
rect 6696 29124 6868 29152
rect 6696 29112 6702 29124
rect 6840 29093 6868 29124
rect 6914 29112 6920 29164
rect 6972 29112 6978 29164
rect 7024 29161 7052 29192
rect 7926 29180 7932 29232
rect 7984 29220 7990 29232
rect 7984 29192 8708 29220
rect 7984 29180 7990 29192
rect 8680 29161 8708 29192
rect 9030 29180 9036 29232
rect 9088 29220 9094 29232
rect 9088 29192 9260 29220
rect 9088 29180 9094 29192
rect 7009 29155 7067 29161
rect 7009 29121 7021 29155
rect 7055 29121 7067 29155
rect 7009 29115 7067 29121
rect 8409 29155 8467 29161
rect 8409 29121 8421 29155
rect 8455 29152 8467 29155
rect 8665 29155 8723 29161
rect 8455 29124 8616 29152
rect 8455 29121 8467 29124
rect 8409 29115 8467 29121
rect 6733 29087 6791 29093
rect 6733 29053 6745 29087
rect 6779 29053 6791 29087
rect 6733 29047 6791 29053
rect 6825 29087 6883 29093
rect 6825 29053 6837 29087
rect 6871 29053 6883 29087
rect 8588 29084 8616 29124
rect 8665 29121 8677 29155
rect 8711 29121 8723 29155
rect 8665 29115 8723 29121
rect 8938 29112 8944 29164
rect 8996 29112 9002 29164
rect 9232 29161 9260 29192
rect 10686 29180 10692 29232
rect 10744 29220 10750 29232
rect 11333 29223 11391 29229
rect 11333 29220 11345 29223
rect 10744 29192 11345 29220
rect 10744 29180 10750 29192
rect 11333 29189 11345 29192
rect 11379 29189 11391 29223
rect 11333 29183 11391 29189
rect 12520 29223 12578 29229
rect 12520 29189 12532 29223
rect 12566 29220 12578 29223
rect 12618 29220 12624 29232
rect 12566 29192 12624 29220
rect 12566 29189 12578 29192
rect 12520 29183 12578 29189
rect 12618 29180 12624 29192
rect 12676 29180 12682 29232
rect 13354 29180 13360 29232
rect 13412 29220 13418 29232
rect 15470 29220 15476 29232
rect 13412 29192 14780 29220
rect 13412 29180 13418 29192
rect 9217 29155 9275 29161
rect 9217 29121 9229 29155
rect 9263 29121 9275 29155
rect 9217 29115 9275 29121
rect 9493 29155 9551 29161
rect 9493 29121 9505 29155
rect 9539 29152 9551 29155
rect 9582 29152 9588 29164
rect 9539 29124 9588 29152
rect 9539 29121 9551 29124
rect 9493 29115 9551 29121
rect 9582 29112 9588 29124
rect 9640 29112 9646 29164
rect 9760 29155 9818 29161
rect 9760 29121 9772 29155
rect 9806 29152 9818 29155
rect 10134 29152 10140 29164
rect 9806 29124 10140 29152
rect 9806 29121 9818 29124
rect 9760 29115 9818 29121
rect 10134 29112 10140 29124
rect 10192 29112 10198 29164
rect 14369 29155 14427 29161
rect 14369 29121 14381 29155
rect 14415 29152 14427 29155
rect 14458 29152 14464 29164
rect 14415 29124 14464 29152
rect 14415 29121 14427 29124
rect 14369 29115 14427 29121
rect 14458 29112 14464 29124
rect 14516 29112 14522 29164
rect 14642 29112 14648 29164
rect 14700 29112 14706 29164
rect 14752 29161 14780 29192
rect 14936 29192 15476 29220
rect 14936 29161 14964 29192
rect 15470 29180 15476 29192
rect 15528 29180 15534 29232
rect 14737 29155 14795 29161
rect 14737 29121 14749 29155
rect 14783 29121 14795 29155
rect 14737 29115 14795 29121
rect 14921 29155 14979 29161
rect 14921 29121 14933 29155
rect 14967 29121 14979 29155
rect 14921 29115 14979 29121
rect 15010 29112 15016 29164
rect 15068 29112 15074 29164
rect 15105 29156 15163 29161
rect 15286 29156 15292 29164
rect 15105 29155 15292 29156
rect 15105 29121 15117 29155
rect 15151 29128 15292 29155
rect 15151 29121 15163 29128
rect 15105 29115 15163 29121
rect 15286 29112 15292 29128
rect 15344 29112 15350 29164
rect 15672 29161 15700 29260
rect 15930 29248 15936 29300
rect 15988 29288 15994 29300
rect 16117 29291 16175 29297
rect 16117 29288 16129 29291
rect 15988 29260 16129 29288
rect 15988 29248 15994 29260
rect 16117 29257 16129 29260
rect 16163 29257 16175 29291
rect 16117 29251 16175 29257
rect 15657 29155 15715 29161
rect 15657 29121 15669 29155
rect 15703 29121 15715 29155
rect 15657 29115 15715 29121
rect 15749 29155 15807 29161
rect 15749 29121 15761 29155
rect 15795 29121 15807 29155
rect 15749 29115 15807 29121
rect 8757 29087 8815 29093
rect 8757 29084 8769 29087
rect 8588 29056 8769 29084
rect 6825 29047 6883 29053
rect 8757 29053 8769 29056
rect 8803 29053 8815 29087
rect 8757 29047 8815 29053
rect 12069 29087 12127 29093
rect 12069 29053 12081 29087
rect 12115 29053 12127 29087
rect 12069 29047 12127 29053
rect 6748 29016 6776 29047
rect 7190 29016 7196 29028
rect 6748 28988 7196 29016
rect 7190 28976 7196 28988
rect 7248 28976 7254 29028
rect 7282 28976 7288 29028
rect 7340 28976 7346 29028
rect 10778 28976 10784 29028
rect 10836 29016 10842 29028
rect 10873 29019 10931 29025
rect 10873 29016 10885 29019
rect 10836 28988 10885 29016
rect 10836 28976 10842 28988
rect 10873 28985 10885 28988
rect 10919 29016 10931 29019
rect 12084 29016 12112 29047
rect 12250 29044 12256 29096
rect 12308 29044 12314 29096
rect 13722 29044 13728 29096
rect 13780 29084 13786 29096
rect 15470 29084 15476 29096
rect 13780 29056 15476 29084
rect 13780 29044 13786 29056
rect 15470 29044 15476 29056
rect 15528 29084 15534 29096
rect 15764 29084 15792 29115
rect 15930 29112 15936 29164
rect 15988 29112 15994 29164
rect 16022 29112 16028 29164
rect 16080 29112 16086 29164
rect 16298 29112 16304 29164
rect 16356 29112 16362 29164
rect 15528 29056 15792 29084
rect 15528 29044 15534 29056
rect 10919 28988 12112 29016
rect 10919 28985 10931 28988
rect 10873 28979 10931 28985
rect 13446 28976 13452 29028
rect 13504 29016 13510 29028
rect 13504 28988 13860 29016
rect 13504 28976 13510 28988
rect 9030 28908 9036 28960
rect 9088 28948 9094 28960
rect 9490 28948 9496 28960
rect 9088 28920 9496 28948
rect 9088 28908 9094 28920
rect 9490 28908 9496 28920
rect 9548 28908 9554 28960
rect 11146 28908 11152 28960
rect 11204 28908 11210 28960
rect 11514 28908 11520 28960
rect 11572 28908 11578 28960
rect 13722 28908 13728 28960
rect 13780 28908 13786 28960
rect 13832 28948 13860 28988
rect 14826 28976 14832 29028
rect 14884 29016 14890 29028
rect 15194 29016 15200 29028
rect 14884 28988 15200 29016
rect 14884 28976 14890 28988
rect 15194 28976 15200 28988
rect 15252 28976 15258 29028
rect 15289 29019 15347 29025
rect 15289 28985 15301 29019
rect 15335 29016 15347 29019
rect 15378 29016 15384 29028
rect 15335 28988 15384 29016
rect 15335 28985 15347 28988
rect 15289 28979 15347 28985
rect 15378 28976 15384 28988
rect 15436 28976 15442 29028
rect 14461 28951 14519 28957
rect 14461 28948 14473 28951
rect 13832 28920 14473 28948
rect 14461 28917 14473 28920
rect 14507 28917 14519 28951
rect 14461 28911 14519 28917
rect 14550 28908 14556 28960
rect 14608 28948 14614 28960
rect 15473 28951 15531 28957
rect 15473 28948 15485 28951
rect 14608 28920 15485 28948
rect 14608 28908 14614 28920
rect 15473 28917 15485 28920
rect 15519 28917 15531 28951
rect 15473 28911 15531 28917
rect 1104 28858 16652 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 16652 28858
rect 1104 28784 16652 28806
rect 6822 28704 6828 28756
rect 6880 28704 6886 28756
rect 7101 28747 7159 28753
rect 7101 28713 7113 28747
rect 7147 28744 7159 28747
rect 8938 28744 8944 28756
rect 7147 28716 8944 28744
rect 7147 28713 7159 28716
rect 7101 28707 7159 28713
rect 8938 28704 8944 28716
rect 8996 28704 9002 28756
rect 9030 28704 9036 28756
rect 9088 28744 9094 28756
rect 9125 28747 9183 28753
rect 9125 28744 9137 28747
rect 9088 28716 9137 28744
rect 9088 28704 9094 28716
rect 9125 28713 9137 28716
rect 9171 28713 9183 28747
rect 9125 28707 9183 28713
rect 9309 28747 9367 28753
rect 9309 28713 9321 28747
rect 9355 28744 9367 28747
rect 10042 28744 10048 28756
rect 9355 28716 10048 28744
rect 9355 28713 9367 28716
rect 9309 28707 9367 28713
rect 10042 28704 10048 28716
rect 10100 28704 10106 28756
rect 10134 28704 10140 28756
rect 10192 28704 10198 28756
rect 13725 28747 13783 28753
rect 13725 28713 13737 28747
rect 13771 28744 13783 28747
rect 14458 28744 14464 28756
rect 13771 28716 14464 28744
rect 13771 28713 13783 28716
rect 13725 28707 13783 28713
rect 14458 28704 14464 28716
rect 14516 28704 14522 28756
rect 15286 28704 15292 28756
rect 15344 28744 15350 28756
rect 16301 28747 16359 28753
rect 16301 28744 16313 28747
rect 15344 28716 16313 28744
rect 15344 28704 15350 28716
rect 16301 28713 16313 28716
rect 16347 28713 16359 28747
rect 16301 28707 16359 28713
rect 8757 28679 8815 28685
rect 8757 28645 8769 28679
rect 8803 28676 8815 28679
rect 9214 28676 9220 28688
rect 8803 28648 9220 28676
rect 8803 28645 8815 28648
rect 8757 28639 8815 28645
rect 9214 28636 9220 28648
rect 9272 28636 9278 28688
rect 9861 28679 9919 28685
rect 9861 28645 9873 28679
rect 9907 28676 9919 28679
rect 9907 28648 11192 28676
rect 9907 28645 9919 28648
rect 9861 28639 9919 28645
rect 7650 28568 7656 28620
rect 7708 28608 7714 28620
rect 8113 28611 8171 28617
rect 8113 28608 8125 28611
rect 7708 28580 8125 28608
rect 7708 28568 7714 28580
rect 8113 28577 8125 28580
rect 8159 28577 8171 28611
rect 8113 28571 8171 28577
rect 10226 28568 10232 28620
rect 10284 28608 10290 28620
rect 10689 28611 10747 28617
rect 10689 28608 10701 28611
rect 10284 28580 10701 28608
rect 10284 28568 10290 28580
rect 10689 28577 10701 28580
rect 10735 28577 10747 28611
rect 11164 28608 11192 28648
rect 13354 28636 13360 28688
rect 13412 28676 13418 28688
rect 14550 28676 14556 28688
rect 13412 28648 14556 28676
rect 13412 28636 13418 28648
rect 14550 28636 14556 28648
rect 14608 28636 14614 28688
rect 14642 28608 14648 28620
rect 11164 28580 12480 28608
rect 10689 28571 10747 28577
rect 5718 28500 5724 28552
rect 5776 28540 5782 28552
rect 6733 28543 6791 28549
rect 6733 28540 6745 28543
rect 5776 28512 6745 28540
rect 5776 28500 5782 28512
rect 6733 28509 6745 28512
rect 6779 28509 6791 28543
rect 6733 28503 6791 28509
rect 6822 28500 6828 28552
rect 6880 28540 6886 28552
rect 7009 28543 7067 28549
rect 7009 28540 7021 28543
rect 6880 28512 7021 28540
rect 6880 28500 6886 28512
rect 7009 28509 7021 28512
rect 7055 28509 7067 28543
rect 7009 28503 7067 28509
rect 7190 28500 7196 28552
rect 7248 28500 7254 28552
rect 8573 28543 8631 28549
rect 8573 28509 8585 28543
rect 8619 28509 8631 28543
rect 8573 28503 8631 28509
rect 8757 28543 8815 28549
rect 8757 28509 8769 28543
rect 8803 28540 8815 28543
rect 9030 28540 9036 28552
rect 8803 28512 9036 28540
rect 8803 28509 8815 28512
rect 8757 28503 8815 28509
rect 2958 28432 2964 28484
rect 3016 28472 3022 28484
rect 3329 28475 3387 28481
rect 3329 28472 3341 28475
rect 3016 28444 3341 28472
rect 3016 28432 3022 28444
rect 3329 28441 3341 28444
rect 3375 28441 3387 28475
rect 3329 28435 3387 28441
rect 3513 28475 3571 28481
rect 3513 28441 3525 28475
rect 3559 28472 3571 28475
rect 8202 28472 8208 28484
rect 3559 28444 8208 28472
rect 3559 28441 3571 28444
rect 3513 28435 3571 28441
rect 8202 28432 8208 28444
rect 8260 28432 8266 28484
rect 8588 28472 8616 28503
rect 9030 28500 9036 28512
rect 9088 28500 9094 28552
rect 10045 28543 10103 28549
rect 10045 28509 10057 28543
rect 10091 28540 10103 28543
rect 10502 28540 10508 28552
rect 10091 28512 10508 28540
rect 10091 28509 10103 28512
rect 10045 28503 10103 28509
rect 10502 28500 10508 28512
rect 10560 28500 10566 28552
rect 10597 28543 10655 28549
rect 10597 28509 10609 28543
rect 10643 28540 10655 28543
rect 11514 28540 11520 28552
rect 10643 28512 11520 28540
rect 10643 28509 10655 28512
rect 10597 28503 10655 28509
rect 11514 28500 11520 28512
rect 11572 28500 11578 28552
rect 11606 28500 11612 28552
rect 11664 28500 11670 28552
rect 12250 28500 12256 28552
rect 12308 28540 12314 28552
rect 12345 28543 12403 28549
rect 12345 28540 12357 28543
rect 12308 28512 12357 28540
rect 12308 28500 12314 28512
rect 12345 28509 12357 28512
rect 12391 28509 12403 28543
rect 12452 28540 12480 28580
rect 14108 28580 14648 28608
rect 14108 28549 14136 28580
rect 14642 28568 14648 28580
rect 14700 28608 14706 28620
rect 14826 28608 14832 28620
rect 14700 28580 14832 28608
rect 14700 28568 14706 28580
rect 14826 28568 14832 28580
rect 14884 28568 14890 28620
rect 14918 28568 14924 28620
rect 14976 28568 14982 28620
rect 14093 28543 14151 28549
rect 12452 28512 13124 28540
rect 12345 28503 12403 28509
rect 8941 28475 8999 28481
rect 8941 28472 8953 28475
rect 8588 28444 8953 28472
rect 8941 28441 8953 28444
rect 8987 28472 8999 28475
rect 9398 28472 9404 28484
rect 8987 28444 9404 28472
rect 8987 28441 8999 28444
rect 8941 28435 8999 28441
rect 9398 28432 9404 28444
rect 9456 28432 9462 28484
rect 9674 28432 9680 28484
rect 9732 28472 9738 28484
rect 10965 28475 11023 28481
rect 10965 28472 10977 28475
rect 9732 28444 10977 28472
rect 9732 28432 9738 28444
rect 10965 28441 10977 28444
rect 11011 28472 11023 28475
rect 12360 28472 12388 28503
rect 11011 28444 12388 28472
rect 12612 28475 12670 28481
rect 11011 28441 11023 28444
rect 10965 28435 11023 28441
rect 12612 28441 12624 28475
rect 12658 28472 12670 28475
rect 12986 28472 12992 28484
rect 12658 28444 12992 28472
rect 12658 28441 12670 28444
rect 12612 28435 12670 28441
rect 12986 28432 12992 28444
rect 13044 28432 13050 28484
rect 13096 28472 13124 28512
rect 14093 28509 14105 28543
rect 14139 28509 14151 28543
rect 14093 28503 14151 28509
rect 14274 28500 14280 28552
rect 14332 28500 14338 28552
rect 14366 28500 14372 28552
rect 14424 28500 14430 28552
rect 14461 28543 14519 28549
rect 14461 28509 14473 28543
rect 14507 28540 14519 28543
rect 15562 28540 15568 28552
rect 14507 28512 15568 28540
rect 14507 28509 14519 28512
rect 14461 28503 14519 28509
rect 15562 28500 15568 28512
rect 15620 28500 15626 28552
rect 15188 28475 15246 28481
rect 13096 28444 14872 28472
rect 7558 28364 7564 28416
rect 7616 28364 7622 28416
rect 8846 28364 8852 28416
rect 8904 28404 8910 28416
rect 9141 28407 9199 28413
rect 9141 28404 9153 28407
rect 8904 28376 9153 28404
rect 8904 28364 8910 28376
rect 9141 28373 9153 28376
rect 9187 28373 9199 28407
rect 9141 28367 9199 28373
rect 10502 28364 10508 28416
rect 10560 28364 10566 28416
rect 12253 28407 12311 28413
rect 12253 28373 12265 28407
rect 12299 28404 12311 28407
rect 12802 28404 12808 28416
rect 12299 28376 12808 28404
rect 12299 28373 12311 28376
rect 12253 28367 12311 28373
rect 12802 28364 12808 28376
rect 12860 28364 12866 28416
rect 14734 28364 14740 28416
rect 14792 28364 14798 28416
rect 14844 28404 14872 28444
rect 15188 28441 15200 28475
rect 15234 28472 15246 28475
rect 15286 28472 15292 28484
rect 15234 28444 15292 28472
rect 15234 28441 15246 28444
rect 15188 28435 15246 28441
rect 15286 28432 15292 28444
rect 15344 28432 15350 28484
rect 15378 28404 15384 28416
rect 14844 28376 15384 28404
rect 15378 28364 15384 28376
rect 15436 28364 15442 28416
rect 1104 28314 16652 28336
rect 1104 28262 4874 28314
rect 4926 28262 4938 28314
rect 4990 28262 5002 28314
rect 5054 28262 5066 28314
rect 5118 28262 5130 28314
rect 5182 28262 16652 28314
rect 1104 28240 16652 28262
rect 7745 28203 7803 28209
rect 7745 28169 7757 28203
rect 7791 28200 7803 28203
rect 7834 28200 7840 28212
rect 7791 28172 7840 28200
rect 7791 28169 7803 28172
rect 7745 28163 7803 28169
rect 7834 28160 7840 28172
rect 7892 28160 7898 28212
rect 8757 28203 8815 28209
rect 8757 28169 8769 28203
rect 8803 28200 8815 28203
rect 9122 28200 9128 28212
rect 8803 28172 9128 28200
rect 8803 28169 8815 28172
rect 8757 28163 8815 28169
rect 9122 28160 9128 28172
rect 9180 28160 9186 28212
rect 10502 28160 10508 28212
rect 10560 28200 10566 28212
rect 10597 28203 10655 28209
rect 10597 28200 10609 28203
rect 10560 28172 10609 28200
rect 10560 28160 10566 28172
rect 10597 28169 10609 28172
rect 10643 28169 10655 28203
rect 10597 28163 10655 28169
rect 10965 28203 11023 28209
rect 10965 28169 10977 28203
rect 11011 28200 11023 28203
rect 11517 28203 11575 28209
rect 11517 28200 11529 28203
rect 11011 28172 11529 28200
rect 11011 28169 11023 28172
rect 10965 28163 11023 28169
rect 11517 28169 11529 28172
rect 11563 28169 11575 28203
rect 11517 28163 11575 28169
rect 6825 28135 6883 28141
rect 6825 28101 6837 28135
rect 6871 28132 6883 28135
rect 7006 28132 7012 28144
rect 6871 28104 7012 28132
rect 6871 28101 6883 28104
rect 6825 28095 6883 28101
rect 7006 28092 7012 28104
rect 7064 28092 7070 28144
rect 8113 28135 8171 28141
rect 8113 28132 8125 28135
rect 7300 28104 8125 28132
rect 7300 28076 7328 28104
rect 8113 28101 8125 28104
rect 8159 28101 8171 28135
rect 8113 28095 8171 28101
rect 2590 28024 2596 28076
rect 2648 28064 2654 28076
rect 3033 28067 3091 28073
rect 3033 28064 3045 28067
rect 2648 28036 3045 28064
rect 2648 28024 2654 28036
rect 3033 28033 3045 28036
rect 3079 28033 3091 28067
rect 3033 28027 3091 28033
rect 3418 28024 3424 28076
rect 3476 28064 3482 28076
rect 4249 28067 4307 28073
rect 4249 28064 4261 28067
rect 3476 28036 4261 28064
rect 3476 28024 3482 28036
rect 4249 28033 4261 28036
rect 4295 28033 4307 28067
rect 4249 28027 4307 28033
rect 4433 28067 4491 28073
rect 4433 28033 4445 28067
rect 4479 28064 4491 28067
rect 4706 28064 4712 28076
rect 4479 28036 4712 28064
rect 4479 28033 4491 28036
rect 4433 28027 4491 28033
rect 4706 28024 4712 28036
rect 4764 28024 4770 28076
rect 6730 28024 6736 28076
rect 6788 28024 6794 28076
rect 6917 28067 6975 28073
rect 6917 28033 6929 28067
rect 6963 28064 6975 28067
rect 7098 28064 7104 28076
rect 6963 28036 7104 28064
rect 6963 28033 6975 28036
rect 6917 28027 6975 28033
rect 7098 28024 7104 28036
rect 7156 28024 7162 28076
rect 7282 28024 7288 28076
rect 7340 28024 7346 28076
rect 7561 28067 7619 28073
rect 7561 28033 7573 28067
rect 7607 28064 7619 28067
rect 7607 28036 7788 28064
rect 7607 28033 7619 28036
rect 7561 28027 7619 28033
rect 2774 27956 2780 28008
rect 2832 27956 2838 28008
rect 7190 27956 7196 28008
rect 7248 27956 7254 28008
rect 3786 27888 3792 27940
rect 3844 27928 3850 27940
rect 4249 27931 4307 27937
rect 4249 27928 4261 27931
rect 3844 27900 4261 27928
rect 3844 27888 3850 27900
rect 4249 27897 4261 27900
rect 4295 27897 4307 27931
rect 4249 27891 4307 27897
rect 5810 27888 5816 27940
rect 5868 27928 5874 27940
rect 7576 27928 7604 28027
rect 7653 27999 7711 28005
rect 7653 27965 7665 27999
rect 7699 27965 7711 27999
rect 7760 27996 7788 28036
rect 7834 28024 7840 28076
rect 7892 28064 7898 28076
rect 7929 28067 7987 28073
rect 7929 28064 7941 28067
rect 7892 28036 7941 28064
rect 7892 28024 7898 28036
rect 7929 28033 7941 28036
rect 7975 28033 7987 28067
rect 7929 28027 7987 28033
rect 8202 28024 8208 28076
rect 8260 28064 8266 28076
rect 8389 28067 8447 28073
rect 8389 28064 8401 28067
rect 8260 28036 8401 28064
rect 8260 28024 8266 28036
rect 8389 28033 8401 28036
rect 8435 28033 8447 28067
rect 8389 28027 8447 28033
rect 8754 28024 8760 28076
rect 8812 28064 8818 28076
rect 9125 28067 9183 28073
rect 9125 28064 9137 28067
rect 8812 28036 9137 28064
rect 8812 28024 8818 28036
rect 9125 28033 9137 28036
rect 9171 28033 9183 28067
rect 9125 28027 9183 28033
rect 7760 27968 8248 27996
rect 7653 27959 7711 27965
rect 5868 27900 7604 27928
rect 5868 27888 5874 27900
rect 3970 27820 3976 27872
rect 4028 27860 4034 27872
rect 4157 27863 4215 27869
rect 4157 27860 4169 27863
rect 4028 27832 4169 27860
rect 4028 27820 4034 27832
rect 4157 27829 4169 27832
rect 4203 27829 4215 27863
rect 4157 27823 4215 27829
rect 6914 27820 6920 27872
rect 6972 27860 6978 27872
rect 7009 27863 7067 27869
rect 7009 27860 7021 27863
rect 6972 27832 7021 27860
rect 6972 27820 6978 27832
rect 7009 27829 7021 27832
rect 7055 27829 7067 27863
rect 7668 27860 7696 27959
rect 8220 27937 8248 27968
rect 9214 27956 9220 28008
rect 9272 27956 9278 28008
rect 9401 27999 9459 28005
rect 9401 27965 9413 27999
rect 9447 27996 9459 27999
rect 9950 27996 9956 28008
rect 9447 27968 9956 27996
rect 9447 27965 9459 27968
rect 9401 27959 9459 27965
rect 9950 27956 9956 27968
rect 10008 27956 10014 28008
rect 10870 27956 10876 28008
rect 10928 27996 10934 28008
rect 11057 27999 11115 28005
rect 11057 27996 11069 27999
rect 10928 27968 11069 27996
rect 10928 27956 10934 27968
rect 11057 27965 11069 27968
rect 11103 27965 11115 27999
rect 11057 27959 11115 27965
rect 11146 27956 11152 28008
rect 11204 27956 11210 28008
rect 8205 27931 8263 27937
rect 8205 27897 8217 27931
rect 8251 27897 8263 27931
rect 8205 27891 8263 27897
rect 10226 27860 10232 27872
rect 7668 27832 10232 27860
rect 7009 27823 7067 27829
rect 10226 27820 10232 27832
rect 10284 27820 10290 27872
rect 11532 27860 11560 28163
rect 11974 28160 11980 28212
rect 12032 28200 12038 28212
rect 12032 28172 12940 28200
rect 12032 28160 12038 28172
rect 12250 28092 12256 28144
rect 12308 28132 12314 28144
rect 12912 28132 12940 28172
rect 12986 28160 12992 28212
rect 13044 28160 13050 28212
rect 13357 28203 13415 28209
rect 13357 28169 13369 28203
rect 13403 28200 13415 28203
rect 13722 28200 13728 28212
rect 13403 28172 13728 28200
rect 13403 28169 13415 28172
rect 13357 28163 13415 28169
rect 13722 28160 13728 28172
rect 13780 28160 13786 28212
rect 15286 28160 15292 28212
rect 15344 28160 15350 28212
rect 12308 28104 12756 28132
rect 12912 28104 14412 28132
rect 12308 28092 12314 28104
rect 12618 28024 12624 28076
rect 12676 28073 12682 28076
rect 12676 28027 12688 28073
rect 12728 28064 12756 28104
rect 12897 28067 12955 28073
rect 12897 28064 12909 28067
rect 12728 28036 12909 28064
rect 12897 28033 12909 28036
rect 12943 28033 12955 28067
rect 12897 28027 12955 28033
rect 12676 28024 12682 28027
rect 12986 28024 12992 28076
rect 13044 28064 13050 28076
rect 14384 28073 14412 28104
rect 15102 28092 15108 28144
rect 15160 28132 15166 28144
rect 15160 28104 15700 28132
rect 15160 28092 15166 28104
rect 14369 28067 14427 28073
rect 13044 28036 13584 28064
rect 13044 28024 13050 28036
rect 13078 27956 13084 28008
rect 13136 27996 13142 28008
rect 13556 28005 13584 28036
rect 14369 28033 14381 28067
rect 14415 28033 14427 28067
rect 14369 28027 14427 28033
rect 15562 28024 15568 28076
rect 15620 28024 15626 28076
rect 15672 28073 15700 28104
rect 15657 28067 15715 28073
rect 15657 28033 15669 28067
rect 15703 28033 15715 28067
rect 15657 28027 15715 28033
rect 15746 28024 15752 28076
rect 15804 28024 15810 28076
rect 15838 28024 15844 28076
rect 15896 28064 15902 28076
rect 15933 28067 15991 28073
rect 15933 28064 15945 28067
rect 15896 28036 15945 28064
rect 15896 28024 15902 28036
rect 15933 28033 15945 28036
rect 15979 28033 15991 28067
rect 15933 28027 15991 28033
rect 16025 28067 16083 28073
rect 16025 28033 16037 28067
rect 16071 28064 16083 28067
rect 16114 28064 16120 28076
rect 16071 28036 16120 28064
rect 16071 28033 16083 28036
rect 16025 28027 16083 28033
rect 16114 28024 16120 28036
rect 16172 28064 16178 28076
rect 16298 28064 16304 28076
rect 16172 28036 16304 28064
rect 16172 28024 16178 28036
rect 16298 28024 16304 28036
rect 16356 28024 16362 28076
rect 13449 27999 13507 28005
rect 13449 27996 13461 27999
rect 13136 27968 13461 27996
rect 13136 27956 13142 27968
rect 13449 27965 13461 27968
rect 13495 27965 13507 27999
rect 13449 27959 13507 27965
rect 13541 27999 13599 28005
rect 13541 27965 13553 27999
rect 13587 27965 13599 27999
rect 13541 27959 13599 27965
rect 15105 27999 15163 28005
rect 15105 27965 15117 27999
rect 15151 27965 15163 27999
rect 15580 27996 15608 28024
rect 15580 27968 15792 27996
rect 15105 27959 15163 27965
rect 15120 27928 15148 27959
rect 15764 27940 15792 27968
rect 13464 27900 15148 27928
rect 13464 27860 13492 27900
rect 15746 27888 15752 27940
rect 15804 27888 15810 27940
rect 11532 27832 13492 27860
rect 13538 27820 13544 27872
rect 13596 27860 13602 27872
rect 13817 27863 13875 27869
rect 13817 27860 13829 27863
rect 13596 27832 13829 27860
rect 13596 27820 13602 27832
rect 13817 27829 13829 27832
rect 13863 27829 13875 27863
rect 13817 27823 13875 27829
rect 14550 27820 14556 27872
rect 14608 27820 14614 27872
rect 16206 27820 16212 27872
rect 16264 27820 16270 27872
rect 1104 27770 16652 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 16652 27770
rect 1104 27696 16652 27718
rect 7006 27616 7012 27668
rect 7064 27656 7070 27668
rect 7374 27656 7380 27668
rect 7064 27628 7380 27656
rect 7064 27616 7070 27628
rect 7374 27616 7380 27628
rect 7432 27616 7438 27668
rect 10965 27659 11023 27665
rect 10965 27625 10977 27659
rect 11011 27656 11023 27659
rect 11606 27656 11612 27668
rect 11011 27628 11612 27656
rect 11011 27625 11023 27628
rect 10965 27619 11023 27625
rect 11606 27616 11612 27628
rect 11664 27616 11670 27668
rect 12250 27616 12256 27668
rect 12308 27656 12314 27668
rect 12308 27628 12480 27656
rect 12308 27616 12314 27628
rect 7098 27548 7104 27600
rect 7156 27588 7162 27600
rect 7834 27588 7840 27600
rect 7156 27560 7840 27588
rect 7156 27548 7162 27560
rect 7834 27548 7840 27560
rect 7892 27548 7898 27600
rect 8938 27548 8944 27600
rect 8996 27548 9002 27600
rect 12345 27591 12403 27597
rect 12345 27588 12357 27591
rect 11072 27560 12357 27588
rect 4065 27523 4123 27529
rect 4065 27520 4077 27523
rect 3712 27492 4077 27520
rect 2041 27455 2099 27461
rect 2041 27421 2053 27455
rect 2087 27452 2099 27455
rect 2774 27452 2780 27464
rect 2087 27424 2780 27452
rect 2087 27421 2099 27424
rect 2041 27415 2099 27421
rect 2774 27412 2780 27424
rect 2832 27452 2838 27464
rect 3712 27452 3740 27492
rect 4065 27489 4077 27492
rect 4111 27520 4123 27523
rect 7852 27520 7880 27548
rect 4111 27492 4200 27520
rect 7852 27492 9168 27520
rect 4111 27489 4123 27492
rect 4065 27483 4123 27489
rect 4172 27464 4200 27492
rect 2832 27424 3740 27452
rect 2832 27412 2838 27424
rect 3786 27412 3792 27464
rect 3844 27412 3850 27464
rect 3973 27455 4031 27461
rect 3973 27421 3985 27455
rect 4019 27452 4031 27455
rect 4019 27424 4108 27452
rect 4019 27421 4031 27424
rect 3973 27415 4031 27421
rect 4080 27396 4108 27424
rect 4154 27412 4160 27464
rect 4212 27412 4218 27464
rect 5537 27455 5595 27461
rect 5537 27421 5549 27455
rect 5583 27452 5595 27455
rect 5626 27452 5632 27464
rect 5583 27424 5632 27452
rect 5583 27421 5595 27424
rect 5537 27415 5595 27421
rect 5626 27412 5632 27424
rect 5684 27412 5690 27464
rect 7561 27455 7619 27461
rect 7561 27452 7573 27455
rect 6932 27424 7573 27452
rect 2308 27387 2366 27393
rect 2308 27353 2320 27387
rect 2354 27384 2366 27387
rect 2406 27384 2412 27396
rect 2354 27356 2412 27384
rect 2354 27353 2366 27356
rect 2308 27347 2366 27353
rect 2406 27344 2412 27356
rect 2464 27344 2470 27396
rect 4062 27344 4068 27396
rect 4120 27344 4126 27396
rect 4332 27387 4390 27393
rect 4332 27353 4344 27387
rect 4378 27384 4390 27387
rect 4614 27384 4620 27396
rect 4378 27356 4620 27384
rect 4378 27353 4390 27356
rect 4332 27347 4390 27353
rect 4614 27344 4620 27356
rect 4672 27344 4678 27396
rect 5804 27387 5862 27393
rect 5804 27353 5816 27387
rect 5850 27384 5862 27387
rect 5994 27384 6000 27396
rect 5850 27356 6000 27384
rect 5850 27353 5862 27356
rect 5804 27347 5862 27353
rect 5994 27344 6000 27356
rect 6052 27344 6058 27396
rect 3326 27276 3332 27328
rect 3384 27316 3390 27328
rect 3421 27319 3479 27325
rect 3421 27316 3433 27319
rect 3384 27288 3433 27316
rect 3384 27276 3390 27288
rect 3421 27285 3433 27288
rect 3467 27285 3479 27319
rect 3421 27279 3479 27285
rect 3878 27276 3884 27328
rect 3936 27276 3942 27328
rect 5258 27276 5264 27328
rect 5316 27316 5322 27328
rect 5445 27319 5503 27325
rect 5445 27316 5457 27319
rect 5316 27288 5457 27316
rect 5316 27276 5322 27288
rect 5445 27285 5457 27288
rect 5491 27285 5503 27319
rect 5445 27279 5503 27285
rect 6270 27276 6276 27328
rect 6328 27316 6334 27328
rect 6730 27316 6736 27328
rect 6328 27288 6736 27316
rect 6328 27276 6334 27288
rect 6730 27276 6736 27288
rect 6788 27316 6794 27328
rect 6932 27325 6960 27424
rect 7561 27421 7573 27424
rect 7607 27421 7619 27455
rect 7561 27415 7619 27421
rect 8754 27412 8760 27464
rect 8812 27412 8818 27464
rect 9140 27461 9168 27492
rect 8941 27455 8999 27461
rect 8941 27421 8953 27455
rect 8987 27421 8999 27455
rect 8941 27415 8999 27421
rect 9125 27455 9183 27461
rect 9125 27421 9137 27455
rect 9171 27421 9183 27455
rect 9125 27415 9183 27421
rect 9585 27455 9643 27461
rect 9585 27421 9597 27455
rect 9631 27452 9643 27455
rect 9674 27452 9680 27464
rect 9631 27424 9680 27452
rect 9631 27421 9643 27424
rect 9585 27415 9643 27421
rect 7282 27344 7288 27396
rect 7340 27384 7346 27396
rect 8956 27384 8984 27415
rect 9674 27412 9680 27424
rect 9732 27412 9738 27464
rect 9852 27455 9910 27461
rect 9852 27421 9864 27455
rect 9898 27452 9910 27455
rect 11072 27452 11100 27560
rect 12345 27557 12357 27560
rect 12391 27557 12403 27591
rect 12452 27588 12480 27628
rect 14274 27616 14280 27668
rect 14332 27656 14338 27668
rect 14826 27656 14832 27668
rect 14332 27628 14832 27656
rect 14332 27616 14338 27628
rect 14826 27616 14832 27628
rect 14884 27656 14890 27668
rect 14884 27628 15148 27656
rect 14884 27616 14890 27628
rect 12452 27560 12940 27588
rect 12345 27551 12403 27557
rect 11146 27480 11152 27532
rect 11204 27520 11210 27532
rect 11609 27523 11667 27529
rect 11609 27520 11621 27523
rect 11204 27492 11621 27520
rect 11204 27480 11210 27492
rect 11609 27489 11621 27492
rect 11655 27489 11667 27523
rect 11882 27520 11888 27532
rect 11609 27483 11667 27489
rect 11716 27492 11888 27520
rect 9898 27424 11100 27452
rect 9898 27421 9910 27424
rect 9852 27415 9910 27421
rect 7340 27356 8984 27384
rect 7340 27344 7346 27356
rect 10594 27344 10600 27396
rect 10652 27384 10658 27396
rect 11164 27384 11192 27480
rect 11425 27455 11483 27461
rect 11425 27421 11437 27455
rect 11471 27452 11483 27455
rect 11716 27452 11744 27492
rect 11882 27480 11888 27492
rect 11940 27480 11946 27532
rect 12802 27480 12808 27532
rect 12860 27480 12866 27532
rect 12912 27529 12940 27560
rect 12897 27523 12955 27529
rect 12897 27489 12909 27523
rect 12943 27489 12955 27523
rect 12897 27483 12955 27489
rect 13446 27480 13452 27532
rect 13504 27520 13510 27532
rect 13725 27523 13783 27529
rect 13725 27520 13737 27523
rect 13504 27492 13737 27520
rect 13504 27480 13510 27492
rect 13725 27489 13737 27492
rect 13771 27489 13783 27523
rect 15120 27520 15148 27628
rect 15120 27492 16252 27520
rect 13725 27483 13783 27489
rect 11471 27424 11744 27452
rect 11793 27455 11851 27461
rect 11471 27421 11483 27424
rect 11425 27415 11483 27421
rect 11793 27421 11805 27455
rect 11839 27452 11851 27455
rect 12986 27452 12992 27464
rect 11839 27424 12992 27452
rect 11839 27421 11851 27424
rect 11793 27415 11851 27421
rect 12986 27412 12992 27424
rect 13044 27412 13050 27464
rect 13538 27412 13544 27464
rect 13596 27412 13602 27464
rect 14093 27455 14151 27461
rect 14093 27421 14105 27455
rect 14139 27452 14151 27455
rect 14918 27452 14924 27464
rect 14139 27424 14924 27452
rect 14139 27421 14151 27424
rect 14093 27415 14151 27421
rect 14918 27412 14924 27424
rect 14976 27412 14982 27464
rect 15746 27412 15752 27464
rect 15804 27452 15810 27464
rect 15841 27455 15899 27461
rect 15841 27452 15853 27455
rect 15804 27424 15853 27452
rect 15804 27412 15810 27424
rect 15841 27421 15853 27424
rect 15887 27421 15899 27455
rect 15841 27415 15899 27421
rect 15933 27455 15991 27461
rect 15933 27421 15945 27455
rect 15979 27421 15991 27455
rect 15933 27415 15991 27421
rect 12713 27387 12771 27393
rect 12713 27384 12725 27387
rect 10652 27356 11192 27384
rect 12268 27356 12725 27384
rect 10652 27344 10658 27356
rect 6917 27319 6975 27325
rect 6917 27316 6929 27319
rect 6788 27288 6929 27316
rect 6788 27276 6794 27288
rect 6917 27285 6929 27288
rect 6963 27285 6975 27319
rect 6917 27279 6975 27285
rect 7006 27276 7012 27328
rect 7064 27276 7070 27328
rect 8113 27319 8171 27325
rect 8113 27285 8125 27319
rect 8159 27316 8171 27319
rect 8478 27316 8484 27328
rect 8159 27288 8484 27316
rect 8159 27285 8171 27288
rect 8113 27279 8171 27285
rect 8478 27276 8484 27288
rect 8536 27276 8542 27328
rect 11238 27276 11244 27328
rect 11296 27276 11302 27328
rect 11882 27276 11888 27328
rect 11940 27276 11946 27328
rect 12268 27325 12296 27356
rect 12713 27353 12725 27356
rect 12759 27353 12771 27387
rect 12713 27347 12771 27353
rect 14360 27387 14418 27393
rect 14360 27353 14372 27387
rect 14406 27384 14418 27387
rect 14734 27384 14740 27396
rect 14406 27356 14740 27384
rect 14406 27353 14418 27356
rect 14360 27347 14418 27353
rect 14734 27344 14740 27356
rect 14792 27344 14798 27396
rect 15378 27344 15384 27396
rect 15436 27384 15442 27396
rect 15654 27384 15660 27396
rect 15436 27356 15660 27384
rect 15436 27344 15442 27356
rect 15654 27344 15660 27356
rect 15712 27384 15718 27396
rect 15948 27384 15976 27415
rect 16022 27412 16028 27464
rect 16080 27412 16086 27464
rect 16114 27412 16120 27464
rect 16172 27452 16178 27464
rect 16224 27461 16252 27492
rect 16209 27455 16267 27461
rect 16209 27452 16221 27455
rect 16172 27424 16221 27452
rect 16172 27412 16178 27424
rect 16209 27421 16221 27424
rect 16255 27421 16267 27455
rect 16209 27415 16267 27421
rect 15712 27356 15976 27384
rect 15712 27344 15718 27356
rect 12253 27319 12311 27325
rect 12253 27285 12265 27319
rect 12299 27285 12311 27319
rect 12253 27279 12311 27285
rect 13170 27276 13176 27328
rect 13228 27276 13234 27328
rect 13633 27319 13691 27325
rect 13633 27285 13645 27319
rect 13679 27316 13691 27319
rect 15102 27316 15108 27328
rect 13679 27288 15108 27316
rect 13679 27285 13691 27288
rect 13633 27279 13691 27285
rect 15102 27276 15108 27288
rect 15160 27276 15166 27328
rect 15286 27276 15292 27328
rect 15344 27316 15350 27328
rect 15470 27316 15476 27328
rect 15344 27288 15476 27316
rect 15344 27276 15350 27288
rect 15470 27276 15476 27288
rect 15528 27276 15534 27328
rect 15562 27276 15568 27328
rect 15620 27276 15626 27328
rect 1104 27226 16652 27248
rect 1104 27174 4874 27226
rect 4926 27174 4938 27226
rect 4990 27174 5002 27226
rect 5054 27174 5066 27226
rect 5118 27174 5130 27226
rect 5182 27174 16652 27226
rect 1104 27152 16652 27174
rect 2130 27072 2136 27124
rect 2188 27112 2194 27124
rect 2866 27112 2872 27124
rect 2188 27084 2452 27112
rect 2188 27072 2194 27084
rect 1581 27047 1639 27053
rect 1581 27013 1593 27047
rect 1627 27044 1639 27047
rect 2314 27044 2320 27056
rect 1627 27016 2320 27044
rect 1627 27013 1639 27016
rect 1581 27007 1639 27013
rect 2314 27004 2320 27016
rect 2372 27004 2378 27056
rect 2424 27044 2452 27084
rect 2700 27084 2872 27112
rect 2700 27044 2728 27084
rect 2866 27072 2872 27084
rect 2924 27072 2930 27124
rect 3878 27112 3884 27124
rect 3160 27084 3884 27112
rect 2424 27016 2728 27044
rect 2774 27004 2780 27056
rect 2832 27004 2838 27056
rect 2986 27047 3044 27053
rect 2986 27013 2998 27047
rect 3032 27044 3044 27047
rect 3160 27044 3188 27084
rect 3878 27072 3884 27084
rect 3936 27072 3942 27124
rect 4617 27115 4675 27121
rect 4617 27081 4629 27115
rect 4663 27112 4675 27115
rect 4706 27112 4712 27124
rect 4663 27084 4712 27112
rect 4663 27081 4675 27084
rect 4617 27075 4675 27081
rect 4706 27072 4712 27084
rect 4764 27072 4770 27124
rect 7745 27115 7803 27121
rect 7745 27081 7757 27115
rect 7791 27112 7803 27115
rect 8202 27112 8208 27124
rect 7791 27084 8208 27112
rect 7791 27081 7803 27084
rect 7745 27075 7803 27081
rect 8202 27072 8208 27084
rect 8260 27072 8266 27124
rect 8754 27072 8760 27124
rect 8812 27112 8818 27124
rect 9401 27115 9459 27121
rect 9401 27112 9413 27115
rect 8812 27084 9413 27112
rect 8812 27072 8818 27084
rect 9401 27081 9413 27084
rect 9447 27081 9459 27115
rect 9401 27075 9459 27081
rect 10226 27072 10232 27124
rect 10284 27112 10290 27124
rect 12250 27112 12256 27124
rect 10284 27084 12256 27112
rect 10284 27072 10290 27084
rect 12250 27072 12256 27084
rect 12308 27072 12314 27124
rect 12529 27115 12587 27121
rect 12529 27081 12541 27115
rect 12575 27112 12587 27115
rect 12618 27112 12624 27124
rect 12575 27084 12624 27112
rect 12575 27081 12587 27084
rect 12529 27075 12587 27081
rect 12618 27072 12624 27084
rect 12676 27072 12682 27124
rect 12897 27115 12955 27121
rect 12897 27081 12909 27115
rect 12943 27112 12955 27115
rect 14550 27112 14556 27124
rect 12943 27084 14556 27112
rect 12943 27081 12955 27084
rect 12897 27075 12955 27081
rect 14550 27072 14556 27084
rect 14608 27072 14614 27124
rect 4154 27044 4160 27056
rect 3032 27016 3188 27044
rect 3343 27016 4160 27044
rect 3032 27013 3044 27016
rect 2986 27007 3044 27013
rect 1489 26979 1547 26985
rect 1489 26945 1501 26979
rect 1535 26945 1547 26979
rect 1489 26939 1547 26945
rect 1504 26840 1532 26939
rect 1670 26936 1676 26988
rect 1728 26936 1734 26988
rect 1765 26979 1823 26985
rect 1765 26945 1777 26979
rect 1811 26976 1823 26979
rect 3226 26979 3284 26985
rect 1811 26948 2544 26976
rect 1811 26945 1823 26948
rect 1765 26939 1823 26945
rect 2038 26868 2044 26920
rect 2096 26868 2102 26920
rect 2222 26868 2228 26920
rect 2280 26917 2286 26920
rect 2516 26917 2544 26948
rect 3226 26945 3238 26979
rect 3272 26976 3284 26979
rect 3343 26976 3371 27016
rect 4154 27004 4160 27016
rect 4212 27004 4218 27056
rect 7098 27044 7104 27056
rect 6380 27016 7104 27044
rect 3510 26985 3516 26988
rect 3504 26976 3516 26985
rect 3272 26948 3371 26976
rect 3471 26948 3516 26976
rect 3272 26945 3284 26948
rect 3226 26939 3284 26945
rect 3504 26939 3516 26948
rect 3510 26936 3516 26939
rect 3568 26936 3574 26988
rect 4982 26985 4988 26988
rect 4976 26939 4988 26985
rect 4982 26936 4988 26939
rect 5040 26936 5046 26988
rect 6380 26985 6408 27016
rect 7098 27004 7104 27016
rect 7156 27044 7162 27056
rect 7926 27044 7932 27056
rect 7156 27016 7932 27044
rect 7156 27004 7162 27016
rect 7926 27004 7932 27016
rect 7984 27044 7990 27056
rect 7984 27016 8064 27044
rect 7984 27004 7990 27016
rect 6365 26979 6423 26985
rect 6365 26945 6377 26979
rect 6411 26945 6423 26979
rect 6365 26939 6423 26945
rect 6632 26979 6690 26985
rect 6632 26945 6644 26979
rect 6678 26976 6690 26979
rect 6914 26976 6920 26988
rect 6678 26948 6920 26976
rect 6678 26945 6690 26948
rect 6632 26939 6690 26945
rect 6914 26936 6920 26948
rect 6972 26936 6978 26988
rect 8036 26985 8064 27016
rect 9674 27004 9680 27056
rect 9732 27044 9738 27056
rect 11609 27047 11667 27053
rect 11609 27044 11621 27047
rect 9732 27016 11621 27044
rect 9732 27004 9738 27016
rect 11609 27013 11621 27016
rect 11655 27013 11667 27047
rect 11609 27007 11667 27013
rect 12437 27047 12495 27053
rect 12437 27013 12449 27047
rect 12483 27044 12495 27047
rect 13262 27044 13268 27056
rect 12483 27016 13268 27044
rect 12483 27013 12495 27016
rect 12437 27007 12495 27013
rect 13262 27004 13268 27016
rect 13320 27004 13326 27056
rect 15188 27047 15246 27053
rect 15188 27013 15200 27047
rect 15234 27044 15246 27047
rect 15562 27044 15568 27056
rect 15234 27016 15568 27044
rect 15234 27013 15246 27016
rect 15188 27007 15246 27013
rect 15562 27004 15568 27016
rect 15620 27004 15626 27056
rect 8021 26979 8079 26985
rect 8021 26945 8033 26979
rect 8067 26945 8079 26979
rect 8021 26939 8079 26945
rect 8110 26936 8116 26988
rect 8168 26976 8174 26988
rect 8277 26979 8335 26985
rect 8277 26976 8289 26979
rect 8168 26948 8289 26976
rect 8168 26936 8174 26948
rect 8277 26945 8289 26948
rect 8323 26945 8335 26979
rect 8277 26939 8335 26945
rect 9953 26979 10011 26985
rect 9953 26945 9965 26979
rect 9999 26945 10011 26979
rect 9953 26939 10011 26945
rect 10045 26979 10103 26985
rect 10045 26945 10057 26979
rect 10091 26976 10103 26979
rect 10413 26979 10471 26985
rect 10413 26976 10425 26979
rect 10091 26948 10425 26976
rect 10091 26945 10103 26948
rect 10045 26939 10103 26945
rect 10413 26945 10425 26948
rect 10459 26945 10471 26979
rect 10413 26939 10471 26945
rect 12989 26979 13047 26985
rect 12989 26945 13001 26979
rect 13035 26976 13047 26979
rect 13354 26976 13360 26988
rect 13035 26948 13360 26976
rect 13035 26945 13047 26948
rect 12989 26939 13047 26945
rect 2280 26911 2308 26917
rect 2296 26877 2308 26911
rect 2280 26871 2308 26877
rect 2501 26911 2559 26917
rect 2501 26877 2513 26911
rect 2547 26908 2559 26911
rect 2958 26908 2964 26920
rect 2547 26880 2964 26908
rect 2547 26877 2559 26880
rect 2501 26871 2559 26877
rect 2280 26868 2286 26871
rect 2958 26868 2964 26880
rect 3016 26868 3022 26920
rect 4709 26911 4767 26917
rect 4709 26877 4721 26911
rect 4755 26877 4767 26911
rect 4709 26871 4767 26877
rect 1504 26812 2084 26840
rect 2056 26772 2084 26812
rect 2406 26800 2412 26852
rect 2464 26800 2470 26852
rect 3050 26800 3056 26852
rect 3108 26840 3114 26852
rect 3145 26843 3203 26849
rect 3145 26840 3157 26843
rect 3108 26812 3157 26840
rect 3108 26800 3114 26812
rect 3145 26809 3157 26812
rect 3191 26809 3203 26843
rect 3145 26803 3203 26809
rect 3418 26772 3424 26784
rect 2056 26744 3424 26772
rect 3418 26732 3424 26744
rect 3476 26732 3482 26784
rect 4154 26732 4160 26784
rect 4212 26772 4218 26784
rect 4724 26772 4752 26871
rect 9968 26840 9996 26939
rect 13354 26936 13360 26948
rect 13412 26936 13418 26988
rect 14573 26979 14631 26985
rect 14573 26945 14585 26979
rect 14619 26976 14631 26979
rect 14734 26976 14740 26988
rect 14619 26948 14740 26976
rect 14619 26945 14631 26948
rect 14573 26939 14631 26945
rect 14734 26936 14740 26948
rect 14792 26936 14798 26988
rect 14829 26979 14887 26985
rect 14829 26945 14841 26979
rect 14875 26976 14887 26979
rect 14918 26976 14924 26988
rect 14875 26948 14924 26976
rect 14875 26945 14887 26948
rect 14829 26939 14887 26945
rect 14918 26936 14924 26948
rect 14976 26936 14982 26988
rect 10226 26868 10232 26920
rect 10284 26868 10290 26920
rect 10318 26868 10324 26920
rect 10376 26908 10382 26920
rect 10965 26911 11023 26917
rect 10965 26908 10977 26911
rect 10376 26880 10977 26908
rect 10376 26868 10382 26880
rect 10965 26877 10977 26880
rect 11011 26877 11023 26911
rect 10965 26871 11023 26877
rect 12618 26868 12624 26920
rect 12676 26908 12682 26920
rect 13081 26911 13139 26917
rect 13081 26908 13093 26911
rect 12676 26880 13093 26908
rect 12676 26868 12682 26880
rect 13081 26877 13093 26880
rect 13127 26877 13139 26911
rect 13081 26871 13139 26877
rect 8956 26812 9996 26840
rect 5626 26772 5632 26784
rect 4212 26744 5632 26772
rect 4212 26732 4218 26744
rect 5626 26732 5632 26744
rect 5684 26732 5690 26784
rect 6086 26732 6092 26784
rect 6144 26732 6150 26784
rect 7466 26732 7472 26784
rect 7524 26772 7530 26784
rect 8956 26772 8984 26812
rect 11238 26800 11244 26852
rect 11296 26840 11302 26852
rect 11296 26812 13952 26840
rect 11296 26800 11302 26812
rect 7524 26744 8984 26772
rect 7524 26732 7530 26744
rect 9582 26732 9588 26784
rect 9640 26732 9646 26784
rect 13446 26732 13452 26784
rect 13504 26732 13510 26784
rect 13924 26772 13952 26812
rect 15286 26772 15292 26784
rect 13924 26744 15292 26772
rect 15286 26732 15292 26744
rect 15344 26732 15350 26784
rect 16298 26732 16304 26784
rect 16356 26732 16362 26784
rect 1104 26682 16652 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 16652 26682
rect 1104 26608 16652 26630
rect 1949 26571 2007 26577
rect 1949 26537 1961 26571
rect 1995 26568 2007 26571
rect 2222 26568 2228 26580
rect 1995 26540 2228 26568
rect 1995 26537 2007 26540
rect 1949 26531 2007 26537
rect 2222 26528 2228 26540
rect 2280 26528 2286 26580
rect 2590 26528 2596 26580
rect 2648 26528 2654 26580
rect 2774 26528 2780 26580
rect 2832 26568 2838 26580
rect 2832 26540 3740 26568
rect 2832 26528 2838 26540
rect 1670 26460 1676 26512
rect 1728 26500 1734 26512
rect 3605 26503 3663 26509
rect 3605 26500 3617 26503
rect 1728 26472 3617 26500
rect 1728 26460 1734 26472
rect 3605 26469 3617 26472
rect 3651 26469 3663 26503
rect 3712 26500 3740 26540
rect 3786 26528 3792 26580
rect 3844 26568 3850 26580
rect 6365 26571 6423 26577
rect 3844 26540 6132 26568
rect 3844 26528 3850 26540
rect 3712 26472 4384 26500
rect 3605 26463 3663 26469
rect 2406 26392 2412 26444
rect 2464 26392 2470 26444
rect 2498 26392 2504 26444
rect 2556 26432 2562 26444
rect 2752 26435 2810 26441
rect 2752 26432 2764 26435
rect 2556 26404 2764 26432
rect 2556 26392 2562 26404
rect 2752 26401 2764 26404
rect 2798 26401 2810 26435
rect 2752 26395 2810 26401
rect 2961 26435 3019 26441
rect 2961 26401 2973 26435
rect 3007 26432 3019 26435
rect 4246 26432 4252 26444
rect 3007 26404 4252 26432
rect 3007 26401 3019 26404
rect 2961 26395 3019 26401
rect 4246 26392 4252 26404
rect 4304 26392 4310 26444
rect 2317 26367 2375 26373
rect 2317 26333 2329 26367
rect 2363 26364 2375 26367
rect 2363 26336 3096 26364
rect 2363 26333 2375 26336
rect 2317 26327 2375 26333
rect 2866 26188 2872 26240
rect 2924 26188 2930 26240
rect 3068 26228 3096 26336
rect 3142 26324 3148 26376
rect 3200 26364 3206 26376
rect 3237 26367 3295 26373
rect 3237 26364 3249 26367
rect 3200 26336 3249 26364
rect 3200 26324 3206 26336
rect 3237 26333 3249 26336
rect 3283 26333 3295 26367
rect 3237 26327 3295 26333
rect 3326 26324 3332 26376
rect 3384 26324 3390 26376
rect 3605 26367 3663 26373
rect 3605 26333 3617 26367
rect 3651 26364 3663 26367
rect 3878 26364 3884 26376
rect 3651 26336 3884 26364
rect 3651 26333 3663 26336
rect 3605 26327 3663 26333
rect 3878 26324 3884 26336
rect 3936 26324 3942 26376
rect 3973 26367 4031 26373
rect 3973 26333 3985 26367
rect 4019 26364 4031 26367
rect 4356 26364 4384 26472
rect 4614 26460 4620 26512
rect 4672 26460 4678 26512
rect 5813 26503 5871 26509
rect 4724 26472 5672 26500
rect 4724 26441 4752 26472
rect 4709 26435 4767 26441
rect 4709 26401 4721 26435
rect 4755 26401 4767 26435
rect 4709 26395 4767 26401
rect 4724 26364 4752 26395
rect 4798 26392 4804 26444
rect 4856 26432 4862 26444
rect 4985 26435 5043 26441
rect 4985 26432 4997 26435
rect 4856 26404 4997 26432
rect 4856 26392 4862 26404
rect 4985 26401 4997 26404
rect 5031 26401 5043 26435
rect 4985 26395 5043 26401
rect 5074 26392 5080 26444
rect 5132 26392 5138 26444
rect 5194 26435 5252 26441
rect 5194 26401 5206 26435
rect 5240 26432 5252 26435
rect 5534 26432 5540 26444
rect 5240 26404 5540 26432
rect 5240 26401 5252 26404
rect 5194 26395 5252 26401
rect 5534 26392 5540 26404
rect 5592 26392 5598 26444
rect 4019 26336 4752 26364
rect 4019 26333 4031 26336
rect 3973 26327 4031 26333
rect 5350 26324 5356 26376
rect 5408 26364 5414 26376
rect 5445 26367 5503 26373
rect 5445 26364 5457 26367
rect 5408 26336 5457 26364
rect 5408 26324 5414 26336
rect 5445 26333 5457 26336
rect 5491 26333 5503 26367
rect 5445 26327 5503 26333
rect 3510 26256 3516 26308
rect 3568 26296 3574 26308
rect 3786 26296 3792 26308
rect 3568 26268 3792 26296
rect 3568 26256 3574 26268
rect 3786 26256 3792 26268
rect 3844 26296 3850 26308
rect 4341 26299 4399 26305
rect 4341 26296 4353 26299
rect 3844 26268 4353 26296
rect 3844 26256 3850 26268
rect 4341 26265 4353 26268
rect 4387 26265 4399 26299
rect 4341 26259 4399 26265
rect 4430 26256 4436 26308
rect 4488 26305 4494 26308
rect 4488 26299 4516 26305
rect 4504 26265 4516 26299
rect 4488 26259 4516 26265
rect 4488 26256 4494 26259
rect 4798 26256 4804 26308
rect 4856 26296 4862 26308
rect 5258 26296 5264 26308
rect 4856 26268 5264 26296
rect 4856 26256 4862 26268
rect 5258 26256 5264 26268
rect 5316 26296 5322 26308
rect 5537 26299 5595 26305
rect 5537 26296 5549 26299
rect 5316 26268 5549 26296
rect 5316 26256 5322 26268
rect 5537 26265 5549 26268
rect 5583 26265 5595 26299
rect 5644 26296 5672 26472
rect 5813 26469 5825 26503
rect 5859 26500 5871 26503
rect 5994 26500 6000 26512
rect 5859 26472 6000 26500
rect 5859 26469 5871 26472
rect 5813 26463 5871 26469
rect 5994 26460 6000 26472
rect 6052 26460 6058 26512
rect 5721 26367 5779 26373
rect 5721 26333 5733 26367
rect 5767 26364 5779 26367
rect 5994 26364 6000 26376
rect 5767 26336 6000 26364
rect 5767 26333 5779 26336
rect 5721 26327 5779 26333
rect 5994 26324 6000 26336
rect 6052 26324 6058 26376
rect 6104 26373 6132 26540
rect 6365 26537 6377 26571
rect 6411 26568 6423 26571
rect 7282 26568 7288 26580
rect 6411 26540 7288 26568
rect 6411 26537 6423 26540
rect 6365 26531 6423 26537
rect 7282 26528 7288 26540
rect 7340 26528 7346 26580
rect 8021 26571 8079 26577
rect 8021 26537 8033 26571
rect 8067 26568 8079 26571
rect 8110 26568 8116 26580
rect 8067 26540 8116 26568
rect 8067 26537 8079 26540
rect 8021 26531 8079 26537
rect 8110 26528 8116 26540
rect 8168 26528 8174 26580
rect 9306 26568 9312 26580
rect 8956 26540 9312 26568
rect 8478 26392 8484 26444
rect 8536 26392 8542 26444
rect 8665 26435 8723 26441
rect 8665 26401 8677 26435
rect 8711 26432 8723 26435
rect 8956 26432 8984 26540
rect 9306 26528 9312 26540
rect 9364 26568 9370 26580
rect 10226 26568 10232 26580
rect 9364 26540 10232 26568
rect 9364 26528 9370 26540
rect 10226 26528 10232 26540
rect 10284 26528 10290 26580
rect 10318 26528 10324 26580
rect 10376 26528 10382 26580
rect 10778 26528 10784 26580
rect 10836 26568 10842 26580
rect 14093 26571 14151 26577
rect 14093 26568 14105 26571
rect 10836 26540 14105 26568
rect 10836 26528 10842 26540
rect 14093 26537 14105 26540
rect 14139 26537 14151 26571
rect 14093 26531 14151 26537
rect 14734 26528 14740 26580
rect 14792 26568 14798 26580
rect 15565 26571 15623 26577
rect 15565 26568 15577 26571
rect 14792 26540 15577 26568
rect 14792 26528 14798 26540
rect 15565 26537 15577 26540
rect 15611 26537 15623 26571
rect 15565 26531 15623 26537
rect 11885 26503 11943 26509
rect 11885 26469 11897 26503
rect 11931 26500 11943 26503
rect 11974 26500 11980 26512
rect 11931 26472 11980 26500
rect 11931 26469 11943 26472
rect 11885 26463 11943 26469
rect 11974 26460 11980 26472
rect 12032 26460 12038 26512
rect 14550 26460 14556 26512
rect 14608 26500 14614 26512
rect 14608 26472 15976 26500
rect 14608 26460 14614 26472
rect 13630 26432 13636 26444
rect 8711 26404 8984 26432
rect 13556 26404 13636 26432
rect 8711 26401 8723 26404
rect 8665 26395 8723 26401
rect 6089 26367 6147 26373
rect 6089 26333 6101 26367
rect 6135 26333 6147 26367
rect 6089 26327 6147 26333
rect 6270 26324 6276 26376
rect 6328 26324 6334 26376
rect 6457 26367 6515 26373
rect 6457 26333 6469 26367
rect 6503 26333 6515 26367
rect 6457 26327 6515 26333
rect 6549 26367 6607 26373
rect 6549 26333 6561 26367
rect 6595 26364 6607 26367
rect 7098 26364 7104 26376
rect 6595 26336 7104 26364
rect 6595 26333 6607 26336
rect 6549 26327 6607 26333
rect 5810 26296 5816 26308
rect 5644 26268 5816 26296
rect 5537 26259 5595 26265
rect 5810 26256 5816 26268
rect 5868 26256 5874 26308
rect 6472 26296 6500 26327
rect 7098 26324 7104 26336
rect 7156 26364 7162 26376
rect 7926 26364 7932 26376
rect 7156 26336 7932 26364
rect 7156 26324 7162 26336
rect 7926 26324 7932 26336
rect 7984 26364 7990 26376
rect 8941 26367 8999 26373
rect 8941 26364 8953 26367
rect 7984 26336 8953 26364
rect 7984 26324 7990 26336
rect 8941 26333 8953 26336
rect 8987 26333 8999 26367
rect 8941 26327 8999 26333
rect 9208 26367 9266 26373
rect 9208 26333 9220 26367
rect 9254 26364 9266 26367
rect 9582 26364 9588 26376
rect 9254 26336 9588 26364
rect 9254 26333 9266 26336
rect 9208 26327 9266 26333
rect 9582 26324 9588 26336
rect 9640 26324 9646 26376
rect 9674 26324 9680 26376
rect 9732 26364 9738 26376
rect 10413 26367 10471 26373
rect 10413 26364 10425 26367
rect 9732 26336 10425 26364
rect 9732 26324 9738 26336
rect 10413 26333 10425 26336
rect 10459 26333 10471 26367
rect 10413 26327 10471 26333
rect 13009 26367 13067 26373
rect 13009 26333 13021 26367
rect 13055 26364 13067 26367
rect 13170 26364 13176 26376
rect 13055 26336 13176 26364
rect 13055 26333 13067 26336
rect 13009 26327 13067 26333
rect 13170 26324 13176 26336
rect 13228 26324 13234 26376
rect 13265 26367 13323 26373
rect 13265 26333 13277 26367
rect 13311 26364 13323 26367
rect 13311 26336 13400 26364
rect 13311 26333 13323 26336
rect 13265 26327 13323 26333
rect 6816 26299 6874 26305
rect 6472 26268 6776 26296
rect 3234 26228 3240 26240
rect 3068 26200 3240 26228
rect 3234 26188 3240 26200
rect 3292 26228 3298 26240
rect 3421 26231 3479 26237
rect 3421 26228 3433 26231
rect 3292 26200 3433 26228
rect 3292 26188 3298 26200
rect 3421 26197 3433 26200
rect 3467 26197 3479 26231
rect 3421 26191 3479 26197
rect 4246 26188 4252 26240
rect 4304 26228 4310 26240
rect 4614 26228 4620 26240
rect 4304 26200 4620 26228
rect 4304 26188 4310 26200
rect 4614 26188 4620 26200
rect 4672 26188 4678 26240
rect 4982 26188 4988 26240
rect 5040 26228 5046 26240
rect 5353 26231 5411 26237
rect 5353 26228 5365 26231
rect 5040 26200 5365 26228
rect 5040 26188 5046 26200
rect 5353 26197 5365 26200
rect 5399 26197 5411 26231
rect 5353 26191 5411 26197
rect 5622 26231 5680 26237
rect 5622 26197 5634 26231
rect 5668 26228 5680 26231
rect 5718 26228 5724 26240
rect 5668 26200 5724 26228
rect 5668 26197 5680 26200
rect 5622 26191 5680 26197
rect 5718 26188 5724 26200
rect 5776 26188 5782 26240
rect 5902 26188 5908 26240
rect 5960 26228 5966 26240
rect 5997 26231 6055 26237
rect 5997 26228 6009 26231
rect 5960 26200 6009 26228
rect 5960 26188 5966 26200
rect 5997 26197 6009 26200
rect 6043 26197 6055 26231
rect 6748 26228 6776 26268
rect 6816 26265 6828 26299
rect 6862 26296 6874 26299
rect 6914 26296 6920 26308
rect 6862 26268 6920 26296
rect 6862 26265 6874 26268
rect 6816 26259 6874 26265
rect 6914 26256 6920 26268
rect 6972 26256 6978 26308
rect 8389 26299 8447 26305
rect 8389 26265 8401 26299
rect 8435 26296 8447 26299
rect 9766 26296 9772 26308
rect 8435 26268 9772 26296
rect 8435 26265 8447 26268
rect 8389 26259 8447 26265
rect 9766 26256 9772 26268
rect 9824 26256 9830 26308
rect 10686 26305 10692 26308
rect 10680 26259 10692 26305
rect 10686 26256 10692 26259
rect 10744 26256 10750 26308
rect 13372 26240 13400 26336
rect 13556 26305 13584 26404
rect 13630 26392 13636 26404
rect 13688 26392 13694 26444
rect 13909 26435 13967 26441
rect 13909 26401 13921 26435
rect 13955 26432 13967 26435
rect 13955 26404 15516 26432
rect 13955 26401 13967 26404
rect 13909 26395 13967 26401
rect 13814 26324 13820 26376
rect 13872 26364 13878 26376
rect 14645 26367 14703 26373
rect 14645 26364 14657 26367
rect 13872 26336 14657 26364
rect 13872 26324 13878 26336
rect 14645 26333 14657 26336
rect 14691 26333 14703 26367
rect 14645 26327 14703 26333
rect 15381 26367 15439 26373
rect 15381 26333 15393 26367
rect 15427 26333 15439 26367
rect 15381 26327 15439 26333
rect 13541 26299 13599 26305
rect 13541 26265 13553 26299
rect 13587 26265 13599 26299
rect 13541 26259 13599 26265
rect 13725 26299 13783 26305
rect 13725 26265 13737 26299
rect 13771 26265 13783 26299
rect 13725 26259 13783 26265
rect 7650 26228 7656 26240
rect 6748 26200 7656 26228
rect 5997 26191 6055 26197
rect 7650 26188 7656 26200
rect 7708 26188 7714 26240
rect 7834 26188 7840 26240
rect 7892 26228 7898 26240
rect 7929 26231 7987 26237
rect 7929 26228 7941 26231
rect 7892 26200 7941 26228
rect 7892 26188 7898 26200
rect 7929 26197 7941 26200
rect 7975 26197 7987 26231
rect 7929 26191 7987 26197
rect 11790 26188 11796 26240
rect 11848 26188 11854 26240
rect 13354 26188 13360 26240
rect 13412 26188 13418 26240
rect 13446 26188 13452 26240
rect 13504 26228 13510 26240
rect 13740 26228 13768 26259
rect 13906 26256 13912 26308
rect 13964 26296 13970 26308
rect 15396 26296 15424 26327
rect 13964 26268 15424 26296
rect 15488 26296 15516 26404
rect 15838 26324 15844 26376
rect 15896 26324 15902 26376
rect 15948 26373 15976 26472
rect 15933 26367 15991 26373
rect 15933 26333 15945 26367
rect 15979 26333 15991 26367
rect 15933 26327 15991 26333
rect 16025 26367 16083 26373
rect 16025 26333 16037 26367
rect 16071 26333 16083 26367
rect 16025 26327 16083 26333
rect 16040 26296 16068 26327
rect 16114 26324 16120 26376
rect 16172 26364 16178 26376
rect 16209 26367 16267 26373
rect 16209 26364 16221 26367
rect 16172 26336 16221 26364
rect 16172 26324 16178 26336
rect 16209 26333 16221 26336
rect 16255 26333 16267 26367
rect 16209 26327 16267 26333
rect 15488 26268 16068 26296
rect 13964 26256 13970 26268
rect 13504 26200 13768 26228
rect 13504 26188 13510 26200
rect 14826 26188 14832 26240
rect 14884 26188 14890 26240
rect 1104 26138 16652 26160
rect 1104 26086 4874 26138
rect 4926 26086 4938 26138
rect 4990 26086 5002 26138
rect 5054 26086 5066 26138
rect 5118 26086 5130 26138
rect 5182 26086 16652 26138
rect 1104 26064 16652 26086
rect 3970 26024 3976 26036
rect 3528 25996 3976 26024
rect 2406 25916 2412 25968
rect 2464 25956 2470 25968
rect 3142 25956 3148 25968
rect 2464 25928 3148 25956
rect 2464 25916 2470 25928
rect 3142 25916 3148 25928
rect 3200 25956 3206 25968
rect 3326 25965 3332 25968
rect 3297 25959 3332 25965
rect 3297 25956 3309 25959
rect 3200 25928 3309 25956
rect 3200 25916 3206 25928
rect 3297 25925 3309 25928
rect 3297 25919 3332 25925
rect 3326 25916 3332 25919
rect 3384 25916 3390 25968
rect 3528 25965 3556 25996
rect 3970 25984 3976 25996
rect 4028 25984 4034 26036
rect 5350 25984 5356 26036
rect 5408 26033 5414 26036
rect 5408 26027 5432 26033
rect 5420 25993 5432 26027
rect 5408 25987 5432 25993
rect 5408 25984 5414 25987
rect 5534 25984 5540 26036
rect 5592 26024 5598 26036
rect 5721 26027 5779 26033
rect 5721 26024 5733 26027
rect 5592 25996 5733 26024
rect 5592 25984 5598 25996
rect 5721 25993 5733 25996
rect 5767 25993 5779 26027
rect 5721 25987 5779 25993
rect 6914 25984 6920 26036
rect 6972 26024 6978 26036
rect 7101 26027 7159 26033
rect 7101 26024 7113 26027
rect 6972 25996 7113 26024
rect 6972 25984 6978 25996
rect 7101 25993 7113 25996
rect 7147 25993 7159 26027
rect 7101 25987 7159 25993
rect 9214 25984 9220 26036
rect 9272 26024 9278 26036
rect 9585 26027 9643 26033
rect 9585 26024 9597 26027
rect 9272 25996 9597 26024
rect 9272 25984 9278 25996
rect 9585 25993 9597 25996
rect 9631 25993 9643 26027
rect 9585 25987 9643 25993
rect 9677 26027 9735 26033
rect 9677 25993 9689 26027
rect 9723 26024 9735 26027
rect 9766 26024 9772 26036
rect 9723 25996 9772 26024
rect 9723 25993 9735 25996
rect 9677 25987 9735 25993
rect 9766 25984 9772 25996
rect 9824 25984 9830 26036
rect 10597 26027 10655 26033
rect 10597 25993 10609 26027
rect 10643 26024 10655 26027
rect 10686 26024 10692 26036
rect 10643 25996 10692 26024
rect 10643 25993 10655 25996
rect 10597 25987 10655 25993
rect 10686 25984 10692 25996
rect 10744 25984 10750 26036
rect 10778 25984 10784 26036
rect 10836 26024 10842 26036
rect 10965 26027 11023 26033
rect 10965 26024 10977 26027
rect 10836 25996 10977 26024
rect 10836 25984 10842 25996
rect 10965 25993 10977 25996
rect 11011 25993 11023 26027
rect 14277 26027 14335 26033
rect 14277 26024 14289 26027
rect 10965 25987 11023 25993
rect 13096 25996 14289 26024
rect 3513 25959 3571 25965
rect 3513 25925 3525 25959
rect 3559 25925 3571 25959
rect 3513 25919 3571 25925
rect 4157 25959 4215 25965
rect 4157 25925 4169 25959
rect 4203 25956 4215 25959
rect 4706 25956 4712 25968
rect 4203 25928 4712 25956
rect 4203 25925 4215 25928
rect 4157 25919 4215 25925
rect 4706 25916 4712 25928
rect 4764 25916 4770 25968
rect 5169 25959 5227 25965
rect 5169 25925 5181 25959
rect 5215 25956 5227 25959
rect 6086 25956 6092 25968
rect 5215 25928 6092 25956
rect 5215 25925 5227 25928
rect 5169 25919 5227 25925
rect 6086 25916 6092 25928
rect 6144 25916 6150 25968
rect 7193 25959 7251 25965
rect 7193 25925 7205 25959
rect 7239 25956 7251 25959
rect 8202 25956 8208 25968
rect 7239 25928 8208 25956
rect 7239 25925 7251 25928
rect 7193 25919 7251 25925
rect 8202 25916 8208 25928
rect 8260 25916 8266 25968
rect 10045 25959 10103 25965
rect 10045 25925 10057 25959
rect 10091 25956 10103 25959
rect 12066 25956 12072 25968
rect 10091 25928 12072 25956
rect 10091 25925 10103 25928
rect 10045 25919 10103 25925
rect 12066 25916 12072 25928
rect 12124 25916 12130 25968
rect 12928 25959 12986 25965
rect 12928 25925 12940 25959
rect 12974 25956 12986 25959
rect 13096 25956 13124 25996
rect 14277 25993 14289 25996
rect 14323 25993 14335 26027
rect 14277 25987 14335 25993
rect 14645 26027 14703 26033
rect 14645 25993 14657 26027
rect 14691 26024 14703 26027
rect 14826 26024 14832 26036
rect 14691 25996 14832 26024
rect 14691 25993 14703 25996
rect 14645 25987 14703 25993
rect 14826 25984 14832 25996
rect 14884 25984 14890 26036
rect 15102 25984 15108 26036
rect 15160 25984 15166 26036
rect 13354 25956 13360 25968
rect 12974 25928 13124 25956
rect 13188 25928 13360 25956
rect 12974 25925 12986 25928
rect 12928 25919 12986 25925
rect 3344 25888 3372 25916
rect 3789 25891 3847 25897
rect 3789 25888 3801 25891
rect 3344 25860 3801 25888
rect 3789 25857 3801 25860
rect 3835 25857 3847 25891
rect 3789 25851 3847 25857
rect 3881 25891 3939 25897
rect 3881 25857 3893 25891
rect 3927 25857 3939 25891
rect 3881 25851 3939 25857
rect 4617 25891 4675 25897
rect 4617 25857 4629 25891
rect 4663 25888 4675 25891
rect 4798 25888 4804 25900
rect 4663 25860 4804 25888
rect 4663 25857 4675 25860
rect 4617 25851 4675 25857
rect 3896 25820 3924 25851
rect 4798 25848 4804 25860
rect 4856 25848 4862 25900
rect 5629 25891 5687 25897
rect 5629 25857 5641 25891
rect 5675 25888 5687 25891
rect 5718 25888 5724 25900
rect 5675 25860 5724 25888
rect 5675 25857 5687 25860
rect 5629 25851 5687 25857
rect 5718 25848 5724 25860
rect 5776 25848 5782 25900
rect 5810 25848 5816 25900
rect 5868 25848 5874 25900
rect 6181 25891 6239 25897
rect 6181 25857 6193 25891
rect 6227 25888 6239 25891
rect 7834 25888 7840 25900
rect 6227 25860 7840 25888
rect 6227 25857 6239 25860
rect 6181 25851 6239 25857
rect 7834 25848 7840 25860
rect 7892 25848 7898 25900
rect 7926 25848 7932 25900
rect 7984 25888 7990 25900
rect 8472 25891 8530 25897
rect 7984 25860 8248 25888
rect 7984 25848 7990 25860
rect 3528 25792 3924 25820
rect 4249 25823 4307 25829
rect 3145 25755 3203 25761
rect 3145 25721 3157 25755
rect 3191 25752 3203 25755
rect 3418 25752 3424 25764
rect 3191 25724 3424 25752
rect 3191 25721 3203 25724
rect 3145 25715 3203 25721
rect 3418 25712 3424 25724
rect 3476 25712 3482 25764
rect 3234 25644 3240 25696
rect 3292 25684 3298 25696
rect 3329 25687 3387 25693
rect 3329 25684 3341 25687
rect 3292 25656 3341 25684
rect 3292 25644 3298 25656
rect 3329 25653 3341 25656
rect 3375 25684 3387 25687
rect 3528 25684 3556 25792
rect 4249 25789 4261 25823
rect 4295 25820 4307 25823
rect 4430 25820 4436 25832
rect 4295 25792 4436 25820
rect 4295 25789 4307 25792
rect 4249 25783 4307 25789
rect 4430 25780 4436 25792
rect 4488 25780 4494 25832
rect 4709 25823 4767 25829
rect 4709 25789 4721 25823
rect 4755 25820 4767 25823
rect 5350 25820 5356 25832
rect 4755 25792 5356 25820
rect 4755 25789 4767 25792
rect 4709 25783 4767 25789
rect 3605 25755 3663 25761
rect 3605 25721 3617 25755
rect 3651 25752 3663 25755
rect 4062 25752 4068 25764
rect 3651 25724 4068 25752
rect 3651 25721 3663 25724
rect 3605 25715 3663 25721
rect 4062 25712 4068 25724
rect 4120 25752 4126 25764
rect 4724 25752 4752 25783
rect 5350 25780 5356 25792
rect 5408 25780 5414 25832
rect 6546 25780 6552 25832
rect 6604 25780 6610 25832
rect 8220 25829 8248 25860
rect 8472 25857 8484 25891
rect 8518 25888 8530 25891
rect 9030 25888 9036 25900
rect 8518 25860 9036 25888
rect 8518 25857 8530 25860
rect 8472 25851 8530 25857
rect 9030 25848 9036 25860
rect 9088 25848 9094 25900
rect 10137 25891 10195 25897
rect 10137 25857 10149 25891
rect 10183 25888 10195 25891
rect 10410 25888 10416 25900
rect 10183 25860 10416 25888
rect 10183 25857 10195 25860
rect 10137 25851 10195 25857
rect 10410 25848 10416 25860
rect 10468 25848 10474 25900
rect 11057 25891 11115 25897
rect 11057 25857 11069 25891
rect 11103 25888 11115 25891
rect 11698 25888 11704 25900
rect 11103 25860 11704 25888
rect 11103 25857 11115 25860
rect 11057 25851 11115 25857
rect 11698 25848 11704 25860
rect 11756 25848 11762 25900
rect 13188 25897 13216 25928
rect 13354 25916 13360 25928
rect 13412 25956 13418 25968
rect 14093 25959 14151 25965
rect 14093 25956 14105 25959
rect 13412 25928 14105 25956
rect 13412 25916 13418 25928
rect 14093 25925 14105 25928
rect 14139 25956 14151 25959
rect 14918 25956 14924 25968
rect 14139 25928 14924 25956
rect 14139 25925 14151 25928
rect 14093 25919 14151 25925
rect 14918 25916 14924 25928
rect 14976 25916 14982 25968
rect 16117 25959 16175 25965
rect 16117 25956 16129 25959
rect 15120 25928 15424 25956
rect 13173 25891 13231 25897
rect 13173 25857 13185 25891
rect 13219 25857 13231 25891
rect 13173 25851 13231 25857
rect 13262 25848 13268 25900
rect 13320 25848 13326 25900
rect 13446 25848 13452 25900
rect 13504 25888 13510 25900
rect 15120 25888 15148 25928
rect 13504 25860 15148 25888
rect 13504 25848 13510 25860
rect 15194 25848 15200 25900
rect 15252 25888 15258 25900
rect 15396 25897 15424 25928
rect 15856 25928 16129 25956
rect 15289 25891 15347 25897
rect 15289 25888 15301 25891
rect 15252 25860 15301 25888
rect 15252 25848 15258 25860
rect 15289 25857 15301 25860
rect 15335 25857 15347 25891
rect 15289 25851 15347 25857
rect 15381 25891 15439 25897
rect 15381 25857 15393 25891
rect 15427 25857 15439 25891
rect 15381 25851 15439 25857
rect 15562 25848 15568 25900
rect 15620 25848 15626 25900
rect 15654 25848 15660 25900
rect 15712 25848 15718 25900
rect 8205 25823 8263 25829
rect 8205 25789 8217 25823
rect 8251 25789 8263 25823
rect 8205 25783 8263 25789
rect 10226 25780 10232 25832
rect 10284 25820 10290 25832
rect 10594 25820 10600 25832
rect 10284 25792 10600 25820
rect 10284 25780 10290 25792
rect 10594 25780 10600 25792
rect 10652 25780 10658 25832
rect 11149 25823 11207 25829
rect 11149 25789 11161 25823
rect 11195 25789 11207 25823
rect 11149 25783 11207 25789
rect 4120 25724 4752 25752
rect 6089 25755 6147 25761
rect 4120 25712 4126 25724
rect 6089 25721 6101 25755
rect 6135 25752 6147 25755
rect 7190 25752 7196 25764
rect 6135 25724 7196 25752
rect 6135 25721 6147 25724
rect 6089 25715 6147 25721
rect 7190 25712 7196 25724
rect 7248 25712 7254 25764
rect 10962 25712 10968 25764
rect 11020 25752 11026 25764
rect 11164 25752 11192 25783
rect 14458 25780 14464 25832
rect 14516 25820 14522 25832
rect 14737 25823 14795 25829
rect 14737 25820 14749 25823
rect 14516 25792 14749 25820
rect 14516 25780 14522 25792
rect 14737 25789 14749 25792
rect 14783 25789 14795 25823
rect 14737 25783 14795 25789
rect 14826 25780 14832 25832
rect 14884 25780 14890 25832
rect 11020 25724 11192 25752
rect 11020 25712 11026 25724
rect 14366 25712 14372 25764
rect 14424 25752 14430 25764
rect 15749 25755 15807 25761
rect 15749 25752 15761 25755
rect 14424 25724 15761 25752
rect 14424 25712 14430 25724
rect 15749 25721 15761 25724
rect 15795 25721 15807 25755
rect 15749 25715 15807 25721
rect 15856 25696 15884 25928
rect 16117 25925 16129 25928
rect 16163 25925 16175 25959
rect 16117 25919 16175 25925
rect 15933 25891 15991 25897
rect 15933 25857 15945 25891
rect 15979 25857 15991 25891
rect 15933 25851 15991 25857
rect 15948 25820 15976 25851
rect 16206 25820 16212 25832
rect 15948 25792 16212 25820
rect 16206 25780 16212 25792
rect 16264 25780 16270 25832
rect 3375 25656 3556 25684
rect 3375 25653 3387 25656
rect 3329 25647 3387 25653
rect 4798 25644 4804 25696
rect 4856 25684 4862 25696
rect 5353 25687 5411 25693
rect 5353 25684 5365 25687
rect 4856 25656 5365 25684
rect 4856 25644 4862 25656
rect 5353 25653 5365 25656
rect 5399 25653 5411 25687
rect 5353 25647 5411 25653
rect 5537 25687 5595 25693
rect 5537 25653 5549 25687
rect 5583 25684 5595 25687
rect 5810 25684 5816 25696
rect 5583 25656 5816 25684
rect 5583 25653 5595 25656
rect 5537 25647 5595 25653
rect 5810 25644 5816 25656
rect 5868 25644 5874 25696
rect 11793 25687 11851 25693
rect 11793 25653 11805 25687
rect 11839 25684 11851 25687
rect 11882 25684 11888 25696
rect 11839 25656 11888 25684
rect 11839 25653 11851 25656
rect 11793 25647 11851 25653
rect 11882 25644 11888 25656
rect 11940 25684 11946 25696
rect 13906 25684 13912 25696
rect 11940 25656 13912 25684
rect 11940 25644 11946 25656
rect 13906 25644 13912 25656
rect 13964 25644 13970 25696
rect 14182 25644 14188 25696
rect 14240 25684 14246 25696
rect 15838 25684 15844 25696
rect 14240 25656 15844 25684
rect 14240 25644 14246 25656
rect 15838 25644 15844 25656
rect 15896 25644 15902 25696
rect 1104 25594 16652 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 16652 25594
rect 1104 25520 16652 25542
rect 6546 25440 6552 25492
rect 6604 25480 6610 25492
rect 6641 25483 6699 25489
rect 6641 25480 6653 25483
rect 6604 25452 6653 25480
rect 6604 25440 6610 25452
rect 6641 25449 6653 25452
rect 6687 25449 6699 25483
rect 6641 25443 6699 25449
rect 7006 25440 7012 25492
rect 7064 25440 7070 25492
rect 7650 25440 7656 25492
rect 7708 25440 7714 25492
rect 7834 25440 7840 25492
rect 7892 25440 7898 25492
rect 8110 25440 8116 25492
rect 8168 25440 8174 25492
rect 9030 25440 9036 25492
rect 9088 25440 9094 25492
rect 11054 25440 11060 25492
rect 11112 25440 11118 25492
rect 12618 25440 12624 25492
rect 12676 25480 12682 25492
rect 14826 25480 14832 25492
rect 12676 25452 14832 25480
rect 12676 25440 12682 25452
rect 14826 25440 14832 25452
rect 14884 25440 14890 25492
rect 6822 25412 6828 25424
rect 6748 25384 6828 25412
rect 4614 25304 4620 25356
rect 4672 25344 4678 25356
rect 6638 25344 6644 25356
rect 4672 25316 6644 25344
rect 4672 25304 4678 25316
rect 6638 25304 6644 25316
rect 6696 25304 6702 25356
rect 6748 25353 6776 25384
rect 6822 25372 6828 25384
rect 6880 25372 6886 25424
rect 8294 25412 8300 25424
rect 7668 25384 8300 25412
rect 6733 25347 6791 25353
rect 6733 25313 6745 25347
rect 6779 25313 6791 25347
rect 7668 25344 7696 25384
rect 8294 25372 8300 25384
rect 8352 25372 8358 25424
rect 8404 25384 14688 25412
rect 6733 25307 6791 25313
rect 6840 25316 7696 25344
rect 842 25236 848 25288
rect 900 25276 906 25288
rect 6840 25285 6868 25316
rect 7742 25304 7748 25356
rect 7800 25344 7806 25356
rect 7929 25347 7987 25353
rect 7929 25344 7941 25347
rect 7800 25316 7941 25344
rect 7800 25304 7806 25316
rect 7929 25313 7941 25316
rect 7975 25313 7987 25347
rect 7929 25307 7987 25313
rect 1397 25279 1455 25285
rect 1397 25276 1409 25279
rect 900 25248 1409 25276
rect 900 25236 906 25248
rect 1397 25245 1409 25248
rect 1443 25245 1455 25279
rect 1397 25239 1455 25245
rect 6825 25279 6883 25285
rect 6825 25245 6837 25279
rect 6871 25245 6883 25279
rect 6825 25239 6883 25245
rect 7101 25279 7159 25285
rect 7101 25245 7113 25279
rect 7147 25276 7159 25279
rect 7190 25276 7196 25288
rect 7147 25248 7196 25276
rect 7147 25245 7159 25248
rect 7101 25239 7159 25245
rect 7190 25236 7196 25248
rect 7248 25236 7254 25288
rect 7469 25279 7527 25285
rect 7469 25245 7481 25279
rect 7515 25276 7527 25279
rect 7834 25276 7840 25288
rect 7515 25248 7840 25276
rect 7515 25245 7527 25248
rect 7469 25239 7527 25245
rect 7834 25236 7840 25248
rect 7892 25236 7898 25288
rect 8018 25236 8024 25288
rect 8076 25236 8082 25288
rect 5626 25168 5632 25220
rect 5684 25168 5690 25220
rect 6457 25211 6515 25217
rect 6457 25177 6469 25211
rect 6503 25208 6515 25211
rect 8202 25208 8208 25220
rect 6503 25180 8208 25208
rect 6503 25177 6515 25180
rect 6457 25171 6515 25177
rect 8202 25168 8208 25180
rect 8260 25168 8266 25220
rect 1581 25143 1639 25149
rect 1581 25109 1593 25143
rect 1627 25140 1639 25143
rect 3510 25140 3516 25152
rect 1627 25112 3516 25140
rect 1627 25109 1639 25112
rect 1581 25103 1639 25109
rect 3510 25100 3516 25112
rect 3568 25100 3574 25152
rect 7926 25100 7932 25152
rect 7984 25140 7990 25152
rect 8404 25140 8432 25384
rect 8757 25347 8815 25353
rect 8757 25313 8769 25347
rect 8803 25344 8815 25347
rect 8846 25344 8852 25356
rect 8803 25316 8852 25344
rect 8803 25313 8815 25316
rect 8757 25307 8815 25313
rect 8846 25304 8852 25316
rect 8904 25304 8910 25356
rect 9306 25304 9312 25356
rect 9364 25344 9370 25356
rect 9585 25347 9643 25353
rect 9585 25344 9597 25347
rect 9364 25316 9597 25344
rect 9364 25304 9370 25316
rect 9585 25313 9597 25316
rect 9631 25313 9643 25347
rect 9585 25307 9643 25313
rect 11330 25304 11336 25356
rect 11388 25304 11394 25356
rect 11974 25304 11980 25356
rect 12032 25344 12038 25356
rect 13173 25347 13231 25353
rect 13173 25344 13185 25347
rect 12032 25316 13185 25344
rect 12032 25304 12038 25316
rect 13173 25313 13185 25316
rect 13219 25313 13231 25347
rect 13173 25307 13231 25313
rect 13814 25304 13820 25356
rect 13872 25344 13878 25356
rect 13872 25316 14412 25344
rect 13872 25304 13878 25316
rect 9214 25236 9220 25288
rect 9272 25276 9278 25288
rect 10413 25279 10471 25285
rect 10413 25276 10425 25279
rect 9272 25248 10425 25276
rect 9272 25236 9278 25248
rect 10413 25245 10425 25248
rect 10459 25245 10471 25279
rect 10413 25239 10471 25245
rect 11238 25236 11244 25288
rect 11296 25236 11302 25288
rect 12345 25279 12403 25285
rect 12345 25245 12357 25279
rect 12391 25245 12403 25279
rect 12345 25239 12403 25245
rect 9401 25211 9459 25217
rect 9401 25177 9413 25211
rect 9447 25208 9459 25211
rect 10134 25208 10140 25220
rect 9447 25180 10140 25208
rect 9447 25177 9459 25180
rect 9401 25171 9459 25177
rect 10134 25168 10140 25180
rect 10192 25168 10198 25220
rect 12360 25208 12388 25239
rect 12986 25236 12992 25288
rect 13044 25236 13050 25288
rect 14090 25236 14096 25288
rect 14148 25276 14154 25288
rect 14384 25285 14412 25316
rect 14458 25304 14464 25356
rect 14516 25304 14522 25356
rect 14277 25279 14335 25285
rect 14277 25276 14289 25279
rect 14148 25248 14289 25276
rect 14148 25236 14154 25248
rect 14277 25245 14289 25248
rect 14323 25245 14335 25279
rect 14277 25239 14335 25245
rect 14369 25279 14427 25285
rect 14369 25245 14381 25279
rect 14415 25245 14427 25279
rect 14369 25239 14427 25245
rect 13998 25208 14004 25220
rect 12360 25180 14004 25208
rect 13998 25168 14004 25180
rect 14056 25168 14062 25220
rect 7984 25112 8432 25140
rect 9493 25143 9551 25149
rect 7984 25100 7990 25112
rect 9493 25109 9505 25143
rect 9539 25140 9551 25143
rect 9861 25143 9919 25149
rect 9861 25140 9873 25143
rect 9539 25112 9873 25140
rect 9539 25109 9551 25112
rect 9493 25103 9551 25109
rect 9861 25109 9873 25112
rect 9907 25109 9919 25143
rect 9861 25103 9919 25109
rect 11977 25143 12035 25149
rect 11977 25109 11989 25143
rect 12023 25140 12035 25143
rect 12066 25140 12072 25152
rect 12023 25112 12072 25140
rect 12023 25109 12035 25112
rect 11977 25103 12035 25109
rect 12066 25100 12072 25112
rect 12124 25100 12130 25152
rect 12158 25100 12164 25152
rect 12216 25100 12222 25152
rect 12250 25100 12256 25152
rect 12308 25140 12314 25152
rect 12437 25143 12495 25149
rect 12437 25140 12449 25143
rect 12308 25112 12449 25140
rect 12308 25100 12314 25112
rect 12437 25109 12449 25112
rect 12483 25109 12495 25143
rect 12437 25103 12495 25109
rect 13354 25100 13360 25152
rect 13412 25140 13418 25152
rect 13817 25143 13875 25149
rect 13817 25140 13829 25143
rect 13412 25112 13829 25140
rect 13412 25100 13418 25112
rect 13817 25109 13829 25112
rect 13863 25109 13875 25143
rect 13817 25103 13875 25109
rect 14093 25143 14151 25149
rect 14093 25109 14105 25143
rect 14139 25140 14151 25143
rect 14476 25140 14504 25304
rect 14660 25285 14688 25384
rect 14918 25304 14924 25356
rect 14976 25304 14982 25356
rect 14553 25279 14611 25285
rect 14553 25245 14565 25279
rect 14599 25245 14611 25279
rect 14553 25239 14611 25245
rect 14645 25279 14703 25285
rect 14645 25245 14657 25279
rect 14691 25245 14703 25279
rect 14645 25239 14703 25245
rect 14139 25112 14504 25140
rect 14568 25140 14596 25239
rect 15194 25217 15200 25220
rect 15188 25171 15200 25217
rect 15194 25168 15200 25171
rect 15252 25168 15258 25220
rect 15562 25140 15568 25152
rect 14568 25112 15568 25140
rect 14139 25109 14151 25112
rect 14093 25103 14151 25109
rect 15562 25100 15568 25112
rect 15620 25100 15626 25152
rect 16206 25100 16212 25152
rect 16264 25140 16270 25152
rect 16301 25143 16359 25149
rect 16301 25140 16313 25143
rect 16264 25112 16313 25140
rect 16264 25100 16270 25112
rect 16301 25109 16313 25112
rect 16347 25109 16359 25143
rect 16301 25103 16359 25109
rect 1104 25050 16652 25072
rect 1104 24998 4874 25050
rect 4926 24998 4938 25050
rect 4990 24998 5002 25050
rect 5054 24998 5066 25050
rect 5118 24998 5130 25050
rect 5182 24998 16652 25050
rect 1104 24976 16652 24998
rect 2038 24896 2044 24948
rect 2096 24936 2102 24948
rect 4614 24936 4620 24948
rect 2096 24908 4620 24936
rect 2096 24896 2102 24908
rect 4614 24896 4620 24908
rect 4672 24896 4678 24948
rect 7650 24896 7656 24948
rect 7708 24936 7714 24948
rect 7708 24908 8064 24936
rect 7708 24896 7714 24908
rect 3602 24828 3608 24880
rect 3660 24868 3666 24880
rect 4706 24868 4712 24880
rect 3660 24840 4016 24868
rect 3660 24828 3666 24840
rect 3988 24812 4016 24840
rect 4172 24840 4712 24868
rect 1949 24803 2007 24809
rect 1949 24769 1961 24803
rect 1995 24800 2007 24803
rect 2866 24800 2872 24812
rect 1995 24772 2872 24800
rect 1995 24769 2007 24772
rect 1949 24763 2007 24769
rect 2866 24760 2872 24772
rect 2924 24800 2930 24812
rect 3418 24800 3424 24812
rect 2924 24772 3424 24800
rect 2924 24760 2930 24772
rect 3418 24760 3424 24772
rect 3476 24760 3482 24812
rect 3510 24760 3516 24812
rect 3568 24760 3574 24812
rect 3970 24760 3976 24812
rect 4028 24760 4034 24812
rect 4172 24809 4200 24840
rect 4706 24828 4712 24840
rect 4764 24828 4770 24880
rect 7834 24868 7840 24880
rect 7024 24840 7840 24868
rect 4157 24803 4215 24809
rect 4157 24769 4169 24803
rect 4203 24769 4215 24803
rect 4617 24803 4675 24809
rect 4617 24800 4629 24803
rect 4157 24763 4215 24769
rect 4264 24772 4629 24800
rect 1854 24741 1860 24744
rect 1832 24735 1860 24741
rect 1832 24701 1844 24735
rect 1832 24695 1860 24701
rect 1854 24692 1860 24695
rect 1912 24692 1918 24744
rect 2317 24735 2375 24741
rect 2317 24701 2329 24735
rect 2363 24732 2375 24735
rect 2590 24732 2596 24744
rect 2363 24704 2596 24732
rect 2363 24701 2375 24704
rect 2317 24695 2375 24701
rect 2590 24692 2596 24704
rect 2648 24692 2654 24744
rect 3878 24692 3884 24744
rect 3936 24692 3942 24744
rect 3786 24624 3792 24676
rect 3844 24664 3850 24676
rect 4264 24664 4292 24772
rect 4617 24769 4629 24772
rect 4663 24769 4675 24803
rect 4617 24763 4675 24769
rect 5261 24803 5319 24809
rect 5261 24769 5273 24803
rect 5307 24769 5319 24803
rect 5261 24763 5319 24769
rect 5445 24803 5503 24809
rect 5445 24769 5457 24803
rect 5491 24769 5503 24803
rect 5445 24763 5503 24769
rect 4801 24735 4859 24741
rect 4801 24701 4813 24735
rect 4847 24732 4859 24735
rect 4890 24732 4896 24744
rect 4847 24704 4896 24732
rect 4847 24701 4859 24704
rect 4801 24695 4859 24701
rect 4890 24692 4896 24704
rect 4948 24692 4954 24744
rect 3844 24636 4292 24664
rect 4341 24667 4399 24673
rect 3844 24624 3850 24636
rect 4341 24633 4353 24667
rect 4387 24664 4399 24667
rect 4614 24664 4620 24676
rect 4387 24636 4620 24664
rect 4387 24633 4399 24636
rect 4341 24627 4399 24633
rect 4614 24624 4620 24636
rect 4672 24624 4678 24676
rect 5276 24664 5304 24763
rect 5460 24732 5488 24763
rect 5626 24760 5632 24812
rect 5684 24760 5690 24812
rect 5810 24760 5816 24812
rect 5868 24800 5874 24812
rect 6365 24803 6423 24809
rect 6365 24800 6377 24803
rect 5868 24772 6377 24800
rect 5868 24760 5874 24772
rect 6365 24769 6377 24772
rect 6411 24769 6423 24803
rect 6365 24763 6423 24769
rect 6549 24803 6607 24809
rect 6549 24769 6561 24803
rect 6595 24769 6607 24803
rect 6549 24763 6607 24769
rect 6825 24803 6883 24809
rect 6825 24769 6837 24803
rect 6871 24800 6883 24803
rect 7024 24800 7052 24840
rect 7834 24828 7840 24840
rect 7892 24828 7898 24880
rect 8036 24868 8064 24908
rect 8110 24896 8116 24948
rect 8168 24936 8174 24948
rect 8757 24939 8815 24945
rect 8757 24936 8769 24939
rect 8168 24908 8769 24936
rect 8168 24896 8174 24908
rect 8757 24905 8769 24908
rect 8803 24905 8815 24939
rect 8757 24899 8815 24905
rect 9306 24896 9312 24948
rect 9364 24896 9370 24948
rect 11330 24896 11336 24948
rect 11388 24896 11394 24948
rect 12897 24939 12955 24945
rect 12897 24905 12909 24939
rect 12943 24936 12955 24939
rect 12986 24936 12992 24948
rect 12943 24908 12992 24936
rect 12943 24905 12955 24908
rect 12897 24899 12955 24905
rect 12986 24896 12992 24908
rect 13044 24896 13050 24948
rect 13354 24896 13360 24948
rect 13412 24896 13418 24948
rect 13538 24896 13544 24948
rect 13596 24936 13602 24948
rect 15746 24936 15752 24948
rect 13596 24908 15752 24936
rect 13596 24896 13602 24908
rect 15746 24896 15752 24908
rect 15804 24896 15810 24948
rect 8036 24840 8340 24868
rect 7098 24809 7104 24812
rect 6871 24772 7052 24800
rect 6871 24769 6883 24772
rect 6825 24763 6883 24769
rect 7092 24763 7104 24809
rect 6457 24735 6515 24741
rect 6457 24732 6469 24735
rect 5460 24704 6469 24732
rect 6457 24701 6469 24704
rect 6503 24701 6515 24735
rect 6457 24695 6515 24701
rect 5810 24664 5816 24676
rect 5276 24636 5816 24664
rect 5810 24624 5816 24636
rect 5868 24664 5874 24676
rect 6178 24664 6184 24676
rect 5868 24636 6184 24664
rect 5868 24624 5874 24636
rect 6178 24624 6184 24636
rect 6236 24624 6242 24676
rect 6270 24624 6276 24676
rect 6328 24664 6334 24676
rect 6564 24664 6592 24763
rect 7098 24760 7104 24763
rect 7156 24760 7162 24812
rect 8312 24800 8340 24840
rect 8662 24828 8668 24880
rect 8720 24828 8726 24880
rect 15010 24868 15016 24880
rect 14476 24840 15016 24868
rect 9217 24803 9275 24809
rect 9217 24800 9229 24803
rect 8312 24772 9229 24800
rect 9217 24769 9229 24772
rect 9263 24769 9275 24803
rect 9217 24763 9275 24769
rect 9674 24760 9680 24812
rect 9732 24800 9738 24812
rect 9953 24803 10011 24809
rect 9953 24800 9965 24803
rect 9732 24772 9965 24800
rect 9732 24760 9738 24772
rect 9953 24769 9965 24772
rect 9999 24769 10011 24803
rect 9953 24763 10011 24769
rect 10220 24803 10278 24809
rect 10220 24769 10232 24803
rect 10266 24800 10278 24803
rect 11238 24800 11244 24812
rect 10266 24772 11244 24800
rect 10266 24769 10278 24772
rect 10220 24763 10278 24769
rect 11238 24760 11244 24772
rect 11296 24760 11302 24812
rect 11606 24760 11612 24812
rect 11664 24800 11670 24812
rect 11773 24803 11831 24809
rect 11773 24800 11785 24803
rect 11664 24772 11785 24800
rect 11664 24760 11670 24772
rect 11773 24769 11785 24772
rect 11819 24769 11831 24803
rect 11773 24763 11831 24769
rect 12342 24760 12348 24812
rect 12400 24800 12406 24812
rect 13449 24803 13507 24809
rect 12400 24772 12572 24800
rect 12400 24760 12406 24772
rect 8294 24692 8300 24744
rect 8352 24732 8358 24744
rect 8941 24735 8999 24741
rect 8941 24732 8953 24735
rect 8352 24704 8953 24732
rect 8352 24692 8358 24704
rect 8941 24701 8953 24704
rect 8987 24732 8999 24735
rect 9306 24732 9312 24744
rect 8987 24704 9312 24732
rect 8987 24701 8999 24704
rect 8941 24695 8999 24701
rect 9306 24692 9312 24704
rect 9364 24692 9370 24744
rect 11514 24692 11520 24744
rect 11572 24692 11578 24744
rect 6328 24636 6592 24664
rect 12544 24664 12572 24772
rect 13449 24769 13461 24803
rect 13495 24800 13507 24803
rect 13722 24800 13728 24812
rect 13495 24772 13728 24800
rect 13495 24769 13507 24772
rect 13449 24763 13507 24769
rect 13722 24760 13728 24772
rect 13780 24760 13786 24812
rect 14093 24803 14151 24809
rect 14093 24769 14105 24803
rect 14139 24769 14151 24803
rect 14093 24763 14151 24769
rect 14185 24803 14243 24809
rect 14185 24769 14197 24803
rect 14231 24800 14243 24803
rect 14274 24800 14280 24812
rect 14231 24772 14280 24800
rect 14231 24769 14243 24772
rect 14185 24763 14243 24769
rect 12618 24692 12624 24744
rect 12676 24732 12682 24744
rect 13541 24735 13599 24741
rect 13541 24732 13553 24735
rect 12676 24704 13553 24732
rect 12676 24692 12682 24704
rect 13541 24701 13553 24704
rect 13587 24701 13599 24735
rect 14108 24732 14136 24763
rect 14274 24760 14280 24772
rect 14332 24760 14338 24812
rect 14366 24760 14372 24812
rect 14424 24760 14430 24812
rect 14476 24809 14504 24840
rect 15010 24828 15016 24840
rect 15068 24828 15074 24880
rect 16206 24868 16212 24880
rect 15120 24840 16212 24868
rect 14461 24803 14519 24809
rect 14461 24769 14473 24803
rect 14507 24769 14519 24803
rect 14461 24763 14519 24769
rect 14550 24760 14556 24812
rect 14608 24760 14614 24812
rect 14918 24760 14924 24812
rect 14976 24760 14982 24812
rect 15120 24800 15148 24840
rect 16206 24828 16212 24840
rect 16264 24828 16270 24880
rect 15028 24772 15148 24800
rect 15188 24803 15246 24809
rect 15028 24732 15056 24772
rect 15188 24769 15200 24803
rect 15234 24800 15246 24803
rect 15470 24800 15476 24812
rect 15234 24772 15476 24800
rect 15234 24769 15246 24772
rect 15188 24763 15246 24769
rect 15470 24760 15476 24772
rect 15528 24760 15534 24812
rect 14108 24704 15056 24732
rect 13541 24695 13599 24701
rect 12544 24636 13860 24664
rect 6328 24624 6334 24636
rect 1673 24599 1731 24605
rect 1673 24565 1685 24599
rect 1719 24596 1731 24599
rect 1762 24596 1768 24608
rect 1719 24568 1768 24596
rect 1719 24565 1731 24568
rect 1673 24559 1731 24565
rect 1762 24556 1768 24568
rect 1820 24556 1826 24608
rect 3418 24556 3424 24608
rect 3476 24596 3482 24608
rect 3697 24599 3755 24605
rect 3697 24596 3709 24599
rect 3476 24568 3709 24596
rect 3476 24556 3482 24568
rect 3697 24565 3709 24568
rect 3743 24596 3755 24599
rect 4062 24596 4068 24608
rect 3743 24568 4068 24596
rect 3743 24565 3755 24568
rect 3697 24559 3755 24565
rect 4062 24556 4068 24568
rect 4120 24556 4126 24608
rect 4433 24599 4491 24605
rect 4433 24565 4445 24599
rect 4479 24596 4491 24599
rect 4706 24596 4712 24608
rect 4479 24568 4712 24596
rect 4479 24565 4491 24568
rect 4433 24559 4491 24565
rect 4706 24556 4712 24568
rect 4764 24556 4770 24608
rect 5442 24556 5448 24608
rect 5500 24556 5506 24608
rect 7742 24556 7748 24608
rect 7800 24596 7806 24608
rect 8205 24599 8263 24605
rect 8205 24596 8217 24599
rect 7800 24568 8217 24596
rect 7800 24556 7806 24568
rect 8205 24565 8217 24568
rect 8251 24565 8263 24599
rect 8205 24559 8263 24565
rect 8297 24599 8355 24605
rect 8297 24565 8309 24599
rect 8343 24596 8355 24599
rect 8478 24596 8484 24608
rect 8343 24568 8484 24596
rect 8343 24565 8355 24568
rect 8297 24559 8355 24565
rect 8478 24556 8484 24568
rect 8536 24556 8542 24608
rect 11422 24556 11428 24608
rect 11480 24596 11486 24608
rect 12802 24596 12808 24608
rect 11480 24568 12808 24596
rect 11480 24556 11486 24568
rect 12802 24556 12808 24568
rect 12860 24556 12866 24608
rect 12986 24556 12992 24608
rect 13044 24556 13050 24608
rect 13832 24596 13860 24636
rect 13906 24624 13912 24676
rect 13964 24624 13970 24676
rect 14090 24624 14096 24676
rect 14148 24664 14154 24676
rect 14366 24664 14372 24676
rect 14148 24636 14372 24664
rect 14148 24624 14154 24636
rect 14366 24624 14372 24636
rect 14424 24624 14430 24676
rect 14734 24624 14740 24676
rect 14792 24664 14798 24676
rect 14918 24664 14924 24676
rect 14792 24636 14924 24664
rect 14792 24624 14798 24636
rect 14918 24624 14924 24636
rect 14976 24624 14982 24676
rect 14642 24596 14648 24608
rect 13832 24568 14648 24596
rect 14642 24556 14648 24568
rect 14700 24556 14706 24608
rect 14829 24599 14887 24605
rect 14829 24565 14841 24599
rect 14875 24596 14887 24599
rect 15194 24596 15200 24608
rect 14875 24568 15200 24596
rect 14875 24565 14887 24568
rect 14829 24559 14887 24565
rect 15194 24556 15200 24568
rect 15252 24556 15258 24608
rect 15286 24556 15292 24608
rect 15344 24596 15350 24608
rect 15654 24596 15660 24608
rect 15344 24568 15660 24596
rect 15344 24556 15350 24568
rect 15654 24556 15660 24568
rect 15712 24556 15718 24608
rect 15838 24556 15844 24608
rect 15896 24596 15902 24608
rect 16301 24599 16359 24605
rect 16301 24596 16313 24599
rect 15896 24568 16313 24596
rect 15896 24556 15902 24568
rect 16301 24565 16313 24568
rect 16347 24565 16359 24599
rect 16301 24559 16359 24565
rect 1104 24506 16652 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 16652 24506
rect 1104 24432 16652 24454
rect 1854 24352 1860 24404
rect 1912 24392 1918 24404
rect 2961 24395 3019 24401
rect 2961 24392 2973 24395
rect 1912 24364 2973 24392
rect 1912 24352 1918 24364
rect 2961 24361 2973 24364
rect 3007 24361 3019 24395
rect 2961 24355 3019 24361
rect 4246 24352 4252 24404
rect 4304 24392 4310 24404
rect 4890 24392 4896 24404
rect 4304 24364 4896 24392
rect 4304 24352 4310 24364
rect 4890 24352 4896 24364
rect 4948 24352 4954 24404
rect 5350 24352 5356 24404
rect 5408 24392 5414 24404
rect 5408 24364 6132 24392
rect 5408 24352 5414 24364
rect 3881 24327 3939 24333
rect 3881 24293 3893 24327
rect 3927 24324 3939 24327
rect 3970 24324 3976 24336
rect 3927 24296 3976 24324
rect 3927 24293 3939 24296
rect 3881 24287 3939 24293
rect 3970 24284 3976 24296
rect 4028 24284 4034 24336
rect 4908 24324 4936 24352
rect 6104 24324 6132 24364
rect 6178 24352 6184 24404
rect 6236 24392 6242 24404
rect 6641 24395 6699 24401
rect 6641 24392 6653 24395
rect 6236 24364 6653 24392
rect 6236 24352 6242 24364
rect 6641 24361 6653 24364
rect 6687 24361 6699 24395
rect 6641 24355 6699 24361
rect 7098 24352 7104 24404
rect 7156 24392 7162 24404
rect 7193 24395 7251 24401
rect 7193 24392 7205 24395
rect 7156 24364 7205 24392
rect 7156 24352 7162 24364
rect 7193 24361 7205 24364
rect 7239 24361 7251 24395
rect 7193 24355 7251 24361
rect 7377 24395 7435 24401
rect 7377 24361 7389 24395
rect 7423 24392 7435 24395
rect 8846 24392 8852 24404
rect 7423 24364 8852 24392
rect 7423 24361 7435 24364
rect 7377 24355 7435 24361
rect 8846 24352 8852 24364
rect 8904 24352 8910 24404
rect 10134 24352 10140 24404
rect 10192 24352 10198 24404
rect 10226 24352 10232 24404
rect 10284 24392 10290 24404
rect 10686 24392 10692 24404
rect 10284 24364 10692 24392
rect 10284 24352 10290 24364
rect 10686 24352 10692 24364
rect 10744 24352 10750 24404
rect 12250 24392 12256 24404
rect 10980 24364 12256 24392
rect 10980 24324 11008 24364
rect 12250 24352 12256 24364
rect 12308 24352 12314 24404
rect 13170 24352 13176 24404
rect 13228 24392 13234 24404
rect 13228 24364 13400 24392
rect 13228 24352 13234 24364
rect 4908 24296 6040 24324
rect 6104 24296 6500 24324
rect 3050 24256 3056 24268
rect 2884 24228 3056 24256
rect 1394 24148 1400 24200
rect 1452 24188 1458 24200
rect 1762 24197 1768 24200
rect 1489 24191 1547 24197
rect 1489 24188 1501 24191
rect 1452 24160 1501 24188
rect 1452 24148 1458 24160
rect 1489 24157 1501 24160
rect 1535 24157 1547 24191
rect 1756 24188 1768 24197
rect 1723 24160 1768 24188
rect 1489 24151 1547 24157
rect 1756 24151 1768 24160
rect 1762 24148 1768 24151
rect 1820 24148 1826 24200
rect 2038 24148 2044 24200
rect 2096 24188 2102 24200
rect 2884 24188 2912 24228
rect 3050 24216 3056 24228
rect 3108 24256 3114 24268
rect 4617 24259 4675 24265
rect 4617 24256 4629 24259
rect 3108 24228 4629 24256
rect 3108 24216 3114 24228
rect 4617 24225 4629 24228
rect 4663 24225 4675 24259
rect 4617 24219 4675 24225
rect 2096 24160 2912 24188
rect 2096 24148 2102 24160
rect 2958 24148 2964 24200
rect 3016 24148 3022 24200
rect 3142 24148 3148 24200
rect 3200 24148 3206 24200
rect 3418 24148 3424 24200
rect 3476 24197 3482 24200
rect 3476 24191 3509 24197
rect 3497 24157 3509 24191
rect 3476 24151 3509 24157
rect 3476 24148 3482 24151
rect 3602 24148 3608 24200
rect 3660 24148 3666 24200
rect 3789 24191 3847 24197
rect 3789 24157 3801 24191
rect 3835 24157 3847 24191
rect 3789 24151 3847 24157
rect 3973 24191 4031 24197
rect 3973 24157 3985 24191
rect 4019 24157 4031 24191
rect 3973 24151 4031 24157
rect 2590 24080 2596 24132
rect 2648 24120 2654 24132
rect 3160 24120 3188 24148
rect 2648 24092 3188 24120
rect 3237 24123 3295 24129
rect 2648 24080 2654 24092
rect 3237 24089 3249 24123
rect 3283 24120 3295 24123
rect 3326 24120 3332 24132
rect 3283 24092 3332 24120
rect 3283 24089 3295 24092
rect 3237 24083 3295 24089
rect 3326 24080 3332 24092
rect 3384 24120 3390 24132
rect 3804 24120 3832 24151
rect 3384 24092 3832 24120
rect 3384 24080 3390 24092
rect 2869 24055 2927 24061
rect 2869 24021 2881 24055
rect 2915 24052 2927 24055
rect 3050 24052 3056 24064
rect 2915 24024 3056 24052
rect 2915 24021 2927 24024
rect 2869 24015 2927 24021
rect 3050 24012 3056 24024
rect 3108 24012 3114 24064
rect 3142 24012 3148 24064
rect 3200 24052 3206 24064
rect 3988 24052 4016 24151
rect 4062 24148 4068 24200
rect 4120 24188 4126 24200
rect 4157 24191 4215 24197
rect 4157 24188 4169 24191
rect 4120 24160 4169 24188
rect 4120 24148 4126 24160
rect 4157 24157 4169 24160
rect 4203 24157 4215 24191
rect 4632 24188 4660 24219
rect 4982 24216 4988 24268
rect 5040 24216 5046 24268
rect 5102 24259 5160 24265
rect 5102 24225 5114 24259
rect 5148 24256 5160 24259
rect 5442 24256 5448 24268
rect 5148 24228 5448 24256
rect 5148 24225 5160 24228
rect 5102 24219 5160 24225
rect 5442 24216 5448 24228
rect 5500 24216 5506 24268
rect 5629 24259 5687 24265
rect 5629 24225 5641 24259
rect 5675 24256 5687 24259
rect 5902 24256 5908 24268
rect 5675 24228 5908 24256
rect 5675 24225 5687 24228
rect 5629 24219 5687 24225
rect 5353 24191 5411 24197
rect 5353 24188 5365 24191
rect 4632 24160 5365 24188
rect 4157 24151 4215 24157
rect 5353 24157 5365 24160
rect 5399 24157 5411 24191
rect 5644 24188 5672 24219
rect 5902 24216 5908 24228
rect 5960 24216 5966 24268
rect 5353 24151 5411 24157
rect 5460 24160 5672 24188
rect 6012 24188 6040 24296
rect 6472 24197 6500 24296
rect 9784 24296 11008 24324
rect 7009 24259 7067 24265
rect 7009 24225 7021 24259
rect 7055 24256 7067 24259
rect 7374 24256 7380 24268
rect 7055 24228 7380 24256
rect 7055 24225 7067 24228
rect 7009 24219 7067 24225
rect 7374 24216 7380 24228
rect 7432 24216 7438 24268
rect 6365 24191 6423 24197
rect 6365 24188 6377 24191
rect 6012 24160 6377 24188
rect 4893 24123 4951 24129
rect 4893 24089 4905 24123
rect 4939 24120 4951 24123
rect 5166 24120 5172 24132
rect 4939 24092 5172 24120
rect 4939 24089 4951 24092
rect 4893 24083 4951 24089
rect 5166 24080 5172 24092
rect 5224 24120 5230 24132
rect 5460 24120 5488 24160
rect 6365 24157 6377 24160
rect 6411 24157 6423 24191
rect 6365 24151 6423 24157
rect 6457 24191 6515 24197
rect 6457 24157 6469 24191
rect 6503 24157 6515 24191
rect 6457 24151 6515 24157
rect 6917 24191 6975 24197
rect 6917 24157 6929 24191
rect 6963 24188 6975 24191
rect 7558 24188 7564 24200
rect 6963 24160 7564 24188
rect 6963 24157 6975 24160
rect 6917 24151 6975 24157
rect 7558 24148 7564 24160
rect 7616 24148 7622 24200
rect 8478 24148 8484 24200
rect 8536 24197 8542 24200
rect 8536 24188 8548 24197
rect 8757 24191 8815 24197
rect 8536 24160 8581 24188
rect 8536 24151 8548 24160
rect 8757 24157 8769 24191
rect 8803 24188 8815 24191
rect 9214 24188 9220 24200
rect 8803 24160 9220 24188
rect 8803 24157 8815 24160
rect 8757 24151 8815 24157
rect 8536 24148 8542 24151
rect 9214 24148 9220 24160
rect 9272 24148 9278 24200
rect 9784 24197 9812 24296
rect 11054 24284 11060 24336
rect 11112 24324 11118 24336
rect 11974 24324 11980 24336
rect 11112 24296 11980 24324
rect 11112 24284 11118 24296
rect 11974 24284 11980 24296
rect 12032 24284 12038 24336
rect 10594 24216 10600 24268
rect 10652 24216 10658 24268
rect 10686 24216 10692 24268
rect 10744 24216 10750 24268
rect 11422 24256 11428 24268
rect 11256 24228 11428 24256
rect 9769 24191 9827 24197
rect 9769 24157 9781 24191
rect 9815 24157 9827 24191
rect 9769 24151 9827 24157
rect 9858 24148 9864 24200
rect 9916 24148 9922 24200
rect 11256 24197 11284 24228
rect 11422 24216 11428 24228
rect 11480 24216 11486 24268
rect 12158 24256 12164 24268
rect 11532 24228 12164 24256
rect 10045 24191 10103 24197
rect 10045 24157 10057 24191
rect 10091 24188 10103 24191
rect 11241 24191 11299 24197
rect 11241 24188 11253 24191
rect 10091 24160 11253 24188
rect 10091 24157 10103 24160
rect 10045 24151 10103 24157
rect 11241 24157 11253 24160
rect 11287 24157 11299 24191
rect 11241 24151 11299 24157
rect 11330 24148 11336 24200
rect 11388 24148 11394 24200
rect 11532 24197 11560 24228
rect 12158 24216 12164 24228
rect 12216 24216 12222 24268
rect 13372 24265 13400 24364
rect 14274 24352 14280 24404
rect 14332 24392 14338 24404
rect 14918 24392 14924 24404
rect 14332 24364 14924 24392
rect 14332 24352 14338 24364
rect 14918 24352 14924 24364
rect 14976 24352 14982 24404
rect 15470 24352 15476 24404
rect 15528 24352 15534 24404
rect 15562 24352 15568 24404
rect 15620 24352 15626 24404
rect 13630 24284 13636 24336
rect 13688 24324 13694 24336
rect 13998 24324 14004 24336
rect 13688 24296 14004 24324
rect 13688 24284 13694 24296
rect 13998 24284 14004 24296
rect 14056 24284 14062 24336
rect 14550 24284 14556 24336
rect 14608 24284 14614 24336
rect 15102 24284 15108 24336
rect 15160 24324 15166 24336
rect 15160 24296 15792 24324
rect 15160 24284 15166 24296
rect 13357 24259 13415 24265
rect 13357 24225 13369 24259
rect 13403 24225 13415 24259
rect 13814 24256 13820 24268
rect 13357 24219 13415 24225
rect 13740 24228 13820 24256
rect 11517 24191 11575 24197
rect 11517 24157 11529 24191
rect 11563 24157 11575 24191
rect 11517 24151 11575 24157
rect 11609 24191 11667 24197
rect 11609 24157 11621 24191
rect 11655 24188 11667 24191
rect 11698 24188 11704 24200
rect 11655 24160 11704 24188
rect 11655 24157 11667 24160
rect 11609 24151 11667 24157
rect 11698 24148 11704 24160
rect 11756 24148 11762 24200
rect 11793 24191 11851 24197
rect 11793 24157 11805 24191
rect 11839 24188 11851 24191
rect 12250 24188 12256 24200
rect 11839 24160 12256 24188
rect 11839 24157 11851 24160
rect 11793 24151 11851 24157
rect 12250 24148 12256 24160
rect 12308 24148 12314 24200
rect 13541 24191 13599 24197
rect 13541 24157 13553 24191
rect 13587 24188 13599 24191
rect 13630 24188 13636 24200
rect 13587 24160 13636 24188
rect 13587 24157 13599 24160
rect 13541 24151 13599 24157
rect 13630 24148 13636 24160
rect 13688 24148 13694 24200
rect 13740 24197 13768 24228
rect 13814 24216 13820 24228
rect 13872 24216 13878 24268
rect 13906 24216 13912 24268
rect 13964 24256 13970 24268
rect 14568 24256 14596 24284
rect 13964 24228 15240 24256
rect 13964 24216 13970 24228
rect 14384 24197 14412 24228
rect 13725 24191 13783 24197
rect 13725 24157 13737 24191
rect 13771 24157 13783 24191
rect 13725 24151 13783 24157
rect 14369 24191 14427 24197
rect 14369 24157 14381 24191
rect 14415 24157 14427 24191
rect 14369 24151 14427 24157
rect 14458 24148 14464 24200
rect 14516 24148 14522 24200
rect 14553 24188 14611 24194
rect 14553 24154 14565 24188
rect 14599 24154 14611 24188
rect 14553 24148 14611 24154
rect 14737 24191 14795 24197
rect 14737 24157 14749 24191
rect 14783 24188 14795 24191
rect 14829 24191 14887 24197
rect 14829 24188 14841 24191
rect 14783 24160 14841 24188
rect 14783 24157 14795 24160
rect 14737 24151 14795 24157
rect 14829 24157 14841 24160
rect 14875 24188 14887 24191
rect 14918 24188 14924 24200
rect 14875 24160 14924 24188
rect 14875 24157 14887 24160
rect 14829 24151 14887 24157
rect 14918 24148 14924 24160
rect 14976 24148 14982 24200
rect 15010 24148 15016 24200
rect 15068 24148 15074 24200
rect 15212 24197 15240 24228
rect 15105 24191 15163 24197
rect 15105 24157 15117 24191
rect 15151 24157 15163 24191
rect 15105 24151 15163 24157
rect 15197 24191 15255 24197
rect 15197 24157 15209 24191
rect 15243 24157 15255 24191
rect 15197 24151 15255 24157
rect 5224 24092 5488 24120
rect 5224 24080 5230 24092
rect 5534 24080 5540 24132
rect 5592 24120 5598 24132
rect 5838 24123 5896 24129
rect 5838 24120 5850 24123
rect 5592 24092 5850 24120
rect 5592 24080 5598 24092
rect 5838 24089 5850 24092
rect 5884 24089 5896 24123
rect 5838 24083 5896 24089
rect 6086 24080 6092 24132
rect 6144 24080 6150 24132
rect 9953 24123 10011 24129
rect 9953 24089 9965 24123
rect 9999 24120 10011 24123
rect 12526 24120 12532 24132
rect 9999 24092 12532 24120
rect 9999 24089 10011 24092
rect 9953 24083 10011 24089
rect 12526 24080 12532 24092
rect 12584 24080 12590 24132
rect 12986 24080 12992 24132
rect 13044 24120 13050 24132
rect 13090 24123 13148 24129
rect 13090 24120 13102 24123
rect 13044 24092 13102 24120
rect 13044 24080 13050 24092
rect 13090 24089 13102 24092
rect 13136 24089 13148 24123
rect 13090 24083 13148 24089
rect 13909 24123 13967 24129
rect 13909 24089 13921 24123
rect 13955 24120 13967 24123
rect 14568 24120 14596 24148
rect 13955 24092 14596 24120
rect 15120 24120 15148 24151
rect 15562 24148 15568 24200
rect 15620 24188 15626 24200
rect 15764 24197 15792 24296
rect 15749 24191 15807 24197
rect 15749 24188 15761 24191
rect 15620 24160 15761 24188
rect 15620 24148 15626 24160
rect 15749 24157 15761 24160
rect 15795 24157 15807 24191
rect 15749 24151 15807 24157
rect 16117 24191 16175 24197
rect 16117 24157 16129 24191
rect 16163 24188 16175 24191
rect 16206 24188 16212 24200
rect 16163 24160 16212 24188
rect 16163 24157 16175 24160
rect 16117 24151 16175 24157
rect 16206 24148 16212 24160
rect 16264 24148 16270 24200
rect 15378 24120 15384 24132
rect 15120 24092 15384 24120
rect 13955 24089 13967 24092
rect 13909 24083 13967 24089
rect 15378 24080 15384 24092
rect 15436 24080 15442 24132
rect 15838 24080 15844 24132
rect 15896 24080 15902 24132
rect 15930 24080 15936 24132
rect 15988 24120 15994 24132
rect 16390 24120 16396 24132
rect 15988 24092 16396 24120
rect 15988 24080 15994 24092
rect 16390 24080 16396 24092
rect 16448 24080 16454 24132
rect 3200 24024 4016 24052
rect 3200 24012 3206 24024
rect 4062 24012 4068 24064
rect 4120 24052 4126 24064
rect 4249 24055 4307 24061
rect 4249 24052 4261 24055
rect 4120 24024 4261 24052
rect 4120 24012 4126 24024
rect 4249 24021 4261 24024
rect 4295 24021 4307 24055
rect 4249 24015 4307 24021
rect 5261 24055 5319 24061
rect 5261 24021 5273 24055
rect 5307 24052 5319 24055
rect 5350 24052 5356 24064
rect 5307 24024 5356 24052
rect 5307 24021 5319 24024
rect 5261 24015 5319 24021
rect 5350 24012 5356 24024
rect 5408 24012 5414 24064
rect 5442 24012 5448 24064
rect 5500 24052 5506 24064
rect 5721 24055 5779 24061
rect 5721 24052 5733 24055
rect 5500 24024 5733 24052
rect 5500 24012 5506 24024
rect 5721 24021 5733 24024
rect 5767 24021 5779 24055
rect 5721 24015 5779 24021
rect 5997 24055 6055 24061
rect 5997 24021 6009 24055
rect 6043 24052 6055 24055
rect 6178 24052 6184 24064
rect 6043 24024 6184 24052
rect 6043 24021 6055 24024
rect 5997 24015 6055 24021
rect 6178 24012 6184 24024
rect 6236 24012 6242 24064
rect 6270 24012 6276 24064
rect 6328 24012 6334 24064
rect 9674 24012 9680 24064
rect 9732 24012 9738 24064
rect 10505 24055 10563 24061
rect 10505 24021 10517 24055
rect 10551 24052 10563 24055
rect 10962 24052 10968 24064
rect 10551 24024 10968 24052
rect 10551 24021 10563 24024
rect 10505 24015 10563 24021
rect 10962 24012 10968 24024
rect 11020 24012 11026 24064
rect 11057 24055 11115 24061
rect 11057 24021 11069 24055
rect 11103 24052 11115 24055
rect 11146 24052 11152 24064
rect 11103 24024 11152 24052
rect 11103 24021 11115 24024
rect 11057 24015 11115 24021
rect 11146 24012 11152 24024
rect 11204 24052 11210 24064
rect 11330 24052 11336 24064
rect 11204 24024 11336 24052
rect 11204 24012 11210 24024
rect 11330 24012 11336 24024
rect 11388 24012 11394 24064
rect 11422 24012 11428 24064
rect 11480 24012 11486 24064
rect 11698 24012 11704 24064
rect 11756 24012 11762 24064
rect 14090 24012 14096 24064
rect 14148 24012 14154 24064
rect 14182 24012 14188 24064
rect 14240 24052 14246 24064
rect 15856 24052 15884 24080
rect 14240 24024 15884 24052
rect 14240 24012 14246 24024
rect 1104 23962 16652 23984
rect 1104 23910 4874 23962
rect 4926 23910 4938 23962
rect 4990 23910 5002 23962
rect 5054 23910 5066 23962
rect 5118 23910 5130 23962
rect 5182 23910 16652 23962
rect 1104 23888 16652 23910
rect 2958 23808 2964 23860
rect 3016 23808 3022 23860
rect 10594 23808 10600 23860
rect 10652 23808 10658 23860
rect 11532 23820 12204 23848
rect 11532 23792 11560 23820
rect 5626 23780 5632 23792
rect 1412 23752 5632 23780
rect 1412 23724 1440 23752
rect 1394 23672 1400 23724
rect 1452 23672 1458 23724
rect 1670 23721 1676 23724
rect 1664 23675 1676 23721
rect 1670 23672 1676 23675
rect 1728 23672 1734 23724
rect 2866 23672 2872 23724
rect 2924 23672 2930 23724
rect 3050 23672 3056 23724
rect 3108 23672 3114 23724
rect 3142 23672 3148 23724
rect 3200 23672 3206 23724
rect 3326 23672 3332 23724
rect 3384 23672 3390 23724
rect 3418 23672 3424 23724
rect 3476 23672 3482 23724
rect 3513 23715 3571 23721
rect 3513 23681 3525 23715
rect 3559 23681 3571 23715
rect 3513 23675 3571 23681
rect 3068 23644 3096 23672
rect 3528 23644 3556 23675
rect 3694 23672 3700 23724
rect 3752 23712 3758 23724
rect 4157 23715 4215 23721
rect 4157 23712 4169 23715
rect 3752 23684 4169 23712
rect 3752 23672 3758 23684
rect 4157 23681 4169 23684
rect 4203 23681 4215 23715
rect 4157 23675 4215 23681
rect 4246 23672 4252 23724
rect 4304 23672 4310 23724
rect 4816 23721 4844 23752
rect 5626 23740 5632 23752
rect 5684 23740 5690 23792
rect 9214 23740 9220 23792
rect 9272 23780 9278 23792
rect 11514 23780 11520 23792
rect 9272 23752 11520 23780
rect 9272 23740 9278 23752
rect 11514 23740 11520 23752
rect 11572 23740 11578 23792
rect 11793 23783 11851 23789
rect 11793 23749 11805 23783
rect 11839 23780 11851 23783
rect 11974 23780 11980 23792
rect 11839 23752 11980 23780
rect 11839 23749 11851 23752
rect 11793 23743 11851 23749
rect 11974 23740 11980 23752
rect 12032 23740 12038 23792
rect 4525 23715 4583 23721
rect 4525 23681 4537 23715
rect 4571 23681 4583 23715
rect 4525 23675 4583 23681
rect 4801 23715 4859 23721
rect 4801 23681 4813 23715
rect 4847 23681 4859 23715
rect 4801 23675 4859 23681
rect 5068 23715 5126 23721
rect 5068 23681 5080 23715
rect 5114 23712 5126 23715
rect 5350 23712 5356 23724
rect 5114 23684 5356 23712
rect 5114 23681 5126 23684
rect 5068 23675 5126 23681
rect 3068 23616 3556 23644
rect 3602 23604 3608 23656
rect 3660 23644 3666 23656
rect 4062 23644 4068 23656
rect 3660 23616 4068 23644
rect 3660 23604 3666 23616
rect 4062 23604 4068 23616
rect 4120 23644 4126 23656
rect 4540 23644 4568 23675
rect 5350 23672 5356 23684
rect 5408 23672 5414 23724
rect 9484 23715 9542 23721
rect 9484 23681 9496 23715
rect 9530 23712 9542 23715
rect 10502 23712 10508 23724
rect 9530 23684 10508 23712
rect 9530 23681 9542 23684
rect 9484 23675 9542 23681
rect 10502 23672 10508 23684
rect 10560 23672 10566 23724
rect 10594 23672 10600 23724
rect 10652 23712 10658 23724
rect 10689 23715 10747 23721
rect 10689 23712 10701 23715
rect 10652 23684 10701 23712
rect 10652 23672 10658 23684
rect 10689 23681 10701 23684
rect 10735 23681 10747 23715
rect 10689 23675 10747 23681
rect 11422 23672 11428 23724
rect 11480 23712 11486 23724
rect 11701 23715 11759 23721
rect 11701 23712 11713 23715
rect 11480 23684 11713 23712
rect 11480 23672 11486 23684
rect 11701 23681 11713 23684
rect 11747 23681 11759 23715
rect 11701 23675 11759 23681
rect 4120 23616 4568 23644
rect 4120 23604 4126 23616
rect 9214 23604 9220 23656
rect 9272 23604 9278 23656
rect 10962 23604 10968 23656
rect 11020 23644 11026 23656
rect 11333 23647 11391 23653
rect 11333 23644 11345 23647
rect 11020 23616 11345 23644
rect 11020 23604 11026 23616
rect 11333 23613 11345 23616
rect 11379 23613 11391 23647
rect 11333 23607 11391 23613
rect 4433 23579 4491 23585
rect 4433 23545 4445 23579
rect 4479 23576 4491 23579
rect 4798 23576 4804 23588
rect 4479 23548 4804 23576
rect 4479 23545 4491 23548
rect 4433 23539 4491 23545
rect 4798 23536 4804 23548
rect 4856 23536 4862 23588
rect 11238 23536 11244 23588
rect 11296 23576 11302 23588
rect 11517 23579 11575 23585
rect 11296 23548 11376 23576
rect 11296 23536 11302 23548
rect 2777 23511 2835 23517
rect 2777 23477 2789 23511
rect 2823 23508 2835 23511
rect 2958 23508 2964 23520
rect 2823 23480 2964 23508
rect 2823 23477 2835 23480
rect 2777 23471 2835 23477
rect 2958 23468 2964 23480
rect 3016 23468 3022 23520
rect 3786 23468 3792 23520
rect 3844 23468 3850 23520
rect 3973 23511 4031 23517
rect 3973 23477 3985 23511
rect 4019 23508 4031 23511
rect 4062 23508 4068 23520
rect 4019 23480 4068 23508
rect 4019 23477 4031 23480
rect 3973 23471 4031 23477
rect 4062 23468 4068 23480
rect 4120 23468 4126 23520
rect 5902 23468 5908 23520
rect 5960 23508 5966 23520
rect 6181 23511 6239 23517
rect 6181 23508 6193 23511
rect 5960 23480 6193 23508
rect 5960 23468 5966 23480
rect 6181 23477 6193 23480
rect 6227 23508 6239 23511
rect 6270 23508 6276 23520
rect 6227 23480 6276 23508
rect 6227 23477 6239 23480
rect 6181 23471 6239 23477
rect 6270 23468 6276 23480
rect 6328 23468 6334 23520
rect 9858 23468 9864 23520
rect 9916 23508 9922 23520
rect 11054 23508 11060 23520
rect 9916 23480 11060 23508
rect 9916 23468 9922 23480
rect 11054 23468 11060 23480
rect 11112 23468 11118 23520
rect 11348 23508 11376 23548
rect 11517 23545 11529 23579
rect 11563 23545 11575 23579
rect 11716 23576 11744 23675
rect 11882 23672 11888 23724
rect 11940 23672 11946 23724
rect 12066 23672 12072 23724
rect 12124 23672 12130 23724
rect 12176 23644 12204 23820
rect 12802 23808 12808 23860
rect 12860 23848 12866 23860
rect 12986 23848 12992 23860
rect 12860 23820 12992 23848
rect 12860 23808 12866 23820
rect 12986 23808 12992 23820
rect 13044 23808 13050 23860
rect 13078 23808 13084 23860
rect 13136 23808 13142 23860
rect 13814 23848 13820 23860
rect 13372 23820 13820 23848
rect 13372 23780 13400 23820
rect 13814 23808 13820 23820
rect 13872 23848 13878 23860
rect 14553 23851 14611 23857
rect 14553 23848 14565 23851
rect 13872 23820 14565 23848
rect 13872 23808 13878 23820
rect 14553 23817 14565 23820
rect 14599 23817 14611 23851
rect 14553 23811 14611 23817
rect 15010 23808 15016 23860
rect 15068 23808 15074 23860
rect 15304 23820 16160 23848
rect 12452 23752 13400 23780
rect 13440 23783 13498 23789
rect 12452 23721 12480 23752
rect 13440 23749 13452 23783
rect 13486 23780 13498 23783
rect 14090 23780 14096 23792
rect 13486 23752 14096 23780
rect 13486 23749 13498 23752
rect 13440 23743 13498 23749
rect 14090 23740 14096 23752
rect 14148 23740 14154 23792
rect 14182 23740 14188 23792
rect 14240 23780 14246 23792
rect 14829 23783 14887 23789
rect 14829 23780 14841 23783
rect 14240 23752 14841 23780
rect 14240 23740 14246 23752
rect 14829 23749 14841 23752
rect 14875 23749 14887 23783
rect 15304 23780 15332 23820
rect 16132 23789 16160 23820
rect 15933 23783 15991 23789
rect 15933 23780 15945 23783
rect 14829 23743 14887 23749
rect 15028 23752 15332 23780
rect 15396 23752 15945 23780
rect 12437 23715 12495 23721
rect 12437 23681 12449 23715
rect 12483 23681 12495 23715
rect 12437 23675 12495 23681
rect 12526 23672 12532 23724
rect 12584 23672 12590 23724
rect 12710 23672 12716 23724
rect 12768 23672 12774 23724
rect 12802 23672 12808 23724
rect 12860 23672 12866 23724
rect 12897 23715 12955 23721
rect 12897 23681 12909 23715
rect 12943 23712 12955 23715
rect 13078 23712 13084 23724
rect 12943 23684 13084 23712
rect 12943 23681 12955 23684
rect 12897 23675 12955 23681
rect 13078 23672 13084 23684
rect 13136 23672 13142 23724
rect 14645 23715 14703 23721
rect 14645 23681 14657 23715
rect 14691 23712 14703 23715
rect 15028 23712 15056 23752
rect 15396 23724 15424 23752
rect 15933 23749 15945 23752
rect 15979 23749 15991 23783
rect 15933 23743 15991 23749
rect 16117 23783 16175 23789
rect 16117 23749 16129 23783
rect 16163 23780 16175 23783
rect 16482 23780 16488 23792
rect 16163 23752 16488 23780
rect 16163 23749 16175 23752
rect 16117 23743 16175 23749
rect 16482 23740 16488 23752
rect 16540 23740 16546 23792
rect 14691 23684 15056 23712
rect 14691 23681 14703 23684
rect 14645 23675 14703 23681
rect 15102 23672 15108 23724
rect 15160 23672 15166 23724
rect 15289 23715 15347 23721
rect 15289 23681 15301 23715
rect 15335 23681 15347 23715
rect 15289 23675 15347 23681
rect 13170 23644 13176 23656
rect 12176 23616 13176 23644
rect 13170 23604 13176 23616
rect 13228 23604 13234 23656
rect 15194 23644 15200 23656
rect 14200 23616 15200 23644
rect 12066 23576 12072 23588
rect 11716 23548 12072 23576
rect 11517 23539 11575 23545
rect 11532 23508 11560 23539
rect 12066 23536 12072 23548
rect 12124 23536 12130 23588
rect 11348 23480 11560 23508
rect 12253 23511 12311 23517
rect 12253 23477 12265 23511
rect 12299 23508 12311 23511
rect 14200 23508 14228 23616
rect 15194 23604 15200 23616
rect 15252 23604 15258 23656
rect 15304 23644 15332 23675
rect 15378 23672 15384 23724
rect 15436 23672 15442 23724
rect 15473 23715 15531 23721
rect 15473 23681 15485 23715
rect 15519 23712 15531 23715
rect 15562 23712 15568 23724
rect 15519 23684 15568 23712
rect 15519 23681 15531 23684
rect 15473 23675 15531 23681
rect 15562 23672 15568 23684
rect 15620 23712 15626 23724
rect 15620 23684 16160 23712
rect 15620 23672 15626 23684
rect 16132 23656 16160 23684
rect 15654 23644 15660 23656
rect 15304 23616 15660 23644
rect 15654 23604 15660 23616
rect 15712 23644 15718 23656
rect 15930 23644 15936 23656
rect 15712 23616 15936 23644
rect 15712 23604 15718 23616
rect 15930 23604 15936 23616
rect 15988 23604 15994 23656
rect 16114 23604 16120 23656
rect 16172 23604 16178 23656
rect 14274 23536 14280 23588
rect 14332 23576 14338 23588
rect 15749 23579 15807 23585
rect 15749 23576 15761 23579
rect 14332 23548 15761 23576
rect 14332 23536 14338 23548
rect 15749 23545 15761 23548
rect 15795 23545 15807 23579
rect 15749 23539 15807 23545
rect 12299 23480 14228 23508
rect 12299 23477 12311 23480
rect 12253 23471 12311 23477
rect 15286 23468 15292 23520
rect 15344 23508 15350 23520
rect 15657 23511 15715 23517
rect 15657 23508 15669 23511
rect 15344 23480 15669 23508
rect 15344 23468 15350 23480
rect 15657 23477 15669 23480
rect 15703 23477 15715 23511
rect 15657 23471 15715 23477
rect 1104 23418 16652 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 16652 23418
rect 1104 23344 16652 23366
rect 1581 23307 1639 23313
rect 1581 23273 1593 23307
rect 1627 23304 1639 23307
rect 1670 23304 1676 23316
rect 1627 23276 1676 23304
rect 1627 23273 1639 23276
rect 1581 23267 1639 23273
rect 1670 23264 1676 23276
rect 1728 23264 1734 23316
rect 2590 23264 2596 23316
rect 2648 23264 2654 23316
rect 2958 23264 2964 23316
rect 3016 23304 3022 23316
rect 3237 23307 3295 23313
rect 3237 23304 3249 23307
rect 3016 23276 3249 23304
rect 3016 23264 3022 23276
rect 3237 23273 3249 23276
rect 3283 23273 3295 23307
rect 3237 23267 3295 23273
rect 8018 23264 8024 23316
rect 8076 23264 8082 23316
rect 8662 23264 8668 23316
rect 8720 23304 8726 23316
rect 9125 23307 9183 23313
rect 9125 23304 9137 23307
rect 8720 23276 9137 23304
rect 8720 23264 8726 23276
rect 9125 23273 9137 23276
rect 9171 23273 9183 23307
rect 10226 23304 10232 23316
rect 9125 23267 9183 23273
rect 9692 23276 10232 23304
rect 2682 23236 2688 23248
rect 1964 23208 2688 23236
rect 1964 23177 1992 23208
rect 2682 23196 2688 23208
rect 2740 23196 2746 23248
rect 3050 23196 3056 23248
rect 3108 23236 3114 23248
rect 3145 23239 3203 23245
rect 3145 23236 3157 23239
rect 3108 23208 3157 23236
rect 3108 23196 3114 23208
rect 3145 23205 3157 23208
rect 3191 23236 3203 23239
rect 3191 23208 3372 23236
rect 3191 23205 3203 23208
rect 3145 23199 3203 23205
rect 3344 23180 3372 23208
rect 1949 23171 2007 23177
rect 1949 23137 1961 23171
rect 1995 23137 2007 23171
rect 1949 23131 2007 23137
rect 2038 23128 2044 23180
rect 2096 23168 2102 23180
rect 2225 23171 2283 23177
rect 2225 23168 2237 23171
rect 2096 23140 2237 23168
rect 2096 23128 2102 23140
rect 2225 23137 2237 23140
rect 2271 23137 2283 23171
rect 2225 23131 2283 23137
rect 3326 23128 3332 23180
rect 3384 23128 3390 23180
rect 7929 23171 7987 23177
rect 7929 23137 7941 23171
rect 7975 23168 7987 23171
rect 8294 23168 8300 23180
rect 7975 23140 8300 23168
rect 7975 23137 7987 23140
rect 7929 23131 7987 23137
rect 8294 23128 8300 23140
rect 8352 23128 8358 23180
rect 9490 23128 9496 23180
rect 9548 23168 9554 23180
rect 9692 23177 9720 23276
rect 10226 23264 10232 23276
rect 10284 23264 10290 23316
rect 10502 23264 10508 23316
rect 10560 23304 10566 23316
rect 10689 23307 10747 23313
rect 10689 23304 10701 23307
rect 10560 23276 10701 23304
rect 10560 23264 10566 23276
rect 10689 23273 10701 23276
rect 10735 23273 10747 23307
rect 10689 23267 10747 23273
rect 11054 23264 11060 23316
rect 11112 23304 11118 23316
rect 11149 23307 11207 23313
rect 11149 23304 11161 23307
rect 11112 23276 11161 23304
rect 11112 23264 11118 23276
rect 11149 23273 11161 23276
rect 11195 23273 11207 23307
rect 11149 23267 11207 23273
rect 11238 23264 11244 23316
rect 11296 23304 11302 23316
rect 11425 23307 11483 23313
rect 11425 23304 11437 23307
rect 11296 23276 11437 23304
rect 11296 23264 11302 23276
rect 11425 23273 11437 23276
rect 11471 23273 11483 23307
rect 11425 23267 11483 23273
rect 11517 23307 11575 23313
rect 11517 23273 11529 23307
rect 11563 23304 11575 23307
rect 11606 23304 11612 23316
rect 11563 23276 11612 23304
rect 11563 23273 11575 23276
rect 11517 23267 11575 23273
rect 11606 23264 11612 23276
rect 11664 23264 11670 23316
rect 11793 23307 11851 23313
rect 11793 23273 11805 23307
rect 11839 23304 11851 23307
rect 11882 23304 11888 23316
rect 11839 23276 11888 23304
rect 11839 23273 11851 23276
rect 11793 23267 11851 23273
rect 11882 23264 11888 23276
rect 11940 23264 11946 23316
rect 12066 23264 12072 23316
rect 12124 23264 12130 23316
rect 13446 23264 13452 23316
rect 13504 23304 13510 23316
rect 13630 23304 13636 23316
rect 13504 23276 13636 23304
rect 13504 23264 13510 23276
rect 13630 23264 13636 23276
rect 13688 23264 13694 23316
rect 15470 23304 15476 23316
rect 14384 23276 15476 23304
rect 12084 23236 12112 23264
rect 13906 23236 13912 23248
rect 11900 23208 12112 23236
rect 12360 23208 13912 23236
rect 9677 23171 9735 23177
rect 9677 23168 9689 23171
rect 9548 23140 9689 23168
rect 9548 23128 9554 23140
rect 9677 23137 9689 23140
rect 9723 23137 9735 23171
rect 9677 23131 9735 23137
rect 10134 23128 10140 23180
rect 10192 23168 10198 23180
rect 10192 23140 11100 23168
rect 10192 23128 10198 23140
rect 1857 23103 1915 23109
rect 1857 23069 1869 23103
rect 1903 23100 1915 23103
rect 2130 23100 2136 23112
rect 1903 23072 2136 23100
rect 1903 23069 1915 23072
rect 1857 23063 1915 23069
rect 2130 23060 2136 23072
rect 2188 23060 2194 23112
rect 2314 23060 2320 23112
rect 2372 23060 2378 23112
rect 2501 23103 2559 23109
rect 2501 23069 2513 23103
rect 2547 23100 2559 23103
rect 2866 23100 2872 23112
rect 2547 23072 2872 23100
rect 2547 23069 2559 23072
rect 2501 23063 2559 23069
rect 2866 23060 2872 23072
rect 2924 23060 2930 23112
rect 2958 23060 2964 23112
rect 3016 23060 3022 23112
rect 3234 23060 3240 23112
rect 3292 23060 3298 23112
rect 3786 23060 3792 23112
rect 3844 23060 3850 23112
rect 3973 23103 4031 23109
rect 3973 23069 3985 23103
rect 4019 23069 4031 23103
rect 3973 23063 4031 23069
rect 4065 23103 4123 23109
rect 4065 23069 4077 23103
rect 4111 23069 4123 23103
rect 4065 23063 4123 23069
rect 1740 23035 1798 23041
rect 1740 23001 1752 23035
rect 1786 23032 1798 23035
rect 2409 23035 2467 23041
rect 2409 23032 2421 23035
rect 1786 23004 2421 23032
rect 1786 23001 1798 23004
rect 1740 22995 1798 23001
rect 2409 23001 2421 23004
rect 2455 23001 2467 23035
rect 3050 23032 3056 23044
rect 2409 22995 2467 23001
rect 2884 23004 3056 23032
rect 2498 22924 2504 22976
rect 2556 22964 2562 22976
rect 2884 22973 2912 23004
rect 3050 22992 3056 23004
rect 3108 22992 3114 23044
rect 3988 23032 4016 23063
rect 3620 23004 4016 23032
rect 4080 23032 4108 23063
rect 4154 23060 4160 23112
rect 4212 23100 4218 23112
rect 4709 23103 4767 23109
rect 4709 23100 4721 23103
rect 4212 23072 4721 23100
rect 4212 23060 4218 23072
rect 4709 23069 4721 23072
rect 4755 23069 4767 23103
rect 4709 23063 4767 23069
rect 6178 23060 6184 23112
rect 6236 23109 6242 23112
rect 6236 23100 6248 23109
rect 6236 23072 6281 23100
rect 6236 23063 6248 23072
rect 6236 23060 6242 23063
rect 6362 23060 6368 23112
rect 6420 23100 6426 23112
rect 6457 23103 6515 23109
rect 6457 23100 6469 23103
rect 6420 23072 6469 23100
rect 6420 23060 6426 23072
rect 6457 23069 6469 23072
rect 6503 23069 6515 23103
rect 6457 23063 6515 23069
rect 8021 23103 8079 23109
rect 8021 23069 8033 23103
rect 8067 23069 8079 23103
rect 8021 23063 8079 23069
rect 8205 23103 8263 23109
rect 8205 23069 8217 23103
rect 8251 23100 8263 23103
rect 8570 23100 8576 23112
rect 8251 23072 8576 23100
rect 8251 23069 8263 23072
rect 8205 23063 8263 23069
rect 4246 23032 4252 23044
rect 4080 23004 4252 23032
rect 3620 22973 3648 23004
rect 4246 22992 4252 23004
rect 4304 23032 4310 23044
rect 4525 23035 4583 23041
rect 4525 23032 4537 23035
rect 4304 23004 4537 23032
rect 4304 22992 4310 23004
rect 4525 23001 4537 23004
rect 4571 23032 4583 23035
rect 7684 23035 7742 23041
rect 4571 23004 4752 23032
rect 4571 23001 4583 23004
rect 4525 22995 4583 23001
rect 4724 22976 4752 23004
rect 7684 23001 7696 23035
rect 7730 23032 7742 23035
rect 8036 23032 8064 23063
rect 8570 23060 8576 23072
rect 8628 23060 8634 23112
rect 9585 23103 9643 23109
rect 9585 23069 9597 23103
rect 9631 23100 9643 23103
rect 9766 23100 9772 23112
rect 9631 23072 9772 23100
rect 9631 23069 9643 23072
rect 9585 23063 9643 23069
rect 9766 23060 9772 23072
rect 9824 23100 9830 23112
rect 9953 23103 10011 23109
rect 9953 23100 9965 23103
rect 9824 23072 9965 23100
rect 9824 23060 9830 23072
rect 9953 23069 9965 23072
rect 9999 23069 10011 23103
rect 9953 23063 10011 23069
rect 10686 23060 10692 23112
rect 10744 23100 10750 23112
rect 10873 23103 10931 23109
rect 10873 23100 10885 23103
rect 10744 23072 10885 23100
rect 10744 23060 10750 23072
rect 10873 23069 10885 23072
rect 10919 23069 10931 23103
rect 10873 23063 10931 23069
rect 10962 23060 10968 23112
rect 11020 23060 11026 23112
rect 11072 23100 11100 23140
rect 11606 23136 11612 23188
rect 11664 23136 11670 23188
rect 11701 23176 11759 23177
rect 11790 23176 11796 23180
rect 11701 23171 11796 23176
rect 11701 23137 11713 23171
rect 11747 23148 11796 23171
rect 11747 23137 11759 23148
rect 11701 23131 11759 23137
rect 11790 23128 11796 23148
rect 11848 23128 11854 23180
rect 11900 23177 11928 23208
rect 11885 23171 11943 23177
rect 11885 23137 11897 23171
rect 11931 23137 11943 23171
rect 11885 23131 11943 23137
rect 12066 23128 12072 23180
rect 12124 23168 12130 23180
rect 12360 23168 12388 23208
rect 13906 23196 13912 23208
rect 13964 23196 13970 23248
rect 12124 23140 12388 23168
rect 12124 23128 12130 23140
rect 11238 23100 11244 23112
rect 11072 23072 11244 23100
rect 11238 23060 11244 23072
rect 11296 23060 11302 23112
rect 11330 23060 11336 23112
rect 11388 23060 11394 23112
rect 11974 23060 11980 23112
rect 12032 23060 12038 23112
rect 12250 23060 12256 23112
rect 12308 23060 12314 23112
rect 12360 23109 12388 23140
rect 12434 23128 12440 23180
rect 12492 23168 12498 23180
rect 12713 23171 12771 23177
rect 12713 23168 12725 23171
rect 12492 23140 12725 23168
rect 12492 23128 12498 23140
rect 12713 23137 12725 23140
rect 12759 23137 12771 23171
rect 12713 23131 12771 23137
rect 12986 23128 12992 23180
rect 13044 23168 13050 23180
rect 13446 23168 13452 23180
rect 13044 23140 13452 23168
rect 13044 23128 13050 23140
rect 13446 23128 13452 23140
rect 13504 23128 13510 23180
rect 12345 23103 12403 23109
rect 12345 23069 12357 23103
rect 12391 23069 12403 23103
rect 12345 23063 12403 23069
rect 12621 23103 12679 23109
rect 12621 23069 12633 23103
rect 12667 23100 12679 23103
rect 12802 23100 12808 23112
rect 12667 23072 12808 23100
rect 12667 23069 12679 23072
rect 12621 23063 12679 23069
rect 12802 23060 12808 23072
rect 12860 23060 12866 23112
rect 14090 23060 14096 23112
rect 14148 23060 14154 23112
rect 14274 23060 14280 23112
rect 14332 23060 14338 23112
rect 14384 23109 14412 23276
rect 15470 23264 15476 23276
rect 15528 23264 15534 23316
rect 14369 23103 14427 23109
rect 14369 23069 14381 23103
rect 14415 23069 14427 23103
rect 14369 23063 14427 23069
rect 14458 23060 14464 23112
rect 14516 23060 14522 23112
rect 14829 23103 14887 23109
rect 14829 23100 14841 23103
rect 14568 23072 14841 23100
rect 8386 23032 8392 23044
rect 7730 23004 7972 23032
rect 8036 23004 8392 23032
rect 7730 23001 7742 23004
rect 7684 22995 7742 23001
rect 2777 22967 2835 22973
rect 2777 22964 2789 22967
rect 2556 22936 2789 22964
rect 2556 22924 2562 22936
rect 2777 22933 2789 22936
rect 2823 22933 2835 22967
rect 2777 22927 2835 22933
rect 2869 22967 2927 22973
rect 2869 22933 2881 22967
rect 2915 22933 2927 22967
rect 2869 22927 2927 22933
rect 3605 22967 3663 22973
rect 3605 22933 3617 22967
rect 3651 22933 3663 22967
rect 3605 22927 3663 22933
rect 4433 22967 4491 22973
rect 4433 22933 4445 22967
rect 4479 22964 4491 22967
rect 4614 22964 4620 22976
rect 4479 22936 4620 22964
rect 4479 22933 4491 22936
rect 4433 22927 4491 22933
rect 4614 22924 4620 22936
rect 4672 22924 4678 22976
rect 4706 22924 4712 22976
rect 4764 22924 4770 22976
rect 4798 22924 4804 22976
rect 4856 22964 4862 22976
rect 4893 22967 4951 22973
rect 4893 22964 4905 22967
rect 4856 22936 4905 22964
rect 4856 22924 4862 22936
rect 4893 22933 4905 22936
rect 4939 22933 4951 22967
rect 4893 22927 4951 22933
rect 5077 22967 5135 22973
rect 5077 22933 5089 22967
rect 5123 22964 5135 22967
rect 5350 22964 5356 22976
rect 5123 22936 5356 22964
rect 5123 22933 5135 22936
rect 5077 22927 5135 22933
rect 5350 22924 5356 22936
rect 5408 22924 5414 22976
rect 6549 22967 6607 22973
rect 6549 22933 6561 22967
rect 6595 22964 6607 22967
rect 6914 22964 6920 22976
rect 6595 22936 6920 22964
rect 6595 22933 6607 22936
rect 6549 22927 6607 22933
rect 6914 22924 6920 22936
rect 6972 22924 6978 22976
rect 7944 22964 7972 23004
rect 8386 22992 8392 23004
rect 8444 22992 8450 23044
rect 12158 23032 12164 23044
rect 9416 23004 12164 23032
rect 9416 22964 9444 23004
rect 12158 22992 12164 23004
rect 12216 22992 12222 23044
rect 12437 23035 12495 23041
rect 12437 23001 12449 23035
rect 12483 23032 12495 23035
rect 12710 23032 12716 23044
rect 12483 23004 12716 23032
rect 12483 23001 12495 23004
rect 12437 22995 12495 23001
rect 12710 22992 12716 23004
rect 12768 22992 12774 23044
rect 13449 23035 13507 23041
rect 13449 23001 13461 23035
rect 13495 23032 13507 23035
rect 13906 23032 13912 23044
rect 13495 23004 13912 23032
rect 13495 23001 13507 23004
rect 13449 22995 13507 23001
rect 13906 22992 13912 23004
rect 13964 23032 13970 23044
rect 14568 23032 14596 23072
rect 14829 23069 14841 23072
rect 14875 23069 14887 23103
rect 14829 23063 14887 23069
rect 13964 23004 14596 23032
rect 14737 23035 14795 23041
rect 13964 22992 13970 23004
rect 14737 23001 14749 23035
rect 14783 23032 14795 23035
rect 15074 23035 15132 23041
rect 15074 23032 15086 23035
rect 14783 23004 15086 23032
rect 14783 23001 14795 23004
rect 14737 22995 14795 23001
rect 15074 23001 15086 23004
rect 15120 23001 15132 23035
rect 15074 22995 15132 23001
rect 7944 22936 9444 22964
rect 9490 22924 9496 22976
rect 9548 22924 9554 22976
rect 10594 22924 10600 22976
rect 10652 22924 10658 22976
rect 11146 22924 11152 22976
rect 11204 22964 11210 22976
rect 11974 22964 11980 22976
rect 11204 22936 11980 22964
rect 11204 22924 11210 22936
rect 11974 22924 11980 22936
rect 12032 22924 12038 22976
rect 12069 22967 12127 22973
rect 12069 22933 12081 22967
rect 12115 22964 12127 22967
rect 13170 22964 13176 22976
rect 12115 22936 13176 22964
rect 12115 22933 12127 22936
rect 12069 22927 12127 22933
rect 13170 22924 13176 22936
rect 13228 22924 13234 22976
rect 13354 22924 13360 22976
rect 13412 22924 13418 22976
rect 14090 22924 14096 22976
rect 14148 22964 14154 22976
rect 14826 22964 14832 22976
rect 14148 22936 14832 22964
rect 14148 22924 14154 22936
rect 14826 22924 14832 22936
rect 14884 22924 14890 22976
rect 15378 22924 15384 22976
rect 15436 22964 15442 22976
rect 16209 22967 16267 22973
rect 16209 22964 16221 22967
rect 15436 22936 16221 22964
rect 15436 22924 15442 22936
rect 16209 22933 16221 22936
rect 16255 22933 16267 22967
rect 16209 22927 16267 22933
rect 1104 22874 16652 22896
rect 1104 22822 4874 22874
rect 4926 22822 4938 22874
rect 4990 22822 5002 22874
rect 5054 22822 5066 22874
rect 5118 22822 5130 22874
rect 5182 22822 16652 22874
rect 1104 22800 16652 22822
rect 2222 22760 2228 22772
rect 1964 22732 2228 22760
rect 1964 22633 1992 22732
rect 2222 22720 2228 22732
rect 2280 22760 2286 22772
rect 2498 22760 2504 22772
rect 2556 22769 2562 22772
rect 2556 22763 2575 22769
rect 2280 22732 2504 22760
rect 2280 22720 2286 22732
rect 2498 22720 2504 22732
rect 2563 22729 2575 22763
rect 2556 22723 2575 22729
rect 2685 22763 2743 22769
rect 2685 22729 2697 22763
rect 2731 22760 2743 22763
rect 2866 22760 2872 22772
rect 2731 22732 2872 22760
rect 2731 22729 2743 22732
rect 2685 22723 2743 22729
rect 2556 22720 2562 22723
rect 2866 22720 2872 22732
rect 2924 22720 2930 22772
rect 3510 22720 3516 22772
rect 3568 22760 3574 22772
rect 3786 22760 3792 22772
rect 3568 22732 3792 22760
rect 3568 22720 3574 22732
rect 3786 22720 3792 22732
rect 3844 22760 3850 22772
rect 3844 22732 6592 22760
rect 3844 22720 3850 22732
rect 2317 22695 2375 22701
rect 2317 22661 2329 22695
rect 2363 22661 2375 22695
rect 2317 22655 2375 22661
rect 1949 22627 2007 22633
rect 1949 22593 1961 22627
rect 1995 22593 2007 22627
rect 1949 22587 2007 22593
rect 2041 22627 2099 22633
rect 2041 22593 2053 22627
rect 2087 22593 2099 22627
rect 2041 22587 2099 22593
rect 2225 22627 2283 22633
rect 2225 22593 2237 22627
rect 2271 22624 2283 22627
rect 2332 22624 2360 22655
rect 5442 22652 5448 22704
rect 5500 22692 5506 22704
rect 6564 22701 6592 22732
rect 9766 22720 9772 22772
rect 9824 22720 9830 22772
rect 11149 22763 11207 22769
rect 11149 22760 11161 22763
rect 10888 22732 11161 22760
rect 6365 22695 6423 22701
rect 6365 22692 6377 22695
rect 5500 22664 6377 22692
rect 5500 22652 5506 22664
rect 6365 22661 6377 22664
rect 6411 22661 6423 22695
rect 6365 22655 6423 22661
rect 6549 22695 6607 22701
rect 6549 22661 6561 22695
rect 6595 22661 6607 22695
rect 8294 22692 8300 22704
rect 6549 22655 6607 22661
rect 6932 22664 8300 22692
rect 3050 22624 3056 22636
rect 2271 22596 3056 22624
rect 2271 22593 2283 22596
rect 2225 22587 2283 22593
rect 2056 22420 2084 22587
rect 3050 22584 3056 22596
rect 3108 22584 3114 22636
rect 3881 22627 3939 22633
rect 3881 22593 3893 22627
rect 3927 22624 3939 22627
rect 4062 22624 4068 22636
rect 3927 22596 4068 22624
rect 3927 22593 3939 22596
rect 3881 22587 3939 22593
rect 4062 22584 4068 22596
rect 4120 22584 4126 22636
rect 4249 22627 4307 22633
rect 4249 22593 4261 22627
rect 4295 22624 4307 22627
rect 4430 22624 4436 22636
rect 4295 22596 4436 22624
rect 4295 22593 4307 22596
rect 4249 22587 4307 22593
rect 4430 22584 4436 22596
rect 4488 22584 4494 22636
rect 4525 22627 4583 22633
rect 4525 22593 4537 22627
rect 4571 22593 4583 22627
rect 4525 22587 4583 22593
rect 2406 22516 2412 22568
rect 2464 22556 2470 22568
rect 3145 22559 3203 22565
rect 3145 22556 3157 22559
rect 2464 22528 3157 22556
rect 2464 22516 2470 22528
rect 3145 22525 3157 22528
rect 3191 22556 3203 22559
rect 3234 22556 3240 22568
rect 3191 22528 3240 22556
rect 3191 22525 3203 22528
rect 3145 22519 3203 22525
rect 3234 22516 3240 22528
rect 3292 22516 3298 22568
rect 4540 22556 4568 22587
rect 4706 22584 4712 22636
rect 4764 22584 4770 22636
rect 5169 22627 5227 22633
rect 5169 22593 5181 22627
rect 5215 22593 5227 22627
rect 5810 22624 5816 22636
rect 5169 22587 5227 22593
rect 5276 22596 5816 22624
rect 4982 22556 4988 22568
rect 3436 22528 4988 22556
rect 2225 22491 2283 22497
rect 2225 22457 2237 22491
rect 2271 22488 2283 22491
rect 2314 22488 2320 22500
rect 2271 22460 2320 22488
rect 2271 22457 2283 22460
rect 2225 22451 2283 22457
rect 2314 22448 2320 22460
rect 2372 22448 2378 22500
rect 3436 22497 3464 22528
rect 4982 22516 4988 22528
rect 5040 22516 5046 22568
rect 3421 22491 3479 22497
rect 3421 22457 3433 22491
rect 3467 22457 3479 22491
rect 4246 22488 4252 22500
rect 3421 22451 3479 22457
rect 4080 22460 4252 22488
rect 2501 22423 2559 22429
rect 2501 22420 2513 22423
rect 2056 22392 2513 22420
rect 2501 22389 2513 22392
rect 2547 22420 2559 22423
rect 3142 22420 3148 22432
rect 2547 22392 3148 22420
rect 2547 22389 2559 22392
rect 2501 22383 2559 22389
rect 3142 22380 3148 22392
rect 3200 22380 3206 22432
rect 4080 22429 4108 22460
rect 4246 22448 4252 22460
rect 4304 22448 4310 22500
rect 4433 22491 4491 22497
rect 4433 22457 4445 22491
rect 4479 22488 4491 22491
rect 4706 22488 4712 22500
rect 4479 22460 4712 22488
rect 4479 22457 4491 22460
rect 4433 22451 4491 22457
rect 4706 22448 4712 22460
rect 4764 22448 4770 22500
rect 5074 22488 5080 22500
rect 4816 22460 5080 22488
rect 4065 22423 4123 22429
rect 4065 22389 4077 22423
rect 4111 22389 4123 22423
rect 4065 22383 4123 22389
rect 4617 22423 4675 22429
rect 4617 22389 4629 22423
rect 4663 22420 4675 22423
rect 4816 22420 4844 22460
rect 5074 22448 5080 22460
rect 5132 22448 5138 22500
rect 5184 22488 5212 22587
rect 5276 22565 5304 22596
rect 5810 22584 5816 22596
rect 5868 22584 5874 22636
rect 5905 22627 5963 22633
rect 5905 22593 5917 22627
rect 5951 22624 5963 22627
rect 6454 22624 6460 22636
rect 5951 22596 6460 22624
rect 5951 22593 5963 22596
rect 5905 22587 5963 22593
rect 6454 22584 6460 22596
rect 6512 22584 6518 22636
rect 6932 22633 6960 22664
rect 8294 22652 8300 22664
rect 8352 22652 8358 22704
rect 8656 22695 8714 22701
rect 8656 22661 8668 22695
rect 8702 22692 8714 22695
rect 10888 22692 10916 22732
rect 11149 22729 11161 22732
rect 11195 22729 11207 22763
rect 11149 22723 11207 22729
rect 12158 22720 12164 22772
rect 12216 22760 12222 22772
rect 12216 22732 13952 22760
rect 12216 22720 12222 22732
rect 8702 22664 10916 22692
rect 8702 22661 8714 22664
rect 8656 22655 8714 22661
rect 11054 22652 11060 22704
rect 11112 22692 11118 22704
rect 13725 22695 13783 22701
rect 13725 22692 13737 22695
rect 11112 22664 13737 22692
rect 11112 22652 11118 22664
rect 13725 22661 13737 22664
rect 13771 22661 13783 22695
rect 13725 22655 13783 22661
rect 6917 22627 6975 22633
rect 6917 22593 6929 22627
rect 6963 22593 6975 22627
rect 6917 22587 6975 22593
rect 7184 22627 7242 22633
rect 7184 22593 7196 22627
rect 7230 22624 7242 22627
rect 8478 22624 8484 22636
rect 7230 22596 8484 22624
rect 7230 22593 7242 22596
rect 7184 22587 7242 22593
rect 8478 22584 8484 22596
rect 8536 22584 8542 22636
rect 10410 22584 10416 22636
rect 10468 22584 10474 22636
rect 10594 22584 10600 22636
rect 10652 22584 10658 22636
rect 10778 22584 10784 22636
rect 10836 22584 10842 22636
rect 10873 22627 10931 22633
rect 10873 22593 10885 22627
rect 10919 22593 10931 22627
rect 10873 22587 10931 22593
rect 5261 22559 5319 22565
rect 5261 22525 5273 22559
rect 5307 22525 5319 22559
rect 5261 22519 5319 22525
rect 5534 22516 5540 22568
rect 5592 22516 5598 22568
rect 5997 22559 6055 22565
rect 5997 22525 6009 22559
rect 6043 22525 6055 22559
rect 5997 22519 6055 22525
rect 6089 22559 6147 22565
rect 6089 22525 6101 22559
rect 6135 22556 6147 22559
rect 6270 22556 6276 22568
rect 6135 22528 6276 22556
rect 6135 22525 6147 22528
rect 6089 22519 6147 22525
rect 5350 22488 5356 22500
rect 5184 22460 5356 22488
rect 5350 22448 5356 22460
rect 5408 22488 5414 22500
rect 6012 22488 6040 22519
rect 6270 22516 6276 22528
rect 6328 22516 6334 22568
rect 8294 22516 8300 22568
rect 8352 22556 8358 22568
rect 8389 22559 8447 22565
rect 8389 22556 8401 22559
rect 8352 22528 8401 22556
rect 8352 22516 8358 22528
rect 8389 22525 8401 22528
rect 8435 22525 8447 22559
rect 10428 22556 10456 22584
rect 8389 22519 8447 22525
rect 9416 22528 10456 22556
rect 6178 22488 6184 22500
rect 5408 22460 6184 22488
rect 5408 22448 5414 22460
rect 6178 22448 6184 22460
rect 6236 22448 6242 22500
rect 4663 22392 4844 22420
rect 4663 22389 4675 22392
rect 4617 22383 4675 22389
rect 4890 22380 4896 22432
rect 4948 22380 4954 22432
rect 5626 22380 5632 22432
rect 5684 22380 5690 22432
rect 8297 22423 8355 22429
rect 8297 22389 8309 22423
rect 8343 22420 8355 22423
rect 9416 22420 9444 22528
rect 10502 22516 10508 22568
rect 10560 22556 10566 22568
rect 10888 22556 10916 22587
rect 10962 22584 10968 22636
rect 11020 22584 11026 22636
rect 11514 22584 11520 22636
rect 11572 22584 11578 22636
rect 12986 22584 12992 22636
rect 13044 22624 13050 22636
rect 13274 22627 13332 22633
rect 13274 22624 13286 22627
rect 13044 22596 13286 22624
rect 13044 22584 13050 22596
rect 13274 22593 13286 22596
rect 13320 22593 13332 22627
rect 13274 22587 13332 22593
rect 13541 22627 13599 22633
rect 13541 22593 13553 22627
rect 13587 22593 13599 22627
rect 13541 22587 13599 22593
rect 13633 22627 13691 22633
rect 13633 22593 13645 22627
rect 13679 22593 13691 22627
rect 13633 22587 13691 22593
rect 13817 22627 13875 22633
rect 13817 22593 13829 22627
rect 13863 22624 13875 22627
rect 13924 22624 13952 22732
rect 15102 22720 15108 22772
rect 15160 22760 15166 22772
rect 15289 22763 15347 22769
rect 15289 22760 15301 22763
rect 15160 22732 15301 22760
rect 15160 22720 15166 22732
rect 15289 22729 15301 22732
rect 15335 22729 15347 22763
rect 15289 22723 15347 22729
rect 15304 22692 15332 22723
rect 16022 22720 16028 22772
rect 16080 22760 16086 22772
rect 16209 22763 16267 22769
rect 16209 22760 16221 22763
rect 16080 22732 16221 22760
rect 16080 22720 16086 22732
rect 16209 22729 16221 22732
rect 16255 22729 16267 22763
rect 16209 22723 16267 22729
rect 15565 22695 15623 22701
rect 15565 22692 15577 22695
rect 15304 22664 15577 22692
rect 15565 22661 15577 22664
rect 15611 22661 15623 22695
rect 15565 22655 15623 22661
rect 15746 22652 15752 22704
rect 15804 22652 15810 22704
rect 15841 22695 15899 22701
rect 15841 22661 15853 22695
rect 15887 22692 15899 22695
rect 16482 22692 16488 22704
rect 15887 22664 16488 22692
rect 15887 22661 15899 22664
rect 15841 22655 15899 22661
rect 16482 22652 16488 22664
rect 16540 22652 16546 22704
rect 13863 22596 13952 22624
rect 14176 22627 14234 22633
rect 13863 22593 13875 22596
rect 13817 22587 13875 22593
rect 14176 22593 14188 22627
rect 14222 22624 14234 22627
rect 14550 22624 14556 22636
rect 14222 22596 14556 22624
rect 14222 22593 14234 22596
rect 14176 22587 14234 22593
rect 10560 22528 10916 22556
rect 10560 22516 10566 22528
rect 9490 22448 9496 22500
rect 9548 22488 9554 22500
rect 12161 22491 12219 22497
rect 12161 22488 12173 22491
rect 9548 22460 12173 22488
rect 9548 22448 9554 22460
rect 12161 22457 12173 22460
rect 12207 22488 12219 22491
rect 12434 22488 12440 22500
rect 12207 22460 12440 22488
rect 12207 22457 12219 22460
rect 12161 22451 12219 22457
rect 12434 22448 12440 22460
rect 12492 22448 12498 22500
rect 8343 22392 9444 22420
rect 8343 22389 8355 22392
rect 8297 22383 8355 22389
rect 9858 22380 9864 22432
rect 9916 22380 9922 22432
rect 10042 22380 10048 22432
rect 10100 22420 10106 22432
rect 11790 22420 11796 22432
rect 10100 22392 11796 22420
rect 10100 22380 10106 22392
rect 11790 22380 11796 22392
rect 11848 22380 11854 22432
rect 13556 22420 13584 22587
rect 13648 22556 13676 22587
rect 14550 22584 14556 22596
rect 14608 22584 14614 22636
rect 16025 22627 16083 22633
rect 16025 22593 16037 22627
rect 16071 22624 16083 22627
rect 16298 22624 16304 22636
rect 16071 22596 16304 22624
rect 16071 22593 16083 22596
rect 16025 22587 16083 22593
rect 16298 22584 16304 22596
rect 16356 22584 16362 22636
rect 13648 22528 13860 22556
rect 13832 22500 13860 22528
rect 13906 22516 13912 22568
rect 13964 22516 13970 22568
rect 13814 22448 13820 22500
rect 13872 22448 13878 22500
rect 13924 22420 13952 22516
rect 15010 22448 15016 22500
rect 15068 22488 15074 22500
rect 15381 22491 15439 22497
rect 15381 22488 15393 22491
rect 15068 22460 15393 22488
rect 15068 22448 15074 22460
rect 15381 22457 15393 22460
rect 15427 22457 15439 22491
rect 15381 22451 15439 22457
rect 14090 22420 14096 22432
rect 13556 22392 14096 22420
rect 14090 22380 14096 22392
rect 14148 22380 14154 22432
rect 1104 22330 16652 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 16652 22330
rect 1104 22256 16652 22278
rect 3326 22176 3332 22228
rect 3384 22176 3390 22228
rect 4430 22176 4436 22228
rect 4488 22216 4494 22228
rect 4982 22216 4988 22228
rect 4488 22188 4988 22216
rect 4488 22176 4494 22188
rect 4982 22176 4988 22188
rect 5040 22176 5046 22228
rect 8297 22219 8355 22225
rect 8297 22185 8309 22219
rect 8343 22216 8355 22219
rect 8386 22216 8392 22228
rect 8343 22188 8392 22216
rect 8343 22185 8355 22188
rect 8297 22179 8355 22185
rect 8386 22176 8392 22188
rect 8444 22176 8450 22228
rect 8478 22176 8484 22228
rect 8536 22216 8542 22228
rect 8941 22219 8999 22225
rect 8941 22216 8953 22219
rect 8536 22188 8953 22216
rect 8536 22176 8542 22188
rect 8941 22185 8953 22188
rect 8987 22185 8999 22219
rect 8941 22179 8999 22185
rect 10321 22219 10379 22225
rect 10321 22185 10333 22219
rect 10367 22216 10379 22219
rect 10778 22216 10784 22228
rect 10367 22188 10784 22216
rect 10367 22185 10379 22188
rect 10321 22179 10379 22185
rect 10778 22176 10784 22188
rect 10836 22176 10842 22228
rect 11606 22176 11612 22228
rect 11664 22216 11670 22228
rect 11977 22219 12035 22225
rect 11977 22216 11989 22219
rect 11664 22188 11989 22216
rect 11664 22176 11670 22188
rect 11977 22185 11989 22188
rect 12023 22185 12035 22219
rect 11977 22179 12035 22185
rect 13446 22176 13452 22228
rect 13504 22216 13510 22228
rect 13541 22219 13599 22225
rect 13541 22216 13553 22219
rect 13504 22188 13553 22216
rect 13504 22176 13510 22188
rect 13541 22185 13553 22188
rect 13587 22185 13599 22219
rect 13541 22179 13599 22185
rect 13630 22176 13636 22228
rect 13688 22176 13694 22228
rect 14366 22176 14372 22228
rect 14424 22216 14430 22228
rect 14918 22216 14924 22228
rect 14424 22188 14924 22216
rect 14424 22176 14430 22188
rect 14918 22176 14924 22188
rect 14976 22176 14982 22228
rect 3344 22148 3372 22176
rect 3252 22120 3372 22148
rect 3605 22151 3663 22157
rect 3252 22021 3280 22120
rect 3605 22117 3617 22151
rect 3651 22148 3663 22151
rect 4338 22148 4344 22160
rect 3651 22120 4344 22148
rect 3651 22117 3663 22120
rect 3605 22111 3663 22117
rect 4338 22108 4344 22120
rect 4396 22148 4402 22160
rect 5074 22148 5080 22160
rect 4396 22120 5080 22148
rect 4396 22108 4402 22120
rect 5074 22108 5080 22120
rect 5132 22108 5138 22160
rect 6362 22108 6368 22160
rect 6420 22148 6426 22160
rect 6420 22120 6960 22148
rect 6420 22108 6426 22120
rect 3326 22040 3332 22092
rect 3384 22040 3390 22092
rect 4614 22080 4620 22092
rect 4356 22052 4620 22080
rect 3237 22015 3295 22021
rect 3237 21981 3249 22015
rect 3283 21981 3295 22015
rect 3237 21975 3295 21981
rect 3970 21972 3976 22024
rect 4028 21972 4034 22024
rect 4121 22015 4179 22021
rect 4121 21981 4133 22015
rect 4167 22012 4179 22015
rect 4356 22012 4384 22052
rect 4614 22040 4620 22052
rect 4672 22040 4678 22092
rect 5810 22040 5816 22092
rect 5868 22080 5874 22092
rect 6932 22089 6960 22120
rect 10594 22108 10600 22160
rect 10652 22148 10658 22160
rect 11882 22148 11888 22160
rect 10652 22120 11888 22148
rect 10652 22108 10658 22120
rect 11882 22108 11888 22120
rect 11940 22148 11946 22160
rect 12986 22148 12992 22160
rect 11940 22120 12388 22148
rect 11940 22108 11946 22120
rect 6917 22083 6975 22089
rect 5868 22052 6684 22080
rect 5868 22040 5874 22052
rect 4167 21984 4384 22012
rect 4479 22015 4537 22021
rect 4167 21981 4179 21984
rect 4121 21975 4179 21981
rect 4479 21981 4491 22015
rect 4525 22012 4537 22015
rect 4798 22012 4804 22024
rect 4525 21984 4804 22012
rect 4525 21981 4537 21984
rect 4479 21975 4537 21981
rect 4798 21972 4804 21984
rect 4856 21972 4862 22024
rect 5442 21972 5448 22024
rect 5500 22012 5506 22024
rect 6362 22012 6368 22024
rect 5500 21984 6368 22012
rect 5500 21972 5506 21984
rect 6362 21972 6368 21984
rect 6420 21972 6426 22024
rect 6656 22021 6684 22052
rect 6917 22049 6929 22083
rect 6963 22049 6975 22083
rect 6917 22043 6975 22049
rect 9398 22040 9404 22092
rect 9456 22080 9462 22092
rect 9493 22083 9551 22089
rect 9493 22080 9505 22083
rect 9456 22052 9505 22080
rect 9456 22040 9462 22052
rect 9493 22049 9505 22052
rect 9539 22049 9551 22083
rect 9493 22043 9551 22049
rect 10410 22040 10416 22092
rect 10468 22080 10474 22092
rect 10505 22083 10563 22089
rect 10505 22080 10517 22083
rect 10468 22052 10517 22080
rect 10468 22040 10474 22052
rect 10505 22049 10517 22052
rect 10551 22049 10563 22083
rect 12066 22080 12072 22092
rect 10505 22043 10563 22049
rect 10704 22052 12072 22080
rect 6641 22015 6699 22021
rect 6641 21981 6653 22015
rect 6687 21981 6699 22015
rect 6641 21975 6699 21981
rect 6822 21972 6828 22024
rect 6880 22012 6886 22024
rect 6880 21984 7788 22012
rect 6880 21972 6886 21984
rect 3878 21904 3884 21956
rect 3936 21944 3942 21956
rect 4249 21947 4307 21953
rect 4249 21944 4261 21947
rect 3936 21916 4261 21944
rect 3936 21904 3942 21916
rect 4249 21913 4261 21916
rect 4295 21913 4307 21947
rect 4249 21907 4307 21913
rect 4341 21947 4399 21953
rect 4341 21913 4353 21947
rect 4387 21944 4399 21947
rect 4706 21944 4712 21956
rect 4387 21916 4712 21944
rect 4387 21913 4399 21916
rect 4341 21907 4399 21913
rect 4706 21904 4712 21916
rect 4764 21904 4770 21956
rect 5629 21947 5687 21953
rect 5629 21913 5641 21947
rect 5675 21944 5687 21947
rect 7006 21944 7012 21956
rect 5675 21916 7012 21944
rect 5675 21913 5687 21916
rect 5629 21907 5687 21913
rect 7006 21904 7012 21916
rect 7064 21904 7070 21956
rect 7184 21947 7242 21953
rect 7184 21913 7196 21947
rect 7230 21944 7242 21947
rect 7558 21944 7564 21956
rect 7230 21916 7564 21944
rect 7230 21913 7242 21916
rect 7184 21907 7242 21913
rect 7558 21904 7564 21916
rect 7616 21904 7622 21956
rect 7760 21944 7788 21984
rect 9306 21972 9312 22024
rect 9364 22012 9370 22024
rect 9769 22015 9827 22021
rect 9769 22012 9781 22015
rect 9364 21984 9781 22012
rect 9364 21972 9370 21984
rect 9769 21981 9781 21984
rect 9815 21981 9827 22015
rect 9769 21975 9827 21981
rect 9861 22015 9919 22021
rect 9861 21981 9873 22015
rect 9907 21981 9919 22015
rect 9861 21975 9919 21981
rect 7834 21944 7840 21956
rect 7760 21916 7840 21944
rect 7834 21904 7840 21916
rect 7892 21904 7898 21956
rect 9490 21904 9496 21956
rect 9548 21944 9554 21956
rect 9876 21944 9904 21975
rect 9950 21972 9956 22024
rect 10008 22012 10014 22024
rect 10045 22015 10103 22021
rect 10045 22012 10057 22015
rect 10008 21984 10057 22012
rect 10008 21972 10014 21984
rect 10045 21981 10057 21984
rect 10091 21981 10103 22015
rect 10045 21975 10103 21981
rect 10137 22015 10195 22021
rect 10137 21981 10149 22015
rect 10183 22012 10195 22015
rect 10318 22012 10324 22024
rect 10183 21984 10324 22012
rect 10183 21981 10195 21984
rect 10137 21975 10195 21981
rect 10318 21972 10324 21984
rect 10376 21972 10382 22024
rect 10704 22021 10732 22052
rect 12066 22040 12072 22052
rect 12124 22040 12130 22092
rect 12360 22089 12388 22120
rect 12912 22120 12992 22148
rect 12345 22083 12403 22089
rect 12345 22049 12357 22083
rect 12391 22049 12403 22083
rect 12345 22043 12403 22049
rect 12434 22040 12440 22092
rect 12492 22040 12498 22092
rect 12912 22089 12940 22120
rect 12986 22108 12992 22120
rect 13044 22148 13050 22160
rect 13648 22148 13676 22176
rect 13044 22120 13676 22148
rect 13044 22108 13050 22120
rect 12897 22083 12955 22089
rect 12897 22049 12909 22083
rect 12943 22049 12955 22083
rect 12897 22043 12955 22049
rect 13081 22083 13139 22089
rect 13081 22049 13093 22083
rect 13127 22080 13139 22083
rect 14182 22080 14188 22092
rect 13127 22052 14188 22080
rect 13127 22049 13139 22052
rect 13081 22043 13139 22049
rect 14182 22040 14188 22052
rect 14240 22040 14246 22092
rect 14274 22040 14280 22092
rect 14332 22080 14338 22092
rect 14734 22080 14740 22092
rect 14332 22052 14740 22080
rect 14332 22040 14338 22052
rect 14734 22040 14740 22052
rect 14792 22040 14798 22092
rect 10689 22015 10747 22021
rect 10689 21981 10701 22015
rect 10735 21981 10747 22015
rect 10689 21975 10747 21981
rect 11698 21972 11704 22024
rect 11756 22012 11762 22024
rect 12161 22015 12219 22021
rect 12161 22012 12173 22015
rect 11756 21984 12173 22012
rect 11756 21972 11762 21984
rect 12161 21981 12173 21984
rect 12207 21981 12219 22015
rect 12161 21975 12219 21981
rect 12250 21972 12256 22024
rect 12308 21972 12314 22024
rect 13173 22015 13231 22021
rect 13173 21981 13185 22015
rect 13219 22012 13231 22015
rect 13354 22012 13360 22024
rect 13219 21984 13360 22012
rect 13219 21981 13231 21984
rect 13173 21975 13231 21981
rect 13354 21972 13360 21984
rect 13412 21972 13418 22024
rect 13909 22015 13967 22021
rect 13909 21981 13921 22015
rect 13955 22012 13967 22015
rect 15102 22012 15108 22024
rect 13955 21984 15108 22012
rect 13955 21981 13967 21984
rect 13909 21975 13967 21981
rect 15102 21972 15108 21984
rect 15160 21972 15166 22024
rect 15378 21972 15384 22024
rect 15436 21972 15442 22024
rect 15657 22015 15715 22021
rect 15657 21981 15669 22015
rect 15703 22012 15715 22015
rect 15930 22012 15936 22024
rect 15703 21984 15936 22012
rect 15703 21981 15715 21984
rect 15657 21975 15715 21981
rect 15930 21972 15936 21984
rect 15988 21972 15994 22024
rect 16022 21972 16028 22024
rect 16080 21972 16086 22024
rect 9548 21916 9904 21944
rect 9548 21904 9554 21916
rect 10226 21904 10232 21956
rect 10284 21944 10290 21956
rect 10965 21947 11023 21953
rect 10965 21944 10977 21947
rect 10284 21916 10977 21944
rect 10284 21904 10290 21916
rect 10965 21913 10977 21916
rect 11011 21913 11023 21947
rect 10965 21907 11023 21913
rect 4614 21836 4620 21888
rect 4672 21836 4678 21888
rect 6730 21836 6736 21888
rect 6788 21836 6794 21888
rect 9122 21836 9128 21888
rect 9180 21876 9186 21888
rect 9309 21879 9367 21885
rect 9309 21876 9321 21879
rect 9180 21848 9321 21876
rect 9180 21836 9186 21848
rect 9309 21845 9321 21848
rect 9355 21845 9367 21879
rect 9309 21839 9367 21845
rect 9401 21879 9459 21885
rect 9401 21845 9413 21879
rect 9447 21876 9459 21879
rect 9858 21876 9864 21888
rect 9447 21848 9864 21876
rect 9447 21845 9459 21848
rect 9401 21839 9459 21845
rect 9858 21836 9864 21848
rect 9916 21836 9922 21888
rect 10778 21836 10784 21888
rect 10836 21876 10842 21888
rect 10873 21879 10931 21885
rect 10873 21876 10885 21879
rect 10836 21848 10885 21876
rect 10836 21836 10842 21848
rect 10873 21845 10885 21848
rect 10919 21845 10931 21879
rect 10980 21876 11008 21907
rect 11514 21904 11520 21956
rect 11572 21944 11578 21956
rect 11793 21947 11851 21953
rect 11793 21944 11805 21947
rect 11572 21916 11805 21944
rect 11572 21904 11578 21916
rect 11793 21913 11805 21916
rect 11839 21944 11851 21947
rect 11974 21944 11980 21956
rect 11839 21916 11980 21944
rect 11839 21913 11851 21916
rect 11793 21907 11851 21913
rect 11974 21904 11980 21916
rect 12032 21904 12038 21956
rect 13262 21944 13268 21956
rect 12406 21916 13268 21944
rect 12406 21876 12434 21916
rect 13262 21904 13268 21916
rect 13320 21944 13326 21956
rect 14093 21947 14151 21953
rect 14093 21944 14105 21947
rect 13320 21916 14105 21944
rect 13320 21904 13326 21916
rect 14093 21913 14105 21916
rect 14139 21913 14151 21947
rect 14093 21907 14151 21913
rect 14458 21904 14464 21956
rect 14516 21944 14522 21956
rect 14829 21947 14887 21953
rect 14829 21944 14841 21947
rect 14516 21916 14841 21944
rect 14516 21904 14522 21916
rect 14829 21913 14841 21916
rect 14875 21913 14887 21947
rect 15286 21944 15292 21956
rect 14829 21907 14887 21913
rect 14936 21916 15292 21944
rect 10980 21848 12434 21876
rect 13725 21879 13783 21885
rect 10873 21839 10931 21845
rect 13725 21845 13737 21879
rect 13771 21876 13783 21879
rect 14936 21876 14964 21916
rect 15286 21904 15292 21916
rect 15344 21904 15350 21956
rect 13771 21848 14964 21876
rect 13771 21845 13783 21848
rect 13725 21839 13783 21845
rect 15194 21836 15200 21888
rect 15252 21836 15258 21888
rect 15838 21836 15844 21888
rect 15896 21836 15902 21888
rect 16206 21836 16212 21888
rect 16264 21836 16270 21888
rect 1104 21786 16652 21808
rect 1104 21734 4874 21786
rect 4926 21734 4938 21786
rect 4990 21734 5002 21786
rect 5054 21734 5066 21786
rect 5118 21734 5130 21786
rect 5182 21734 16652 21786
rect 1104 21712 16652 21734
rect 3602 21672 3608 21684
rect 2976 21644 3608 21672
rect 842 21496 848 21548
rect 900 21536 906 21548
rect 1397 21539 1455 21545
rect 1397 21536 1409 21539
rect 900 21508 1409 21536
rect 900 21496 906 21508
rect 1397 21505 1409 21508
rect 1443 21505 1455 21539
rect 1397 21499 1455 21505
rect 2869 21539 2927 21545
rect 2869 21505 2881 21539
rect 2915 21536 2927 21539
rect 2976 21536 3004 21644
rect 3602 21632 3608 21644
rect 3660 21632 3666 21684
rect 3878 21632 3884 21684
rect 3936 21632 3942 21684
rect 5258 21632 5264 21684
rect 5316 21632 5322 21684
rect 5350 21632 5356 21684
rect 5408 21632 5414 21684
rect 7558 21632 7564 21684
rect 7616 21632 7622 21684
rect 10870 21632 10876 21684
rect 10928 21632 10934 21684
rect 12066 21632 12072 21684
rect 12124 21672 12130 21684
rect 12342 21672 12348 21684
rect 12124 21644 12348 21672
rect 12124 21632 12130 21644
rect 12342 21632 12348 21644
rect 12400 21632 12406 21684
rect 14090 21632 14096 21684
rect 14148 21672 14154 21684
rect 14458 21672 14464 21684
rect 14148 21644 14464 21672
rect 14148 21632 14154 21644
rect 14458 21632 14464 21644
rect 14516 21632 14522 21684
rect 14550 21632 14556 21684
rect 14608 21632 14614 21684
rect 15473 21675 15531 21681
rect 15473 21641 15485 21675
rect 15519 21672 15531 21675
rect 16022 21672 16028 21684
rect 15519 21644 16028 21672
rect 15519 21641 15531 21644
rect 15473 21635 15531 21641
rect 16022 21632 16028 21644
rect 16080 21632 16086 21684
rect 3513 21607 3571 21613
rect 3513 21604 3525 21607
rect 3160 21576 3525 21604
rect 3160 21548 3188 21576
rect 3513 21573 3525 21576
rect 3559 21573 3571 21607
rect 3513 21567 3571 21573
rect 4709 21607 4767 21613
rect 4709 21573 4721 21607
rect 4755 21604 4767 21607
rect 4982 21604 4988 21616
rect 4755 21576 4988 21604
rect 4755 21573 4767 21576
rect 4709 21567 4767 21573
rect 4982 21564 4988 21576
rect 5040 21564 5046 21616
rect 5470 21607 5528 21613
rect 5470 21573 5482 21607
rect 5516 21604 5528 21607
rect 5626 21604 5632 21616
rect 5516 21576 5632 21604
rect 5516 21573 5528 21576
rect 5470 21567 5528 21573
rect 5626 21564 5632 21576
rect 5684 21564 5690 21616
rect 5810 21564 5816 21616
rect 5868 21604 5874 21616
rect 6089 21607 6147 21613
rect 6089 21604 6101 21607
rect 5868 21576 6101 21604
rect 5868 21564 5874 21576
rect 6089 21573 6101 21576
rect 6135 21604 6147 21607
rect 6178 21604 6184 21616
rect 6135 21576 6184 21604
rect 6135 21573 6147 21576
rect 6089 21567 6147 21573
rect 6178 21564 6184 21576
rect 6236 21604 6242 21616
rect 6822 21604 6828 21616
rect 6236 21576 6828 21604
rect 6236 21564 6242 21576
rect 6822 21564 6828 21576
rect 6880 21564 6886 21616
rect 7006 21564 7012 21616
rect 7064 21604 7070 21616
rect 8202 21604 8208 21616
rect 7064 21576 8208 21604
rect 7064 21564 7070 21576
rect 8202 21564 8208 21576
rect 8260 21604 8266 21616
rect 10226 21604 10232 21616
rect 8260 21576 10232 21604
rect 8260 21564 8266 21576
rect 10226 21564 10232 21576
rect 10284 21564 10290 21616
rect 10410 21564 10416 21616
rect 10468 21604 10474 21616
rect 11238 21604 11244 21616
rect 10468 21576 11244 21604
rect 10468 21564 10474 21576
rect 11238 21564 11244 21576
rect 11296 21564 11302 21616
rect 12250 21604 12256 21616
rect 11900 21576 12256 21604
rect 2915 21508 3004 21536
rect 3053 21539 3111 21545
rect 2915 21505 2927 21508
rect 2869 21499 2927 21505
rect 3053 21505 3065 21539
rect 3099 21536 3111 21539
rect 3142 21536 3148 21548
rect 3099 21508 3148 21536
rect 3099 21505 3111 21508
rect 3053 21499 3111 21505
rect 3142 21496 3148 21508
rect 3200 21496 3206 21548
rect 3237 21539 3295 21545
rect 3237 21505 3249 21539
rect 3283 21505 3295 21539
rect 3237 21499 3295 21505
rect 2961 21471 3019 21477
rect 2961 21437 2973 21471
rect 3007 21468 3019 21471
rect 3252 21468 3280 21499
rect 3326 21496 3332 21548
rect 3384 21536 3390 21548
rect 3421 21539 3479 21545
rect 3421 21536 3433 21539
rect 3384 21508 3433 21536
rect 3384 21496 3390 21508
rect 3421 21505 3433 21508
rect 3467 21505 3479 21539
rect 3421 21499 3479 21505
rect 3605 21539 3663 21545
rect 3605 21505 3617 21539
rect 3651 21505 3663 21539
rect 3605 21499 3663 21505
rect 3007 21440 3280 21468
rect 3620 21468 3648 21499
rect 3878 21496 3884 21548
rect 3936 21536 3942 21548
rect 4065 21539 4123 21545
rect 4065 21536 4077 21539
rect 3936 21508 4077 21536
rect 3936 21496 3942 21508
rect 4065 21505 4077 21508
rect 4111 21505 4123 21539
rect 4065 21499 4123 21505
rect 4157 21539 4215 21545
rect 4157 21505 4169 21539
rect 4203 21505 4215 21539
rect 4157 21499 4215 21505
rect 4172 21468 4200 21499
rect 4338 21496 4344 21548
rect 4396 21496 4402 21548
rect 4430 21496 4436 21548
rect 4488 21496 4494 21548
rect 4890 21496 4896 21548
rect 4948 21536 4954 21548
rect 4948 21508 5212 21536
rect 4948 21496 4954 21508
rect 4908 21468 4936 21496
rect 3620 21440 4936 21468
rect 4985 21471 5043 21477
rect 3007 21437 3019 21440
rect 2961 21431 3019 21437
rect 4985 21437 4997 21471
rect 5031 21468 5043 21471
rect 5074 21468 5080 21480
rect 5031 21440 5080 21468
rect 5031 21437 5043 21440
rect 4985 21431 5043 21437
rect 5074 21428 5080 21440
rect 5132 21428 5138 21480
rect 5184 21468 5212 21508
rect 5902 21496 5908 21548
rect 5960 21496 5966 21548
rect 6549 21539 6607 21545
rect 6012 21529 6316 21536
rect 6012 21508 6190 21529
rect 6012 21468 6040 21508
rect 6178 21495 6190 21508
rect 6224 21508 6316 21529
rect 6224 21495 6236 21508
rect 6178 21489 6236 21495
rect 5184 21440 6040 21468
rect 6288 21468 6316 21508
rect 6549 21505 6561 21539
rect 6595 21536 6607 21539
rect 6638 21536 6644 21548
rect 6595 21508 6644 21536
rect 6595 21505 6607 21508
rect 6549 21499 6607 21505
rect 6638 21496 6644 21508
rect 6696 21496 6702 21548
rect 6914 21496 6920 21548
rect 6972 21496 6978 21548
rect 7653 21539 7711 21545
rect 7653 21505 7665 21539
rect 7699 21505 7711 21539
rect 7653 21499 7711 21505
rect 7668 21468 7696 21499
rect 7834 21496 7840 21548
rect 7892 21496 7898 21548
rect 9214 21496 9220 21548
rect 9272 21536 9278 21548
rect 9766 21545 9772 21548
rect 9493 21539 9551 21545
rect 9493 21536 9505 21539
rect 9272 21508 9505 21536
rect 9272 21496 9278 21508
rect 9493 21505 9505 21508
rect 9539 21505 9551 21539
rect 9493 21499 9551 21505
rect 9760 21499 9772 21545
rect 9766 21496 9772 21499
rect 9824 21496 9830 21548
rect 10778 21496 10784 21548
rect 10836 21536 10842 21548
rect 10965 21539 11023 21545
rect 10965 21536 10977 21539
rect 10836 21508 10977 21536
rect 10836 21496 10842 21508
rect 10965 21505 10977 21508
rect 11011 21536 11023 21539
rect 11422 21536 11428 21548
rect 11011 21508 11428 21536
rect 11011 21505 11023 21508
rect 10965 21499 11023 21505
rect 11422 21496 11428 21508
rect 11480 21496 11486 21548
rect 11514 21496 11520 21548
rect 11572 21496 11578 21548
rect 11698 21496 11704 21548
rect 11756 21496 11762 21548
rect 11900 21480 11928 21576
rect 12250 21564 12256 21576
rect 12308 21564 12314 21616
rect 14366 21564 14372 21616
rect 14424 21564 14430 21616
rect 14734 21564 14740 21616
rect 14792 21604 14798 21616
rect 15562 21604 15568 21616
rect 14792 21576 15568 21604
rect 14792 21564 14798 21576
rect 12069 21539 12127 21545
rect 12069 21505 12081 21539
rect 12115 21536 12127 21539
rect 12342 21536 12348 21558
rect 12115 21508 12348 21536
rect 12115 21505 12127 21508
rect 12342 21506 12348 21508
rect 12400 21506 12406 21558
rect 12618 21545 12624 21548
rect 12069 21499 12127 21505
rect 12612 21499 12624 21545
rect 12618 21496 12624 21499
rect 12676 21496 12682 21548
rect 14384 21536 14412 21564
rect 14829 21539 14887 21545
rect 14829 21536 14841 21539
rect 14384 21508 14841 21536
rect 14829 21505 14841 21508
rect 14875 21505 14887 21539
rect 14829 21499 14887 21505
rect 14918 21496 14924 21548
rect 14976 21496 14982 21548
rect 15010 21496 15016 21548
rect 15068 21496 15074 21548
rect 15212 21545 15240 21576
rect 15562 21564 15568 21576
rect 15620 21564 15626 21616
rect 15197 21539 15255 21545
rect 15197 21505 15209 21539
rect 15243 21505 15255 21539
rect 15197 21499 15255 21505
rect 15289 21539 15347 21545
rect 15289 21505 15301 21539
rect 15335 21505 15347 21539
rect 15289 21499 15347 21505
rect 15749 21539 15807 21545
rect 15749 21505 15761 21539
rect 15795 21536 15807 21539
rect 15838 21536 15844 21548
rect 15795 21508 15844 21536
rect 15795 21505 15807 21508
rect 15749 21499 15807 21505
rect 6288 21440 7696 21468
rect 8938 21428 8944 21480
rect 8996 21428 9002 21480
rect 11057 21471 11115 21477
rect 11057 21437 11069 21471
rect 11103 21468 11115 21471
rect 11146 21468 11152 21480
rect 11103 21440 11152 21468
rect 11103 21437 11115 21440
rect 11057 21431 11115 21437
rect 11146 21428 11152 21440
rect 11204 21428 11210 21480
rect 11330 21428 11336 21480
rect 11388 21428 11394 21480
rect 11793 21471 11851 21477
rect 11793 21437 11805 21471
rect 11839 21437 11851 21471
rect 11793 21431 11851 21437
rect 5258 21360 5264 21412
rect 5316 21400 5322 21412
rect 6365 21403 6423 21409
rect 6365 21400 6377 21403
rect 5316 21372 6377 21400
rect 5316 21360 5322 21372
rect 6365 21369 6377 21372
rect 6411 21369 6423 21403
rect 11348 21400 11376 21428
rect 11808 21400 11836 21431
rect 11882 21428 11888 21480
rect 11940 21428 11946 21480
rect 11974 21428 11980 21480
rect 12032 21468 12038 21480
rect 12345 21471 12403 21477
rect 12345 21468 12357 21471
rect 12032 21440 12357 21468
rect 12032 21428 12038 21440
rect 12345 21437 12357 21440
rect 12391 21437 12403 21471
rect 12345 21431 12403 21437
rect 14369 21471 14427 21477
rect 14369 21437 14381 21471
rect 14415 21468 14427 21471
rect 15304 21468 15332 21499
rect 15838 21496 15844 21508
rect 15896 21496 15902 21548
rect 15933 21539 15991 21545
rect 15933 21505 15945 21539
rect 15979 21505 15991 21539
rect 15933 21499 15991 21505
rect 15948 21468 15976 21499
rect 16022 21496 16028 21548
rect 16080 21496 16086 21548
rect 16482 21468 16488 21480
rect 14415 21440 15332 21468
rect 15856 21440 16488 21468
rect 14415 21437 14427 21440
rect 14369 21431 14427 21437
rect 6365 21363 6423 21369
rect 10980 21372 11836 21400
rect 13725 21403 13783 21409
rect 1581 21335 1639 21341
rect 1581 21301 1593 21335
rect 1627 21332 1639 21335
rect 3418 21332 3424 21344
rect 1627 21304 3424 21332
rect 1627 21301 1639 21304
rect 1581 21295 1639 21301
rect 3418 21292 3424 21304
rect 3476 21292 3482 21344
rect 3789 21335 3847 21341
rect 3789 21301 3801 21335
rect 3835 21332 3847 21335
rect 3878 21332 3884 21344
rect 3835 21304 3884 21332
rect 3835 21301 3847 21304
rect 3789 21295 3847 21301
rect 3878 21292 3884 21304
rect 3936 21292 3942 21344
rect 4525 21335 4583 21341
rect 4525 21301 4537 21335
rect 4571 21332 4583 21335
rect 4706 21332 4712 21344
rect 4571 21304 4712 21332
rect 4571 21301 4583 21304
rect 4525 21295 4583 21301
rect 4706 21292 4712 21304
rect 4764 21292 4770 21344
rect 5626 21292 5632 21344
rect 5684 21292 5690 21344
rect 5721 21335 5779 21341
rect 5721 21301 5733 21335
rect 5767 21332 5779 21335
rect 5810 21332 5816 21344
rect 5767 21304 5816 21332
rect 5767 21301 5779 21304
rect 5721 21295 5779 21301
rect 5810 21292 5816 21304
rect 5868 21292 5874 21344
rect 6546 21292 6552 21344
rect 6604 21332 6610 21344
rect 7653 21335 7711 21341
rect 7653 21332 7665 21335
rect 6604 21304 7665 21332
rect 6604 21292 6610 21304
rect 7653 21301 7665 21304
rect 7699 21301 7711 21335
rect 7653 21295 7711 21301
rect 8662 21292 8668 21344
rect 8720 21332 8726 21344
rect 9490 21332 9496 21344
rect 8720 21304 9496 21332
rect 8720 21292 8726 21304
rect 9490 21292 9496 21304
rect 9548 21332 9554 21344
rect 10980 21341 11008 21372
rect 13725 21369 13737 21403
rect 13771 21400 13783 21403
rect 14384 21400 14412 21431
rect 15856 21412 15884 21440
rect 16482 21428 16488 21440
rect 16540 21428 16546 21480
rect 13771 21372 14412 21400
rect 13771 21369 13783 21372
rect 13725 21363 13783 21369
rect 15378 21360 15384 21412
rect 15436 21400 15442 21412
rect 15565 21403 15623 21409
rect 15565 21400 15577 21403
rect 15436 21372 15577 21400
rect 15436 21360 15442 21372
rect 15565 21369 15577 21372
rect 15611 21369 15623 21403
rect 15565 21363 15623 21369
rect 15838 21360 15844 21412
rect 15896 21360 15902 21412
rect 10965 21335 11023 21341
rect 10965 21332 10977 21335
rect 9548 21304 10977 21332
rect 9548 21292 9554 21304
rect 10965 21301 10977 21304
rect 11011 21301 11023 21335
rect 10965 21295 11023 21301
rect 11333 21335 11391 21341
rect 11333 21301 11345 21335
rect 11379 21332 11391 21335
rect 11882 21332 11888 21344
rect 11379 21304 11888 21332
rect 11379 21301 11391 21304
rect 11333 21295 11391 21301
rect 11882 21292 11888 21304
rect 11940 21292 11946 21344
rect 12253 21335 12311 21341
rect 12253 21301 12265 21335
rect 12299 21332 12311 21335
rect 13262 21332 13268 21344
rect 12299 21304 13268 21332
rect 12299 21301 12311 21304
rect 12253 21295 12311 21301
rect 13262 21292 13268 21304
rect 13320 21292 13326 21344
rect 13814 21292 13820 21344
rect 13872 21292 13878 21344
rect 14274 21292 14280 21344
rect 14332 21332 14338 21344
rect 14918 21332 14924 21344
rect 14332 21304 14924 21332
rect 14332 21292 14338 21304
rect 14918 21292 14924 21304
rect 14976 21292 14982 21344
rect 16209 21335 16267 21341
rect 16209 21301 16221 21335
rect 16255 21332 16267 21335
rect 16298 21332 16304 21344
rect 16255 21304 16304 21332
rect 16255 21301 16267 21304
rect 16209 21295 16267 21301
rect 16298 21292 16304 21304
rect 16356 21292 16362 21344
rect 1104 21242 16652 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 16652 21242
rect 1104 21168 16652 21190
rect 3326 21088 3332 21140
rect 3384 21088 3390 21140
rect 3786 21088 3792 21140
rect 3844 21088 3850 21140
rect 6181 21131 6239 21137
rect 4264 21100 5028 21128
rect 2038 21020 2044 21072
rect 2096 21060 2102 21072
rect 2225 21063 2283 21069
rect 2225 21060 2237 21063
rect 2096 21032 2237 21060
rect 2096 21020 2102 21032
rect 2225 21029 2237 21032
rect 2271 21060 2283 21063
rect 2271 21032 3096 21060
rect 2271 21029 2283 21032
rect 2225 21023 2283 21029
rect 1673 20995 1731 21001
rect 1673 20961 1685 20995
rect 1719 20992 1731 20995
rect 2130 20992 2136 21004
rect 1719 20964 2136 20992
rect 1719 20961 1731 20964
rect 1673 20955 1731 20961
rect 2130 20952 2136 20964
rect 2188 20992 2194 21004
rect 2685 20995 2743 21001
rect 2685 20992 2697 20995
rect 2188 20964 2697 20992
rect 2188 20952 2194 20964
rect 2685 20961 2697 20964
rect 2731 20961 2743 20995
rect 2685 20955 2743 20961
rect 2774 20952 2780 21004
rect 2832 20952 2838 21004
rect 3068 21001 3096 21032
rect 3053 20995 3111 21001
rect 3053 20961 3065 20995
rect 3099 20992 3111 20995
rect 3099 20964 3556 20992
rect 3099 20961 3111 20964
rect 3053 20955 3111 20961
rect 1765 20927 1823 20933
rect 1765 20893 1777 20927
rect 1811 20924 1823 20927
rect 2406 20924 2412 20936
rect 1811 20896 2412 20924
rect 1811 20893 1823 20896
rect 1765 20887 1823 20893
rect 2406 20884 2412 20896
rect 2464 20884 2470 20936
rect 2568 20927 2626 20933
rect 2568 20893 2580 20927
rect 2614 20893 2626 20927
rect 2568 20887 2626 20893
rect 2222 20816 2228 20868
rect 2280 20816 2286 20868
rect 2583 20856 2611 20887
rect 2866 20884 2872 20936
rect 2924 20924 2930 20936
rect 3145 20927 3203 20933
rect 3145 20924 3157 20927
rect 2924 20896 3157 20924
rect 2924 20884 2930 20896
rect 3145 20893 3157 20896
rect 3191 20893 3203 20927
rect 3145 20887 3203 20893
rect 3299 20927 3357 20933
rect 3299 20893 3311 20927
rect 3345 20924 3357 20927
rect 3418 20924 3424 20936
rect 3345 20896 3424 20924
rect 3345 20893 3357 20896
rect 3299 20887 3357 20893
rect 3418 20884 3424 20896
rect 3476 20884 3482 20936
rect 2958 20856 2964 20868
rect 2583 20828 2964 20856
rect 2958 20816 2964 20828
rect 3016 20816 3022 20868
rect 3528 20856 3556 20964
rect 3970 20927 4028 20933
rect 3970 20893 3982 20927
rect 4016 20924 4028 20927
rect 4264 20924 4292 21100
rect 5000 21072 5028 21100
rect 6181 21097 6193 21131
rect 6227 21128 6239 21131
rect 7282 21128 7288 21140
rect 6227 21100 7288 21128
rect 6227 21097 6239 21100
rect 6181 21091 6239 21097
rect 7282 21088 7288 21100
rect 7340 21088 7346 21140
rect 8297 21131 8355 21137
rect 8297 21097 8309 21131
rect 8343 21128 8355 21131
rect 8478 21128 8484 21140
rect 8343 21100 8484 21128
rect 8343 21097 8355 21100
rect 8297 21091 8355 21097
rect 8478 21088 8484 21100
rect 8536 21088 8542 21140
rect 9766 21088 9772 21140
rect 9824 21088 9830 21140
rect 10781 21131 10839 21137
rect 10781 21097 10793 21131
rect 10827 21128 10839 21131
rect 11698 21128 11704 21140
rect 10827 21100 11704 21128
rect 10827 21097 10839 21100
rect 10781 21091 10839 21097
rect 11698 21088 11704 21100
rect 11756 21088 11762 21140
rect 12342 21088 12348 21140
rect 12400 21088 12406 21140
rect 12618 21088 12624 21140
rect 12676 21128 12682 21140
rect 12713 21131 12771 21137
rect 12713 21128 12725 21131
rect 12676 21100 12725 21128
rect 12676 21088 12682 21100
rect 12713 21097 12725 21100
rect 12759 21097 12771 21131
rect 12713 21091 12771 21097
rect 13722 21088 13728 21140
rect 13780 21128 13786 21140
rect 15102 21128 15108 21140
rect 13780 21100 15108 21128
rect 13780 21088 13786 21100
rect 15102 21088 15108 21100
rect 15160 21088 15166 21140
rect 4798 21060 4804 21072
rect 4448 21032 4804 21060
rect 4448 21001 4476 21032
rect 4798 21020 4804 21032
rect 4856 21020 4862 21072
rect 4982 21020 4988 21072
rect 5040 21060 5046 21072
rect 6270 21060 6276 21072
rect 5040 21032 6276 21060
rect 5040 21020 5046 21032
rect 6270 21020 6276 21032
rect 6328 21020 6334 21072
rect 6362 21020 6368 21072
rect 6420 21060 6426 21072
rect 6420 21032 6960 21060
rect 6420 21020 6426 21032
rect 4433 20995 4491 21001
rect 4433 20961 4445 20995
rect 4479 20961 4491 20995
rect 5074 20992 5080 21004
rect 4433 20955 4491 20961
rect 4632 20964 5080 20992
rect 4016 20896 4292 20924
rect 4016 20893 4028 20896
rect 3970 20887 4028 20893
rect 4338 20884 4344 20936
rect 4396 20884 4402 20936
rect 4522 20884 4528 20936
rect 4580 20884 4586 20936
rect 4632 20856 4660 20964
rect 5074 20952 5080 20964
rect 5132 20992 5138 21004
rect 5537 20995 5595 21001
rect 5537 20992 5549 20995
rect 5132 20964 5549 20992
rect 5132 20952 5138 20964
rect 5537 20961 5549 20964
rect 5583 20961 5595 20995
rect 5537 20955 5595 20961
rect 6730 20952 6736 21004
rect 6788 20952 6794 21004
rect 6932 21001 6960 21032
rect 10134 21020 10140 21072
rect 10192 21020 10198 21072
rect 10318 21020 10324 21072
rect 10376 21060 10382 21072
rect 10376 21032 10732 21060
rect 10376 21020 10382 21032
rect 6917 20995 6975 21001
rect 6917 20961 6929 20995
rect 6963 20961 6975 20995
rect 6917 20955 6975 20961
rect 9306 20952 9312 21004
rect 9364 20992 9370 21004
rect 10045 20995 10103 21001
rect 10045 20992 10057 20995
rect 9364 20964 10057 20992
rect 9364 20952 9370 20964
rect 10045 20961 10057 20964
rect 10091 20992 10103 20995
rect 10091 20964 10456 20992
rect 10091 20961 10103 20964
rect 10045 20955 10103 20961
rect 4801 20927 4859 20933
rect 4801 20893 4813 20927
rect 4847 20924 4859 20927
rect 4890 20924 4896 20936
rect 4847 20896 4896 20924
rect 4847 20893 4859 20896
rect 4801 20887 4859 20893
rect 3528 20828 4660 20856
rect 4816 20800 4844 20887
rect 4890 20884 4896 20896
rect 4948 20884 4954 20936
rect 5258 20884 5264 20936
rect 5316 20924 5322 20936
rect 5813 20927 5871 20933
rect 5813 20924 5825 20927
rect 5316 20896 5825 20924
rect 5316 20884 5322 20896
rect 5813 20893 5825 20896
rect 5859 20893 5871 20927
rect 5813 20887 5871 20893
rect 6454 20884 6460 20936
rect 6512 20924 6518 20936
rect 6641 20927 6699 20933
rect 6641 20924 6653 20927
rect 6512 20896 6653 20924
rect 6512 20884 6518 20896
rect 6641 20893 6653 20896
rect 6687 20893 6699 20927
rect 6641 20887 6699 20893
rect 8294 20884 8300 20936
rect 8352 20924 8358 20936
rect 8938 20924 8944 20936
rect 8352 20896 8944 20924
rect 8352 20884 8358 20896
rect 8938 20884 8944 20896
rect 8996 20884 9002 20936
rect 9950 20884 9956 20936
rect 10008 20884 10014 20936
rect 10229 20927 10287 20933
rect 10229 20893 10241 20927
rect 10275 20924 10287 20927
rect 10318 20924 10324 20936
rect 10275 20896 10324 20924
rect 10275 20893 10287 20896
rect 10229 20887 10287 20893
rect 10318 20884 10324 20896
rect 10376 20884 10382 20936
rect 10428 20933 10456 20964
rect 10413 20927 10471 20933
rect 10413 20893 10425 20927
rect 10459 20893 10471 20927
rect 10413 20887 10471 20893
rect 10594 20884 10600 20936
rect 10652 20884 10658 20936
rect 10704 20933 10732 21032
rect 10870 21020 10876 21072
rect 10928 21060 10934 21072
rect 10928 21032 11008 21060
rect 10928 21020 10934 21032
rect 10980 21001 11008 21032
rect 11606 21020 11612 21072
rect 11664 21060 11670 21072
rect 12529 21063 12587 21069
rect 11664 21032 12480 21060
rect 11664 21020 11670 21032
rect 10965 20995 11023 21001
rect 10965 20961 10977 20995
rect 11011 20961 11023 20995
rect 10965 20955 11023 20961
rect 10689 20927 10747 20933
rect 10689 20893 10701 20927
rect 10735 20924 10747 20927
rect 10778 20924 10784 20936
rect 10735 20896 10784 20924
rect 10735 20893 10747 20896
rect 10689 20887 10747 20893
rect 10778 20884 10784 20896
rect 10836 20884 10842 20936
rect 10873 20927 10931 20933
rect 10873 20893 10885 20927
rect 10919 20924 10931 20927
rect 11624 20924 11652 21020
rect 12158 20992 12164 21004
rect 11992 20964 12164 20992
rect 10919 20896 11652 20924
rect 10919 20893 10931 20896
rect 10873 20887 10931 20893
rect 11698 20884 11704 20936
rect 11756 20884 11762 20936
rect 11882 20884 11888 20936
rect 11940 20884 11946 20936
rect 11992 20933 12020 20964
rect 12158 20952 12164 20964
rect 12216 20952 12222 21004
rect 11977 20927 12035 20933
rect 11977 20893 11989 20927
rect 12023 20893 12035 20927
rect 11977 20887 12035 20893
rect 12069 20927 12127 20933
rect 12069 20893 12081 20927
rect 12115 20924 12127 20927
rect 12250 20924 12256 20936
rect 12115 20896 12256 20924
rect 12115 20893 12127 20896
rect 12069 20887 12127 20893
rect 12250 20884 12256 20896
rect 12308 20884 12314 20936
rect 12452 20933 12480 21032
rect 12529 21029 12541 21063
rect 12575 21060 12587 21063
rect 12802 21060 12808 21072
rect 12575 21032 12808 21060
rect 12575 21029 12587 21032
rect 12529 21023 12587 21029
rect 12802 21020 12808 21032
rect 12860 21020 12866 21072
rect 12986 21020 12992 21072
rect 13044 21060 13050 21072
rect 14366 21060 14372 21072
rect 13044 21032 14372 21060
rect 13044 21020 13050 21032
rect 14366 21020 14372 21032
rect 14424 21020 14430 21072
rect 13170 20952 13176 21004
rect 13228 20952 13234 21004
rect 13262 20952 13268 21004
rect 13320 20952 13326 21004
rect 12437 20927 12495 20933
rect 12437 20893 12449 20927
rect 12483 20893 12495 20927
rect 12437 20887 12495 20893
rect 12618 20884 12624 20936
rect 12676 20924 12682 20936
rect 12894 20924 12900 20936
rect 12676 20896 12900 20924
rect 12676 20884 12682 20896
rect 12894 20884 12900 20896
rect 12952 20884 12958 20936
rect 13081 20927 13139 20933
rect 13081 20893 13093 20927
rect 13127 20924 13139 20927
rect 13814 20924 13820 20936
rect 13127 20896 13820 20924
rect 13127 20893 13139 20896
rect 13081 20887 13139 20893
rect 13814 20884 13820 20896
rect 13872 20884 13878 20936
rect 14182 20884 14188 20936
rect 14240 20924 14246 20936
rect 14458 20924 14464 20936
rect 14240 20896 14464 20924
rect 14240 20884 14246 20896
rect 14458 20884 14464 20896
rect 14516 20924 14522 20936
rect 14921 20927 14979 20933
rect 14921 20924 14933 20927
rect 14516 20896 14933 20924
rect 14516 20884 14522 20896
rect 14921 20893 14933 20896
rect 14967 20893 14979 20927
rect 14921 20887 14979 20893
rect 5350 20816 5356 20868
rect 5408 20856 5414 20868
rect 5905 20859 5963 20865
rect 5905 20856 5917 20859
rect 5408 20828 5917 20856
rect 5408 20816 5414 20828
rect 5905 20825 5917 20828
rect 5951 20825 5963 20859
rect 5905 20819 5963 20825
rect 6022 20859 6080 20865
rect 6022 20825 6034 20859
rect 6068 20856 6080 20859
rect 7184 20859 7242 20865
rect 6068 20828 6316 20856
rect 6068 20825 6080 20828
rect 6022 20819 6080 20825
rect 1486 20748 1492 20800
rect 1544 20748 1550 20800
rect 2406 20748 2412 20800
rect 2464 20748 2470 20800
rect 3973 20791 4031 20797
rect 3973 20757 3985 20791
rect 4019 20788 4031 20791
rect 4798 20788 4804 20800
rect 4019 20760 4804 20788
rect 4019 20757 4031 20760
rect 3973 20751 4031 20757
rect 4798 20748 4804 20760
rect 4856 20748 4862 20800
rect 6288 20797 6316 20828
rect 7184 20825 7196 20859
rect 7230 20856 7242 20859
rect 8846 20856 8852 20868
rect 7230 20828 8852 20856
rect 7230 20825 7242 20828
rect 7184 20819 7242 20825
rect 8846 20816 8852 20828
rect 8904 20816 8910 20868
rect 10505 20859 10563 20865
rect 10505 20825 10517 20859
rect 10551 20856 10563 20859
rect 10962 20856 10968 20868
rect 10551 20828 10968 20856
rect 10551 20825 10563 20828
rect 10505 20819 10563 20825
rect 10962 20816 10968 20828
rect 11020 20856 11026 20868
rect 11020 20828 12480 20856
rect 11020 20816 11026 20828
rect 12452 20800 12480 20828
rect 13998 20816 14004 20868
rect 14056 20856 14062 20868
rect 14056 20828 14320 20856
rect 14056 20816 14062 20828
rect 6273 20791 6331 20797
rect 6273 20757 6285 20791
rect 6319 20757 6331 20791
rect 6273 20751 6331 20757
rect 11054 20748 11060 20800
rect 11112 20788 11118 20800
rect 11609 20791 11667 20797
rect 11609 20788 11621 20791
rect 11112 20760 11621 20788
rect 11112 20748 11118 20760
rect 11609 20757 11621 20760
rect 11655 20757 11667 20791
rect 11609 20751 11667 20757
rect 12434 20748 12440 20800
rect 12492 20748 12498 20800
rect 12894 20748 12900 20800
rect 12952 20788 12958 20800
rect 14185 20791 14243 20797
rect 14185 20788 14197 20791
rect 12952 20760 14197 20788
rect 12952 20748 12958 20760
rect 14185 20757 14197 20760
rect 14231 20757 14243 20791
rect 14292 20788 14320 20828
rect 14366 20816 14372 20868
rect 14424 20816 14430 20868
rect 14553 20859 14611 20865
rect 14553 20825 14565 20859
rect 14599 20825 14611 20859
rect 14553 20819 14611 20825
rect 14568 20788 14596 20819
rect 15010 20816 15016 20868
rect 15068 20856 15074 20868
rect 15166 20859 15224 20865
rect 15166 20856 15178 20859
rect 15068 20828 15178 20856
rect 15068 20816 15074 20828
rect 15166 20825 15178 20828
rect 15212 20825 15224 20859
rect 15166 20819 15224 20825
rect 14292 20760 14596 20788
rect 14185 20751 14243 20757
rect 15930 20748 15936 20800
rect 15988 20788 15994 20800
rect 16301 20791 16359 20797
rect 16301 20788 16313 20791
rect 15988 20760 16313 20788
rect 15988 20748 15994 20760
rect 16301 20757 16313 20760
rect 16347 20757 16359 20791
rect 16301 20751 16359 20757
rect 1104 20698 16652 20720
rect 1104 20646 4874 20698
rect 4926 20646 4938 20698
rect 4990 20646 5002 20698
rect 5054 20646 5066 20698
rect 5118 20646 5130 20698
rect 5182 20646 16652 20698
rect 1104 20624 16652 20646
rect 2869 20587 2927 20593
rect 2869 20553 2881 20587
rect 2915 20584 2927 20587
rect 3142 20584 3148 20596
rect 2915 20556 3148 20584
rect 2915 20553 2927 20556
rect 2869 20547 2927 20553
rect 3142 20544 3148 20556
rect 3200 20544 3206 20596
rect 4338 20544 4344 20596
rect 4396 20584 4402 20596
rect 4433 20587 4491 20593
rect 4433 20584 4445 20587
rect 4396 20556 4445 20584
rect 4396 20544 4402 20556
rect 4433 20553 4445 20556
rect 4479 20553 4491 20587
rect 4433 20547 4491 20553
rect 6365 20587 6423 20593
rect 6365 20553 6377 20587
rect 6411 20584 6423 20587
rect 6454 20584 6460 20596
rect 6411 20556 6460 20584
rect 6411 20553 6423 20556
rect 6365 20547 6423 20553
rect 6454 20544 6460 20556
rect 6512 20544 6518 20596
rect 8846 20544 8852 20596
rect 8904 20544 8910 20596
rect 10318 20544 10324 20596
rect 10376 20584 10382 20596
rect 10597 20587 10655 20593
rect 10597 20584 10609 20587
rect 10376 20556 10609 20584
rect 10376 20544 10382 20556
rect 10597 20553 10609 20556
rect 10643 20553 10655 20587
rect 10597 20547 10655 20553
rect 11238 20544 11244 20596
rect 11296 20584 11302 20596
rect 11609 20587 11667 20593
rect 11609 20584 11621 20587
rect 11296 20556 11621 20584
rect 11296 20544 11302 20556
rect 11609 20553 11621 20556
rect 11655 20553 11667 20587
rect 11609 20547 11667 20553
rect 12820 20556 13860 20584
rect 1756 20519 1814 20525
rect 1756 20485 1768 20519
rect 1802 20516 1814 20519
rect 2406 20516 2412 20528
rect 1802 20488 2412 20516
rect 1802 20485 1814 20488
rect 1756 20479 1814 20485
rect 2406 20476 2412 20488
rect 2464 20476 2470 20528
rect 3970 20476 3976 20528
rect 4028 20516 4034 20528
rect 4028 20488 4292 20516
rect 4028 20476 4034 20488
rect 2866 20408 2872 20460
rect 2924 20448 2930 20460
rect 2924 20420 3096 20448
rect 2924 20408 2930 20420
rect 1394 20340 1400 20392
rect 1452 20380 1458 20392
rect 1489 20383 1547 20389
rect 1489 20380 1501 20383
rect 1452 20352 1501 20380
rect 1452 20340 1458 20352
rect 1489 20349 1501 20352
rect 1535 20349 1547 20383
rect 1489 20343 1547 20349
rect 2958 20340 2964 20392
rect 3016 20340 3022 20392
rect 3068 20380 3096 20420
rect 3142 20408 3148 20460
rect 3200 20448 3206 20460
rect 3329 20451 3387 20457
rect 3329 20448 3341 20451
rect 3200 20420 3341 20448
rect 3200 20408 3206 20420
rect 3329 20417 3341 20420
rect 3375 20417 3387 20451
rect 3329 20411 3387 20417
rect 3602 20408 3608 20460
rect 3660 20448 3666 20460
rect 3789 20451 3847 20457
rect 3789 20448 3801 20451
rect 3660 20420 3801 20448
rect 3660 20408 3666 20420
rect 3789 20417 3801 20420
rect 3835 20417 3847 20451
rect 3789 20411 3847 20417
rect 4154 20408 4160 20460
rect 4212 20408 4218 20460
rect 4264 20457 4292 20488
rect 7282 20476 7288 20528
rect 7340 20516 7346 20528
rect 7478 20519 7536 20525
rect 7478 20516 7490 20519
rect 7340 20488 7490 20516
rect 7340 20476 7346 20488
rect 7478 20485 7490 20488
rect 7524 20485 7536 20519
rect 7478 20479 7536 20485
rect 9950 20476 9956 20528
rect 10008 20516 10014 20528
rect 10502 20516 10508 20528
rect 10008 20488 10508 20516
rect 10008 20476 10014 20488
rect 10502 20476 10508 20488
rect 10560 20516 10566 20528
rect 10560 20488 11192 20516
rect 10560 20476 10566 20488
rect 4249 20451 4307 20457
rect 4249 20417 4261 20451
rect 4295 20417 4307 20451
rect 4249 20411 4307 20417
rect 4614 20408 4620 20460
rect 4672 20448 4678 20460
rect 4985 20451 5043 20457
rect 4985 20448 4997 20451
rect 4672 20420 4997 20448
rect 4672 20408 4678 20420
rect 4985 20417 4997 20420
rect 5031 20417 5043 20451
rect 5629 20451 5687 20457
rect 5629 20448 5641 20451
rect 4985 20411 5043 20417
rect 5083 20420 5641 20448
rect 3237 20383 3295 20389
rect 3237 20380 3249 20383
rect 3068 20352 3249 20380
rect 3237 20349 3249 20352
rect 3283 20349 3295 20383
rect 3237 20343 3295 20349
rect 4062 20340 4068 20392
rect 4120 20380 4126 20392
rect 5083 20380 5111 20420
rect 5629 20417 5641 20420
rect 5675 20417 5687 20451
rect 5629 20411 5687 20417
rect 8478 20408 8484 20460
rect 8536 20448 8542 20460
rect 8665 20451 8723 20457
rect 8665 20448 8677 20451
rect 8536 20420 8677 20448
rect 8536 20408 8542 20420
rect 8665 20417 8677 20420
rect 8711 20417 8723 20451
rect 8665 20411 8723 20417
rect 10410 20408 10416 20460
rect 10468 20448 10474 20460
rect 10468 20420 11008 20448
rect 10468 20408 10474 20420
rect 4120 20352 5111 20380
rect 4120 20340 4126 20352
rect 5258 20340 5264 20392
rect 5316 20340 5322 20392
rect 5537 20383 5595 20389
rect 5537 20380 5549 20383
rect 5384 20352 5549 20380
rect 4890 20272 4896 20324
rect 4948 20312 4954 20324
rect 5384 20312 5412 20352
rect 5537 20349 5549 20352
rect 5583 20380 5595 20383
rect 6086 20380 6092 20392
rect 5583 20352 6092 20380
rect 5583 20349 5595 20352
rect 5537 20343 5595 20349
rect 6086 20340 6092 20352
rect 6144 20340 6150 20392
rect 7745 20383 7803 20389
rect 7745 20349 7757 20383
rect 7791 20380 7803 20383
rect 8294 20380 8300 20392
rect 7791 20352 8300 20380
rect 7791 20349 7803 20352
rect 7745 20343 7803 20349
rect 8294 20340 8300 20352
rect 8352 20340 8358 20392
rect 8386 20340 8392 20392
rect 8444 20380 8450 20392
rect 9401 20383 9459 20389
rect 9401 20380 9413 20383
rect 8444 20352 9413 20380
rect 8444 20340 8450 20352
rect 9401 20349 9413 20352
rect 9447 20349 9459 20383
rect 9401 20343 9459 20349
rect 10781 20383 10839 20389
rect 10781 20349 10793 20383
rect 10827 20349 10839 20383
rect 10781 20343 10839 20349
rect 4948 20284 5412 20312
rect 5445 20315 5503 20321
rect 4948 20272 4954 20284
rect 5445 20281 5457 20315
rect 5491 20312 5503 20315
rect 6638 20312 6644 20324
rect 5491 20284 6644 20312
rect 5491 20281 5503 20284
rect 5445 20275 5503 20281
rect 6638 20272 6644 20284
rect 6696 20272 6702 20324
rect 10796 20312 10824 20343
rect 10870 20340 10876 20392
rect 10928 20340 10934 20392
rect 10980 20389 11008 20420
rect 11054 20408 11060 20460
rect 11112 20408 11118 20460
rect 11164 20448 11192 20488
rect 11330 20476 11336 20528
rect 11388 20516 11394 20528
rect 12158 20516 12164 20528
rect 11388 20488 12164 20516
rect 11388 20476 11394 20488
rect 12158 20476 12164 20488
rect 12216 20476 12222 20528
rect 11517 20451 11575 20457
rect 11517 20448 11529 20451
rect 11164 20420 11529 20448
rect 11517 20417 11529 20420
rect 11563 20417 11575 20451
rect 11517 20411 11575 20417
rect 12713 20451 12771 20457
rect 12713 20417 12725 20451
rect 12759 20448 12771 20451
rect 12820 20448 12848 20556
rect 13170 20516 13176 20528
rect 13004 20488 13176 20516
rect 12759 20420 12848 20448
rect 12759 20417 12771 20420
rect 12713 20411 12771 20417
rect 12894 20408 12900 20460
rect 12952 20408 12958 20460
rect 13004 20457 13032 20488
rect 13170 20476 13176 20488
rect 13228 20476 13234 20528
rect 13357 20519 13415 20525
rect 13357 20485 13369 20519
rect 13403 20516 13415 20519
rect 13694 20519 13752 20525
rect 13694 20516 13706 20519
rect 13403 20488 13706 20516
rect 13403 20485 13415 20488
rect 13357 20479 13415 20485
rect 13694 20485 13706 20488
rect 13740 20485 13752 20519
rect 13832 20516 13860 20556
rect 14366 20544 14372 20596
rect 14424 20584 14430 20596
rect 14826 20584 14832 20596
rect 14424 20556 14832 20584
rect 14424 20544 14430 20556
rect 14826 20544 14832 20556
rect 14884 20544 14890 20596
rect 14921 20587 14979 20593
rect 14921 20553 14933 20587
rect 14967 20584 14979 20587
rect 15010 20584 15016 20596
rect 14967 20556 15016 20584
rect 14967 20553 14979 20556
rect 14921 20547 14979 20553
rect 15010 20544 15016 20556
rect 15068 20544 15074 20596
rect 15102 20544 15108 20596
rect 15160 20584 15166 20596
rect 15657 20587 15715 20593
rect 15657 20584 15669 20587
rect 15160 20556 15669 20584
rect 15160 20544 15166 20556
rect 15657 20553 15669 20556
rect 15703 20553 15715 20587
rect 15657 20547 15715 20553
rect 14642 20516 14648 20528
rect 13832 20488 14648 20516
rect 13694 20479 13752 20485
rect 14642 20476 14648 20488
rect 14700 20476 14706 20528
rect 14734 20476 14740 20528
rect 14792 20516 14798 20528
rect 14792 20488 15884 20516
rect 14792 20476 14798 20488
rect 12989 20451 13047 20457
rect 12989 20417 13001 20451
rect 13035 20417 13047 20451
rect 12989 20411 13047 20417
rect 13081 20451 13139 20457
rect 13081 20417 13093 20451
rect 13127 20448 13139 20451
rect 15197 20451 15255 20457
rect 15197 20448 15209 20451
rect 13127 20420 15209 20448
rect 13127 20417 13139 20420
rect 13081 20411 13139 20417
rect 15197 20417 15209 20420
rect 15243 20417 15255 20451
rect 15197 20411 15255 20417
rect 15289 20451 15347 20457
rect 15289 20417 15301 20451
rect 15335 20417 15347 20451
rect 15289 20411 15347 20417
rect 10965 20383 11023 20389
rect 10965 20349 10977 20383
rect 11011 20380 11023 20383
rect 11011 20352 11100 20380
rect 11011 20349 11023 20352
rect 10965 20343 11023 20349
rect 11072 20324 11100 20352
rect 12158 20340 12164 20392
rect 12216 20380 12222 20392
rect 13096 20380 13124 20411
rect 12216 20352 13124 20380
rect 13449 20383 13507 20389
rect 12216 20340 12222 20352
rect 13449 20349 13461 20383
rect 13495 20349 13507 20383
rect 15304 20380 15332 20411
rect 15378 20408 15384 20460
rect 15436 20408 15442 20460
rect 15562 20408 15568 20460
rect 15620 20408 15626 20460
rect 15856 20457 15884 20488
rect 15841 20451 15899 20457
rect 15841 20417 15853 20451
rect 15887 20417 15899 20451
rect 15841 20411 15899 20417
rect 15933 20451 15991 20457
rect 15933 20417 15945 20451
rect 15979 20448 15991 20451
rect 16022 20448 16028 20460
rect 15979 20420 16028 20448
rect 15979 20417 15991 20420
rect 15933 20411 15991 20417
rect 15470 20380 15476 20392
rect 15304 20352 15476 20380
rect 13449 20343 13507 20349
rect 10796 20284 11008 20312
rect 10980 20256 11008 20284
rect 11054 20272 11060 20324
rect 11112 20272 11118 20324
rect 3878 20204 3884 20256
rect 3936 20204 3942 20256
rect 7926 20204 7932 20256
rect 7984 20244 7990 20256
rect 8113 20247 8171 20253
rect 8113 20244 8125 20247
rect 7984 20216 8125 20244
rect 7984 20204 7990 20216
rect 8113 20213 8125 20216
rect 8159 20213 8171 20247
rect 8113 20207 8171 20213
rect 10962 20204 10968 20256
rect 11020 20204 11026 20256
rect 13464 20244 13492 20343
rect 15470 20340 15476 20352
rect 15528 20340 15534 20392
rect 15378 20272 15384 20324
rect 15436 20312 15442 20324
rect 15856 20312 15884 20411
rect 16022 20408 16028 20420
rect 16080 20408 16086 20460
rect 16114 20408 16120 20460
rect 16172 20408 16178 20460
rect 16209 20451 16267 20457
rect 16209 20417 16221 20451
rect 16255 20448 16267 20451
rect 16255 20420 16344 20448
rect 16255 20417 16267 20420
rect 16209 20411 16267 20417
rect 16316 20392 16344 20420
rect 16298 20340 16304 20392
rect 16356 20340 16362 20392
rect 15436 20284 15884 20312
rect 15436 20272 15442 20284
rect 14182 20244 14188 20256
rect 13464 20216 14188 20244
rect 14182 20204 14188 20216
rect 14240 20204 14246 20256
rect 1104 20154 16652 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 16652 20154
rect 1104 20080 16652 20102
rect 1394 20000 1400 20052
rect 1452 20040 1458 20052
rect 1452 20012 3556 20040
rect 1452 20000 1458 20012
rect 2777 19975 2835 19981
rect 2777 19941 2789 19975
rect 2823 19972 2835 19975
rect 2866 19972 2872 19984
rect 2823 19944 2872 19972
rect 2823 19941 2835 19944
rect 2777 19935 2835 19941
rect 2866 19932 2872 19944
rect 2924 19932 2930 19984
rect 3528 19972 3556 20012
rect 3602 20000 3608 20052
rect 3660 20000 3666 20052
rect 4154 20000 4160 20052
rect 4212 20000 4218 20052
rect 4338 20000 4344 20052
rect 4396 20000 4402 20052
rect 4522 20000 4528 20052
rect 4580 20040 4586 20052
rect 4798 20040 4804 20052
rect 4580 20012 4804 20040
rect 4580 20000 4586 20012
rect 4798 20000 4804 20012
rect 4856 20000 4862 20052
rect 6270 20000 6276 20052
rect 6328 20040 6334 20052
rect 6733 20043 6791 20049
rect 6733 20040 6745 20043
rect 6328 20012 6745 20040
rect 6328 20000 6334 20012
rect 6733 20009 6745 20012
rect 6779 20009 6791 20043
rect 6733 20003 6791 20009
rect 8202 20000 8208 20052
rect 8260 20040 8266 20052
rect 8481 20043 8539 20049
rect 8481 20040 8493 20043
rect 8260 20012 8493 20040
rect 8260 20000 8266 20012
rect 8481 20009 8493 20012
rect 8527 20009 8539 20043
rect 8481 20003 8539 20009
rect 10778 20000 10784 20052
rect 10836 20000 10842 20052
rect 11514 20040 11520 20052
rect 11164 20012 11520 20040
rect 8754 19972 8760 19984
rect 3528 19944 5304 19972
rect 1394 19864 1400 19916
rect 1452 19864 1458 19916
rect 2884 19904 2912 19932
rect 3145 19907 3203 19913
rect 3145 19904 3157 19907
rect 2884 19876 3157 19904
rect 3145 19873 3157 19876
rect 3191 19873 3203 19907
rect 4706 19904 4712 19916
rect 3145 19867 3203 19873
rect 3436 19876 4712 19904
rect 1486 19796 1492 19848
rect 1544 19836 1550 19848
rect 3436 19845 3464 19876
rect 4706 19864 4712 19876
rect 4764 19864 4770 19916
rect 4985 19907 5043 19913
rect 4985 19873 4997 19907
rect 5031 19904 5043 19907
rect 5166 19904 5172 19916
rect 5031 19876 5172 19904
rect 5031 19873 5043 19876
rect 4985 19867 5043 19873
rect 5166 19864 5172 19876
rect 5224 19864 5230 19916
rect 1653 19839 1711 19845
rect 1653 19836 1665 19839
rect 1544 19808 1665 19836
rect 1544 19796 1550 19808
rect 1653 19805 1665 19808
rect 1699 19805 1711 19839
rect 1653 19799 1711 19805
rect 3237 19839 3295 19845
rect 3237 19805 3249 19839
rect 3283 19805 3295 19839
rect 3237 19799 3295 19805
rect 3421 19839 3479 19845
rect 3421 19805 3433 19839
rect 3467 19805 3479 19839
rect 3421 19799 3479 19805
rect 3252 19768 3280 19799
rect 4246 19796 4252 19848
rect 4304 19836 4310 19848
rect 4341 19839 4399 19845
rect 4341 19836 4353 19839
rect 4304 19808 4353 19836
rect 4304 19796 4310 19808
rect 4341 19805 4353 19808
rect 4387 19805 4399 19839
rect 4341 19799 4399 19805
rect 4430 19796 4436 19848
rect 4488 19796 4494 19848
rect 4890 19796 4896 19848
rect 4948 19796 4954 19848
rect 5276 19836 5304 19944
rect 8496 19944 8760 19972
rect 8205 19907 8263 19913
rect 8205 19873 8217 19907
rect 8251 19904 8263 19907
rect 8386 19904 8392 19916
rect 8251 19876 8392 19904
rect 8251 19873 8263 19876
rect 8205 19867 8263 19873
rect 8386 19864 8392 19876
rect 8444 19864 8450 19916
rect 8496 19913 8524 19944
rect 8754 19932 8760 19944
rect 8812 19932 8818 19984
rect 9033 19975 9091 19981
rect 9033 19941 9045 19975
rect 9079 19972 9091 19975
rect 9306 19972 9312 19984
rect 9079 19944 9312 19972
rect 9079 19941 9091 19944
rect 9033 19935 9091 19941
rect 8481 19907 8539 19913
rect 8481 19873 8493 19907
rect 8527 19873 8539 19907
rect 8481 19867 8539 19873
rect 8573 19907 8631 19913
rect 8573 19873 8585 19907
rect 8619 19904 8631 19907
rect 9048 19904 9076 19935
rect 9306 19932 9312 19944
rect 9364 19932 9370 19984
rect 10796 19972 10824 20000
rect 11164 19972 11192 20012
rect 11514 20000 11520 20012
rect 11572 20000 11578 20052
rect 12342 20040 12348 20052
rect 11624 20012 12348 20040
rect 10796 19944 11192 19972
rect 8619 19876 9076 19904
rect 9217 19907 9275 19913
rect 8619 19873 8631 19876
rect 8573 19867 8631 19873
rect 9217 19873 9229 19907
rect 9263 19904 9275 19907
rect 9398 19904 9404 19916
rect 9263 19876 9404 19904
rect 9263 19873 9275 19876
rect 9217 19867 9275 19873
rect 9398 19864 9404 19876
rect 9456 19864 9462 19916
rect 11164 19913 11192 19944
rect 11149 19907 11207 19913
rect 11149 19873 11161 19907
rect 11195 19873 11207 19907
rect 11149 19867 11207 19873
rect 11238 19864 11244 19916
rect 11296 19904 11302 19916
rect 11517 19907 11575 19913
rect 11517 19904 11529 19907
rect 11296 19876 11529 19904
rect 11296 19864 11302 19876
rect 11517 19873 11529 19876
rect 11563 19904 11575 19907
rect 11624 19904 11652 20012
rect 12342 20000 12348 20012
rect 12400 20000 12406 20052
rect 14734 20040 14740 20052
rect 14016 20012 14740 20040
rect 11701 19975 11759 19981
rect 11701 19941 11713 19975
rect 11747 19941 11759 19975
rect 11701 19935 11759 19941
rect 11563 19876 11652 19904
rect 11563 19873 11575 19876
rect 11517 19867 11575 19873
rect 5353 19839 5411 19845
rect 5353 19836 5365 19839
rect 5276 19808 5365 19836
rect 5353 19805 5365 19808
rect 5399 19836 5411 19839
rect 5442 19836 5448 19848
rect 5399 19808 5448 19836
rect 5399 19805 5411 19808
rect 5353 19799 5411 19805
rect 5442 19796 5448 19808
rect 5500 19796 5506 19848
rect 5626 19845 5632 19848
rect 5620 19836 5632 19845
rect 5587 19808 5632 19836
rect 5620 19799 5632 19808
rect 5626 19796 5632 19799
rect 5684 19796 5690 19848
rect 7561 19839 7619 19845
rect 7561 19805 7573 19839
rect 7607 19805 7619 19839
rect 7561 19799 7619 19805
rect 7745 19839 7803 19845
rect 7745 19805 7757 19839
rect 7791 19805 7803 19839
rect 7745 19799 7803 19805
rect 4154 19768 4160 19780
rect 3252 19740 4160 19768
rect 4154 19728 4160 19740
rect 4212 19728 4218 19780
rect 4617 19771 4675 19777
rect 4617 19737 4629 19771
rect 4663 19768 4675 19771
rect 5810 19768 5816 19780
rect 4663 19740 5816 19768
rect 4663 19737 4675 19740
rect 4617 19731 4675 19737
rect 5810 19728 5816 19740
rect 5868 19728 5874 19780
rect 3418 19660 3424 19712
rect 3476 19700 3482 19712
rect 4338 19700 4344 19712
rect 3476 19672 4344 19700
rect 3476 19660 3482 19672
rect 4338 19660 4344 19672
rect 4396 19660 4402 19712
rect 5261 19703 5319 19709
rect 5261 19669 5273 19703
rect 5307 19700 5319 19703
rect 5902 19700 5908 19712
rect 5307 19672 5908 19700
rect 5307 19669 5319 19672
rect 5261 19663 5319 19669
rect 5902 19660 5908 19672
rect 5960 19660 5966 19712
rect 7576 19700 7604 19799
rect 7760 19768 7788 19799
rect 7834 19796 7840 19848
rect 7892 19796 7898 19848
rect 7926 19796 7932 19848
rect 7984 19796 7990 19848
rect 8662 19796 8668 19848
rect 8720 19796 8726 19848
rect 8938 19796 8944 19848
rect 8996 19796 9002 19848
rect 9677 19839 9735 19845
rect 9677 19836 9689 19839
rect 9232 19808 9689 19836
rect 9232 19780 9260 19808
rect 9677 19805 9689 19808
rect 9723 19805 9735 19839
rect 9677 19799 9735 19805
rect 9769 19839 9827 19845
rect 9769 19805 9781 19839
rect 9815 19836 9827 19839
rect 9858 19836 9864 19848
rect 9815 19808 9864 19836
rect 9815 19805 9827 19808
rect 9769 19799 9827 19805
rect 9858 19796 9864 19808
rect 9916 19796 9922 19848
rect 9953 19839 10011 19845
rect 9953 19805 9965 19839
rect 9999 19805 10011 19839
rect 9953 19799 10011 19805
rect 8110 19768 8116 19780
rect 7760 19740 8116 19768
rect 8110 19728 8116 19740
rect 8168 19728 8174 19780
rect 8297 19771 8355 19777
rect 8297 19737 8309 19771
rect 8343 19768 8355 19771
rect 8846 19768 8852 19780
rect 8343 19740 8852 19768
rect 8343 19737 8355 19740
rect 8297 19731 8355 19737
rect 8846 19728 8852 19740
rect 8904 19728 8910 19780
rect 9214 19728 9220 19780
rect 9272 19728 9278 19780
rect 9968 19768 9996 19799
rect 10042 19796 10048 19848
rect 10100 19796 10106 19848
rect 10778 19796 10784 19848
rect 10836 19836 10842 19848
rect 11054 19836 11060 19848
rect 10836 19808 11060 19836
rect 10836 19796 10842 19808
rect 11054 19796 11060 19808
rect 11112 19796 11118 19848
rect 11422 19796 11428 19848
rect 11480 19796 11486 19848
rect 11716 19836 11744 19935
rect 12250 19932 12256 19984
rect 12308 19972 12314 19984
rect 12894 19972 12900 19984
rect 12308 19944 12900 19972
rect 12308 19932 12314 19944
rect 12894 19932 12900 19944
rect 12952 19972 12958 19984
rect 13078 19972 13084 19984
rect 12952 19944 13084 19972
rect 12952 19932 12958 19944
rect 13078 19932 13084 19944
rect 13136 19932 13142 19984
rect 11793 19839 11851 19845
rect 11793 19836 11805 19839
rect 11716 19808 11805 19836
rect 11793 19805 11805 19808
rect 11839 19805 11851 19839
rect 11793 19799 11851 19805
rect 12253 19839 12311 19845
rect 12253 19805 12265 19839
rect 12299 19805 12311 19839
rect 12253 19799 12311 19805
rect 13909 19839 13967 19845
rect 13909 19805 13921 19839
rect 13955 19836 13967 19839
rect 14016 19836 14044 20012
rect 14734 20000 14740 20012
rect 14792 20040 14798 20052
rect 15473 20043 15531 20049
rect 15473 20040 15485 20043
rect 14792 20012 15485 20040
rect 14792 20000 14798 20012
rect 15473 20009 15485 20012
rect 15519 20009 15531 20043
rect 15473 20003 15531 20009
rect 16114 20000 16120 20052
rect 16172 20040 16178 20052
rect 16209 20043 16267 20049
rect 16209 20040 16221 20043
rect 16172 20012 16221 20040
rect 16172 20000 16178 20012
rect 16209 20009 16221 20012
rect 16255 20009 16267 20043
rect 16209 20003 16267 20009
rect 16298 19904 16304 19916
rect 15120 19876 16304 19904
rect 13955 19808 14044 19836
rect 14093 19839 14151 19845
rect 13955 19805 13967 19808
rect 13909 19799 13967 19805
rect 14093 19805 14105 19839
rect 14139 19836 14151 19839
rect 14182 19836 14188 19848
rect 14139 19808 14188 19836
rect 14139 19805 14151 19808
rect 14093 19799 14151 19805
rect 10686 19768 10692 19780
rect 9968 19740 10692 19768
rect 10686 19728 10692 19740
rect 10744 19728 10750 19780
rect 11698 19768 11704 19780
rect 11440 19740 11704 19768
rect 11440 19712 11468 19740
rect 11698 19728 11704 19740
rect 11756 19768 11762 19780
rect 12268 19768 12296 19799
rect 14182 19796 14188 19808
rect 14240 19796 14246 19848
rect 15120 19836 15148 19876
rect 16298 19864 16304 19876
rect 16356 19864 16362 19916
rect 14292 19808 15148 19836
rect 11756 19740 12296 19768
rect 11756 19728 11762 19740
rect 13538 19728 13544 19780
rect 13596 19768 13602 19780
rect 14292 19768 14320 19808
rect 15654 19796 15660 19848
rect 15712 19796 15718 19848
rect 15930 19796 15936 19848
rect 15988 19796 15994 19848
rect 16025 19839 16083 19845
rect 16025 19805 16037 19839
rect 16071 19836 16083 19839
rect 16206 19836 16212 19848
rect 16071 19808 16212 19836
rect 16071 19805 16083 19808
rect 16025 19799 16083 19805
rect 16206 19796 16212 19808
rect 16264 19796 16270 19848
rect 14366 19777 14372 19780
rect 13596 19740 14320 19768
rect 13596 19728 13602 19740
rect 14360 19731 14372 19777
rect 14366 19728 14372 19731
rect 14424 19728 14430 19780
rect 15841 19771 15899 19777
rect 15841 19737 15853 19771
rect 15887 19737 15899 19771
rect 15841 19731 15899 19737
rect 8386 19700 8392 19712
rect 7576 19672 8392 19700
rect 8386 19660 8392 19672
rect 8444 19660 8450 19712
rect 9490 19660 9496 19712
rect 9548 19660 9554 19712
rect 10502 19660 10508 19712
rect 10560 19700 10566 19712
rect 11054 19700 11060 19712
rect 10560 19672 11060 19700
rect 10560 19660 10566 19672
rect 11054 19660 11060 19672
rect 11112 19660 11118 19712
rect 11422 19660 11428 19712
rect 11480 19660 11486 19712
rect 11606 19660 11612 19712
rect 11664 19700 11670 19712
rect 11885 19703 11943 19709
rect 11885 19700 11897 19703
rect 11664 19672 11897 19700
rect 11664 19660 11670 19672
rect 11885 19669 11897 19672
rect 11931 19669 11943 19703
rect 11885 19663 11943 19669
rect 11977 19703 12035 19709
rect 11977 19669 11989 19703
rect 12023 19700 12035 19703
rect 13078 19700 13084 19712
rect 12023 19672 13084 19700
rect 12023 19669 12035 19672
rect 11977 19663 12035 19669
rect 13078 19660 13084 19672
rect 13136 19660 13142 19712
rect 13725 19703 13783 19709
rect 13725 19669 13737 19703
rect 13771 19700 13783 19703
rect 15194 19700 15200 19712
rect 13771 19672 15200 19700
rect 13771 19669 13783 19672
rect 13725 19663 13783 19669
rect 15194 19660 15200 19672
rect 15252 19660 15258 19712
rect 15856 19700 15884 19731
rect 16022 19700 16028 19712
rect 15856 19672 16028 19700
rect 16022 19660 16028 19672
rect 16080 19660 16086 19712
rect 1104 19610 16652 19632
rect 1104 19558 4874 19610
rect 4926 19558 4938 19610
rect 4990 19558 5002 19610
rect 5054 19558 5066 19610
rect 5118 19558 5130 19610
rect 5182 19558 16652 19610
rect 1104 19536 16652 19558
rect 3418 19496 3424 19508
rect 2516 19468 3424 19496
rect 2516 19437 2544 19468
rect 3418 19456 3424 19468
rect 3476 19456 3482 19508
rect 4065 19499 4123 19505
rect 4065 19465 4077 19499
rect 4111 19496 4123 19499
rect 4154 19496 4160 19508
rect 4111 19468 4160 19496
rect 4111 19465 4123 19468
rect 4065 19459 4123 19465
rect 4154 19456 4160 19468
rect 4212 19496 4218 19508
rect 4798 19496 4804 19508
rect 4212 19468 4804 19496
rect 4212 19456 4218 19468
rect 4798 19456 4804 19468
rect 4856 19456 4862 19508
rect 5258 19456 5264 19508
rect 5316 19496 5322 19508
rect 5353 19499 5411 19505
rect 5353 19496 5365 19499
rect 5316 19468 5365 19496
rect 5316 19456 5322 19468
rect 5353 19465 5365 19468
rect 5399 19465 5411 19499
rect 5353 19459 5411 19465
rect 5445 19499 5503 19505
rect 5445 19465 5457 19499
rect 5491 19465 5503 19499
rect 6454 19496 6460 19508
rect 5445 19459 5503 19465
rect 5736 19468 6460 19496
rect 2501 19431 2559 19437
rect 2501 19397 2513 19431
rect 2547 19397 2559 19431
rect 3605 19431 3663 19437
rect 3605 19428 3617 19431
rect 2501 19391 2559 19397
rect 2746 19400 3617 19428
rect 1949 19363 2007 19369
rect 1949 19329 1961 19363
rect 1995 19360 2007 19363
rect 2746 19360 2774 19400
rect 3605 19397 3617 19400
rect 3651 19428 3663 19431
rect 3694 19428 3700 19440
rect 3651 19400 3700 19428
rect 3651 19397 3663 19400
rect 3605 19391 3663 19397
rect 1995 19332 2774 19360
rect 2869 19363 2927 19369
rect 1995 19329 2007 19332
rect 1949 19323 2007 19329
rect 2869 19329 2881 19363
rect 2915 19360 2927 19363
rect 3328 19363 3386 19369
rect 3328 19360 3340 19363
rect 2915 19332 3340 19360
rect 2915 19329 2927 19332
rect 2869 19323 2927 19329
rect 3328 19329 3340 19332
rect 3374 19329 3386 19363
rect 3328 19323 3386 19329
rect 3421 19363 3479 19369
rect 3421 19329 3433 19363
rect 3467 19360 3479 19363
rect 3620 19360 3648 19391
rect 3694 19388 3700 19400
rect 3752 19388 3758 19440
rect 3970 19388 3976 19440
rect 4028 19428 4034 19440
rect 5460 19428 5488 19459
rect 5736 19428 5764 19468
rect 6454 19456 6460 19468
rect 6512 19456 6518 19508
rect 8297 19499 8355 19505
rect 8297 19465 8309 19499
rect 8343 19496 8355 19499
rect 8386 19496 8392 19508
rect 8343 19468 8392 19496
rect 8343 19465 8355 19468
rect 8297 19459 8355 19465
rect 8386 19456 8392 19468
rect 8444 19456 8450 19508
rect 10686 19456 10692 19508
rect 10744 19456 10750 19508
rect 10870 19456 10876 19508
rect 10928 19456 10934 19508
rect 11054 19456 11060 19508
rect 11112 19496 11118 19508
rect 11241 19499 11299 19505
rect 11241 19496 11253 19499
rect 11112 19468 11253 19496
rect 11112 19456 11118 19468
rect 11241 19465 11253 19468
rect 11287 19465 11299 19499
rect 11241 19459 11299 19465
rect 11606 19456 11612 19508
rect 11664 19456 11670 19508
rect 12437 19499 12495 19505
rect 12437 19465 12449 19499
rect 12483 19496 12495 19499
rect 12989 19499 13047 19505
rect 12989 19496 13001 19499
rect 12483 19468 13001 19496
rect 12483 19465 12495 19468
rect 12437 19459 12495 19465
rect 12989 19465 13001 19468
rect 13035 19465 13047 19499
rect 12989 19459 13047 19465
rect 14093 19499 14151 19505
rect 14093 19465 14105 19499
rect 14139 19496 14151 19499
rect 14366 19496 14372 19508
rect 14139 19468 14372 19496
rect 14139 19465 14151 19468
rect 14093 19459 14151 19465
rect 14366 19456 14372 19468
rect 14424 19456 14430 19508
rect 14550 19496 14556 19508
rect 14476 19468 14556 19496
rect 4028 19400 5488 19428
rect 5644 19400 5764 19428
rect 4028 19388 4034 19400
rect 4062 19360 4068 19372
rect 3467 19332 4068 19360
rect 3467 19329 3479 19332
rect 3421 19323 3479 19329
rect 2041 19295 2099 19301
rect 2041 19261 2053 19295
rect 2087 19292 2099 19295
rect 2884 19292 2912 19323
rect 2087 19264 2912 19292
rect 3344 19292 3372 19323
rect 4062 19320 4068 19332
rect 4120 19360 4126 19372
rect 4157 19363 4215 19369
rect 4157 19360 4169 19363
rect 4120 19332 4169 19360
rect 4120 19320 4126 19332
rect 4157 19329 4169 19332
rect 4203 19329 4215 19363
rect 4157 19323 4215 19329
rect 4246 19320 4252 19372
rect 4304 19320 4310 19372
rect 4706 19320 4712 19372
rect 4764 19360 4770 19372
rect 4893 19363 4951 19369
rect 4893 19360 4905 19363
rect 4764 19332 4905 19360
rect 4764 19320 4770 19332
rect 4893 19329 4905 19332
rect 4939 19329 4951 19363
rect 4893 19323 4951 19329
rect 5166 19320 5172 19372
rect 5224 19320 5230 19372
rect 5644 19369 5672 19400
rect 5902 19388 5908 19440
rect 5960 19388 5966 19440
rect 5629 19363 5687 19369
rect 5629 19360 5641 19363
rect 5460 19332 5641 19360
rect 3344 19264 4016 19292
rect 2087 19261 2099 19264
rect 2041 19255 2099 19261
rect 3988 19236 4016 19264
rect 4430 19252 4436 19304
rect 4488 19292 4494 19304
rect 5077 19295 5135 19301
rect 5077 19292 5089 19295
rect 4488 19264 5089 19292
rect 4488 19252 4494 19264
rect 5077 19261 5089 19264
rect 5123 19292 5135 19295
rect 5460 19292 5488 19332
rect 5629 19329 5641 19332
rect 5675 19329 5687 19363
rect 5629 19323 5687 19329
rect 5721 19363 5779 19369
rect 5721 19329 5733 19363
rect 5767 19360 5779 19363
rect 5810 19360 5816 19372
rect 5767 19332 5816 19360
rect 5767 19329 5779 19332
rect 5721 19323 5779 19329
rect 5810 19320 5816 19332
rect 5868 19320 5874 19372
rect 7184 19363 7242 19369
rect 7184 19329 7196 19363
rect 7230 19360 7242 19363
rect 7558 19360 7564 19372
rect 7230 19332 7564 19360
rect 7230 19329 7242 19332
rect 7184 19323 7242 19329
rect 7558 19320 7564 19332
rect 7616 19320 7622 19372
rect 8404 19369 8432 19456
rect 8662 19388 8668 19440
rect 8720 19428 8726 19440
rect 8757 19431 8815 19437
rect 8757 19428 8769 19431
rect 8720 19400 8769 19428
rect 8720 19388 8726 19400
rect 8757 19397 8769 19400
rect 8803 19397 8815 19431
rect 8757 19391 8815 19397
rect 9300 19431 9358 19437
rect 9300 19397 9312 19431
rect 9346 19428 9358 19431
rect 9490 19428 9496 19440
rect 9346 19400 9496 19428
rect 9346 19397 9358 19400
rect 9300 19391 9358 19397
rect 9490 19388 9496 19400
rect 9548 19388 9554 19440
rect 11624 19428 11652 19456
rect 10796 19400 11652 19428
rect 12069 19431 12127 19437
rect 8389 19363 8447 19369
rect 8389 19329 8401 19363
rect 8435 19329 8447 19363
rect 8389 19323 8447 19329
rect 10597 19363 10655 19369
rect 10597 19329 10609 19363
rect 10643 19360 10655 19363
rect 10686 19360 10692 19372
rect 10643 19332 10692 19360
rect 10643 19329 10655 19332
rect 10597 19323 10655 19329
rect 10686 19320 10692 19332
rect 10744 19320 10750 19372
rect 10796 19369 10824 19400
rect 12069 19397 12081 19431
rect 12115 19428 12127 19431
rect 12342 19428 12348 19440
rect 12115 19400 12348 19428
rect 12115 19397 12127 19400
rect 12069 19391 12127 19397
rect 12342 19388 12348 19400
rect 12400 19428 12406 19440
rect 12400 19388 12434 19428
rect 13170 19388 13176 19440
rect 13228 19428 13234 19440
rect 13722 19428 13728 19440
rect 13228 19400 13728 19428
rect 13228 19388 13234 19400
rect 13722 19388 13728 19400
rect 13780 19428 13786 19440
rect 14476 19428 14504 19468
rect 14550 19456 14556 19468
rect 14608 19456 14614 19508
rect 14918 19428 14924 19440
rect 13780 19400 14504 19428
rect 13780 19388 13786 19400
rect 10781 19363 10839 19369
rect 10781 19329 10793 19363
rect 10827 19329 10839 19363
rect 10781 19323 10839 19329
rect 11057 19363 11115 19369
rect 11057 19329 11069 19363
rect 11103 19360 11115 19363
rect 11146 19360 11152 19372
rect 11103 19332 11152 19360
rect 11103 19329 11115 19332
rect 11057 19323 11115 19329
rect 11146 19320 11152 19332
rect 11204 19320 11210 19372
rect 11330 19360 11336 19372
rect 11311 19332 11336 19360
rect 11330 19320 11336 19332
rect 11388 19320 11394 19372
rect 11517 19363 11575 19369
rect 11517 19358 11529 19363
rect 11440 19330 11529 19358
rect 5123 19264 5488 19292
rect 5123 19261 5135 19264
rect 5077 19255 5135 19261
rect 6914 19252 6920 19304
rect 6972 19252 6978 19304
rect 8294 19252 8300 19304
rect 8352 19292 8358 19304
rect 9033 19295 9091 19301
rect 9033 19292 9045 19295
rect 8352 19264 9045 19292
rect 8352 19252 8358 19264
rect 9033 19261 9045 19264
rect 9079 19261 9091 19295
rect 9033 19255 9091 19261
rect 10318 19252 10324 19304
rect 10376 19292 10382 19304
rect 11348 19292 11376 19320
rect 10376 19264 11376 19292
rect 10376 19252 10382 19264
rect 3970 19184 3976 19236
rect 4028 19184 4034 19236
rect 4522 19184 4528 19236
rect 4580 19224 4586 19236
rect 4985 19227 5043 19233
rect 4985 19224 4997 19227
rect 4580 19196 4997 19224
rect 4580 19184 4586 19196
rect 4985 19193 4997 19196
rect 5031 19193 5043 19227
rect 4985 19187 5043 19193
rect 10042 19184 10048 19236
rect 10100 19224 10106 19236
rect 10594 19224 10600 19236
rect 10100 19196 10600 19224
rect 10100 19184 10106 19196
rect 10594 19184 10600 19196
rect 10652 19224 10658 19236
rect 11440 19224 11468 19330
rect 11517 19329 11529 19330
rect 11563 19329 11575 19363
rect 11517 19323 11575 19329
rect 11698 19320 11704 19372
rect 11756 19320 11762 19372
rect 11882 19320 11888 19372
rect 11940 19320 11946 19372
rect 12158 19320 12164 19372
rect 12216 19320 12222 19372
rect 12250 19320 12256 19372
rect 12308 19320 12314 19372
rect 12406 19360 12434 19388
rect 12710 19360 12716 19372
rect 12406 19332 12716 19360
rect 12710 19320 12716 19332
rect 12768 19320 12774 19372
rect 14476 19369 14504 19400
rect 14752 19400 14924 19428
rect 12897 19363 12955 19369
rect 12897 19329 12909 19363
rect 12943 19360 12955 19363
rect 13357 19363 13415 19369
rect 13357 19360 13369 19363
rect 12943 19332 13369 19360
rect 12943 19329 12955 19332
rect 12897 19323 12955 19329
rect 13357 19329 13369 19332
rect 13403 19329 13415 19363
rect 14369 19363 14427 19369
rect 14369 19360 14381 19363
rect 13357 19323 13415 19329
rect 14200 19332 14381 19360
rect 13078 19252 13084 19304
rect 13136 19252 13142 19304
rect 13906 19252 13912 19304
rect 13964 19252 13970 19304
rect 10652 19196 11468 19224
rect 14200 19224 14228 19332
rect 14369 19329 14381 19332
rect 14415 19329 14427 19363
rect 14369 19323 14427 19329
rect 14461 19363 14519 19369
rect 14461 19329 14473 19363
rect 14507 19329 14519 19363
rect 14461 19323 14519 19329
rect 14550 19320 14556 19372
rect 14608 19320 14614 19372
rect 14752 19369 14780 19400
rect 14918 19388 14924 19400
rect 14976 19428 14982 19440
rect 15562 19428 15568 19440
rect 14976 19400 15568 19428
rect 14976 19388 14982 19400
rect 15562 19388 15568 19400
rect 15620 19388 15626 19440
rect 14737 19363 14795 19369
rect 14737 19329 14749 19363
rect 14783 19329 14795 19363
rect 14737 19323 14795 19329
rect 15010 19320 15016 19372
rect 15068 19360 15074 19372
rect 15177 19363 15235 19369
rect 15177 19360 15189 19363
rect 15068 19332 15189 19360
rect 15068 19320 15074 19332
rect 15177 19329 15189 19332
rect 15223 19329 15235 19363
rect 15177 19323 15235 19329
rect 14274 19252 14280 19304
rect 14332 19292 14338 19304
rect 14921 19295 14979 19301
rect 14921 19292 14933 19295
rect 14332 19264 14933 19292
rect 14332 19252 14338 19264
rect 14921 19261 14933 19264
rect 14967 19261 14979 19295
rect 14921 19255 14979 19261
rect 14200 19196 14320 19224
rect 10652 19184 10658 19196
rect 2314 19116 2320 19168
rect 2372 19156 2378 19168
rect 2682 19156 2688 19168
rect 2372 19128 2688 19156
rect 2372 19116 2378 19128
rect 2682 19116 2688 19128
rect 2740 19116 2746 19168
rect 3142 19116 3148 19168
rect 3200 19156 3206 19168
rect 3237 19159 3295 19165
rect 3237 19156 3249 19159
rect 3200 19128 3249 19156
rect 3200 19116 3206 19128
rect 3237 19125 3249 19128
rect 3283 19125 3295 19159
rect 3237 19119 3295 19125
rect 4338 19116 4344 19168
rect 4396 19156 4402 19168
rect 4706 19156 4712 19168
rect 4396 19128 4712 19156
rect 4396 19116 4402 19128
rect 4706 19116 4712 19128
rect 4764 19116 4770 19168
rect 5905 19159 5963 19165
rect 5905 19125 5917 19159
rect 5951 19156 5963 19159
rect 6546 19156 6552 19168
rect 5951 19128 6552 19156
rect 5951 19125 5963 19128
rect 5905 19119 5963 19125
rect 6546 19116 6552 19128
rect 6604 19116 6610 19168
rect 6638 19116 6644 19168
rect 6696 19156 6702 19168
rect 8110 19156 8116 19168
rect 6696 19128 8116 19156
rect 6696 19116 6702 19128
rect 8110 19116 8116 19128
rect 8168 19116 8174 19168
rect 8754 19116 8760 19168
rect 8812 19116 8818 19168
rect 8941 19159 8999 19165
rect 8941 19125 8953 19159
rect 8987 19156 8999 19159
rect 9398 19156 9404 19168
rect 8987 19128 9404 19156
rect 8987 19125 8999 19128
rect 8941 19119 8999 19125
rect 9398 19116 9404 19128
rect 9456 19116 9462 19168
rect 9950 19116 9956 19168
rect 10008 19156 10014 19168
rect 10413 19159 10471 19165
rect 10413 19156 10425 19159
rect 10008 19128 10425 19156
rect 10008 19116 10014 19128
rect 10413 19125 10425 19128
rect 10459 19125 10471 19159
rect 10413 19119 10471 19125
rect 12526 19116 12532 19168
rect 12584 19116 12590 19168
rect 14292 19156 14320 19196
rect 15102 19156 15108 19168
rect 14292 19128 15108 19156
rect 15102 19116 15108 19128
rect 15160 19116 15166 19168
rect 15930 19116 15936 19168
rect 15988 19156 15994 19168
rect 16301 19159 16359 19165
rect 16301 19156 16313 19159
rect 15988 19128 16313 19156
rect 15988 19116 15994 19128
rect 16301 19125 16313 19128
rect 16347 19125 16359 19159
rect 16301 19119 16359 19125
rect 1104 19066 16652 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 16652 19066
rect 1104 18992 16652 19014
rect 6104 18924 8524 18952
rect 6104 18757 6132 18924
rect 8496 18816 8524 18924
rect 8846 18912 8852 18964
rect 8904 18952 8910 18964
rect 8941 18955 8999 18961
rect 8941 18952 8953 18955
rect 8904 18924 8953 18952
rect 8904 18912 8910 18924
rect 8941 18921 8953 18924
rect 8987 18921 8999 18955
rect 8941 18915 8999 18921
rect 9030 18912 9036 18964
rect 9088 18952 9094 18964
rect 10042 18952 10048 18964
rect 9088 18924 10048 18952
rect 9088 18912 9094 18924
rect 10042 18912 10048 18924
rect 10100 18912 10106 18964
rect 10137 18955 10195 18961
rect 10137 18921 10149 18955
rect 10183 18952 10195 18955
rect 10318 18952 10324 18964
rect 10183 18924 10324 18952
rect 10183 18921 10195 18924
rect 10137 18915 10195 18921
rect 10318 18912 10324 18924
rect 10376 18912 10382 18964
rect 10689 18955 10747 18961
rect 10689 18921 10701 18955
rect 10735 18952 10747 18955
rect 11698 18952 11704 18964
rect 10735 18924 11704 18952
rect 10735 18921 10747 18924
rect 10689 18915 10747 18921
rect 11698 18912 11704 18924
rect 11756 18912 11762 18964
rect 11882 18912 11888 18964
rect 11940 18912 11946 18964
rect 12618 18952 12624 18964
rect 11992 18924 12624 18952
rect 8570 18844 8576 18896
rect 8628 18884 8634 18896
rect 8665 18887 8723 18893
rect 8665 18884 8677 18887
rect 8628 18856 8677 18884
rect 8628 18844 8634 18856
rect 8665 18853 8677 18856
rect 8711 18884 8723 18887
rect 9766 18884 9772 18896
rect 8711 18856 9772 18884
rect 8711 18853 8723 18856
rect 8665 18847 8723 18853
rect 9766 18844 9772 18856
rect 9824 18844 9830 18896
rect 9950 18844 9956 18896
rect 10008 18844 10014 18896
rect 10505 18887 10563 18893
rect 10505 18853 10517 18887
rect 10551 18853 10563 18887
rect 11146 18884 11152 18896
rect 10505 18847 10563 18853
rect 10796 18856 11152 18884
rect 9309 18819 9367 18825
rect 9309 18816 9321 18819
rect 8496 18788 9321 18816
rect 8496 18760 8524 18788
rect 9309 18785 9321 18788
rect 9355 18785 9367 18819
rect 9309 18779 9367 18785
rect 9674 18776 9680 18828
rect 9732 18816 9738 18828
rect 10520 18816 10548 18847
rect 9732 18788 10548 18816
rect 9732 18776 9738 18788
rect 5905 18751 5963 18757
rect 5905 18717 5917 18751
rect 5951 18717 5963 18751
rect 5905 18711 5963 18717
rect 6089 18751 6147 18757
rect 6089 18717 6101 18751
rect 6135 18717 6147 18751
rect 6089 18711 6147 18717
rect 6273 18751 6331 18757
rect 6273 18717 6285 18751
rect 6319 18717 6331 18751
rect 6273 18711 6331 18717
rect 5920 18680 5948 18711
rect 6288 18680 6316 18711
rect 6914 18708 6920 18760
rect 6972 18748 6978 18760
rect 8294 18748 8300 18760
rect 6972 18720 8300 18748
rect 6972 18708 6978 18720
rect 8294 18708 8300 18720
rect 8352 18708 8358 18760
rect 8478 18708 8484 18760
rect 8536 18708 8542 18760
rect 8757 18751 8815 18757
rect 8757 18717 8769 18751
rect 8803 18748 8815 18751
rect 9490 18748 9496 18760
rect 8803 18720 9496 18748
rect 8803 18717 8815 18720
rect 8757 18711 8815 18717
rect 9490 18708 9496 18720
rect 9548 18708 9554 18760
rect 9582 18708 9588 18760
rect 9640 18708 9646 18760
rect 10410 18708 10416 18760
rect 10468 18748 10474 18760
rect 10796 18748 10824 18856
rect 11146 18844 11152 18856
rect 11204 18844 11210 18896
rect 10870 18776 10876 18828
rect 10928 18816 10934 18828
rect 11333 18819 11391 18825
rect 11333 18816 11345 18819
rect 10928 18788 11345 18816
rect 10928 18776 10934 18788
rect 11333 18785 11345 18788
rect 11379 18785 11391 18819
rect 11333 18779 11391 18785
rect 10468 18720 10824 18748
rect 10965 18751 11023 18757
rect 10468 18708 10474 18720
rect 10965 18717 10977 18751
rect 11011 18717 11023 18751
rect 10965 18711 11023 18717
rect 5920 18652 6316 18680
rect 5994 18572 6000 18624
rect 6052 18572 6058 18624
rect 6288 18612 6316 18652
rect 6825 18683 6883 18689
rect 6825 18649 6837 18683
rect 6871 18680 6883 18683
rect 7006 18680 7012 18692
rect 6871 18652 7012 18680
rect 6871 18649 6883 18652
rect 6825 18643 6883 18649
rect 7006 18640 7012 18652
rect 7064 18680 7070 18692
rect 8052 18683 8110 18689
rect 7064 18652 7880 18680
rect 7064 18640 7070 18652
rect 7852 18624 7880 18652
rect 8052 18649 8064 18683
rect 8098 18680 8110 18683
rect 8202 18680 8208 18692
rect 8098 18652 8208 18680
rect 8098 18649 8110 18652
rect 8052 18643 8110 18649
rect 8202 18640 8208 18652
rect 8260 18640 8266 18692
rect 9122 18689 9128 18692
rect 9100 18683 9128 18689
rect 9100 18649 9112 18683
rect 9180 18680 9186 18692
rect 9306 18680 9312 18692
rect 9180 18652 9312 18680
rect 9100 18643 9128 18649
rect 9122 18640 9128 18643
rect 9180 18640 9186 18652
rect 9306 18640 9312 18652
rect 9364 18640 9370 18692
rect 9950 18640 9956 18692
rect 10008 18680 10014 18692
rect 10229 18683 10287 18689
rect 10229 18680 10241 18683
rect 10008 18652 10241 18680
rect 10008 18640 10014 18652
rect 10229 18649 10241 18652
rect 10275 18649 10287 18683
rect 10229 18643 10287 18649
rect 10594 18640 10600 18692
rect 10652 18680 10658 18692
rect 10980 18680 11008 18711
rect 11054 18708 11060 18760
rect 11112 18748 11118 18760
rect 11149 18751 11207 18757
rect 11149 18748 11161 18751
rect 11112 18720 11161 18748
rect 11112 18708 11118 18720
rect 11149 18717 11161 18720
rect 11195 18717 11207 18751
rect 11149 18711 11207 18717
rect 11238 18708 11244 18760
rect 11296 18708 11302 18760
rect 11517 18751 11575 18757
rect 11517 18717 11529 18751
rect 11563 18717 11575 18751
rect 11517 18711 11575 18717
rect 11422 18680 11428 18692
rect 10652 18652 11428 18680
rect 10652 18640 10658 18652
rect 11422 18640 11428 18652
rect 11480 18640 11486 18692
rect 6917 18615 6975 18621
rect 6917 18612 6929 18615
rect 6288 18584 6929 18612
rect 6917 18581 6929 18584
rect 6963 18612 6975 18615
rect 7098 18612 7104 18624
rect 6963 18584 7104 18612
rect 6963 18581 6975 18584
rect 6917 18575 6975 18581
rect 7098 18572 7104 18584
rect 7156 18572 7162 18624
rect 7834 18572 7840 18624
rect 7892 18572 7898 18624
rect 8294 18572 8300 18624
rect 8352 18612 8358 18624
rect 8662 18612 8668 18624
rect 8352 18584 8668 18612
rect 8352 18572 8358 18584
rect 8662 18572 8668 18584
rect 8720 18612 8726 18624
rect 9217 18615 9275 18621
rect 9217 18612 9229 18615
rect 8720 18584 9229 18612
rect 8720 18572 8726 18584
rect 9217 18581 9229 18584
rect 9263 18581 9275 18615
rect 9217 18575 9275 18581
rect 9766 18572 9772 18624
rect 9824 18612 9830 18624
rect 10686 18612 10692 18624
rect 9824 18584 10692 18612
rect 9824 18572 9830 18584
rect 10686 18572 10692 18584
rect 10744 18612 10750 18624
rect 10870 18612 10876 18624
rect 10744 18584 10876 18612
rect 10744 18572 10750 18584
rect 10870 18572 10876 18584
rect 10928 18612 10934 18624
rect 11532 18612 11560 18711
rect 11606 18708 11612 18760
rect 11664 18748 11670 18760
rect 11992 18757 12020 18924
rect 12618 18912 12624 18924
rect 12676 18912 12682 18964
rect 14090 18912 14096 18964
rect 14148 18952 14154 18964
rect 14277 18955 14335 18961
rect 14277 18952 14289 18955
rect 14148 18924 14289 18952
rect 14148 18912 14154 18924
rect 14277 18921 14289 18924
rect 14323 18921 14335 18955
rect 14277 18915 14335 18921
rect 14921 18955 14979 18961
rect 14921 18921 14933 18955
rect 14967 18952 14979 18955
rect 15010 18952 15016 18964
rect 14967 18924 15016 18952
rect 14967 18921 14979 18924
rect 14921 18915 14979 18921
rect 15010 18912 15016 18924
rect 15068 18912 15074 18964
rect 15378 18952 15384 18964
rect 15120 18924 15384 18952
rect 13633 18887 13691 18893
rect 13633 18853 13645 18887
rect 13679 18884 13691 18887
rect 13906 18884 13912 18896
rect 13679 18856 13912 18884
rect 13679 18853 13691 18856
rect 13633 18847 13691 18853
rect 13906 18844 13912 18856
rect 13964 18844 13970 18896
rect 15120 18816 15148 18924
rect 15378 18912 15384 18924
rect 15436 18912 15442 18964
rect 15194 18844 15200 18896
rect 15252 18884 15258 18896
rect 15252 18856 15884 18884
rect 15252 18844 15258 18856
rect 15470 18816 15476 18828
rect 14476 18788 15148 18816
rect 15304 18788 15476 18816
rect 11793 18751 11851 18757
rect 11793 18748 11805 18751
rect 11664 18720 11805 18748
rect 11664 18708 11670 18720
rect 11793 18717 11805 18720
rect 11839 18717 11851 18751
rect 11793 18711 11851 18717
rect 11977 18751 12035 18757
rect 11977 18717 11989 18751
rect 12023 18717 12035 18751
rect 11977 18711 12035 18717
rect 12250 18708 12256 18760
rect 12308 18708 12314 18760
rect 12526 18757 12532 18760
rect 12520 18748 12532 18757
rect 12487 18720 12532 18748
rect 12520 18711 12532 18720
rect 12526 18708 12532 18711
rect 12584 18708 12590 18760
rect 13906 18708 13912 18760
rect 13964 18708 13970 18760
rect 14476 18757 14504 18788
rect 14461 18751 14519 18757
rect 14461 18717 14473 18751
rect 14507 18717 14519 18751
rect 14461 18711 14519 18717
rect 14553 18751 14611 18757
rect 14553 18717 14565 18751
rect 14599 18748 14611 18751
rect 14642 18748 14648 18760
rect 14599 18720 14648 18748
rect 14599 18717 14611 18720
rect 14553 18711 14611 18717
rect 14642 18708 14648 18720
rect 14700 18708 14706 18760
rect 14734 18708 14740 18760
rect 14792 18708 14798 18760
rect 14829 18751 14887 18757
rect 14829 18717 14841 18751
rect 14875 18717 14887 18751
rect 14829 18711 14887 18717
rect 14844 18680 14872 18711
rect 15102 18708 15108 18760
rect 15160 18748 15166 18760
rect 15304 18757 15332 18788
rect 15470 18776 15476 18788
rect 15528 18776 15534 18828
rect 15197 18751 15255 18757
rect 15197 18748 15209 18751
rect 15160 18720 15209 18748
rect 15160 18708 15166 18720
rect 15197 18717 15209 18720
rect 15243 18717 15255 18751
rect 15197 18711 15255 18717
rect 15289 18751 15347 18757
rect 15289 18717 15301 18751
rect 15335 18717 15347 18751
rect 15289 18711 15347 18717
rect 15378 18708 15384 18760
rect 15436 18708 15442 18760
rect 15562 18708 15568 18760
rect 15620 18708 15626 18760
rect 15856 18757 15884 18856
rect 15841 18751 15899 18757
rect 15841 18717 15853 18751
rect 15887 18748 15899 18751
rect 16114 18748 16120 18760
rect 15887 18720 16120 18748
rect 15887 18717 15899 18720
rect 15841 18711 15899 18717
rect 16114 18708 16120 18720
rect 16172 18708 16178 18760
rect 16209 18751 16267 18757
rect 16209 18717 16221 18751
rect 16255 18748 16267 18751
rect 16298 18748 16304 18760
rect 16255 18720 16304 18748
rect 16255 18717 16267 18720
rect 16209 18711 16267 18717
rect 16298 18708 16304 18720
rect 16356 18708 16362 18760
rect 14844 18652 15700 18680
rect 10928 18584 11560 18612
rect 10928 18572 10934 18584
rect 11698 18572 11704 18624
rect 11756 18572 11762 18624
rect 13262 18572 13268 18624
rect 13320 18612 13326 18624
rect 15672 18621 15700 18652
rect 15746 18640 15752 18692
rect 15804 18680 15810 18692
rect 15930 18680 15936 18692
rect 15804 18652 15936 18680
rect 15804 18640 15810 18652
rect 15930 18640 15936 18652
rect 15988 18640 15994 18692
rect 16022 18640 16028 18692
rect 16080 18640 16086 18692
rect 13725 18615 13783 18621
rect 13725 18612 13737 18615
rect 13320 18584 13737 18612
rect 13320 18572 13326 18584
rect 13725 18581 13737 18584
rect 13771 18581 13783 18615
rect 13725 18575 13783 18581
rect 15657 18615 15715 18621
rect 15657 18581 15669 18615
rect 15703 18581 15715 18615
rect 15657 18575 15715 18581
rect 1104 18522 16652 18544
rect 1104 18470 4874 18522
rect 4926 18470 4938 18522
rect 4990 18470 5002 18522
rect 5054 18470 5066 18522
rect 5118 18470 5130 18522
rect 5182 18470 16652 18522
rect 1104 18448 16652 18470
rect 3970 18368 3976 18420
rect 4028 18408 4034 18420
rect 6549 18411 6607 18417
rect 4028 18380 5212 18408
rect 4028 18368 4034 18380
rect 3234 18300 3240 18352
rect 3292 18340 3298 18352
rect 3786 18340 3792 18352
rect 3292 18312 3792 18340
rect 3292 18300 3298 18312
rect 3786 18300 3792 18312
rect 3844 18340 3850 18352
rect 3881 18343 3939 18349
rect 3881 18340 3893 18343
rect 3844 18312 3893 18340
rect 3844 18300 3850 18312
rect 3881 18309 3893 18312
rect 3927 18309 3939 18343
rect 3881 18303 3939 18309
rect 4154 18300 4160 18352
rect 4212 18340 4218 18352
rect 4212 18312 4844 18340
rect 4212 18300 4218 18312
rect 2317 18275 2375 18281
rect 2317 18241 2329 18275
rect 2363 18272 2375 18275
rect 2406 18272 2412 18284
rect 2363 18244 2412 18272
rect 2363 18241 2375 18244
rect 2317 18235 2375 18241
rect 2406 18232 2412 18244
rect 2464 18232 2470 18284
rect 2501 18275 2559 18281
rect 2501 18241 2513 18275
rect 2547 18272 2559 18275
rect 3050 18272 3056 18284
rect 2547 18244 3056 18272
rect 2547 18241 2559 18244
rect 2501 18235 2559 18241
rect 3050 18232 3056 18244
rect 3108 18232 3114 18284
rect 4816 18281 4844 18312
rect 5184 18284 5212 18380
rect 6549 18377 6561 18411
rect 6595 18408 6607 18411
rect 7926 18408 7932 18420
rect 6595 18380 7932 18408
rect 6595 18377 6607 18380
rect 6549 18371 6607 18377
rect 7926 18368 7932 18380
rect 7984 18368 7990 18420
rect 8478 18368 8484 18420
rect 8536 18408 8542 18420
rect 9122 18408 9128 18420
rect 8536 18380 9128 18408
rect 8536 18368 8542 18380
rect 9122 18368 9128 18380
rect 9180 18408 9186 18420
rect 9180 18380 9812 18408
rect 9180 18368 9186 18380
rect 7006 18340 7012 18352
rect 6840 18312 7012 18340
rect 4801 18275 4859 18281
rect 4801 18241 4813 18275
rect 4847 18272 4859 18275
rect 4982 18272 4988 18284
rect 4847 18244 4988 18272
rect 4847 18241 4859 18244
rect 4801 18235 4859 18241
rect 4982 18232 4988 18244
rect 5040 18232 5046 18284
rect 5166 18232 5172 18284
rect 5224 18272 5230 18284
rect 5537 18275 5595 18281
rect 5537 18272 5549 18275
rect 5224 18244 5549 18272
rect 5224 18232 5230 18244
rect 5537 18241 5549 18244
rect 5583 18241 5595 18275
rect 5537 18235 5595 18241
rect 5994 18232 6000 18284
rect 6052 18272 6058 18284
rect 6365 18275 6423 18281
rect 6365 18272 6377 18275
rect 6052 18244 6377 18272
rect 6052 18232 6058 18244
rect 6365 18241 6377 18244
rect 6411 18241 6423 18275
rect 6365 18235 6423 18241
rect 6549 18275 6607 18281
rect 6549 18241 6561 18275
rect 6595 18272 6607 18275
rect 6638 18272 6644 18284
rect 6595 18244 6644 18272
rect 6595 18241 6607 18244
rect 6549 18235 6607 18241
rect 6380 18204 6408 18235
rect 6638 18232 6644 18244
rect 6696 18232 6702 18284
rect 6840 18281 6868 18312
rect 7006 18300 7012 18312
rect 7064 18300 7070 18352
rect 7374 18349 7380 18352
rect 7368 18303 7380 18349
rect 7374 18300 7380 18303
rect 7432 18300 7438 18352
rect 8386 18300 8392 18352
rect 8444 18340 8450 18352
rect 8573 18343 8631 18349
rect 8573 18340 8585 18343
rect 8444 18312 8585 18340
rect 8444 18300 8450 18312
rect 8573 18309 8585 18312
rect 8619 18340 8631 18343
rect 9582 18340 9588 18352
rect 8619 18312 9588 18340
rect 8619 18309 8631 18312
rect 8573 18303 8631 18309
rect 9582 18300 9588 18312
rect 9640 18300 9646 18352
rect 9784 18349 9812 18380
rect 10134 18368 10140 18420
rect 10192 18368 10198 18420
rect 10502 18368 10508 18420
rect 10560 18408 10566 18420
rect 10965 18411 11023 18417
rect 10965 18408 10977 18411
rect 10560 18380 10977 18408
rect 10560 18368 10566 18380
rect 10965 18377 10977 18380
rect 11011 18377 11023 18411
rect 10965 18371 11023 18377
rect 11333 18411 11391 18417
rect 11333 18377 11345 18411
rect 11379 18408 11391 18411
rect 13906 18408 13912 18420
rect 11379 18380 13912 18408
rect 11379 18377 11391 18380
rect 11333 18371 11391 18377
rect 13906 18368 13912 18380
rect 13964 18368 13970 18420
rect 14182 18368 14188 18420
rect 14240 18368 14246 18420
rect 15378 18368 15384 18420
rect 15436 18408 15442 18420
rect 16301 18411 16359 18417
rect 16301 18408 16313 18411
rect 15436 18380 16313 18408
rect 15436 18368 15442 18380
rect 16301 18377 16313 18380
rect 16347 18377 16359 18411
rect 16301 18371 16359 18377
rect 9769 18343 9827 18349
rect 9769 18309 9781 18343
rect 9815 18309 9827 18343
rect 9769 18303 9827 18309
rect 9985 18343 10043 18349
rect 9985 18309 9997 18343
rect 10031 18340 10043 18343
rect 10318 18340 10324 18352
rect 10031 18312 10324 18340
rect 10031 18309 10043 18312
rect 9985 18303 10043 18309
rect 10318 18300 10324 18312
rect 10376 18340 10382 18352
rect 12250 18340 12256 18352
rect 10376 18312 10916 18340
rect 10376 18300 10382 18312
rect 6825 18275 6883 18281
rect 6825 18241 6837 18275
rect 6871 18241 6883 18275
rect 6825 18235 6883 18241
rect 6914 18232 6920 18284
rect 6972 18272 6978 18284
rect 7101 18275 7159 18281
rect 7101 18272 7113 18275
rect 6972 18244 7113 18272
rect 6972 18232 6978 18244
rect 7101 18241 7113 18244
rect 7147 18241 7159 18275
rect 7742 18272 7748 18284
rect 7101 18235 7159 18241
rect 7208 18270 7420 18272
rect 7484 18270 7748 18272
rect 7208 18244 7748 18270
rect 7208 18204 7236 18244
rect 7392 18242 7512 18244
rect 7742 18232 7748 18244
rect 7800 18272 7806 18284
rect 9401 18275 9459 18281
rect 7800 18244 8892 18272
rect 7800 18232 7806 18244
rect 6380 18176 7236 18204
rect 8754 18136 8760 18148
rect 8404 18108 8760 18136
rect 2130 18028 2136 18080
rect 2188 18068 2194 18080
rect 2317 18071 2375 18077
rect 2317 18068 2329 18071
rect 2188 18040 2329 18068
rect 2188 18028 2194 18040
rect 2317 18037 2329 18040
rect 2363 18037 2375 18071
rect 2317 18031 2375 18037
rect 6733 18071 6791 18077
rect 6733 18037 6745 18071
rect 6779 18068 6791 18071
rect 8404 18068 8432 18108
rect 8754 18096 8760 18108
rect 8812 18096 8818 18148
rect 8864 18145 8892 18244
rect 9401 18241 9413 18275
rect 9447 18241 9459 18275
rect 9401 18235 9459 18241
rect 9493 18275 9551 18281
rect 9493 18241 9505 18275
rect 9539 18272 9551 18275
rect 9674 18272 9680 18284
rect 9539 18244 9680 18272
rect 9539 18241 9551 18244
rect 9493 18235 9551 18241
rect 9416 18204 9444 18235
rect 9674 18232 9680 18244
rect 9732 18232 9738 18284
rect 9858 18232 9864 18284
rect 9916 18232 9922 18284
rect 10229 18275 10287 18281
rect 10229 18272 10241 18275
rect 9968 18244 10241 18272
rect 9876 18204 9904 18232
rect 9416 18176 9904 18204
rect 8849 18139 8907 18145
rect 8849 18105 8861 18139
rect 8895 18105 8907 18139
rect 8849 18099 8907 18105
rect 9033 18139 9091 18145
rect 9033 18105 9045 18139
rect 9079 18136 9091 18139
rect 9858 18136 9864 18148
rect 9079 18108 9864 18136
rect 9079 18105 9091 18108
rect 9033 18099 9091 18105
rect 9858 18096 9864 18108
rect 9916 18096 9922 18148
rect 6779 18040 8432 18068
rect 6779 18037 6791 18040
rect 6733 18031 6791 18037
rect 9398 18028 9404 18080
rect 9456 18028 9462 18080
rect 9582 18028 9588 18080
rect 9640 18068 9646 18080
rect 9968 18077 9996 18244
rect 10229 18241 10241 18244
rect 10275 18241 10287 18275
rect 10229 18235 10287 18241
rect 10413 18275 10471 18281
rect 10413 18241 10425 18275
rect 10459 18241 10471 18275
rect 10413 18235 10471 18241
rect 10428 18204 10456 18235
rect 10594 18232 10600 18284
rect 10652 18232 10658 18284
rect 10888 18281 10916 18312
rect 11900 18312 12256 18340
rect 10873 18275 10931 18281
rect 10873 18241 10885 18275
rect 10919 18241 10931 18275
rect 10873 18235 10931 18241
rect 11149 18275 11207 18281
rect 11149 18241 11161 18275
rect 11195 18272 11207 18275
rect 11514 18272 11520 18284
rect 11195 18244 11520 18272
rect 11195 18241 11207 18244
rect 11149 18235 11207 18241
rect 11514 18232 11520 18244
rect 11572 18232 11578 18284
rect 11900 18281 11928 18312
rect 12250 18300 12256 18312
rect 12308 18340 12314 18352
rect 15746 18340 15752 18352
rect 12308 18312 12434 18340
rect 12308 18300 12314 18312
rect 12158 18281 12164 18284
rect 11885 18275 11943 18281
rect 11885 18241 11897 18275
rect 11931 18241 11943 18275
rect 11885 18235 11943 18241
rect 12152 18235 12164 18281
rect 12158 18232 12164 18235
rect 12216 18232 12222 18284
rect 12406 18272 12434 18312
rect 14384 18312 15752 18340
rect 14274 18272 14280 18284
rect 12406 18244 14280 18272
rect 14274 18232 14280 18244
rect 14332 18232 14338 18284
rect 14384 18281 14412 18312
rect 15746 18300 15752 18312
rect 15804 18340 15810 18352
rect 16117 18343 16175 18349
rect 16117 18340 16129 18343
rect 15804 18312 16129 18340
rect 15804 18300 15810 18312
rect 16117 18309 16129 18312
rect 16163 18309 16175 18343
rect 16117 18303 16175 18309
rect 14369 18275 14427 18281
rect 14369 18241 14381 18275
rect 14415 18241 14427 18275
rect 14369 18235 14427 18241
rect 14550 18232 14556 18284
rect 14608 18272 14614 18284
rect 14717 18275 14775 18281
rect 14717 18272 14729 18275
rect 14608 18244 14729 18272
rect 14608 18232 14614 18244
rect 14717 18241 14729 18244
rect 14763 18241 14775 18275
rect 14717 18235 14775 18241
rect 15654 18232 15660 18284
rect 15712 18272 15718 18284
rect 15838 18272 15844 18284
rect 15712 18244 15844 18272
rect 15712 18232 15718 18244
rect 15838 18232 15844 18244
rect 15896 18272 15902 18284
rect 15933 18275 15991 18281
rect 15933 18272 15945 18275
rect 15896 18244 15945 18272
rect 15896 18232 15902 18244
rect 15933 18241 15945 18244
rect 15979 18241 15991 18275
rect 15933 18235 15991 18241
rect 10686 18204 10692 18216
rect 10428 18176 10692 18204
rect 10686 18164 10692 18176
rect 10744 18164 10750 18216
rect 13909 18207 13967 18213
rect 13909 18173 13921 18207
rect 13955 18173 13967 18207
rect 14292 18204 14320 18232
rect 14461 18207 14519 18213
rect 14461 18204 14473 18207
rect 14292 18176 14473 18204
rect 13909 18167 13967 18173
rect 14461 18173 14473 18176
rect 14507 18173 14519 18207
rect 14461 18167 14519 18173
rect 13265 18139 13323 18145
rect 13265 18105 13277 18139
rect 13311 18136 13323 18139
rect 13924 18136 13952 18167
rect 14090 18136 14096 18148
rect 13311 18108 14096 18136
rect 13311 18105 13323 18108
rect 13265 18099 13323 18105
rect 14090 18096 14096 18108
rect 14148 18096 14154 18148
rect 9953 18071 10011 18077
rect 9953 18068 9965 18071
rect 9640 18040 9965 18068
rect 9640 18028 9646 18040
rect 9953 18037 9965 18040
rect 9999 18037 10011 18071
rect 9953 18031 10011 18037
rect 10594 18028 10600 18080
rect 10652 18068 10658 18080
rect 10962 18068 10968 18080
rect 10652 18040 10968 18068
rect 10652 18028 10658 18040
rect 10962 18028 10968 18040
rect 11020 18028 11026 18080
rect 13354 18028 13360 18080
rect 13412 18028 13418 18080
rect 15378 18028 15384 18080
rect 15436 18068 15442 18080
rect 15841 18071 15899 18077
rect 15841 18068 15853 18071
rect 15436 18040 15853 18068
rect 15436 18028 15442 18040
rect 15841 18037 15853 18040
rect 15887 18037 15899 18071
rect 15841 18031 15899 18037
rect 1104 17978 16652 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 16652 17978
rect 1104 17904 16652 17926
rect 1581 17867 1639 17873
rect 1581 17833 1593 17867
rect 1627 17864 1639 17867
rect 1946 17864 1952 17876
rect 1627 17836 1952 17864
rect 1627 17833 1639 17836
rect 1581 17827 1639 17833
rect 1946 17824 1952 17836
rect 2004 17824 2010 17876
rect 2041 17867 2099 17873
rect 2041 17833 2053 17867
rect 2087 17864 2099 17867
rect 2866 17864 2872 17876
rect 2087 17836 2872 17864
rect 2087 17833 2099 17836
rect 2041 17827 2099 17833
rect 2866 17824 2872 17836
rect 2924 17824 2930 17876
rect 3326 17824 3332 17876
rect 3384 17864 3390 17876
rect 3513 17867 3571 17873
rect 3513 17864 3525 17867
rect 3384 17836 3525 17864
rect 3384 17824 3390 17836
rect 3513 17833 3525 17836
rect 3559 17833 3571 17867
rect 3513 17827 3571 17833
rect 4525 17867 4583 17873
rect 4525 17833 4537 17867
rect 4571 17864 4583 17867
rect 4614 17864 4620 17876
rect 4571 17836 4620 17864
rect 4571 17833 4583 17836
rect 4525 17827 4583 17833
rect 4614 17824 4620 17836
rect 4672 17824 4678 17876
rect 5350 17824 5356 17876
rect 5408 17824 5414 17876
rect 7285 17867 7343 17873
rect 7285 17833 7297 17867
rect 7331 17864 7343 17867
rect 7374 17864 7380 17876
rect 7331 17836 7380 17864
rect 7331 17833 7343 17836
rect 7285 17827 7343 17833
rect 7374 17824 7380 17836
rect 7432 17824 7438 17876
rect 7558 17824 7564 17876
rect 7616 17824 7622 17876
rect 10226 17824 10232 17876
rect 10284 17824 10290 17876
rect 12158 17824 12164 17876
rect 12216 17864 12222 17876
rect 12253 17867 12311 17873
rect 12253 17864 12265 17867
rect 12216 17836 12265 17864
rect 12216 17824 12222 17836
rect 12253 17833 12265 17836
rect 12299 17833 12311 17867
rect 12253 17827 12311 17833
rect 12342 17824 12348 17876
rect 12400 17864 12406 17876
rect 14369 17867 14427 17873
rect 12400 17836 13676 17864
rect 12400 17824 12406 17836
rect 2777 17799 2835 17805
rect 2777 17765 2789 17799
rect 2823 17796 2835 17799
rect 2958 17796 2964 17808
rect 2823 17768 2964 17796
rect 2823 17765 2835 17768
rect 2777 17759 2835 17765
rect 2958 17756 2964 17768
rect 3016 17796 3022 17808
rect 3786 17796 3792 17808
rect 3016 17768 3792 17796
rect 3016 17756 3022 17768
rect 3786 17756 3792 17768
rect 3844 17756 3850 17808
rect 8573 17799 8631 17805
rect 8573 17765 8585 17799
rect 8619 17796 8631 17799
rect 8754 17796 8760 17808
rect 8619 17768 8760 17796
rect 8619 17765 8631 17768
rect 8573 17759 8631 17765
rect 8754 17756 8760 17768
rect 8812 17756 8818 17808
rect 13648 17796 13676 17836
rect 14369 17833 14381 17867
rect 14415 17864 14427 17867
rect 14550 17864 14556 17876
rect 14415 17836 14556 17864
rect 14415 17833 14427 17836
rect 14369 17827 14427 17833
rect 14550 17824 14556 17836
rect 14608 17824 14614 17876
rect 15102 17864 15108 17876
rect 14660 17836 15108 17864
rect 13648 17768 13768 17796
rect 106 17688 112 17740
rect 164 17728 170 17740
rect 164 17700 8984 17728
rect 164 17688 170 17700
rect 2406 17620 2412 17672
rect 2464 17620 2470 17672
rect 2593 17663 2651 17669
rect 2593 17662 2605 17663
rect 2536 17634 2605 17662
rect 1762 17552 1768 17604
rect 1820 17552 1826 17604
rect 2225 17595 2283 17601
rect 2225 17561 2237 17595
rect 2271 17592 2283 17595
rect 2314 17592 2320 17604
rect 2271 17564 2320 17592
rect 2271 17561 2283 17564
rect 2225 17555 2283 17561
rect 2314 17552 2320 17564
rect 2372 17552 2378 17604
rect 2536 17592 2564 17634
rect 2593 17629 2605 17634
rect 2639 17629 2651 17663
rect 2593 17623 2651 17629
rect 2682 17620 2688 17672
rect 2740 17620 2746 17672
rect 3050 17620 3056 17672
rect 3108 17660 3114 17672
rect 3148 17663 3206 17669
rect 3148 17660 3160 17663
rect 3108 17632 3160 17660
rect 3108 17620 3114 17632
rect 3148 17629 3160 17632
rect 3194 17629 3206 17663
rect 3148 17623 3206 17629
rect 3326 17620 3332 17672
rect 3384 17620 3390 17672
rect 3418 17620 3424 17672
rect 3476 17620 3482 17672
rect 3605 17663 3663 17669
rect 3605 17629 3617 17663
rect 3651 17629 3663 17663
rect 3605 17623 3663 17629
rect 3344 17592 3372 17620
rect 2536 17564 3372 17592
rect 3510 17552 3516 17604
rect 3568 17592 3574 17604
rect 3620 17592 3648 17623
rect 3786 17620 3792 17672
rect 3844 17620 3850 17672
rect 3878 17620 3884 17672
rect 3936 17620 3942 17672
rect 4709 17663 4767 17669
rect 4709 17629 4721 17663
rect 4755 17660 4767 17663
rect 4982 17660 4988 17672
rect 4755 17632 4988 17660
rect 4755 17629 4767 17632
rect 4709 17623 4767 17629
rect 4982 17620 4988 17632
rect 5040 17620 5046 17672
rect 5166 17620 5172 17672
rect 5224 17620 5230 17672
rect 5262 17663 5320 17669
rect 5262 17629 5274 17663
rect 5308 17629 5320 17663
rect 5262 17623 5320 17629
rect 7285 17663 7343 17669
rect 7285 17629 7297 17663
rect 7331 17629 7343 17663
rect 7285 17623 7343 17629
rect 7469 17663 7527 17669
rect 7469 17629 7481 17663
rect 7515 17660 7527 17663
rect 7745 17663 7803 17669
rect 7745 17660 7757 17663
rect 7515 17632 7757 17660
rect 7515 17629 7527 17632
rect 7469 17623 7527 17629
rect 7745 17629 7757 17632
rect 7791 17629 7803 17663
rect 7745 17623 7803 17629
rect 4062 17592 4068 17604
rect 3568 17564 4068 17592
rect 3568 17552 3574 17564
rect 4062 17552 4068 17564
rect 4120 17552 4126 17604
rect 4893 17595 4951 17601
rect 4893 17561 4905 17595
rect 4939 17561 4951 17595
rect 5000 17592 5028 17620
rect 5276 17592 5304 17623
rect 5000 17564 5304 17592
rect 4893 17555 4951 17561
rect 1394 17484 1400 17536
rect 1452 17484 1458 17536
rect 1578 17533 1584 17536
rect 1565 17527 1584 17533
rect 1565 17493 1577 17527
rect 1565 17487 1584 17493
rect 1578 17484 1584 17487
rect 1636 17484 1642 17536
rect 1854 17484 1860 17536
rect 1912 17484 1918 17536
rect 2025 17527 2083 17533
rect 2025 17493 2037 17527
rect 2071 17524 2083 17527
rect 2406 17524 2412 17536
rect 2071 17496 2412 17524
rect 2071 17493 2083 17496
rect 2025 17487 2083 17493
rect 2406 17484 2412 17496
rect 2464 17484 2470 17536
rect 2498 17484 2504 17536
rect 2556 17484 2562 17536
rect 3142 17484 3148 17536
rect 3200 17484 3206 17536
rect 3329 17527 3387 17533
rect 3329 17493 3341 17527
rect 3375 17524 3387 17527
rect 3418 17524 3424 17536
rect 3375 17496 3424 17524
rect 3375 17493 3387 17496
rect 3329 17487 3387 17493
rect 3418 17484 3424 17496
rect 3476 17484 3482 17536
rect 4908 17524 4936 17555
rect 5166 17524 5172 17536
rect 4908 17496 5172 17524
rect 5166 17484 5172 17496
rect 5224 17524 5230 17536
rect 6086 17524 6092 17536
rect 5224 17496 6092 17524
rect 5224 17484 5230 17496
rect 6086 17484 6092 17496
rect 6144 17484 6150 17536
rect 7300 17524 7328 17623
rect 7760 17592 7788 17623
rect 7834 17620 7840 17672
rect 7892 17620 7898 17672
rect 7926 17620 7932 17672
rect 7984 17620 7990 17672
rect 8113 17663 8171 17669
rect 8113 17629 8125 17663
rect 8159 17660 8171 17663
rect 8294 17660 8300 17672
rect 8159 17632 8300 17660
rect 8159 17629 8171 17632
rect 8113 17623 8171 17629
rect 8294 17620 8300 17632
rect 8352 17620 8358 17672
rect 8386 17620 8392 17672
rect 8444 17620 8450 17672
rect 8662 17620 8668 17672
rect 8720 17620 8726 17672
rect 8956 17669 8984 17700
rect 11698 17688 11704 17740
rect 11756 17728 11762 17740
rect 12805 17731 12863 17737
rect 12805 17728 12817 17731
rect 11756 17700 12817 17728
rect 11756 17688 11762 17700
rect 12805 17697 12817 17700
rect 12851 17697 12863 17731
rect 12805 17691 12863 17697
rect 8941 17663 8999 17669
rect 8941 17629 8953 17663
rect 8987 17629 8999 17663
rect 8941 17623 8999 17629
rect 12621 17663 12679 17669
rect 12621 17629 12633 17663
rect 12667 17660 12679 17663
rect 13354 17660 13360 17672
rect 12667 17632 13360 17660
rect 12667 17629 12679 17632
rect 12621 17623 12679 17629
rect 13354 17620 13360 17632
rect 13412 17620 13418 17672
rect 13541 17663 13599 17669
rect 13541 17629 13553 17663
rect 13587 17629 13599 17663
rect 13541 17623 13599 17629
rect 8846 17592 8852 17604
rect 7760 17564 8852 17592
rect 8846 17552 8852 17564
rect 8904 17552 8910 17604
rect 12894 17552 12900 17604
rect 12952 17592 12958 17604
rect 13556 17592 13584 17623
rect 13630 17620 13636 17672
rect 13688 17620 13694 17672
rect 13740 17669 13768 17768
rect 13725 17663 13783 17669
rect 13725 17629 13737 17663
rect 13771 17629 13783 17663
rect 13725 17623 13783 17629
rect 13906 17620 13912 17672
rect 13964 17620 13970 17672
rect 14090 17620 14096 17672
rect 14148 17620 14154 17672
rect 14274 17620 14280 17672
rect 14332 17660 14338 17672
rect 14660 17669 14688 17836
rect 15102 17824 15108 17836
rect 15160 17824 15166 17876
rect 14826 17796 14832 17808
rect 14752 17768 14832 17796
rect 14752 17669 14780 17768
rect 14826 17756 14832 17768
rect 14884 17756 14890 17808
rect 15105 17731 15163 17737
rect 15105 17728 15117 17731
rect 14844 17700 15117 17728
rect 14844 17669 14872 17700
rect 15105 17697 15117 17700
rect 15151 17697 15163 17731
rect 15562 17728 15568 17740
rect 15105 17691 15163 17697
rect 15488 17700 15568 17728
rect 14645 17663 14703 17669
rect 14645 17660 14657 17663
rect 14332 17632 14657 17660
rect 14332 17620 14338 17632
rect 14645 17629 14657 17632
rect 14691 17629 14703 17663
rect 14645 17623 14703 17629
rect 14737 17663 14795 17669
rect 14737 17629 14749 17663
rect 14783 17629 14795 17663
rect 14737 17623 14795 17629
rect 14829 17663 14887 17669
rect 14829 17629 14841 17663
rect 14875 17629 14887 17663
rect 14829 17623 14887 17629
rect 14918 17620 14924 17672
rect 14976 17660 14982 17672
rect 15488 17669 15516 17700
rect 15562 17688 15568 17700
rect 15620 17728 15626 17740
rect 16206 17728 16212 17740
rect 15620 17700 16212 17728
rect 15620 17688 15626 17700
rect 16206 17688 16212 17700
rect 16264 17688 16270 17740
rect 15013 17663 15071 17669
rect 15013 17660 15025 17663
rect 14976 17632 15025 17660
rect 14976 17620 14982 17632
rect 15013 17629 15025 17632
rect 15059 17629 15071 17663
rect 15013 17623 15071 17629
rect 15473 17663 15531 17669
rect 15473 17629 15485 17663
rect 15519 17629 15531 17663
rect 15473 17623 15531 17629
rect 16298 17620 16304 17672
rect 16356 17620 16362 17672
rect 12952 17564 13584 17592
rect 12952 17552 12958 17564
rect 15286 17552 15292 17604
rect 15344 17552 15350 17604
rect 15565 17595 15623 17601
rect 15565 17561 15577 17595
rect 15611 17592 15623 17595
rect 15654 17592 15660 17604
rect 15611 17564 15660 17592
rect 15611 17561 15623 17564
rect 15565 17555 15623 17561
rect 15654 17552 15660 17564
rect 15712 17552 15718 17604
rect 15749 17595 15807 17601
rect 15749 17561 15761 17595
rect 15795 17592 15807 17595
rect 15838 17592 15844 17604
rect 15795 17564 15844 17592
rect 15795 17561 15807 17564
rect 15749 17555 15807 17561
rect 15838 17552 15844 17564
rect 15896 17552 15902 17604
rect 8205 17527 8263 17533
rect 8205 17524 8217 17527
rect 7300 17496 8217 17524
rect 8205 17493 8217 17496
rect 8251 17493 8263 17527
rect 8205 17487 8263 17493
rect 12713 17527 12771 17533
rect 12713 17493 12725 17527
rect 12759 17524 12771 17527
rect 13357 17527 13415 17533
rect 13357 17524 13369 17527
rect 12759 17496 13369 17524
rect 12759 17493 12771 17496
rect 12713 17487 12771 17493
rect 13357 17493 13369 17496
rect 13403 17493 13415 17527
rect 13357 17487 13415 17493
rect 14277 17527 14335 17533
rect 14277 17493 14289 17527
rect 14323 17524 14335 17527
rect 15010 17524 15016 17536
rect 14323 17496 15016 17524
rect 14323 17493 14335 17496
rect 14277 17487 14335 17493
rect 15010 17484 15016 17496
rect 15068 17484 15074 17536
rect 15933 17527 15991 17533
rect 15933 17493 15945 17527
rect 15979 17524 15991 17527
rect 16022 17524 16028 17536
rect 15979 17496 16028 17524
rect 15979 17493 15991 17496
rect 15933 17487 15991 17493
rect 16022 17484 16028 17496
rect 16080 17484 16086 17536
rect 16117 17527 16175 17533
rect 16117 17493 16129 17527
rect 16163 17524 16175 17527
rect 16298 17524 16304 17536
rect 16163 17496 16304 17524
rect 16163 17493 16175 17496
rect 16117 17487 16175 17493
rect 16298 17484 16304 17496
rect 16356 17484 16362 17536
rect 1104 17434 16652 17456
rect 1104 17382 4874 17434
rect 4926 17382 4938 17434
rect 4990 17382 5002 17434
rect 5054 17382 5066 17434
rect 5118 17382 5130 17434
rect 5182 17382 16652 17434
rect 1104 17360 16652 17382
rect 2958 17280 2964 17332
rect 3016 17280 3022 17332
rect 8386 17280 8392 17332
rect 8444 17320 8450 17332
rect 8938 17320 8944 17332
rect 8444 17292 8944 17320
rect 8444 17280 8450 17292
rect 5074 17252 5080 17264
rect 1596 17224 2774 17252
rect 1394 17144 1400 17196
rect 1452 17184 1458 17196
rect 1596 17193 1624 17224
rect 1854 17193 1860 17196
rect 1581 17187 1639 17193
rect 1581 17184 1593 17187
rect 1452 17156 1593 17184
rect 1452 17144 1458 17156
rect 1581 17153 1593 17156
rect 1627 17153 1639 17187
rect 1848 17184 1860 17193
rect 1815 17156 1860 17184
rect 1581 17147 1639 17153
rect 1848 17147 1860 17156
rect 1854 17144 1860 17147
rect 1912 17144 1918 17196
rect 2746 17116 2774 17224
rect 3252 17224 5080 17252
rect 3142 17144 3148 17196
rect 3200 17144 3206 17196
rect 3252 17116 3280 17224
rect 3436 17193 3464 17224
rect 5074 17212 5080 17224
rect 5132 17212 5138 17264
rect 5169 17255 5227 17261
rect 5169 17221 5181 17255
rect 5215 17221 5227 17255
rect 5169 17215 5227 17221
rect 3329 17187 3387 17193
rect 3329 17153 3341 17187
rect 3375 17153 3387 17187
rect 3329 17147 3387 17153
rect 3421 17187 3479 17193
rect 3421 17153 3433 17187
rect 3467 17153 3479 17187
rect 3421 17147 3479 17153
rect 2746 17088 3280 17116
rect 3344 17116 3372 17147
rect 3510 17144 3516 17196
rect 3568 17144 3574 17196
rect 3694 17193 3700 17196
rect 3688 17147 3700 17193
rect 3694 17144 3700 17147
rect 3752 17144 3758 17196
rect 3528 17116 3556 17144
rect 3344 17088 3556 17116
rect 5184 17116 5212 17215
rect 5350 17212 5356 17264
rect 5408 17261 5414 17264
rect 5408 17255 5427 17261
rect 5415 17221 5427 17255
rect 5408 17215 5427 17221
rect 5721 17255 5779 17261
rect 5721 17221 5733 17255
rect 5767 17252 5779 17255
rect 6270 17252 6276 17264
rect 5767 17224 6276 17252
rect 5767 17221 5779 17224
rect 5721 17215 5779 17221
rect 5408 17212 5414 17215
rect 6270 17212 6276 17224
rect 6328 17212 6334 17264
rect 5626 17144 5632 17196
rect 5684 17144 5690 17196
rect 5902 17144 5908 17196
rect 5960 17144 5966 17196
rect 8496 17193 8524 17292
rect 8938 17280 8944 17292
rect 8996 17320 9002 17332
rect 9033 17323 9091 17329
rect 9033 17320 9045 17323
rect 8996 17292 9045 17320
rect 8996 17280 9002 17292
rect 9033 17289 9045 17292
rect 9079 17289 9091 17323
rect 9033 17283 9091 17289
rect 9217 17323 9275 17329
rect 9217 17289 9229 17323
rect 9263 17320 9275 17323
rect 9306 17320 9312 17332
rect 9263 17292 9312 17320
rect 9263 17289 9275 17292
rect 9217 17283 9275 17289
rect 9306 17280 9312 17292
rect 9364 17280 9370 17332
rect 10689 17323 10747 17329
rect 10689 17289 10701 17323
rect 10735 17320 10747 17323
rect 10778 17320 10784 17332
rect 10735 17292 10784 17320
rect 10735 17289 10747 17292
rect 10689 17283 10747 17289
rect 10778 17280 10784 17292
rect 10836 17320 10842 17332
rect 11422 17320 11428 17332
rect 10836 17292 11428 17320
rect 10836 17280 10842 17292
rect 11422 17280 11428 17292
rect 11480 17280 11486 17332
rect 13078 17280 13084 17332
rect 13136 17280 13142 17332
rect 13814 17280 13820 17332
rect 13872 17280 13878 17332
rect 14458 17280 14464 17332
rect 14516 17280 14522 17332
rect 14734 17280 14740 17332
rect 14792 17320 14798 17332
rect 15473 17323 15531 17329
rect 15473 17320 15485 17323
rect 14792 17292 15485 17320
rect 14792 17280 14798 17292
rect 15473 17289 15485 17292
rect 15519 17289 15531 17323
rect 15473 17283 15531 17289
rect 8754 17212 8760 17264
rect 8812 17252 8818 17264
rect 8812 17224 9720 17252
rect 8812 17212 8818 17224
rect 8481 17187 8539 17193
rect 8481 17153 8493 17187
rect 8527 17153 8539 17187
rect 8481 17147 8539 17153
rect 9122 17144 9128 17196
rect 9180 17144 9186 17196
rect 9398 17144 9404 17196
rect 9456 17193 9462 17196
rect 9456 17187 9489 17193
rect 9477 17153 9489 17187
rect 9456 17147 9489 17153
rect 9585 17187 9643 17193
rect 9585 17153 9597 17187
rect 9631 17153 9643 17187
rect 9692 17184 9720 17224
rect 9858 17212 9864 17264
rect 9916 17252 9922 17264
rect 9953 17255 10011 17261
rect 9953 17252 9965 17255
rect 9916 17224 9965 17252
rect 9916 17212 9922 17224
rect 9953 17221 9965 17224
rect 9999 17252 10011 17255
rect 10318 17252 10324 17264
rect 9999 17224 10324 17252
rect 9999 17221 10011 17224
rect 9953 17215 10011 17221
rect 10318 17212 10324 17224
rect 10376 17252 10382 17264
rect 15286 17252 15292 17264
rect 10376 17224 10916 17252
rect 10376 17212 10382 17224
rect 10888 17193 10916 17224
rect 14016 17224 15292 17252
rect 10137 17187 10195 17193
rect 10137 17184 10149 17187
rect 9692 17156 10149 17184
rect 9585 17147 9643 17153
rect 10137 17153 10149 17156
rect 10183 17184 10195 17187
rect 10413 17187 10471 17193
rect 10413 17184 10425 17187
rect 10183 17156 10425 17184
rect 10183 17153 10195 17156
rect 10137 17147 10195 17153
rect 10413 17153 10425 17156
rect 10459 17153 10471 17187
rect 10413 17147 10471 17153
rect 10597 17187 10655 17193
rect 10597 17153 10609 17187
rect 10643 17153 10655 17187
rect 10597 17147 10655 17153
rect 10873 17187 10931 17193
rect 10873 17153 10885 17187
rect 10919 17153 10931 17187
rect 10873 17147 10931 17153
rect 11149 17187 11207 17193
rect 11149 17153 11161 17187
rect 11195 17184 11207 17187
rect 12250 17184 12256 17196
rect 11195 17156 12256 17184
rect 11195 17153 11207 17156
rect 11149 17147 11207 17153
rect 9456 17144 9462 17147
rect 5718 17116 5724 17128
rect 5184 17088 5724 17116
rect 5718 17076 5724 17088
rect 5776 17076 5782 17128
rect 8573 17119 8631 17125
rect 8573 17085 8585 17119
rect 8619 17116 8631 17119
rect 8662 17116 8668 17128
rect 8619 17088 8668 17116
rect 8619 17085 8631 17088
rect 8573 17079 8631 17085
rect 8662 17076 8668 17088
rect 8720 17076 8726 17128
rect 9600 17116 9628 17147
rect 9674 17116 9680 17128
rect 8864 17088 9680 17116
rect 8864 17057 8892 17088
rect 9674 17076 9680 17088
rect 9732 17116 9738 17128
rect 10612 17116 10640 17147
rect 9732 17088 10640 17116
rect 9732 17076 9738 17088
rect 10686 17076 10692 17128
rect 10744 17116 10750 17128
rect 11164 17116 11192 17147
rect 12250 17144 12256 17156
rect 12308 17184 12314 17196
rect 12894 17184 12900 17196
rect 12308 17156 12900 17184
rect 12308 17144 12314 17156
rect 12894 17144 12900 17156
rect 12952 17144 12958 17196
rect 13262 17144 13268 17196
rect 13320 17144 13326 17196
rect 13633 17187 13691 17193
rect 13633 17153 13645 17187
rect 13679 17184 13691 17187
rect 13906 17184 13912 17196
rect 13679 17156 13912 17184
rect 13679 17153 13691 17156
rect 13633 17147 13691 17153
rect 13906 17144 13912 17156
rect 13964 17144 13970 17196
rect 14016 17193 14044 17224
rect 15286 17212 15292 17224
rect 15344 17252 15350 17264
rect 15344 17224 16068 17252
rect 15344 17212 15350 17224
rect 14001 17187 14059 17193
rect 14001 17153 14013 17187
rect 14047 17153 14059 17187
rect 14001 17147 14059 17153
rect 14090 17144 14096 17196
rect 14148 17144 14154 17196
rect 14277 17187 14335 17193
rect 14277 17153 14289 17187
rect 14323 17184 14335 17187
rect 14550 17184 14556 17196
rect 14323 17156 14556 17184
rect 14323 17153 14335 17156
rect 14277 17147 14335 17153
rect 14550 17144 14556 17156
rect 14608 17144 14614 17196
rect 14645 17187 14703 17193
rect 14645 17153 14657 17187
rect 14691 17153 14703 17187
rect 14645 17147 14703 17153
rect 10744 17088 11192 17116
rect 11241 17119 11299 17125
rect 10744 17076 10750 17088
rect 11241 17085 11253 17119
rect 11287 17116 11299 17119
rect 11606 17116 11612 17128
rect 11287 17088 11612 17116
rect 11287 17085 11299 17088
rect 11241 17079 11299 17085
rect 11606 17076 11612 17088
rect 11664 17116 11670 17128
rect 12342 17116 12348 17128
rect 11664 17088 12348 17116
rect 11664 17076 11670 17088
rect 12342 17076 12348 17088
rect 12400 17076 12406 17128
rect 14660 17116 14688 17147
rect 14826 17144 14832 17196
rect 14884 17144 14890 17196
rect 15010 17144 15016 17196
rect 15068 17144 15074 17196
rect 15378 17144 15384 17196
rect 15436 17184 15442 17196
rect 15657 17187 15715 17193
rect 15657 17184 15669 17187
rect 15436 17156 15669 17184
rect 15436 17144 15442 17156
rect 15657 17153 15669 17156
rect 15703 17153 15715 17187
rect 15657 17147 15715 17153
rect 15746 17144 15752 17196
rect 15804 17144 15810 17196
rect 16040 17193 16068 17224
rect 15841 17187 15899 17193
rect 15841 17153 15853 17187
rect 15887 17153 15899 17187
rect 15841 17147 15899 17153
rect 16025 17187 16083 17193
rect 16025 17153 16037 17187
rect 16071 17153 16083 17187
rect 16025 17147 16083 17153
rect 14734 17116 14740 17128
rect 14660 17088 14740 17116
rect 14734 17076 14740 17088
rect 14792 17076 14798 17128
rect 15562 17076 15568 17128
rect 15620 17116 15626 17128
rect 15856 17116 15884 17147
rect 16390 17116 16396 17128
rect 15620 17088 16396 17116
rect 15620 17076 15626 17088
rect 16390 17076 16396 17088
rect 16448 17076 16454 17128
rect 8849 17051 8907 17057
rect 8849 17017 8861 17051
rect 8895 17017 8907 17051
rect 8849 17011 8907 17017
rect 10321 17051 10379 17057
rect 10321 17017 10333 17051
rect 10367 17048 10379 17051
rect 11146 17048 11152 17060
rect 10367 17020 11152 17048
rect 10367 17017 10379 17020
rect 10321 17011 10379 17017
rect 11146 17008 11152 17020
rect 11204 17048 11210 17060
rect 11790 17048 11796 17060
rect 11204 17020 11796 17048
rect 11204 17008 11210 17020
rect 11790 17008 11796 17020
rect 11848 17008 11854 17060
rect 13449 17051 13507 17057
rect 13449 17017 13461 17051
rect 13495 17048 13507 17051
rect 15010 17048 15016 17060
rect 13495 17020 15016 17048
rect 13495 17017 13507 17020
rect 13449 17011 13507 17017
rect 15010 17008 15016 17020
rect 15068 17008 15074 17060
rect 15194 17008 15200 17060
rect 15252 17008 15258 17060
rect 3329 16983 3387 16989
rect 3329 16949 3341 16983
rect 3375 16980 3387 16983
rect 3786 16980 3792 16992
rect 3375 16952 3792 16980
rect 3375 16949 3387 16952
rect 3329 16943 3387 16949
rect 3786 16940 3792 16952
rect 3844 16940 3850 16992
rect 4062 16940 4068 16992
rect 4120 16980 4126 16992
rect 4801 16983 4859 16989
rect 4801 16980 4813 16983
rect 4120 16952 4813 16980
rect 4120 16940 4126 16952
rect 4801 16949 4813 16952
rect 4847 16949 4859 16983
rect 4801 16943 4859 16949
rect 5258 16940 5264 16992
rect 5316 16980 5322 16992
rect 5353 16983 5411 16989
rect 5353 16980 5365 16983
rect 5316 16952 5365 16980
rect 5316 16940 5322 16952
rect 5353 16949 5365 16952
rect 5399 16949 5411 16983
rect 5353 16943 5411 16949
rect 5534 16940 5540 16992
rect 5592 16940 5598 16992
rect 5810 16940 5816 16992
rect 5868 16980 5874 16992
rect 6089 16983 6147 16989
rect 6089 16980 6101 16983
rect 5868 16952 6101 16980
rect 5868 16940 5874 16952
rect 6089 16949 6101 16952
rect 6135 16949 6147 16983
rect 6089 16943 6147 16949
rect 7098 16940 7104 16992
rect 7156 16980 7162 16992
rect 8481 16983 8539 16989
rect 8481 16980 8493 16983
rect 7156 16952 8493 16980
rect 7156 16940 7162 16952
rect 8481 16949 8493 16952
rect 8527 16949 8539 16983
rect 8481 16943 8539 16949
rect 12618 16940 12624 16992
rect 12676 16980 12682 16992
rect 14274 16980 14280 16992
rect 12676 16952 14280 16980
rect 12676 16940 12682 16952
rect 14274 16940 14280 16952
rect 14332 16940 14338 16992
rect 14829 16983 14887 16989
rect 14829 16949 14841 16983
rect 14875 16980 14887 16983
rect 15470 16980 15476 16992
rect 14875 16952 15476 16980
rect 14875 16949 14887 16952
rect 14829 16943 14887 16949
rect 15470 16940 15476 16952
rect 15528 16940 15534 16992
rect 1104 16890 16652 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 16652 16890
rect 1104 16816 16652 16838
rect 2314 16736 2320 16788
rect 2372 16776 2378 16788
rect 3605 16779 3663 16785
rect 2372 16748 3096 16776
rect 2372 16736 2378 16748
rect 3068 16717 3096 16748
rect 3605 16745 3617 16779
rect 3651 16776 3663 16779
rect 3694 16776 3700 16788
rect 3651 16748 3700 16776
rect 3651 16745 3663 16748
rect 3605 16739 3663 16745
rect 3694 16736 3700 16748
rect 3752 16736 3758 16788
rect 5077 16779 5135 16785
rect 5077 16745 5089 16779
rect 5123 16776 5135 16779
rect 5258 16776 5264 16788
rect 5123 16748 5264 16776
rect 5123 16745 5135 16748
rect 5077 16739 5135 16745
rect 5258 16736 5264 16748
rect 5316 16736 5322 16788
rect 5902 16736 5908 16788
rect 5960 16776 5966 16788
rect 6733 16779 6791 16785
rect 6733 16776 6745 16779
rect 5960 16748 6745 16776
rect 5960 16736 5966 16748
rect 6733 16745 6745 16748
rect 6779 16745 6791 16779
rect 6733 16739 6791 16745
rect 8938 16736 8944 16788
rect 8996 16776 9002 16788
rect 9306 16776 9312 16788
rect 8996 16748 9312 16776
rect 8996 16736 9002 16748
rect 9306 16736 9312 16748
rect 9364 16736 9370 16788
rect 9766 16736 9772 16788
rect 9824 16736 9830 16788
rect 10413 16779 10471 16785
rect 10413 16745 10425 16779
rect 10459 16776 10471 16779
rect 10870 16776 10876 16788
rect 10459 16748 10876 16776
rect 10459 16745 10471 16748
rect 10413 16739 10471 16745
rect 10870 16736 10876 16748
rect 10928 16736 10934 16788
rect 12986 16736 12992 16788
rect 13044 16776 13050 16788
rect 15378 16776 15384 16788
rect 13044 16748 15384 16776
rect 13044 16736 13050 16748
rect 15378 16736 15384 16748
rect 15436 16736 15442 16788
rect 3053 16711 3111 16717
rect 3053 16677 3065 16711
rect 3099 16677 3111 16711
rect 10502 16708 10508 16720
rect 3053 16671 3111 16677
rect 9876 16680 10508 16708
rect 1394 16600 1400 16652
rect 1452 16600 1458 16652
rect 4706 16640 4712 16652
rect 4540 16612 4712 16640
rect 1486 16532 1492 16584
rect 1544 16572 1550 16584
rect 1653 16575 1711 16581
rect 1653 16572 1665 16575
rect 1544 16544 1665 16572
rect 1544 16532 1550 16544
rect 1653 16541 1665 16544
rect 1699 16541 1711 16575
rect 1653 16535 1711 16541
rect 3786 16532 3792 16584
rect 3844 16532 3850 16584
rect 4062 16532 4068 16584
rect 4120 16532 4126 16584
rect 4157 16575 4215 16581
rect 4157 16541 4169 16575
rect 4203 16541 4215 16575
rect 4157 16535 4215 16541
rect 2866 16464 2872 16516
rect 2924 16504 2930 16516
rect 3237 16507 3295 16513
rect 3237 16504 3249 16507
rect 2924 16476 3249 16504
rect 2924 16464 2930 16476
rect 3237 16473 3249 16476
rect 3283 16473 3295 16507
rect 3237 16467 3295 16473
rect 3970 16464 3976 16516
rect 4028 16464 4034 16516
rect 4172 16504 4200 16535
rect 4246 16532 4252 16584
rect 4304 16572 4310 16584
rect 4540 16572 4568 16612
rect 4706 16600 4712 16612
rect 4764 16600 4770 16652
rect 5074 16600 5080 16652
rect 5132 16640 5138 16652
rect 5258 16640 5264 16652
rect 5132 16612 5264 16640
rect 5132 16600 5138 16612
rect 5258 16600 5264 16612
rect 5316 16600 5322 16652
rect 9766 16640 9772 16652
rect 9508 16612 9772 16640
rect 4304 16544 4568 16572
rect 4304 16532 4310 16544
rect 4614 16532 4620 16584
rect 4672 16572 4678 16584
rect 5534 16581 5540 16584
rect 4801 16575 4859 16581
rect 4801 16572 4813 16575
rect 4672 16544 4813 16572
rect 4672 16532 4678 16544
rect 4801 16541 4813 16544
rect 4847 16541 4859 16575
rect 4801 16535 4859 16541
rect 4985 16575 5043 16581
rect 4985 16541 4997 16575
rect 5031 16541 5043 16575
rect 4985 16535 5043 16541
rect 5169 16575 5227 16581
rect 5169 16541 5181 16575
rect 5215 16541 5227 16575
rect 5528 16572 5540 16581
rect 5495 16544 5540 16572
rect 5169 16535 5227 16541
rect 5528 16535 5540 16544
rect 4172 16476 4568 16504
rect 4540 16448 4568 16476
rect 4706 16464 4712 16516
rect 4764 16504 4770 16516
rect 5000 16504 5028 16535
rect 4764 16476 5028 16504
rect 4764 16464 4770 16476
rect 2777 16439 2835 16445
rect 2777 16405 2789 16439
rect 2823 16436 2835 16439
rect 3050 16436 3056 16448
rect 2823 16408 3056 16436
rect 2823 16405 2835 16408
rect 2777 16399 2835 16405
rect 3050 16396 3056 16408
rect 3108 16396 3114 16448
rect 3326 16396 3332 16448
rect 3384 16396 3390 16448
rect 3421 16439 3479 16445
rect 3421 16405 3433 16439
rect 3467 16436 3479 16439
rect 3510 16436 3516 16448
rect 3467 16408 3516 16436
rect 3467 16405 3479 16408
rect 3421 16399 3479 16405
rect 3510 16396 3516 16408
rect 3568 16396 3574 16448
rect 4154 16396 4160 16448
rect 4212 16436 4218 16448
rect 4341 16439 4399 16445
rect 4341 16436 4353 16439
rect 4212 16408 4353 16436
rect 4212 16396 4218 16408
rect 4341 16405 4353 16408
rect 4387 16405 4399 16439
rect 4341 16399 4399 16405
rect 4522 16396 4528 16448
rect 4580 16396 4586 16448
rect 5184 16436 5212 16535
rect 5534 16532 5540 16535
rect 5592 16532 5598 16584
rect 8110 16532 8116 16584
rect 8168 16532 8174 16584
rect 9309 16575 9367 16581
rect 9309 16541 9321 16575
rect 9355 16572 9367 16575
rect 9398 16572 9404 16584
rect 9355 16544 9404 16572
rect 9355 16541 9367 16544
rect 9309 16535 9367 16541
rect 9398 16532 9404 16544
rect 9456 16532 9462 16584
rect 9508 16581 9536 16612
rect 9766 16600 9772 16612
rect 9824 16600 9830 16652
rect 9493 16575 9551 16581
rect 9493 16541 9505 16575
rect 9539 16541 9551 16575
rect 9876 16572 9904 16680
rect 10502 16668 10508 16680
rect 10560 16668 10566 16720
rect 10781 16711 10839 16717
rect 10781 16677 10793 16711
rect 10827 16708 10839 16711
rect 11698 16708 11704 16720
rect 10827 16680 11704 16708
rect 10827 16677 10839 16680
rect 10781 16671 10839 16677
rect 11698 16668 11704 16680
rect 11756 16668 11762 16720
rect 13814 16708 13820 16720
rect 13188 16680 13820 16708
rect 10134 16600 10140 16652
rect 10192 16640 10198 16652
rect 10873 16643 10931 16649
rect 10192 16612 10640 16640
rect 10192 16600 10198 16612
rect 9493 16535 9551 16541
rect 9600 16544 9904 16572
rect 5994 16464 6000 16516
rect 6052 16504 6058 16516
rect 7846 16507 7904 16513
rect 7846 16504 7858 16507
rect 6052 16476 7858 16504
rect 6052 16464 6058 16476
rect 7846 16473 7858 16476
rect 7892 16473 7904 16507
rect 7846 16467 7904 16473
rect 9030 16464 9036 16516
rect 9088 16504 9094 16516
rect 9600 16513 9628 16544
rect 9950 16532 9956 16584
rect 10008 16572 10014 16584
rect 10152 16572 10180 16600
rect 10008 16544 10180 16572
rect 10008 16532 10014 16544
rect 10410 16532 10416 16584
rect 10468 16532 10474 16584
rect 10612 16581 10640 16612
rect 10873 16609 10885 16643
rect 10919 16640 10931 16643
rect 11330 16640 11336 16652
rect 10919 16612 11336 16640
rect 10919 16609 10931 16612
rect 10873 16603 10931 16609
rect 11330 16600 11336 16612
rect 11388 16600 11394 16652
rect 10505 16575 10563 16581
rect 10505 16541 10517 16575
rect 10551 16541 10563 16575
rect 10505 16535 10563 16541
rect 10597 16575 10655 16581
rect 10597 16541 10609 16575
rect 10643 16541 10655 16575
rect 10597 16535 10655 16541
rect 10689 16575 10747 16581
rect 10689 16541 10701 16575
rect 10735 16572 10747 16575
rect 10778 16572 10784 16584
rect 10735 16544 10784 16572
rect 10735 16541 10747 16544
rect 10689 16535 10747 16541
rect 9585 16507 9643 16513
rect 9585 16504 9597 16507
rect 9088 16476 9597 16504
rect 9088 16464 9094 16476
rect 9585 16473 9597 16476
rect 9631 16473 9643 16507
rect 9801 16507 9859 16513
rect 9801 16504 9813 16507
rect 9759 16476 9813 16504
rect 9585 16467 9643 16473
rect 9784 16473 9813 16476
rect 9847 16504 9859 16507
rect 9968 16504 9996 16532
rect 9847 16476 9996 16504
rect 9847 16473 9859 16476
rect 9784 16467 9859 16473
rect 6270 16436 6276 16448
rect 5184 16408 6276 16436
rect 6270 16396 6276 16408
rect 6328 16436 6334 16448
rect 6641 16439 6699 16445
rect 6641 16436 6653 16439
rect 6328 16408 6653 16436
rect 6328 16396 6334 16408
rect 6641 16405 6653 16408
rect 6687 16405 6699 16439
rect 6641 16399 6699 16405
rect 9306 16396 9312 16448
rect 9364 16436 9370 16448
rect 9401 16439 9459 16445
rect 9401 16436 9413 16439
rect 9364 16408 9413 16436
rect 9364 16396 9370 16408
rect 9401 16405 9413 16408
rect 9447 16405 9459 16439
rect 9401 16399 9459 16405
rect 9490 16396 9496 16448
rect 9548 16436 9554 16448
rect 9784 16436 9812 16467
rect 10042 16464 10048 16516
rect 10100 16504 10106 16516
rect 10428 16504 10456 16532
rect 10100 16476 10456 16504
rect 10520 16504 10548 16535
rect 10778 16532 10784 16544
rect 10836 16532 10842 16584
rect 12434 16572 12440 16584
rect 10888 16544 12440 16572
rect 10888 16504 10916 16544
rect 12434 16532 12440 16544
rect 12492 16532 12498 16584
rect 13078 16532 13084 16584
rect 13136 16532 13142 16584
rect 13188 16581 13216 16680
rect 13814 16668 13820 16680
rect 13872 16668 13878 16720
rect 15470 16600 15476 16652
rect 15528 16640 15534 16652
rect 15528 16612 15976 16640
rect 15528 16600 15534 16612
rect 13173 16575 13231 16581
rect 13173 16541 13185 16575
rect 13219 16541 13231 16575
rect 13173 16535 13231 16541
rect 13262 16532 13268 16584
rect 13320 16532 13326 16584
rect 13446 16532 13452 16584
rect 13504 16532 13510 16584
rect 13541 16575 13599 16581
rect 13541 16541 13553 16575
rect 13587 16541 13599 16575
rect 13541 16535 13599 16541
rect 13633 16575 13691 16581
rect 13633 16541 13645 16575
rect 13679 16572 13691 16575
rect 13998 16572 14004 16584
rect 13679 16544 14004 16572
rect 13679 16541 13691 16544
rect 13633 16535 13691 16541
rect 10520 16476 10916 16504
rect 10965 16507 11023 16513
rect 10100 16464 10106 16476
rect 10965 16473 10977 16507
rect 11011 16473 11023 16507
rect 10965 16467 11023 16473
rect 9548 16408 9812 16436
rect 9548 16396 9554 16408
rect 9950 16396 9956 16448
rect 10008 16396 10014 16448
rect 10137 16439 10195 16445
rect 10137 16405 10149 16439
rect 10183 16436 10195 16439
rect 10410 16436 10416 16448
rect 10183 16408 10416 16436
rect 10183 16405 10195 16408
rect 10137 16399 10195 16405
rect 10410 16396 10416 16408
rect 10468 16396 10474 16448
rect 10594 16396 10600 16448
rect 10652 16436 10658 16448
rect 10980 16436 11008 16467
rect 11146 16464 11152 16516
rect 11204 16464 11210 16516
rect 13096 16504 13124 16532
rect 13556 16504 13584 16535
rect 13998 16532 14004 16544
rect 14056 16532 14062 16584
rect 14093 16575 14151 16581
rect 14093 16541 14105 16575
rect 14139 16572 14151 16575
rect 14139 16544 14596 16572
rect 14139 16541 14151 16544
rect 14093 16535 14151 16541
rect 14568 16516 14596 16544
rect 14734 16532 14740 16584
rect 14792 16572 14798 16584
rect 15948 16581 15976 16612
rect 15841 16575 15899 16581
rect 15841 16572 15853 16575
rect 14792 16544 15853 16572
rect 14792 16532 14798 16544
rect 15841 16541 15853 16544
rect 15887 16541 15899 16575
rect 15841 16535 15899 16541
rect 15933 16575 15991 16581
rect 15933 16541 15945 16575
rect 15979 16541 15991 16575
rect 15933 16535 15991 16541
rect 16022 16532 16028 16584
rect 16080 16532 16086 16584
rect 16209 16575 16267 16581
rect 16209 16541 16221 16575
rect 16255 16572 16267 16575
rect 16298 16572 16304 16584
rect 16255 16544 16304 16572
rect 16255 16541 16267 16544
rect 16209 16535 16267 16541
rect 13722 16504 13728 16516
rect 13096 16476 13728 16504
rect 13722 16464 13728 16476
rect 13780 16464 13786 16516
rect 13909 16507 13967 16513
rect 13909 16473 13921 16507
rect 13955 16504 13967 16507
rect 14338 16507 14396 16513
rect 14338 16504 14350 16507
rect 13955 16476 14350 16504
rect 13955 16473 13967 16476
rect 13909 16467 13967 16473
rect 14338 16473 14350 16476
rect 14384 16473 14396 16507
rect 14338 16467 14396 16473
rect 14550 16464 14556 16516
rect 14608 16464 14614 16516
rect 14826 16464 14832 16516
rect 14884 16504 14890 16516
rect 15102 16504 15108 16516
rect 14884 16476 15108 16504
rect 14884 16464 14890 16476
rect 15102 16464 15108 16476
rect 15160 16464 15166 16516
rect 15746 16464 15752 16516
rect 15804 16504 15810 16516
rect 16224 16504 16252 16535
rect 16298 16532 16304 16544
rect 16356 16532 16362 16584
rect 15804 16476 16252 16504
rect 15804 16464 15810 16476
rect 10652 16408 11008 16436
rect 11333 16439 11391 16445
rect 10652 16396 10658 16408
rect 11333 16405 11345 16439
rect 11379 16436 11391 16439
rect 11882 16436 11888 16448
rect 11379 16408 11888 16436
rect 11379 16405 11391 16408
rect 11333 16399 11391 16405
rect 11882 16396 11888 16408
rect 11940 16396 11946 16448
rect 12526 16396 12532 16448
rect 12584 16436 12590 16448
rect 12894 16436 12900 16448
rect 12584 16408 12900 16436
rect 12584 16396 12590 16408
rect 12894 16396 12900 16408
rect 12952 16396 12958 16448
rect 13081 16439 13139 16445
rect 13081 16405 13093 16439
rect 13127 16436 13139 16439
rect 13354 16436 13360 16448
rect 13127 16408 13360 16436
rect 13127 16405 13139 16408
rect 13081 16399 13139 16405
rect 13354 16396 13360 16408
rect 13412 16396 13418 16448
rect 13998 16396 14004 16448
rect 14056 16436 14062 16448
rect 15010 16436 15016 16448
rect 14056 16408 15016 16436
rect 14056 16396 14062 16408
rect 15010 16396 15016 16408
rect 15068 16436 15074 16448
rect 15473 16439 15531 16445
rect 15473 16436 15485 16439
rect 15068 16408 15485 16436
rect 15068 16396 15074 16408
rect 15473 16405 15485 16408
rect 15519 16405 15531 16439
rect 15473 16399 15531 16405
rect 15562 16396 15568 16448
rect 15620 16396 15626 16448
rect 1104 16346 16652 16368
rect 1104 16294 4874 16346
rect 4926 16294 4938 16346
rect 4990 16294 5002 16346
rect 5054 16294 5066 16346
rect 5118 16294 5130 16346
rect 5182 16294 16652 16346
rect 1104 16272 16652 16294
rect 2958 16192 2964 16244
rect 3016 16232 3022 16244
rect 3145 16235 3203 16241
rect 3145 16232 3157 16235
rect 3016 16204 3157 16232
rect 3016 16192 3022 16204
rect 3145 16201 3157 16204
rect 3191 16201 3203 16235
rect 3145 16195 3203 16201
rect 3510 16192 3516 16244
rect 3568 16192 3574 16244
rect 3970 16192 3976 16244
rect 4028 16192 4034 16244
rect 4433 16235 4491 16241
rect 4433 16201 4445 16235
rect 4479 16232 4491 16235
rect 4614 16232 4620 16244
rect 4479 16204 4620 16232
rect 4479 16201 4491 16204
rect 4433 16195 4491 16201
rect 4614 16192 4620 16204
rect 4672 16192 4678 16244
rect 5902 16232 5908 16244
rect 5000 16204 5908 16232
rect 3326 16124 3332 16176
rect 3384 16164 3390 16176
rect 5000 16173 5028 16204
rect 5902 16192 5908 16204
rect 5960 16192 5966 16244
rect 5994 16192 6000 16244
rect 6052 16192 6058 16244
rect 9030 16192 9036 16244
rect 9088 16232 9094 16244
rect 9125 16235 9183 16241
rect 9125 16232 9137 16235
rect 9088 16204 9137 16232
rect 9088 16192 9094 16204
rect 9125 16201 9137 16204
rect 9171 16201 9183 16235
rect 9125 16195 9183 16201
rect 9398 16192 9404 16244
rect 9456 16192 9462 16244
rect 9582 16192 9588 16244
rect 9640 16192 9646 16244
rect 9766 16192 9772 16244
rect 9824 16232 9830 16244
rect 10873 16235 10931 16241
rect 10873 16232 10885 16235
rect 9824 16204 10885 16232
rect 9824 16192 9830 16204
rect 10873 16201 10885 16204
rect 10919 16201 10931 16235
rect 10873 16195 10931 16201
rect 11054 16192 11060 16244
rect 11112 16232 11118 16244
rect 11333 16235 11391 16241
rect 11333 16232 11345 16235
rect 11112 16204 11345 16232
rect 11112 16192 11118 16204
rect 11333 16201 11345 16204
rect 11379 16201 11391 16235
rect 11333 16195 11391 16201
rect 11514 16192 11520 16244
rect 11572 16192 11578 16244
rect 12621 16235 12679 16241
rect 12621 16201 12633 16235
rect 12667 16232 12679 16235
rect 15286 16232 15292 16244
rect 12667 16204 15292 16232
rect 12667 16201 12679 16204
rect 12621 16195 12679 16201
rect 15286 16192 15292 16204
rect 15344 16192 15350 16244
rect 4985 16167 5043 16173
rect 3384 16136 4660 16164
rect 3384 16124 3390 16136
rect 1394 16056 1400 16108
rect 1452 16056 1458 16108
rect 1670 16105 1676 16108
rect 1664 16059 1676 16105
rect 1670 16056 1676 16059
rect 1728 16056 1734 16108
rect 2038 16056 2044 16108
rect 2096 16096 2102 16108
rect 2869 16099 2927 16105
rect 2869 16096 2881 16099
rect 2096 16068 2881 16096
rect 2096 16056 2102 16068
rect 2869 16065 2881 16068
rect 2915 16065 2927 16099
rect 2869 16059 2927 16065
rect 3053 16099 3111 16105
rect 3053 16065 3065 16099
rect 3099 16065 3111 16099
rect 3053 16059 3111 16065
rect 3068 16028 3096 16059
rect 3142 16056 3148 16108
rect 3200 16096 3206 16108
rect 3237 16099 3295 16105
rect 3237 16096 3249 16099
rect 3200 16068 3249 16096
rect 3200 16056 3206 16068
rect 3237 16065 3249 16068
rect 3283 16065 3295 16099
rect 3237 16059 3295 16065
rect 3421 16099 3479 16105
rect 3421 16065 3433 16099
rect 3467 16096 3479 16099
rect 3602 16096 3608 16108
rect 3467 16068 3608 16096
rect 3467 16065 3479 16068
rect 3421 16059 3479 16065
rect 3602 16056 3608 16068
rect 3660 16096 3666 16108
rect 3697 16099 3755 16105
rect 3697 16096 3709 16099
rect 3660 16068 3709 16096
rect 3660 16056 3666 16068
rect 3697 16065 3709 16068
rect 3743 16065 3755 16099
rect 3697 16059 3755 16065
rect 3881 16099 3939 16105
rect 3881 16065 3893 16099
rect 3927 16096 3939 16099
rect 4062 16096 4068 16108
rect 3927 16068 4068 16096
rect 3927 16065 3939 16068
rect 3881 16059 3939 16065
rect 3896 16028 3924 16059
rect 4062 16056 4068 16068
rect 4120 16056 4126 16108
rect 4246 16056 4252 16108
rect 4304 16056 4310 16108
rect 4338 16056 4344 16108
rect 4396 16056 4402 16108
rect 4632 16105 4660 16136
rect 4985 16133 4997 16167
rect 5031 16133 5043 16167
rect 4985 16127 5043 16133
rect 5074 16124 5080 16176
rect 5132 16164 5138 16176
rect 5185 16167 5243 16173
rect 5185 16164 5197 16167
rect 5132 16136 5197 16164
rect 5132 16124 5138 16136
rect 5185 16133 5197 16136
rect 5231 16164 5243 16167
rect 5626 16164 5632 16176
rect 5231 16136 5632 16164
rect 5231 16133 5243 16136
rect 5185 16127 5243 16133
rect 5626 16124 5632 16136
rect 5684 16124 5690 16176
rect 5718 16124 5724 16176
rect 5776 16164 5782 16176
rect 5813 16167 5871 16173
rect 5813 16164 5825 16167
rect 5776 16136 5825 16164
rect 5776 16124 5782 16136
rect 5813 16133 5825 16136
rect 5859 16164 5871 16167
rect 6454 16164 6460 16176
rect 5859 16136 6460 16164
rect 5859 16133 5871 16136
rect 5813 16127 5871 16133
rect 6454 16124 6460 16136
rect 6512 16164 6518 16176
rect 7009 16167 7067 16173
rect 7009 16164 7021 16167
rect 6512 16136 7021 16164
rect 6512 16124 6518 16136
rect 7009 16133 7021 16136
rect 7055 16133 7067 16167
rect 9600 16164 9628 16192
rect 9600 16136 9904 16164
rect 7009 16127 7067 16133
rect 4617 16099 4675 16105
rect 4617 16065 4629 16099
rect 4663 16065 4675 16099
rect 4617 16059 4675 16065
rect 4706 16056 4712 16108
rect 4764 16096 4770 16108
rect 5092 16096 5120 16124
rect 4764 16068 5120 16096
rect 5445 16099 5503 16105
rect 4764 16056 4770 16068
rect 5445 16065 5457 16099
rect 5491 16096 5503 16099
rect 7285 16099 7343 16105
rect 7285 16096 7297 16099
rect 5491 16068 7297 16096
rect 5491 16065 5503 16068
rect 5445 16059 5503 16065
rect 7285 16065 7297 16068
rect 7331 16065 7343 16099
rect 7285 16059 7343 16065
rect 3068 16000 3924 16028
rect 3970 15988 3976 16040
rect 4028 16028 4034 16040
rect 4801 16031 4859 16037
rect 4801 16028 4813 16031
rect 4028 16000 4813 16028
rect 4028 15988 4034 16000
rect 4801 15997 4813 16000
rect 4847 15997 4859 16031
rect 4801 15991 4859 15997
rect 2774 15920 2780 15972
rect 2832 15960 2838 15972
rect 3602 15960 3608 15972
rect 2832 15932 3608 15960
rect 2832 15920 2838 15932
rect 3602 15920 3608 15932
rect 3660 15960 3666 15972
rect 4338 15960 4344 15972
rect 3660 15932 4344 15960
rect 3660 15920 3666 15932
rect 4338 15920 4344 15932
rect 4396 15920 4402 15972
rect 4982 15960 4988 15972
rect 4448 15932 4988 15960
rect 2958 15852 2964 15904
rect 3016 15892 3022 15904
rect 4448 15892 4476 15932
rect 4982 15920 4988 15932
rect 5040 15920 5046 15972
rect 5353 15963 5411 15969
rect 5353 15929 5365 15963
rect 5399 15960 5411 15963
rect 5460 15960 5488 16059
rect 7374 16056 7380 16108
rect 7432 16096 7438 16108
rect 7469 16099 7527 16105
rect 7469 16096 7481 16099
rect 7432 16068 7481 16096
rect 7432 16056 7438 16068
rect 7469 16065 7481 16068
rect 7515 16065 7527 16099
rect 7469 16059 7527 16065
rect 8754 16056 8760 16108
rect 8812 16056 8818 16108
rect 8938 16056 8944 16108
rect 8996 16056 9002 16108
rect 9122 16056 9128 16108
rect 9180 16096 9186 16108
rect 9309 16099 9367 16105
rect 9309 16096 9321 16099
rect 9180 16068 9321 16096
rect 9180 16056 9186 16068
rect 9309 16065 9321 16068
rect 9355 16065 9367 16099
rect 9309 16059 9367 16065
rect 9582 16056 9588 16108
rect 9640 16056 9646 16108
rect 9674 16056 9680 16108
rect 9732 16056 9738 16108
rect 9876 16105 9904 16136
rect 10134 16124 10140 16176
rect 10192 16164 10198 16176
rect 10965 16167 11023 16173
rect 10965 16164 10977 16167
rect 10192 16136 10977 16164
rect 10192 16124 10198 16136
rect 10965 16133 10977 16136
rect 11011 16133 11023 16167
rect 10965 16127 11023 16133
rect 11195 16133 11253 16139
rect 11195 16130 11207 16133
rect 9861 16099 9919 16105
rect 9861 16065 9873 16099
rect 9907 16065 9919 16099
rect 10413 16099 10471 16105
rect 10413 16096 10425 16099
rect 9861 16059 9919 16065
rect 9968 16068 10425 16096
rect 5534 15960 5540 15972
rect 5399 15932 5540 15960
rect 5399 15929 5411 15932
rect 5353 15923 5411 15929
rect 5534 15920 5540 15932
rect 5592 15920 5598 15972
rect 5718 15920 5724 15972
rect 5776 15960 5782 15972
rect 6641 15963 6699 15969
rect 6641 15960 6653 15963
rect 5776 15932 6653 15960
rect 5776 15920 5782 15932
rect 6641 15929 6653 15932
rect 6687 15929 6699 15963
rect 7653 15963 7711 15969
rect 7653 15960 7665 15963
rect 6641 15923 6699 15929
rect 7024 15932 7665 15960
rect 3016 15864 4476 15892
rect 3016 15852 3022 15864
rect 4522 15852 4528 15904
rect 4580 15892 4586 15904
rect 4890 15892 4896 15904
rect 4580 15864 4896 15892
rect 4580 15852 4586 15864
rect 4890 15852 4896 15864
rect 4948 15852 4954 15904
rect 5169 15895 5227 15901
rect 5169 15861 5181 15895
rect 5215 15892 5227 15895
rect 5626 15892 5632 15904
rect 5215 15864 5632 15892
rect 5215 15861 5227 15864
rect 5169 15855 5227 15861
rect 5626 15852 5632 15864
rect 5684 15852 5690 15904
rect 5810 15852 5816 15904
rect 5868 15852 5874 15904
rect 7024 15901 7052 15932
rect 7653 15929 7665 15932
rect 7699 15929 7711 15963
rect 8956 15960 8984 16056
rect 9692 15960 9720 16056
rect 9968 16040 9996 16068
rect 10413 16065 10425 16068
rect 10459 16096 10471 16099
rect 10505 16099 10563 16105
rect 10505 16096 10517 16099
rect 10459 16068 10517 16096
rect 10459 16065 10471 16068
rect 10413 16059 10471 16065
rect 10505 16065 10517 16068
rect 10551 16065 10563 16099
rect 10505 16059 10563 16065
rect 10686 16056 10692 16108
rect 10744 16096 10750 16108
rect 11184 16099 11207 16130
rect 11241 16099 11253 16133
rect 11422 16124 11428 16176
rect 11480 16164 11486 16176
rect 11669 16167 11727 16173
rect 11669 16164 11681 16167
rect 11480 16136 11681 16164
rect 11480 16124 11486 16136
rect 11669 16133 11681 16136
rect 11715 16133 11727 16167
rect 11669 16127 11727 16133
rect 11882 16124 11888 16176
rect 11940 16124 11946 16176
rect 12345 16167 12403 16173
rect 12345 16133 12357 16167
rect 12391 16164 12403 16167
rect 13081 16167 13139 16173
rect 13081 16164 13093 16167
rect 12391 16136 13093 16164
rect 12391 16133 12403 16136
rect 12345 16127 12403 16133
rect 13081 16133 13093 16136
rect 13127 16164 13139 16167
rect 13127 16136 13400 16164
rect 13127 16133 13139 16136
rect 13081 16127 13139 16133
rect 11184 16096 11253 16099
rect 10744 16093 11253 16096
rect 10744 16068 11212 16093
rect 10744 16056 10750 16068
rect 12250 16056 12256 16108
rect 12308 16056 12314 16108
rect 12805 16099 12863 16105
rect 12805 16065 12817 16099
rect 12851 16065 12863 16099
rect 12805 16059 12863 16065
rect 12897 16099 12955 16105
rect 12897 16065 12909 16099
rect 12943 16065 12955 16099
rect 12897 16059 12955 16065
rect 9769 16031 9827 16037
rect 9769 15997 9781 16031
rect 9815 16028 9827 16031
rect 9950 16028 9956 16040
rect 9815 16000 9956 16028
rect 9815 15997 9827 16000
rect 9769 15991 9827 15997
rect 9950 15988 9956 16000
rect 10008 15988 10014 16040
rect 10134 15988 10140 16040
rect 10192 16028 10198 16040
rect 10321 16031 10379 16037
rect 10321 16028 10333 16031
rect 10192 16000 10333 16028
rect 10192 15988 10198 16000
rect 10321 15997 10333 16000
rect 10367 16028 10379 16031
rect 10367 16000 10548 16028
rect 10367 15997 10379 16000
rect 10321 15991 10379 15997
rect 10520 15960 10548 16000
rect 10594 15988 10600 16040
rect 10652 15988 10658 16040
rect 10870 15988 10876 16040
rect 10928 16028 10934 16040
rect 11514 16028 11520 16040
rect 10928 16000 11520 16028
rect 10928 15988 10934 16000
rect 11514 15988 11520 16000
rect 11572 15988 11578 16040
rect 12526 16028 12532 16040
rect 12406 16000 12532 16028
rect 11330 15960 11336 15972
rect 8956 15932 9628 15960
rect 9692 15932 10456 15960
rect 10520 15932 11336 15960
rect 7653 15923 7711 15929
rect 7009 15895 7067 15901
rect 7009 15861 7021 15895
rect 7055 15861 7067 15895
rect 7009 15855 7067 15861
rect 7190 15852 7196 15904
rect 7248 15852 7254 15904
rect 8938 15852 8944 15904
rect 8996 15852 9002 15904
rect 9600 15892 9628 15932
rect 9950 15892 9956 15904
rect 9600 15864 9956 15892
rect 9950 15852 9956 15864
rect 10008 15852 10014 15904
rect 10042 15852 10048 15904
rect 10100 15852 10106 15904
rect 10318 15852 10324 15904
rect 10376 15852 10382 15904
rect 10428 15892 10456 15932
rect 11330 15920 11336 15932
rect 11388 15960 11394 15972
rect 12406 15960 12434 16000
rect 12526 15988 12532 16000
rect 12584 15988 12590 16040
rect 11388 15932 12434 15960
rect 12820 15960 12848 16059
rect 12912 16028 12940 16059
rect 13262 16056 13268 16108
rect 13320 16096 13326 16108
rect 13372 16105 13400 16136
rect 13446 16124 13452 16176
rect 13504 16164 13510 16176
rect 14001 16167 14059 16173
rect 14001 16164 14013 16167
rect 13504 16136 14013 16164
rect 13504 16124 13510 16136
rect 14001 16133 14013 16136
rect 14047 16133 14059 16167
rect 14001 16127 14059 16133
rect 14090 16124 14096 16176
rect 14148 16164 14154 16176
rect 14369 16167 14427 16173
rect 14369 16164 14381 16167
rect 14148 16136 14381 16164
rect 14148 16124 14154 16136
rect 14369 16133 14381 16136
rect 14415 16133 14427 16167
rect 14918 16164 14924 16176
rect 14369 16127 14427 16133
rect 14752 16136 14924 16164
rect 13357 16099 13415 16105
rect 13357 16096 13369 16099
rect 13320 16068 13369 16096
rect 13320 16056 13326 16068
rect 13357 16065 13369 16068
rect 13403 16065 13415 16099
rect 13357 16059 13415 16065
rect 13541 16099 13599 16105
rect 13541 16065 13553 16099
rect 13587 16065 13599 16099
rect 13541 16059 13599 16065
rect 13446 16028 13452 16040
rect 12912 16000 13452 16028
rect 13446 15988 13452 16000
rect 13504 16028 13510 16040
rect 13556 16028 13584 16059
rect 13906 16056 13912 16108
rect 13964 16096 13970 16108
rect 14185 16099 14243 16105
rect 14185 16096 14197 16099
rect 13964 16068 14197 16096
rect 13964 16056 13970 16068
rect 14185 16065 14197 16068
rect 14231 16065 14243 16099
rect 14185 16059 14243 16065
rect 14642 16056 14648 16108
rect 14700 16056 14706 16108
rect 14752 16105 14780 16136
rect 14918 16124 14924 16136
rect 14976 16124 14982 16176
rect 15188 16167 15246 16173
rect 15188 16133 15200 16167
rect 15234 16164 15246 16167
rect 15562 16164 15568 16176
rect 15234 16136 15568 16164
rect 15234 16133 15246 16136
rect 15188 16127 15246 16133
rect 15562 16124 15568 16136
rect 15620 16124 15626 16176
rect 14737 16099 14795 16105
rect 14737 16065 14749 16099
rect 14783 16065 14795 16099
rect 15654 16096 15660 16108
rect 14737 16059 14795 16065
rect 14844 16068 15660 16096
rect 13504 16000 13584 16028
rect 14461 16031 14519 16037
rect 13504 15988 13510 16000
rect 14461 15997 14473 16031
rect 14507 16028 14519 16031
rect 14844 16028 14872 16068
rect 15654 16056 15660 16068
rect 15712 16056 15718 16108
rect 14507 16000 14872 16028
rect 14921 16031 14979 16037
rect 14507 15997 14519 16000
rect 14461 15991 14519 15997
rect 14921 15997 14933 16031
rect 14967 15997 14979 16031
rect 14921 15991 14979 15997
rect 13633 15963 13691 15969
rect 12820 15932 13584 15960
rect 11388 15920 11394 15932
rect 10505 15895 10563 15901
rect 10505 15892 10517 15895
rect 10428 15864 10517 15892
rect 10505 15861 10517 15864
rect 10551 15861 10563 15895
rect 10505 15855 10563 15861
rect 10778 15852 10784 15904
rect 10836 15892 10842 15904
rect 11149 15895 11207 15901
rect 11149 15892 11161 15895
rect 10836 15864 11161 15892
rect 10836 15852 10842 15864
rect 11149 15861 11161 15864
rect 11195 15861 11207 15895
rect 11149 15855 11207 15861
rect 11698 15852 11704 15904
rect 11756 15852 11762 15904
rect 13170 15852 13176 15904
rect 13228 15852 13234 15904
rect 13556 15892 13584 15932
rect 13633 15929 13645 15963
rect 13679 15960 13691 15963
rect 14090 15960 14096 15972
rect 13679 15932 14096 15960
rect 13679 15929 13691 15932
rect 13633 15923 13691 15929
rect 14090 15920 14096 15932
rect 14148 15920 14154 15972
rect 14550 15920 14556 15972
rect 14608 15960 14614 15972
rect 14936 15960 14964 15991
rect 14608 15932 14964 15960
rect 14608 15920 14614 15932
rect 15838 15892 15844 15904
rect 13556 15864 15844 15892
rect 15838 15852 15844 15864
rect 15896 15892 15902 15904
rect 16022 15892 16028 15904
rect 15896 15864 16028 15892
rect 15896 15852 15902 15864
rect 16022 15852 16028 15864
rect 16080 15892 16086 15904
rect 16301 15895 16359 15901
rect 16301 15892 16313 15895
rect 16080 15864 16313 15892
rect 16080 15852 16086 15864
rect 16301 15861 16313 15864
rect 16347 15861 16359 15895
rect 16301 15855 16359 15861
rect 1104 15802 16652 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 16652 15802
rect 1104 15728 16652 15750
rect 1581 15691 1639 15697
rect 1581 15657 1593 15691
rect 1627 15688 1639 15691
rect 1670 15688 1676 15700
rect 1627 15660 1676 15688
rect 1627 15657 1639 15660
rect 1581 15651 1639 15657
rect 1670 15648 1676 15660
rect 1728 15648 1734 15700
rect 1762 15648 1768 15700
rect 1820 15688 1826 15700
rect 2682 15688 2688 15700
rect 1820 15660 2688 15688
rect 1820 15648 1826 15660
rect 2682 15648 2688 15660
rect 2740 15648 2746 15700
rect 2777 15691 2835 15697
rect 2777 15657 2789 15691
rect 2823 15688 2835 15691
rect 3421 15691 3479 15697
rect 2823 15660 3080 15688
rect 2823 15657 2835 15660
rect 2777 15651 2835 15657
rect 3052 15632 3080 15660
rect 3421 15657 3433 15691
rect 3467 15688 3479 15691
rect 3878 15688 3884 15700
rect 3467 15660 3884 15688
rect 3467 15657 3479 15660
rect 3421 15651 3479 15657
rect 3878 15648 3884 15660
rect 3936 15648 3942 15700
rect 4614 15648 4620 15700
rect 4672 15688 4678 15700
rect 4709 15691 4767 15697
rect 4709 15688 4721 15691
rect 4672 15660 4721 15688
rect 4672 15648 4678 15660
rect 4709 15657 4721 15660
rect 4755 15657 4767 15691
rect 4709 15651 4767 15657
rect 4798 15648 4804 15700
rect 4856 15648 4862 15700
rect 5350 15648 5356 15700
rect 5408 15688 5414 15700
rect 5445 15691 5503 15697
rect 5445 15688 5457 15691
rect 5408 15660 5457 15688
rect 5408 15648 5414 15660
rect 5445 15657 5457 15660
rect 5491 15657 5503 15691
rect 5445 15651 5503 15657
rect 5626 15648 5632 15700
rect 5684 15688 5690 15700
rect 6270 15688 6276 15700
rect 5684 15660 6276 15688
rect 5684 15648 5690 15660
rect 6270 15648 6276 15660
rect 6328 15648 6334 15700
rect 6641 15691 6699 15697
rect 6641 15657 6653 15691
rect 6687 15688 6699 15691
rect 6914 15688 6920 15700
rect 6687 15660 6920 15688
rect 6687 15657 6699 15660
rect 6641 15651 6699 15657
rect 6914 15648 6920 15660
rect 6972 15688 6978 15700
rect 7374 15688 7380 15700
rect 6972 15660 7380 15688
rect 6972 15648 6978 15660
rect 7374 15648 7380 15660
rect 7432 15648 7438 15700
rect 8113 15691 8171 15697
rect 8113 15657 8125 15691
rect 8159 15688 8171 15691
rect 8202 15688 8208 15700
rect 8159 15660 8208 15688
rect 8159 15657 8171 15660
rect 8113 15651 8171 15657
rect 8202 15648 8208 15660
rect 8260 15648 8266 15700
rect 8297 15691 8355 15697
rect 8297 15657 8309 15691
rect 8343 15688 8355 15691
rect 8570 15688 8576 15700
rect 8343 15660 8576 15688
rect 8343 15657 8355 15660
rect 8297 15651 8355 15657
rect 8570 15648 8576 15660
rect 8628 15648 8634 15700
rect 9674 15688 9680 15700
rect 8772 15660 9680 15688
rect 2961 15623 3019 15629
rect 2961 15589 2973 15623
rect 3007 15589 3019 15623
rect 2961 15583 3019 15589
rect 2133 15555 2191 15561
rect 2133 15521 2145 15555
rect 2179 15552 2191 15555
rect 2774 15552 2780 15564
rect 2179 15524 2780 15552
rect 2179 15521 2191 15524
rect 2133 15515 2191 15521
rect 2774 15512 2780 15524
rect 2832 15512 2838 15564
rect 2976 15552 3004 15583
rect 3050 15580 3056 15632
rect 3108 15580 3114 15632
rect 3602 15580 3608 15632
rect 3660 15620 3666 15632
rect 4525 15623 4583 15629
rect 3660 15592 4108 15620
rect 3660 15580 3666 15592
rect 3326 15552 3332 15564
rect 2976 15524 3332 15552
rect 3326 15512 3332 15524
rect 3384 15552 3390 15564
rect 4080 15552 4108 15592
rect 4525 15589 4537 15623
rect 4571 15620 4583 15623
rect 4816 15620 4844 15648
rect 4571 15592 4844 15620
rect 5460 15592 6408 15620
rect 4571 15589 4583 15592
rect 4525 15583 4583 15589
rect 5460 15564 5488 15592
rect 4709 15555 4767 15561
rect 4709 15552 4721 15555
rect 3384 15524 4016 15552
rect 4080 15524 4721 15552
rect 3384 15512 3390 15524
rect 2409 15487 2467 15493
rect 2409 15453 2421 15487
rect 2455 15453 2467 15487
rect 2409 15447 2467 15453
rect 2685 15487 2743 15493
rect 2685 15453 2697 15487
rect 2731 15484 2743 15487
rect 2866 15484 2872 15496
rect 2731 15456 2872 15484
rect 2731 15453 2743 15456
rect 2685 15447 2743 15453
rect 1765 15419 1823 15425
rect 1765 15385 1777 15419
rect 1811 15416 1823 15419
rect 1946 15416 1952 15428
rect 1811 15388 1952 15416
rect 1811 15385 1823 15388
rect 1765 15379 1823 15385
rect 1946 15376 1952 15388
rect 2004 15376 2010 15428
rect 2424 15416 2452 15447
rect 2866 15444 2872 15456
rect 2924 15444 2930 15496
rect 3418 15444 3424 15496
rect 3476 15484 3482 15496
rect 3789 15487 3847 15493
rect 3789 15484 3801 15487
rect 3476 15456 3801 15484
rect 3476 15444 3482 15456
rect 3789 15453 3801 15456
rect 3835 15453 3847 15487
rect 3789 15447 3847 15453
rect 3878 15444 3884 15496
rect 3936 15444 3942 15496
rect 3988 15493 4016 15524
rect 4709 15521 4721 15524
rect 4755 15521 4767 15555
rect 4709 15515 4767 15521
rect 4798 15512 4804 15564
rect 4856 15552 4862 15564
rect 4856 15524 5304 15552
rect 4856 15512 4862 15524
rect 3973 15487 4031 15493
rect 3973 15453 3985 15487
rect 4019 15453 4031 15487
rect 3973 15447 4031 15453
rect 4062 15444 4068 15496
rect 4120 15444 4126 15496
rect 4157 15487 4215 15493
rect 4157 15453 4169 15487
rect 4203 15453 4215 15487
rect 4157 15447 4215 15453
rect 3694 15416 3700 15428
rect 2424 15388 3700 15416
rect 3694 15376 3700 15388
rect 3752 15376 3758 15428
rect 3896 15416 3924 15444
rect 4172 15416 4200 15447
rect 4890 15444 4896 15496
rect 4948 15444 4954 15496
rect 4982 15444 4988 15496
rect 5040 15444 5046 15496
rect 5166 15444 5172 15496
rect 5224 15444 5230 15496
rect 5276 15484 5304 15524
rect 5442 15512 5448 15564
rect 5500 15512 5506 15564
rect 5552 15552 5764 15560
rect 5552 15532 6041 15552
rect 5552 15484 5580 15532
rect 5736 15524 6041 15532
rect 5276 15456 5580 15484
rect 5626 15444 5632 15496
rect 5684 15444 5690 15496
rect 5902 15444 5908 15496
rect 5960 15444 5966 15496
rect 6013 15493 6041 15524
rect 5998 15487 6056 15493
rect 5998 15453 6010 15487
rect 6044 15453 6056 15487
rect 5998 15447 6056 15453
rect 6270 15444 6276 15496
rect 6328 15444 6334 15496
rect 6380 15493 6408 15592
rect 8021 15555 8079 15561
rect 8021 15521 8033 15555
rect 8067 15552 8079 15555
rect 8110 15552 8116 15564
rect 8067 15524 8116 15552
rect 8067 15521 8079 15524
rect 8021 15515 8079 15521
rect 8110 15512 8116 15524
rect 8168 15512 8174 15564
rect 6370 15487 6428 15493
rect 6370 15453 6382 15487
rect 6416 15453 6428 15487
rect 6370 15447 6428 15453
rect 7190 15444 7196 15496
rect 7248 15484 7254 15496
rect 7754 15487 7812 15493
rect 7754 15484 7766 15487
rect 7248 15456 7766 15484
rect 7248 15444 7254 15456
rect 7754 15453 7766 15456
rect 7800 15453 7812 15487
rect 7754 15447 7812 15453
rect 8386 15444 8392 15496
rect 8444 15484 8450 15496
rect 8665 15487 8723 15493
rect 8665 15484 8677 15487
rect 8444 15456 8677 15484
rect 8444 15444 8450 15456
rect 8665 15453 8677 15456
rect 8711 15453 8723 15487
rect 8772 15484 8800 15660
rect 9674 15648 9680 15660
rect 9732 15648 9738 15700
rect 9766 15648 9772 15700
rect 9824 15648 9830 15700
rect 9950 15648 9956 15700
rect 10008 15688 10014 15700
rect 10502 15688 10508 15700
rect 10008 15660 10508 15688
rect 10008 15648 10014 15660
rect 10502 15648 10508 15660
rect 10560 15648 10566 15700
rect 12989 15691 13047 15697
rect 12989 15688 13001 15691
rect 12084 15660 13001 15688
rect 9125 15623 9183 15629
rect 9125 15589 9137 15623
rect 9171 15620 9183 15623
rect 10594 15620 10600 15632
rect 9171 15592 10600 15620
rect 9171 15589 9183 15592
rect 9125 15583 9183 15589
rect 10594 15580 10600 15592
rect 10652 15620 10658 15632
rect 10870 15620 10876 15632
rect 10652 15592 10876 15620
rect 10652 15580 10658 15592
rect 10870 15580 10876 15592
rect 10928 15580 10934 15632
rect 11698 15620 11704 15632
rect 11348 15592 11704 15620
rect 8846 15512 8852 15564
rect 8904 15552 8910 15564
rect 9217 15555 9275 15561
rect 8904 15541 9168 15552
rect 9217 15541 9229 15555
rect 8904 15524 9229 15541
rect 8904 15512 8910 15524
rect 9140 15521 9229 15524
rect 9263 15521 9275 15555
rect 9446 15552 9628 15560
rect 10778 15552 10784 15564
rect 9140 15515 9275 15521
rect 9350 15532 10784 15552
rect 9350 15524 9474 15532
rect 9600 15524 10784 15532
rect 9140 15513 9260 15515
rect 8941 15487 8999 15493
rect 8941 15484 8953 15487
rect 8772 15456 8953 15484
rect 8665 15447 8723 15453
rect 8941 15453 8953 15456
rect 8987 15453 8999 15487
rect 8941 15447 8999 15453
rect 9033 15487 9091 15493
rect 9033 15453 9045 15487
rect 9079 15484 9091 15487
rect 9350 15484 9378 15524
rect 10778 15512 10784 15524
rect 10836 15512 10842 15564
rect 9490 15484 9496 15496
rect 9079 15456 9378 15484
rect 9452 15456 9496 15484
rect 9079 15453 9091 15456
rect 9033 15447 9091 15453
rect 9490 15444 9496 15456
rect 9548 15444 9554 15496
rect 9631 15487 9689 15493
rect 9631 15453 9643 15487
rect 9677 15453 9689 15487
rect 9631 15447 9689 15453
rect 3896 15388 4200 15416
rect 5810 15376 5816 15428
rect 5868 15376 5874 15428
rect 6178 15376 6184 15428
rect 6236 15376 6242 15428
rect 9646 15416 9674 15447
rect 9766 15444 9772 15496
rect 9824 15484 9830 15496
rect 9861 15487 9919 15493
rect 9861 15484 9873 15487
rect 9824 15456 9873 15484
rect 9824 15444 9830 15456
rect 9861 15453 9873 15456
rect 9907 15453 9919 15487
rect 9861 15447 9919 15453
rect 9950 15444 9956 15496
rect 10008 15444 10014 15496
rect 10045 15487 10103 15493
rect 10045 15453 10057 15487
rect 10091 15484 10103 15487
rect 10134 15484 10140 15496
rect 10091 15456 10140 15484
rect 10091 15453 10103 15456
rect 10045 15447 10103 15453
rect 10134 15444 10140 15456
rect 10192 15444 10198 15496
rect 10229 15487 10287 15493
rect 10229 15453 10241 15487
rect 10275 15484 10287 15487
rect 10318 15484 10324 15496
rect 10275 15456 10324 15484
rect 10275 15453 10287 15456
rect 10229 15447 10287 15453
rect 10318 15444 10324 15456
rect 10376 15444 10382 15496
rect 10410 15444 10416 15496
rect 10468 15444 10474 15496
rect 10502 15444 10508 15496
rect 10560 15444 10566 15496
rect 10594 15444 10600 15496
rect 10652 15444 10658 15496
rect 10962 15444 10968 15496
rect 11020 15484 11026 15496
rect 11348 15493 11376 15592
rect 11698 15580 11704 15592
rect 11756 15580 11762 15632
rect 11517 15555 11575 15561
rect 11517 15521 11529 15555
rect 11563 15552 11575 15555
rect 11882 15552 11888 15564
rect 11563 15524 11888 15552
rect 11563 15521 11575 15524
rect 11517 15515 11575 15521
rect 11882 15512 11888 15524
rect 11940 15512 11946 15564
rect 11149 15487 11207 15493
rect 11149 15484 11161 15487
rect 11020 15456 11161 15484
rect 11020 15444 11026 15456
rect 11149 15453 11161 15456
rect 11195 15453 11207 15487
rect 11149 15447 11207 15453
rect 11333 15487 11391 15493
rect 11333 15453 11345 15487
rect 11379 15453 11391 15487
rect 11333 15447 11391 15453
rect 11425 15487 11483 15493
rect 11425 15453 11437 15487
rect 11471 15453 11483 15487
rect 11425 15447 11483 15453
rect 11701 15487 11759 15493
rect 11701 15453 11713 15487
rect 11747 15484 11759 15487
rect 11790 15484 11796 15496
rect 11747 15456 11796 15484
rect 11747 15453 11759 15456
rect 11701 15447 11759 15453
rect 10980 15416 11008 15444
rect 9646 15388 9812 15416
rect 9784 15360 9812 15388
rect 10704 15388 11008 15416
rect 3142 15308 3148 15360
rect 3200 15348 3206 15360
rect 3421 15351 3479 15357
rect 3421 15348 3433 15351
rect 3200 15320 3433 15348
rect 3200 15308 3206 15320
rect 3421 15317 3433 15320
rect 3467 15317 3479 15351
rect 3421 15311 3479 15317
rect 3605 15351 3663 15357
rect 3605 15317 3617 15351
rect 3651 15348 3663 15351
rect 3878 15348 3884 15360
rect 3651 15320 3884 15348
rect 3651 15317 3663 15320
rect 3605 15311 3663 15317
rect 3878 15308 3884 15320
rect 3936 15308 3942 15360
rect 3970 15308 3976 15360
rect 4028 15348 4034 15360
rect 4433 15351 4491 15357
rect 4433 15348 4445 15351
rect 4028 15320 4445 15348
rect 4028 15308 4034 15320
rect 4433 15317 4445 15320
rect 4479 15317 4491 15351
rect 4433 15311 4491 15317
rect 5169 15351 5227 15357
rect 5169 15317 5181 15351
rect 5215 15348 5227 15351
rect 6362 15348 6368 15360
rect 5215 15320 6368 15348
rect 5215 15317 5227 15320
rect 5169 15311 5227 15317
rect 6362 15308 6368 15320
rect 6420 15308 6426 15360
rect 6546 15308 6552 15360
rect 6604 15308 6610 15360
rect 8294 15308 8300 15360
rect 8352 15308 8358 15360
rect 9306 15308 9312 15360
rect 9364 15308 9370 15360
rect 9766 15308 9772 15360
rect 9824 15308 9830 15360
rect 10318 15308 10324 15360
rect 10376 15348 10382 15360
rect 10704 15348 10732 15388
rect 10376 15320 10732 15348
rect 10873 15351 10931 15357
rect 10376 15308 10382 15320
rect 10873 15317 10885 15351
rect 10919 15348 10931 15351
rect 10962 15348 10968 15360
rect 10919 15320 10968 15348
rect 10919 15317 10931 15320
rect 10873 15311 10931 15317
rect 10962 15308 10968 15320
rect 11020 15308 11026 15360
rect 11330 15308 11336 15360
rect 11388 15348 11394 15360
rect 11440 15348 11468 15447
rect 11790 15444 11796 15456
rect 11848 15444 11854 15496
rect 11977 15487 12035 15493
rect 11977 15453 11989 15487
rect 12023 15484 12035 15487
rect 12084 15484 12112 15660
rect 12989 15657 13001 15660
rect 13035 15657 13047 15691
rect 12989 15651 13047 15657
rect 13449 15691 13507 15697
rect 13449 15657 13461 15691
rect 13495 15688 13507 15691
rect 13998 15688 14004 15700
rect 13495 15660 14004 15688
rect 13495 15657 13507 15660
rect 13449 15651 13507 15657
rect 13998 15648 14004 15660
rect 14056 15688 14062 15700
rect 14277 15691 14335 15697
rect 14277 15688 14289 15691
rect 14056 15660 14289 15688
rect 14056 15648 14062 15660
rect 14277 15657 14289 15660
rect 14323 15657 14335 15691
rect 14277 15651 14335 15657
rect 14461 15691 14519 15697
rect 14461 15657 14473 15691
rect 14507 15688 14519 15691
rect 14642 15688 14648 15700
rect 14507 15660 14648 15688
rect 14507 15657 14519 15660
rect 14461 15651 14519 15657
rect 14642 15648 14648 15660
rect 14700 15648 14706 15700
rect 14737 15691 14795 15697
rect 14737 15657 14749 15691
rect 14783 15688 14795 15691
rect 14826 15688 14832 15700
rect 14783 15660 14832 15688
rect 14783 15657 14795 15660
rect 14737 15651 14795 15657
rect 14826 15648 14832 15660
rect 14884 15648 14890 15700
rect 13722 15580 13728 15632
rect 13780 15620 13786 15632
rect 15105 15623 15163 15629
rect 15105 15620 15117 15623
rect 13780 15592 15117 15620
rect 13780 15580 13786 15592
rect 15105 15589 15117 15592
rect 15151 15589 15163 15623
rect 15105 15583 15163 15589
rect 15749 15623 15807 15629
rect 15749 15589 15761 15623
rect 15795 15589 15807 15623
rect 15749 15583 15807 15589
rect 15010 15512 15016 15564
rect 15068 15552 15074 15564
rect 15068 15524 15424 15552
rect 15068 15512 15074 15524
rect 12023 15456 12112 15484
rect 12023 15453 12035 15456
rect 11977 15447 12035 15453
rect 12342 15444 12348 15496
rect 12400 15444 12406 15496
rect 12526 15444 12532 15496
rect 12584 15484 12590 15496
rect 12621 15487 12679 15493
rect 12621 15484 12633 15487
rect 12584 15456 12633 15484
rect 12584 15444 12590 15456
rect 12621 15453 12633 15456
rect 12667 15453 12679 15487
rect 12621 15447 12679 15453
rect 13280 15456 14136 15484
rect 13280 15428 13308 15456
rect 11606 15376 11612 15428
rect 11664 15416 11670 15428
rect 12161 15419 12219 15425
rect 12161 15416 12173 15419
rect 11664 15388 12173 15416
rect 11664 15376 11670 15388
rect 12161 15385 12173 15388
rect 12207 15385 12219 15419
rect 12161 15379 12219 15385
rect 12253 15419 12311 15425
rect 12253 15385 12265 15419
rect 12299 15416 12311 15419
rect 12805 15419 12863 15425
rect 12299 15388 12664 15416
rect 12299 15385 12311 15388
rect 12253 15379 12311 15385
rect 12636 15360 12664 15388
rect 12805 15385 12817 15419
rect 12851 15416 12863 15419
rect 12894 15416 12900 15428
rect 12851 15388 12900 15416
rect 12851 15385 12863 15388
rect 12805 15379 12863 15385
rect 12894 15376 12900 15388
rect 12952 15376 12958 15428
rect 13262 15376 13268 15428
rect 13320 15376 13326 15428
rect 13354 15376 13360 15428
rect 13412 15416 13418 15428
rect 14108 15425 14136 15456
rect 14182 15444 14188 15496
rect 14240 15484 14246 15496
rect 14645 15487 14703 15493
rect 14645 15484 14657 15487
rect 14240 15456 14657 15484
rect 14240 15444 14246 15456
rect 14645 15453 14657 15456
rect 14691 15453 14703 15487
rect 14645 15447 14703 15453
rect 14918 15444 14924 15496
rect 14976 15444 14982 15496
rect 15286 15444 15292 15496
rect 15344 15444 15350 15496
rect 15396 15493 15424 15524
rect 15381 15487 15439 15493
rect 15381 15453 15393 15487
rect 15427 15453 15439 15487
rect 15381 15447 15439 15453
rect 15562 15444 15568 15496
rect 15620 15444 15626 15496
rect 15657 15487 15715 15493
rect 15657 15453 15669 15487
rect 15703 15484 15715 15487
rect 15764 15484 15792 15583
rect 15703 15456 15792 15484
rect 15933 15487 15991 15493
rect 15703 15453 15715 15456
rect 15657 15447 15715 15453
rect 15933 15453 15945 15487
rect 15979 15453 15991 15487
rect 15933 15447 15991 15453
rect 13449 15419 13507 15425
rect 13449 15416 13461 15419
rect 13412 15388 13461 15416
rect 13412 15376 13418 15388
rect 13449 15385 13461 15388
rect 13495 15385 13507 15419
rect 13449 15379 13507 15385
rect 14093 15419 14151 15425
rect 14093 15385 14105 15419
rect 14139 15385 14151 15419
rect 15948 15416 15976 15447
rect 16022 15444 16028 15496
rect 16080 15444 16086 15496
rect 16114 15444 16120 15496
rect 16172 15444 16178 15496
rect 16301 15487 16359 15493
rect 16301 15453 16313 15487
rect 16347 15484 16359 15487
rect 16390 15484 16396 15496
rect 16347 15456 16396 15484
rect 16347 15453 16359 15456
rect 16301 15447 16359 15453
rect 16390 15444 16396 15456
rect 16448 15444 16454 15496
rect 14093 15379 14151 15385
rect 14660 15388 15976 15416
rect 14660 15360 14688 15388
rect 11514 15348 11520 15360
rect 11388 15320 11520 15348
rect 11388 15308 11394 15320
rect 11514 15308 11520 15320
rect 11572 15308 11578 15360
rect 11885 15351 11943 15357
rect 11885 15317 11897 15351
rect 11931 15348 11943 15351
rect 12066 15348 12072 15360
rect 11931 15320 12072 15348
rect 11931 15317 11943 15320
rect 11885 15311 11943 15317
rect 12066 15308 12072 15320
rect 12124 15308 12130 15360
rect 12526 15308 12532 15360
rect 12584 15308 12590 15360
rect 12618 15308 12624 15360
rect 12676 15308 12682 15360
rect 12986 15308 12992 15360
rect 13044 15348 13050 15360
rect 13633 15351 13691 15357
rect 13633 15348 13645 15351
rect 13044 15320 13645 15348
rect 13044 15308 13050 15320
rect 13633 15317 13645 15320
rect 13679 15317 13691 15351
rect 13633 15311 13691 15317
rect 13814 15308 13820 15360
rect 13872 15348 13878 15360
rect 14277 15351 14335 15357
rect 14277 15348 14289 15351
rect 13872 15320 14289 15348
rect 13872 15308 13878 15320
rect 14277 15317 14289 15320
rect 14323 15348 14335 15351
rect 14366 15348 14372 15360
rect 14323 15320 14372 15348
rect 14323 15317 14335 15320
rect 14277 15311 14335 15317
rect 14366 15308 14372 15320
rect 14424 15308 14430 15360
rect 14642 15308 14648 15360
rect 14700 15308 14706 15360
rect 1104 15258 16652 15280
rect 1104 15206 4874 15258
rect 4926 15206 4938 15258
rect 4990 15206 5002 15258
rect 5054 15206 5066 15258
rect 5118 15206 5130 15258
rect 5182 15206 16652 15258
rect 1104 15184 16652 15206
rect 1578 15104 1584 15156
rect 1636 15144 1642 15156
rect 2041 15147 2099 15153
rect 2041 15144 2053 15147
rect 1636 15116 2053 15144
rect 1636 15104 1642 15116
rect 2041 15113 2053 15116
rect 2087 15113 2099 15147
rect 2041 15107 2099 15113
rect 2406 15104 2412 15156
rect 2464 15144 2470 15156
rect 2593 15147 2651 15153
rect 2593 15144 2605 15147
rect 2464 15116 2605 15144
rect 2464 15104 2470 15116
rect 2593 15113 2605 15116
rect 2639 15113 2651 15147
rect 2593 15107 2651 15113
rect 3694 15104 3700 15156
rect 3752 15144 3758 15156
rect 4890 15144 4896 15156
rect 3752 15116 4896 15144
rect 3752 15104 3758 15116
rect 4890 15104 4896 15116
rect 4948 15104 4954 15156
rect 5718 15104 5724 15156
rect 5776 15104 5782 15156
rect 6178 15104 6184 15156
rect 6236 15104 6242 15156
rect 6914 15144 6920 15156
rect 6380 15116 6920 15144
rect 5077 15079 5135 15085
rect 5077 15045 5089 15079
rect 5123 15076 5135 15079
rect 5442 15076 5448 15088
rect 5123 15048 5448 15076
rect 5123 15045 5135 15048
rect 5077 15039 5135 15045
rect 5442 15036 5448 15048
rect 5500 15036 5506 15088
rect 5813 15079 5871 15085
rect 5813 15045 5825 15079
rect 5859 15076 5871 15079
rect 6380 15076 6408 15116
rect 6914 15104 6920 15116
rect 6972 15104 6978 15156
rect 7837 15147 7895 15153
rect 7837 15113 7849 15147
rect 7883 15144 7895 15147
rect 8294 15144 8300 15156
rect 7883 15116 8300 15144
rect 7883 15113 7895 15116
rect 7837 15107 7895 15113
rect 8294 15104 8300 15116
rect 8352 15104 8358 15156
rect 9585 15147 9643 15153
rect 9585 15113 9597 15147
rect 9631 15144 9643 15147
rect 9858 15144 9864 15156
rect 9631 15116 9864 15144
rect 9631 15113 9643 15116
rect 9585 15107 9643 15113
rect 9858 15104 9864 15116
rect 9916 15104 9922 15156
rect 10597 15147 10655 15153
rect 10597 15144 10609 15147
rect 9968 15116 10609 15144
rect 5859 15048 6408 15076
rect 6472 15048 8156 15076
rect 5859 15045 5871 15048
rect 5813 15039 5871 15045
rect 1949 15011 2007 15017
rect 1949 14977 1961 15011
rect 1995 15008 2007 15011
rect 2038 15008 2044 15020
rect 1995 14980 2044 15008
rect 1995 14977 2007 14980
rect 1949 14971 2007 14977
rect 2038 14968 2044 14980
rect 2096 14968 2102 15020
rect 2130 14968 2136 15020
rect 2188 14968 2194 15020
rect 2498 14968 2504 15020
rect 2556 14968 2562 15020
rect 2685 15011 2743 15017
rect 2685 14977 2697 15011
rect 2731 15008 2743 15011
rect 4706 15008 4712 15020
rect 2731 14980 4712 15008
rect 2731 14977 2743 14980
rect 2685 14971 2743 14977
rect 4706 14968 4712 14980
rect 4764 14968 4770 15020
rect 5166 14968 5172 15020
rect 5224 15008 5230 15020
rect 5261 15011 5319 15017
rect 5261 15008 5273 15011
rect 5224 14980 5273 15008
rect 5224 14968 5230 14980
rect 5261 14977 5273 14980
rect 5307 14977 5319 15011
rect 5261 14971 5319 14977
rect 5534 14968 5540 15020
rect 5592 14968 5598 15020
rect 5353 14943 5411 14949
rect 5353 14909 5365 14943
rect 5399 14940 5411 14943
rect 5828 14940 5856 15039
rect 5994 14968 6000 15020
rect 6052 14968 6058 15020
rect 6472 15017 6500 15048
rect 8128 15020 8156 15048
rect 8938 15036 8944 15088
rect 8996 15076 9002 15088
rect 9968 15085 9996 15116
rect 10597 15113 10609 15116
rect 10643 15144 10655 15147
rect 10686 15144 10692 15156
rect 10643 15116 10692 15144
rect 10643 15113 10655 15116
rect 10597 15107 10655 15113
rect 10686 15104 10692 15116
rect 10744 15104 10750 15156
rect 10778 15104 10784 15156
rect 10836 15104 10842 15156
rect 10870 15104 10876 15156
rect 10928 15104 10934 15156
rect 11054 15104 11060 15156
rect 11112 15144 11118 15156
rect 11790 15144 11796 15156
rect 11112 15116 11796 15144
rect 11112 15104 11118 15116
rect 11790 15104 11796 15116
rect 11848 15104 11854 15156
rect 12069 15147 12127 15153
rect 12069 15113 12081 15147
rect 12115 15144 12127 15147
rect 12621 15147 12679 15153
rect 12621 15144 12633 15147
rect 12115 15116 12633 15144
rect 12115 15113 12127 15116
rect 12069 15107 12127 15113
rect 12621 15113 12633 15116
rect 12667 15113 12679 15147
rect 12621 15107 12679 15113
rect 14185 15147 14243 15153
rect 14185 15113 14197 15147
rect 14231 15144 14243 15147
rect 14231 15116 16252 15144
rect 14231 15113 14243 15116
rect 14185 15107 14243 15113
rect 9953 15079 10011 15085
rect 8996 15048 9904 15076
rect 8996 15036 9002 15048
rect 6457 15011 6515 15017
rect 6457 14977 6469 15011
rect 6503 14977 6515 15011
rect 6713 15011 6771 15017
rect 6713 15008 6725 15011
rect 6457 14971 6515 14977
rect 6564 14980 6725 15008
rect 5399 14912 5856 14940
rect 5399 14909 5411 14912
rect 5353 14903 5411 14909
rect 6362 14900 6368 14952
rect 6420 14940 6426 14952
rect 6564 14940 6592 14980
rect 6713 14977 6725 14980
rect 6759 14977 6771 15011
rect 6713 14971 6771 14977
rect 8110 14968 8116 15020
rect 8168 15008 8174 15020
rect 9876 15017 9904 15048
rect 9953 15045 9965 15079
rect 9999 15045 10011 15079
rect 9953 15039 10011 15045
rect 10045 15079 10103 15085
rect 10045 15045 10057 15079
rect 10091 15076 10103 15079
rect 10502 15076 10508 15088
rect 10091 15048 10508 15076
rect 10091 15045 10103 15048
rect 10045 15039 10103 15045
rect 10502 15036 10508 15048
rect 10560 15076 10566 15088
rect 10796 15076 10824 15104
rect 10560 15048 10824 15076
rect 10888 15076 10916 15104
rect 16224 15088 16252 15116
rect 10888 15048 11192 15076
rect 10560 15036 10566 15048
rect 8205 15011 8263 15017
rect 8205 15008 8217 15011
rect 8168 14980 8217 15008
rect 8168 14968 8174 14980
rect 8205 14977 8217 14980
rect 8251 14977 8263 15011
rect 8205 14971 8263 14977
rect 8472 15011 8530 15017
rect 8472 14977 8484 15011
rect 8518 15008 8530 15011
rect 9677 15011 9735 15017
rect 9677 15008 9689 15011
rect 8518 14980 9689 15008
rect 8518 14977 8530 14980
rect 8472 14971 8530 14977
rect 9677 14977 9689 14980
rect 9723 14977 9735 15011
rect 9677 14971 9735 14977
rect 9861 15011 9919 15017
rect 9861 14977 9873 15011
rect 9907 14977 9919 15011
rect 10163 15011 10221 15017
rect 10163 15008 10175 15011
rect 9861 14971 9919 14977
rect 10152 14977 10175 15008
rect 10209 14977 10221 15011
rect 10152 14971 10221 14977
rect 10413 15011 10471 15017
rect 10413 14977 10425 15011
rect 10459 14977 10471 15011
rect 10413 14971 10471 14977
rect 6420 14912 6592 14940
rect 6420 14900 6426 14912
rect 9214 14900 9220 14952
rect 9272 14940 9278 14952
rect 10152 14940 10180 14971
rect 9272 14912 10180 14940
rect 10321 14943 10379 14949
rect 9272 14900 9278 14912
rect 10321 14909 10333 14943
rect 10367 14940 10379 14943
rect 10428 14940 10456 14971
rect 10594 14968 10600 15020
rect 10652 14968 10658 15020
rect 10689 15011 10747 15017
rect 10689 14977 10701 15011
rect 10735 15008 10747 15011
rect 10778 15008 10784 15020
rect 10735 14980 10784 15008
rect 10735 14977 10747 14980
rect 10689 14971 10747 14977
rect 10778 14968 10784 14980
rect 10836 14968 10842 15020
rect 10873 15011 10931 15017
rect 10873 14977 10885 15011
rect 10919 14977 10931 15011
rect 10873 14971 10931 14977
rect 10965 15011 11023 15017
rect 10965 14977 10977 15011
rect 11011 14977 11023 15011
rect 10965 14971 11023 14977
rect 10888 14940 10916 14971
rect 10367 14912 10456 14940
rect 10520 14912 10916 14940
rect 10367 14909 10379 14912
rect 10321 14903 10379 14909
rect 9858 14832 9864 14884
rect 9916 14872 9922 14884
rect 10134 14872 10140 14884
rect 9916 14844 10140 14872
rect 9916 14832 9922 14844
rect 10134 14832 10140 14844
rect 10192 14872 10198 14884
rect 10336 14872 10364 14903
rect 10192 14844 10364 14872
rect 10192 14832 10198 14844
rect 10410 14832 10416 14884
rect 10468 14872 10474 14884
rect 10520 14872 10548 14912
rect 10468 14844 10548 14872
rect 10468 14832 10474 14844
rect 10870 14832 10876 14884
rect 10928 14872 10934 14884
rect 10980 14872 11008 14971
rect 11054 14968 11060 15020
rect 11112 14968 11118 15020
rect 11164 15008 11192 15048
rect 11422 15036 11428 15088
rect 11480 15076 11486 15088
rect 11480 15048 14504 15076
rect 11480 15036 11486 15048
rect 14476 15020 14504 15048
rect 14752 15048 15516 15076
rect 14752 15020 14780 15048
rect 11517 15011 11575 15017
rect 11517 15008 11529 15011
rect 11164 14980 11529 15008
rect 11517 14977 11529 14980
rect 11563 14977 11575 15011
rect 11517 14971 11575 14977
rect 11698 14968 11704 15020
rect 11756 14968 11762 15020
rect 11790 14968 11796 15020
rect 11848 14968 11854 15020
rect 11885 15011 11943 15017
rect 11885 14977 11897 15011
rect 11931 15008 11943 15011
rect 12342 15008 12348 15020
rect 11931 14980 12348 15008
rect 11931 14977 11943 14980
rect 11885 14971 11943 14977
rect 11606 14900 11612 14952
rect 11664 14940 11670 14952
rect 11900 14940 11928 14971
rect 12342 14968 12348 14980
rect 12400 14968 12406 15020
rect 12529 15011 12587 15017
rect 12529 14977 12541 15011
rect 12575 15008 12587 15011
rect 12989 15011 13047 15017
rect 12989 15008 13001 15011
rect 12575 14980 13001 15008
rect 12575 14977 12587 14980
rect 12529 14971 12587 14977
rect 12989 14977 13001 14980
rect 13035 14977 13047 15011
rect 12989 14971 13047 14977
rect 14001 15011 14059 15017
rect 14001 14977 14013 15011
rect 14047 15008 14059 15011
rect 14090 15008 14096 15020
rect 14047 14980 14096 15008
rect 14047 14977 14059 14980
rect 14001 14971 14059 14977
rect 14090 14968 14096 14980
rect 14148 14968 14154 15020
rect 14458 14968 14464 15020
rect 14516 15008 14522 15020
rect 14645 15011 14703 15017
rect 14645 15008 14657 15011
rect 14516 14980 14657 15008
rect 14516 14968 14522 14980
rect 14645 14977 14657 14980
rect 14691 14977 14703 15011
rect 14645 14971 14703 14977
rect 11664 14912 11928 14940
rect 11664 14900 11670 14912
rect 12066 14900 12072 14952
rect 12124 14940 12130 14952
rect 12713 14943 12771 14949
rect 12124 14912 12572 14940
rect 12124 14900 12130 14912
rect 10928 14844 11008 14872
rect 11333 14875 11391 14881
rect 10928 14832 10934 14844
rect 11333 14841 11345 14875
rect 11379 14872 11391 14875
rect 12434 14872 12440 14884
rect 11379 14844 12440 14872
rect 11379 14841 11391 14844
rect 11333 14835 11391 14841
rect 12434 14832 12440 14844
rect 12492 14832 12498 14884
rect 12544 14872 12572 14912
rect 12713 14909 12725 14943
rect 12759 14909 12771 14943
rect 12713 14903 12771 14909
rect 12728 14872 12756 14903
rect 13262 14900 13268 14952
rect 13320 14940 13326 14952
rect 13541 14943 13599 14949
rect 13541 14940 13553 14943
rect 13320 14912 13553 14940
rect 13320 14900 13326 14912
rect 13541 14909 13553 14912
rect 13587 14909 13599 14943
rect 13541 14903 13599 14909
rect 13814 14900 13820 14952
rect 13872 14900 13878 14952
rect 12544 14844 12756 14872
rect 14660 14872 14688 14971
rect 14734 14968 14740 15020
rect 14792 14968 14798 15020
rect 14829 15011 14887 15017
rect 14829 14977 14841 15011
rect 14875 14977 14887 15011
rect 14829 14971 14887 14977
rect 14844 14940 14872 14971
rect 15010 14968 15016 15020
rect 15068 14968 15074 15020
rect 15378 14968 15384 15020
rect 15436 14968 15442 15020
rect 15488 15017 15516 15048
rect 16206 15036 16212 15088
rect 16264 15036 16270 15088
rect 15473 15011 15531 15017
rect 15473 14977 15485 15011
rect 15519 14977 15531 15011
rect 15473 14971 15531 14977
rect 15565 15011 15623 15017
rect 15565 14977 15577 15011
rect 15611 15008 15623 15011
rect 15654 15008 15660 15020
rect 15611 14980 15660 15008
rect 15611 14977 15623 14980
rect 15565 14971 15623 14977
rect 15654 14968 15660 14980
rect 15712 14968 15718 15020
rect 15749 15011 15807 15017
rect 15749 14977 15761 15011
rect 15795 15008 15807 15011
rect 15930 15008 15936 15020
rect 15795 14980 15936 15008
rect 15795 14977 15807 14980
rect 15749 14971 15807 14977
rect 15930 14968 15936 14980
rect 15988 14968 15994 15020
rect 16022 14968 16028 15020
rect 16080 14968 16086 15020
rect 15841 14943 15899 14949
rect 15841 14940 15853 14943
rect 14844 14912 15853 14940
rect 15841 14909 15853 14912
rect 15887 14909 15899 14943
rect 15841 14903 15899 14909
rect 14826 14872 14832 14884
rect 14660 14844 14832 14872
rect 14826 14832 14832 14844
rect 14884 14832 14890 14884
rect 15010 14832 15016 14884
rect 15068 14872 15074 14884
rect 15930 14872 15936 14884
rect 15068 14844 15936 14872
rect 15068 14832 15074 14844
rect 15930 14832 15936 14844
rect 15988 14832 15994 14884
rect 4706 14764 4712 14816
rect 4764 14804 4770 14816
rect 4893 14807 4951 14813
rect 4893 14804 4905 14807
rect 4764 14776 4905 14804
rect 4764 14764 4770 14776
rect 4893 14773 4905 14776
rect 4939 14773 4951 14807
rect 4893 14767 4951 14773
rect 9490 14764 9496 14816
rect 9548 14804 9554 14816
rect 10594 14804 10600 14816
rect 9548 14776 10600 14804
rect 9548 14764 9554 14776
rect 10594 14764 10600 14776
rect 10652 14764 10658 14816
rect 12158 14764 12164 14816
rect 12216 14764 12222 14816
rect 12342 14764 12348 14816
rect 12400 14804 12406 14816
rect 13722 14804 13728 14816
rect 12400 14776 13728 14804
rect 12400 14764 12406 14776
rect 13722 14764 13728 14776
rect 13780 14764 13786 14816
rect 14369 14807 14427 14813
rect 14369 14773 14381 14807
rect 14415 14804 14427 14807
rect 14734 14804 14740 14816
rect 14415 14776 14740 14804
rect 14415 14773 14427 14776
rect 14369 14767 14427 14773
rect 14734 14764 14740 14776
rect 14792 14764 14798 14816
rect 15102 14764 15108 14816
rect 15160 14764 15166 14816
rect 1104 14714 16652 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 16652 14714
rect 1104 14640 16652 14662
rect 5626 14560 5632 14612
rect 5684 14560 5690 14612
rect 10413 14603 10471 14609
rect 10413 14569 10425 14603
rect 10459 14600 10471 14603
rect 10502 14600 10508 14612
rect 10459 14572 10508 14600
rect 10459 14569 10471 14572
rect 10413 14563 10471 14569
rect 10502 14560 10508 14572
rect 10560 14560 10566 14612
rect 10689 14603 10747 14609
rect 10689 14569 10701 14603
rect 10735 14569 10747 14603
rect 10689 14563 10747 14569
rect 6270 14492 6276 14544
rect 6328 14492 6334 14544
rect 8754 14492 8760 14544
rect 8812 14492 8818 14544
rect 9030 14492 9036 14544
rect 9088 14532 9094 14544
rect 9490 14532 9496 14544
rect 9088 14504 9496 14532
rect 9088 14492 9094 14504
rect 9490 14492 9496 14504
rect 9548 14532 9554 14544
rect 9548 14504 9628 14532
rect 9548 14492 9554 14504
rect 4062 14424 4068 14476
rect 4120 14464 4126 14476
rect 4249 14467 4307 14473
rect 4249 14464 4261 14467
rect 4120 14436 4261 14464
rect 4120 14424 4126 14436
rect 4249 14433 4261 14436
rect 4295 14433 4307 14467
rect 4249 14427 4307 14433
rect 4890 14424 4896 14476
rect 4948 14464 4954 14476
rect 5721 14467 5779 14473
rect 5721 14464 5733 14467
rect 4948 14436 5733 14464
rect 4948 14424 4954 14436
rect 5721 14433 5733 14436
rect 5767 14464 5779 14467
rect 6288 14464 6316 14492
rect 6914 14464 6920 14476
rect 5767 14436 6316 14464
rect 6472 14436 6920 14464
rect 5767 14433 5779 14436
rect 5721 14427 5779 14433
rect 3326 14356 3332 14408
rect 3384 14356 3390 14408
rect 4338 14356 4344 14408
rect 4396 14396 4402 14408
rect 4433 14399 4491 14405
rect 4433 14396 4445 14399
rect 4396 14368 4445 14396
rect 4396 14356 4402 14368
rect 4433 14365 4445 14368
rect 4479 14365 4491 14399
rect 4433 14359 4491 14365
rect 4525 14399 4583 14405
rect 4525 14365 4537 14399
rect 4571 14396 4583 14399
rect 4614 14396 4620 14408
rect 4571 14368 4620 14396
rect 4571 14365 4583 14368
rect 4525 14359 4583 14365
rect 4614 14356 4620 14368
rect 4672 14356 4678 14408
rect 5077 14399 5135 14405
rect 5077 14365 5089 14399
rect 5123 14396 5135 14399
rect 5258 14396 5264 14408
rect 5123 14368 5264 14396
rect 5123 14365 5135 14368
rect 5077 14359 5135 14365
rect 5258 14356 5264 14368
rect 5316 14356 5322 14408
rect 5442 14356 5448 14408
rect 5500 14356 5506 14408
rect 5997 14399 6055 14405
rect 5997 14365 6009 14399
rect 6043 14396 6055 14399
rect 6086 14396 6092 14408
rect 6043 14368 6092 14396
rect 6043 14365 6055 14368
rect 5997 14359 6055 14365
rect 6086 14356 6092 14368
rect 6144 14356 6150 14408
rect 6178 14356 6184 14408
rect 6236 14356 6242 14408
rect 6273 14399 6331 14405
rect 6273 14365 6285 14399
rect 6319 14396 6331 14399
rect 6362 14396 6368 14408
rect 6319 14368 6368 14396
rect 6319 14365 6331 14368
rect 6273 14359 6331 14365
rect 6362 14356 6368 14368
rect 6420 14356 6426 14408
rect 6472 14405 6500 14436
rect 6914 14424 6920 14436
rect 6972 14464 6978 14476
rect 7190 14464 7196 14476
rect 6972 14436 7196 14464
rect 6972 14424 6978 14436
rect 7190 14424 7196 14436
rect 7248 14424 7254 14476
rect 9214 14424 9220 14476
rect 9272 14464 9278 14476
rect 9600 14473 9628 14504
rect 9674 14492 9680 14544
rect 9732 14532 9738 14544
rect 10045 14535 10103 14541
rect 10045 14532 10057 14535
rect 9732 14504 10057 14532
rect 9732 14492 9738 14504
rect 10045 14501 10057 14504
rect 10091 14501 10103 14535
rect 10045 14495 10103 14501
rect 10594 14492 10600 14544
rect 10652 14492 10658 14544
rect 10704 14532 10732 14563
rect 10778 14560 10784 14612
rect 10836 14600 10842 14612
rect 11057 14603 11115 14609
rect 11057 14600 11069 14603
rect 10836 14572 11069 14600
rect 10836 14560 10842 14572
rect 11057 14569 11069 14572
rect 11103 14569 11115 14603
rect 13633 14603 13691 14609
rect 13633 14600 13645 14603
rect 11057 14563 11115 14569
rect 11164 14572 13645 14600
rect 10704 14504 11100 14532
rect 11072 14476 11100 14504
rect 9401 14467 9459 14473
rect 9401 14464 9413 14467
rect 9272 14436 9413 14464
rect 9272 14424 9278 14436
rect 9401 14433 9413 14436
rect 9447 14433 9459 14467
rect 9401 14427 9459 14433
rect 9585 14467 9643 14473
rect 9585 14433 9597 14467
rect 9631 14433 9643 14467
rect 9585 14427 9643 14433
rect 9950 14424 9956 14476
rect 10008 14464 10014 14476
rect 10781 14467 10839 14473
rect 10781 14464 10793 14467
rect 10008 14436 10793 14464
rect 10008 14424 10014 14436
rect 10781 14433 10793 14436
rect 10827 14433 10839 14467
rect 10781 14427 10839 14433
rect 11054 14424 11060 14476
rect 11112 14424 11118 14476
rect 6457 14399 6515 14405
rect 6457 14365 6469 14399
rect 6503 14365 6515 14399
rect 6457 14359 6515 14365
rect 6733 14399 6791 14405
rect 6733 14365 6745 14399
rect 6779 14365 6791 14399
rect 6733 14359 6791 14365
rect 7837 14399 7895 14405
rect 7837 14365 7849 14399
rect 7883 14396 7895 14399
rect 8018 14396 8024 14408
rect 7883 14368 8024 14396
rect 7883 14365 7895 14368
rect 7837 14359 7895 14365
rect 4798 14288 4804 14340
rect 4856 14328 4862 14340
rect 6748 14328 6776 14359
rect 8018 14356 8024 14368
rect 8076 14356 8082 14408
rect 8113 14399 8171 14405
rect 8113 14365 8125 14399
rect 8159 14365 8171 14399
rect 8113 14359 8171 14365
rect 7282 14328 7288 14340
rect 4856 14300 7288 14328
rect 4856 14288 4862 14300
rect 7282 14288 7288 14300
rect 7340 14288 7346 14340
rect 8128 14328 8156 14359
rect 8294 14356 8300 14408
rect 8352 14356 8358 14408
rect 8570 14356 8576 14408
rect 8628 14356 8634 14408
rect 8938 14356 8944 14408
rect 8996 14396 9002 14408
rect 11164 14405 11192 14572
rect 13633 14569 13645 14572
rect 13679 14569 13691 14603
rect 13633 14563 13691 14569
rect 14277 14603 14335 14609
rect 14277 14569 14289 14603
rect 14323 14600 14335 14603
rect 15194 14600 15200 14612
rect 14323 14572 15200 14600
rect 14323 14569 14335 14572
rect 14277 14563 14335 14569
rect 15194 14560 15200 14572
rect 15252 14600 15258 14612
rect 15252 14572 15424 14600
rect 15252 14560 15258 14572
rect 11330 14532 11336 14544
rect 11256 14504 11336 14532
rect 9309 14399 9367 14405
rect 9309 14396 9321 14399
rect 8996 14368 9321 14396
rect 8996 14356 9002 14368
rect 9309 14365 9321 14368
rect 9355 14365 9367 14399
rect 9309 14359 9367 14365
rect 10689 14399 10747 14405
rect 10689 14365 10701 14399
rect 10735 14365 10747 14399
rect 10689 14359 10747 14365
rect 11149 14399 11207 14405
rect 11149 14365 11161 14399
rect 11195 14365 11207 14399
rect 11149 14359 11207 14365
rect 8386 14328 8392 14340
rect 8128 14300 8392 14328
rect 8386 14288 8392 14300
rect 8444 14288 8450 14340
rect 10704 14328 10732 14359
rect 11256 14328 11284 14504
rect 11330 14492 11336 14504
rect 11388 14492 11394 14544
rect 13998 14492 14004 14544
rect 14056 14532 14062 14544
rect 14185 14535 14243 14541
rect 14185 14532 14197 14535
rect 14056 14504 14197 14532
rect 14056 14492 14062 14504
rect 14185 14501 14197 14504
rect 14231 14501 14243 14535
rect 15396 14532 15424 14572
rect 15654 14560 15660 14612
rect 15712 14600 15718 14612
rect 16301 14603 16359 14609
rect 16301 14600 16313 14603
rect 15712 14572 16313 14600
rect 15712 14560 15718 14572
rect 16301 14569 16313 14572
rect 16347 14569 16359 14603
rect 16301 14563 16359 14569
rect 16114 14532 16120 14544
rect 15396 14504 16120 14532
rect 14185 14495 14243 14501
rect 16114 14492 16120 14504
rect 16172 14492 16178 14544
rect 11698 14464 11704 14476
rect 11348 14436 11704 14464
rect 11348 14405 11376 14436
rect 11698 14424 11704 14436
rect 11756 14424 11762 14476
rect 13354 14424 13360 14476
rect 13412 14464 13418 14476
rect 13412 14436 13860 14464
rect 13412 14424 13418 14436
rect 11333 14399 11391 14405
rect 11333 14365 11345 14399
rect 11379 14365 11391 14399
rect 11333 14359 11391 14365
rect 11422 14356 11428 14408
rect 11480 14356 11486 14408
rect 11517 14399 11575 14405
rect 11517 14365 11529 14399
rect 11563 14396 11575 14399
rect 11606 14396 11612 14408
rect 11563 14368 11612 14396
rect 11563 14365 11575 14368
rect 11517 14359 11575 14365
rect 11606 14356 11612 14368
rect 11664 14356 11670 14408
rect 11793 14399 11851 14405
rect 11793 14365 11805 14399
rect 11839 14396 11851 14399
rect 11882 14396 11888 14408
rect 11839 14368 11888 14396
rect 11839 14365 11851 14368
rect 11793 14359 11851 14365
rect 11882 14356 11888 14368
rect 11940 14356 11946 14408
rect 13265 14399 13323 14405
rect 13265 14396 13277 14399
rect 11992 14368 13277 14396
rect 11992 14328 12020 14368
rect 13265 14365 13277 14368
rect 13311 14365 13323 14399
rect 13725 14399 13783 14405
rect 13725 14396 13737 14399
rect 13265 14359 13323 14365
rect 13556 14368 13737 14396
rect 10704 14300 11284 14328
rect 11624 14300 12020 14328
rect 12060 14331 12118 14337
rect 3418 14220 3424 14272
rect 3476 14220 3482 14272
rect 4246 14220 4252 14272
rect 4304 14260 4310 14272
rect 4525 14263 4583 14269
rect 4525 14260 4537 14263
rect 4304 14232 4537 14260
rect 4304 14220 4310 14232
rect 4525 14229 4537 14232
rect 4571 14229 4583 14263
rect 4525 14223 4583 14229
rect 4614 14220 4620 14272
rect 4672 14260 4678 14272
rect 5166 14260 5172 14272
rect 4672 14232 5172 14260
rect 4672 14220 4678 14232
rect 5166 14220 5172 14232
rect 5224 14220 5230 14272
rect 5261 14263 5319 14269
rect 5261 14229 5273 14263
rect 5307 14260 5319 14263
rect 5534 14260 5540 14272
rect 5307 14232 5540 14260
rect 5307 14229 5319 14232
rect 5261 14223 5319 14229
rect 5534 14220 5540 14232
rect 5592 14220 5598 14272
rect 5626 14220 5632 14272
rect 5684 14260 5690 14272
rect 5813 14263 5871 14269
rect 5813 14260 5825 14263
rect 5684 14232 5825 14260
rect 5684 14220 5690 14232
rect 5813 14229 5825 14232
rect 5859 14229 5871 14263
rect 5813 14223 5871 14229
rect 5994 14220 6000 14272
rect 6052 14260 6058 14272
rect 6549 14263 6607 14269
rect 6549 14260 6561 14263
rect 6052 14232 6561 14260
rect 6052 14220 6058 14232
rect 6549 14229 6561 14232
rect 6595 14229 6607 14263
rect 6549 14223 6607 14229
rect 6914 14220 6920 14272
rect 6972 14220 6978 14272
rect 8294 14220 8300 14272
rect 8352 14260 8358 14272
rect 8941 14263 8999 14269
rect 8941 14260 8953 14263
rect 8352 14232 8953 14260
rect 8352 14220 8358 14232
rect 8941 14229 8953 14232
rect 8987 14229 8999 14263
rect 8941 14223 8999 14229
rect 10413 14263 10471 14269
rect 10413 14229 10425 14263
rect 10459 14260 10471 14263
rect 10686 14260 10692 14272
rect 10459 14232 10692 14260
rect 10459 14229 10471 14232
rect 10413 14223 10471 14229
rect 10686 14220 10692 14232
rect 10744 14220 10750 14272
rect 11054 14220 11060 14272
rect 11112 14260 11118 14272
rect 11624 14260 11652 14300
rect 12060 14297 12072 14331
rect 12106 14328 12118 14331
rect 12158 14328 12164 14340
rect 12106 14300 12164 14328
rect 12106 14297 12118 14300
rect 12060 14291 12118 14297
rect 12158 14288 12164 14300
rect 12216 14288 12222 14340
rect 12894 14288 12900 14340
rect 12952 14328 12958 14340
rect 13449 14331 13507 14337
rect 13449 14328 13461 14331
rect 12952 14300 13461 14328
rect 12952 14288 12958 14300
rect 13449 14297 13461 14300
rect 13495 14297 13507 14331
rect 13449 14291 13507 14297
rect 11112 14232 11652 14260
rect 11701 14263 11759 14269
rect 11112 14220 11118 14232
rect 11701 14229 11713 14263
rect 11747 14260 11759 14263
rect 12802 14260 12808 14272
rect 11747 14232 12808 14260
rect 11747 14229 11759 14232
rect 11701 14223 11759 14229
rect 12802 14220 12808 14232
rect 12860 14220 12866 14272
rect 13173 14263 13231 14269
rect 13173 14229 13185 14263
rect 13219 14260 13231 14263
rect 13262 14260 13268 14272
rect 13219 14232 13268 14260
rect 13219 14229 13231 14232
rect 13173 14223 13231 14229
rect 13262 14220 13268 14232
rect 13320 14220 13326 14272
rect 13354 14220 13360 14272
rect 13412 14260 13418 14272
rect 13556 14260 13584 14368
rect 13725 14365 13737 14368
rect 13771 14365 13783 14399
rect 13832 14396 13860 14436
rect 13906 14424 13912 14476
rect 13964 14464 13970 14476
rect 13964 14436 14412 14464
rect 13964 14424 13970 14436
rect 13832 14390 14044 14396
rect 14082 14393 14140 14399
rect 14082 14390 14094 14393
rect 13832 14368 14094 14390
rect 13725 14359 13783 14365
rect 14016 14362 14094 14368
rect 14082 14359 14094 14362
rect 14128 14359 14140 14393
rect 14082 14353 14140 14359
rect 14384 14337 14412 14436
rect 14461 14399 14519 14405
rect 14461 14365 14473 14399
rect 14507 14396 14519 14399
rect 14550 14396 14556 14408
rect 14507 14368 14556 14396
rect 14507 14365 14519 14368
rect 14461 14359 14519 14365
rect 14550 14356 14556 14368
rect 14608 14356 14614 14408
rect 14734 14405 14740 14408
rect 14728 14396 14740 14405
rect 14695 14368 14740 14396
rect 14728 14359 14740 14368
rect 14734 14356 14740 14359
rect 14792 14356 14798 14408
rect 15654 14356 15660 14408
rect 15712 14396 15718 14408
rect 16117 14399 16175 14405
rect 16117 14396 16129 14399
rect 15712 14368 16129 14396
rect 15712 14356 15718 14368
rect 16117 14365 16129 14368
rect 16163 14365 16175 14399
rect 16117 14359 16175 14365
rect 14369 14331 14427 14337
rect 14369 14297 14381 14331
rect 14415 14328 14427 14331
rect 15286 14328 15292 14340
rect 14415 14300 15292 14328
rect 14415 14297 14427 14300
rect 14369 14291 14427 14297
rect 15286 14288 15292 14300
rect 15344 14288 15350 14340
rect 15933 14331 15991 14337
rect 15933 14297 15945 14331
rect 15979 14328 15991 14331
rect 16206 14328 16212 14340
rect 15979 14300 16212 14328
rect 15979 14297 15991 14300
rect 15933 14291 15991 14297
rect 16206 14288 16212 14300
rect 16264 14288 16270 14340
rect 13412 14232 13584 14260
rect 13412 14220 13418 14232
rect 13814 14220 13820 14272
rect 13872 14260 13878 14272
rect 14918 14260 14924 14272
rect 13872 14232 14924 14260
rect 13872 14220 13878 14232
rect 14918 14220 14924 14232
rect 14976 14220 14982 14272
rect 15841 14263 15899 14269
rect 15841 14229 15853 14263
rect 15887 14260 15899 14263
rect 16022 14260 16028 14272
rect 15887 14232 16028 14260
rect 15887 14229 15899 14232
rect 15841 14223 15899 14229
rect 16022 14220 16028 14232
rect 16080 14220 16086 14272
rect 1104 14170 16652 14192
rect 1104 14118 4874 14170
rect 4926 14118 4938 14170
rect 4990 14118 5002 14170
rect 5054 14118 5066 14170
rect 5118 14118 5130 14170
rect 5182 14118 16652 14170
rect 1104 14096 16652 14118
rect 2866 14016 2872 14068
rect 2924 14056 2930 14068
rect 3142 14056 3148 14068
rect 2924 14028 3148 14056
rect 2924 14016 2930 14028
rect 3142 14016 3148 14028
rect 3200 14056 3206 14068
rect 4617 14059 4675 14065
rect 3200 14028 4384 14056
rect 3200 14016 3206 14028
rect 3697 13991 3755 13997
rect 3697 13957 3709 13991
rect 3743 13988 3755 13991
rect 3786 13988 3792 14000
rect 3743 13960 3792 13988
rect 3743 13957 3755 13960
rect 3697 13951 3755 13957
rect 3786 13948 3792 13960
rect 3844 13948 3850 14000
rect 3927 13957 3985 13963
rect 3927 13954 3939 13957
rect 1857 13923 1915 13929
rect 1857 13889 1869 13923
rect 1903 13889 1915 13923
rect 1857 13883 1915 13889
rect 1872 13852 1900 13883
rect 2038 13880 2044 13932
rect 2096 13880 2102 13932
rect 3421 13923 3479 13929
rect 3421 13889 3433 13923
rect 3467 13889 3479 13923
rect 3421 13883 3479 13889
rect 2406 13852 2412 13864
rect 1872 13824 2412 13852
rect 2406 13812 2412 13824
rect 2464 13812 2470 13864
rect 3436 13852 3464 13883
rect 3602 13880 3608 13932
rect 3660 13880 3666 13932
rect 3922 13923 3939 13954
rect 3973 13923 3985 13957
rect 3922 13920 3985 13923
rect 4246 13920 4252 13932
rect 3922 13892 4252 13920
rect 4246 13880 4252 13892
rect 4304 13880 4310 13932
rect 4356 13929 4384 14028
rect 4617 14025 4629 14059
rect 4663 14056 4675 14059
rect 5166 14056 5172 14068
rect 4663 14028 5172 14056
rect 4663 14025 4675 14028
rect 4617 14019 4675 14025
rect 5166 14016 5172 14028
rect 5224 14056 5230 14068
rect 5442 14056 5448 14068
rect 5224 14028 5448 14056
rect 5224 14016 5230 14028
rect 5442 14016 5448 14028
rect 5500 14016 5506 14068
rect 6917 14059 6975 14065
rect 6917 14025 6929 14059
rect 6963 14056 6975 14059
rect 7098 14056 7104 14068
rect 6963 14028 7104 14056
rect 6963 14025 6975 14028
rect 6917 14019 6975 14025
rect 7098 14016 7104 14028
rect 7156 14016 7162 14068
rect 9122 14016 9128 14068
rect 9180 14056 9186 14068
rect 9401 14059 9459 14065
rect 9401 14056 9413 14059
rect 9180 14028 9413 14056
rect 9180 14016 9186 14028
rect 9401 14025 9413 14028
rect 9447 14025 9459 14059
rect 9401 14019 9459 14025
rect 9769 14059 9827 14065
rect 9769 14025 9781 14059
rect 9815 14056 9827 14059
rect 10502 14056 10508 14068
rect 9815 14028 10508 14056
rect 9815 14025 9827 14028
rect 9769 14019 9827 14025
rect 10502 14016 10508 14028
rect 10560 14016 10566 14068
rect 10781 14059 10839 14065
rect 10781 14025 10793 14059
rect 10827 14056 10839 14059
rect 11054 14056 11060 14068
rect 10827 14028 11060 14056
rect 10827 14025 10839 14028
rect 10781 14019 10839 14025
rect 11054 14016 11060 14028
rect 11112 14016 11118 14068
rect 12802 14016 12808 14068
rect 12860 14016 12866 14068
rect 14182 14016 14188 14068
rect 14240 14016 14246 14068
rect 14461 14059 14519 14065
rect 14461 14025 14473 14059
rect 14507 14056 14519 14059
rect 15194 14056 15200 14068
rect 14507 14028 15200 14056
rect 14507 14025 14519 14028
rect 14461 14019 14519 14025
rect 15194 14016 15200 14028
rect 15252 14016 15258 14068
rect 16206 14016 16212 14068
rect 16264 14016 16270 14068
rect 4540 13960 5856 13988
rect 4341 13923 4399 13929
rect 4341 13889 4353 13923
rect 4387 13920 4399 13923
rect 4430 13920 4436 13932
rect 4387 13892 4436 13920
rect 4387 13889 4399 13892
rect 4341 13883 4399 13889
rect 4430 13880 4436 13892
rect 4488 13880 4494 13932
rect 4540 13929 4568 13960
rect 4525 13923 4583 13929
rect 4525 13889 4537 13923
rect 4571 13889 4583 13923
rect 5166 13920 5172 13932
rect 4525 13883 4583 13889
rect 4724 13892 5172 13920
rect 4062 13852 4068 13864
rect 3436 13824 4068 13852
rect 4062 13812 4068 13824
rect 4120 13812 4126 13864
rect 4157 13855 4215 13861
rect 4157 13821 4169 13855
rect 4203 13852 4215 13855
rect 4724 13852 4752 13892
rect 5166 13880 5172 13892
rect 5224 13880 5230 13932
rect 5718 13880 5724 13932
rect 5776 13929 5782 13932
rect 5776 13883 5788 13929
rect 5828 13920 5856 13960
rect 6012 13960 7880 13988
rect 6012 13929 6040 13960
rect 5997 13923 6055 13929
rect 5828 13892 5948 13920
rect 5776 13880 5782 13883
rect 4203 13824 4752 13852
rect 5920 13852 5948 13892
rect 5997 13889 6009 13923
rect 6043 13889 6055 13923
rect 5997 13883 6055 13889
rect 6365 13923 6423 13929
rect 6365 13889 6377 13923
rect 6411 13920 6423 13923
rect 6822 13920 6828 13932
rect 6411 13892 6828 13920
rect 6411 13889 6423 13892
rect 6365 13883 6423 13889
rect 6822 13880 6828 13892
rect 6880 13880 6886 13932
rect 6914 13880 6920 13932
rect 6972 13880 6978 13932
rect 7006 13880 7012 13932
rect 7064 13880 7070 13932
rect 7852 13929 7880 13960
rect 8110 13948 8116 14000
rect 8168 13988 8174 14000
rect 10226 13988 10232 14000
rect 8168 13960 10232 13988
rect 8168 13948 8174 13960
rect 10226 13948 10232 13960
rect 10284 13948 10290 14000
rect 13262 13948 13268 14000
rect 13320 13988 13326 14000
rect 14820 13991 14878 13997
rect 13320 13960 14320 13988
rect 13320 13948 13326 13960
rect 7837 13923 7895 13929
rect 7837 13889 7849 13923
rect 7883 13920 7895 13923
rect 8018 13920 8024 13932
rect 7883 13892 8024 13920
rect 7883 13889 7895 13892
rect 7837 13883 7895 13889
rect 8018 13880 8024 13892
rect 8076 13880 8082 13932
rect 8294 13929 8300 13932
rect 8288 13920 8300 13929
rect 8255 13892 8300 13920
rect 8288 13883 8300 13892
rect 8294 13880 8300 13883
rect 8352 13880 8358 13932
rect 9490 13880 9496 13932
rect 9548 13920 9554 13932
rect 9953 13923 10011 13929
rect 9953 13920 9965 13923
rect 9548 13892 9965 13920
rect 9548 13880 9554 13892
rect 9953 13889 9965 13892
rect 9999 13889 10011 13923
rect 9953 13883 10011 13889
rect 9968 13852 9996 13883
rect 10134 13880 10140 13932
rect 10192 13880 10198 13932
rect 10594 13880 10600 13932
rect 10652 13880 10658 13932
rect 10965 13923 11023 13929
rect 10965 13920 10977 13923
rect 10704 13892 10977 13920
rect 10413 13855 10471 13861
rect 10413 13852 10425 13855
rect 5920 13824 6776 13852
rect 9968 13824 10425 13852
rect 4203 13821 4215 13824
rect 4157 13815 4215 13821
rect 3602 13744 3608 13796
rect 3660 13784 3666 13796
rect 4338 13784 4344 13796
rect 3660 13756 4344 13784
rect 3660 13744 3666 13756
rect 4338 13744 4344 13756
rect 4396 13784 4402 13796
rect 4890 13784 4896 13796
rect 4396 13756 4896 13784
rect 4396 13744 4402 13756
rect 4890 13744 4896 13756
rect 4948 13744 4954 13796
rect 6638 13744 6644 13796
rect 6696 13744 6702 13796
rect 6748 13793 6776 13824
rect 10413 13821 10425 13824
rect 10459 13821 10471 13855
rect 10413 13815 10471 13821
rect 10502 13812 10508 13864
rect 10560 13852 10566 13864
rect 10704 13852 10732 13892
rect 10965 13889 10977 13892
rect 11011 13920 11023 13923
rect 11238 13920 11244 13932
rect 11011 13892 11244 13920
rect 11011 13889 11023 13892
rect 10965 13883 11023 13889
rect 11238 13880 11244 13892
rect 11296 13880 11302 13932
rect 11333 13923 11391 13929
rect 11333 13889 11345 13923
rect 11379 13920 11391 13923
rect 12066 13920 12072 13932
rect 11379 13892 12072 13920
rect 11379 13889 11391 13892
rect 11333 13883 11391 13889
rect 12066 13880 12072 13892
rect 12124 13880 12130 13932
rect 12713 13923 12771 13929
rect 12713 13889 12725 13923
rect 12759 13920 12771 13923
rect 13173 13923 13231 13929
rect 13173 13920 13185 13923
rect 12759 13892 13185 13920
rect 12759 13889 12771 13892
rect 12713 13883 12771 13889
rect 13173 13889 13185 13892
rect 13219 13889 13231 13923
rect 13173 13883 13231 13889
rect 13906 13880 13912 13932
rect 13964 13880 13970 13932
rect 14292 13929 14320 13960
rect 14820 13957 14832 13991
rect 14866 13988 14878 13991
rect 15102 13988 15108 14000
rect 14866 13960 15108 13988
rect 14866 13957 14878 13960
rect 14820 13951 14878 13957
rect 15102 13948 15108 13960
rect 15160 13948 15166 14000
rect 14185 13923 14243 13929
rect 14185 13889 14197 13923
rect 14231 13889 14243 13923
rect 14185 13883 14243 13889
rect 14277 13923 14335 13929
rect 14277 13889 14289 13923
rect 14323 13889 14335 13923
rect 14277 13883 14335 13889
rect 10560 13824 10732 13852
rect 10560 13812 10566 13824
rect 10778 13812 10784 13864
rect 10836 13852 10842 13864
rect 11517 13855 11575 13861
rect 11517 13852 11529 13855
rect 10836 13824 11529 13852
rect 10836 13812 10842 13824
rect 11517 13821 11529 13824
rect 11563 13821 11575 13855
rect 11517 13815 11575 13821
rect 12434 13812 12440 13864
rect 12492 13852 12498 13864
rect 12897 13855 12955 13861
rect 12897 13852 12909 13855
rect 12492 13824 12909 13852
rect 12492 13812 12498 13824
rect 12897 13821 12909 13824
rect 12943 13821 12955 13855
rect 12897 13815 12955 13821
rect 13814 13812 13820 13864
rect 13872 13812 13878 13864
rect 14200 13852 14228 13883
rect 16022 13880 16028 13932
rect 16080 13880 16086 13932
rect 14366 13852 14372 13864
rect 14200 13824 14372 13852
rect 14366 13812 14372 13824
rect 14424 13812 14430 13864
rect 14550 13812 14556 13864
rect 14608 13812 14614 13864
rect 6733 13787 6791 13793
rect 6733 13753 6745 13787
rect 6779 13753 6791 13787
rect 6733 13747 6791 13753
rect 13998 13744 14004 13796
rect 14056 13784 14062 13796
rect 14093 13787 14151 13793
rect 14093 13784 14105 13787
rect 14056 13756 14105 13784
rect 14056 13744 14062 13756
rect 14093 13753 14105 13756
rect 14139 13753 14151 13787
rect 14093 13747 14151 13753
rect 1946 13676 1952 13728
rect 2004 13676 2010 13728
rect 3513 13719 3571 13725
rect 3513 13685 3525 13719
rect 3559 13716 3571 13719
rect 3694 13716 3700 13728
rect 3559 13688 3700 13716
rect 3559 13685 3571 13688
rect 3513 13679 3571 13685
rect 3694 13676 3700 13688
rect 3752 13676 3758 13728
rect 3881 13719 3939 13725
rect 3881 13685 3893 13719
rect 3927 13716 3939 13719
rect 3970 13716 3976 13728
rect 3927 13688 3976 13716
rect 3927 13685 3939 13688
rect 3881 13679 3939 13685
rect 3970 13676 3976 13688
rect 4028 13676 4034 13728
rect 4062 13676 4068 13728
rect 4120 13676 4126 13728
rect 4430 13676 4436 13728
rect 4488 13716 4494 13728
rect 5350 13716 5356 13728
rect 4488 13688 5356 13716
rect 4488 13676 4494 13688
rect 5350 13676 5356 13688
rect 5408 13676 5414 13728
rect 5810 13676 5816 13728
rect 5868 13716 5874 13728
rect 6503 13719 6561 13725
rect 6503 13716 6515 13719
rect 5868 13688 6515 13716
rect 5868 13676 5874 13688
rect 6503 13685 6515 13688
rect 6549 13685 6561 13719
rect 6503 13679 6561 13685
rect 12158 13676 12164 13728
rect 12216 13676 12222 13728
rect 12250 13676 12256 13728
rect 12308 13716 12314 13728
rect 12345 13719 12403 13725
rect 12345 13716 12357 13719
rect 12308 13688 12357 13716
rect 12308 13676 12314 13688
rect 12345 13685 12357 13688
rect 12391 13685 12403 13719
rect 12345 13679 12403 13685
rect 15654 13676 15660 13728
rect 15712 13716 15718 13728
rect 15933 13719 15991 13725
rect 15933 13716 15945 13719
rect 15712 13688 15945 13716
rect 15712 13676 15718 13688
rect 15933 13685 15945 13688
rect 15979 13685 15991 13719
rect 15933 13679 15991 13685
rect 1104 13626 16652 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 16652 13626
rect 1104 13552 16652 13574
rect 4798 13512 4804 13524
rect 1412 13484 4804 13512
rect 1412 13385 1440 13484
rect 4798 13472 4804 13484
rect 4856 13512 4862 13524
rect 5258 13512 5264 13524
rect 4856 13484 5264 13512
rect 4856 13472 4862 13484
rect 5258 13472 5264 13484
rect 5316 13472 5322 13524
rect 7190 13472 7196 13524
rect 7248 13472 7254 13524
rect 12986 13472 12992 13524
rect 13044 13512 13050 13524
rect 13906 13512 13912 13524
rect 13044 13484 13912 13512
rect 13044 13472 13050 13484
rect 13906 13472 13912 13484
rect 13964 13512 13970 13524
rect 15102 13512 15108 13524
rect 13964 13484 15108 13512
rect 13964 13472 13970 13484
rect 15102 13472 15108 13484
rect 15160 13512 15166 13524
rect 15160 13484 15332 13512
rect 15160 13472 15166 13484
rect 2406 13404 2412 13456
rect 2464 13444 2470 13456
rect 2777 13447 2835 13453
rect 2777 13444 2789 13447
rect 2464 13416 2789 13444
rect 2464 13404 2470 13416
rect 2777 13413 2789 13416
rect 2823 13413 2835 13447
rect 2777 13407 2835 13413
rect 1397 13379 1455 13385
rect 1397 13345 1409 13379
rect 1443 13345 1455 13379
rect 2792 13376 2820 13407
rect 3142 13404 3148 13456
rect 3200 13444 3206 13456
rect 3237 13447 3295 13453
rect 3237 13444 3249 13447
rect 3200 13416 3249 13444
rect 3200 13404 3206 13416
rect 3237 13413 3249 13416
rect 3283 13444 3295 13447
rect 4157 13447 4215 13453
rect 3283 13416 4016 13444
rect 3283 13413 3295 13416
rect 3237 13407 3295 13413
rect 3329 13379 3387 13385
rect 3329 13376 3341 13379
rect 2792 13348 3341 13376
rect 1397 13339 1455 13345
rect 3329 13345 3341 13348
rect 3375 13345 3387 13379
rect 3329 13339 3387 13345
rect 2866 13268 2872 13320
rect 2924 13308 2930 13320
rect 2961 13311 3019 13317
rect 2961 13308 2973 13311
rect 2924 13280 2973 13308
rect 2924 13268 2930 13280
rect 2961 13277 2973 13280
rect 3007 13277 3019 13311
rect 2961 13271 3019 13277
rect 3050 13268 3056 13320
rect 3108 13308 3114 13320
rect 3513 13311 3571 13317
rect 3513 13308 3525 13311
rect 3108 13280 3525 13308
rect 3108 13268 3114 13280
rect 3513 13277 3525 13280
rect 3559 13277 3571 13311
rect 3513 13271 3571 13277
rect 3602 13268 3608 13320
rect 3660 13268 3666 13320
rect 3988 13317 4016 13416
rect 4157 13413 4169 13447
rect 4203 13444 4215 13447
rect 4246 13444 4252 13456
rect 4203 13416 4252 13444
rect 4203 13413 4215 13416
rect 4157 13407 4215 13413
rect 4246 13404 4252 13416
rect 4304 13404 4310 13456
rect 7282 13444 7288 13456
rect 7208 13416 7288 13444
rect 4065 13379 4123 13385
rect 4065 13345 4077 13379
rect 4111 13376 4123 13379
rect 4890 13376 4896 13388
rect 4111 13348 4896 13376
rect 4111 13345 4123 13348
rect 4065 13339 4123 13345
rect 4890 13336 4896 13348
rect 4948 13336 4954 13388
rect 5258 13336 5264 13388
rect 5316 13376 5322 13388
rect 5353 13379 5411 13385
rect 5353 13376 5365 13379
rect 5316 13348 5365 13376
rect 5316 13336 5322 13348
rect 5353 13345 5365 13348
rect 5399 13345 5411 13379
rect 5353 13339 5411 13345
rect 5994 13336 6000 13388
rect 6052 13376 6058 13388
rect 7208 13385 7236 13416
rect 7282 13404 7288 13416
rect 7340 13404 7346 13456
rect 11514 13444 11520 13456
rect 10980 13416 11520 13444
rect 6089 13379 6147 13385
rect 6089 13376 6101 13379
rect 6052 13348 6101 13376
rect 6052 13336 6058 13348
rect 6089 13345 6101 13348
rect 6135 13345 6147 13379
rect 6089 13339 6147 13345
rect 7193 13379 7251 13385
rect 7193 13345 7205 13379
rect 7239 13345 7251 13379
rect 7193 13339 7251 13345
rect 3789 13311 3847 13317
rect 3789 13308 3801 13311
rect 3703 13280 3801 13308
rect 1670 13249 1676 13252
rect 1664 13203 1676 13249
rect 1670 13200 1676 13203
rect 1728 13200 1734 13252
rect 3234 13200 3240 13252
rect 3292 13200 3298 13252
rect 3329 13243 3387 13249
rect 3329 13209 3341 13243
rect 3375 13240 3387 13243
rect 3418 13240 3424 13252
rect 3375 13212 3424 13240
rect 3375 13209 3387 13212
rect 3329 13203 3387 13209
rect 3418 13200 3424 13212
rect 3476 13200 3482 13252
rect 2866 13132 2872 13184
rect 2924 13172 2930 13184
rect 3053 13175 3111 13181
rect 3053 13172 3065 13175
rect 2924 13144 3065 13172
rect 2924 13132 2930 13144
rect 3053 13141 3065 13144
rect 3099 13141 3111 13175
rect 3053 13135 3111 13141
rect 3510 13132 3516 13184
rect 3568 13172 3574 13184
rect 3703 13172 3731 13280
rect 3789 13277 3801 13280
rect 3835 13277 3847 13311
rect 3789 13271 3847 13277
rect 3973 13311 4031 13317
rect 3973 13277 3985 13311
rect 4019 13277 4031 13311
rect 3973 13271 4031 13277
rect 4246 13268 4252 13320
rect 4304 13268 4310 13320
rect 4617 13311 4675 13317
rect 4617 13277 4629 13311
rect 4663 13308 4675 13311
rect 7006 13308 7012 13320
rect 4663 13280 7012 13308
rect 4663 13277 4675 13280
rect 4617 13271 4675 13277
rect 7006 13268 7012 13280
rect 7064 13268 7070 13320
rect 7282 13268 7288 13320
rect 7340 13268 7346 13320
rect 7466 13268 7472 13320
rect 7524 13308 7530 13320
rect 8202 13308 8208 13320
rect 7524 13280 8208 13308
rect 7524 13268 7530 13280
rect 8202 13268 8208 13280
rect 8260 13268 8266 13320
rect 8294 13268 8300 13320
rect 8352 13308 8358 13320
rect 8389 13311 8447 13317
rect 8389 13308 8401 13311
rect 8352 13280 8401 13308
rect 8352 13268 8358 13280
rect 8389 13277 8401 13280
rect 8435 13277 8447 13311
rect 8389 13271 8447 13277
rect 9674 13268 9680 13320
rect 9732 13308 9738 13320
rect 9858 13308 9864 13320
rect 9732 13280 9864 13308
rect 9732 13268 9738 13280
rect 9858 13268 9864 13280
rect 9916 13268 9922 13320
rect 9950 13268 9956 13320
rect 10008 13308 10014 13320
rect 10229 13311 10287 13317
rect 10229 13308 10241 13311
rect 10008 13280 10241 13308
rect 10008 13268 10014 13280
rect 10229 13277 10241 13280
rect 10275 13277 10287 13311
rect 10229 13271 10287 13277
rect 10321 13311 10379 13317
rect 10321 13277 10333 13311
rect 10367 13308 10379 13311
rect 10594 13308 10600 13320
rect 10367 13280 10600 13308
rect 10367 13277 10379 13280
rect 10321 13271 10379 13277
rect 10594 13268 10600 13280
rect 10652 13268 10658 13320
rect 10686 13268 10692 13320
rect 10744 13268 10750 13320
rect 6822 13200 6828 13252
rect 6880 13200 6886 13252
rect 10505 13243 10563 13249
rect 10505 13209 10517 13243
rect 10551 13240 10563 13243
rect 10980 13240 11008 13416
rect 11514 13404 11520 13416
rect 11572 13444 11578 13456
rect 13357 13447 13415 13453
rect 11572 13416 11744 13444
rect 11572 13404 11578 13416
rect 11054 13336 11060 13388
rect 11112 13376 11118 13388
rect 11112 13348 11652 13376
rect 11112 13336 11118 13348
rect 11624 13317 11652 13348
rect 11716 13317 11744 13416
rect 13357 13413 13369 13447
rect 13403 13444 13415 13447
rect 13814 13444 13820 13456
rect 13403 13416 13820 13444
rect 13403 13413 13415 13416
rect 13357 13407 13415 13413
rect 13814 13404 13820 13416
rect 13872 13444 13878 13456
rect 14182 13444 14188 13456
rect 13872 13416 14188 13444
rect 13872 13404 13878 13416
rect 14182 13404 14188 13416
rect 14240 13404 14246 13456
rect 15304 13444 15332 13484
rect 15378 13472 15384 13524
rect 15436 13472 15442 13524
rect 15562 13472 15568 13524
rect 15620 13472 15626 13524
rect 15304 13416 15424 13444
rect 14366 13336 14372 13388
rect 14424 13376 14430 13388
rect 14645 13379 14703 13385
rect 14645 13376 14657 13379
rect 14424 13348 14657 13376
rect 14424 13336 14430 13348
rect 14645 13345 14657 13348
rect 14691 13345 14703 13379
rect 15286 13376 15292 13388
rect 14645 13339 14703 13345
rect 15028 13348 15292 13376
rect 11241 13311 11299 13317
rect 11241 13277 11253 13311
rect 11287 13308 11299 13311
rect 11333 13311 11391 13317
rect 11333 13308 11345 13311
rect 11287 13280 11345 13308
rect 11287 13277 11299 13280
rect 11241 13271 11299 13277
rect 11333 13277 11345 13280
rect 11379 13277 11391 13311
rect 11333 13271 11391 13277
rect 11609 13311 11667 13317
rect 11609 13277 11621 13311
rect 11655 13277 11667 13311
rect 11609 13271 11667 13277
rect 11701 13311 11759 13317
rect 11701 13277 11713 13311
rect 11747 13277 11759 13311
rect 11701 13271 11759 13277
rect 11974 13268 11980 13320
rect 12032 13268 12038 13320
rect 12250 13317 12256 13320
rect 12244 13308 12256 13317
rect 12211 13280 12256 13308
rect 12244 13271 12256 13280
rect 12250 13268 12256 13271
rect 12308 13268 12314 13320
rect 13909 13311 13967 13317
rect 13909 13277 13921 13311
rect 13955 13308 13967 13311
rect 14090 13308 14096 13320
rect 13955 13280 14096 13308
rect 13955 13277 13967 13280
rect 13909 13271 13967 13277
rect 14090 13268 14096 13280
rect 14148 13268 14154 13320
rect 15028 13317 15056 13348
rect 15286 13336 15292 13348
rect 15344 13336 15350 13388
rect 15013 13311 15071 13317
rect 15013 13277 15025 13311
rect 15059 13277 15071 13311
rect 15013 13271 15071 13277
rect 15194 13268 15200 13320
rect 15252 13268 15258 13320
rect 15396 13308 15424 13416
rect 15749 13311 15807 13317
rect 15749 13308 15761 13311
rect 15396 13280 15761 13308
rect 15749 13277 15761 13280
rect 15795 13277 15807 13311
rect 15749 13271 15807 13277
rect 16114 13268 16120 13320
rect 16172 13268 16178 13320
rect 10551 13212 11008 13240
rect 11517 13243 11575 13249
rect 10551 13209 10563 13212
rect 10505 13203 10563 13209
rect 11517 13209 11529 13243
rect 11563 13209 11575 13243
rect 11517 13203 11575 13209
rect 13740 13212 14688 13240
rect 3568 13144 3731 13172
rect 3568 13132 3574 13144
rect 4154 13132 4160 13184
rect 4212 13172 4218 13184
rect 4433 13175 4491 13181
rect 4433 13172 4445 13175
rect 4212 13144 4445 13172
rect 4212 13132 4218 13144
rect 4433 13141 4445 13144
rect 4479 13141 4491 13175
rect 4433 13135 4491 13141
rect 6546 13132 6552 13184
rect 6604 13172 6610 13184
rect 6733 13175 6791 13181
rect 6733 13172 6745 13175
rect 6604 13144 6745 13172
rect 6604 13132 6610 13144
rect 6733 13141 6745 13144
rect 6779 13141 6791 13175
rect 6733 13135 6791 13141
rect 7374 13132 7380 13184
rect 7432 13172 7438 13184
rect 7469 13175 7527 13181
rect 7469 13172 7481 13175
rect 7432 13144 7481 13172
rect 7432 13132 7438 13144
rect 7469 13141 7481 13144
rect 7515 13141 7527 13175
rect 7469 13135 7527 13141
rect 7742 13132 7748 13184
rect 7800 13172 7806 13184
rect 7837 13175 7895 13181
rect 7837 13172 7849 13175
rect 7800 13144 7849 13172
rect 7800 13132 7806 13144
rect 7837 13141 7849 13144
rect 7883 13141 7895 13175
rect 7837 13135 7895 13141
rect 9766 13132 9772 13184
rect 9824 13172 9830 13184
rect 10045 13175 10103 13181
rect 10045 13172 10057 13175
rect 9824 13144 10057 13172
rect 9824 13132 9830 13144
rect 10045 13141 10057 13144
rect 10091 13141 10103 13175
rect 10045 13135 10103 13141
rect 10413 13175 10471 13181
rect 10413 13141 10425 13175
rect 10459 13172 10471 13175
rect 11532 13172 11560 13203
rect 10459 13144 11560 13172
rect 10459 13141 10471 13144
rect 10413 13135 10471 13141
rect 11790 13132 11796 13184
rect 11848 13172 11854 13184
rect 13740 13181 13768 13212
rect 14660 13184 14688 13212
rect 14734 13200 14740 13252
rect 14792 13240 14798 13252
rect 14829 13243 14887 13249
rect 14829 13240 14841 13243
rect 14792 13212 14841 13240
rect 14792 13200 14798 13212
rect 14829 13209 14841 13212
rect 14875 13209 14887 13243
rect 14829 13203 14887 13209
rect 15286 13200 15292 13252
rect 15344 13240 15350 13252
rect 15841 13243 15899 13249
rect 15841 13240 15853 13243
rect 15344 13212 15853 13240
rect 15344 13200 15350 13212
rect 15841 13209 15853 13212
rect 15887 13209 15899 13243
rect 15841 13203 15899 13209
rect 15933 13243 15991 13249
rect 15933 13209 15945 13243
rect 15979 13209 15991 13243
rect 15933 13203 15991 13209
rect 11885 13175 11943 13181
rect 11885 13172 11897 13175
rect 11848 13144 11897 13172
rect 11848 13132 11854 13144
rect 11885 13141 11897 13144
rect 11931 13141 11943 13175
rect 11885 13135 11943 13141
rect 13725 13175 13783 13181
rect 13725 13141 13737 13175
rect 13771 13141 13783 13175
rect 13725 13135 13783 13141
rect 14090 13132 14096 13184
rect 14148 13132 14154 13184
rect 14642 13132 14648 13184
rect 14700 13172 14706 13184
rect 15746 13172 15752 13184
rect 14700 13144 15752 13172
rect 14700 13132 14706 13144
rect 15746 13132 15752 13144
rect 15804 13172 15810 13184
rect 15948 13172 15976 13203
rect 15804 13144 15976 13172
rect 15804 13132 15810 13144
rect 1104 13082 16652 13104
rect 1104 13030 4874 13082
rect 4926 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 16652 13082
rect 1104 13008 16652 13030
rect 1581 12971 1639 12977
rect 1581 12937 1593 12971
rect 1627 12968 1639 12971
rect 1670 12968 1676 12980
rect 1627 12940 1676 12968
rect 1627 12937 1639 12940
rect 1581 12931 1639 12937
rect 1670 12928 1676 12940
rect 1728 12928 1734 12980
rect 1857 12971 1915 12977
rect 1857 12937 1869 12971
rect 1903 12968 1915 12971
rect 1946 12968 1952 12980
rect 1903 12940 1952 12968
rect 1903 12937 1915 12940
rect 1857 12931 1915 12937
rect 1946 12928 1952 12940
rect 2004 12928 2010 12980
rect 3421 12971 3479 12977
rect 3421 12937 3433 12971
rect 3467 12968 3479 12971
rect 3786 12968 3792 12980
rect 3467 12940 3792 12968
rect 3467 12937 3479 12940
rect 3421 12931 3479 12937
rect 3786 12928 3792 12940
rect 3844 12968 3850 12980
rect 4985 12971 5043 12977
rect 3844 12940 3924 12968
rect 3844 12928 3850 12940
rect 1765 12903 1823 12909
rect 1765 12869 1777 12903
rect 1811 12900 1823 12903
rect 2225 12903 2283 12909
rect 2225 12900 2237 12903
rect 1811 12872 2237 12900
rect 1811 12869 1823 12872
rect 1765 12863 1823 12869
rect 2225 12869 2237 12872
rect 2271 12869 2283 12903
rect 2225 12863 2283 12869
rect 2406 12860 2412 12912
rect 2464 12860 2470 12912
rect 2777 12903 2835 12909
rect 2777 12869 2789 12903
rect 2823 12900 2835 12903
rect 2866 12900 2872 12912
rect 2823 12872 2872 12900
rect 2823 12869 2835 12872
rect 2777 12863 2835 12869
rect 2866 12860 2872 12872
rect 2924 12900 2930 12912
rect 3896 12909 3924 12940
rect 4985 12937 4997 12971
rect 5031 12968 5043 12971
rect 5718 12968 5724 12980
rect 5031 12940 5724 12968
rect 5031 12937 5043 12940
rect 4985 12931 5043 12937
rect 5718 12928 5724 12940
rect 5776 12928 5782 12980
rect 5810 12928 5816 12980
rect 5868 12928 5874 12980
rect 6457 12971 6515 12977
rect 6457 12937 6469 12971
rect 6503 12968 6515 12971
rect 7282 12968 7288 12980
rect 6503 12940 7288 12968
rect 6503 12937 6515 12940
rect 6457 12931 6515 12937
rect 7282 12928 7288 12940
rect 7340 12968 7346 12980
rect 8205 12971 8263 12977
rect 8205 12968 8217 12971
rect 7340 12940 8217 12968
rect 7340 12928 7346 12940
rect 8205 12937 8217 12940
rect 8251 12937 8263 12971
rect 8205 12931 8263 12937
rect 8294 12928 8300 12980
rect 8352 12928 8358 12980
rect 10413 12971 10471 12977
rect 10413 12937 10425 12971
rect 10459 12937 10471 12971
rect 10413 12931 10471 12937
rect 3881 12903 3939 12909
rect 2924 12872 3372 12900
rect 2924 12860 2930 12872
rect 1854 12792 1860 12844
rect 1912 12832 1918 12844
rect 1949 12835 2007 12841
rect 1949 12832 1961 12835
rect 1912 12804 1961 12832
rect 1912 12792 1918 12804
rect 1949 12801 1961 12804
rect 1995 12801 2007 12835
rect 1949 12795 2007 12801
rect 2038 12792 2044 12844
rect 2096 12832 2102 12844
rect 2593 12835 2651 12841
rect 2593 12832 2605 12835
rect 2096 12804 2605 12832
rect 2096 12792 2102 12804
rect 2516 12776 2544 12804
rect 2593 12801 2605 12804
rect 2639 12801 2651 12835
rect 2593 12795 2651 12801
rect 2685 12835 2743 12841
rect 2685 12801 2697 12835
rect 2731 12832 2743 12835
rect 2961 12835 3019 12841
rect 2731 12804 2820 12832
rect 2731 12801 2743 12804
rect 2685 12795 2743 12801
rect 2792 12776 2820 12804
rect 2961 12801 2973 12835
rect 3007 12832 3019 12835
rect 3007 12804 3041 12832
rect 3007 12801 3019 12804
rect 2961 12795 3019 12801
rect 2133 12767 2191 12773
rect 2133 12733 2145 12767
rect 2179 12764 2191 12767
rect 2314 12764 2320 12776
rect 2179 12736 2320 12764
rect 2179 12733 2191 12736
rect 2133 12727 2191 12733
rect 2314 12724 2320 12736
rect 2372 12724 2378 12776
rect 2498 12724 2504 12776
rect 2556 12724 2562 12776
rect 2774 12724 2780 12776
rect 2832 12724 2838 12776
rect 2976 12764 3004 12795
rect 3142 12792 3148 12844
rect 3200 12832 3206 12844
rect 3237 12835 3295 12841
rect 3237 12832 3249 12835
rect 3200 12804 3249 12832
rect 3200 12792 3206 12804
rect 3237 12801 3249 12804
rect 3283 12801 3295 12835
rect 3237 12795 3295 12801
rect 3053 12767 3111 12773
rect 3053 12764 3065 12767
rect 2884 12736 3065 12764
rect 2332 12696 2360 12724
rect 2590 12696 2596 12708
rect 2332 12668 2596 12696
rect 2590 12656 2596 12668
rect 2648 12656 2654 12708
rect 2884 12628 2912 12736
rect 3053 12733 3065 12736
rect 3099 12733 3111 12767
rect 3344 12764 3372 12872
rect 3881 12869 3893 12903
rect 3927 12869 3939 12903
rect 3881 12863 3939 12869
rect 4801 12903 4859 12909
rect 4801 12869 4813 12903
rect 4847 12900 4859 12903
rect 6822 12900 6828 12912
rect 4847 12872 5028 12900
rect 4847 12869 4859 12872
rect 4801 12863 4859 12869
rect 5000 12844 5028 12872
rect 5092 12872 5764 12900
rect 3694 12792 3700 12844
rect 3752 12792 3758 12844
rect 3789 12835 3847 12841
rect 3789 12801 3801 12835
rect 3835 12832 3847 12835
rect 3970 12832 3976 12844
rect 3835 12804 3976 12832
rect 3835 12801 3847 12804
rect 3789 12795 3847 12801
rect 3970 12792 3976 12804
rect 4028 12792 4034 12844
rect 4065 12835 4123 12841
rect 4065 12801 4077 12835
rect 4111 12801 4123 12835
rect 4065 12795 4123 12801
rect 3878 12764 3884 12776
rect 3344 12736 3884 12764
rect 3053 12727 3111 12733
rect 3878 12724 3884 12736
rect 3936 12724 3942 12776
rect 2961 12699 3019 12705
rect 2961 12665 2973 12699
rect 3007 12696 3019 12699
rect 4080 12696 4108 12795
rect 4154 12792 4160 12844
rect 4212 12792 4218 12844
rect 4982 12792 4988 12844
rect 5040 12792 5046 12844
rect 5092 12841 5120 12872
rect 5736 12844 5764 12872
rect 6196 12872 6828 12900
rect 5077 12835 5135 12841
rect 5077 12801 5089 12835
rect 5123 12801 5135 12835
rect 5077 12795 5135 12801
rect 5261 12835 5319 12841
rect 5261 12801 5273 12835
rect 5307 12832 5319 12835
rect 5534 12832 5540 12844
rect 5307 12804 5540 12832
rect 5307 12801 5319 12804
rect 5261 12795 5319 12801
rect 5534 12792 5540 12804
rect 5592 12792 5598 12844
rect 5626 12792 5632 12844
rect 5684 12792 5690 12844
rect 5718 12792 5724 12844
rect 5776 12792 5782 12844
rect 5902 12792 5908 12844
rect 5960 12832 5966 12844
rect 6196 12841 6224 12872
rect 6822 12860 6828 12872
rect 6880 12860 6886 12912
rect 10428 12900 10456 12931
rect 10686 12928 10692 12980
rect 10744 12968 10750 12980
rect 10873 12971 10931 12977
rect 10873 12968 10885 12971
rect 10744 12940 10885 12968
rect 10744 12928 10750 12940
rect 10873 12937 10885 12940
rect 10919 12937 10931 12971
rect 10873 12931 10931 12937
rect 11885 12971 11943 12977
rect 11885 12937 11897 12971
rect 11931 12968 11943 12971
rect 12158 12968 12164 12980
rect 11931 12940 12164 12968
rect 11931 12937 11943 12940
rect 11885 12931 11943 12937
rect 12158 12928 12164 12940
rect 12216 12928 12222 12980
rect 12805 12971 12863 12977
rect 12805 12937 12817 12971
rect 12851 12968 12863 12971
rect 13633 12971 13691 12977
rect 12851 12940 13492 12968
rect 12851 12937 12863 12940
rect 12805 12931 12863 12937
rect 7024 12872 8156 12900
rect 5997 12835 6055 12841
rect 5997 12832 6009 12835
rect 5960 12804 6009 12832
rect 5960 12792 5966 12804
rect 5997 12801 6009 12804
rect 6043 12801 6055 12835
rect 5997 12795 6055 12801
rect 6181 12835 6239 12841
rect 6181 12801 6193 12835
rect 6227 12801 6239 12835
rect 6181 12795 6239 12801
rect 6546 12792 6552 12844
rect 6604 12792 6610 12844
rect 5350 12724 5356 12776
rect 5408 12724 5414 12776
rect 5445 12767 5503 12773
rect 5445 12733 5457 12767
rect 5491 12733 5503 12767
rect 5445 12727 5503 12733
rect 6089 12767 6147 12773
rect 6089 12733 6101 12767
rect 6135 12764 6147 12767
rect 6914 12764 6920 12776
rect 6135 12736 6920 12764
rect 6135 12733 6147 12736
rect 6089 12727 6147 12733
rect 3007 12668 4108 12696
rect 4433 12699 4491 12705
rect 3007 12665 3019 12668
rect 2961 12659 3019 12665
rect 4433 12665 4445 12699
rect 4479 12696 4491 12699
rect 4890 12696 4896 12708
rect 4479 12668 4896 12696
rect 4479 12665 4491 12668
rect 4433 12659 4491 12665
rect 4890 12656 4896 12668
rect 4948 12656 4954 12708
rect 3142 12628 3148 12640
rect 2884 12600 3148 12628
rect 3142 12588 3148 12600
rect 3200 12628 3206 12640
rect 3418 12628 3424 12640
rect 3200 12600 3424 12628
rect 3200 12588 3206 12600
rect 3418 12588 3424 12600
rect 3476 12588 3482 12640
rect 3513 12631 3571 12637
rect 3513 12597 3525 12631
rect 3559 12628 3571 12631
rect 3602 12628 3608 12640
rect 3559 12600 3608 12628
rect 3559 12597 3571 12600
rect 3513 12591 3571 12597
rect 3602 12588 3608 12600
rect 3660 12588 3666 12640
rect 4706 12588 4712 12640
rect 4764 12628 4770 12640
rect 4801 12631 4859 12637
rect 4801 12628 4813 12631
rect 4764 12600 4813 12628
rect 4764 12588 4770 12600
rect 4801 12597 4813 12600
rect 4847 12597 4859 12631
rect 4801 12591 4859 12597
rect 5350 12588 5356 12640
rect 5408 12628 5414 12640
rect 5460 12628 5488 12727
rect 6914 12724 6920 12736
rect 6972 12764 6978 12776
rect 7024 12764 7052 12872
rect 7742 12792 7748 12844
rect 7800 12841 7806 12844
rect 7800 12832 7812 12841
rect 7800 12804 7845 12832
rect 7800 12795 7812 12804
rect 7800 12792 7806 12795
rect 8018 12792 8024 12844
rect 8076 12792 8082 12844
rect 8128 12841 8156 12872
rect 8220 12872 10456 12900
rect 8220 12844 8248 12872
rect 10778 12860 10784 12912
rect 10836 12860 10842 12912
rect 12066 12860 12072 12912
rect 12124 12900 12130 12912
rect 13464 12900 13492 12940
rect 13633 12937 13645 12971
rect 13679 12968 13691 12971
rect 14090 12968 14096 12980
rect 13679 12940 14096 12968
rect 13679 12937 13691 12940
rect 13633 12931 13691 12937
rect 14090 12928 14096 12940
rect 14148 12928 14154 12980
rect 15102 12928 15108 12980
rect 15160 12968 15166 12980
rect 15473 12971 15531 12977
rect 15160 12940 15424 12968
rect 15160 12928 15166 12940
rect 12124 12872 13124 12900
rect 13464 12872 14136 12900
rect 12124 12860 12130 12872
rect 8113 12835 8171 12841
rect 8113 12801 8125 12835
rect 8159 12801 8171 12835
rect 8113 12795 8171 12801
rect 8202 12792 8208 12844
rect 8260 12792 8266 12844
rect 9033 12835 9091 12841
rect 9033 12801 9045 12835
rect 9079 12832 9091 12835
rect 9493 12835 9551 12841
rect 9493 12832 9505 12835
rect 9079 12804 9505 12832
rect 9079 12801 9091 12804
rect 9033 12795 9091 12801
rect 9493 12801 9505 12804
rect 9539 12801 9551 12835
rect 9493 12795 9551 12801
rect 11977 12835 12035 12841
rect 11977 12801 11989 12835
rect 12023 12832 12035 12835
rect 12342 12832 12348 12844
rect 12023 12804 12348 12832
rect 12023 12801 12035 12804
rect 11977 12795 12035 12801
rect 12342 12792 12348 12804
rect 12400 12792 12406 12844
rect 13096 12832 13124 12872
rect 14108 12841 14136 12872
rect 14182 12860 14188 12912
rect 14240 12900 14246 12912
rect 15396 12900 15424 12940
rect 15473 12937 15485 12971
rect 15519 12968 15531 12971
rect 16022 12968 16028 12980
rect 15519 12940 16028 12968
rect 15519 12937 15531 12940
rect 15473 12931 15531 12937
rect 16022 12928 16028 12940
rect 16080 12928 16086 12980
rect 14240 12872 15332 12900
rect 15396 12872 15976 12900
rect 14240 12860 14246 12872
rect 14093 12835 14151 12841
rect 13096 12804 13860 12832
rect 8573 12767 8631 12773
rect 8573 12764 8585 12767
rect 6972 12736 7052 12764
rect 8220 12736 8585 12764
rect 6972 12724 6978 12736
rect 8220 12708 8248 12736
rect 8573 12733 8585 12736
rect 8619 12733 8631 12767
rect 8573 12727 8631 12733
rect 9122 12724 9128 12776
rect 9180 12724 9186 12776
rect 9306 12724 9312 12776
rect 9364 12724 9370 12776
rect 9950 12724 9956 12776
rect 10008 12764 10014 12776
rect 10045 12767 10103 12773
rect 10045 12764 10057 12767
rect 10008 12736 10057 12764
rect 10008 12724 10014 12736
rect 10045 12733 10057 12736
rect 10091 12733 10103 12767
rect 10045 12727 10103 12733
rect 10965 12767 11023 12773
rect 10965 12733 10977 12767
rect 11011 12733 11023 12767
rect 10965 12727 11023 12733
rect 5994 12656 6000 12708
rect 6052 12696 6058 12708
rect 6641 12699 6699 12705
rect 6641 12696 6653 12699
rect 6052 12668 6653 12696
rect 6052 12656 6058 12668
rect 6641 12665 6653 12668
rect 6687 12665 6699 12699
rect 6641 12659 6699 12665
rect 8202 12656 8208 12708
rect 8260 12656 8266 12708
rect 9858 12656 9864 12708
rect 9916 12696 9922 12708
rect 10980 12696 11008 12727
rect 12066 12724 12072 12776
rect 12124 12724 12130 12776
rect 12618 12724 12624 12776
rect 12676 12764 12682 12776
rect 13096 12773 13124 12804
rect 12897 12767 12955 12773
rect 12897 12764 12909 12767
rect 12676 12736 12909 12764
rect 12676 12724 12682 12736
rect 12897 12733 12909 12736
rect 12943 12733 12955 12767
rect 12897 12727 12955 12733
rect 13081 12767 13139 12773
rect 13081 12733 13093 12767
rect 13127 12733 13139 12767
rect 13081 12727 13139 12733
rect 13630 12724 13636 12776
rect 13688 12764 13694 12776
rect 13832 12773 13860 12804
rect 14093 12801 14105 12835
rect 14139 12801 14151 12835
rect 14093 12795 14151 12801
rect 14366 12792 14372 12844
rect 14424 12832 14430 12844
rect 14829 12835 14887 12841
rect 14829 12832 14841 12835
rect 14424 12804 14841 12832
rect 14424 12792 14430 12804
rect 14829 12801 14841 12804
rect 14875 12801 14887 12835
rect 14829 12795 14887 12801
rect 14918 12792 14924 12844
rect 14976 12792 14982 12844
rect 15304 12841 15332 12872
rect 15105 12835 15163 12841
rect 15105 12801 15117 12835
rect 15151 12801 15163 12835
rect 15105 12795 15163 12801
rect 15289 12835 15347 12841
rect 15289 12801 15301 12835
rect 15335 12801 15347 12835
rect 15289 12795 15347 12801
rect 15565 12835 15623 12841
rect 15565 12801 15577 12835
rect 15611 12832 15623 12835
rect 15654 12832 15660 12844
rect 15611 12804 15660 12832
rect 15611 12801 15623 12804
rect 15565 12795 15623 12801
rect 13725 12767 13783 12773
rect 13725 12764 13737 12767
rect 13688 12736 13737 12764
rect 13688 12724 13694 12736
rect 13725 12733 13737 12736
rect 13771 12733 13783 12767
rect 13725 12727 13783 12733
rect 13817 12767 13875 12773
rect 13817 12733 13829 12767
rect 13863 12733 13875 12767
rect 13817 12727 13875 12733
rect 14642 12724 14648 12776
rect 14700 12724 14706 12776
rect 14734 12724 14740 12776
rect 14792 12764 14798 12776
rect 15120 12764 15148 12795
rect 14792 12736 15148 12764
rect 14792 12724 14798 12736
rect 15194 12724 15200 12776
rect 15252 12764 15258 12776
rect 15580 12764 15608 12795
rect 15654 12792 15660 12804
rect 15712 12792 15718 12844
rect 15746 12792 15752 12844
rect 15804 12792 15810 12844
rect 15838 12792 15844 12844
rect 15896 12792 15902 12844
rect 15948 12841 15976 12872
rect 15933 12835 15991 12841
rect 15933 12801 15945 12835
rect 15979 12801 15991 12835
rect 15933 12795 15991 12801
rect 15252 12736 15608 12764
rect 15252 12724 15258 12736
rect 9916 12668 11008 12696
rect 9916 12656 9922 12668
rect 12342 12656 12348 12708
rect 12400 12696 12406 12708
rect 13265 12699 13323 12705
rect 13265 12696 13277 12699
rect 12400 12668 13277 12696
rect 12400 12656 12406 12668
rect 13265 12665 13277 12668
rect 13311 12665 13323 12699
rect 13265 12659 13323 12665
rect 13538 12656 13544 12708
rect 13596 12696 13602 12708
rect 16117 12699 16175 12705
rect 16117 12696 16129 12699
rect 13596 12668 16129 12696
rect 13596 12656 13602 12668
rect 16117 12665 16129 12668
rect 16163 12665 16175 12699
rect 16117 12659 16175 12665
rect 5408 12600 5488 12628
rect 5408 12588 5414 12600
rect 5534 12588 5540 12640
rect 5592 12628 5598 12640
rect 7006 12628 7012 12640
rect 5592 12600 7012 12628
rect 5592 12588 5598 12600
rect 7006 12588 7012 12600
rect 7064 12628 7070 12640
rect 8110 12628 8116 12640
rect 7064 12600 8116 12628
rect 7064 12588 7070 12600
rect 8110 12588 8116 12600
rect 8168 12588 8174 12640
rect 8294 12588 8300 12640
rect 8352 12628 8358 12640
rect 8665 12631 8723 12637
rect 8665 12628 8677 12631
rect 8352 12600 8677 12628
rect 8352 12588 8358 12600
rect 8665 12597 8677 12600
rect 8711 12597 8723 12631
rect 8665 12591 8723 12597
rect 11514 12588 11520 12640
rect 11572 12588 11578 12640
rect 12250 12588 12256 12640
rect 12308 12628 12314 12640
rect 12437 12631 12495 12637
rect 12437 12628 12449 12631
rect 12308 12600 12449 12628
rect 12308 12588 12314 12600
rect 12437 12597 12449 12600
rect 12483 12597 12495 12631
rect 12437 12591 12495 12597
rect 14182 12588 14188 12640
rect 14240 12628 14246 12640
rect 14826 12628 14832 12640
rect 14240 12600 14832 12628
rect 14240 12588 14246 12600
rect 14826 12588 14832 12600
rect 14884 12588 14890 12640
rect 1104 12538 16652 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 16652 12538
rect 1104 12464 16652 12486
rect 2041 12427 2099 12433
rect 2041 12393 2053 12427
rect 2087 12424 2099 12427
rect 3145 12427 3203 12433
rect 2087 12396 2636 12424
rect 2087 12393 2099 12396
rect 2041 12387 2099 12393
rect 2056 12288 2084 12387
rect 1688 12260 2084 12288
rect 2608 12288 2636 12396
rect 3145 12393 3157 12427
rect 3191 12424 3203 12427
rect 3234 12424 3240 12436
rect 3191 12396 3240 12424
rect 3191 12393 3203 12396
rect 3145 12387 3203 12393
rect 3234 12384 3240 12396
rect 3292 12384 3298 12436
rect 5166 12424 5172 12436
rect 4816 12396 5172 12424
rect 3050 12316 3056 12368
rect 3108 12356 3114 12368
rect 3513 12359 3571 12365
rect 3513 12356 3525 12359
rect 3108 12328 3525 12356
rect 3108 12316 3114 12328
rect 3513 12325 3525 12328
rect 3559 12325 3571 12359
rect 3513 12319 3571 12325
rect 4157 12359 4215 12365
rect 4157 12325 4169 12359
rect 4203 12356 4215 12359
rect 4816 12356 4844 12396
rect 5166 12384 5172 12396
rect 5224 12384 5230 12436
rect 5718 12384 5724 12436
rect 5776 12424 5782 12436
rect 6273 12427 6331 12433
rect 6273 12424 6285 12427
rect 5776 12396 6285 12424
rect 5776 12384 5782 12396
rect 6273 12393 6285 12396
rect 6319 12393 6331 12427
rect 6273 12387 6331 12393
rect 6822 12384 6828 12436
rect 6880 12424 6886 12436
rect 8205 12427 8263 12433
rect 8205 12424 8217 12427
rect 6880 12396 8217 12424
rect 6880 12384 6886 12396
rect 8205 12393 8217 12396
rect 8251 12393 8263 12427
rect 8205 12387 8263 12393
rect 4203 12328 4844 12356
rect 4203 12325 4215 12328
rect 4157 12319 4215 12325
rect 2682 12288 2688 12300
rect 2608 12260 2688 12288
rect 1688 12229 1716 12260
rect 1673 12223 1731 12229
rect 1673 12189 1685 12223
rect 1719 12189 1731 12223
rect 1673 12183 1731 12189
rect 1765 12223 1823 12229
rect 1765 12189 1777 12223
rect 1811 12220 1823 12223
rect 2498 12220 2504 12232
rect 1811 12192 2504 12220
rect 1811 12189 1823 12192
rect 1765 12183 1823 12189
rect 1486 12112 1492 12164
rect 1544 12152 1550 12164
rect 2056 12161 2084 12192
rect 2498 12180 2504 12192
rect 2556 12180 2562 12232
rect 2608 12229 2636 12260
rect 2682 12248 2688 12260
rect 2740 12248 2746 12300
rect 2593 12223 2651 12229
rect 2593 12189 2605 12223
rect 2639 12189 2651 12223
rect 3068 12220 3096 12316
rect 3418 12248 3424 12300
rect 3476 12288 3482 12300
rect 3605 12291 3663 12297
rect 3605 12288 3617 12291
rect 3476 12260 3617 12288
rect 3476 12248 3482 12260
rect 3605 12257 3617 12260
rect 3651 12257 3663 12291
rect 3605 12251 3663 12257
rect 6178 12248 6184 12300
rect 6236 12288 6242 12300
rect 6236 12260 6776 12288
rect 6236 12248 6242 12260
rect 2593 12183 2651 12189
rect 2700 12192 3096 12220
rect 3329 12223 3387 12229
rect 2700 12161 2728 12192
rect 3329 12189 3341 12223
rect 3375 12189 3387 12223
rect 3329 12183 3387 12189
rect 4525 12223 4583 12229
rect 4525 12189 4537 12223
rect 4571 12220 4583 12223
rect 4614 12220 4620 12232
rect 4571 12192 4620 12220
rect 4571 12189 4583 12192
rect 4525 12183 4583 12189
rect 1857 12155 1915 12161
rect 1857 12152 1869 12155
rect 1544 12124 1869 12152
rect 1544 12112 1550 12124
rect 1857 12121 1869 12124
rect 1903 12121 1915 12155
rect 2056 12155 2115 12161
rect 2056 12124 2069 12155
rect 1857 12115 1915 12121
rect 2057 12121 2069 12124
rect 2103 12121 2115 12155
rect 2685 12155 2743 12161
rect 2685 12152 2697 12155
rect 2057 12115 2115 12121
rect 2148 12124 2697 12152
rect 1587 12087 1645 12093
rect 1587 12053 1599 12087
rect 1633 12084 1645 12087
rect 1762 12084 1768 12096
rect 1633 12056 1768 12084
rect 1633 12053 1645 12056
rect 1587 12047 1645 12053
rect 1762 12044 1768 12056
rect 1820 12044 1826 12096
rect 1872 12084 1900 12115
rect 2148 12084 2176 12124
rect 2685 12121 2697 12124
rect 2731 12121 2743 12155
rect 2685 12115 2743 12121
rect 2774 12112 2780 12164
rect 2832 12152 2838 12164
rect 2869 12155 2927 12161
rect 2869 12152 2881 12155
rect 2832 12124 2881 12152
rect 2832 12112 2838 12124
rect 2869 12121 2881 12124
rect 2915 12152 2927 12155
rect 3344 12152 3372 12183
rect 4614 12180 4620 12192
rect 4672 12180 4678 12232
rect 4798 12180 4804 12232
rect 4856 12180 4862 12232
rect 6086 12220 6092 12232
rect 5920 12192 6092 12220
rect 3878 12152 3884 12164
rect 2915 12124 3884 12152
rect 2915 12121 2927 12124
rect 2869 12115 2927 12121
rect 3878 12112 3884 12124
rect 3936 12112 3942 12164
rect 4341 12155 4399 12161
rect 4341 12121 4353 12155
rect 4387 12152 4399 12155
rect 4709 12155 4767 12161
rect 4387 12124 4660 12152
rect 4387 12121 4399 12124
rect 4341 12115 4399 12121
rect 1872 12056 2176 12084
rect 2222 12044 2228 12096
rect 2280 12044 2286 12096
rect 2314 12044 2320 12096
rect 2372 12044 2378 12096
rect 3142 12044 3148 12096
rect 3200 12084 3206 12096
rect 3970 12084 3976 12096
rect 3200 12056 3976 12084
rect 3200 12044 3206 12056
rect 3970 12044 3976 12056
rect 4028 12044 4034 12096
rect 4430 12044 4436 12096
rect 4488 12044 4494 12096
rect 4632 12084 4660 12124
rect 4709 12121 4721 12155
rect 4755 12152 4767 12155
rect 4890 12152 4896 12164
rect 4755 12124 4896 12152
rect 4755 12121 4767 12124
rect 4709 12115 4767 12121
rect 4890 12112 4896 12124
rect 4948 12112 4954 12164
rect 5068 12155 5126 12161
rect 5068 12121 5080 12155
rect 5114 12152 5126 12155
rect 5258 12152 5264 12164
rect 5114 12124 5264 12152
rect 5114 12121 5126 12124
rect 5068 12115 5126 12121
rect 5258 12112 5264 12124
rect 5316 12112 5322 12164
rect 5810 12084 5816 12096
rect 4632 12056 5816 12084
rect 5810 12044 5816 12056
rect 5868 12084 5874 12096
rect 5920 12084 5948 12192
rect 6086 12180 6092 12192
rect 6144 12220 6150 12232
rect 6748 12229 6776 12260
rect 6457 12223 6515 12229
rect 6457 12220 6469 12223
rect 6144 12192 6469 12220
rect 6144 12180 6150 12192
rect 6457 12189 6469 12192
rect 6503 12189 6515 12223
rect 6457 12183 6515 12189
rect 6733 12223 6791 12229
rect 6733 12189 6745 12223
rect 6779 12189 6791 12223
rect 6733 12183 6791 12189
rect 6825 12223 6883 12229
rect 6825 12189 6837 12223
rect 6871 12220 6883 12223
rect 8018 12220 8024 12232
rect 6871 12192 8024 12220
rect 6871 12189 6883 12192
rect 6825 12183 6883 12189
rect 8018 12180 8024 12192
rect 8076 12180 8082 12232
rect 8220 12220 8248 12387
rect 9122 12384 9128 12436
rect 9180 12424 9186 12436
rect 9217 12427 9275 12433
rect 9217 12424 9229 12427
rect 9180 12396 9229 12424
rect 9180 12384 9186 12396
rect 9217 12393 9229 12396
rect 9263 12393 9275 12427
rect 9217 12387 9275 12393
rect 10045 12427 10103 12433
rect 10045 12393 10057 12427
rect 10091 12424 10103 12427
rect 10686 12424 10692 12436
rect 10091 12396 10692 12424
rect 10091 12393 10103 12396
rect 10045 12387 10103 12393
rect 10686 12384 10692 12396
rect 10744 12384 10750 12436
rect 11701 12427 11759 12433
rect 11701 12393 11713 12427
rect 11747 12424 11759 12427
rect 15010 12424 15016 12436
rect 11747 12396 15016 12424
rect 11747 12393 11759 12396
rect 11701 12387 11759 12393
rect 15010 12384 15016 12396
rect 15068 12384 15074 12436
rect 13357 12359 13415 12365
rect 13357 12325 13369 12359
rect 13403 12356 13415 12359
rect 13998 12356 14004 12368
rect 13403 12328 14004 12356
rect 13403 12325 13415 12328
rect 13357 12319 13415 12325
rect 13998 12316 14004 12328
rect 14056 12356 14062 12368
rect 14642 12356 14648 12368
rect 14056 12328 14648 12356
rect 14056 12316 14062 12328
rect 14642 12316 14648 12328
rect 14700 12316 14706 12368
rect 9766 12248 9772 12300
rect 9824 12248 9830 12300
rect 11790 12288 11796 12300
rect 11348 12260 11796 12288
rect 8481 12223 8539 12229
rect 8481 12220 8493 12223
rect 8220 12192 8493 12220
rect 8481 12189 8493 12192
rect 8527 12189 8539 12223
rect 8481 12183 8539 12189
rect 9122 12180 9128 12232
rect 9180 12180 9186 12232
rect 9585 12223 9643 12229
rect 9585 12189 9597 12223
rect 9631 12220 9643 12223
rect 10042 12220 10048 12232
rect 9631 12192 10048 12220
rect 9631 12189 9643 12192
rect 9585 12183 9643 12189
rect 10042 12180 10048 12192
rect 10100 12180 10106 12232
rect 11169 12223 11227 12229
rect 11169 12189 11181 12223
rect 11215 12220 11227 12223
rect 11348 12220 11376 12260
rect 11790 12248 11796 12260
rect 11848 12248 11854 12300
rect 11974 12248 11980 12300
rect 12032 12248 12038 12300
rect 13538 12248 13544 12300
rect 13596 12288 13602 12300
rect 15286 12288 15292 12300
rect 13596 12260 15292 12288
rect 13596 12248 13602 12260
rect 15286 12248 15292 12260
rect 15344 12288 15350 12300
rect 15930 12288 15936 12300
rect 15344 12260 15936 12288
rect 15344 12248 15350 12260
rect 15930 12248 15936 12260
rect 15988 12248 15994 12300
rect 11215 12192 11376 12220
rect 11215 12189 11227 12192
rect 11169 12183 11227 12189
rect 11422 12180 11428 12232
rect 11480 12180 11486 12232
rect 11882 12180 11888 12232
rect 11940 12180 11946 12232
rect 11992 12220 12020 12248
rect 13449 12223 13507 12229
rect 13449 12220 13461 12223
rect 11992 12192 13461 12220
rect 13449 12189 13461 12192
rect 13495 12220 13507 12223
rect 13495 12192 13768 12220
rect 13495 12189 13507 12192
rect 13449 12183 13507 12189
rect 5994 12112 6000 12164
rect 6052 12152 6058 12164
rect 7092 12155 7150 12161
rect 6052 12124 6776 12152
rect 6052 12112 6058 12124
rect 6181 12087 6239 12093
rect 6181 12084 6193 12087
rect 5868 12056 6193 12084
rect 5868 12044 5874 12056
rect 6181 12053 6193 12056
rect 6227 12053 6239 12087
rect 6181 12047 6239 12053
rect 6638 12044 6644 12096
rect 6696 12044 6702 12096
rect 6748 12084 6776 12124
rect 7092 12121 7104 12155
rect 7138 12152 7150 12155
rect 7282 12152 7288 12164
rect 7138 12124 7288 12152
rect 7138 12121 7150 12124
rect 7092 12115 7150 12121
rect 7282 12112 7288 12124
rect 7340 12112 7346 12164
rect 12250 12161 12256 12164
rect 8297 12155 8355 12161
rect 8297 12121 8309 12155
rect 8343 12121 8355 12155
rect 8297 12115 8355 12121
rect 12244 12115 12256 12161
rect 8312 12084 8340 12115
rect 12250 12112 12256 12115
rect 12308 12112 12314 12164
rect 13740 12152 13768 12192
rect 13906 12180 13912 12232
rect 13964 12220 13970 12232
rect 14093 12223 14151 12229
rect 14093 12220 14105 12223
rect 13964 12192 14105 12220
rect 13964 12180 13970 12192
rect 14093 12189 14105 12192
rect 14139 12189 14151 12223
rect 14093 12183 14151 12189
rect 14182 12180 14188 12232
rect 14240 12220 14246 12232
rect 15381 12223 15439 12229
rect 15381 12220 15393 12223
rect 14240 12192 15393 12220
rect 14240 12180 14246 12192
rect 15381 12189 15393 12192
rect 15427 12189 15439 12223
rect 15381 12183 15439 12189
rect 15470 12180 15476 12232
rect 15528 12180 15534 12232
rect 15565 12223 15623 12229
rect 15565 12189 15577 12223
rect 15611 12220 15623 12223
rect 15654 12220 15660 12232
rect 15611 12192 15660 12220
rect 15611 12189 15623 12192
rect 15565 12183 15623 12189
rect 15654 12180 15660 12192
rect 15712 12180 15718 12232
rect 15746 12180 15752 12232
rect 15804 12180 15810 12232
rect 14550 12152 14556 12164
rect 13740 12124 14556 12152
rect 14550 12112 14556 12124
rect 14608 12152 14614 12164
rect 14829 12155 14887 12161
rect 14829 12152 14841 12155
rect 14608 12124 14841 12152
rect 14608 12112 14614 12124
rect 14829 12121 14841 12124
rect 14875 12152 14887 12155
rect 14918 12152 14924 12164
rect 14875 12124 14924 12152
rect 14875 12121 14887 12124
rect 14829 12115 14887 12121
rect 14918 12112 14924 12124
rect 14976 12112 14982 12164
rect 15841 12155 15899 12161
rect 15841 12121 15853 12155
rect 15887 12121 15899 12155
rect 15841 12115 15899 12121
rect 6748 12056 8340 12084
rect 8662 12044 8668 12096
rect 8720 12044 8726 12096
rect 9030 12044 9036 12096
rect 9088 12044 9094 12096
rect 9677 12087 9735 12093
rect 9677 12053 9689 12087
rect 9723 12084 9735 12087
rect 10686 12084 10692 12096
rect 9723 12056 10692 12084
rect 9723 12053 9735 12056
rect 9677 12047 9735 12053
rect 10686 12044 10692 12056
rect 10744 12044 10750 12096
rect 11698 12044 11704 12096
rect 11756 12084 11762 12096
rect 13906 12084 13912 12096
rect 11756 12056 13912 12084
rect 11756 12044 11762 12056
rect 13906 12044 13912 12056
rect 13964 12044 13970 12096
rect 14090 12044 14096 12096
rect 14148 12084 14154 12096
rect 14734 12084 14740 12096
rect 14148 12056 14740 12084
rect 14148 12044 14154 12056
rect 14734 12044 14740 12056
rect 14792 12044 14798 12096
rect 15105 12087 15163 12093
rect 15105 12053 15117 12087
rect 15151 12084 15163 12087
rect 15194 12084 15200 12096
rect 15151 12056 15200 12084
rect 15151 12053 15163 12056
rect 15105 12047 15163 12053
rect 15194 12044 15200 12056
rect 15252 12044 15258 12096
rect 15562 12044 15568 12096
rect 15620 12084 15626 12096
rect 15856 12084 15884 12115
rect 16022 12112 16028 12164
rect 16080 12152 16086 12164
rect 16390 12152 16396 12164
rect 16080 12124 16396 12152
rect 16080 12112 16086 12124
rect 16390 12112 16396 12124
rect 16448 12112 16454 12164
rect 15620 12056 15884 12084
rect 15620 12044 15626 12056
rect 16206 12044 16212 12096
rect 16264 12044 16270 12096
rect 1104 11994 16652 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 16652 11994
rect 1104 11920 16652 11942
rect 1397 11883 1455 11889
rect 1397 11849 1409 11883
rect 1443 11880 1455 11883
rect 1486 11880 1492 11892
rect 1443 11852 1492 11880
rect 1443 11849 1455 11852
rect 1397 11843 1455 11849
rect 1486 11840 1492 11852
rect 1544 11840 1550 11892
rect 2222 11840 2228 11892
rect 2280 11880 2286 11892
rect 2866 11880 2872 11892
rect 2280 11852 2872 11880
rect 2280 11840 2286 11852
rect 2866 11840 2872 11852
rect 2924 11840 2930 11892
rect 3513 11883 3571 11889
rect 3513 11880 3525 11883
rect 2976 11852 3525 11880
rect 1854 11772 1860 11824
rect 1912 11812 1918 11824
rect 2976 11812 3004 11852
rect 3513 11849 3525 11852
rect 3559 11849 3571 11883
rect 3513 11843 3571 11849
rect 3970 11840 3976 11892
rect 4028 11880 4034 11892
rect 4341 11883 4399 11889
rect 4341 11880 4353 11883
rect 4028 11852 4353 11880
rect 4028 11840 4034 11852
rect 4341 11849 4353 11852
rect 4387 11849 4399 11883
rect 4341 11843 4399 11849
rect 4430 11840 4436 11892
rect 4488 11880 4494 11892
rect 4890 11880 4896 11892
rect 4488 11852 4896 11880
rect 4488 11840 4494 11852
rect 4890 11840 4896 11852
rect 4948 11840 4954 11892
rect 4985 11883 5043 11889
rect 4985 11849 4997 11883
rect 5031 11880 5043 11883
rect 5258 11880 5264 11892
rect 5031 11852 5264 11880
rect 5031 11849 5043 11852
rect 4985 11843 5043 11849
rect 5258 11840 5264 11852
rect 5316 11840 5322 11892
rect 5997 11883 6055 11889
rect 5997 11849 6009 11883
rect 6043 11880 6055 11883
rect 6178 11880 6184 11892
rect 6043 11852 6184 11880
rect 6043 11849 6055 11852
rect 5997 11843 6055 11849
rect 6178 11840 6184 11852
rect 6236 11840 6242 11892
rect 7127 11883 7185 11889
rect 7127 11849 7139 11883
rect 7173 11880 7185 11883
rect 8662 11880 8668 11892
rect 7173 11852 8668 11880
rect 7173 11849 7185 11852
rect 7127 11843 7185 11849
rect 8662 11840 8668 11852
rect 8720 11840 8726 11892
rect 9953 11883 10011 11889
rect 9953 11849 9965 11883
rect 9999 11880 10011 11883
rect 10778 11880 10784 11892
rect 9999 11852 10784 11880
rect 9999 11849 10011 11852
rect 9953 11843 10011 11849
rect 10778 11840 10784 11852
rect 10836 11840 10842 11892
rect 11882 11840 11888 11892
rect 11940 11880 11946 11892
rect 13538 11880 13544 11892
rect 11940 11852 13544 11880
rect 11940 11840 11946 11852
rect 13538 11840 13544 11852
rect 13596 11840 13602 11892
rect 13633 11883 13691 11889
rect 13633 11849 13645 11883
rect 13679 11880 13691 11883
rect 13722 11880 13728 11892
rect 13679 11852 13728 11880
rect 13679 11849 13691 11852
rect 13633 11843 13691 11849
rect 13722 11840 13728 11852
rect 13780 11840 13786 11892
rect 15102 11880 15108 11892
rect 13832 11852 15108 11880
rect 1912 11784 3004 11812
rect 3037 11815 3095 11821
rect 1912 11772 1918 11784
rect 3037 11781 3049 11815
rect 3083 11812 3095 11815
rect 3142 11812 3148 11824
rect 3083 11784 3148 11812
rect 3083 11781 3095 11784
rect 3037 11775 3095 11781
rect 3142 11772 3148 11784
rect 3200 11772 3206 11824
rect 3234 11772 3240 11824
rect 3292 11772 3298 11824
rect 4798 11812 4804 11824
rect 3344 11784 4804 11812
rect 2521 11747 2579 11753
rect 2521 11713 2533 11747
rect 2567 11744 2579 11747
rect 2777 11748 2835 11753
rect 2777 11747 3004 11748
rect 2567 11716 2728 11744
rect 2567 11713 2579 11716
rect 2521 11707 2579 11713
rect 2700 11676 2728 11716
rect 2777 11713 2789 11747
rect 2823 11744 3004 11747
rect 3344 11744 3372 11784
rect 4798 11772 4804 11784
rect 4856 11772 4862 11824
rect 5074 11772 5080 11824
rect 5132 11812 5138 11824
rect 5169 11815 5227 11821
rect 5169 11812 5181 11815
rect 5132 11784 5181 11812
rect 5132 11772 5138 11784
rect 5169 11781 5181 11784
rect 5215 11781 5227 11815
rect 5169 11775 5227 11781
rect 6454 11772 6460 11824
rect 6512 11812 6518 11824
rect 6917 11815 6975 11821
rect 6917 11812 6929 11815
rect 6512 11784 6929 11812
rect 6512 11772 6518 11784
rect 6917 11781 6929 11784
rect 6963 11781 6975 11815
rect 6917 11775 6975 11781
rect 8104 11815 8162 11821
rect 8104 11781 8116 11815
rect 8150 11812 8162 11815
rect 8294 11812 8300 11824
rect 8150 11784 8300 11812
rect 8150 11781 8162 11784
rect 8104 11775 8162 11781
rect 8294 11772 8300 11784
rect 8352 11772 8358 11824
rect 9858 11772 9864 11824
rect 9916 11772 9922 11824
rect 11088 11815 11146 11821
rect 11088 11781 11100 11815
rect 11134 11812 11146 11815
rect 11514 11812 11520 11824
rect 11134 11784 11520 11812
rect 11134 11781 11146 11784
rect 11088 11775 11146 11781
rect 11514 11772 11520 11784
rect 11572 11772 11578 11824
rect 12342 11821 12348 11824
rect 12336 11812 12348 11821
rect 12303 11784 12348 11812
rect 12336 11775 12348 11784
rect 12342 11772 12348 11775
rect 12400 11772 12406 11824
rect 2823 11720 3372 11744
rect 2823 11713 2835 11720
rect 2976 11716 3372 11720
rect 2777 11707 2835 11713
rect 3418 11704 3424 11756
rect 3476 11704 3482 11756
rect 3510 11704 3516 11756
rect 3568 11744 3574 11756
rect 3789 11747 3847 11753
rect 3789 11744 3801 11747
rect 3568 11716 3801 11744
rect 3568 11704 3574 11716
rect 3789 11713 3801 11716
rect 3835 11713 3847 11747
rect 3789 11707 3847 11713
rect 3970 11704 3976 11756
rect 4028 11744 4034 11756
rect 4065 11747 4123 11753
rect 4065 11744 4077 11747
rect 4028 11716 4077 11744
rect 4028 11704 4034 11716
rect 4065 11713 4077 11716
rect 4111 11713 4123 11747
rect 4065 11707 4123 11713
rect 4154 11704 4160 11756
rect 4212 11704 4218 11756
rect 4433 11747 4491 11753
rect 4433 11713 4445 11747
rect 4479 11713 4491 11747
rect 4617 11747 4675 11753
rect 4617 11744 4629 11747
rect 4433 11707 4491 11713
rect 4540 11716 4629 11744
rect 4448 11676 4476 11707
rect 2700 11648 2912 11676
rect 2884 11617 2912 11648
rect 2976 11648 4476 11676
rect 2869 11611 2927 11617
rect 2869 11577 2881 11611
rect 2915 11577 2927 11611
rect 2869 11571 2927 11577
rect 2976 11552 3004 11648
rect 3878 11568 3884 11620
rect 3936 11608 3942 11620
rect 4540 11608 4568 11716
rect 4617 11713 4629 11716
rect 4663 11713 4675 11747
rect 4617 11707 4675 11713
rect 4706 11704 4712 11756
rect 4764 11704 4770 11756
rect 5537 11747 5595 11753
rect 5537 11744 5549 11747
rect 5276 11716 5549 11744
rect 3936 11580 4568 11608
rect 4724 11608 4752 11704
rect 5276 11620 5304 11716
rect 5537 11713 5549 11716
rect 5583 11713 5595 11747
rect 5537 11707 5595 11713
rect 5810 11704 5816 11756
rect 5868 11704 5874 11756
rect 6089 11747 6147 11753
rect 6089 11713 6101 11747
rect 6135 11713 6147 11747
rect 6089 11707 6147 11713
rect 6641 11747 6699 11753
rect 6641 11713 6653 11747
rect 6687 11744 6699 11747
rect 7098 11744 7104 11756
rect 6687 11716 7104 11744
rect 6687 11713 6699 11716
rect 6641 11707 6699 11713
rect 5626 11636 5632 11688
rect 5684 11676 5690 11688
rect 6104 11676 6132 11707
rect 7098 11704 7104 11716
rect 7156 11704 7162 11756
rect 7837 11747 7895 11753
rect 7837 11713 7849 11747
rect 7883 11744 7895 11747
rect 7926 11744 7932 11756
rect 7883 11716 7932 11744
rect 7883 11713 7895 11716
rect 7837 11707 7895 11713
rect 7926 11704 7932 11716
rect 7984 11704 7990 11756
rect 8386 11704 8392 11756
rect 8444 11744 8450 11756
rect 8444 11716 8892 11744
rect 8444 11704 8450 11716
rect 8864 11688 8892 11716
rect 9306 11704 9312 11756
rect 9364 11704 9370 11756
rect 9490 11704 9496 11756
rect 9548 11704 9554 11756
rect 11333 11747 11391 11753
rect 11333 11713 11345 11747
rect 11379 11744 11391 11747
rect 11422 11744 11428 11756
rect 11379 11716 11428 11744
rect 11379 11713 11391 11716
rect 11333 11707 11391 11713
rect 11422 11704 11428 11716
rect 11480 11744 11486 11756
rect 12066 11744 12072 11756
rect 11480 11716 12072 11744
rect 11480 11704 11486 11716
rect 12066 11704 12072 11716
rect 12124 11704 12130 11756
rect 13832 11753 13860 11852
rect 15102 11840 15108 11852
rect 15160 11840 15166 11892
rect 14826 11812 14832 11824
rect 14016 11784 14832 11812
rect 13817 11747 13875 11753
rect 13817 11713 13829 11747
rect 13863 11713 13875 11747
rect 13817 11707 13875 11713
rect 13906 11704 13912 11756
rect 13964 11744 13970 11756
rect 14016 11753 14044 11784
rect 14826 11772 14832 11784
rect 14884 11772 14890 11824
rect 14001 11747 14059 11753
rect 14001 11744 14013 11747
rect 13964 11716 14013 11744
rect 13964 11704 13970 11716
rect 14001 11713 14013 11716
rect 14047 11713 14059 11747
rect 14001 11707 14059 11713
rect 14090 11704 14096 11756
rect 14148 11704 14154 11756
rect 14366 11744 14372 11756
rect 14200 11716 14372 11744
rect 5684 11648 6132 11676
rect 5684 11636 5690 11648
rect 8846 11636 8852 11688
rect 8904 11676 8910 11688
rect 9508 11676 9536 11704
rect 8904 11648 9536 11676
rect 8904 11636 8910 11648
rect 5258 11608 5264 11620
rect 4724 11580 5264 11608
rect 3936 11568 3942 11580
rect 5258 11568 5264 11580
rect 5316 11568 5322 11620
rect 6825 11611 6883 11617
rect 6825 11577 6837 11611
rect 6871 11608 6883 11611
rect 7190 11608 7196 11620
rect 6871 11580 7196 11608
rect 6871 11577 6883 11580
rect 6825 11571 6883 11577
rect 7190 11568 7196 11580
rect 7248 11568 7254 11620
rect 7282 11568 7288 11620
rect 7340 11568 7346 11620
rect 13449 11611 13507 11617
rect 13449 11577 13461 11611
rect 13495 11608 13507 11611
rect 13998 11608 14004 11620
rect 13495 11580 14004 11608
rect 13495 11577 13507 11580
rect 13449 11571 13507 11577
rect 13998 11568 14004 11580
rect 14056 11568 14062 11620
rect 2958 11500 2964 11552
rect 3016 11500 3022 11552
rect 3050 11500 3056 11552
rect 3108 11540 3114 11552
rect 3418 11540 3424 11552
rect 3108 11512 3424 11540
rect 3108 11500 3114 11512
rect 3418 11500 3424 11512
rect 3476 11500 3482 11552
rect 3510 11500 3516 11552
rect 3568 11540 3574 11552
rect 4433 11543 4491 11549
rect 4433 11540 4445 11543
rect 3568 11512 4445 11540
rect 3568 11500 3574 11512
rect 4433 11509 4445 11512
rect 4479 11509 4491 11543
rect 4433 11503 4491 11509
rect 5169 11543 5227 11549
rect 5169 11509 5181 11543
rect 5215 11540 5227 11543
rect 5629 11543 5687 11549
rect 5629 11540 5641 11543
rect 5215 11512 5641 11540
rect 5215 11509 5227 11512
rect 5169 11503 5227 11509
rect 5629 11509 5641 11512
rect 5675 11509 5687 11543
rect 5629 11503 5687 11509
rect 6914 11500 6920 11552
rect 6972 11540 6978 11552
rect 7101 11543 7159 11549
rect 7101 11540 7113 11543
rect 6972 11512 7113 11540
rect 6972 11500 6978 11512
rect 7101 11509 7113 11512
rect 7147 11509 7159 11543
rect 7101 11503 7159 11509
rect 9214 11500 9220 11552
rect 9272 11540 9278 11552
rect 9950 11540 9956 11552
rect 9272 11512 9956 11540
rect 9272 11500 9278 11512
rect 9950 11500 9956 11512
rect 10008 11500 10014 11552
rect 14200 11540 14228 11716
rect 14366 11704 14372 11716
rect 14424 11704 14430 11756
rect 14553 11747 14611 11753
rect 14553 11713 14565 11747
rect 14599 11713 14611 11747
rect 14553 11707 14611 11713
rect 14274 11636 14280 11688
rect 14332 11676 14338 11688
rect 14568 11676 14596 11707
rect 14918 11704 14924 11756
rect 14976 11704 14982 11756
rect 15177 11747 15235 11753
rect 15177 11744 15189 11747
rect 15028 11716 15189 11744
rect 14332 11648 14596 11676
rect 14332 11636 14338 11648
rect 14826 11636 14832 11688
rect 14884 11676 14890 11688
rect 15028 11676 15056 11716
rect 15177 11713 15189 11716
rect 15223 11713 15235 11747
rect 15177 11707 15235 11713
rect 14884 11648 15056 11676
rect 14884 11636 14890 11648
rect 14277 11543 14335 11549
rect 14277 11540 14289 11543
rect 14200 11512 14289 11540
rect 14277 11509 14289 11512
rect 14323 11509 14335 11543
rect 14277 11503 14335 11509
rect 14366 11500 14372 11552
rect 14424 11540 14430 11552
rect 14737 11543 14795 11549
rect 14737 11540 14749 11543
rect 14424 11512 14749 11540
rect 14424 11500 14430 11512
rect 14737 11509 14749 11512
rect 14783 11509 14795 11543
rect 14737 11503 14795 11509
rect 15102 11500 15108 11552
rect 15160 11540 15166 11552
rect 16022 11540 16028 11552
rect 15160 11512 16028 11540
rect 15160 11500 15166 11512
rect 16022 11500 16028 11512
rect 16080 11540 16086 11552
rect 16301 11543 16359 11549
rect 16301 11540 16313 11543
rect 16080 11512 16313 11540
rect 16080 11500 16086 11512
rect 16301 11509 16313 11512
rect 16347 11509 16359 11543
rect 16301 11503 16359 11509
rect 1104 11450 16652 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 16652 11450
rect 1104 11376 16652 11398
rect 1762 11296 1768 11348
rect 1820 11336 1826 11348
rect 1820 11308 2452 11336
rect 1820 11296 1826 11308
rect 2424 11200 2452 11308
rect 2774 11296 2780 11348
rect 2832 11296 2838 11348
rect 2869 11339 2927 11345
rect 2869 11305 2881 11339
rect 2915 11336 2927 11339
rect 3142 11336 3148 11348
rect 2915 11308 3148 11336
rect 2915 11305 2927 11308
rect 2869 11299 2927 11305
rect 3142 11296 3148 11308
rect 3200 11296 3206 11348
rect 5258 11296 5264 11348
rect 5316 11296 5322 11348
rect 5445 11339 5503 11345
rect 5445 11305 5457 11339
rect 5491 11336 5503 11339
rect 5718 11336 5724 11348
rect 5491 11308 5724 11336
rect 5491 11305 5503 11308
rect 5445 11299 5503 11305
rect 5718 11296 5724 11308
rect 5776 11336 5782 11348
rect 6178 11336 6184 11348
rect 5776 11308 6184 11336
rect 5776 11296 5782 11308
rect 6178 11296 6184 11308
rect 6236 11296 6242 11348
rect 8570 11296 8576 11348
rect 8628 11336 8634 11348
rect 8628 11308 8708 11336
rect 8628 11296 8634 11308
rect 4433 11271 4491 11277
rect 4433 11237 4445 11271
rect 4479 11268 4491 11271
rect 4614 11268 4620 11280
rect 4479 11240 4620 11268
rect 4479 11237 4491 11240
rect 4433 11231 4491 11237
rect 4614 11228 4620 11240
rect 4672 11228 4678 11280
rect 4709 11203 4767 11209
rect 2424 11172 2912 11200
rect 1397 11135 1455 11141
rect 1397 11101 1409 11135
rect 1443 11132 1455 11135
rect 2774 11132 2780 11144
rect 1443 11104 2780 11132
rect 1443 11101 1455 11104
rect 1397 11095 1455 11101
rect 2774 11092 2780 11104
rect 2832 11092 2838 11144
rect 2884 11141 2912 11172
rect 4709 11169 4721 11203
rect 4755 11200 4767 11203
rect 6546 11200 6552 11212
rect 4755 11172 6552 11200
rect 4755 11169 4767 11172
rect 4709 11163 4767 11169
rect 6546 11160 6552 11172
rect 6604 11160 6610 11212
rect 8680 11200 8708 11308
rect 8938 11296 8944 11348
rect 8996 11296 9002 11348
rect 9122 11296 9128 11348
rect 9180 11336 9186 11348
rect 9769 11339 9827 11345
rect 9769 11336 9781 11339
rect 9180 11308 9781 11336
rect 9180 11296 9186 11308
rect 9769 11305 9781 11308
rect 9815 11305 9827 11339
rect 9769 11299 9827 11305
rect 9953 11339 10011 11345
rect 9953 11305 9965 11339
rect 9999 11336 10011 11339
rect 10502 11336 10508 11348
rect 9999 11308 10508 11336
rect 9999 11305 10011 11308
rect 9953 11299 10011 11305
rect 10502 11296 10508 11308
rect 10560 11296 10566 11348
rect 13262 11336 13268 11348
rect 10888 11308 13268 11336
rect 8757 11271 8815 11277
rect 8757 11237 8769 11271
rect 8803 11268 8815 11271
rect 9674 11268 9680 11280
rect 8803 11240 9680 11268
rect 8803 11237 8815 11240
rect 8757 11231 8815 11237
rect 9674 11228 9680 11240
rect 9732 11228 9738 11280
rect 9335 11203 9393 11209
rect 8680 11172 9168 11200
rect 2869 11135 2927 11141
rect 2869 11101 2881 11135
rect 2915 11101 2927 11135
rect 2869 11095 2927 11101
rect 3053 11135 3111 11141
rect 3053 11101 3065 11135
rect 3099 11101 3111 11135
rect 3053 11095 3111 11101
rect 1670 11073 1676 11076
rect 1664 11027 1676 11073
rect 1670 11024 1676 11027
rect 1728 11024 1734 11076
rect 2222 11024 2228 11076
rect 2280 11064 2286 11076
rect 3068 11064 3096 11095
rect 4154 11092 4160 11144
rect 4212 11132 4218 11144
rect 4341 11135 4399 11141
rect 4341 11132 4353 11135
rect 4212 11104 4353 11132
rect 4212 11092 4218 11104
rect 4341 11101 4353 11104
rect 4387 11101 4399 11135
rect 4341 11095 4399 11101
rect 4522 11092 4528 11144
rect 4580 11092 4586 11144
rect 4617 11135 4675 11141
rect 4617 11101 4629 11135
rect 4663 11101 4675 11135
rect 4617 11095 4675 11101
rect 4801 11135 4859 11141
rect 4801 11101 4813 11135
rect 4847 11132 4859 11135
rect 4890 11132 4896 11144
rect 4847 11104 4896 11132
rect 4847 11101 4859 11104
rect 4801 11095 4859 11101
rect 2280 11036 3096 11064
rect 2280 11024 2286 11036
rect 3142 11024 3148 11076
rect 3200 11064 3206 11076
rect 3786 11064 3792 11076
rect 3200 11036 3792 11064
rect 3200 11024 3206 11036
rect 3786 11024 3792 11036
rect 3844 11024 3850 11076
rect 4632 11064 4660 11095
rect 4890 11092 4896 11104
rect 4948 11132 4954 11144
rect 5718 11132 5724 11144
rect 4948 11104 5724 11132
rect 4948 11092 4954 11104
rect 5718 11092 5724 11104
rect 5776 11092 5782 11144
rect 9140 11141 9168 11172
rect 9335 11169 9347 11203
rect 9381 11200 9393 11203
rect 10888 11200 10916 11308
rect 13262 11296 13268 11308
rect 13320 11296 13326 11348
rect 13357 11339 13415 11345
rect 13357 11305 13369 11339
rect 13403 11336 13415 11339
rect 13446 11336 13452 11348
rect 13403 11308 13452 11336
rect 13403 11305 13415 11308
rect 13357 11299 13415 11305
rect 13446 11296 13452 11308
rect 13504 11296 13510 11348
rect 14182 11296 14188 11348
rect 14240 11336 14246 11348
rect 14550 11336 14556 11348
rect 14240 11308 14556 11336
rect 14240 11296 14246 11308
rect 14550 11296 14556 11308
rect 14608 11296 14614 11348
rect 14826 11296 14832 11348
rect 14884 11296 14890 11348
rect 16206 11336 16212 11348
rect 14936 11308 16212 11336
rect 14936 11268 14964 11308
rect 16206 11296 16212 11308
rect 16264 11296 16270 11348
rect 14384 11240 14964 11268
rect 13906 11200 13912 11212
rect 9381 11172 10916 11200
rect 13280 11172 13912 11200
rect 9381 11169 9393 11172
rect 9335 11163 9393 11169
rect 9125 11135 9183 11141
rect 9125 11101 9137 11135
rect 9171 11132 9183 11135
rect 9214 11132 9220 11144
rect 9171 11104 9220 11132
rect 9171 11101 9183 11104
rect 9125 11095 9183 11101
rect 9214 11092 9220 11104
rect 9272 11092 9278 11144
rect 9490 11092 9496 11144
rect 9548 11092 9554 11144
rect 10226 11092 10232 11144
rect 10284 11132 10290 11144
rect 11698 11132 11704 11144
rect 10284 11104 11704 11132
rect 10284 11092 10290 11104
rect 11698 11092 11704 11104
rect 11756 11092 11762 11144
rect 13280 11141 13308 11172
rect 13906 11160 13912 11172
rect 13964 11160 13970 11212
rect 13265 11135 13323 11141
rect 13265 11101 13277 11135
rect 13311 11101 13323 11135
rect 13265 11095 13323 11101
rect 13449 11135 13507 11141
rect 13449 11101 13461 11135
rect 13495 11132 13507 11135
rect 13725 11135 13783 11141
rect 13725 11132 13737 11135
rect 13495 11104 13737 11132
rect 13495 11101 13507 11104
rect 13449 11095 13507 11101
rect 13725 11101 13737 11104
rect 13771 11132 13783 11135
rect 13814 11132 13820 11144
rect 13771 11104 13820 11132
rect 13771 11101 13783 11104
rect 13725 11095 13783 11101
rect 13814 11092 13820 11104
rect 13872 11092 13878 11144
rect 14384 11141 14412 11240
rect 15930 11228 15936 11280
rect 15988 11268 15994 11280
rect 16301 11271 16359 11277
rect 16301 11268 16313 11271
rect 15988 11240 16313 11268
rect 15988 11228 15994 11240
rect 16301 11237 16313 11240
rect 16347 11237 16359 11271
rect 16301 11231 16359 11237
rect 14918 11160 14924 11212
rect 14976 11160 14982 11212
rect 14185 11135 14243 11141
rect 14185 11101 14197 11135
rect 14231 11101 14243 11135
rect 14185 11095 14243 11101
rect 14369 11135 14427 11141
rect 14369 11101 14381 11135
rect 14415 11101 14427 11135
rect 14369 11095 14427 11101
rect 4706 11064 4712 11076
rect 4632 11036 4712 11064
rect 4706 11024 4712 11036
rect 4764 11064 4770 11076
rect 5429 11067 5487 11073
rect 5429 11064 5441 11067
rect 4764 11036 5441 11064
rect 4764 11024 4770 11036
rect 5429 11033 5441 11036
rect 5475 11064 5487 11067
rect 5534 11064 5540 11076
rect 5475 11036 5540 11064
rect 5475 11033 5487 11036
rect 5429 11027 5487 11033
rect 5534 11024 5540 11036
rect 5592 11024 5598 11076
rect 5629 11067 5687 11073
rect 5629 11033 5641 11067
rect 5675 11064 5687 11067
rect 5810 11064 5816 11076
rect 5675 11036 5816 11064
rect 5675 11033 5687 11036
rect 5629 11027 5687 11033
rect 5810 11024 5816 11036
rect 5868 11024 5874 11076
rect 8389 11067 8447 11073
rect 8389 11033 8401 11067
rect 8435 11064 8447 11067
rect 8846 11064 8852 11076
rect 8435 11036 8852 11064
rect 8435 11033 8447 11036
rect 8389 11027 8447 11033
rect 8846 11024 8852 11036
rect 8904 11024 8910 11076
rect 9030 11024 9036 11076
rect 9088 11064 9094 11076
rect 9585 11067 9643 11073
rect 9088 11036 9536 11064
rect 9088 11024 9094 11036
rect 2038 10956 2044 11008
rect 2096 10996 2102 11008
rect 2590 10996 2596 11008
rect 2096 10968 2596 10996
rect 2096 10956 2102 10968
rect 2590 10956 2596 10968
rect 2648 10956 2654 11008
rect 4798 10956 4804 11008
rect 4856 10996 4862 11008
rect 5074 10996 5080 11008
rect 4856 10968 5080 10996
rect 4856 10956 4862 10968
rect 5074 10956 5080 10968
rect 5132 10996 5138 11008
rect 8110 10996 8116 11008
rect 5132 10968 8116 10996
rect 5132 10956 5138 10968
rect 8110 10956 8116 10968
rect 8168 10956 8174 11008
rect 8599 10999 8657 11005
rect 8599 10965 8611 10999
rect 8645 10996 8657 10999
rect 8754 10996 8760 11008
rect 8645 10968 8760 10996
rect 8645 10965 8657 10968
rect 8599 10959 8657 10965
rect 8754 10956 8760 10968
rect 8812 10996 8818 11008
rect 9122 10996 9128 11008
rect 8812 10968 9128 10996
rect 8812 10956 8818 10968
rect 9122 10956 9128 10968
rect 9180 10956 9186 11008
rect 9508 10996 9536 11036
rect 9585 11033 9597 11067
rect 9631 11064 9643 11067
rect 9631 11036 11652 11064
rect 9631 11033 9643 11036
rect 9585 11027 9643 11033
rect 9785 10999 9843 11005
rect 9785 10996 9797 10999
rect 9508 10968 9797 10996
rect 9785 10965 9797 10968
rect 9831 10965 9843 10999
rect 11624 10996 11652 11036
rect 12066 11024 12072 11076
rect 12124 11064 12130 11076
rect 12437 11067 12495 11073
rect 12437 11064 12449 11067
rect 12124 11036 12449 11064
rect 12124 11024 12130 11036
rect 12437 11033 12449 11036
rect 12483 11033 12495 11067
rect 12437 11027 12495 11033
rect 13541 11067 13599 11073
rect 13541 11033 13553 11067
rect 13587 11064 13599 11067
rect 13906 11064 13912 11076
rect 13587 11036 13912 11064
rect 13587 11033 13599 11036
rect 13541 11027 13599 11033
rect 13906 11024 13912 11036
rect 13964 11024 13970 11076
rect 12710 10996 12716 11008
rect 11624 10968 12716 10996
rect 9785 10959 9843 10965
rect 12710 10956 12716 10968
rect 12768 10996 12774 11008
rect 14090 10996 14096 11008
rect 12768 10968 14096 10996
rect 12768 10956 12774 10968
rect 14090 10956 14096 10968
rect 14148 10996 14154 11008
rect 14200 10996 14228 11095
rect 14458 11092 14464 11144
rect 14516 11092 14522 11144
rect 14550 11092 14556 11144
rect 14608 11092 14614 11144
rect 15194 11141 15200 11144
rect 15188 11132 15200 11141
rect 15155 11104 15200 11132
rect 15188 11095 15200 11104
rect 15194 11092 15200 11095
rect 15252 11092 15258 11144
rect 14274 11024 14280 11076
rect 14332 11064 14338 11076
rect 15286 11064 15292 11076
rect 14332 11036 15292 11064
rect 14332 11024 14338 11036
rect 15286 11024 15292 11036
rect 15344 11024 15350 11076
rect 15746 10996 15752 11008
rect 14148 10968 15752 10996
rect 14148 10956 14154 10968
rect 15746 10956 15752 10968
rect 15804 10956 15810 11008
rect 1104 10906 16652 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 16652 10906
rect 1104 10832 16652 10854
rect 1670 10752 1676 10804
rect 1728 10752 1734 10804
rect 3234 10792 3240 10804
rect 2240 10764 3240 10792
rect 1841 10727 1899 10733
rect 1841 10693 1853 10727
rect 1887 10724 1899 10727
rect 1887 10696 1992 10724
rect 1887 10693 1899 10696
rect 1841 10687 1899 10693
rect 1964 10588 1992 10696
rect 2038 10684 2044 10736
rect 2096 10684 2102 10736
rect 2240 10665 2268 10764
rect 3234 10752 3240 10764
rect 3292 10752 3298 10804
rect 7190 10752 7196 10804
rect 7248 10792 7254 10804
rect 7469 10795 7527 10801
rect 7469 10792 7481 10795
rect 7248 10764 7481 10792
rect 7248 10752 7254 10764
rect 7469 10761 7481 10764
rect 7515 10761 7527 10795
rect 7469 10755 7527 10761
rect 13630 10752 13636 10804
rect 13688 10752 13694 10804
rect 15010 10792 15016 10804
rect 13832 10764 15016 10792
rect 2409 10727 2467 10733
rect 2409 10693 2421 10727
rect 2455 10724 2467 10727
rect 2590 10724 2596 10736
rect 2455 10696 2596 10724
rect 2455 10693 2467 10696
rect 2409 10687 2467 10693
rect 2590 10684 2596 10696
rect 2648 10684 2654 10736
rect 5718 10684 5724 10736
rect 5776 10684 5782 10736
rect 7653 10727 7711 10733
rect 7653 10693 7665 10727
rect 7699 10724 7711 10727
rect 8662 10724 8668 10736
rect 7699 10696 8668 10724
rect 7699 10693 7711 10696
rect 7653 10687 7711 10693
rect 8662 10684 8668 10696
rect 8720 10684 8726 10736
rect 9125 10727 9183 10733
rect 9125 10693 9137 10727
rect 9171 10724 9183 10727
rect 9171 10696 9720 10724
rect 9171 10693 9183 10696
rect 9125 10687 9183 10693
rect 2225 10659 2283 10665
rect 2225 10625 2237 10659
rect 2271 10625 2283 10659
rect 2225 10619 2283 10625
rect 2314 10616 2320 10668
rect 2372 10656 2378 10668
rect 2501 10659 2559 10665
rect 2501 10656 2513 10659
rect 2372 10628 2513 10656
rect 2372 10616 2378 10628
rect 2501 10625 2513 10628
rect 2547 10625 2559 10659
rect 2501 10619 2559 10625
rect 2685 10659 2743 10665
rect 2685 10625 2697 10659
rect 2731 10656 2743 10659
rect 3510 10656 3516 10668
rect 2731 10628 3516 10656
rect 2731 10625 2743 10628
rect 2685 10619 2743 10625
rect 3510 10616 3516 10628
rect 3568 10616 3574 10668
rect 4062 10616 4068 10668
rect 4120 10616 4126 10668
rect 4706 10616 4712 10668
rect 4764 10616 4770 10668
rect 4982 10616 4988 10668
rect 5040 10616 5046 10668
rect 5353 10659 5411 10665
rect 5353 10625 5365 10659
rect 5399 10625 5411 10659
rect 5353 10619 5411 10625
rect 5537 10659 5595 10665
rect 5537 10625 5549 10659
rect 5583 10656 5595 10659
rect 5626 10656 5632 10668
rect 5583 10628 5632 10656
rect 5583 10625 5595 10628
rect 5537 10619 5595 10625
rect 2593 10591 2651 10597
rect 2593 10588 2605 10591
rect 1964 10560 2605 10588
rect 2593 10557 2605 10560
rect 2639 10557 2651 10591
rect 5000 10588 5028 10616
rect 5258 10588 5264 10600
rect 5000 10560 5264 10588
rect 2593 10551 2651 10557
rect 5258 10548 5264 10560
rect 5316 10548 5322 10600
rect 3418 10480 3424 10532
rect 3476 10520 3482 10532
rect 4065 10523 4123 10529
rect 4065 10520 4077 10523
rect 3476 10492 4077 10520
rect 3476 10480 3482 10492
rect 4065 10489 4077 10492
rect 4111 10489 4123 10523
rect 4065 10483 4123 10489
rect 4522 10480 4528 10532
rect 4580 10520 4586 10532
rect 4798 10520 4804 10532
rect 4580 10492 4804 10520
rect 4580 10480 4586 10492
rect 4798 10480 4804 10492
rect 4856 10520 4862 10532
rect 5368 10520 5396 10619
rect 5626 10616 5632 10628
rect 5684 10616 5690 10668
rect 7374 10616 7380 10668
rect 7432 10616 7438 10668
rect 8297 10659 8355 10665
rect 8297 10625 8309 10659
rect 8343 10625 8355 10659
rect 8297 10619 8355 10625
rect 8481 10659 8539 10665
rect 8481 10625 8493 10659
rect 8527 10656 8539 10659
rect 9030 10656 9036 10668
rect 8527 10628 9036 10656
rect 8527 10625 8539 10628
rect 8481 10619 8539 10625
rect 8312 10588 8340 10619
rect 9030 10616 9036 10628
rect 9088 10616 9094 10668
rect 9692 10665 9720 10696
rect 9309 10659 9367 10665
rect 9309 10625 9321 10659
rect 9355 10656 9367 10659
rect 9677 10659 9735 10665
rect 9355 10628 9628 10656
rect 9355 10625 9367 10628
rect 9309 10619 9367 10625
rect 8570 10588 8576 10600
rect 8312 10560 8576 10588
rect 8570 10548 8576 10560
rect 8628 10548 8634 10600
rect 8846 10548 8852 10600
rect 8904 10588 8910 10600
rect 9401 10591 9459 10597
rect 9401 10588 9413 10591
rect 8904 10560 9413 10588
rect 8904 10548 8910 10560
rect 9401 10557 9413 10560
rect 9447 10557 9459 10591
rect 9600 10588 9628 10628
rect 9677 10625 9689 10659
rect 9723 10656 9735 10659
rect 9766 10656 9772 10668
rect 9723 10628 9772 10656
rect 9723 10625 9735 10628
rect 9677 10619 9735 10625
rect 9766 10616 9772 10628
rect 9824 10616 9830 10668
rect 12066 10616 12072 10668
rect 12124 10616 12130 10668
rect 13832 10665 13860 10764
rect 15010 10752 15016 10764
rect 15068 10752 15074 10804
rect 15286 10752 15292 10804
rect 15344 10792 15350 10804
rect 15838 10792 15844 10804
rect 15344 10764 15844 10792
rect 15344 10752 15350 10764
rect 15838 10752 15844 10764
rect 15896 10792 15902 10804
rect 16301 10795 16359 10801
rect 16301 10792 16313 10795
rect 15896 10764 16313 10792
rect 15896 10752 15902 10764
rect 16301 10761 16313 10764
rect 16347 10761 16359 10795
rect 16301 10755 16359 10761
rect 14829 10727 14887 10733
rect 14829 10693 14841 10727
rect 14875 10724 14887 10727
rect 15166 10727 15224 10733
rect 15166 10724 15178 10727
rect 14875 10696 15178 10724
rect 14875 10693 14887 10696
rect 14829 10687 14887 10693
rect 15166 10693 15178 10696
rect 15212 10693 15224 10727
rect 15166 10687 15224 10693
rect 13449 10659 13507 10665
rect 13449 10625 13461 10659
rect 13495 10625 13507 10659
rect 13449 10619 13507 10625
rect 13817 10659 13875 10665
rect 13817 10625 13829 10659
rect 13863 10625 13875 10659
rect 13817 10619 13875 10625
rect 10502 10588 10508 10600
rect 9600 10560 10508 10588
rect 9401 10551 9459 10557
rect 10502 10548 10508 10560
rect 10560 10548 10566 10600
rect 13464 10588 13492 10619
rect 14090 10616 14096 10668
rect 14148 10656 14154 10668
rect 14185 10659 14243 10665
rect 14185 10656 14197 10659
rect 14148 10628 14197 10656
rect 14148 10616 14154 10628
rect 14185 10625 14197 10628
rect 14231 10625 14243 10659
rect 14185 10619 14243 10625
rect 14366 10616 14372 10668
rect 14424 10616 14430 10668
rect 14458 10616 14464 10668
rect 14516 10616 14522 10668
rect 14553 10659 14611 10665
rect 14553 10625 14565 10659
rect 14599 10656 14611 10659
rect 15470 10656 15476 10668
rect 14599 10628 15476 10656
rect 14599 10625 14611 10628
rect 14553 10619 14611 10625
rect 15470 10616 15476 10628
rect 15528 10616 15534 10668
rect 14826 10588 14832 10600
rect 13464 10560 14832 10588
rect 14826 10548 14832 10560
rect 14884 10548 14890 10600
rect 14918 10548 14924 10600
rect 14976 10548 14982 10600
rect 4856 10492 5396 10520
rect 4856 10480 4862 10492
rect 8202 10480 8208 10532
rect 8260 10520 8266 10532
rect 9493 10523 9551 10529
rect 9493 10520 9505 10523
rect 8260 10492 9505 10520
rect 8260 10480 8266 10492
rect 9493 10489 9505 10492
rect 9539 10489 9551 10523
rect 9493 10483 9551 10489
rect 13265 10523 13323 10529
rect 13265 10489 13277 10523
rect 13311 10520 13323 10523
rect 13311 10492 14964 10520
rect 13311 10489 13323 10492
rect 13265 10483 13323 10489
rect 1854 10412 1860 10464
rect 1912 10412 1918 10464
rect 5902 10412 5908 10464
rect 5960 10412 5966 10464
rect 7650 10412 7656 10464
rect 7708 10412 7714 10464
rect 8478 10412 8484 10464
rect 8536 10412 8542 10464
rect 8941 10455 8999 10461
rect 8941 10421 8953 10455
rect 8987 10452 8999 10455
rect 9122 10452 9128 10464
rect 8987 10424 9128 10452
rect 8987 10421 8999 10424
rect 8941 10415 8999 10421
rect 9122 10412 9128 10424
rect 9180 10412 9186 10464
rect 9585 10455 9643 10461
rect 9585 10421 9597 10455
rect 9631 10452 9643 10455
rect 10962 10452 10968 10464
rect 9631 10424 10968 10452
rect 9631 10421 9643 10424
rect 9585 10415 9643 10421
rect 10962 10412 10968 10424
rect 11020 10412 11026 10464
rect 13909 10455 13967 10461
rect 13909 10421 13921 10455
rect 13955 10452 13967 10455
rect 13998 10452 14004 10464
rect 13955 10424 14004 10452
rect 13955 10421 13967 10424
rect 13909 10415 13967 10421
rect 13998 10412 14004 10424
rect 14056 10412 14062 10464
rect 14936 10452 14964 10492
rect 15194 10452 15200 10464
rect 14936 10424 15200 10452
rect 15194 10412 15200 10424
rect 15252 10412 15258 10464
rect 1104 10362 16652 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 16652 10362
rect 1104 10288 16652 10310
rect 3145 10251 3203 10257
rect 3145 10217 3157 10251
rect 3191 10248 3203 10251
rect 3234 10248 3240 10260
rect 3191 10220 3240 10248
rect 3191 10217 3203 10220
rect 3145 10211 3203 10217
rect 3234 10208 3240 10220
rect 3292 10208 3298 10260
rect 5261 10251 5319 10257
rect 5261 10217 5273 10251
rect 5307 10248 5319 10251
rect 5718 10248 5724 10260
rect 5307 10220 5724 10248
rect 5307 10217 5319 10220
rect 5261 10211 5319 10217
rect 5718 10208 5724 10220
rect 5776 10208 5782 10260
rect 7101 10251 7159 10257
rect 7101 10217 7113 10251
rect 7147 10248 7159 10251
rect 7190 10248 7196 10260
rect 7147 10220 7196 10248
rect 7147 10217 7159 10220
rect 7101 10211 7159 10217
rect 7190 10208 7196 10220
rect 7248 10208 7254 10260
rect 7285 10251 7343 10257
rect 7285 10217 7297 10251
rect 7331 10248 7343 10251
rect 7926 10248 7932 10260
rect 7331 10220 7932 10248
rect 7331 10217 7343 10220
rect 7285 10211 7343 10217
rect 7926 10208 7932 10220
rect 7984 10208 7990 10260
rect 8021 10251 8079 10257
rect 8021 10217 8033 10251
rect 8067 10248 8079 10251
rect 8662 10248 8668 10260
rect 8067 10220 8668 10248
rect 8067 10217 8079 10220
rect 8021 10211 8079 10217
rect 8662 10208 8668 10220
rect 8720 10208 8726 10260
rect 8754 10208 8760 10260
rect 8812 10208 8818 10260
rect 12989 10251 13047 10257
rect 12989 10217 13001 10251
rect 13035 10248 13047 10251
rect 15286 10248 15292 10260
rect 13035 10220 15292 10248
rect 13035 10217 13047 10220
rect 12989 10211 13047 10217
rect 15286 10208 15292 10220
rect 15344 10208 15350 10260
rect 16209 10251 16267 10257
rect 16209 10217 16221 10251
rect 16255 10248 16267 10251
rect 16298 10248 16304 10260
rect 16255 10220 16304 10248
rect 16255 10217 16267 10220
rect 16209 10211 16267 10217
rect 16298 10208 16304 10220
rect 16356 10208 16362 10260
rect 8110 10140 8116 10192
rect 8168 10140 8174 10192
rect 8941 10183 8999 10189
rect 8941 10180 8953 10183
rect 8404 10152 8953 10180
rect 2774 10072 2780 10124
rect 2832 10112 2838 10124
rect 3970 10112 3976 10124
rect 2832 10084 3976 10112
rect 2832 10072 2838 10084
rect 3970 10072 3976 10084
rect 4028 10112 4034 10124
rect 4341 10115 4399 10121
rect 4341 10112 4353 10115
rect 4028 10084 4353 10112
rect 4028 10072 4034 10084
rect 4341 10081 4353 10084
rect 4387 10081 4399 10115
rect 4341 10075 4399 10081
rect 3326 10004 3332 10056
rect 3384 10004 3390 10056
rect 3602 10004 3608 10056
rect 3660 10004 3666 10056
rect 4706 10044 4712 10056
rect 3896 10016 4712 10044
rect 3513 9979 3571 9985
rect 3513 9945 3525 9979
rect 3559 9976 3571 9979
rect 3896 9976 3924 10016
rect 4706 10004 4712 10016
rect 4764 10004 4770 10056
rect 5169 10047 5227 10053
rect 5169 10013 5181 10047
rect 5215 10044 5227 10047
rect 5442 10044 5448 10056
rect 5215 10016 5448 10044
rect 5215 10013 5227 10016
rect 5169 10007 5227 10013
rect 5442 10004 5448 10016
rect 5500 10004 5506 10056
rect 6638 10004 6644 10056
rect 6696 10004 6702 10056
rect 6733 10047 6791 10053
rect 6733 10013 6745 10047
rect 6779 10044 6791 10047
rect 6914 10044 6920 10056
rect 6779 10016 6920 10044
rect 6779 10013 6791 10016
rect 6733 10007 6791 10013
rect 6914 10004 6920 10016
rect 6972 10044 6978 10056
rect 7377 10047 7435 10053
rect 7377 10044 7389 10047
rect 6972 10016 7389 10044
rect 6972 10004 6978 10016
rect 7377 10013 7389 10016
rect 7423 10013 7435 10047
rect 7377 10007 7435 10013
rect 8113 10047 8171 10053
rect 8113 10013 8125 10047
rect 8159 10044 8171 10047
rect 8294 10044 8300 10056
rect 8159 10016 8300 10044
rect 8159 10013 8171 10016
rect 8113 10007 8171 10013
rect 8294 10004 8300 10016
rect 8352 10004 8358 10056
rect 8404 10053 8432 10152
rect 8941 10149 8953 10152
rect 8987 10149 8999 10183
rect 14090 10180 14096 10192
rect 8941 10143 8999 10149
rect 13648 10152 14096 10180
rect 8478 10072 8484 10124
rect 8536 10112 8542 10124
rect 9493 10115 9551 10121
rect 9493 10112 9505 10115
rect 8536 10084 9505 10112
rect 8536 10072 8542 10084
rect 9493 10081 9505 10084
rect 9539 10081 9551 10115
rect 9493 10075 9551 10081
rect 12894 10072 12900 10124
rect 12952 10112 12958 10124
rect 12952 10084 13584 10112
rect 12952 10072 12958 10084
rect 8389 10047 8447 10053
rect 8389 10013 8401 10047
rect 8435 10013 8447 10047
rect 8389 10007 8447 10013
rect 8570 10004 8576 10056
rect 8628 10004 8634 10056
rect 8757 10047 8815 10053
rect 8757 10044 8769 10047
rect 8680 10016 8769 10044
rect 3559 9948 3924 9976
rect 3973 9979 4031 9985
rect 3559 9945 3571 9948
rect 3513 9939 3571 9945
rect 3973 9945 3985 9979
rect 4019 9976 4031 9979
rect 4890 9976 4896 9988
rect 4019 9948 4896 9976
rect 4019 9945 4031 9948
rect 3973 9939 4031 9945
rect 4890 9936 4896 9948
rect 4948 9936 4954 9988
rect 6362 9936 6368 9988
rect 6420 9985 6426 9988
rect 6420 9939 6432 9985
rect 7101 9979 7159 9985
rect 7101 9945 7113 9979
rect 7147 9976 7159 9979
rect 7147 9948 7420 9976
rect 7147 9945 7159 9948
rect 7101 9939 7159 9945
rect 6420 9936 6426 9939
rect 7392 9920 7420 9948
rect 4065 9911 4123 9917
rect 4065 9877 4077 9911
rect 4111 9908 4123 9911
rect 4522 9908 4528 9920
rect 4111 9880 4528 9908
rect 4111 9877 4123 9880
rect 4065 9871 4123 9877
rect 4522 9868 4528 9880
rect 4580 9908 4586 9920
rect 6454 9908 6460 9920
rect 4580 9880 6460 9908
rect 4580 9868 4586 9880
rect 6454 9868 6460 9880
rect 6512 9868 6518 9920
rect 7374 9868 7380 9920
rect 7432 9868 7438 9920
rect 8297 9911 8355 9917
rect 8297 9877 8309 9911
rect 8343 9908 8355 9911
rect 8680 9908 8708 10016
rect 8757 10013 8769 10016
rect 8803 10044 8815 10047
rect 9122 10044 9128 10056
rect 8803 10016 9128 10044
rect 8803 10013 8815 10016
rect 8757 10007 8815 10013
rect 9122 10004 9128 10016
rect 9180 10004 9186 10056
rect 10502 10004 10508 10056
rect 10560 10004 10566 10056
rect 11149 10047 11207 10053
rect 11149 10013 11161 10047
rect 11195 10044 11207 10047
rect 11195 10016 12112 10044
rect 11195 10013 11207 10016
rect 11149 10007 11207 10013
rect 11532 9988 11560 10016
rect 12084 9988 12112 10016
rect 13170 10004 13176 10056
rect 13228 10004 13234 10056
rect 13556 10053 13584 10084
rect 13648 10053 13676 10152
rect 14090 10140 14096 10152
rect 14148 10140 14154 10192
rect 13740 10084 14228 10112
rect 13740 10053 13768 10084
rect 13541 10047 13599 10053
rect 13541 10013 13553 10047
rect 13587 10013 13599 10047
rect 13541 10007 13599 10013
rect 13633 10047 13691 10053
rect 13633 10013 13645 10047
rect 13679 10013 13691 10047
rect 13633 10007 13691 10013
rect 13725 10047 13783 10053
rect 13725 10013 13737 10047
rect 13771 10013 13783 10047
rect 13725 10007 13783 10013
rect 13909 10047 13967 10053
rect 13909 10013 13921 10047
rect 13955 10044 13967 10047
rect 13998 10044 14004 10056
rect 13955 10016 14004 10044
rect 13955 10013 13967 10016
rect 13909 10007 13967 10013
rect 13998 10004 14004 10016
rect 14056 10004 14062 10056
rect 14093 10047 14151 10053
rect 14093 10013 14105 10047
rect 14139 10013 14151 10047
rect 14200 10044 14228 10084
rect 15565 10047 15623 10053
rect 15565 10044 15577 10047
rect 14200 10016 15577 10044
rect 14093 10007 14151 10013
rect 15565 10013 15577 10016
rect 15611 10013 15623 10047
rect 15565 10007 15623 10013
rect 16025 10047 16083 10053
rect 16025 10013 16037 10047
rect 16071 10044 16083 10047
rect 16114 10044 16120 10056
rect 16071 10016 16120 10044
rect 16071 10013 16083 10016
rect 16025 10007 16083 10013
rect 11422 9985 11428 9988
rect 11416 9939 11428 9985
rect 11422 9936 11428 9939
rect 11480 9936 11486 9988
rect 11514 9936 11520 9988
rect 11572 9936 11578 9988
rect 12066 9936 12072 9988
rect 12124 9976 12130 9988
rect 13078 9976 13084 9988
rect 12124 9948 13084 9976
rect 12124 9936 12130 9948
rect 13078 9936 13084 9948
rect 13136 9976 13142 9988
rect 14108 9976 14136 10007
rect 16114 10004 16120 10016
rect 16172 10004 16178 10056
rect 14338 9979 14396 9985
rect 14338 9976 14350 9979
rect 13136 9948 14136 9976
rect 14200 9948 14350 9976
rect 13136 9936 13142 9948
rect 8343 9880 8708 9908
rect 8343 9877 8355 9880
rect 8297 9871 8355 9877
rect 8754 9868 8760 9920
rect 8812 9908 8818 9920
rect 9861 9911 9919 9917
rect 9861 9908 9873 9911
rect 8812 9880 9873 9908
rect 8812 9868 8818 9880
rect 9861 9877 9873 9880
rect 9907 9877 9919 9911
rect 9861 9871 9919 9877
rect 12434 9868 12440 9920
rect 12492 9908 12498 9920
rect 12529 9911 12587 9917
rect 12529 9908 12541 9911
rect 12492 9880 12541 9908
rect 12492 9868 12498 9880
rect 12529 9877 12541 9880
rect 12575 9877 12587 9911
rect 12529 9871 12587 9877
rect 13265 9911 13323 9917
rect 13265 9877 13277 9911
rect 13311 9908 13323 9911
rect 14200 9908 14228 9948
rect 14338 9945 14350 9948
rect 14384 9945 14396 9979
rect 15749 9979 15807 9985
rect 15749 9976 15761 9979
rect 14338 9939 14396 9945
rect 15488 9948 15761 9976
rect 13311 9880 14228 9908
rect 13311 9877 13323 9880
rect 13265 9871 13323 9877
rect 14826 9868 14832 9920
rect 14884 9908 14890 9920
rect 15488 9917 15516 9948
rect 15749 9945 15761 9948
rect 15795 9945 15807 9979
rect 15749 9939 15807 9945
rect 15933 9979 15991 9985
rect 15933 9945 15945 9979
rect 15979 9945 15991 9979
rect 15933 9939 15991 9945
rect 15473 9911 15531 9917
rect 15473 9908 15485 9911
rect 14884 9880 15485 9908
rect 14884 9868 14890 9880
rect 15473 9877 15485 9880
rect 15519 9877 15531 9911
rect 15473 9871 15531 9877
rect 15562 9868 15568 9920
rect 15620 9908 15626 9920
rect 15948 9908 15976 9939
rect 16114 9908 16120 9920
rect 15620 9880 16120 9908
rect 15620 9868 15626 9880
rect 16114 9868 16120 9880
rect 16172 9868 16178 9920
rect 1104 9818 16652 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 16652 9818
rect 1104 9744 16652 9766
rect 3053 9707 3111 9713
rect 3053 9673 3065 9707
rect 3099 9704 3111 9707
rect 3326 9704 3332 9716
rect 3099 9676 3332 9704
rect 3099 9673 3111 9676
rect 3053 9667 3111 9673
rect 3326 9664 3332 9676
rect 3384 9664 3390 9716
rect 3697 9707 3755 9713
rect 3697 9673 3709 9707
rect 3743 9704 3755 9707
rect 4157 9707 4215 9713
rect 4157 9704 4169 9707
rect 3743 9676 4169 9704
rect 3743 9673 3755 9676
rect 3697 9667 3755 9673
rect 4157 9673 4169 9676
rect 4203 9673 4215 9707
rect 4157 9667 4215 9673
rect 4433 9707 4491 9713
rect 4433 9673 4445 9707
rect 4479 9704 4491 9707
rect 4706 9704 4712 9716
rect 4479 9676 4712 9704
rect 4479 9673 4491 9676
rect 4433 9667 4491 9673
rect 4706 9664 4712 9676
rect 4764 9664 4770 9716
rect 6362 9664 6368 9716
rect 6420 9664 6426 9716
rect 6914 9664 6920 9716
rect 6972 9664 6978 9716
rect 8570 9664 8576 9716
rect 8628 9704 8634 9716
rect 9030 9704 9036 9716
rect 8628 9676 9036 9704
rect 8628 9664 8634 9676
rect 9030 9664 9036 9676
rect 9088 9664 9094 9716
rect 12894 9664 12900 9716
rect 12952 9664 12958 9716
rect 14550 9704 14556 9716
rect 13740 9676 14556 9704
rect 3878 9636 3884 9648
rect 2884 9608 3884 9636
rect 2884 9577 2912 9608
rect 3878 9596 3884 9608
rect 3936 9636 3942 9648
rect 4065 9639 4123 9645
rect 4065 9636 4077 9639
rect 3936 9608 4077 9636
rect 3936 9596 3942 9608
rect 4065 9605 4077 9608
rect 4111 9605 4123 9639
rect 4065 9599 4123 9605
rect 4274 9639 4332 9645
rect 4274 9605 4286 9639
rect 4320 9636 4332 9639
rect 4614 9636 4620 9648
rect 4320 9608 4620 9636
rect 4320 9605 4332 9608
rect 4274 9599 4332 9605
rect 4614 9596 4620 9608
rect 4672 9596 4678 9648
rect 5902 9596 5908 9648
rect 5960 9636 5966 9648
rect 6517 9639 6575 9645
rect 6517 9636 6529 9639
rect 5960 9608 6529 9636
rect 5960 9596 5966 9608
rect 6517 9605 6529 9608
rect 6563 9605 6575 9639
rect 6517 9599 6575 9605
rect 6733 9639 6791 9645
rect 6733 9605 6745 9639
rect 6779 9605 6791 9639
rect 6733 9599 6791 9605
rect 8312 9608 9812 9636
rect 2777 9571 2835 9577
rect 2777 9537 2789 9571
rect 2823 9537 2835 9571
rect 2777 9531 2835 9537
rect 2869 9571 2927 9577
rect 2869 9537 2881 9571
rect 2915 9537 2927 9571
rect 2869 9531 2927 9537
rect 2792 9500 2820 9531
rect 3326 9528 3332 9580
rect 3384 9528 3390 9580
rect 3436 9540 3924 9568
rect 2958 9500 2964 9512
rect 2792 9472 2964 9500
rect 2958 9460 2964 9472
rect 3016 9460 3022 9512
rect 3436 9509 3464 9540
rect 3053 9503 3111 9509
rect 3053 9469 3065 9503
rect 3099 9469 3111 9503
rect 3053 9463 3111 9469
rect 3421 9503 3479 9509
rect 3421 9469 3433 9503
rect 3467 9469 3479 9503
rect 3421 9463 3479 9469
rect 3068 9364 3096 9463
rect 3602 9460 3608 9512
rect 3660 9500 3666 9512
rect 3789 9503 3847 9509
rect 3789 9500 3801 9503
rect 3660 9472 3801 9500
rect 3660 9460 3666 9472
rect 3789 9469 3801 9472
rect 3835 9469 3847 9503
rect 3896 9500 3924 9540
rect 3970 9528 3976 9580
rect 4028 9568 4034 9580
rect 4801 9571 4859 9577
rect 4801 9568 4813 9571
rect 4028 9540 4813 9568
rect 4028 9528 4034 9540
rect 4801 9537 4813 9540
rect 4847 9537 4859 9571
rect 4801 9531 4859 9537
rect 5997 9571 6055 9577
rect 5997 9537 6009 9571
rect 6043 9568 6055 9571
rect 6270 9568 6276 9580
rect 6043 9540 6276 9568
rect 6043 9537 6055 9540
rect 5997 9531 6055 9537
rect 6270 9528 6276 9540
rect 6328 9528 6334 9580
rect 6748 9568 6776 9599
rect 8312 9577 8340 9608
rect 6472 9540 6776 9568
rect 8041 9571 8099 9577
rect 6472 9512 6500 9540
rect 8041 9537 8053 9571
rect 8087 9568 8099 9571
rect 8297 9571 8355 9577
rect 8087 9540 8248 9568
rect 8087 9537 8099 9540
rect 8041 9531 8099 9537
rect 5442 9500 5448 9512
rect 3896 9472 5448 9500
rect 3789 9463 3847 9469
rect 5442 9460 5448 9472
rect 5500 9500 5506 9512
rect 5537 9503 5595 9509
rect 5537 9500 5549 9503
rect 5500 9472 5549 9500
rect 5500 9460 5506 9472
rect 5537 9469 5549 9472
rect 5583 9469 5595 9503
rect 5537 9463 5595 9469
rect 6454 9460 6460 9512
rect 6512 9460 6518 9512
rect 8220 9500 8248 9540
rect 8297 9537 8309 9571
rect 8343 9537 8355 9571
rect 8297 9531 8355 9537
rect 8662 9528 8668 9580
rect 8720 9568 8726 9580
rect 9784 9577 9812 9608
rect 12434 9596 12440 9648
rect 12492 9636 12498 9648
rect 13740 9636 13768 9676
rect 14550 9664 14556 9676
rect 14608 9664 14614 9716
rect 14752 9676 14964 9704
rect 12492 9608 13768 9636
rect 12492 9596 12498 9608
rect 13814 9596 13820 9648
rect 13872 9636 13878 9648
rect 14182 9636 14188 9648
rect 13872 9608 14188 9636
rect 13872 9596 13878 9608
rect 14182 9596 14188 9608
rect 14240 9636 14246 9648
rect 14752 9636 14780 9676
rect 14240 9608 14780 9636
rect 14240 9596 14246 9608
rect 14826 9596 14832 9648
rect 14884 9596 14890 9648
rect 14936 9636 14964 9676
rect 15381 9639 15439 9645
rect 15381 9636 15393 9639
rect 14936 9608 14970 9636
rect 9309 9571 9367 9577
rect 9309 9568 9321 9571
rect 8720 9540 9321 9568
rect 8720 9528 8726 9540
rect 9309 9537 9321 9540
rect 9355 9537 9367 9571
rect 9309 9531 9367 9537
rect 9769 9571 9827 9577
rect 9769 9537 9781 9571
rect 9815 9568 9827 9571
rect 9858 9568 9864 9580
rect 9815 9540 9864 9568
rect 9815 9537 9827 9540
rect 9769 9531 9827 9537
rect 9858 9528 9864 9540
rect 9916 9528 9922 9580
rect 10036 9571 10094 9577
rect 10036 9537 10048 9571
rect 10082 9568 10094 9571
rect 10410 9568 10416 9580
rect 10082 9540 10416 9568
rect 10082 9537 10094 9540
rect 10036 9531 10094 9537
rect 10410 9528 10416 9540
rect 10468 9528 10474 9580
rect 11514 9528 11520 9580
rect 11572 9528 11578 9580
rect 11784 9571 11842 9577
rect 11784 9537 11796 9571
rect 11830 9568 11842 9571
rect 12618 9568 12624 9580
rect 11830 9540 12624 9568
rect 11830 9537 11842 9540
rect 11784 9531 11842 9537
rect 12618 9528 12624 9540
rect 12676 9528 12682 9580
rect 13078 9528 13084 9580
rect 13136 9528 13142 9580
rect 13354 9577 13360 9580
rect 13348 9531 13360 9577
rect 13354 9528 13360 9531
rect 13412 9528 13418 9580
rect 14734 9528 14740 9580
rect 14792 9528 14798 9580
rect 14942 9577 14970 9608
rect 15028 9608 15393 9636
rect 15028 9580 15056 9608
rect 15381 9605 15393 9608
rect 15427 9605 15439 9639
rect 15381 9599 15439 9605
rect 15654 9596 15660 9648
rect 15712 9636 15718 9648
rect 15749 9639 15807 9645
rect 15749 9636 15761 9639
rect 15712 9608 15761 9636
rect 15712 9596 15718 9608
rect 15749 9605 15761 9608
rect 15795 9605 15807 9639
rect 15749 9599 15807 9605
rect 15841 9639 15899 9645
rect 15841 9605 15853 9639
rect 15887 9636 15899 9639
rect 16114 9636 16120 9648
rect 15887 9608 16120 9636
rect 15887 9605 15899 9608
rect 15841 9599 15899 9605
rect 16114 9596 16120 9608
rect 16172 9596 16178 9648
rect 14921 9571 14979 9577
rect 14921 9537 14933 9571
rect 14967 9537 14979 9571
rect 14921 9531 14979 9537
rect 15010 9528 15016 9580
rect 15068 9528 15074 9580
rect 15105 9571 15163 9577
rect 15105 9537 15117 9571
rect 15151 9537 15163 9571
rect 15105 9531 15163 9537
rect 15565 9571 15623 9577
rect 15565 9537 15577 9571
rect 15611 9537 15623 9571
rect 15565 9531 15623 9537
rect 8220 9472 8340 9500
rect 5721 9435 5779 9441
rect 5721 9401 5733 9435
rect 5767 9432 5779 9435
rect 6730 9432 6736 9444
rect 5767 9404 6736 9432
rect 5767 9401 5779 9404
rect 5721 9395 5779 9401
rect 6730 9392 6736 9404
rect 6788 9392 6794 9444
rect 8312 9432 8340 9472
rect 8386 9460 8392 9512
rect 8444 9460 8450 9512
rect 9582 9460 9588 9512
rect 9640 9460 9646 9512
rect 15120 9500 15148 9531
rect 14476 9472 15148 9500
rect 15580 9500 15608 9531
rect 16022 9528 16028 9580
rect 16080 9528 16086 9580
rect 15930 9500 15936 9512
rect 15580 9472 15936 9500
rect 9125 9435 9183 9441
rect 9125 9432 9137 9435
rect 8312 9404 9137 9432
rect 9125 9401 9137 9404
rect 9171 9401 9183 9435
rect 9125 9395 9183 9401
rect 14476 9376 14504 9472
rect 15930 9460 15936 9472
rect 15988 9460 15994 9512
rect 14550 9392 14556 9444
rect 14608 9392 14614 9444
rect 4062 9364 4068 9376
rect 3068 9336 4068 9364
rect 4062 9324 4068 9336
rect 4120 9324 4126 9376
rect 6546 9324 6552 9376
rect 6604 9324 6610 9376
rect 9214 9324 9220 9376
rect 9272 9364 9278 9376
rect 9493 9367 9551 9373
rect 9493 9364 9505 9367
rect 9272 9336 9505 9364
rect 9272 9324 9278 9336
rect 9493 9333 9505 9336
rect 9539 9333 9551 9367
rect 9493 9327 9551 9333
rect 10778 9324 10784 9376
rect 10836 9364 10842 9376
rect 11149 9367 11207 9373
rect 11149 9364 11161 9367
rect 10836 9336 11161 9364
rect 10836 9324 10842 9336
rect 11149 9333 11161 9336
rect 11195 9364 11207 9367
rect 12250 9364 12256 9376
rect 11195 9336 12256 9364
rect 11195 9333 11207 9336
rect 11149 9327 11207 9333
rect 12250 9324 12256 9336
rect 12308 9364 12314 9376
rect 13262 9364 13268 9376
rect 12308 9336 13268 9364
rect 12308 9324 12314 9336
rect 13262 9324 13268 9336
rect 13320 9324 13326 9376
rect 14458 9324 14464 9376
rect 14516 9324 14522 9376
rect 14642 9324 14648 9376
rect 14700 9364 14706 9376
rect 16209 9367 16267 9373
rect 16209 9364 16221 9367
rect 14700 9336 16221 9364
rect 14700 9324 14706 9336
rect 16209 9333 16221 9336
rect 16255 9333 16267 9367
rect 16209 9327 16267 9333
rect 1104 9274 16652 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 16652 9274
rect 1104 9200 16652 9222
rect 1854 9120 1860 9172
rect 1912 9160 1918 9172
rect 1949 9163 2007 9169
rect 1949 9160 1961 9163
rect 1912 9132 1961 9160
rect 1912 9120 1918 9132
rect 1949 9129 1961 9132
rect 1995 9129 2007 9163
rect 1949 9123 2007 9129
rect 3602 9120 3608 9172
rect 3660 9120 3666 9172
rect 3973 9163 4031 9169
rect 3973 9129 3985 9163
rect 4019 9129 4031 9163
rect 3973 9123 4031 9129
rect 1578 9052 1584 9104
rect 1636 9092 1642 9104
rect 2501 9095 2559 9101
rect 2501 9092 2513 9095
rect 1636 9064 2513 9092
rect 1636 9052 1642 9064
rect 2501 9061 2513 9064
rect 2547 9061 2559 9095
rect 2501 9055 2559 9061
rect 2314 9024 2320 9036
rect 2240 8996 2320 9024
rect 2240 8965 2268 8996
rect 2314 8984 2320 8996
rect 2372 8984 2378 9036
rect 2225 8959 2283 8965
rect 2225 8925 2237 8959
rect 2271 8925 2283 8959
rect 3142 8956 3148 8968
rect 2225 8919 2283 8925
rect 2332 8928 3148 8956
rect 1486 8848 1492 8900
rect 1544 8888 1550 8900
rect 1917 8891 1975 8897
rect 1917 8888 1929 8891
rect 1544 8860 1929 8888
rect 1544 8848 1550 8860
rect 1917 8857 1929 8860
rect 1963 8857 1975 8891
rect 1917 8851 1975 8857
rect 2038 8848 2044 8900
rect 2096 8888 2102 8900
rect 2133 8891 2191 8897
rect 2133 8888 2145 8891
rect 2096 8860 2145 8888
rect 2096 8848 2102 8860
rect 2133 8857 2145 8860
rect 2179 8857 2191 8891
rect 2133 8851 2191 8857
rect 2332 8832 2360 8928
rect 3142 8916 3148 8928
rect 3200 8916 3206 8968
rect 3237 8959 3295 8965
rect 3237 8925 3249 8959
rect 3283 8956 3295 8959
rect 3510 8956 3516 8968
rect 3283 8928 3516 8956
rect 3283 8925 3295 8928
rect 3237 8919 3295 8925
rect 3510 8916 3516 8928
rect 3568 8916 3574 8968
rect 3620 8956 3648 9120
rect 3988 9092 4016 9123
rect 4062 9120 4068 9172
rect 4120 9160 4126 9172
rect 4525 9163 4583 9169
rect 4525 9160 4537 9163
rect 4120 9132 4537 9160
rect 4120 9120 4126 9132
rect 4525 9129 4537 9132
rect 4571 9129 4583 9163
rect 4525 9123 4583 9129
rect 4798 9120 4804 9172
rect 4856 9160 4862 9172
rect 4985 9163 5043 9169
rect 4985 9160 4997 9163
rect 4856 9132 4997 9160
rect 4856 9120 4862 9132
rect 4985 9129 4997 9132
rect 5031 9129 5043 9163
rect 4985 9123 5043 9129
rect 8297 9163 8355 9169
rect 8297 9129 8309 9163
rect 8343 9160 8355 9163
rect 8386 9160 8392 9172
rect 8343 9132 8392 9160
rect 8343 9129 8355 9132
rect 8297 9123 8355 9129
rect 8386 9120 8392 9132
rect 8444 9120 8450 9172
rect 8570 9120 8576 9172
rect 8628 9120 8634 9172
rect 11422 9120 11428 9172
rect 11480 9120 11486 9172
rect 13446 9120 13452 9172
rect 13504 9120 13510 9172
rect 16206 9120 16212 9172
rect 16264 9120 16270 9172
rect 6270 9092 6276 9104
rect 3988 9064 6276 9092
rect 6270 9052 6276 9064
rect 6328 9052 6334 9104
rect 8757 9095 8815 9101
rect 8757 9061 8769 9095
rect 8803 9061 8815 9095
rect 8757 9055 8815 9061
rect 3694 8984 3700 9036
rect 3752 9024 3758 9036
rect 3752 8996 3924 9024
rect 3752 8984 3758 8996
rect 3789 8959 3847 8965
rect 3789 8956 3801 8959
rect 3620 8928 3801 8956
rect 3789 8925 3801 8928
rect 3835 8925 3847 8959
rect 3896 8956 3924 8996
rect 3970 8984 3976 9036
rect 4028 8984 4034 9036
rect 4172 8996 4844 9024
rect 4065 8959 4123 8965
rect 4065 8956 4077 8959
rect 3896 8928 4077 8956
rect 3789 8919 3847 8925
rect 4065 8925 4077 8928
rect 4111 8925 4123 8959
rect 4065 8919 4123 8925
rect 2501 8891 2559 8897
rect 2501 8857 2513 8891
rect 2547 8888 2559 8891
rect 2547 8860 2774 8888
rect 2547 8857 2559 8860
rect 2501 8851 2559 8857
rect 1762 8780 1768 8832
rect 1820 8780 1826 8832
rect 2314 8780 2320 8832
rect 2372 8780 2378 8832
rect 2746 8820 2774 8860
rect 2958 8848 2964 8900
rect 3016 8888 3022 8900
rect 3418 8888 3424 8900
rect 3016 8860 3424 8888
rect 3016 8848 3022 8860
rect 3418 8848 3424 8860
rect 3476 8848 3482 8900
rect 2866 8820 2872 8832
rect 2746 8792 2872 8820
rect 2866 8780 2872 8792
rect 2924 8820 2930 8832
rect 3326 8820 3332 8832
rect 2924 8792 3332 8820
rect 2924 8780 2930 8792
rect 3326 8780 3332 8792
rect 3384 8820 3390 8832
rect 4172 8820 4200 8996
rect 4816 8965 4844 8996
rect 8294 8984 8300 9036
rect 8352 9024 8358 9036
rect 8772 9024 8800 9055
rect 12250 9052 12256 9104
rect 12308 9092 12314 9104
rect 14458 9092 14464 9104
rect 12308 9064 14464 9092
rect 12308 9052 12314 9064
rect 8352 8996 8800 9024
rect 8352 8984 8358 8996
rect 4709 8959 4767 8965
rect 4709 8956 4721 8959
rect 4264 8928 4721 8956
rect 4264 8829 4292 8928
rect 4709 8925 4721 8928
rect 4755 8925 4767 8959
rect 4709 8919 4767 8925
rect 4801 8959 4859 8965
rect 4801 8925 4813 8959
rect 4847 8925 4859 8959
rect 4801 8919 4859 8925
rect 5077 8959 5135 8965
rect 5077 8925 5089 8959
rect 5123 8956 5135 8959
rect 5258 8956 5264 8968
rect 5123 8928 5264 8956
rect 5123 8925 5135 8928
rect 5077 8919 5135 8925
rect 5258 8916 5264 8928
rect 5316 8916 5322 8968
rect 5445 8959 5503 8965
rect 5445 8925 5457 8959
rect 5491 8925 5503 8959
rect 5445 8919 5503 8925
rect 5460 8888 5488 8919
rect 5534 8916 5540 8968
rect 5592 8956 5598 8968
rect 6825 8959 6883 8965
rect 6825 8956 6837 8959
rect 5592 8928 6837 8956
rect 5592 8916 5598 8928
rect 6825 8925 6837 8928
rect 6871 8925 6883 8959
rect 6825 8919 6883 8925
rect 6917 8959 6975 8965
rect 6917 8925 6929 8959
rect 6963 8925 6975 8959
rect 6917 8919 6975 8925
rect 7184 8959 7242 8965
rect 7184 8925 7196 8959
rect 7230 8956 7242 8959
rect 7650 8956 7656 8968
rect 7230 8928 7656 8956
rect 7230 8925 7242 8928
rect 7184 8919 7242 8925
rect 6089 8891 6147 8897
rect 6089 8888 6101 8891
rect 5460 8860 6101 8888
rect 6089 8857 6101 8860
rect 6135 8888 6147 8891
rect 6362 8888 6368 8900
rect 6135 8860 6368 8888
rect 6135 8857 6147 8860
rect 6089 8851 6147 8857
rect 6362 8848 6368 8860
rect 6420 8888 6426 8900
rect 6638 8888 6644 8900
rect 6420 8860 6644 8888
rect 6420 8848 6426 8860
rect 6638 8848 6644 8860
rect 6696 8888 6702 8900
rect 6932 8888 6960 8919
rect 7650 8916 7656 8928
rect 7708 8916 7714 8968
rect 6696 8860 6960 8888
rect 6696 8848 6702 8860
rect 8386 8848 8392 8900
rect 8444 8848 8450 8900
rect 8772 8888 8800 8996
rect 11974 8984 11980 9036
rect 12032 8984 12038 9036
rect 12158 8984 12164 9036
rect 12216 9024 12222 9036
rect 12216 8996 13492 9024
rect 12216 8984 12222 8996
rect 8941 8959 8999 8965
rect 8941 8925 8953 8959
rect 8987 8956 8999 8959
rect 11333 8959 11391 8965
rect 8987 8928 9904 8956
rect 8987 8925 8999 8928
rect 8941 8919 8999 8925
rect 9876 8900 9904 8928
rect 11333 8925 11345 8959
rect 11379 8956 11391 8959
rect 11698 8956 11704 8968
rect 11379 8928 11704 8956
rect 11379 8925 11391 8928
rect 11333 8919 11391 8925
rect 11698 8916 11704 8928
rect 11756 8956 11762 8968
rect 13464 8965 13492 8996
rect 13357 8959 13415 8965
rect 13357 8956 13369 8959
rect 11756 8928 13369 8956
rect 11756 8916 11762 8928
rect 13357 8925 13369 8928
rect 13403 8925 13415 8959
rect 13357 8919 13415 8925
rect 13449 8959 13507 8965
rect 13449 8925 13461 8959
rect 13495 8925 13507 8959
rect 13449 8919 13507 8925
rect 13538 8916 13544 8968
rect 13596 8916 13602 8968
rect 13814 8916 13820 8968
rect 13872 8916 13878 8968
rect 14292 8965 14320 9064
rect 14458 9052 14464 9064
rect 14516 9052 14522 9104
rect 14277 8959 14335 8965
rect 14277 8925 14289 8959
rect 14323 8925 14335 8959
rect 14277 8919 14335 8925
rect 14918 8916 14924 8968
rect 14976 8956 14982 8968
rect 15105 8959 15163 8965
rect 15105 8956 15117 8959
rect 14976 8928 15117 8956
rect 14976 8916 14982 8928
rect 15105 8925 15117 8928
rect 15151 8925 15163 8959
rect 15105 8919 15163 8925
rect 15194 8916 15200 8968
rect 15252 8916 15258 8968
rect 15289 8959 15347 8965
rect 15289 8925 15301 8959
rect 15335 8925 15347 8959
rect 15289 8919 15347 8925
rect 9186 8891 9244 8897
rect 9186 8888 9198 8891
rect 8772 8860 9198 8888
rect 9186 8857 9198 8860
rect 9232 8857 9244 8891
rect 9186 8851 9244 8857
rect 9858 8848 9864 8900
rect 9916 8888 9922 8900
rect 10505 8891 10563 8897
rect 10505 8888 10517 8891
rect 9916 8860 10517 8888
rect 9916 8848 9922 8860
rect 10505 8857 10517 8860
rect 10551 8857 10563 8891
rect 10505 8851 10563 8857
rect 11793 8891 11851 8897
rect 11793 8857 11805 8891
rect 11839 8888 11851 8891
rect 12434 8888 12440 8900
rect 11839 8860 12440 8888
rect 11839 8857 11851 8860
rect 11793 8851 11851 8857
rect 12434 8848 12440 8860
rect 12492 8848 12498 8900
rect 12526 8848 12532 8900
rect 12584 8848 12590 8900
rect 13832 8888 13860 8916
rect 14461 8891 14519 8897
rect 14461 8888 14473 8891
rect 13832 8860 14473 8888
rect 14461 8857 14473 8860
rect 14507 8888 14519 8891
rect 15010 8888 15016 8900
rect 14507 8860 15016 8888
rect 14507 8857 14519 8860
rect 14461 8851 14519 8857
rect 15010 8848 15016 8860
rect 15068 8848 15074 8900
rect 15304 8888 15332 8919
rect 15378 8916 15384 8968
rect 15436 8956 15442 8968
rect 15473 8959 15531 8965
rect 15473 8956 15485 8959
rect 15436 8928 15485 8956
rect 15436 8916 15442 8928
rect 15473 8925 15485 8928
rect 15519 8925 15531 8959
rect 15473 8919 15531 8925
rect 15746 8916 15752 8968
rect 15804 8916 15810 8968
rect 15838 8916 15844 8968
rect 15896 8956 15902 8968
rect 16025 8959 16083 8965
rect 16025 8956 16037 8959
rect 15896 8928 16037 8956
rect 15896 8916 15902 8928
rect 16025 8925 16037 8928
rect 16071 8925 16083 8959
rect 16025 8919 16083 8925
rect 15565 8891 15623 8897
rect 15565 8888 15577 8891
rect 15304 8860 15577 8888
rect 15565 8857 15577 8860
rect 15611 8857 15623 8891
rect 15565 8851 15623 8857
rect 15930 8848 15936 8900
rect 15988 8888 15994 8900
rect 16114 8888 16120 8900
rect 15988 8860 16120 8888
rect 15988 8848 15994 8860
rect 16114 8848 16120 8860
rect 16172 8848 16178 8900
rect 3384 8792 4200 8820
rect 4249 8823 4307 8829
rect 3384 8780 3390 8792
rect 4249 8789 4261 8823
rect 4295 8789 4307 8823
rect 4249 8783 4307 8789
rect 8294 8780 8300 8832
rect 8352 8820 8358 8832
rect 8589 8823 8647 8829
rect 8589 8820 8601 8823
rect 8352 8792 8601 8820
rect 8352 8780 8358 8792
rect 8589 8789 8601 8792
rect 8635 8820 8647 8823
rect 9030 8820 9036 8832
rect 8635 8792 9036 8820
rect 8635 8789 8647 8792
rect 8589 8783 8647 8789
rect 9030 8780 9036 8792
rect 9088 8780 9094 8832
rect 10321 8823 10379 8829
rect 10321 8789 10333 8823
rect 10367 8820 10379 8823
rect 11146 8820 11152 8832
rect 10367 8792 11152 8820
rect 10367 8789 10379 8792
rect 10321 8783 10379 8789
rect 11146 8780 11152 8792
rect 11204 8780 11210 8832
rect 11882 8780 11888 8832
rect 11940 8780 11946 8832
rect 12342 8780 12348 8832
rect 12400 8820 12406 8832
rect 13817 8823 13875 8829
rect 13817 8820 13829 8823
rect 12400 8792 13829 8820
rect 12400 8780 12406 8792
rect 13817 8789 13829 8792
rect 13863 8789 13875 8823
rect 13817 8783 13875 8789
rect 13906 8780 13912 8832
rect 13964 8820 13970 8832
rect 14093 8823 14151 8829
rect 14093 8820 14105 8823
rect 13964 8792 14105 8820
rect 13964 8780 13970 8792
rect 14093 8789 14105 8792
rect 14139 8789 14151 8823
rect 14093 8783 14151 8789
rect 14826 8780 14832 8832
rect 14884 8780 14890 8832
rect 1104 8730 16652 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 16652 8730
rect 1104 8656 16652 8678
rect 1397 8619 1455 8625
rect 1397 8585 1409 8619
rect 1443 8616 1455 8619
rect 2314 8616 2320 8628
rect 1443 8588 2320 8616
rect 1443 8585 1455 8588
rect 1397 8579 1455 8585
rect 2314 8576 2320 8588
rect 2372 8576 2378 8628
rect 3878 8576 3884 8628
rect 3936 8616 3942 8628
rect 4341 8619 4399 8625
rect 4341 8616 4353 8619
rect 3936 8588 4353 8616
rect 3936 8576 3942 8588
rect 4341 8585 4353 8588
rect 4387 8585 4399 8619
rect 4341 8579 4399 8585
rect 4706 8576 4712 8628
rect 4764 8616 4770 8628
rect 5001 8619 5059 8625
rect 5001 8616 5013 8619
rect 4764 8588 5013 8616
rect 4764 8576 4770 8588
rect 5001 8585 5013 8588
rect 5047 8585 5059 8619
rect 5001 8579 5059 8585
rect 5261 8619 5319 8625
rect 5261 8585 5273 8619
rect 5307 8616 5319 8619
rect 5350 8616 5356 8628
rect 5307 8588 5356 8616
rect 5307 8585 5319 8588
rect 5261 8579 5319 8585
rect 5350 8576 5356 8588
rect 5408 8576 5414 8628
rect 8297 8619 8355 8625
rect 8297 8585 8309 8619
rect 8343 8616 8355 8619
rect 8478 8616 8484 8628
rect 8343 8588 8484 8616
rect 8343 8585 8355 8588
rect 8297 8579 8355 8585
rect 8478 8576 8484 8588
rect 8536 8576 8542 8628
rect 9766 8576 9772 8628
rect 9824 8576 9830 8628
rect 10410 8576 10416 8628
rect 10468 8576 10474 8628
rect 10778 8576 10784 8628
rect 10836 8576 10842 8628
rect 12529 8619 12587 8625
rect 12529 8585 12541 8619
rect 12575 8616 12587 8619
rect 12618 8616 12624 8628
rect 12575 8588 12624 8616
rect 12575 8585 12587 8588
rect 12529 8579 12587 8585
rect 12618 8576 12624 8588
rect 12676 8576 12682 8628
rect 12894 8576 12900 8628
rect 12952 8616 12958 8628
rect 12989 8619 13047 8625
rect 12989 8616 13001 8619
rect 12952 8588 13001 8616
rect 12952 8576 12958 8588
rect 12989 8585 13001 8588
rect 13035 8585 13047 8619
rect 12989 8579 13047 8585
rect 2406 8508 2412 8560
rect 2464 8548 2470 8560
rect 2464 8520 2728 8548
rect 2464 8508 2470 8520
rect 2498 8440 2504 8492
rect 2556 8489 2562 8492
rect 2556 8443 2568 8489
rect 2556 8440 2562 8443
rect 2700 8412 2728 8520
rect 2866 8508 2872 8560
rect 2924 8508 2930 8560
rect 3069 8551 3127 8557
rect 3069 8548 3081 8551
rect 2976 8520 3081 8548
rect 2774 8440 2780 8492
rect 2832 8440 2838 8492
rect 2976 8412 3004 8520
rect 3069 8517 3081 8520
rect 3115 8517 3127 8551
rect 3069 8511 3127 8517
rect 3970 8508 3976 8560
rect 4028 8548 4034 8560
rect 4525 8551 4583 8557
rect 4525 8548 4537 8551
rect 4028 8520 4537 8548
rect 4028 8508 4034 8520
rect 4525 8517 4537 8520
rect 4571 8517 4583 8551
rect 4525 8511 4583 8517
rect 4801 8551 4859 8557
rect 4801 8517 4813 8551
rect 4847 8548 4859 8551
rect 5534 8548 5540 8560
rect 4847 8520 5540 8548
rect 4847 8517 4859 8520
rect 4801 8511 4859 8517
rect 5534 8508 5540 8520
rect 5592 8508 5598 8560
rect 6365 8551 6423 8557
rect 6365 8548 6377 8551
rect 5644 8520 6377 8548
rect 3329 8483 3387 8489
rect 3329 8480 3341 8483
rect 2700 8384 3004 8412
rect 3252 8452 3341 8480
rect 2958 8304 2964 8356
rect 3016 8344 3022 8356
rect 3252 8353 3280 8452
rect 3329 8449 3341 8452
rect 3375 8449 3387 8483
rect 3329 8443 3387 8449
rect 3510 8440 3516 8492
rect 3568 8440 3574 8492
rect 4709 8483 4767 8489
rect 4709 8449 4721 8483
rect 4755 8449 4767 8483
rect 4709 8443 4767 8449
rect 4724 8412 4752 8443
rect 5442 8440 5448 8492
rect 5500 8440 5506 8492
rect 5644 8489 5672 8520
rect 6365 8517 6377 8520
rect 6411 8517 6423 8551
rect 6365 8511 6423 8517
rect 7184 8551 7242 8557
rect 7184 8517 7196 8551
rect 7230 8548 7242 8551
rect 8110 8548 8116 8560
rect 7230 8520 8116 8548
rect 7230 8517 7242 8520
rect 7184 8511 7242 8517
rect 8110 8508 8116 8520
rect 8168 8508 8174 8560
rect 12161 8551 12219 8557
rect 8404 8520 9904 8548
rect 5629 8483 5687 8489
rect 5629 8449 5641 8483
rect 5675 8449 5687 8483
rect 5629 8443 5687 8449
rect 5718 8440 5724 8492
rect 5776 8440 5782 8492
rect 6270 8440 6276 8492
rect 6328 8480 6334 8492
rect 8404 8489 8432 8520
rect 9876 8492 9904 8520
rect 12161 8517 12173 8551
rect 12207 8548 12219 8551
rect 12802 8548 12808 8560
rect 12207 8520 12808 8548
rect 12207 8517 12219 8520
rect 12161 8511 12219 8517
rect 12802 8508 12808 8520
rect 12860 8508 12866 8560
rect 6549 8483 6607 8489
rect 6549 8480 6561 8483
rect 6328 8452 6561 8480
rect 6328 8440 6334 8452
rect 6549 8449 6561 8452
rect 6595 8449 6607 8483
rect 6549 8443 6607 8449
rect 8389 8483 8447 8489
rect 8389 8449 8401 8483
rect 8435 8449 8447 8483
rect 8389 8443 8447 8449
rect 8478 8440 8484 8492
rect 8536 8480 8542 8492
rect 8645 8483 8703 8489
rect 8645 8480 8657 8483
rect 8536 8452 8657 8480
rect 8536 8440 8542 8452
rect 8645 8449 8657 8452
rect 8691 8449 8703 8483
rect 8645 8443 8703 8449
rect 9858 8440 9864 8492
rect 9916 8440 9922 8492
rect 10873 8483 10931 8489
rect 10873 8449 10885 8483
rect 10919 8480 10931 8483
rect 11882 8480 11888 8492
rect 10919 8452 11888 8480
rect 10919 8449 10931 8452
rect 10873 8443 10931 8449
rect 4798 8412 4804 8424
rect 4724 8384 4804 8412
rect 4798 8372 4804 8384
rect 4856 8372 4862 8424
rect 5902 8412 5908 8424
rect 5184 8384 5908 8412
rect 3237 8347 3295 8353
rect 3237 8344 3249 8347
rect 3016 8316 3249 8344
rect 3016 8304 3022 8316
rect 3237 8313 3249 8316
rect 3283 8313 3295 8347
rect 3237 8307 3295 8313
rect 3329 8347 3387 8353
rect 3329 8313 3341 8347
rect 3375 8344 3387 8347
rect 4062 8344 4068 8356
rect 3375 8316 4068 8344
rect 3375 8313 3387 8316
rect 3329 8307 3387 8313
rect 4062 8304 4068 8316
rect 4120 8304 4126 8356
rect 5184 8353 5212 8384
rect 5902 8372 5908 8384
rect 5960 8372 5966 8424
rect 6730 8372 6736 8424
rect 6788 8372 6794 8424
rect 6917 8415 6975 8421
rect 6917 8381 6929 8415
rect 6963 8381 6975 8415
rect 6917 8375 6975 8381
rect 5169 8347 5227 8353
rect 5169 8313 5181 8347
rect 5215 8313 5227 8347
rect 5169 8307 5227 8313
rect 5534 8304 5540 8356
rect 5592 8304 5598 8356
rect 6362 8304 6368 8356
rect 6420 8344 6426 8356
rect 6932 8344 6960 8375
rect 9582 8372 9588 8424
rect 9640 8412 9646 8424
rect 10888 8412 10916 8443
rect 11882 8440 11888 8452
rect 11940 8480 11946 8492
rect 12069 8483 12127 8489
rect 12069 8480 12081 8483
rect 11940 8452 12081 8480
rect 11940 8440 11946 8452
rect 12069 8449 12081 8452
rect 12115 8480 12127 8483
rect 12897 8483 12955 8489
rect 12897 8480 12909 8483
rect 12115 8452 12909 8480
rect 12115 8449 12127 8452
rect 12069 8443 12127 8449
rect 12897 8449 12909 8452
rect 12943 8449 12955 8483
rect 13004 8480 13032 8579
rect 13354 8576 13360 8628
rect 13412 8576 13418 8628
rect 13722 8576 13728 8628
rect 13780 8616 13786 8628
rect 13780 8588 14780 8616
rect 13780 8576 13786 8588
rect 14642 8548 14648 8560
rect 14384 8520 14648 8548
rect 13633 8483 13691 8489
rect 13633 8480 13645 8483
rect 13004 8452 13645 8480
rect 12897 8443 12955 8449
rect 13633 8449 13645 8452
rect 13679 8449 13691 8483
rect 13633 8443 13691 8449
rect 13722 8440 13728 8492
rect 13780 8440 13786 8492
rect 13817 8483 13875 8489
rect 13817 8449 13829 8483
rect 13863 8480 13875 8483
rect 13906 8480 13912 8492
rect 13863 8452 13912 8480
rect 13863 8449 13875 8452
rect 13817 8443 13875 8449
rect 13906 8440 13912 8452
rect 13964 8440 13970 8492
rect 13998 8440 14004 8492
rect 14056 8480 14062 8492
rect 14384 8489 14412 8520
rect 14642 8508 14648 8520
rect 14700 8508 14706 8560
rect 14185 8483 14243 8489
rect 14185 8480 14197 8483
rect 14056 8452 14197 8480
rect 14056 8440 14062 8452
rect 14185 8449 14197 8452
rect 14231 8449 14243 8483
rect 14185 8443 14243 8449
rect 14369 8483 14427 8489
rect 14369 8449 14381 8483
rect 14415 8449 14427 8483
rect 14369 8443 14427 8449
rect 14461 8483 14519 8489
rect 14461 8449 14473 8483
rect 14507 8449 14519 8483
rect 14461 8443 14519 8449
rect 14553 8483 14611 8489
rect 14553 8449 14565 8483
rect 14599 8480 14611 8483
rect 14752 8480 14780 8588
rect 15746 8576 15752 8628
rect 15804 8616 15810 8628
rect 16301 8619 16359 8625
rect 16301 8616 16313 8619
rect 15804 8588 16313 8616
rect 15804 8576 15810 8588
rect 16301 8585 16313 8588
rect 16347 8585 16359 8619
rect 16301 8579 16359 8585
rect 14826 8508 14832 8560
rect 14884 8548 14890 8560
rect 15166 8551 15224 8557
rect 15166 8548 15178 8551
rect 14884 8520 15178 8548
rect 14884 8508 14890 8520
rect 15166 8517 15178 8520
rect 15212 8517 15224 8551
rect 15166 8511 15224 8517
rect 15746 8480 15752 8492
rect 14599 8452 15752 8480
rect 14599 8449 14611 8452
rect 14553 8443 14611 8449
rect 9640 8384 10916 8412
rect 9640 8372 9646 8384
rect 10962 8372 10968 8424
rect 11020 8372 11026 8424
rect 12342 8372 12348 8424
rect 12400 8372 12406 8424
rect 13078 8372 13084 8424
rect 13136 8372 13142 8424
rect 13354 8372 13360 8424
rect 13412 8412 13418 8424
rect 13740 8412 13768 8440
rect 14476 8412 14504 8443
rect 13412 8384 13768 8412
rect 14384 8384 14504 8412
rect 13412 8372 13418 8384
rect 14384 8356 14412 8384
rect 6420 8316 6960 8344
rect 6420 8304 6426 8316
rect 14366 8304 14372 8356
rect 14424 8304 14430 8356
rect 3053 8279 3111 8285
rect 3053 8245 3065 8279
rect 3099 8276 3111 8279
rect 3142 8276 3148 8288
rect 3099 8248 3148 8276
rect 3099 8245 3111 8248
rect 3053 8239 3111 8245
rect 3142 8236 3148 8248
rect 3200 8236 3206 8288
rect 4614 8236 4620 8288
rect 4672 8276 4678 8288
rect 4985 8279 5043 8285
rect 4985 8276 4997 8279
rect 4672 8248 4997 8276
rect 4672 8236 4678 8248
rect 4985 8245 4997 8248
rect 5031 8276 5043 8279
rect 5350 8276 5356 8288
rect 5031 8248 5356 8276
rect 5031 8245 5043 8248
rect 4985 8239 5043 8245
rect 5350 8236 5356 8248
rect 5408 8236 5414 8288
rect 9766 8236 9772 8288
rect 9824 8276 9830 8288
rect 10686 8276 10692 8288
rect 9824 8248 10692 8276
rect 9824 8236 9830 8248
rect 10686 8236 10692 8248
rect 10744 8276 10750 8288
rect 11238 8276 11244 8288
rect 10744 8248 11244 8276
rect 10744 8236 10750 8248
rect 11238 8236 11244 8248
rect 11296 8236 11302 8288
rect 11701 8279 11759 8285
rect 11701 8245 11713 8279
rect 11747 8276 11759 8279
rect 11790 8276 11796 8288
rect 11747 8248 11796 8276
rect 11747 8245 11759 8248
rect 11701 8239 11759 8245
rect 11790 8236 11796 8248
rect 11848 8236 11854 8288
rect 12986 8236 12992 8288
rect 13044 8276 13050 8288
rect 14568 8276 14596 8443
rect 15746 8440 15752 8452
rect 15804 8440 15810 8492
rect 14918 8372 14924 8424
rect 14976 8372 14982 8424
rect 14829 8347 14887 8353
rect 14829 8313 14841 8347
rect 14875 8344 14887 8347
rect 14875 8316 14964 8344
rect 14875 8313 14887 8316
rect 14829 8307 14887 8313
rect 13044 8248 14596 8276
rect 14936 8276 14964 8316
rect 15194 8276 15200 8288
rect 14936 8248 15200 8276
rect 13044 8236 13050 8248
rect 15194 8236 15200 8248
rect 15252 8236 15258 8288
rect 1104 8186 16652 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 16652 8186
rect 1104 8112 16652 8134
rect 2774 8072 2780 8084
rect 1596 8044 2780 8072
rect 1596 7945 1624 8044
rect 2774 8032 2780 8044
rect 2832 8032 2838 8084
rect 2866 8032 2872 8084
rect 2924 8072 2930 8084
rect 2961 8075 3019 8081
rect 2961 8072 2973 8075
rect 2924 8044 2973 8072
rect 2924 8032 2930 8044
rect 2961 8041 2973 8044
rect 3007 8072 3019 8075
rect 5353 8075 5411 8081
rect 3007 8044 3648 8072
rect 3007 8041 3019 8044
rect 2961 8035 3019 8041
rect 2590 7964 2596 8016
rect 2648 8004 2654 8016
rect 3620 8013 3648 8044
rect 5353 8041 5365 8075
rect 5399 8072 5411 8075
rect 6457 8075 6515 8081
rect 6457 8072 6469 8075
rect 5399 8044 6469 8072
rect 5399 8041 5411 8044
rect 5353 8035 5411 8041
rect 6457 8041 6469 8044
rect 6503 8041 6515 8075
rect 6457 8035 6515 8041
rect 8113 8075 8171 8081
rect 8113 8041 8125 8075
rect 8159 8072 8171 8075
rect 8386 8072 8392 8084
rect 8159 8044 8392 8072
rect 8159 8041 8171 8044
rect 8113 8035 8171 8041
rect 8386 8032 8392 8044
rect 8444 8032 8450 8084
rect 8938 8032 8944 8084
rect 8996 8032 9002 8084
rect 9309 8075 9367 8081
rect 9309 8041 9321 8075
rect 9355 8041 9367 8075
rect 9309 8035 9367 8041
rect 9493 8075 9551 8081
rect 9493 8041 9505 8075
rect 9539 8072 9551 8075
rect 11054 8072 11060 8084
rect 9539 8044 11060 8072
rect 9539 8041 9551 8044
rect 9493 8035 9551 8041
rect 3053 8007 3111 8013
rect 3053 8004 3065 8007
rect 2648 7976 3065 8004
rect 2648 7964 2654 7976
rect 3053 7973 3065 7976
rect 3099 7973 3111 8007
rect 3053 7967 3111 7973
rect 3605 8007 3663 8013
rect 3605 7973 3617 8007
rect 3651 7973 3663 8007
rect 3605 7967 3663 7973
rect 4065 8007 4123 8013
rect 4065 7973 4077 8007
rect 4111 8004 4123 8007
rect 5442 8004 5448 8016
rect 4111 7976 5448 8004
rect 4111 7973 4123 7976
rect 4065 7967 4123 7973
rect 1581 7939 1639 7945
rect 1581 7905 1593 7939
rect 1627 7905 1639 7939
rect 3068 7936 3096 7967
rect 5442 7964 5448 7976
rect 5500 7964 5506 8016
rect 5626 7964 5632 8016
rect 5684 8004 5690 8016
rect 5721 8007 5779 8013
rect 5721 8004 5733 8007
rect 5684 7976 5733 8004
rect 5684 7964 5690 7976
rect 5721 7973 5733 7976
rect 5767 8004 5779 8007
rect 5813 8007 5871 8013
rect 5813 8004 5825 8007
rect 5767 7976 5825 8004
rect 5767 7973 5779 7976
rect 5721 7967 5779 7973
rect 5813 7973 5825 7976
rect 5859 7973 5871 8007
rect 5813 7967 5871 7973
rect 6270 7964 6276 8016
rect 6328 8004 6334 8016
rect 9324 8004 9352 8035
rect 11054 8032 11060 8044
rect 11112 8032 11118 8084
rect 11333 8075 11391 8081
rect 11333 8041 11345 8075
rect 11379 8072 11391 8075
rect 11698 8072 11704 8084
rect 11379 8044 11704 8072
rect 11379 8041 11391 8044
rect 11333 8035 11391 8041
rect 11698 8032 11704 8044
rect 11756 8072 11762 8084
rect 12158 8072 12164 8084
rect 11756 8044 12164 8072
rect 11756 8032 11762 8044
rect 12158 8032 12164 8044
rect 12216 8032 12222 8084
rect 12710 8032 12716 8084
rect 12768 8072 12774 8084
rect 13265 8075 13323 8081
rect 13265 8072 13277 8075
rect 12768 8044 13277 8072
rect 12768 8032 12774 8044
rect 13265 8041 13277 8044
rect 13311 8072 13323 8075
rect 13446 8072 13452 8084
rect 13311 8044 13452 8072
rect 13311 8041 13323 8044
rect 13265 8035 13323 8041
rect 13446 8032 13452 8044
rect 13504 8032 13510 8084
rect 16022 8032 16028 8084
rect 16080 8072 16086 8084
rect 16301 8075 16359 8081
rect 16301 8072 16313 8075
rect 16080 8044 16313 8072
rect 16080 8032 16086 8044
rect 16301 8041 16313 8044
rect 16347 8041 16359 8075
rect 16301 8035 16359 8041
rect 9766 8004 9772 8016
rect 6328 7976 7512 8004
rect 9324 7976 9772 8004
rect 6328 7964 6334 7976
rect 6917 7939 6975 7945
rect 6917 7936 6929 7939
rect 3068 7908 4384 7936
rect 1581 7899 1639 7905
rect 1596 7868 1624 7899
rect 1670 7868 1676 7880
rect 1596 7840 1676 7868
rect 1670 7828 1676 7840
rect 1728 7828 1734 7880
rect 1854 7877 1860 7880
rect 1848 7868 1860 7877
rect 1815 7840 1860 7868
rect 1848 7831 1860 7840
rect 1854 7828 1860 7831
rect 1912 7828 1918 7880
rect 3050 7828 3056 7880
rect 3108 7868 3114 7880
rect 3421 7871 3479 7877
rect 3421 7868 3433 7871
rect 3108 7840 3433 7868
rect 3108 7828 3114 7840
rect 3421 7837 3433 7840
rect 3467 7868 3479 7871
rect 3510 7868 3516 7880
rect 3467 7840 3516 7868
rect 3467 7837 3479 7840
rect 3421 7831 3479 7837
rect 3510 7828 3516 7840
rect 3568 7828 3574 7880
rect 3804 7877 3832 7908
rect 3789 7871 3847 7877
rect 3789 7837 3801 7871
rect 3835 7837 3847 7871
rect 3789 7831 3847 7837
rect 3881 7871 3939 7877
rect 3881 7837 3893 7871
rect 3927 7868 3939 7871
rect 3970 7868 3976 7880
rect 3927 7840 3976 7868
rect 3927 7837 3939 7840
rect 3881 7831 3939 7837
rect 3970 7828 3976 7840
rect 4028 7828 4034 7880
rect 4154 7828 4160 7880
rect 4212 7828 4218 7880
rect 4356 7877 4384 7908
rect 6196 7908 6929 7936
rect 4341 7871 4399 7877
rect 4341 7837 4353 7871
rect 4387 7837 4399 7871
rect 4341 7831 4399 7837
rect 5718 7828 5724 7880
rect 5776 7868 5782 7880
rect 6086 7868 6092 7880
rect 5776 7840 6092 7868
rect 5776 7828 5782 7840
rect 6086 7828 6092 7840
rect 6144 7868 6150 7880
rect 6196 7877 6224 7908
rect 6917 7905 6929 7908
rect 6963 7905 6975 7939
rect 6917 7899 6975 7905
rect 6181 7871 6239 7877
rect 6181 7868 6193 7871
rect 6144 7840 6193 7868
rect 6144 7828 6150 7840
rect 6181 7837 6193 7840
rect 6227 7837 6239 7871
rect 6181 7831 6239 7837
rect 6270 7828 6276 7880
rect 6328 7868 6334 7880
rect 6641 7871 6699 7877
rect 6641 7868 6653 7871
rect 6328 7840 6653 7868
rect 6328 7828 6334 7840
rect 6641 7837 6653 7840
rect 6687 7837 6699 7871
rect 6641 7831 6699 7837
rect 6730 7828 6736 7880
rect 6788 7828 6794 7880
rect 7484 7877 7512 7976
rect 9766 7964 9772 7976
rect 9824 7964 9830 8016
rect 12802 7964 12808 8016
rect 12860 8004 12866 8016
rect 12897 8007 12955 8013
rect 12897 8004 12909 8007
rect 12860 7976 12909 8004
rect 12860 7964 12866 7976
rect 12897 7973 12909 7976
rect 12943 8004 12955 8007
rect 14826 8004 14832 8016
rect 12943 7976 14832 8004
rect 12943 7973 12955 7976
rect 12897 7967 12955 7973
rect 14826 7964 14832 7976
rect 14884 7964 14890 8016
rect 8570 7896 8576 7948
rect 8628 7936 8634 7948
rect 8665 7939 8723 7945
rect 8665 7936 8677 7939
rect 8628 7908 8677 7936
rect 8628 7896 8634 7908
rect 8665 7905 8677 7908
rect 8711 7936 8723 7939
rect 9217 7939 9275 7945
rect 9217 7936 9229 7939
rect 8711 7908 9229 7936
rect 8711 7905 8723 7908
rect 8665 7899 8723 7905
rect 9217 7905 9229 7908
rect 9263 7905 9275 7939
rect 11517 7939 11575 7945
rect 11517 7936 11529 7939
rect 9217 7899 9275 7905
rect 10888 7908 11529 7936
rect 6825 7871 6883 7877
rect 6825 7837 6837 7871
rect 6871 7837 6883 7871
rect 6825 7831 6883 7837
rect 7469 7871 7527 7877
rect 7469 7837 7481 7871
rect 7515 7837 7527 7871
rect 7469 7831 7527 7837
rect 7837 7871 7895 7877
rect 7837 7837 7849 7871
rect 7883 7837 7895 7871
rect 7837 7831 7895 7837
rect 8021 7871 8079 7877
rect 8021 7837 8033 7871
rect 8067 7868 8079 7871
rect 9309 7871 9367 7877
rect 9309 7868 9321 7871
rect 8067 7840 9321 7868
rect 8067 7837 8079 7840
rect 8021 7831 8079 7837
rect 9309 7837 9321 7840
rect 9355 7837 9367 7871
rect 9309 7831 9367 7837
rect 2406 7760 2412 7812
rect 2464 7800 2470 7812
rect 3237 7803 3295 7809
rect 3237 7800 3249 7803
rect 2464 7772 3249 7800
rect 2464 7760 2470 7772
rect 3237 7769 3249 7772
rect 3283 7769 3295 7803
rect 4065 7803 4123 7809
rect 4065 7800 4077 7803
rect 3237 7763 3295 7769
rect 3436 7772 4077 7800
rect 3436 7744 3464 7772
rect 4065 7769 4077 7772
rect 4111 7769 4123 7803
rect 4065 7763 4123 7769
rect 4798 7760 4804 7812
rect 4856 7800 4862 7812
rect 6365 7803 6423 7809
rect 6365 7800 6377 7803
rect 4856 7772 6377 7800
rect 4856 7760 4862 7772
rect 6365 7769 6377 7772
rect 6411 7800 6423 7803
rect 6840 7800 6868 7831
rect 6914 7800 6920 7812
rect 6411 7772 6920 7800
rect 6411 7769 6423 7772
rect 6365 7763 6423 7769
rect 6914 7760 6920 7772
rect 6972 7800 6978 7812
rect 7285 7803 7343 7809
rect 7285 7800 7297 7803
rect 6972 7772 7297 7800
rect 6972 7760 6978 7772
rect 7285 7769 7297 7772
rect 7331 7769 7343 7803
rect 7852 7800 7880 7831
rect 9122 7800 9128 7812
rect 7852 7772 9128 7800
rect 7285 7763 7343 7769
rect 9122 7760 9128 7772
rect 9180 7760 9186 7812
rect 9324 7800 9352 7831
rect 9858 7828 9864 7880
rect 9916 7868 9922 7880
rect 10888 7877 10916 7908
rect 11517 7905 11529 7908
rect 11563 7905 11575 7939
rect 11517 7899 11575 7905
rect 12526 7896 12532 7948
rect 12584 7936 12590 7948
rect 14918 7936 14924 7948
rect 12584 7908 14924 7936
rect 12584 7896 12590 7908
rect 14918 7896 14924 7908
rect 14976 7896 14982 7948
rect 10873 7871 10931 7877
rect 10873 7868 10885 7871
rect 9916 7840 10885 7868
rect 9916 7828 9922 7840
rect 10873 7837 10885 7840
rect 10919 7837 10931 7871
rect 10873 7831 10931 7837
rect 10965 7871 11023 7877
rect 10965 7837 10977 7871
rect 11011 7837 11023 7871
rect 10965 7831 11023 7837
rect 11149 7871 11207 7877
rect 11149 7837 11161 7871
rect 11195 7868 11207 7871
rect 11238 7868 11244 7880
rect 11195 7840 11244 7868
rect 11195 7837 11207 7840
rect 11149 7831 11207 7837
rect 10410 7800 10416 7812
rect 9324 7772 10416 7800
rect 10410 7760 10416 7772
rect 10468 7760 10474 7812
rect 10594 7760 10600 7812
rect 10652 7809 10658 7812
rect 10652 7800 10664 7809
rect 10652 7772 10697 7800
rect 10652 7763 10664 7772
rect 10652 7760 10658 7763
rect 2866 7692 2872 7744
rect 2924 7732 2930 7744
rect 3142 7732 3148 7744
rect 2924 7704 3148 7732
rect 2924 7692 2930 7704
rect 3142 7692 3148 7704
rect 3200 7732 3206 7744
rect 3329 7735 3387 7741
rect 3329 7732 3341 7735
rect 3200 7704 3341 7732
rect 3200 7692 3206 7704
rect 3329 7701 3341 7704
rect 3375 7701 3387 7735
rect 3329 7695 3387 7701
rect 3418 7692 3424 7744
rect 3476 7692 3482 7744
rect 4246 7692 4252 7744
rect 4304 7692 4310 7744
rect 5169 7735 5227 7741
rect 5169 7701 5181 7735
rect 5215 7732 5227 7735
rect 5258 7732 5264 7744
rect 5215 7704 5264 7732
rect 5215 7701 5227 7704
rect 5169 7695 5227 7701
rect 5258 7692 5264 7704
rect 5316 7692 5322 7744
rect 5350 7692 5356 7744
rect 5408 7732 5414 7744
rect 5718 7732 5724 7744
rect 5408 7704 5724 7732
rect 5408 7692 5414 7704
rect 5718 7692 5724 7704
rect 5776 7692 5782 7744
rect 5994 7692 6000 7744
rect 6052 7692 6058 7744
rect 6086 7692 6092 7744
rect 6144 7732 6150 7744
rect 6730 7732 6736 7744
rect 6144 7704 6736 7732
rect 6144 7692 6150 7704
rect 6730 7692 6736 7704
rect 6788 7692 6794 7744
rect 7098 7692 7104 7744
rect 7156 7692 7162 7744
rect 8021 7735 8079 7741
rect 8021 7701 8033 7735
rect 8067 7732 8079 7735
rect 9950 7732 9956 7744
rect 8067 7704 9956 7732
rect 8067 7701 8079 7704
rect 8021 7695 8079 7701
rect 9950 7692 9956 7704
rect 10008 7732 10014 7744
rect 10980 7732 11008 7831
rect 11238 7828 11244 7840
rect 11296 7828 11302 7880
rect 11790 7877 11796 7880
rect 11784 7868 11796 7877
rect 11751 7840 11796 7868
rect 11784 7831 11796 7840
rect 11790 7828 11796 7831
rect 11848 7828 11854 7880
rect 12894 7828 12900 7880
rect 12952 7868 12958 7880
rect 13265 7871 13323 7877
rect 13265 7868 13277 7871
rect 12952 7840 13277 7868
rect 12952 7828 12958 7840
rect 13265 7837 13277 7840
rect 13311 7868 13323 7871
rect 13538 7868 13544 7880
rect 13311 7840 13544 7868
rect 13311 7837 13323 7840
rect 13265 7831 13323 7837
rect 13538 7828 13544 7840
rect 13596 7828 13602 7880
rect 13630 7828 13636 7880
rect 13688 7828 13694 7880
rect 13722 7828 13728 7880
rect 13780 7868 13786 7880
rect 13998 7868 14004 7880
rect 13780 7840 14004 7868
rect 13780 7828 13786 7840
rect 13998 7828 14004 7840
rect 14056 7868 14062 7880
rect 14093 7871 14151 7877
rect 14093 7868 14105 7871
rect 14056 7840 14105 7868
rect 14056 7828 14062 7840
rect 14093 7837 14105 7840
rect 14139 7837 14151 7871
rect 14093 7831 14151 7837
rect 14274 7828 14280 7880
rect 14332 7828 14338 7880
rect 14366 7828 14372 7880
rect 14424 7828 14430 7880
rect 14458 7828 14464 7880
rect 14516 7828 14522 7880
rect 15194 7877 15200 7880
rect 15188 7868 15200 7877
rect 15155 7840 15200 7868
rect 15188 7831 15200 7840
rect 15194 7828 15200 7831
rect 15252 7828 15258 7880
rect 12158 7760 12164 7812
rect 12216 7800 12222 7812
rect 14384 7800 14412 7828
rect 15102 7800 15108 7812
rect 12216 7772 13124 7800
rect 14384 7772 15108 7800
rect 12216 7760 12222 7772
rect 13096 7741 13124 7772
rect 15102 7760 15108 7772
rect 15160 7760 15166 7812
rect 10008 7704 11008 7732
rect 13081 7735 13139 7741
rect 10008 7692 10014 7704
rect 13081 7701 13093 7735
rect 13127 7701 13139 7735
rect 13081 7695 13139 7701
rect 14734 7692 14740 7744
rect 14792 7692 14798 7744
rect 14826 7692 14832 7744
rect 14884 7732 14890 7744
rect 15010 7732 15016 7744
rect 14884 7704 15016 7732
rect 14884 7692 14890 7704
rect 15010 7692 15016 7704
rect 15068 7732 15074 7744
rect 16298 7732 16304 7744
rect 15068 7704 16304 7732
rect 15068 7692 15074 7704
rect 16298 7692 16304 7704
rect 16356 7692 16362 7744
rect 1104 7642 16652 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 16652 7642
rect 1104 7568 16652 7590
rect 2958 7528 2964 7540
rect 1412 7500 2964 7528
rect 1412 7401 1440 7500
rect 2958 7488 2964 7500
rect 3016 7488 3022 7540
rect 3050 7488 3056 7540
rect 3108 7488 3114 7540
rect 3145 7531 3203 7537
rect 3145 7497 3157 7531
rect 3191 7497 3203 7531
rect 3145 7491 3203 7497
rect 3313 7531 3371 7537
rect 3313 7497 3325 7531
rect 3359 7528 3371 7531
rect 4246 7528 4252 7540
rect 3359 7500 4252 7528
rect 3359 7497 3371 7500
rect 3313 7491 3371 7497
rect 1486 7420 1492 7472
rect 1544 7420 1550 7472
rect 1940 7463 1998 7469
rect 1940 7429 1952 7463
rect 1986 7460 1998 7463
rect 3160 7460 3188 7491
rect 4246 7488 4252 7500
rect 4304 7488 4310 7540
rect 4706 7488 4712 7540
rect 4764 7488 4770 7540
rect 6086 7528 6092 7540
rect 4908 7500 6092 7528
rect 1986 7432 3188 7460
rect 3513 7463 3571 7469
rect 1986 7429 1998 7432
rect 1940 7423 1998 7429
rect 3513 7429 3525 7463
rect 3559 7429 3571 7463
rect 3513 7423 3571 7429
rect 4617 7463 4675 7469
rect 4617 7429 4629 7463
rect 4663 7460 4675 7463
rect 4908 7460 4936 7500
rect 6086 7488 6092 7500
rect 6144 7488 6150 7540
rect 6178 7488 6184 7540
rect 6236 7488 6242 7540
rect 8113 7531 8171 7537
rect 8113 7497 8125 7531
rect 8159 7528 8171 7531
rect 8478 7528 8484 7540
rect 8159 7500 8484 7528
rect 8159 7497 8171 7500
rect 8113 7491 8171 7497
rect 8478 7488 8484 7500
rect 8536 7488 8542 7540
rect 9582 7528 9588 7540
rect 8588 7500 9588 7528
rect 8588 7460 8616 7500
rect 9582 7488 9588 7500
rect 9640 7488 9646 7540
rect 11330 7488 11336 7540
rect 11388 7528 11394 7540
rect 13630 7528 13636 7540
rect 11388 7500 13636 7528
rect 11388 7488 11394 7500
rect 13630 7488 13636 7500
rect 13688 7488 13694 7540
rect 16206 7488 16212 7540
rect 16264 7488 16270 7540
rect 9858 7460 9864 7472
rect 4663 7432 4936 7460
rect 5000 7432 5672 7460
rect 4663 7429 4675 7432
rect 4617 7423 4675 7429
rect 1397 7395 1455 7401
rect 1397 7361 1409 7395
rect 1443 7361 1455 7395
rect 1397 7355 1455 7361
rect 1578 7352 1584 7404
rect 1636 7352 1642 7404
rect 1670 7352 1676 7404
rect 1728 7352 1734 7404
rect 2222 7352 2228 7404
rect 2280 7392 2286 7404
rect 3528 7392 3556 7423
rect 3697 7395 3755 7401
rect 3697 7392 3709 7395
rect 2280 7364 3709 7392
rect 2280 7352 2286 7364
rect 3697 7361 3709 7364
rect 3743 7361 3755 7395
rect 3697 7355 3755 7361
rect 3881 7395 3939 7401
rect 3881 7361 3893 7395
rect 3927 7361 3939 7395
rect 3881 7355 3939 7361
rect 3896 7324 3924 7355
rect 3970 7352 3976 7404
rect 4028 7352 4034 7404
rect 4062 7352 4068 7404
rect 4120 7352 4126 7404
rect 4433 7395 4491 7401
rect 4433 7361 4445 7395
rect 4479 7361 4491 7395
rect 4433 7355 4491 7361
rect 3344 7296 3924 7324
rect 4448 7324 4476 7355
rect 4706 7352 4712 7404
rect 4764 7352 4770 7404
rect 4801 7395 4859 7401
rect 4801 7361 4813 7395
rect 4847 7392 4859 7395
rect 5000 7392 5028 7432
rect 5644 7404 5672 7432
rect 7852 7432 8616 7460
rect 9048 7432 9864 7460
rect 4847 7364 5028 7392
rect 5068 7395 5126 7401
rect 4847 7361 4859 7364
rect 4801 7355 4859 7361
rect 5068 7361 5080 7395
rect 5114 7392 5126 7395
rect 5350 7392 5356 7404
rect 5114 7364 5356 7392
rect 5114 7361 5126 7364
rect 5068 7355 5126 7361
rect 5350 7352 5356 7364
rect 5408 7352 5414 7404
rect 5626 7352 5632 7404
rect 5684 7392 5690 7404
rect 6362 7392 6368 7404
rect 5684 7364 6368 7392
rect 5684 7352 5690 7364
rect 6362 7352 6368 7364
rect 6420 7352 6426 7404
rect 6632 7395 6690 7401
rect 6632 7361 6644 7395
rect 6678 7392 6690 7395
rect 7006 7392 7012 7404
rect 6678 7364 7012 7392
rect 6678 7361 6690 7364
rect 6632 7355 6690 7361
rect 7006 7352 7012 7364
rect 7064 7352 7070 7404
rect 7852 7401 7880 7432
rect 7837 7395 7895 7401
rect 7837 7361 7849 7395
rect 7883 7361 7895 7395
rect 7837 7355 7895 7361
rect 7929 7395 7987 7401
rect 7929 7361 7941 7395
rect 7975 7392 7987 7395
rect 8294 7392 8300 7404
rect 7975 7364 8300 7392
rect 7975 7361 7987 7364
rect 7929 7355 7987 7361
rect 8294 7352 8300 7364
rect 8352 7352 8358 7404
rect 8389 7395 8447 7401
rect 8389 7361 8401 7395
rect 8435 7392 8447 7395
rect 8754 7392 8760 7404
rect 8435 7364 8760 7392
rect 8435 7361 8447 7364
rect 8389 7355 8447 7361
rect 8754 7352 8760 7364
rect 8812 7352 8818 7404
rect 9048 7401 9076 7432
rect 9858 7420 9864 7432
rect 9916 7420 9922 7472
rect 12526 7460 12532 7472
rect 11532 7432 12532 7460
rect 9033 7395 9091 7401
rect 9033 7361 9045 7395
rect 9079 7361 9091 7395
rect 9289 7395 9347 7401
rect 9289 7392 9301 7395
rect 9033 7355 9091 7361
rect 9140 7364 9301 7392
rect 8113 7327 8171 7333
rect 4448 7296 4844 7324
rect 1946 7148 1952 7200
rect 2004 7188 2010 7200
rect 2314 7188 2320 7200
rect 2004 7160 2320 7188
rect 2004 7148 2010 7160
rect 2314 7148 2320 7160
rect 2372 7188 2378 7200
rect 3344 7197 3372 7296
rect 4341 7259 4399 7265
rect 4341 7225 4353 7259
rect 4387 7256 4399 7259
rect 4614 7256 4620 7268
rect 4387 7228 4620 7256
rect 4387 7225 4399 7228
rect 4341 7219 4399 7225
rect 4614 7216 4620 7228
rect 4672 7216 4678 7268
rect 3329 7191 3387 7197
rect 3329 7188 3341 7191
rect 2372 7160 3341 7188
rect 2372 7148 2378 7160
rect 3329 7157 3341 7160
rect 3375 7157 3387 7191
rect 4816 7188 4844 7296
rect 8113 7293 8125 7327
rect 8159 7324 8171 7327
rect 8202 7324 8208 7336
rect 8159 7296 8208 7324
rect 8159 7293 8171 7296
rect 8113 7287 8171 7293
rect 8202 7284 8208 7296
rect 8260 7284 8266 7336
rect 8481 7327 8539 7333
rect 8481 7293 8493 7327
rect 8527 7324 8539 7327
rect 8662 7324 8668 7336
rect 8527 7296 8668 7324
rect 8527 7293 8539 7296
rect 8481 7287 8539 7293
rect 8662 7284 8668 7296
rect 8720 7284 8726 7336
rect 9140 7324 9168 7364
rect 9289 7361 9301 7364
rect 9335 7361 9347 7395
rect 9289 7355 9347 7361
rect 9674 7352 9680 7404
rect 9732 7392 9738 7404
rect 10505 7395 10563 7401
rect 10505 7392 10517 7395
rect 9732 7364 10517 7392
rect 9732 7352 9738 7364
rect 10505 7361 10517 7364
rect 10551 7361 10563 7395
rect 10505 7355 10563 7361
rect 11146 7352 11152 7404
rect 11204 7352 11210 7404
rect 11532 7401 11560 7432
rect 12526 7420 12532 7432
rect 12584 7460 12590 7472
rect 12584 7432 13124 7460
rect 12584 7420 12590 7432
rect 11517 7395 11575 7401
rect 11517 7361 11529 7395
rect 11563 7361 11575 7395
rect 11517 7355 11575 7361
rect 11606 7352 11612 7404
rect 11664 7392 11670 7404
rect 13096 7401 13124 7432
rect 14918 7420 14924 7472
rect 14976 7460 14982 7472
rect 14976 7432 15976 7460
rect 14976 7420 14982 7432
rect 11773 7395 11831 7401
rect 11773 7392 11785 7395
rect 11664 7364 11785 7392
rect 11664 7352 11670 7364
rect 11773 7361 11785 7364
rect 11819 7361 11831 7395
rect 11773 7355 11831 7361
rect 13081 7395 13139 7401
rect 13081 7361 13093 7395
rect 13127 7361 13139 7395
rect 13081 7355 13139 7361
rect 13170 7352 13176 7404
rect 13228 7392 13234 7404
rect 13337 7395 13395 7401
rect 13337 7392 13349 7395
rect 13228 7364 13349 7392
rect 13228 7352 13234 7364
rect 13337 7361 13349 7364
rect 13383 7361 13395 7395
rect 13337 7355 13395 7361
rect 14734 7352 14740 7404
rect 14792 7392 14798 7404
rect 15948 7401 15976 7432
rect 15666 7395 15724 7401
rect 15666 7392 15678 7395
rect 14792 7364 15678 7392
rect 14792 7352 14798 7364
rect 15666 7361 15678 7364
rect 15712 7361 15724 7395
rect 15666 7355 15724 7361
rect 15933 7395 15991 7401
rect 15933 7361 15945 7395
rect 15979 7361 15991 7395
rect 15933 7355 15991 7361
rect 16022 7352 16028 7404
rect 16080 7352 16086 7404
rect 8772 7296 9168 7324
rect 8772 7265 8800 7296
rect 8757 7259 8815 7265
rect 8757 7225 8769 7259
rect 8803 7225 8815 7259
rect 8757 7219 8815 7225
rect 12897 7259 12955 7265
rect 12897 7225 12909 7259
rect 12943 7256 12955 7259
rect 12986 7256 12992 7268
rect 12943 7228 12992 7256
rect 12943 7225 12955 7228
rect 12897 7219 12955 7225
rect 12986 7216 12992 7228
rect 13044 7216 13050 7268
rect 5994 7188 6000 7200
rect 4816 7160 6000 7188
rect 3329 7151 3387 7157
rect 5994 7148 6000 7160
rect 6052 7188 6058 7200
rect 6638 7188 6644 7200
rect 6052 7160 6644 7188
rect 6052 7148 6058 7160
rect 6638 7148 6644 7160
rect 6696 7188 6702 7200
rect 7745 7191 7803 7197
rect 7745 7188 7757 7191
rect 6696 7160 7757 7188
rect 6696 7148 6702 7160
rect 7745 7157 7757 7160
rect 7791 7188 7803 7191
rect 8018 7188 8024 7200
rect 7791 7160 8024 7188
rect 7791 7157 7803 7160
rect 7745 7151 7803 7157
rect 8018 7148 8024 7160
rect 8076 7148 8082 7200
rect 10410 7148 10416 7200
rect 10468 7188 10474 7200
rect 10778 7188 10784 7200
rect 10468 7160 10784 7188
rect 10468 7148 10474 7160
rect 10778 7148 10784 7160
rect 10836 7148 10842 7200
rect 13998 7148 14004 7200
rect 14056 7188 14062 7200
rect 14461 7191 14519 7197
rect 14461 7188 14473 7191
rect 14056 7160 14473 7188
rect 14056 7148 14062 7160
rect 14461 7157 14473 7160
rect 14507 7157 14519 7191
rect 14461 7151 14519 7157
rect 14550 7148 14556 7200
rect 14608 7148 14614 7200
rect 1104 7098 16652 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 16652 7098
rect 1104 7024 16652 7046
rect 2314 6944 2320 6996
rect 2372 6984 2378 6996
rect 2961 6987 3019 6993
rect 2961 6984 2973 6987
rect 2372 6956 2973 6984
rect 2372 6944 2378 6956
rect 2961 6953 2973 6956
rect 3007 6953 3019 6987
rect 2961 6947 3019 6953
rect 2406 6916 2412 6928
rect 1780 6888 2412 6916
rect 1780 6857 1808 6888
rect 2406 6876 2412 6888
rect 2464 6876 2470 6928
rect 2976 6916 3004 6947
rect 3142 6944 3148 6996
rect 3200 6944 3206 6996
rect 3418 6944 3424 6996
rect 3476 6944 3482 6996
rect 4798 6984 4804 6996
rect 3528 6956 4804 6984
rect 3528 6916 3556 6956
rect 4798 6944 4804 6956
rect 4856 6944 4862 6996
rect 5166 6944 5172 6996
rect 5224 6944 5230 6996
rect 5718 6944 5724 6996
rect 5776 6984 5782 6996
rect 6178 6984 6184 6996
rect 5776 6956 6184 6984
rect 5776 6944 5782 6956
rect 6178 6944 6184 6956
rect 6236 6984 6242 6996
rect 6236 6956 6684 6984
rect 6236 6944 6242 6956
rect 2976 6888 3556 6916
rect 6656 6916 6684 6956
rect 6730 6944 6736 6996
rect 6788 6984 6794 6996
rect 6917 6987 6975 6993
rect 6917 6984 6929 6987
rect 6788 6956 6929 6984
rect 6788 6944 6794 6956
rect 6917 6953 6929 6956
rect 6963 6953 6975 6987
rect 6917 6947 6975 6953
rect 7006 6944 7012 6996
rect 7064 6944 7070 6996
rect 7193 6987 7251 6993
rect 7193 6953 7205 6987
rect 7239 6953 7251 6987
rect 7193 6947 7251 6953
rect 7208 6916 7236 6947
rect 11330 6944 11336 6996
rect 11388 6944 11394 6996
rect 11517 6987 11575 6993
rect 11517 6953 11529 6987
rect 11563 6984 11575 6987
rect 11606 6984 11612 6996
rect 11563 6956 11612 6984
rect 11563 6953 11575 6956
rect 11517 6947 11575 6953
rect 11606 6944 11612 6956
rect 11664 6944 11670 6996
rect 12989 6987 13047 6993
rect 12989 6953 13001 6987
rect 13035 6984 13047 6987
rect 13170 6984 13176 6996
rect 13035 6956 13176 6984
rect 13035 6953 13047 6956
rect 12989 6947 13047 6953
rect 13170 6944 13176 6956
rect 13228 6944 13234 6996
rect 14458 6944 14464 6996
rect 14516 6984 14522 6996
rect 14645 6987 14703 6993
rect 14645 6984 14657 6987
rect 14516 6956 14657 6984
rect 14516 6944 14522 6956
rect 14645 6953 14657 6956
rect 14691 6953 14703 6987
rect 14645 6947 14703 6953
rect 6656 6888 7236 6916
rect 1765 6851 1823 6857
rect 1765 6817 1777 6851
rect 1811 6817 1823 6851
rect 1765 6811 1823 6817
rect 2041 6851 2099 6857
rect 2041 6817 2053 6851
rect 2087 6848 2099 6851
rect 2314 6848 2320 6860
rect 2087 6820 2320 6848
rect 2087 6817 2099 6820
rect 2041 6811 2099 6817
rect 2314 6808 2320 6820
rect 2372 6808 2378 6860
rect 2774 6808 2780 6860
rect 2832 6848 2838 6860
rect 3234 6848 3240 6860
rect 2832 6820 3240 6848
rect 2832 6808 2838 6820
rect 3234 6808 3240 6820
rect 3292 6848 3298 6860
rect 3789 6851 3847 6857
rect 3789 6848 3801 6851
rect 3292 6820 3801 6848
rect 3292 6808 3298 6820
rect 3789 6817 3801 6820
rect 3835 6817 3847 6851
rect 3789 6811 3847 6817
rect 9122 6808 9128 6860
rect 9180 6848 9186 6860
rect 9217 6851 9275 6857
rect 9217 6848 9229 6851
rect 9180 6820 9229 6848
rect 9180 6808 9186 6820
rect 9217 6817 9229 6820
rect 9263 6817 9275 6851
rect 9217 6811 9275 6817
rect 10597 6851 10655 6857
rect 10597 6817 10609 6851
rect 10643 6848 10655 6851
rect 11054 6848 11060 6860
rect 10643 6820 11060 6848
rect 10643 6817 10655 6820
rect 10597 6811 10655 6817
rect 11054 6808 11060 6820
rect 11112 6848 11118 6860
rect 11174 6851 11232 6857
rect 11174 6848 11186 6851
rect 11112 6820 11186 6848
rect 11112 6808 11118 6820
rect 11174 6817 11186 6820
rect 11220 6817 11232 6851
rect 11174 6811 11232 6817
rect 12158 6808 12164 6860
rect 12216 6808 12222 6860
rect 14918 6808 14924 6860
rect 14976 6808 14982 6860
rect 1673 6783 1731 6789
rect 1673 6749 1685 6783
rect 1719 6780 1731 6783
rect 2866 6780 2872 6792
rect 1719 6752 2872 6780
rect 1719 6749 1731 6752
rect 1673 6743 1731 6749
rect 2866 6740 2872 6752
rect 2924 6740 2930 6792
rect 3878 6780 3884 6792
rect 3278 6752 3884 6780
rect 3278 6746 3306 6752
rect 2133 6715 2191 6721
rect 2133 6681 2145 6715
rect 2179 6712 2191 6715
rect 2222 6712 2228 6724
rect 2179 6684 2228 6712
rect 2179 6681 2191 6684
rect 2133 6675 2191 6681
rect 2222 6672 2228 6684
rect 2280 6672 2286 6724
rect 2314 6672 2320 6724
rect 2372 6721 2378 6724
rect 2372 6715 2391 6721
rect 2379 6681 2391 6715
rect 2682 6712 2688 6724
rect 2372 6675 2391 6681
rect 2424 6684 2688 6712
rect 2372 6672 2378 6675
rect 2240 6644 2268 6672
rect 2424 6644 2452 6684
rect 2682 6672 2688 6684
rect 2740 6712 2746 6724
rect 2777 6715 2835 6721
rect 2777 6712 2789 6715
rect 2740 6684 2789 6712
rect 2740 6672 2746 6684
rect 2777 6681 2789 6684
rect 2823 6681 2835 6715
rect 2777 6675 2835 6681
rect 2958 6672 2964 6724
rect 3016 6721 3022 6724
rect 3252 6721 3306 6746
rect 3878 6740 3884 6752
rect 3936 6740 3942 6792
rect 4056 6783 4114 6789
rect 4056 6749 4068 6783
rect 4102 6780 4114 6783
rect 4614 6780 4620 6792
rect 4102 6752 4620 6780
rect 4102 6749 4114 6752
rect 4056 6743 4114 6749
rect 4614 6740 4620 6752
rect 4672 6740 4678 6792
rect 5261 6783 5319 6789
rect 5261 6780 5273 6783
rect 4908 6752 5273 6780
rect 3016 6715 3035 6721
rect 3023 6681 3035 6715
rect 3016 6675 3035 6681
rect 3237 6718 3306 6721
rect 3237 6715 3295 6718
rect 3237 6681 3249 6715
rect 3283 6681 3295 6715
rect 3237 6675 3295 6681
rect 3016 6672 3022 6675
rect 2240 6616 2452 6644
rect 2498 6604 2504 6656
rect 2556 6604 2562 6656
rect 2590 6604 2596 6656
rect 2648 6644 2654 6656
rect 2866 6644 2872 6656
rect 2648 6616 2872 6644
rect 2648 6604 2654 6616
rect 2866 6604 2872 6616
rect 2924 6644 2930 6656
rect 3437 6647 3495 6653
rect 3437 6644 3449 6647
rect 2924 6616 3449 6644
rect 2924 6604 2930 6616
rect 3437 6613 3449 6616
rect 3483 6613 3495 6647
rect 3437 6607 3495 6613
rect 3605 6647 3663 6653
rect 3605 6613 3617 6647
rect 3651 6644 3663 6647
rect 3970 6644 3976 6656
rect 3651 6616 3976 6644
rect 3651 6613 3663 6616
rect 3605 6607 3663 6613
rect 3970 6604 3976 6616
rect 4028 6644 4034 6656
rect 4908 6644 4936 6752
rect 5261 6749 5273 6752
rect 5307 6749 5319 6783
rect 5261 6743 5319 6749
rect 5442 6740 5448 6792
rect 5500 6740 5506 6792
rect 5537 6783 5595 6789
rect 5537 6749 5549 6783
rect 5583 6780 5595 6783
rect 5626 6780 5632 6792
rect 5583 6752 5632 6780
rect 5583 6749 5595 6752
rect 5537 6743 5595 6749
rect 5626 6740 5632 6752
rect 5684 6740 5690 6792
rect 6914 6740 6920 6792
rect 6972 6780 6978 6792
rect 7837 6783 7895 6789
rect 7837 6780 7849 6783
rect 6972 6752 7849 6780
rect 6972 6740 6978 6752
rect 7837 6749 7849 6752
rect 7883 6749 7895 6783
rect 7837 6743 7895 6749
rect 8018 6740 8024 6792
rect 8076 6740 8082 6792
rect 9861 6783 9919 6789
rect 9861 6749 9873 6783
rect 9907 6749 9919 6783
rect 9861 6743 9919 6749
rect 5350 6672 5356 6724
rect 5408 6672 5414 6724
rect 5804 6715 5862 6721
rect 5804 6681 5816 6715
rect 5850 6712 5862 6715
rect 5902 6712 5908 6724
rect 5850 6684 5908 6712
rect 5850 6681 5862 6684
rect 5804 6675 5862 6681
rect 5902 6672 5908 6684
rect 5960 6672 5966 6724
rect 7098 6672 7104 6724
rect 7156 6721 7162 6724
rect 7156 6715 7219 6721
rect 7156 6681 7173 6715
rect 7207 6681 7219 6715
rect 7156 6675 7219 6681
rect 7377 6715 7435 6721
rect 7377 6681 7389 6715
rect 7423 6712 7435 6715
rect 7929 6715 7987 6721
rect 7929 6712 7941 6715
rect 7423 6684 7941 6712
rect 7423 6681 7435 6684
rect 7377 6675 7435 6681
rect 7929 6681 7941 6684
rect 7975 6681 7987 6715
rect 9876 6712 9904 6743
rect 10686 6740 10692 6792
rect 10744 6740 10750 6792
rect 10778 6740 10784 6792
rect 10836 6780 10842 6792
rect 10965 6783 11023 6789
rect 10965 6780 10977 6783
rect 10836 6752 10977 6780
rect 10836 6740 10842 6752
rect 10965 6749 10977 6752
rect 11011 6749 11023 6783
rect 10965 6743 11023 6749
rect 12618 6740 12624 6792
rect 12676 6780 12682 6792
rect 12897 6783 12955 6789
rect 12897 6780 12909 6783
rect 12676 6752 12909 6780
rect 12676 6740 12682 6752
rect 12897 6749 12909 6752
rect 12943 6749 12955 6783
rect 12897 6743 12955 6749
rect 13262 6740 13268 6792
rect 13320 6740 13326 6792
rect 13354 6740 13360 6792
rect 13412 6740 13418 6792
rect 13449 6783 13507 6789
rect 13449 6749 13461 6783
rect 13495 6780 13507 6783
rect 13538 6780 13544 6792
rect 13495 6752 13544 6780
rect 13495 6749 13507 6752
rect 13449 6743 13507 6749
rect 13538 6740 13544 6752
rect 13596 6740 13602 6792
rect 13633 6783 13691 6789
rect 13633 6749 13645 6783
rect 13679 6780 13691 6783
rect 13722 6780 13728 6792
rect 13679 6752 13728 6780
rect 13679 6749 13691 6752
rect 13633 6743 13691 6749
rect 13722 6740 13728 6752
rect 13780 6740 13786 6792
rect 13998 6740 14004 6792
rect 14056 6780 14062 6792
rect 14093 6783 14151 6789
rect 14093 6780 14105 6783
rect 14056 6752 14105 6780
rect 14056 6740 14062 6752
rect 14093 6749 14105 6752
rect 14139 6749 14151 6783
rect 14093 6743 14151 6749
rect 14182 6740 14188 6792
rect 14240 6780 14246 6792
rect 14277 6783 14335 6789
rect 14277 6780 14289 6783
rect 14240 6752 14289 6780
rect 14240 6740 14246 6752
rect 14277 6749 14289 6752
rect 14323 6749 14335 6783
rect 14277 6743 14335 6749
rect 14461 6783 14519 6789
rect 14461 6749 14473 6783
rect 14507 6780 14519 6783
rect 14642 6780 14648 6792
rect 14507 6752 14648 6780
rect 14507 6749 14519 6752
rect 14461 6743 14519 6749
rect 14642 6740 14648 6752
rect 14700 6740 14706 6792
rect 11057 6715 11115 6721
rect 11057 6712 11069 6715
rect 9876 6684 11069 6712
rect 7929 6675 7987 6681
rect 11057 6681 11069 6684
rect 11103 6712 11115 6715
rect 11146 6712 11152 6724
rect 11103 6684 11152 6712
rect 11103 6681 11115 6684
rect 11057 6675 11115 6681
rect 7156 6672 7162 6675
rect 11146 6672 11152 6684
rect 11204 6672 11210 6724
rect 11977 6715 12035 6721
rect 11977 6681 11989 6715
rect 12023 6712 12035 6715
rect 12986 6712 12992 6724
rect 12023 6684 12992 6712
rect 12023 6681 12035 6684
rect 11977 6675 12035 6681
rect 12986 6672 12992 6684
rect 13044 6672 13050 6724
rect 14366 6672 14372 6724
rect 14424 6712 14430 6724
rect 14550 6712 14556 6724
rect 14424 6684 14556 6712
rect 14424 6672 14430 6684
rect 14550 6672 14556 6684
rect 14608 6672 14614 6724
rect 15188 6715 15246 6721
rect 15188 6681 15200 6715
rect 15234 6712 15246 6715
rect 15562 6712 15568 6724
rect 15234 6684 15568 6712
rect 15234 6681 15246 6684
rect 15188 6675 15246 6681
rect 15562 6672 15568 6684
rect 15620 6672 15626 6724
rect 4028 6616 4936 6644
rect 9953 6647 10011 6653
rect 4028 6604 4034 6616
rect 9953 6613 9965 6647
rect 9999 6644 10011 6647
rect 10042 6644 10048 6656
rect 9999 6616 10048 6644
rect 9999 6613 10011 6616
rect 9953 6607 10011 6613
rect 10042 6604 10048 6616
rect 10100 6604 10106 6656
rect 11882 6604 11888 6656
rect 11940 6604 11946 6656
rect 12713 6647 12771 6653
rect 12713 6613 12725 6647
rect 12759 6644 12771 6647
rect 13170 6644 13176 6656
rect 12759 6616 13176 6644
rect 12759 6613 12771 6616
rect 12713 6607 12771 6613
rect 13170 6604 13176 6616
rect 13228 6604 13234 6656
rect 13630 6604 13636 6656
rect 13688 6644 13694 6656
rect 14458 6644 14464 6656
rect 13688 6616 14464 6644
rect 13688 6604 13694 6616
rect 14458 6604 14464 6616
rect 14516 6644 14522 6656
rect 15930 6644 15936 6656
rect 14516 6616 15936 6644
rect 14516 6604 14522 6616
rect 15930 6604 15936 6616
rect 15988 6604 15994 6656
rect 16206 6604 16212 6656
rect 16264 6644 16270 6656
rect 16301 6647 16359 6653
rect 16301 6644 16313 6647
rect 16264 6616 16313 6644
rect 16264 6604 16270 6616
rect 16301 6613 16313 6616
rect 16347 6613 16359 6647
rect 16301 6607 16359 6613
rect 1104 6554 16652 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 16652 6554
rect 1104 6480 16652 6502
rect 3878 6440 3884 6452
rect 3084 6412 3884 6440
rect 2777 6307 2835 6313
rect 2777 6273 2789 6307
rect 2823 6304 2835 6307
rect 3084 6304 3112 6412
rect 3878 6400 3884 6412
rect 3936 6400 3942 6452
rect 5534 6400 5540 6452
rect 5592 6440 5598 6452
rect 6365 6443 6423 6449
rect 6365 6440 6377 6443
rect 5592 6412 6377 6440
rect 5592 6400 5598 6412
rect 6365 6409 6377 6412
rect 6411 6409 6423 6443
rect 6365 6403 6423 6409
rect 6733 6443 6791 6449
rect 6733 6409 6745 6443
rect 6779 6440 6791 6443
rect 6914 6440 6920 6452
rect 6779 6412 6920 6440
rect 6779 6409 6791 6412
rect 6733 6403 6791 6409
rect 3142 6332 3148 6384
rect 3200 6372 3206 6384
rect 3482 6375 3540 6381
rect 3482 6372 3494 6375
rect 3200 6344 3494 6372
rect 3200 6332 3206 6344
rect 3482 6341 3494 6344
rect 3528 6341 3540 6375
rect 4861 6375 4919 6381
rect 4861 6372 4873 6375
rect 3482 6335 3540 6341
rect 3620 6344 4873 6372
rect 2823 6276 3112 6304
rect 2823 6273 2835 6276
rect 2777 6267 2835 6273
rect 3234 6264 3240 6316
rect 3292 6264 3298 6316
rect 3620 6304 3648 6344
rect 4861 6341 4873 6344
rect 4907 6341 4919 6375
rect 4861 6335 4919 6341
rect 5077 6375 5135 6381
rect 5077 6341 5089 6375
rect 5123 6341 5135 6375
rect 5077 6335 5135 6341
rect 5905 6375 5963 6381
rect 5905 6341 5917 6375
rect 5951 6372 5963 6375
rect 6748 6372 6776 6403
rect 6914 6400 6920 6412
rect 6972 6400 6978 6452
rect 8846 6400 8852 6452
rect 8904 6440 8910 6452
rect 9493 6443 9551 6449
rect 9493 6440 9505 6443
rect 8904 6412 9505 6440
rect 8904 6400 8910 6412
rect 9493 6409 9505 6412
rect 9539 6409 9551 6443
rect 9493 6403 9551 6409
rect 10321 6443 10379 6449
rect 10321 6409 10333 6443
rect 10367 6440 10379 6443
rect 10962 6440 10968 6452
rect 10367 6412 10968 6440
rect 10367 6409 10379 6412
rect 10321 6403 10379 6409
rect 10962 6400 10968 6412
rect 11020 6400 11026 6452
rect 11149 6443 11207 6449
rect 11149 6409 11161 6443
rect 11195 6440 11207 6443
rect 11238 6440 11244 6452
rect 11195 6412 11244 6440
rect 11195 6409 11207 6412
rect 11149 6403 11207 6409
rect 11238 6400 11244 6412
rect 11296 6400 11302 6452
rect 11333 6443 11391 6449
rect 11333 6409 11345 6443
rect 11379 6440 11391 6443
rect 11974 6440 11980 6452
rect 11379 6412 11980 6440
rect 11379 6409 11391 6412
rect 11333 6403 11391 6409
rect 11974 6400 11980 6412
rect 12032 6400 12038 6452
rect 12069 6443 12127 6449
rect 12069 6409 12081 6443
rect 12115 6440 12127 6443
rect 13078 6440 13084 6452
rect 12115 6412 13084 6440
rect 12115 6409 12127 6412
rect 12069 6403 12127 6409
rect 13078 6400 13084 6412
rect 13136 6400 13142 6452
rect 13538 6400 13544 6452
rect 13596 6400 13602 6452
rect 14093 6443 14151 6449
rect 14093 6409 14105 6443
rect 14139 6440 14151 6443
rect 14274 6440 14280 6452
rect 14139 6412 14280 6440
rect 14139 6409 14151 6412
rect 14093 6403 14151 6409
rect 14274 6400 14280 6412
rect 14332 6400 14338 6452
rect 14737 6443 14795 6449
rect 14737 6409 14749 6443
rect 14783 6440 14795 6443
rect 15194 6440 15200 6452
rect 14783 6412 15200 6440
rect 14783 6409 14795 6412
rect 14737 6403 14795 6409
rect 15194 6400 15200 6412
rect 15252 6400 15258 6452
rect 15562 6400 15568 6452
rect 15620 6400 15626 6452
rect 15654 6400 15660 6452
rect 15712 6400 15718 6452
rect 16022 6440 16028 6452
rect 15948 6412 16028 6440
rect 5951 6344 6776 6372
rect 10489 6375 10547 6381
rect 5951 6341 5963 6344
rect 5905 6335 5963 6341
rect 10489 6341 10501 6375
rect 10535 6372 10547 6375
rect 10689 6375 10747 6381
rect 10535 6344 10640 6372
rect 10535 6341 10547 6344
rect 10489 6335 10547 6341
rect 3344 6276 3648 6304
rect 2866 6196 2872 6248
rect 2924 6196 2930 6248
rect 3145 6239 3203 6245
rect 3145 6205 3157 6239
rect 3191 6236 3203 6239
rect 3344 6236 3372 6276
rect 4062 6264 4068 6316
rect 4120 6304 4126 6316
rect 5092 6304 5120 6335
rect 4120 6276 5120 6304
rect 6549 6307 6607 6313
rect 4120 6264 4126 6276
rect 6549 6273 6561 6307
rect 6595 6304 6607 6307
rect 6730 6304 6736 6316
rect 6595 6276 6736 6304
rect 6595 6273 6607 6276
rect 6549 6267 6607 6273
rect 6730 6264 6736 6276
rect 6788 6264 6794 6316
rect 6825 6307 6883 6313
rect 6825 6273 6837 6307
rect 6871 6273 6883 6307
rect 6825 6267 6883 6273
rect 9493 6307 9551 6313
rect 9493 6273 9505 6307
rect 9539 6273 9551 6307
rect 9493 6267 9551 6273
rect 3191 6208 3372 6236
rect 3191 6205 3203 6208
rect 3145 6199 3203 6205
rect 6638 6196 6644 6248
rect 6696 6236 6702 6248
rect 6840 6236 6868 6267
rect 6696 6208 6868 6236
rect 9508 6236 9536 6267
rect 9674 6264 9680 6316
rect 9732 6264 9738 6316
rect 9766 6264 9772 6316
rect 9824 6264 9830 6316
rect 9861 6307 9919 6313
rect 9861 6273 9873 6307
rect 9907 6304 9919 6307
rect 9950 6304 9956 6316
rect 9907 6276 9956 6304
rect 9907 6273 9919 6276
rect 9861 6267 9919 6273
rect 9950 6264 9956 6276
rect 10008 6264 10014 6316
rect 9784 6236 9812 6264
rect 9508 6208 9812 6236
rect 6696 6196 6702 6208
rect 10042 6196 10048 6248
rect 10100 6196 10106 6248
rect 10612 6236 10640 6344
rect 10689 6341 10701 6375
rect 10735 6341 10747 6375
rect 12894 6372 12900 6384
rect 10689 6335 10747 6341
rect 12406 6344 12900 6372
rect 10704 6304 10732 6335
rect 10781 6307 10839 6313
rect 10781 6304 10793 6307
rect 10704 6276 10793 6304
rect 10781 6273 10793 6276
rect 10827 6304 10839 6307
rect 11146 6304 11152 6316
rect 10827 6276 11152 6304
rect 10827 6273 10839 6276
rect 10781 6267 10839 6273
rect 11146 6264 11152 6276
rect 11204 6304 11210 6316
rect 11517 6307 11575 6313
rect 11517 6304 11529 6307
rect 11204 6276 11529 6304
rect 11204 6264 11210 6276
rect 11517 6273 11529 6276
rect 11563 6304 11575 6307
rect 12406 6304 12434 6344
rect 12894 6332 12900 6344
rect 12952 6332 12958 6384
rect 13004 6344 14320 6372
rect 13004 6313 13032 6344
rect 11563 6276 12434 6304
rect 12621 6307 12679 6313
rect 11563 6273 11575 6276
rect 11517 6267 11575 6273
rect 12621 6273 12633 6307
rect 12667 6304 12679 6307
rect 12989 6307 13047 6313
rect 12667 6276 12940 6304
rect 12667 6273 12679 6276
rect 12621 6267 12679 6273
rect 11054 6236 11060 6248
rect 10612 6208 11060 6236
rect 11054 6196 11060 6208
rect 11112 6236 11118 6248
rect 11238 6236 11244 6248
rect 11112 6208 11244 6236
rect 11112 6196 11118 6208
rect 11238 6196 11244 6208
rect 11296 6196 11302 6248
rect 11793 6239 11851 6245
rect 11793 6205 11805 6239
rect 11839 6205 11851 6239
rect 12912 6236 12940 6276
rect 12989 6273 13001 6307
rect 13035 6273 13047 6307
rect 12989 6267 13047 6273
rect 13265 6307 13323 6313
rect 13265 6273 13277 6307
rect 13311 6273 13323 6307
rect 13265 6267 13323 6273
rect 13449 6307 13507 6313
rect 13449 6273 13461 6307
rect 13495 6304 13507 6307
rect 13538 6304 13544 6316
rect 13495 6276 13544 6304
rect 13495 6273 13507 6276
rect 13449 6267 13507 6273
rect 13280 6236 13308 6267
rect 13538 6264 13544 6276
rect 13596 6264 13602 6316
rect 13725 6307 13783 6313
rect 13725 6273 13737 6307
rect 13771 6273 13783 6307
rect 13725 6267 13783 6273
rect 13630 6236 13636 6248
rect 12912 6208 13636 6236
rect 11793 6199 11851 6205
rect 5629 6171 5687 6177
rect 5629 6137 5641 6171
rect 5675 6168 5687 6171
rect 6178 6168 6184 6180
rect 5675 6140 6184 6168
rect 5675 6137 5687 6140
rect 5629 6131 5687 6137
rect 6178 6128 6184 6140
rect 6236 6128 6242 6180
rect 11808 6168 11836 6199
rect 13630 6196 13636 6208
rect 13688 6196 13694 6248
rect 13740 6236 13768 6267
rect 13906 6264 13912 6316
rect 13964 6264 13970 6316
rect 14292 6313 14320 6344
rect 14458 6332 14464 6384
rect 14516 6332 14522 6384
rect 14642 6332 14648 6384
rect 14700 6372 14706 6384
rect 15948 6381 15976 6412
rect 16022 6400 16028 6412
rect 16080 6400 16086 6452
rect 15933 6375 15991 6381
rect 14700 6344 15884 6372
rect 14700 6332 14706 6344
rect 14277 6307 14335 6313
rect 14277 6273 14289 6307
rect 14323 6304 14335 6307
rect 14366 6304 14372 6316
rect 14323 6276 14372 6304
rect 14323 6273 14335 6276
rect 14277 6267 14335 6273
rect 14366 6264 14372 6276
rect 14424 6264 14430 6316
rect 14550 6264 14556 6316
rect 14608 6264 14614 6316
rect 14921 6310 14979 6313
rect 15010 6310 15016 6314
rect 14921 6307 15016 6310
rect 14921 6273 14933 6307
rect 14967 6282 15016 6307
rect 14967 6273 14979 6282
rect 14921 6267 14979 6273
rect 15010 6262 15016 6282
rect 15068 6262 15074 6314
rect 15105 6310 15163 6316
rect 15203 6313 15209 6316
rect 15105 6276 15117 6310
rect 15151 6276 15163 6310
rect 15105 6270 15163 6276
rect 13998 6236 14004 6248
rect 13740 6208 14004 6236
rect 13998 6196 14004 6208
rect 14056 6196 14062 6248
rect 14090 6196 14096 6248
rect 14148 6236 14154 6248
rect 14148 6228 14780 6236
rect 15120 6228 15148 6270
rect 15200 6267 15209 6313
rect 15261 6304 15267 6316
rect 15335 6307 15393 6313
rect 15261 6276 15300 6304
rect 15203 6264 15209 6267
rect 15261 6264 15267 6276
rect 15335 6273 15347 6307
rect 15381 6304 15393 6307
rect 15746 6304 15752 6316
rect 15381 6276 15752 6304
rect 15381 6273 15393 6276
rect 15335 6267 15393 6273
rect 15746 6264 15752 6276
rect 15804 6264 15810 6316
rect 15856 6313 15884 6344
rect 15933 6341 15945 6375
rect 15979 6341 15991 6375
rect 15933 6335 15991 6341
rect 15841 6307 15899 6313
rect 15841 6273 15853 6307
rect 15887 6273 15899 6307
rect 15841 6267 15899 6273
rect 16022 6264 16028 6316
rect 16080 6264 16086 6316
rect 16206 6264 16212 6316
rect 16264 6264 16270 6316
rect 14148 6208 15148 6228
rect 14148 6196 14154 6208
rect 14752 6200 15148 6208
rect 11164 6140 11836 6168
rect 3418 6060 3424 6112
rect 3476 6100 3482 6112
rect 4617 6103 4675 6109
rect 4617 6100 4629 6103
rect 3476 6072 4629 6100
rect 3476 6060 3482 6072
rect 4617 6069 4629 6072
rect 4663 6069 4675 6103
rect 4617 6063 4675 6069
rect 4706 6060 4712 6112
rect 4764 6060 4770 6112
rect 4798 6060 4804 6112
rect 4856 6100 4862 6112
rect 4893 6103 4951 6109
rect 4893 6100 4905 6103
rect 4856 6072 4905 6100
rect 4856 6060 4862 6072
rect 4893 6069 4905 6072
rect 4939 6069 4951 6103
rect 4893 6063 4951 6069
rect 5442 6060 5448 6112
rect 5500 6060 5506 6112
rect 9950 6060 9956 6112
rect 10008 6060 10014 6112
rect 10505 6103 10563 6109
rect 10505 6069 10517 6103
rect 10551 6100 10563 6103
rect 10870 6100 10876 6112
rect 10551 6072 10876 6100
rect 10551 6069 10563 6072
rect 10505 6063 10563 6069
rect 10870 6060 10876 6072
rect 10928 6100 10934 6112
rect 11164 6109 11192 6140
rect 11149 6103 11207 6109
rect 11149 6100 11161 6103
rect 10928 6072 11161 6100
rect 10928 6060 10934 6072
rect 11149 6069 11161 6072
rect 11195 6069 11207 6103
rect 11149 6063 11207 6069
rect 11698 6060 11704 6112
rect 11756 6060 11762 6112
rect 11808 6100 11836 6140
rect 12437 6171 12495 6177
rect 12437 6137 12449 6171
rect 12483 6168 12495 6171
rect 15194 6168 15200 6180
rect 12483 6140 15200 6168
rect 12483 6137 12495 6140
rect 12437 6131 12495 6137
rect 15194 6128 15200 6140
rect 15252 6128 15258 6180
rect 12710 6100 12716 6112
rect 11808 6072 12716 6100
rect 12710 6060 12716 6072
rect 12768 6060 12774 6112
rect 12802 6060 12808 6112
rect 12860 6060 12866 6112
rect 13081 6103 13139 6109
rect 13081 6069 13093 6103
rect 13127 6100 13139 6103
rect 13722 6100 13728 6112
rect 13127 6072 13728 6100
rect 13127 6069 13139 6072
rect 13081 6063 13139 6069
rect 13722 6060 13728 6072
rect 13780 6060 13786 6112
rect 13814 6060 13820 6112
rect 13872 6100 13878 6112
rect 15010 6100 15016 6112
rect 13872 6072 15016 6100
rect 13872 6060 13878 6072
rect 15010 6060 15016 6072
rect 15068 6060 15074 6112
rect 1104 6010 16652 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 16652 6010
rect 1104 5936 16652 5958
rect 3789 5899 3847 5905
rect 3789 5865 3801 5899
rect 3835 5896 3847 5899
rect 3878 5896 3884 5908
rect 3835 5868 3884 5896
rect 3835 5865 3847 5868
rect 3789 5859 3847 5865
rect 3878 5856 3884 5868
rect 3936 5856 3942 5908
rect 6641 5899 6699 5905
rect 6641 5865 6653 5899
rect 6687 5896 6699 5899
rect 6914 5896 6920 5908
rect 6687 5868 6920 5896
rect 6687 5865 6699 5868
rect 6641 5859 6699 5865
rect 6914 5856 6920 5868
rect 6972 5856 6978 5908
rect 10594 5856 10600 5908
rect 10652 5856 10658 5908
rect 11977 5899 12035 5905
rect 11977 5865 11989 5899
rect 12023 5896 12035 5899
rect 12066 5896 12072 5908
rect 12023 5868 12072 5896
rect 12023 5865 12035 5868
rect 11977 5859 12035 5865
rect 12066 5856 12072 5868
rect 12124 5856 12130 5908
rect 12621 5899 12679 5905
rect 12621 5865 12633 5899
rect 12667 5896 12679 5899
rect 14090 5896 14096 5908
rect 12667 5868 14096 5896
rect 12667 5865 12679 5868
rect 12621 5859 12679 5865
rect 14090 5856 14096 5868
rect 14148 5856 14154 5908
rect 16022 5896 16028 5908
rect 15120 5868 16028 5896
rect 2682 5788 2688 5840
rect 2740 5828 2746 5840
rect 4062 5828 4068 5840
rect 2740 5800 4068 5828
rect 2740 5788 2746 5800
rect 4062 5788 4068 5800
rect 4120 5788 4126 5840
rect 14182 5788 14188 5840
rect 14240 5788 14246 5840
rect 14734 5788 14740 5840
rect 14792 5788 14798 5840
rect 13906 5760 13912 5772
rect 10704 5732 11376 5760
rect 5169 5695 5227 5701
rect 5169 5661 5181 5695
rect 5215 5692 5227 5695
rect 5261 5695 5319 5701
rect 5261 5692 5273 5695
rect 5215 5664 5273 5692
rect 5215 5661 5227 5664
rect 5169 5655 5227 5661
rect 5261 5661 5273 5664
rect 5307 5692 5319 5695
rect 5528 5695 5586 5701
rect 5307 5664 5396 5692
rect 5307 5661 5319 5664
rect 5261 5655 5319 5661
rect 4706 5584 4712 5636
rect 4764 5624 4770 5636
rect 4902 5627 4960 5633
rect 4902 5624 4914 5627
rect 4764 5596 4914 5624
rect 4764 5584 4770 5596
rect 4902 5593 4914 5596
rect 4948 5593 4960 5627
rect 4902 5587 4960 5593
rect 5368 5556 5396 5664
rect 5528 5661 5540 5695
rect 5574 5661 5586 5695
rect 5528 5655 5586 5661
rect 5442 5584 5448 5636
rect 5500 5624 5506 5636
rect 5552 5624 5580 5655
rect 9950 5652 9956 5704
rect 10008 5692 10014 5704
rect 10704 5701 10732 5732
rect 10505 5695 10563 5701
rect 10505 5692 10517 5695
rect 10008 5664 10517 5692
rect 10008 5652 10014 5664
rect 10505 5661 10517 5664
rect 10551 5661 10563 5695
rect 10505 5655 10563 5661
rect 10689 5695 10747 5701
rect 10689 5661 10701 5695
rect 10735 5661 10747 5695
rect 10689 5655 10747 5661
rect 10778 5652 10784 5704
rect 10836 5652 10842 5704
rect 10870 5652 10876 5704
rect 10928 5692 10934 5704
rect 11348 5701 11376 5732
rect 13096 5732 13912 5760
rect 10965 5695 11023 5701
rect 10965 5692 10977 5695
rect 10928 5664 10977 5692
rect 10928 5652 10934 5664
rect 10965 5661 10977 5664
rect 11011 5661 11023 5695
rect 10965 5655 11023 5661
rect 11333 5695 11391 5701
rect 11333 5661 11345 5695
rect 11379 5692 11391 5695
rect 11698 5692 11704 5704
rect 11379 5664 11704 5692
rect 11379 5661 11391 5664
rect 11333 5655 11391 5661
rect 11698 5652 11704 5664
rect 11756 5652 11762 5704
rect 12161 5695 12219 5701
rect 12161 5661 12173 5695
rect 12207 5692 12219 5695
rect 12250 5692 12256 5704
rect 12207 5664 12256 5692
rect 12207 5661 12219 5664
rect 12161 5655 12219 5661
rect 12250 5652 12256 5664
rect 12308 5652 12314 5704
rect 12529 5695 12587 5701
rect 12529 5661 12541 5695
rect 12575 5692 12587 5695
rect 12802 5692 12808 5704
rect 12575 5664 12808 5692
rect 12575 5661 12587 5664
rect 12529 5655 12587 5661
rect 12802 5652 12808 5664
rect 12860 5652 12866 5704
rect 13096 5636 13124 5732
rect 13906 5720 13912 5732
rect 13964 5720 13970 5772
rect 14200 5760 14228 5788
rect 15120 5760 15148 5868
rect 16022 5856 16028 5868
rect 16080 5856 16086 5908
rect 15286 5788 15292 5840
rect 15344 5788 15350 5840
rect 14200 5732 15148 5760
rect 15304 5760 15332 5788
rect 15304 5732 15884 5760
rect 13265 5695 13323 5701
rect 13265 5661 13277 5695
rect 13311 5692 13323 5695
rect 14093 5695 14151 5701
rect 14093 5692 14105 5695
rect 13311 5664 14105 5692
rect 13311 5661 13323 5664
rect 13265 5655 13323 5661
rect 14093 5661 14105 5664
rect 14139 5692 14151 5695
rect 14182 5692 14188 5704
rect 14139 5664 14188 5692
rect 14139 5661 14151 5664
rect 14093 5655 14151 5661
rect 14182 5652 14188 5664
rect 14240 5652 14246 5704
rect 14292 5701 14320 5732
rect 14277 5695 14335 5701
rect 14277 5661 14289 5695
rect 14323 5661 14335 5695
rect 14277 5655 14335 5661
rect 14369 5695 14427 5701
rect 14369 5661 14381 5695
rect 14415 5661 14427 5695
rect 14369 5655 14427 5661
rect 14461 5695 14519 5701
rect 14461 5661 14473 5695
rect 14507 5692 14519 5695
rect 14642 5692 14648 5704
rect 14507 5664 14648 5692
rect 14507 5661 14519 5664
rect 14461 5655 14519 5661
rect 5500 5596 5580 5624
rect 12989 5627 13047 5633
rect 5500 5584 5506 5596
rect 12989 5593 13001 5627
rect 13035 5624 13047 5627
rect 13078 5624 13084 5636
rect 13035 5596 13084 5624
rect 13035 5593 13047 5596
rect 12989 5587 13047 5593
rect 13078 5584 13084 5596
rect 13136 5584 13142 5636
rect 13538 5584 13544 5636
rect 13596 5584 13602 5636
rect 13725 5627 13783 5633
rect 13725 5593 13737 5627
rect 13771 5593 13783 5627
rect 13725 5587 13783 5593
rect 5534 5556 5540 5568
rect 5368 5528 5540 5556
rect 5534 5516 5540 5528
rect 5592 5516 5598 5568
rect 10873 5559 10931 5565
rect 10873 5525 10885 5559
rect 10919 5556 10931 5559
rect 10962 5556 10968 5568
rect 10919 5528 10968 5556
rect 10919 5525 10931 5528
rect 10873 5519 10931 5525
rect 10962 5516 10968 5528
rect 11020 5516 11026 5568
rect 11425 5559 11483 5565
rect 11425 5525 11437 5559
rect 11471 5556 11483 5559
rect 11514 5556 11520 5568
rect 11471 5528 11520 5556
rect 11471 5525 11483 5528
rect 11425 5519 11483 5525
rect 11514 5516 11520 5528
rect 11572 5516 11578 5568
rect 12342 5516 12348 5568
rect 12400 5516 12406 5568
rect 13449 5559 13507 5565
rect 13449 5525 13461 5559
rect 13495 5556 13507 5559
rect 13630 5556 13636 5568
rect 13495 5528 13636 5556
rect 13495 5525 13507 5528
rect 13449 5519 13507 5525
rect 13630 5516 13636 5528
rect 13688 5516 13694 5568
rect 13740 5556 13768 5587
rect 13814 5584 13820 5636
rect 13872 5624 13878 5636
rect 13909 5627 13967 5633
rect 13909 5624 13921 5627
rect 13872 5596 13921 5624
rect 13872 5584 13878 5596
rect 13909 5593 13921 5596
rect 13955 5593 13967 5627
rect 14384 5624 14412 5655
rect 14642 5652 14648 5664
rect 14700 5692 14706 5704
rect 15120 5701 15148 5732
rect 15856 5704 15884 5732
rect 14921 5695 14979 5701
rect 14921 5692 14933 5695
rect 14700 5664 14933 5692
rect 14700 5652 14706 5664
rect 14921 5661 14933 5664
rect 14967 5661 14979 5695
rect 14921 5655 14979 5661
rect 15105 5695 15163 5701
rect 15105 5661 15117 5695
rect 15151 5661 15163 5695
rect 15105 5655 15163 5661
rect 15289 5695 15347 5701
rect 15289 5661 15301 5695
rect 15335 5661 15347 5695
rect 15289 5655 15347 5661
rect 14550 5624 14556 5636
rect 14384 5596 14556 5624
rect 13909 5587 13967 5593
rect 14182 5556 14188 5568
rect 13740 5528 14188 5556
rect 14182 5516 14188 5528
rect 14240 5516 14246 5568
rect 14366 5516 14372 5568
rect 14424 5556 14430 5568
rect 14476 5556 14504 5596
rect 14550 5584 14556 5596
rect 14608 5584 14614 5636
rect 14734 5624 14740 5636
rect 14660 5596 14740 5624
rect 14660 5565 14688 5596
rect 14734 5584 14740 5596
rect 14792 5584 14798 5636
rect 15010 5584 15016 5636
rect 15068 5584 15074 5636
rect 15304 5624 15332 5655
rect 15654 5652 15660 5704
rect 15712 5692 15718 5704
rect 15749 5695 15807 5701
rect 15749 5692 15761 5695
rect 15712 5664 15761 5692
rect 15712 5652 15718 5664
rect 15749 5661 15761 5664
rect 15795 5661 15807 5695
rect 15749 5655 15807 5661
rect 15838 5652 15844 5704
rect 15896 5652 15902 5704
rect 15930 5652 15936 5704
rect 15988 5652 15994 5704
rect 16114 5652 16120 5704
rect 16172 5652 16178 5704
rect 15120 5596 15332 5624
rect 14424 5528 14504 5556
rect 14645 5559 14703 5565
rect 14424 5516 14430 5528
rect 14645 5525 14657 5559
rect 14691 5525 14703 5559
rect 14645 5519 14703 5525
rect 14826 5516 14832 5568
rect 14884 5556 14890 5568
rect 15120 5556 15148 5596
rect 14884 5528 15148 5556
rect 14884 5516 14890 5528
rect 15286 5516 15292 5568
rect 15344 5556 15350 5568
rect 15473 5559 15531 5565
rect 15473 5556 15485 5559
rect 15344 5528 15485 5556
rect 15344 5516 15350 5528
rect 15473 5525 15485 5528
rect 15519 5525 15531 5559
rect 15473 5519 15531 5525
rect 1104 5466 16652 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 16652 5466
rect 1104 5392 16652 5414
rect 9398 5312 9404 5364
rect 9456 5352 9462 5364
rect 10045 5355 10103 5361
rect 10045 5352 10057 5355
rect 9456 5324 10057 5352
rect 9456 5312 9462 5324
rect 10045 5321 10057 5324
rect 10091 5352 10103 5355
rect 10778 5352 10784 5364
rect 10091 5324 10784 5352
rect 10091 5321 10103 5324
rect 10045 5315 10103 5321
rect 10778 5312 10784 5324
rect 10836 5312 10842 5364
rect 11974 5312 11980 5364
rect 12032 5352 12038 5364
rect 12710 5352 12716 5364
rect 12032 5324 12716 5352
rect 12032 5312 12038 5324
rect 12710 5312 12716 5324
rect 12768 5312 12774 5364
rect 12805 5355 12863 5361
rect 12805 5321 12817 5355
rect 12851 5352 12863 5355
rect 14001 5355 14059 5361
rect 14001 5352 14013 5355
rect 12851 5324 14013 5352
rect 12851 5321 12863 5324
rect 12805 5315 12863 5321
rect 14001 5321 14013 5324
rect 14047 5321 14059 5355
rect 14001 5315 14059 5321
rect 15378 5312 15384 5364
rect 15436 5352 15442 5364
rect 15436 5324 16068 5352
rect 15436 5312 15442 5324
rect 9214 5244 9220 5296
rect 9272 5284 9278 5296
rect 9490 5284 9496 5296
rect 9272 5256 9496 5284
rect 9272 5244 9278 5256
rect 9490 5244 9496 5256
rect 9548 5244 9554 5296
rect 10597 5287 10655 5293
rect 10597 5284 10609 5287
rect 10152 5256 10609 5284
rect 10152 5225 10180 5256
rect 10597 5253 10609 5256
rect 10643 5284 10655 5287
rect 11054 5284 11060 5296
rect 10643 5256 11060 5284
rect 10643 5253 10655 5256
rect 10597 5247 10655 5253
rect 11054 5244 11060 5256
rect 11112 5244 11118 5296
rect 12728 5284 12756 5312
rect 12728 5256 13124 5284
rect 9953 5219 10011 5225
rect 9953 5185 9965 5219
rect 9999 5185 10011 5219
rect 9953 5179 10011 5185
rect 10137 5219 10195 5225
rect 10137 5185 10149 5219
rect 10183 5185 10195 5219
rect 10137 5179 10195 5185
rect 10413 5219 10471 5225
rect 10413 5185 10425 5219
rect 10459 5185 10471 5219
rect 10413 5179 10471 5185
rect 10781 5219 10839 5225
rect 10781 5185 10793 5219
rect 10827 5216 10839 5219
rect 10870 5216 10876 5228
rect 10827 5188 10876 5216
rect 10827 5185 10839 5188
rect 10781 5179 10839 5185
rect 9968 5148 9996 5179
rect 10428 5148 10456 5179
rect 10870 5176 10876 5188
rect 10928 5176 10934 5228
rect 11149 5219 11207 5225
rect 11149 5185 11161 5219
rect 11195 5216 11207 5219
rect 11698 5216 11704 5228
rect 11195 5188 11704 5216
rect 11195 5185 11207 5188
rect 11149 5179 11207 5185
rect 11698 5176 11704 5188
rect 11756 5176 11762 5228
rect 12894 5176 12900 5228
rect 12952 5176 12958 5228
rect 13096 5216 13124 5256
rect 13354 5244 13360 5296
rect 13412 5284 13418 5296
rect 13412 5256 13676 5284
rect 13412 5244 13418 5256
rect 13648 5225 13676 5256
rect 13814 5244 13820 5296
rect 13872 5284 13878 5296
rect 13872 5256 15976 5284
rect 13872 5244 13878 5256
rect 13541 5219 13599 5225
rect 13541 5216 13553 5219
rect 13096 5188 13553 5216
rect 13541 5185 13553 5188
rect 13587 5185 13599 5219
rect 13541 5179 13599 5185
rect 13633 5219 13691 5225
rect 13633 5185 13645 5219
rect 13679 5185 13691 5219
rect 13633 5179 13691 5185
rect 13725 5219 13783 5225
rect 13725 5185 13737 5219
rect 13771 5216 13783 5219
rect 13771 5188 13860 5216
rect 13771 5185 13783 5188
rect 13725 5179 13783 5185
rect 9968 5120 11192 5148
rect 9490 5040 9496 5092
rect 9548 5080 9554 5092
rect 10229 5083 10287 5089
rect 10229 5080 10241 5083
rect 9548 5052 10241 5080
rect 9548 5040 9554 5052
rect 10229 5049 10241 5052
rect 10275 5049 10287 5083
rect 10229 5043 10287 5049
rect 11164 5024 11192 5120
rect 12066 5108 12072 5160
rect 12124 5108 12130 5160
rect 12158 5108 12164 5160
rect 12216 5108 12222 5160
rect 12986 5108 12992 5160
rect 13044 5108 13050 5160
rect 11333 5083 11391 5089
rect 11333 5049 11345 5083
rect 11379 5080 11391 5083
rect 12894 5080 12900 5092
rect 11379 5052 12900 5080
rect 11379 5049 11391 5052
rect 11333 5043 11391 5049
rect 12894 5040 12900 5052
rect 12952 5040 12958 5092
rect 11146 4972 11152 5024
rect 11204 4972 11210 5024
rect 11609 5015 11667 5021
rect 11609 4981 11621 5015
rect 11655 5012 11667 5015
rect 11698 5012 11704 5024
rect 11655 4984 11704 5012
rect 11655 4981 11667 4984
rect 11609 4975 11667 4981
rect 11698 4972 11704 4984
rect 11756 4972 11762 5024
rect 12434 4972 12440 5024
rect 12492 4972 12498 5024
rect 13265 5015 13323 5021
rect 13265 4981 13277 5015
rect 13311 5012 13323 5015
rect 13354 5012 13360 5024
rect 13311 4984 13360 5012
rect 13311 4981 13323 4984
rect 13265 4975 13323 4981
rect 13354 4972 13360 4984
rect 13412 4972 13418 5024
rect 13556 5012 13584 5179
rect 13630 5040 13636 5092
rect 13688 5080 13694 5092
rect 13832 5080 13860 5188
rect 13906 5176 13912 5228
rect 13964 5176 13970 5228
rect 14366 5176 14372 5228
rect 14424 5216 14430 5228
rect 15013 5219 15071 5225
rect 15013 5216 15025 5219
rect 14424 5188 15025 5216
rect 14424 5176 14430 5188
rect 15013 5185 15025 5188
rect 15059 5185 15071 5219
rect 15013 5179 15071 5185
rect 15102 5176 15108 5228
rect 15160 5176 15166 5228
rect 15194 5176 15200 5228
rect 15252 5176 15258 5228
rect 15378 5176 15384 5228
rect 15436 5176 15442 5228
rect 15948 5225 15976 5256
rect 15749 5219 15807 5225
rect 15749 5185 15761 5219
rect 15795 5185 15807 5219
rect 15749 5179 15807 5185
rect 15841 5219 15899 5225
rect 15841 5185 15853 5219
rect 15887 5185 15899 5219
rect 15841 5179 15899 5185
rect 15933 5219 15991 5225
rect 15933 5185 15945 5219
rect 15979 5185 15991 5219
rect 16040 5216 16068 5324
rect 16114 5216 16120 5228
rect 16040 5188 16120 5216
rect 15933 5179 15991 5185
rect 14182 5108 14188 5160
rect 14240 5148 14246 5160
rect 14553 5151 14611 5157
rect 14553 5148 14565 5151
rect 14240 5120 14565 5148
rect 14240 5108 14246 5120
rect 14553 5117 14565 5120
rect 14599 5117 14611 5151
rect 14553 5111 14611 5117
rect 14642 5108 14648 5160
rect 14700 5148 14706 5160
rect 15764 5148 15792 5179
rect 14700 5120 15792 5148
rect 14700 5108 14706 5120
rect 13688 5052 13860 5080
rect 13688 5040 13694 5052
rect 13906 5040 13912 5092
rect 13964 5080 13970 5092
rect 13964 5052 15056 5080
rect 13964 5040 13970 5052
rect 14366 5012 14372 5024
rect 13556 4984 14372 5012
rect 14366 4972 14372 4984
rect 14424 4972 14430 5024
rect 14734 4972 14740 5024
rect 14792 4972 14798 5024
rect 15028 5012 15056 5052
rect 15102 5040 15108 5092
rect 15160 5080 15166 5092
rect 15856 5080 15884 5179
rect 16114 5176 16120 5188
rect 16172 5176 16178 5228
rect 15160 5052 15884 5080
rect 15160 5040 15166 5052
rect 15378 5012 15384 5024
rect 15028 4984 15384 5012
rect 15378 4972 15384 4984
rect 15436 4972 15442 5024
rect 15470 4972 15476 5024
rect 15528 4972 15534 5024
rect 1104 4922 16652 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 16652 4922
rect 1104 4848 16652 4870
rect 8938 4768 8944 4820
rect 8996 4808 9002 4820
rect 9033 4811 9091 4817
rect 9033 4808 9045 4811
rect 8996 4780 9045 4808
rect 8996 4768 9002 4780
rect 9033 4777 9045 4780
rect 9079 4777 9091 4811
rect 9033 4771 9091 4777
rect 11146 4768 11152 4820
rect 11204 4768 11210 4820
rect 12710 4768 12716 4820
rect 12768 4808 12774 4820
rect 12805 4811 12863 4817
rect 12805 4808 12817 4811
rect 12768 4780 12817 4808
rect 12768 4768 12774 4780
rect 12805 4777 12817 4780
rect 12851 4777 12863 4811
rect 12805 4771 12863 4777
rect 14093 4811 14151 4817
rect 14093 4777 14105 4811
rect 14139 4808 14151 4811
rect 14274 4808 14280 4820
rect 14139 4780 14280 4808
rect 14139 4777 14151 4780
rect 14093 4771 14151 4777
rect 14274 4768 14280 4780
rect 14332 4768 14338 4820
rect 15838 4700 15844 4752
rect 15896 4700 15902 4752
rect 9122 4632 9128 4684
rect 9180 4672 9186 4684
rect 9217 4675 9275 4681
rect 9217 4672 9229 4675
rect 9180 4644 9229 4672
rect 9180 4632 9186 4644
rect 9217 4641 9229 4644
rect 9263 4641 9275 4675
rect 9217 4635 9275 4641
rect 12894 4632 12900 4684
rect 12952 4672 12958 4684
rect 13541 4675 13599 4681
rect 13541 4672 13553 4675
rect 12952 4644 13553 4672
rect 12952 4632 12958 4644
rect 13541 4641 13553 4644
rect 13587 4641 13599 4675
rect 15856 4672 15884 4700
rect 15856 4644 15976 4672
rect 13541 4635 13599 4641
rect 8846 4564 8852 4616
rect 8904 4604 8910 4616
rect 8941 4607 8999 4613
rect 8941 4604 8953 4607
rect 8904 4576 8953 4604
rect 8904 4564 8910 4576
rect 8941 4573 8953 4576
rect 8987 4604 8999 4607
rect 9306 4604 9312 4616
rect 8987 4576 9312 4604
rect 8987 4573 8999 4576
rect 8941 4567 8999 4573
rect 9306 4564 9312 4576
rect 9364 4564 9370 4616
rect 9398 4564 9404 4616
rect 9456 4564 9462 4616
rect 9490 4564 9496 4616
rect 9548 4564 9554 4616
rect 9769 4607 9827 4613
rect 9769 4573 9781 4607
rect 9815 4604 9827 4607
rect 9858 4604 9864 4616
rect 9815 4576 9864 4604
rect 9815 4573 9827 4576
rect 9769 4567 9827 4573
rect 9858 4564 9864 4576
rect 9916 4564 9922 4616
rect 11422 4564 11428 4616
rect 11480 4564 11486 4616
rect 11698 4613 11704 4616
rect 11692 4604 11704 4613
rect 11659 4576 11704 4604
rect 11692 4567 11704 4576
rect 11698 4564 11704 4567
rect 11756 4564 11762 4616
rect 13449 4607 13507 4613
rect 13449 4604 13461 4607
rect 11808 4576 13461 4604
rect 9677 4539 9735 4545
rect 9677 4505 9689 4539
rect 9723 4536 9735 4539
rect 10014 4539 10072 4545
rect 10014 4536 10026 4539
rect 9723 4508 10026 4536
rect 9723 4505 9735 4508
rect 9677 4499 9735 4505
rect 10014 4505 10026 4508
rect 10060 4505 10072 4539
rect 10014 4499 10072 4505
rect 11606 4496 11612 4548
rect 11664 4536 11670 4548
rect 11808 4536 11836 4576
rect 13449 4573 13461 4576
rect 13495 4604 13507 4607
rect 14366 4604 14372 4616
rect 13495 4576 14372 4604
rect 13495 4573 13507 4576
rect 13449 4567 13507 4573
rect 14366 4564 14372 4576
rect 14424 4604 14430 4616
rect 14642 4604 14648 4616
rect 14424 4576 14648 4604
rect 14424 4564 14430 4576
rect 14642 4564 14648 4576
rect 14700 4564 14706 4616
rect 14918 4564 14924 4616
rect 14976 4604 14982 4616
rect 15948 4613 15976 4644
rect 15473 4607 15531 4613
rect 15473 4604 15485 4607
rect 14976 4576 15485 4604
rect 14976 4564 14982 4576
rect 15473 4573 15485 4576
rect 15519 4573 15531 4607
rect 15473 4567 15531 4573
rect 15841 4607 15899 4613
rect 15841 4573 15853 4607
rect 15887 4573 15899 4607
rect 15841 4567 15899 4573
rect 15933 4607 15991 4613
rect 15933 4573 15945 4607
rect 15979 4573 15991 4607
rect 15933 4567 15991 4573
rect 13357 4539 13415 4545
rect 13357 4536 13369 4539
rect 11664 4508 11836 4536
rect 12406 4508 13369 4536
rect 11664 4496 11670 4508
rect 9217 4471 9275 4477
rect 9217 4437 9229 4471
rect 9263 4468 9275 4471
rect 9582 4468 9588 4480
rect 9263 4440 9588 4468
rect 9263 4437 9275 4440
rect 9217 4431 9275 4437
rect 9582 4428 9588 4440
rect 9640 4428 9646 4480
rect 10778 4428 10784 4480
rect 10836 4468 10842 4480
rect 12066 4468 12072 4480
rect 10836 4440 12072 4468
rect 10836 4428 10842 4440
rect 12066 4428 12072 4440
rect 12124 4468 12130 4480
rect 12406 4468 12434 4508
rect 13357 4505 13369 4508
rect 13403 4505 13415 4539
rect 13357 4499 13415 4505
rect 14734 4496 14740 4548
rect 14792 4536 14798 4548
rect 15206 4539 15264 4545
rect 15206 4536 15218 4539
rect 14792 4508 15218 4536
rect 14792 4496 14798 4508
rect 15206 4505 15218 4508
rect 15252 4505 15264 4539
rect 15856 4536 15884 4567
rect 16022 4564 16028 4616
rect 16080 4564 16086 4616
rect 16114 4564 16120 4616
rect 16172 4604 16178 4616
rect 16209 4607 16267 4613
rect 16209 4604 16221 4607
rect 16172 4576 16221 4604
rect 16172 4564 16178 4576
rect 16209 4573 16221 4576
rect 16255 4573 16267 4607
rect 16209 4567 16267 4573
rect 16298 4536 16304 4548
rect 15856 4508 16304 4536
rect 15206 4499 15264 4505
rect 16298 4496 16304 4508
rect 16356 4496 16362 4548
rect 12124 4440 12434 4468
rect 12124 4428 12130 4440
rect 12894 4428 12900 4480
rect 12952 4468 12958 4480
rect 12989 4471 13047 4477
rect 12989 4468 13001 4471
rect 12952 4440 13001 4468
rect 12952 4428 12958 4440
rect 12989 4437 13001 4440
rect 13035 4437 13047 4471
rect 12989 4431 13047 4437
rect 15562 4428 15568 4480
rect 15620 4428 15626 4480
rect 1104 4378 16652 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 16652 4378
rect 1104 4304 16652 4326
rect 10962 4264 10968 4276
rect 8220 4236 10968 4264
rect 8220 4205 8248 4236
rect 10962 4224 10968 4236
rect 11020 4224 11026 4276
rect 11606 4224 11612 4276
rect 11664 4224 11670 4276
rect 8205 4199 8263 4205
rect 8205 4165 8217 4199
rect 8251 4165 8263 4199
rect 8205 4159 8263 4165
rect 8846 4156 8852 4208
rect 8904 4196 8910 4208
rect 9217 4199 9275 4205
rect 9217 4196 9229 4199
rect 8904 4168 9229 4196
rect 8904 4156 8910 4168
rect 9217 4165 9229 4168
rect 9263 4165 9275 4199
rect 9217 4159 9275 4165
rect 9306 4156 9312 4208
rect 9364 4156 9370 4208
rect 9447 4199 9505 4205
rect 9447 4165 9459 4199
rect 9493 4196 9505 4199
rect 9766 4196 9772 4208
rect 9493 4168 9772 4196
rect 9493 4165 9505 4168
rect 9447 4159 9505 4165
rect 9766 4156 9772 4168
rect 9824 4156 9830 4208
rect 12744 4199 12802 4205
rect 12744 4165 12756 4199
rect 12790 4196 12802 4199
rect 12894 4196 12900 4208
rect 12790 4168 12900 4196
rect 12790 4165 12802 4168
rect 12744 4159 12802 4165
rect 12894 4156 12900 4168
rect 12952 4156 12958 4208
rect 13814 4196 13820 4208
rect 13280 4168 13820 4196
rect 8389 4131 8447 4137
rect 8389 4097 8401 4131
rect 8435 4128 8447 4131
rect 8481 4131 8539 4137
rect 8481 4128 8493 4131
rect 8435 4100 8493 4128
rect 8435 4097 8447 4100
rect 8389 4091 8447 4097
rect 8481 4097 8493 4100
rect 8527 4097 8539 4131
rect 8481 4091 8539 4097
rect 8665 4131 8723 4137
rect 8665 4097 8677 4131
rect 8711 4128 8723 4131
rect 8711 4100 9076 4128
rect 8711 4097 8723 4100
rect 8665 4091 8723 4097
rect 8849 4063 8907 4069
rect 8849 4029 8861 4063
rect 8895 4029 8907 4063
rect 9048 4060 9076 4100
rect 9122 4088 9128 4140
rect 9180 4088 9186 4140
rect 9582 4088 9588 4140
rect 9640 4088 9646 4140
rect 10128 4131 10186 4137
rect 10128 4097 10140 4131
rect 10174 4128 10186 4131
rect 10410 4128 10416 4140
rect 10174 4100 10416 4128
rect 10174 4097 10186 4100
rect 10128 4091 10186 4097
rect 10410 4088 10416 4100
rect 10468 4088 10474 4140
rect 12989 4131 13047 4137
rect 12989 4097 13001 4131
rect 13035 4128 13047 4131
rect 13081 4131 13139 4137
rect 13081 4128 13093 4131
rect 13035 4100 13093 4128
rect 13035 4097 13047 4100
rect 12989 4091 13047 4097
rect 13081 4097 13093 4100
rect 13127 4128 13139 4131
rect 13280 4128 13308 4168
rect 13814 4156 13820 4168
rect 13872 4196 13878 4208
rect 14918 4196 14924 4208
rect 13872 4168 14924 4196
rect 13872 4156 13878 4168
rect 14918 4156 14924 4168
rect 14976 4196 14982 4208
rect 14976 4168 16068 4196
rect 14976 4156 14982 4168
rect 13354 4137 13360 4140
rect 13127 4100 13308 4128
rect 13127 4097 13139 4100
rect 13081 4091 13139 4097
rect 13348 4091 13360 4137
rect 13412 4128 13418 4140
rect 13412 4100 13448 4128
rect 13354 4088 13360 4091
rect 13412 4088 13418 4100
rect 15470 4088 15476 4140
rect 15528 4128 15534 4140
rect 16040 4137 16068 4168
rect 15758 4131 15816 4137
rect 15758 4128 15770 4131
rect 15528 4100 15770 4128
rect 15528 4088 15534 4100
rect 15758 4097 15770 4100
rect 15804 4097 15816 4131
rect 15758 4091 15816 4097
rect 16025 4131 16083 4137
rect 16025 4097 16037 4131
rect 16071 4097 16083 4131
rect 16025 4091 16083 4097
rect 9398 4060 9404 4072
rect 9048 4032 9404 4060
rect 8849 4023 8907 4029
rect 8864 3992 8892 4023
rect 9398 4020 9404 4032
rect 9456 4020 9462 4072
rect 9858 4020 9864 4072
rect 9916 4020 9922 4072
rect 8864 3964 9904 3992
rect 8018 3884 8024 3936
rect 8076 3884 8082 3936
rect 8938 3884 8944 3936
rect 8996 3884 9002 3936
rect 9876 3924 9904 3964
rect 11238 3952 11244 4004
rect 11296 3952 11302 4004
rect 14645 3995 14703 4001
rect 14645 3961 14657 3995
rect 14691 3992 14703 3995
rect 15010 3992 15016 4004
rect 14691 3964 15016 3992
rect 14691 3961 14703 3964
rect 14645 3955 14703 3961
rect 15010 3952 15016 3964
rect 15068 3952 15074 4004
rect 10870 3924 10876 3936
rect 9876 3896 10876 3924
rect 10870 3884 10876 3896
rect 10928 3884 10934 3936
rect 14458 3884 14464 3936
rect 14516 3884 14522 3936
rect 1104 3834 16652 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 16652 3834
rect 1104 3760 16652 3782
rect 9766 3680 9772 3732
rect 9824 3680 9830 3732
rect 10870 3680 10876 3732
rect 10928 3720 10934 3732
rect 11241 3723 11299 3729
rect 11241 3720 11253 3723
rect 10928 3692 11253 3720
rect 10928 3680 10934 3692
rect 11241 3689 11253 3692
rect 11287 3720 11299 3723
rect 11517 3723 11575 3729
rect 11517 3720 11529 3723
rect 11287 3692 11529 3720
rect 11287 3689 11299 3692
rect 11241 3683 11299 3689
rect 11517 3689 11529 3692
rect 11563 3689 11575 3723
rect 11517 3683 11575 3689
rect 11701 3723 11759 3729
rect 11701 3689 11713 3723
rect 11747 3720 11759 3723
rect 12158 3720 12164 3732
rect 11747 3692 12164 3720
rect 11747 3689 11759 3692
rect 11701 3683 11759 3689
rect 12158 3680 12164 3692
rect 12216 3680 12222 3732
rect 13357 3723 13415 3729
rect 13357 3689 13369 3723
rect 13403 3720 13415 3723
rect 14182 3720 14188 3732
rect 13403 3692 14188 3720
rect 13403 3689 13415 3692
rect 13357 3683 13415 3689
rect 14182 3680 14188 3692
rect 14240 3680 14246 3732
rect 14292 3692 14688 3720
rect 13906 3652 13912 3664
rect 13004 3624 13912 3652
rect 8018 3544 8024 3596
rect 8076 3584 8082 3596
rect 8076 3556 9352 3584
rect 8076 3544 8082 3556
rect 8754 3476 8760 3528
rect 8812 3476 8818 3528
rect 9214 3476 9220 3528
rect 9272 3476 9278 3528
rect 9324 3516 9352 3556
rect 9858 3544 9864 3596
rect 9916 3544 9922 3596
rect 11422 3544 11428 3596
rect 11480 3584 11486 3596
rect 11974 3584 11980 3596
rect 11480 3556 11980 3584
rect 11480 3544 11486 3556
rect 11974 3544 11980 3556
rect 12032 3544 12038 3596
rect 10117 3519 10175 3525
rect 10117 3516 10129 3519
rect 9324 3488 10129 3516
rect 10117 3485 10129 3488
rect 10163 3485 10175 3519
rect 13004 3516 13032 3624
rect 13906 3612 13912 3624
rect 13964 3652 13970 3664
rect 14292 3652 14320 3692
rect 13964 3624 14320 3652
rect 14384 3624 14596 3652
rect 13964 3612 13970 3624
rect 13817 3587 13875 3593
rect 13817 3553 13829 3587
rect 13863 3584 13875 3587
rect 14384 3584 14412 3624
rect 13863 3556 14412 3584
rect 13863 3553 13875 3556
rect 13817 3547 13875 3553
rect 10117 3479 10175 3485
rect 11072 3488 13032 3516
rect 9122 3408 9128 3460
rect 9180 3448 9186 3460
rect 11072 3448 11100 3488
rect 13078 3476 13084 3528
rect 13136 3516 13142 3528
rect 13449 3519 13507 3525
rect 13449 3516 13461 3519
rect 13136 3488 13461 3516
rect 13136 3476 13142 3488
rect 13449 3485 13461 3488
rect 13495 3516 13507 3519
rect 14274 3516 14280 3528
rect 13495 3488 14280 3516
rect 13495 3485 13507 3488
rect 13449 3479 13507 3485
rect 14274 3476 14280 3488
rect 14332 3476 14338 3528
rect 14366 3476 14372 3528
rect 14424 3476 14430 3528
rect 14568 3525 14596 3624
rect 14461 3519 14519 3525
rect 14461 3485 14473 3519
rect 14507 3485 14519 3519
rect 14461 3479 14519 3485
rect 14553 3519 14611 3525
rect 14553 3485 14565 3519
rect 14599 3485 14611 3519
rect 14660 3516 14688 3692
rect 15654 3680 15660 3732
rect 15712 3720 15718 3732
rect 16301 3723 16359 3729
rect 16301 3720 16313 3723
rect 15712 3692 16313 3720
rect 15712 3680 15718 3692
rect 16301 3689 16313 3692
rect 16347 3689 16359 3723
rect 16301 3683 16359 3689
rect 14918 3544 14924 3596
rect 14976 3544 14982 3596
rect 14737 3519 14795 3525
rect 14737 3516 14749 3519
rect 14660 3488 14749 3516
rect 14553 3479 14611 3485
rect 14737 3485 14749 3488
rect 14783 3485 14795 3519
rect 14737 3479 14795 3485
rect 15188 3519 15246 3525
rect 15188 3485 15200 3519
rect 15234 3516 15246 3519
rect 15562 3516 15568 3528
rect 15234 3488 15568 3516
rect 15234 3485 15246 3488
rect 15188 3479 15246 3485
rect 9180 3420 11100 3448
rect 9180 3408 9186 3420
rect 11146 3408 11152 3460
rect 11204 3448 11210 3460
rect 11333 3451 11391 3457
rect 11333 3448 11345 3451
rect 11204 3420 11345 3448
rect 11204 3408 11210 3420
rect 11333 3417 11345 3420
rect 11379 3417 11391 3451
rect 11333 3411 11391 3417
rect 11514 3408 11520 3460
rect 11572 3457 11578 3460
rect 11572 3451 11591 3457
rect 11579 3417 11591 3451
rect 11572 3411 11591 3417
rect 12244 3451 12302 3457
rect 12244 3417 12256 3451
rect 12290 3448 12302 3451
rect 12434 3448 12440 3460
rect 12290 3420 12440 3448
rect 12290 3417 12302 3420
rect 12244 3411 12302 3417
rect 11572 3408 11578 3411
rect 12434 3408 12440 3420
rect 12492 3408 12498 3460
rect 13633 3451 13691 3457
rect 13633 3417 13645 3451
rect 13679 3448 13691 3451
rect 13906 3448 13912 3460
rect 13679 3420 13912 3448
rect 13679 3417 13691 3420
rect 13633 3411 13691 3417
rect 13906 3408 13912 3420
rect 13964 3408 13970 3460
rect 14476 3448 14504 3479
rect 15562 3476 15568 3488
rect 15620 3476 15626 3528
rect 15838 3448 15844 3460
rect 14476 3420 15844 3448
rect 15838 3408 15844 3420
rect 15896 3408 15902 3460
rect 8573 3383 8631 3389
rect 8573 3349 8585 3383
rect 8619 3380 8631 3383
rect 8754 3380 8760 3392
rect 8619 3352 8760 3380
rect 8619 3349 8631 3352
rect 8573 3343 8631 3349
rect 8754 3340 8760 3352
rect 8812 3340 8818 3392
rect 14090 3340 14096 3392
rect 14148 3340 14154 3392
rect 1104 3290 16652 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 16652 3290
rect 1104 3216 16652 3238
rect 9214 3136 9220 3188
rect 9272 3176 9278 3188
rect 9401 3179 9459 3185
rect 9401 3176 9413 3179
rect 9272 3148 9413 3176
rect 9272 3136 9278 3148
rect 9401 3145 9413 3148
rect 9447 3145 9459 3179
rect 9401 3139 9459 3145
rect 10410 3136 10416 3188
rect 10468 3136 10474 3188
rect 10781 3179 10839 3185
rect 10781 3145 10793 3179
rect 10827 3176 10839 3179
rect 11238 3176 11244 3188
rect 10827 3148 11244 3176
rect 10827 3145 10839 3148
rect 10781 3139 10839 3145
rect 11238 3136 11244 3148
rect 11296 3136 11302 3188
rect 13906 3136 13912 3188
rect 13964 3176 13970 3188
rect 14093 3179 14151 3185
rect 14093 3176 14105 3179
rect 13964 3148 14105 3176
rect 13964 3136 13970 3148
rect 14093 3145 14105 3148
rect 14139 3176 14151 3179
rect 14550 3176 14556 3188
rect 14139 3148 14556 3176
rect 14139 3145 14151 3148
rect 14093 3139 14151 3145
rect 14550 3136 14556 3148
rect 14608 3136 14614 3188
rect 14829 3179 14887 3185
rect 14829 3145 14841 3179
rect 14875 3176 14887 3179
rect 15930 3176 15936 3188
rect 14875 3148 15936 3176
rect 14875 3145 14887 3148
rect 14829 3139 14887 3145
rect 15930 3136 15936 3148
rect 15988 3136 15994 3188
rect 8288 3111 8346 3117
rect 8288 3077 8300 3111
rect 8334 3108 8346 3111
rect 8938 3108 8944 3120
rect 8334 3080 8944 3108
rect 8334 3077 8346 3080
rect 8288 3071 8346 3077
rect 8938 3068 8944 3080
rect 8996 3068 9002 3120
rect 11974 3068 11980 3120
rect 12032 3108 12038 3120
rect 13814 3108 13820 3120
rect 12032 3080 13820 3108
rect 12032 3068 12038 3080
rect 5534 3000 5540 3052
rect 5592 3040 5598 3052
rect 12728 3049 12756 3080
rect 13814 3068 13820 3080
rect 13872 3068 13878 3120
rect 14645 3111 14703 3117
rect 14645 3077 14657 3111
rect 14691 3108 14703 3111
rect 14734 3108 14740 3120
rect 14691 3080 14740 3108
rect 14691 3077 14703 3080
rect 14645 3071 14703 3077
rect 14734 3068 14740 3080
rect 14792 3068 14798 3120
rect 15188 3111 15246 3117
rect 15188 3077 15200 3111
rect 15234 3108 15246 3111
rect 15286 3108 15292 3120
rect 15234 3080 15292 3108
rect 15234 3077 15246 3080
rect 15188 3071 15246 3077
rect 15286 3068 15292 3080
rect 15344 3068 15350 3120
rect 8021 3043 8079 3049
rect 8021 3040 8033 3043
rect 5592 3012 8033 3040
rect 5592 3000 5598 3012
rect 8021 3009 8033 3012
rect 8067 3009 8079 3043
rect 8021 3003 8079 3009
rect 12713 3043 12771 3049
rect 12713 3009 12725 3043
rect 12759 3040 12771 3043
rect 12980 3043 13038 3049
rect 12759 3012 12793 3040
rect 12759 3009 12771 3012
rect 12713 3003 12771 3009
rect 12980 3009 12992 3043
rect 13026 3040 13038 3043
rect 14090 3040 14096 3052
rect 13026 3012 14096 3040
rect 13026 3009 13038 3012
rect 12980 3003 13038 3009
rect 14090 3000 14096 3012
rect 14148 3000 14154 3052
rect 14182 3000 14188 3052
rect 14240 3000 14246 3052
rect 14274 3000 14280 3052
rect 14332 3040 14338 3052
rect 14461 3043 14519 3049
rect 14461 3040 14473 3043
rect 14332 3012 14473 3040
rect 14332 3000 14338 3012
rect 14461 3009 14473 3012
rect 14507 3040 14519 3043
rect 14550 3040 14556 3052
rect 14507 3012 14556 3040
rect 14507 3009 14519 3012
rect 14461 3003 14519 3009
rect 14550 3000 14556 3012
rect 14608 3000 14614 3052
rect 14918 3000 14924 3052
rect 14976 3000 14982 3052
rect 10870 2932 10876 2984
rect 10928 2932 10934 2984
rect 10962 2932 10968 2984
rect 11020 2932 11026 2984
rect 13814 2864 13820 2916
rect 13872 2904 13878 2916
rect 14458 2904 14464 2916
rect 13872 2876 14464 2904
rect 13872 2864 13878 2876
rect 14458 2864 14464 2876
rect 14516 2864 14522 2916
rect 14369 2839 14427 2845
rect 14369 2805 14381 2839
rect 14415 2836 14427 2839
rect 14642 2836 14648 2848
rect 14415 2808 14648 2836
rect 14415 2805 14427 2808
rect 14369 2799 14427 2805
rect 14642 2796 14648 2808
rect 14700 2796 14706 2848
rect 14734 2796 14740 2848
rect 14792 2836 14798 2848
rect 16301 2839 16359 2845
rect 16301 2836 16313 2839
rect 14792 2808 16313 2836
rect 14792 2796 14798 2808
rect 16301 2805 16313 2808
rect 16347 2805 16359 2839
rect 16301 2799 16359 2805
rect 1104 2746 16652 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 16652 2746
rect 1104 2672 16652 2694
rect 14826 2592 14832 2644
rect 14884 2592 14890 2644
rect 15194 2592 15200 2644
rect 15252 2592 15258 2644
rect 15749 2635 15807 2641
rect 15749 2601 15761 2635
rect 15795 2632 15807 2635
rect 16022 2632 16028 2644
rect 15795 2604 16028 2632
rect 15795 2601 15807 2604
rect 15749 2595 15807 2601
rect 16022 2592 16028 2604
rect 16080 2592 16086 2644
rect 16206 2592 16212 2644
rect 16264 2592 16270 2644
rect 8389 2567 8447 2573
rect 8389 2533 8401 2567
rect 8435 2564 8447 2567
rect 8846 2564 8852 2576
rect 8435 2536 8852 2564
rect 8435 2533 8447 2536
rect 8389 2527 8447 2533
rect 8846 2524 8852 2536
rect 8904 2524 8910 2576
rect 10045 2567 10103 2573
rect 10045 2533 10057 2567
rect 10091 2564 10103 2567
rect 10870 2564 10876 2576
rect 10091 2536 10876 2564
rect 10091 2533 10103 2536
rect 10045 2527 10103 2533
rect 10870 2524 10876 2536
rect 10928 2524 10934 2576
rect 14550 2524 14556 2576
rect 14608 2564 14614 2576
rect 14608 2536 15424 2564
rect 14608 2524 14614 2536
rect 7469 2499 7527 2505
rect 7469 2465 7481 2499
rect 7515 2496 7527 2499
rect 9306 2496 9312 2508
rect 7515 2468 9312 2496
rect 7515 2465 7527 2468
rect 7469 2459 7527 2465
rect 9306 2456 9312 2468
rect 9364 2456 9370 2508
rect 7098 2388 7104 2440
rect 7156 2428 7162 2440
rect 7193 2431 7251 2437
rect 7193 2428 7205 2431
rect 7156 2400 7205 2428
rect 7156 2388 7162 2400
rect 7193 2397 7205 2400
rect 7239 2397 7251 2431
rect 7193 2391 7251 2397
rect 8754 2388 8760 2440
rect 8812 2388 8818 2440
rect 9214 2388 9220 2440
rect 9272 2428 9278 2440
rect 9401 2431 9459 2437
rect 9401 2428 9413 2431
rect 9272 2400 9413 2428
rect 9272 2388 9278 2400
rect 9401 2397 9413 2400
rect 9447 2397 9459 2431
rect 9401 2391 9459 2397
rect 13265 2431 13323 2437
rect 13265 2397 13277 2431
rect 13311 2428 13323 2431
rect 13814 2428 13820 2440
rect 13311 2400 13820 2428
rect 13311 2397 13323 2400
rect 13265 2391 13323 2397
rect 13814 2388 13820 2400
rect 13872 2388 13878 2440
rect 13906 2388 13912 2440
rect 13964 2388 13970 2440
rect 13998 2388 14004 2440
rect 14056 2428 14062 2440
rect 14553 2431 14611 2437
rect 14553 2428 14565 2431
rect 14056 2400 14565 2428
rect 14056 2388 14062 2400
rect 14553 2397 14565 2400
rect 14599 2397 14611 2431
rect 14553 2391 14611 2397
rect 14642 2388 14648 2440
rect 14700 2388 14706 2440
rect 14734 2388 14740 2440
rect 14792 2428 14798 2440
rect 15396 2437 15424 2536
rect 15013 2431 15071 2437
rect 15013 2428 15025 2431
rect 14792 2400 15025 2428
rect 14792 2388 14798 2400
rect 15013 2397 15025 2400
rect 15059 2397 15071 2431
rect 15013 2391 15071 2397
rect 15381 2431 15439 2437
rect 15381 2397 15393 2431
rect 15427 2397 15439 2431
rect 15381 2391 15439 2397
rect 15565 2431 15623 2437
rect 15565 2397 15577 2431
rect 15611 2428 15623 2431
rect 15654 2428 15660 2440
rect 15611 2400 15660 2428
rect 15611 2397 15623 2400
rect 15565 2391 15623 2397
rect 15654 2388 15660 2400
rect 15712 2428 15718 2440
rect 16025 2431 16083 2437
rect 16025 2428 16037 2431
rect 15712 2400 16037 2428
rect 15712 2388 15718 2400
rect 16025 2397 16037 2400
rect 16071 2397 16083 2431
rect 16025 2391 16083 2397
rect 7742 2320 7748 2372
rect 7800 2360 7806 2372
rect 8205 2363 8263 2369
rect 8205 2360 8217 2363
rect 7800 2332 8217 2360
rect 7800 2320 7806 2332
rect 8205 2329 8217 2332
rect 8251 2329 8263 2363
rect 8205 2323 8263 2329
rect 9674 2320 9680 2372
rect 9732 2360 9738 2372
rect 9861 2363 9919 2369
rect 9861 2360 9873 2363
rect 9732 2332 9873 2360
rect 9732 2320 9738 2332
rect 9861 2329 9873 2332
rect 9907 2329 9919 2363
rect 9861 2323 9919 2329
rect 8386 2252 8392 2304
rect 8444 2292 8450 2304
rect 8573 2295 8631 2301
rect 8573 2292 8585 2295
rect 8444 2264 8585 2292
rect 8444 2252 8450 2264
rect 8573 2261 8585 2264
rect 8619 2261 8631 2295
rect 8573 2255 8631 2261
rect 9030 2252 9036 2304
rect 9088 2292 9094 2304
rect 9217 2295 9275 2301
rect 9217 2292 9229 2295
rect 9088 2264 9229 2292
rect 9088 2252 9094 2264
rect 9217 2261 9229 2264
rect 9263 2261 9275 2295
rect 9217 2255 9275 2261
rect 12894 2252 12900 2304
rect 12952 2292 12958 2304
rect 13081 2295 13139 2301
rect 13081 2292 13093 2295
rect 12952 2264 13093 2292
rect 12952 2252 12958 2264
rect 13081 2261 13093 2264
rect 13127 2261 13139 2295
rect 13081 2255 13139 2261
rect 13538 2252 13544 2304
rect 13596 2292 13602 2304
rect 13725 2295 13783 2301
rect 13725 2292 13737 2295
rect 13596 2264 13737 2292
rect 13596 2252 13602 2264
rect 13725 2261 13737 2264
rect 13771 2261 13783 2295
rect 13725 2255 13783 2261
rect 14182 2252 14188 2304
rect 14240 2292 14246 2304
rect 14369 2295 14427 2301
rect 14369 2292 14381 2295
rect 14240 2264 14381 2292
rect 14240 2252 14246 2264
rect 14369 2261 14381 2264
rect 14415 2261 14427 2295
rect 14369 2255 14427 2261
rect 1104 2202 16652 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 16652 2202
rect 1104 2128 16652 2150
<< via1 >>
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 7748 33056 7800 33108
rect 12900 33056 12952 33108
rect 12992 33056 13044 33108
rect 13544 32988 13596 33040
rect 14832 33056 14884 33108
rect 15292 33056 15344 33108
rect 16488 33056 16540 33108
rect 8116 32895 8168 32904
rect 8116 32861 8125 32895
rect 8125 32861 8159 32895
rect 8159 32861 8168 32895
rect 8116 32852 8168 32861
rect 10600 32895 10652 32904
rect 10600 32861 10609 32895
rect 10609 32861 10643 32895
rect 10643 32861 10652 32895
rect 10600 32852 10652 32861
rect 10876 32852 10928 32904
rect 11336 32895 11388 32904
rect 11336 32861 11345 32895
rect 11345 32861 11379 32895
rect 11379 32861 11388 32895
rect 11336 32852 11388 32861
rect 11520 32895 11572 32904
rect 11520 32861 11529 32895
rect 11529 32861 11563 32895
rect 11563 32861 11572 32895
rect 11520 32852 11572 32861
rect 10416 32759 10468 32768
rect 10416 32725 10425 32759
rect 10425 32725 10459 32759
rect 10459 32725 10468 32759
rect 10416 32716 10468 32725
rect 10784 32759 10836 32768
rect 10784 32725 10793 32759
rect 10793 32725 10827 32759
rect 10827 32725 10836 32759
rect 10784 32716 10836 32725
rect 15476 32920 15528 32972
rect 12256 32759 12308 32768
rect 12256 32725 12265 32759
rect 12265 32725 12299 32759
rect 12299 32725 12308 32759
rect 12256 32716 12308 32725
rect 12532 32784 12584 32836
rect 12808 32784 12860 32836
rect 12992 32784 13044 32836
rect 13176 32759 13228 32768
rect 13176 32725 13185 32759
rect 13185 32725 13219 32759
rect 13219 32725 13228 32759
rect 13176 32716 13228 32725
rect 13360 32827 13412 32836
rect 13360 32793 13369 32827
rect 13369 32793 13403 32827
rect 13403 32793 13412 32827
rect 13360 32784 13412 32793
rect 13452 32784 13504 32836
rect 13912 32895 13964 32904
rect 13912 32861 13921 32895
rect 13921 32861 13955 32895
rect 13955 32861 13964 32895
rect 13912 32852 13964 32861
rect 14924 32852 14976 32904
rect 15292 32852 15344 32904
rect 15384 32852 15436 32904
rect 16120 32852 16172 32904
rect 14188 32784 14240 32836
rect 14280 32827 14332 32836
rect 14280 32793 14289 32827
rect 14289 32793 14323 32827
rect 14323 32793 14332 32827
rect 14280 32784 14332 32793
rect 14372 32784 14424 32836
rect 14648 32784 14700 32836
rect 15660 32784 15712 32836
rect 15752 32827 15804 32836
rect 15752 32793 15761 32827
rect 15761 32793 15795 32827
rect 15795 32793 15804 32827
rect 15752 32784 15804 32793
rect 15844 32827 15896 32836
rect 15844 32793 15853 32827
rect 15853 32793 15887 32827
rect 15887 32793 15896 32827
rect 15844 32784 15896 32793
rect 16212 32784 16264 32836
rect 14464 32759 14516 32768
rect 14464 32725 14473 32759
rect 14473 32725 14507 32759
rect 14507 32725 14516 32759
rect 14464 32716 14516 32725
rect 14832 32716 14884 32768
rect 15292 32716 15344 32768
rect 15476 32716 15528 32768
rect 4874 32614 4926 32666
rect 4938 32614 4990 32666
rect 5002 32614 5054 32666
rect 5066 32614 5118 32666
rect 5130 32614 5182 32666
rect 11336 32512 11388 32564
rect 13360 32512 13412 32564
rect 13452 32512 13504 32564
rect 14372 32512 14424 32564
rect 14464 32512 14516 32564
rect 10784 32444 10836 32496
rect 14004 32444 14056 32496
rect 7196 32419 7248 32428
rect 7196 32385 7205 32419
rect 7205 32385 7239 32419
rect 7239 32385 7248 32419
rect 7196 32376 7248 32385
rect 7380 32419 7432 32428
rect 7380 32385 7389 32419
rect 7389 32385 7423 32419
rect 7423 32385 7432 32419
rect 7380 32376 7432 32385
rect 7472 32376 7524 32428
rect 9128 32419 9180 32428
rect 9128 32385 9137 32419
rect 9137 32385 9171 32419
rect 9171 32385 9180 32419
rect 9128 32376 9180 32385
rect 7656 32308 7708 32360
rect 10784 32351 10836 32360
rect 10784 32317 10793 32351
rect 10793 32317 10827 32351
rect 10827 32317 10836 32351
rect 10784 32308 10836 32317
rect 7012 32283 7064 32292
rect 7012 32249 7021 32283
rect 7021 32249 7055 32283
rect 7055 32249 7064 32283
rect 7012 32240 7064 32249
rect 7104 32283 7156 32292
rect 7104 32249 7113 32283
rect 7113 32249 7147 32283
rect 7147 32249 7156 32283
rect 7104 32240 7156 32249
rect 11060 32240 11112 32292
rect 12072 32351 12124 32360
rect 12072 32317 12081 32351
rect 12081 32317 12115 32351
rect 12115 32317 12124 32351
rect 12072 32308 12124 32317
rect 12624 32240 12676 32292
rect 6736 32215 6788 32224
rect 6736 32181 6745 32215
rect 6745 32181 6779 32215
rect 6779 32181 6788 32215
rect 6736 32172 6788 32181
rect 8392 32172 8444 32224
rect 11336 32215 11388 32224
rect 11336 32181 11345 32215
rect 11345 32181 11379 32215
rect 11379 32181 11388 32215
rect 11336 32172 11388 32181
rect 13544 32419 13596 32428
rect 13544 32385 13562 32419
rect 13562 32385 13596 32419
rect 13544 32376 13596 32385
rect 13728 32376 13780 32428
rect 13912 32308 13964 32360
rect 14464 32419 14516 32428
rect 14464 32385 14473 32419
rect 14473 32385 14507 32419
rect 14507 32385 14516 32419
rect 14464 32376 14516 32385
rect 14924 32444 14976 32496
rect 14648 32308 14700 32360
rect 15016 32376 15068 32428
rect 15660 32444 15712 32496
rect 14832 32308 14884 32360
rect 15108 32240 15160 32292
rect 15936 32419 15988 32428
rect 15936 32385 15945 32419
rect 15945 32385 15979 32419
rect 15979 32385 15988 32419
rect 15936 32376 15988 32385
rect 15660 32308 15712 32360
rect 15844 32308 15896 32360
rect 14096 32215 14148 32224
rect 14096 32181 14105 32215
rect 14105 32181 14139 32215
rect 14139 32181 14148 32215
rect 14096 32172 14148 32181
rect 14372 32172 14424 32224
rect 14924 32172 14976 32224
rect 15568 32215 15620 32224
rect 15568 32181 15577 32215
rect 15577 32181 15611 32215
rect 15611 32181 15620 32215
rect 15568 32172 15620 32181
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 8116 31968 8168 32020
rect 8392 31875 8444 31884
rect 8392 31841 8401 31875
rect 8401 31841 8435 31875
rect 8435 31841 8444 31875
rect 8392 31832 8444 31841
rect 8116 31807 8168 31816
rect 8116 31773 8125 31807
rect 8125 31773 8159 31807
rect 8159 31773 8168 31807
rect 8116 31764 8168 31773
rect 8484 31764 8536 31816
rect 9128 31968 9180 32020
rect 11520 31968 11572 32020
rect 13728 31968 13780 32020
rect 13820 32011 13872 32020
rect 13820 31977 13829 32011
rect 13829 31977 13863 32011
rect 13863 31977 13872 32011
rect 13820 31968 13872 31977
rect 15384 31968 15436 32020
rect 10784 31900 10836 31952
rect 10968 31900 11020 31952
rect 9404 31764 9456 31816
rect 9680 31807 9732 31816
rect 9680 31773 9689 31807
rect 9689 31773 9723 31807
rect 9723 31773 9732 31807
rect 9680 31764 9732 31773
rect 16028 31900 16080 31952
rect 11336 31832 11388 31884
rect 6736 31739 6788 31748
rect 6736 31705 6770 31739
rect 6770 31705 6788 31739
rect 6736 31696 6788 31705
rect 6920 31696 6972 31748
rect 8852 31696 8904 31748
rect 10692 31696 10744 31748
rect 13084 31696 13136 31748
rect 13728 31764 13780 31816
rect 13912 31764 13964 31816
rect 14924 31764 14976 31816
rect 14372 31739 14424 31748
rect 14372 31705 14406 31739
rect 14406 31705 14424 31739
rect 14372 31696 14424 31705
rect 14464 31696 14516 31748
rect 15108 31764 15160 31816
rect 15200 31764 15252 31816
rect 15936 31832 15988 31884
rect 16396 31832 16448 31884
rect 16120 31764 16172 31816
rect 7932 31671 7984 31680
rect 7932 31637 7941 31671
rect 7941 31637 7975 31671
rect 7975 31637 7984 31671
rect 7932 31628 7984 31637
rect 8484 31628 8536 31680
rect 11520 31671 11572 31680
rect 11520 31637 11529 31671
rect 11529 31637 11563 31671
rect 11563 31637 11572 31671
rect 11520 31628 11572 31637
rect 13636 31628 13688 31680
rect 16120 31628 16172 31680
rect 4874 31526 4926 31578
rect 4938 31526 4990 31578
rect 5002 31526 5054 31578
rect 5066 31526 5118 31578
rect 5130 31526 5182 31578
rect 7380 31424 7432 31476
rect 11244 31424 11296 31476
rect 12072 31424 12124 31476
rect 14280 31424 14332 31476
rect 7932 31356 7984 31408
rect 7104 31288 7156 31340
rect 7564 31288 7616 31340
rect 8484 31331 8536 31340
rect 8484 31297 8518 31331
rect 8518 31297 8536 31331
rect 8484 31288 8536 31297
rect 9680 31331 9732 31340
rect 9680 31297 9689 31331
rect 9689 31297 9723 31331
rect 9723 31297 9732 31331
rect 9680 31288 9732 31297
rect 9956 31331 10008 31340
rect 9956 31297 9990 31331
rect 9990 31297 10008 31331
rect 9956 31288 10008 31297
rect 12348 31288 12400 31340
rect 12992 31331 13044 31340
rect 12992 31297 13001 31331
rect 13001 31297 13035 31331
rect 13035 31297 13044 31331
rect 12992 31288 13044 31297
rect 13728 31356 13780 31408
rect 14188 31356 14240 31408
rect 6092 31220 6144 31272
rect 7656 31263 7708 31272
rect 7656 31229 7665 31263
rect 7665 31229 7699 31263
rect 7699 31229 7708 31263
rect 7656 31220 7708 31229
rect 8024 31263 8076 31272
rect 8024 31229 8033 31263
rect 8033 31229 8067 31263
rect 8067 31229 8076 31263
rect 8024 31220 8076 31229
rect 13636 31288 13688 31340
rect 14096 31288 14148 31340
rect 15200 31331 15252 31340
rect 15200 31297 15209 31331
rect 15209 31297 15243 31331
rect 15243 31297 15252 31331
rect 15200 31288 15252 31297
rect 16304 31331 16356 31340
rect 16304 31297 16313 31331
rect 16313 31297 16347 31331
rect 16347 31297 16356 31331
rect 16304 31288 16356 31297
rect 6920 31152 6972 31204
rect 15384 31220 15436 31272
rect 6736 31127 6788 31136
rect 6736 31093 6745 31127
rect 6745 31093 6779 31127
rect 6779 31093 6788 31127
rect 6736 31084 6788 31093
rect 9404 31084 9456 31136
rect 11888 31084 11940 31136
rect 11980 31084 12032 31136
rect 15844 31152 15896 31204
rect 16304 31152 16356 31204
rect 15752 31084 15804 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 6092 30923 6144 30932
rect 6092 30889 6101 30923
rect 6101 30889 6135 30923
rect 6135 30889 6144 30923
rect 6092 30880 6144 30889
rect 8024 30880 8076 30932
rect 9864 30923 9916 30932
rect 9864 30889 9873 30923
rect 9873 30889 9907 30923
rect 9907 30889 9916 30923
rect 9864 30880 9916 30889
rect 9956 30880 10008 30932
rect 11888 30880 11940 30932
rect 6460 30676 6512 30728
rect 6920 30676 6972 30728
rect 7472 30719 7524 30728
rect 7472 30685 7481 30719
rect 7481 30685 7515 30719
rect 7515 30685 7524 30719
rect 7472 30676 7524 30685
rect 8484 30812 8536 30864
rect 9680 30812 9732 30864
rect 9956 30787 10008 30796
rect 9956 30753 9965 30787
rect 9965 30753 9999 30787
rect 9999 30753 10008 30787
rect 9956 30744 10008 30753
rect 10232 30744 10284 30796
rect 10692 30787 10744 30796
rect 10692 30753 10701 30787
rect 10701 30753 10735 30787
rect 10735 30753 10744 30787
rect 10692 30744 10744 30753
rect 7012 30608 7064 30660
rect 8392 30719 8444 30728
rect 8392 30685 8401 30719
rect 8401 30685 8435 30719
rect 8435 30685 8444 30719
rect 8392 30676 8444 30685
rect 8484 30719 8536 30728
rect 8484 30685 8493 30719
rect 8493 30685 8527 30719
rect 8527 30685 8536 30719
rect 8484 30676 8536 30685
rect 8852 30676 8904 30728
rect 9128 30719 9180 30728
rect 9128 30685 9137 30719
rect 9137 30685 9171 30719
rect 9171 30685 9180 30719
rect 9128 30676 9180 30685
rect 9220 30719 9272 30728
rect 9220 30685 9229 30719
rect 9229 30685 9263 30719
rect 9263 30685 9272 30719
rect 9220 30676 9272 30685
rect 9496 30719 9548 30728
rect 9496 30685 9505 30719
rect 9505 30685 9539 30719
rect 9539 30685 9548 30719
rect 9496 30676 9548 30685
rect 10140 30676 10192 30728
rect 12716 30744 12768 30796
rect 16304 30923 16356 30932
rect 16304 30889 16313 30923
rect 16313 30889 16347 30923
rect 16347 30889 16356 30923
rect 16304 30880 16356 30889
rect 14556 30812 14608 30864
rect 12624 30676 12676 30728
rect 14004 30676 14056 30728
rect 14372 30719 14424 30728
rect 14372 30685 14381 30719
rect 14381 30685 14415 30719
rect 14415 30685 14424 30719
rect 14372 30676 14424 30685
rect 8024 30583 8076 30592
rect 8024 30549 8033 30583
rect 8033 30549 8067 30583
rect 8067 30549 8076 30583
rect 8024 30540 8076 30549
rect 10416 30608 10468 30660
rect 11060 30608 11112 30660
rect 11796 30608 11848 30660
rect 12808 30651 12860 30660
rect 9404 30540 9456 30592
rect 9772 30540 9824 30592
rect 12808 30617 12817 30651
rect 12817 30617 12851 30651
rect 12851 30617 12860 30651
rect 12808 30608 12860 30617
rect 13084 30608 13136 30660
rect 14280 30608 14332 30660
rect 14648 30676 14700 30728
rect 14924 30719 14976 30728
rect 14924 30685 14933 30719
rect 14933 30685 14967 30719
rect 14967 30685 14976 30719
rect 14924 30676 14976 30685
rect 14832 30608 14884 30660
rect 12440 30540 12492 30592
rect 13268 30583 13320 30592
rect 13268 30549 13277 30583
rect 13277 30549 13311 30583
rect 13311 30549 13320 30583
rect 13268 30540 13320 30549
rect 4874 30438 4926 30490
rect 4938 30438 4990 30490
rect 5002 30438 5054 30490
rect 5066 30438 5118 30490
rect 5130 30438 5182 30490
rect 6736 30336 6788 30388
rect 6828 30336 6880 30388
rect 8484 30336 8536 30388
rect 9588 30336 9640 30388
rect 9864 30336 9916 30388
rect 10876 30336 10928 30388
rect 11520 30379 11572 30388
rect 11520 30345 11529 30379
rect 11529 30345 11563 30379
rect 11563 30345 11572 30379
rect 11520 30336 11572 30345
rect 11888 30379 11940 30388
rect 11888 30345 11897 30379
rect 11897 30345 11931 30379
rect 11931 30345 11940 30379
rect 11888 30336 11940 30345
rect 12348 30379 12400 30388
rect 12348 30345 12357 30379
rect 12357 30345 12391 30379
rect 12391 30345 12400 30379
rect 12348 30336 12400 30345
rect 13268 30336 13320 30388
rect 16212 30336 16264 30388
rect 5908 30243 5960 30252
rect 5908 30209 5917 30243
rect 5917 30209 5951 30243
rect 5951 30209 5960 30243
rect 5908 30200 5960 30209
rect 6184 30243 6236 30252
rect 6184 30209 6193 30243
rect 6193 30209 6227 30243
rect 6227 30209 6236 30243
rect 6184 30200 6236 30209
rect 6092 30132 6144 30184
rect 6460 30268 6512 30320
rect 8024 30268 8076 30320
rect 10140 30268 10192 30320
rect 10784 30268 10836 30320
rect 12808 30268 12860 30320
rect 7472 30200 7524 30252
rect 7932 30243 7984 30252
rect 7932 30209 7941 30243
rect 7941 30209 7975 30243
rect 7975 30209 7984 30243
rect 7932 30200 7984 30209
rect 10048 30200 10100 30252
rect 10600 30200 10652 30252
rect 13544 30268 13596 30320
rect 5540 30039 5592 30048
rect 5540 30005 5549 30039
rect 5549 30005 5583 30039
rect 5583 30005 5592 30039
rect 5540 29996 5592 30005
rect 7012 29996 7064 30048
rect 7748 30039 7800 30048
rect 7748 30005 7757 30039
rect 7757 30005 7791 30039
rect 7791 30005 7800 30039
rect 7748 29996 7800 30005
rect 8852 29996 8904 30048
rect 10692 30107 10744 30116
rect 10692 30073 10701 30107
rect 10701 30073 10735 30107
rect 10735 30073 10744 30107
rect 10692 30064 10744 30073
rect 9864 29996 9916 30048
rect 10324 30039 10376 30048
rect 10324 30005 10333 30039
rect 10333 30005 10367 30039
rect 10367 30005 10376 30039
rect 11336 30132 11388 30184
rect 10968 30107 11020 30116
rect 10968 30073 10977 30107
rect 10977 30073 11011 30107
rect 11011 30073 11020 30107
rect 10968 30064 11020 30073
rect 11060 30064 11112 30116
rect 12716 30132 12768 30184
rect 12348 30064 12400 30116
rect 14096 30200 14148 30252
rect 14280 30243 14332 30252
rect 14280 30209 14289 30243
rect 14289 30209 14323 30243
rect 14323 30209 14332 30243
rect 14280 30200 14332 30209
rect 13084 30132 13136 30184
rect 13176 30132 13228 30184
rect 14556 30243 14608 30252
rect 14556 30209 14565 30243
rect 14565 30209 14599 30243
rect 14599 30209 14608 30243
rect 14556 30200 14608 30209
rect 14464 30132 14516 30184
rect 14924 30243 14976 30252
rect 14924 30209 14933 30243
rect 14933 30209 14967 30243
rect 14967 30209 14976 30243
rect 14924 30200 14976 30209
rect 15016 30200 15068 30252
rect 15568 30200 15620 30252
rect 10324 29996 10376 30005
rect 12164 29996 12216 30048
rect 14096 29996 14148 30048
rect 15844 29996 15896 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 6092 29835 6144 29844
rect 6092 29801 6101 29835
rect 6101 29801 6135 29835
rect 6135 29801 6144 29835
rect 6092 29792 6144 29801
rect 7104 29835 7156 29844
rect 7104 29801 7113 29835
rect 7113 29801 7147 29835
rect 7147 29801 7156 29835
rect 7104 29792 7156 29801
rect 7380 29792 7432 29844
rect 7840 29792 7892 29844
rect 9496 29792 9548 29844
rect 9956 29835 10008 29844
rect 9956 29801 9965 29835
rect 9965 29801 9999 29835
rect 9999 29801 10008 29835
rect 9956 29792 10008 29801
rect 7196 29724 7248 29776
rect 9588 29724 9640 29776
rect 10324 29792 10376 29844
rect 10416 29792 10468 29844
rect 7748 29656 7800 29708
rect 8116 29699 8168 29708
rect 8116 29665 8125 29699
rect 8125 29665 8159 29699
rect 8159 29665 8168 29699
rect 8116 29656 8168 29665
rect 9956 29656 10008 29708
rect 10140 29656 10192 29708
rect 11244 29724 11296 29776
rect 11152 29656 11204 29708
rect 6184 29631 6236 29640
rect 6184 29597 6193 29631
rect 6193 29597 6227 29631
rect 6227 29597 6236 29631
rect 6184 29588 6236 29597
rect 6920 29631 6972 29640
rect 6920 29597 6929 29631
rect 6929 29597 6963 29631
rect 6963 29597 6972 29631
rect 6920 29588 6972 29597
rect 5724 29495 5776 29504
rect 5724 29461 5733 29495
rect 5733 29461 5767 29495
rect 5767 29461 5776 29495
rect 5724 29452 5776 29461
rect 6092 29452 6144 29504
rect 7104 29520 7156 29572
rect 8852 29588 8904 29640
rect 9220 29588 9272 29640
rect 9404 29588 9456 29640
rect 9588 29631 9640 29640
rect 9588 29597 9597 29631
rect 9597 29597 9631 29631
rect 9631 29597 9640 29631
rect 9588 29588 9640 29597
rect 9772 29588 9824 29640
rect 9864 29631 9916 29640
rect 9864 29597 9873 29631
rect 9873 29597 9907 29631
rect 9907 29597 9916 29631
rect 9864 29588 9916 29597
rect 10692 29588 10744 29640
rect 12992 29792 13044 29844
rect 14096 29792 14148 29844
rect 14832 29835 14884 29844
rect 14832 29801 14841 29835
rect 14841 29801 14875 29835
rect 14875 29801 14884 29835
rect 14832 29792 14884 29801
rect 15568 29835 15620 29844
rect 15568 29801 15577 29835
rect 15577 29801 15611 29835
rect 15611 29801 15620 29835
rect 15568 29792 15620 29801
rect 11796 29767 11848 29776
rect 11796 29733 11805 29767
rect 11805 29733 11839 29767
rect 11839 29733 11848 29767
rect 11796 29724 11848 29733
rect 12256 29724 12308 29776
rect 11428 29631 11480 29640
rect 11428 29597 11437 29631
rect 11437 29597 11471 29631
rect 11471 29597 11480 29631
rect 11428 29588 11480 29597
rect 11612 29631 11664 29640
rect 11612 29597 11621 29631
rect 11621 29597 11655 29631
rect 11655 29597 11664 29631
rect 11612 29588 11664 29597
rect 11704 29631 11756 29640
rect 11704 29597 11713 29631
rect 11713 29597 11747 29631
rect 11747 29597 11756 29631
rect 11704 29588 11756 29597
rect 12348 29656 12400 29708
rect 12716 29656 12768 29708
rect 13084 29656 13136 29708
rect 13268 29656 13320 29708
rect 14372 29656 14424 29708
rect 12164 29631 12216 29640
rect 12164 29597 12173 29631
rect 12173 29597 12207 29631
rect 12207 29597 12216 29631
rect 12164 29588 12216 29597
rect 13452 29520 13504 29572
rect 13544 29563 13596 29572
rect 13544 29529 13553 29563
rect 13553 29529 13587 29563
rect 13587 29529 13596 29563
rect 13544 29520 13596 29529
rect 13728 29563 13780 29572
rect 13728 29529 13737 29563
rect 13737 29529 13771 29563
rect 13771 29529 13780 29563
rect 13728 29520 13780 29529
rect 14832 29588 14884 29640
rect 15660 29656 15712 29708
rect 15292 29631 15344 29640
rect 15292 29597 15301 29631
rect 15301 29597 15335 29631
rect 15335 29597 15344 29631
rect 15292 29588 15344 29597
rect 15844 29631 15896 29640
rect 15844 29597 15853 29631
rect 15853 29597 15887 29631
rect 15887 29597 15896 29631
rect 15844 29588 15896 29597
rect 6736 29452 6788 29504
rect 6920 29452 6972 29504
rect 8668 29495 8720 29504
rect 8668 29461 8677 29495
rect 8677 29461 8711 29495
rect 8711 29461 8720 29495
rect 8668 29452 8720 29461
rect 9036 29495 9088 29504
rect 9036 29461 9045 29495
rect 9045 29461 9079 29495
rect 9079 29461 9088 29495
rect 9036 29452 9088 29461
rect 10324 29452 10376 29504
rect 10508 29452 10560 29504
rect 12532 29452 12584 29504
rect 12624 29495 12676 29504
rect 12624 29461 12633 29495
rect 12633 29461 12667 29495
rect 12667 29461 12676 29495
rect 12624 29452 12676 29461
rect 12900 29452 12952 29504
rect 13268 29452 13320 29504
rect 13636 29452 13688 29504
rect 14280 29452 14332 29504
rect 14556 29452 14608 29504
rect 4874 29350 4926 29402
rect 4938 29350 4990 29402
rect 5002 29350 5054 29402
rect 5066 29350 5118 29402
rect 5130 29350 5182 29402
rect 6644 29248 6696 29300
rect 6736 29248 6788 29300
rect 8392 29248 8444 29300
rect 8668 29248 8720 29300
rect 10876 29248 10928 29300
rect 11612 29248 11664 29300
rect 13636 29291 13688 29300
rect 13636 29257 13645 29291
rect 13645 29257 13679 29291
rect 13679 29257 13688 29291
rect 13636 29248 13688 29257
rect 14096 29248 14148 29300
rect 14648 29248 14700 29300
rect 5908 29180 5960 29232
rect 6828 29180 6880 29232
rect 5540 29112 5592 29164
rect 6644 29112 6696 29164
rect 6920 29155 6972 29164
rect 6920 29121 6929 29155
rect 6929 29121 6963 29155
rect 6963 29121 6972 29155
rect 6920 29112 6972 29121
rect 7932 29180 7984 29232
rect 9036 29180 9088 29232
rect 8944 29155 8996 29164
rect 8944 29121 8953 29155
rect 8953 29121 8987 29155
rect 8987 29121 8996 29155
rect 8944 29112 8996 29121
rect 10692 29180 10744 29232
rect 12624 29180 12676 29232
rect 13360 29180 13412 29232
rect 9588 29112 9640 29164
rect 10140 29112 10192 29164
rect 14464 29112 14516 29164
rect 14648 29155 14700 29164
rect 14648 29121 14657 29155
rect 14657 29121 14691 29155
rect 14691 29121 14700 29155
rect 14648 29112 14700 29121
rect 15476 29180 15528 29232
rect 15016 29155 15068 29164
rect 15016 29121 15025 29155
rect 15025 29121 15059 29155
rect 15059 29121 15068 29155
rect 15016 29112 15068 29121
rect 15292 29112 15344 29164
rect 15936 29248 15988 29300
rect 7196 28976 7248 29028
rect 7288 29019 7340 29028
rect 7288 28985 7297 29019
rect 7297 28985 7331 29019
rect 7331 28985 7340 29019
rect 7288 28976 7340 28985
rect 10784 28976 10836 29028
rect 12256 29087 12308 29096
rect 12256 29053 12265 29087
rect 12265 29053 12299 29087
rect 12299 29053 12308 29087
rect 12256 29044 12308 29053
rect 13728 29044 13780 29096
rect 15476 29044 15528 29096
rect 15936 29155 15988 29164
rect 15936 29121 15945 29155
rect 15945 29121 15979 29155
rect 15979 29121 15988 29155
rect 15936 29112 15988 29121
rect 16028 29155 16080 29164
rect 16028 29121 16037 29155
rect 16037 29121 16071 29155
rect 16071 29121 16080 29155
rect 16028 29112 16080 29121
rect 16304 29155 16356 29164
rect 16304 29121 16313 29155
rect 16313 29121 16347 29155
rect 16347 29121 16356 29155
rect 16304 29112 16356 29121
rect 13452 28976 13504 29028
rect 9036 28908 9088 28960
rect 9496 28908 9548 28960
rect 11152 28951 11204 28960
rect 11152 28917 11161 28951
rect 11161 28917 11195 28951
rect 11195 28917 11204 28951
rect 11152 28908 11204 28917
rect 11520 28951 11572 28960
rect 11520 28917 11529 28951
rect 11529 28917 11563 28951
rect 11563 28917 11572 28951
rect 11520 28908 11572 28917
rect 13728 28951 13780 28960
rect 13728 28917 13737 28951
rect 13737 28917 13771 28951
rect 13771 28917 13780 28951
rect 13728 28908 13780 28917
rect 14832 28976 14884 29028
rect 15200 28976 15252 29028
rect 15384 28976 15436 29028
rect 14556 28908 14608 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 6828 28747 6880 28756
rect 6828 28713 6837 28747
rect 6837 28713 6871 28747
rect 6871 28713 6880 28747
rect 6828 28704 6880 28713
rect 8944 28704 8996 28756
rect 9036 28704 9088 28756
rect 10048 28704 10100 28756
rect 10140 28747 10192 28756
rect 10140 28713 10149 28747
rect 10149 28713 10183 28747
rect 10183 28713 10192 28747
rect 10140 28704 10192 28713
rect 14464 28704 14516 28756
rect 15292 28704 15344 28756
rect 9220 28636 9272 28688
rect 7656 28568 7708 28620
rect 10232 28568 10284 28620
rect 13360 28636 13412 28688
rect 14556 28636 14608 28688
rect 5724 28500 5776 28552
rect 6828 28500 6880 28552
rect 7196 28543 7248 28552
rect 7196 28509 7205 28543
rect 7205 28509 7239 28543
rect 7239 28509 7248 28543
rect 7196 28500 7248 28509
rect 2964 28432 3016 28484
rect 8208 28432 8260 28484
rect 9036 28500 9088 28552
rect 10508 28500 10560 28552
rect 11520 28500 11572 28552
rect 11612 28543 11664 28552
rect 11612 28509 11621 28543
rect 11621 28509 11655 28543
rect 11655 28509 11664 28543
rect 11612 28500 11664 28509
rect 12256 28500 12308 28552
rect 14648 28568 14700 28620
rect 14832 28568 14884 28620
rect 14924 28611 14976 28620
rect 14924 28577 14933 28611
rect 14933 28577 14967 28611
rect 14967 28577 14976 28611
rect 14924 28568 14976 28577
rect 9404 28432 9456 28484
rect 9680 28432 9732 28484
rect 12992 28432 13044 28484
rect 14280 28543 14332 28552
rect 14280 28509 14289 28543
rect 14289 28509 14323 28543
rect 14323 28509 14332 28543
rect 14280 28500 14332 28509
rect 14372 28543 14424 28552
rect 14372 28509 14381 28543
rect 14381 28509 14415 28543
rect 14415 28509 14424 28543
rect 14372 28500 14424 28509
rect 15568 28500 15620 28552
rect 7564 28407 7616 28416
rect 7564 28373 7573 28407
rect 7573 28373 7607 28407
rect 7607 28373 7616 28407
rect 7564 28364 7616 28373
rect 8852 28364 8904 28416
rect 10508 28407 10560 28416
rect 10508 28373 10517 28407
rect 10517 28373 10551 28407
rect 10551 28373 10560 28407
rect 10508 28364 10560 28373
rect 12808 28364 12860 28416
rect 14740 28407 14792 28416
rect 14740 28373 14749 28407
rect 14749 28373 14783 28407
rect 14783 28373 14792 28407
rect 14740 28364 14792 28373
rect 15292 28432 15344 28484
rect 15384 28364 15436 28416
rect 4874 28262 4926 28314
rect 4938 28262 4990 28314
rect 5002 28262 5054 28314
rect 5066 28262 5118 28314
rect 5130 28262 5182 28314
rect 7840 28160 7892 28212
rect 9128 28160 9180 28212
rect 10508 28160 10560 28212
rect 7012 28092 7064 28144
rect 2596 28024 2648 28076
rect 3424 28024 3476 28076
rect 4712 28024 4764 28076
rect 6736 28067 6788 28076
rect 6736 28033 6745 28067
rect 6745 28033 6779 28067
rect 6779 28033 6788 28067
rect 6736 28024 6788 28033
rect 7104 28024 7156 28076
rect 7288 28067 7340 28076
rect 7288 28033 7297 28067
rect 7297 28033 7331 28067
rect 7331 28033 7340 28067
rect 7288 28024 7340 28033
rect 2780 27999 2832 28008
rect 2780 27965 2789 27999
rect 2789 27965 2823 27999
rect 2823 27965 2832 27999
rect 2780 27956 2832 27965
rect 7196 27999 7248 28008
rect 7196 27965 7205 27999
rect 7205 27965 7239 27999
rect 7239 27965 7248 27999
rect 7196 27956 7248 27965
rect 3792 27888 3844 27940
rect 5816 27888 5868 27940
rect 7840 28024 7892 28076
rect 8208 28024 8260 28076
rect 8760 28024 8812 28076
rect 3976 27820 4028 27872
rect 6920 27820 6972 27872
rect 9220 27999 9272 28008
rect 9220 27965 9229 27999
rect 9229 27965 9263 27999
rect 9263 27965 9272 27999
rect 9220 27956 9272 27965
rect 9956 27956 10008 28008
rect 10876 27956 10928 28008
rect 11152 27999 11204 28008
rect 11152 27965 11161 27999
rect 11161 27965 11195 27999
rect 11195 27965 11204 27999
rect 11152 27956 11204 27965
rect 10232 27820 10284 27872
rect 11980 28160 12032 28212
rect 12256 28092 12308 28144
rect 12992 28203 13044 28212
rect 12992 28169 13001 28203
rect 13001 28169 13035 28203
rect 13035 28169 13044 28203
rect 12992 28160 13044 28169
rect 13728 28160 13780 28212
rect 15292 28203 15344 28212
rect 15292 28169 15301 28203
rect 15301 28169 15335 28203
rect 15335 28169 15344 28203
rect 15292 28160 15344 28169
rect 12624 28067 12676 28076
rect 12624 28033 12642 28067
rect 12642 28033 12676 28067
rect 12624 28024 12676 28033
rect 12992 28024 13044 28076
rect 15108 28092 15160 28144
rect 13084 27956 13136 28008
rect 15568 28067 15620 28076
rect 15568 28033 15577 28067
rect 15577 28033 15611 28067
rect 15611 28033 15620 28067
rect 15568 28024 15620 28033
rect 15752 28067 15804 28076
rect 15752 28033 15761 28067
rect 15761 28033 15795 28067
rect 15795 28033 15804 28067
rect 15752 28024 15804 28033
rect 15844 28024 15896 28076
rect 16120 28024 16172 28076
rect 16304 28024 16356 28076
rect 15752 27888 15804 27940
rect 13544 27820 13596 27872
rect 14556 27863 14608 27872
rect 14556 27829 14565 27863
rect 14565 27829 14599 27863
rect 14599 27829 14608 27863
rect 14556 27820 14608 27829
rect 16212 27863 16264 27872
rect 16212 27829 16221 27863
rect 16221 27829 16255 27863
rect 16255 27829 16264 27863
rect 16212 27820 16264 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 7012 27616 7064 27668
rect 7380 27616 7432 27668
rect 11612 27616 11664 27668
rect 12256 27616 12308 27668
rect 7104 27548 7156 27600
rect 7840 27548 7892 27600
rect 8944 27591 8996 27600
rect 8944 27557 8953 27591
rect 8953 27557 8987 27591
rect 8987 27557 8996 27591
rect 8944 27548 8996 27557
rect 2780 27412 2832 27464
rect 3792 27455 3844 27464
rect 3792 27421 3801 27455
rect 3801 27421 3835 27455
rect 3835 27421 3844 27455
rect 3792 27412 3844 27421
rect 4160 27412 4212 27464
rect 5632 27412 5684 27464
rect 2412 27344 2464 27396
rect 4068 27344 4120 27396
rect 4620 27344 4672 27396
rect 6000 27344 6052 27396
rect 3332 27276 3384 27328
rect 3884 27319 3936 27328
rect 3884 27285 3893 27319
rect 3893 27285 3927 27319
rect 3927 27285 3936 27319
rect 3884 27276 3936 27285
rect 5264 27276 5316 27328
rect 6276 27276 6328 27328
rect 6736 27276 6788 27328
rect 8760 27455 8812 27464
rect 8760 27421 8769 27455
rect 8769 27421 8803 27455
rect 8803 27421 8812 27455
rect 8760 27412 8812 27421
rect 7288 27344 7340 27396
rect 9680 27412 9732 27464
rect 14280 27616 14332 27668
rect 14832 27616 14884 27668
rect 11152 27480 11204 27532
rect 10600 27344 10652 27396
rect 11888 27480 11940 27532
rect 12808 27523 12860 27532
rect 12808 27489 12817 27523
rect 12817 27489 12851 27523
rect 12851 27489 12860 27523
rect 12808 27480 12860 27489
rect 13452 27480 13504 27532
rect 12992 27412 13044 27464
rect 13544 27455 13596 27464
rect 13544 27421 13553 27455
rect 13553 27421 13587 27455
rect 13587 27421 13596 27455
rect 13544 27412 13596 27421
rect 14924 27412 14976 27464
rect 15752 27412 15804 27464
rect 7012 27319 7064 27328
rect 7012 27285 7021 27319
rect 7021 27285 7055 27319
rect 7055 27285 7064 27319
rect 7012 27276 7064 27285
rect 8484 27276 8536 27328
rect 11244 27319 11296 27328
rect 11244 27285 11253 27319
rect 11253 27285 11287 27319
rect 11287 27285 11296 27319
rect 11244 27276 11296 27285
rect 11888 27319 11940 27328
rect 11888 27285 11897 27319
rect 11897 27285 11931 27319
rect 11931 27285 11940 27319
rect 11888 27276 11940 27285
rect 14740 27344 14792 27396
rect 15384 27344 15436 27396
rect 15660 27344 15712 27396
rect 16028 27455 16080 27464
rect 16028 27421 16037 27455
rect 16037 27421 16071 27455
rect 16071 27421 16080 27455
rect 16028 27412 16080 27421
rect 16120 27412 16172 27464
rect 13176 27319 13228 27328
rect 13176 27285 13185 27319
rect 13185 27285 13219 27319
rect 13219 27285 13228 27319
rect 13176 27276 13228 27285
rect 15108 27276 15160 27328
rect 15292 27276 15344 27328
rect 15476 27319 15528 27328
rect 15476 27285 15485 27319
rect 15485 27285 15519 27319
rect 15519 27285 15528 27319
rect 15476 27276 15528 27285
rect 15568 27319 15620 27328
rect 15568 27285 15577 27319
rect 15577 27285 15611 27319
rect 15611 27285 15620 27319
rect 15568 27276 15620 27285
rect 4874 27174 4926 27226
rect 4938 27174 4990 27226
rect 5002 27174 5054 27226
rect 5066 27174 5118 27226
rect 5130 27174 5182 27226
rect 2136 27115 2188 27124
rect 2136 27081 2145 27115
rect 2145 27081 2179 27115
rect 2179 27081 2188 27115
rect 2872 27115 2924 27124
rect 2136 27072 2188 27081
rect 2320 27004 2372 27056
rect 2872 27081 2881 27115
rect 2881 27081 2915 27115
rect 2915 27081 2924 27115
rect 2872 27072 2924 27081
rect 2780 27047 2832 27056
rect 2780 27013 2789 27047
rect 2789 27013 2823 27047
rect 2823 27013 2832 27047
rect 2780 27004 2832 27013
rect 3884 27072 3936 27124
rect 4712 27072 4764 27124
rect 8208 27072 8260 27124
rect 8760 27072 8812 27124
rect 10232 27072 10284 27124
rect 12256 27072 12308 27124
rect 12624 27072 12676 27124
rect 14556 27072 14608 27124
rect 1676 26979 1728 26988
rect 1676 26945 1685 26979
rect 1685 26945 1719 26979
rect 1719 26945 1728 26979
rect 1676 26936 1728 26945
rect 2044 26911 2096 26920
rect 2044 26877 2053 26911
rect 2053 26877 2087 26911
rect 2087 26877 2096 26911
rect 2044 26868 2096 26877
rect 2228 26911 2280 26920
rect 4160 27004 4212 27056
rect 3516 26979 3568 26988
rect 3516 26945 3550 26979
rect 3550 26945 3568 26979
rect 3516 26936 3568 26945
rect 4988 26979 5040 26988
rect 4988 26945 5022 26979
rect 5022 26945 5040 26979
rect 4988 26936 5040 26945
rect 7104 27004 7156 27056
rect 7932 27004 7984 27056
rect 6920 26936 6972 26988
rect 9680 27004 9732 27056
rect 13268 27004 13320 27056
rect 15568 27004 15620 27056
rect 8116 26936 8168 26988
rect 2228 26877 2262 26911
rect 2262 26877 2280 26911
rect 2228 26868 2280 26877
rect 2964 26868 3016 26920
rect 2412 26843 2464 26852
rect 2412 26809 2421 26843
rect 2421 26809 2455 26843
rect 2455 26809 2464 26843
rect 2412 26800 2464 26809
rect 3056 26800 3108 26852
rect 3424 26732 3476 26784
rect 4160 26732 4212 26784
rect 13360 26936 13412 26988
rect 14740 26936 14792 26988
rect 14924 26979 14976 26988
rect 14924 26945 14933 26979
rect 14933 26945 14967 26979
rect 14967 26945 14976 26979
rect 14924 26936 14976 26945
rect 10232 26911 10284 26920
rect 10232 26877 10241 26911
rect 10241 26877 10275 26911
rect 10275 26877 10284 26911
rect 10232 26868 10284 26877
rect 10324 26868 10376 26920
rect 12624 26868 12676 26920
rect 5632 26732 5684 26784
rect 6092 26775 6144 26784
rect 6092 26741 6101 26775
rect 6101 26741 6135 26775
rect 6135 26741 6144 26775
rect 6092 26732 6144 26741
rect 7472 26732 7524 26784
rect 11244 26800 11296 26852
rect 9588 26775 9640 26784
rect 9588 26741 9597 26775
rect 9597 26741 9631 26775
rect 9631 26741 9640 26775
rect 9588 26732 9640 26741
rect 13452 26775 13504 26784
rect 13452 26741 13461 26775
rect 13461 26741 13495 26775
rect 13495 26741 13504 26775
rect 13452 26732 13504 26741
rect 15292 26732 15344 26784
rect 16304 26775 16356 26784
rect 16304 26741 16313 26775
rect 16313 26741 16347 26775
rect 16347 26741 16356 26775
rect 16304 26732 16356 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 2228 26528 2280 26580
rect 2596 26571 2648 26580
rect 2596 26537 2605 26571
rect 2605 26537 2639 26571
rect 2639 26537 2648 26571
rect 2596 26528 2648 26537
rect 2780 26528 2832 26580
rect 1676 26460 1728 26512
rect 3792 26528 3844 26580
rect 2412 26435 2464 26444
rect 2412 26401 2421 26435
rect 2421 26401 2455 26435
rect 2455 26401 2464 26435
rect 2412 26392 2464 26401
rect 2504 26392 2556 26444
rect 4252 26392 4304 26444
rect 2872 26231 2924 26240
rect 2872 26197 2881 26231
rect 2881 26197 2915 26231
rect 2915 26197 2924 26231
rect 2872 26188 2924 26197
rect 3148 26324 3200 26376
rect 3332 26367 3384 26376
rect 3332 26333 3341 26367
rect 3341 26333 3375 26367
rect 3375 26333 3384 26367
rect 3332 26324 3384 26333
rect 3884 26324 3936 26376
rect 4620 26503 4672 26512
rect 4620 26469 4629 26503
rect 4629 26469 4663 26503
rect 4663 26469 4672 26503
rect 4620 26460 4672 26469
rect 4804 26392 4856 26444
rect 5080 26435 5132 26444
rect 5080 26401 5089 26435
rect 5089 26401 5123 26435
rect 5123 26401 5132 26435
rect 5080 26392 5132 26401
rect 5540 26392 5592 26444
rect 5356 26324 5408 26376
rect 3516 26256 3568 26308
rect 3792 26256 3844 26308
rect 4436 26299 4488 26308
rect 4436 26265 4470 26299
rect 4470 26265 4488 26299
rect 4436 26256 4488 26265
rect 4804 26256 4856 26308
rect 5264 26256 5316 26308
rect 6000 26460 6052 26512
rect 6000 26324 6052 26376
rect 7288 26528 7340 26580
rect 8116 26528 8168 26580
rect 8484 26435 8536 26444
rect 8484 26401 8493 26435
rect 8493 26401 8527 26435
rect 8527 26401 8536 26435
rect 8484 26392 8536 26401
rect 9312 26528 9364 26580
rect 10232 26528 10284 26580
rect 10324 26571 10376 26580
rect 10324 26537 10333 26571
rect 10333 26537 10367 26571
rect 10367 26537 10376 26571
rect 10324 26528 10376 26537
rect 10784 26528 10836 26580
rect 14740 26528 14792 26580
rect 11980 26460 12032 26512
rect 14556 26460 14608 26512
rect 6276 26367 6328 26376
rect 6276 26333 6285 26367
rect 6285 26333 6319 26367
rect 6319 26333 6328 26367
rect 6276 26324 6328 26333
rect 5816 26299 5868 26308
rect 5816 26265 5825 26299
rect 5825 26265 5859 26299
rect 5859 26265 5868 26299
rect 5816 26256 5868 26265
rect 7104 26324 7156 26376
rect 7932 26324 7984 26376
rect 9588 26324 9640 26376
rect 9680 26324 9732 26376
rect 13176 26324 13228 26376
rect 3240 26188 3292 26240
rect 4252 26231 4304 26240
rect 4252 26197 4261 26231
rect 4261 26197 4295 26231
rect 4295 26197 4304 26231
rect 4252 26188 4304 26197
rect 4620 26188 4672 26240
rect 4988 26188 5040 26240
rect 5724 26188 5776 26240
rect 5908 26188 5960 26240
rect 6920 26256 6972 26308
rect 9772 26256 9824 26308
rect 10692 26299 10744 26308
rect 10692 26265 10726 26299
rect 10726 26265 10744 26299
rect 10692 26256 10744 26265
rect 13636 26392 13688 26444
rect 13820 26324 13872 26376
rect 7656 26188 7708 26240
rect 7840 26188 7892 26240
rect 11796 26231 11848 26240
rect 11796 26197 11805 26231
rect 11805 26197 11839 26231
rect 11839 26197 11848 26231
rect 11796 26188 11848 26197
rect 13360 26188 13412 26240
rect 13452 26188 13504 26240
rect 13912 26256 13964 26308
rect 15844 26367 15896 26376
rect 15844 26333 15853 26367
rect 15853 26333 15887 26367
rect 15887 26333 15896 26367
rect 15844 26324 15896 26333
rect 16120 26324 16172 26376
rect 14832 26231 14884 26240
rect 14832 26197 14841 26231
rect 14841 26197 14875 26231
rect 14875 26197 14884 26231
rect 14832 26188 14884 26197
rect 4874 26086 4926 26138
rect 4938 26086 4990 26138
rect 5002 26086 5054 26138
rect 5066 26086 5118 26138
rect 5130 26086 5182 26138
rect 3976 26027 4028 26036
rect 2412 25916 2464 25968
rect 3148 25916 3200 25968
rect 3332 25959 3384 25968
rect 3332 25925 3343 25959
rect 3343 25925 3384 25959
rect 3332 25916 3384 25925
rect 3976 25993 3985 26027
rect 3985 25993 4019 26027
rect 4019 25993 4028 26027
rect 3976 25984 4028 25993
rect 5356 26027 5408 26036
rect 5356 25993 5386 26027
rect 5386 25993 5408 26027
rect 5356 25984 5408 25993
rect 5540 25984 5592 26036
rect 6920 25984 6972 26036
rect 9220 25984 9272 26036
rect 9772 25984 9824 26036
rect 10692 25984 10744 26036
rect 10784 25984 10836 26036
rect 4712 25916 4764 25968
rect 6092 25916 6144 25968
rect 8208 25916 8260 25968
rect 12072 25916 12124 25968
rect 14832 25984 14884 26036
rect 15108 26027 15160 26036
rect 15108 25993 15117 26027
rect 15117 25993 15151 26027
rect 15151 25993 15160 26027
rect 15108 25984 15160 25993
rect 4804 25848 4856 25900
rect 5724 25848 5776 25900
rect 5816 25891 5868 25900
rect 5816 25857 5825 25891
rect 5825 25857 5859 25891
rect 5859 25857 5868 25891
rect 5816 25848 5868 25857
rect 7840 25848 7892 25900
rect 7932 25891 7984 25900
rect 7932 25857 7941 25891
rect 7941 25857 7975 25891
rect 7975 25857 7984 25891
rect 7932 25848 7984 25857
rect 3424 25712 3476 25764
rect 3240 25644 3292 25696
rect 4436 25780 4488 25832
rect 4068 25712 4120 25764
rect 5356 25780 5408 25832
rect 6552 25823 6604 25832
rect 6552 25789 6561 25823
rect 6561 25789 6595 25823
rect 6595 25789 6604 25823
rect 6552 25780 6604 25789
rect 9036 25848 9088 25900
rect 10416 25848 10468 25900
rect 11704 25848 11756 25900
rect 13360 25916 13412 25968
rect 14924 25916 14976 25968
rect 13268 25891 13320 25900
rect 13268 25857 13277 25891
rect 13277 25857 13311 25891
rect 13311 25857 13320 25891
rect 13268 25848 13320 25857
rect 13452 25848 13504 25900
rect 15200 25848 15252 25900
rect 15568 25891 15620 25900
rect 15568 25857 15577 25891
rect 15577 25857 15611 25891
rect 15611 25857 15620 25891
rect 15568 25848 15620 25857
rect 15660 25891 15712 25900
rect 15660 25857 15669 25891
rect 15669 25857 15703 25891
rect 15703 25857 15712 25891
rect 15660 25848 15712 25857
rect 10232 25823 10284 25832
rect 10232 25789 10241 25823
rect 10241 25789 10275 25823
rect 10275 25789 10284 25823
rect 10232 25780 10284 25789
rect 10600 25780 10652 25832
rect 7196 25712 7248 25764
rect 10968 25712 11020 25764
rect 14464 25780 14516 25832
rect 14832 25823 14884 25832
rect 14832 25789 14841 25823
rect 14841 25789 14875 25823
rect 14875 25789 14884 25823
rect 14832 25780 14884 25789
rect 14372 25712 14424 25764
rect 16212 25780 16264 25832
rect 4804 25644 4856 25696
rect 5816 25644 5868 25696
rect 11888 25644 11940 25696
rect 13912 25644 13964 25696
rect 14188 25644 14240 25696
rect 15844 25644 15896 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 6552 25440 6604 25492
rect 7012 25483 7064 25492
rect 7012 25449 7021 25483
rect 7021 25449 7055 25483
rect 7055 25449 7064 25483
rect 7012 25440 7064 25449
rect 7656 25483 7708 25492
rect 7656 25449 7665 25483
rect 7665 25449 7699 25483
rect 7699 25449 7708 25483
rect 7656 25440 7708 25449
rect 7840 25483 7892 25492
rect 7840 25449 7849 25483
rect 7849 25449 7883 25483
rect 7883 25449 7892 25483
rect 7840 25440 7892 25449
rect 8116 25483 8168 25492
rect 8116 25449 8125 25483
rect 8125 25449 8159 25483
rect 8159 25449 8168 25483
rect 8116 25440 8168 25449
rect 9036 25483 9088 25492
rect 9036 25449 9045 25483
rect 9045 25449 9079 25483
rect 9079 25449 9088 25483
rect 9036 25440 9088 25449
rect 11060 25483 11112 25492
rect 11060 25449 11069 25483
rect 11069 25449 11103 25483
rect 11103 25449 11112 25483
rect 11060 25440 11112 25449
rect 12624 25440 12676 25492
rect 14832 25440 14884 25492
rect 4620 25304 4672 25356
rect 6644 25304 6696 25356
rect 6828 25372 6880 25424
rect 8300 25372 8352 25424
rect 848 25236 900 25288
rect 7748 25304 7800 25356
rect 7196 25236 7248 25288
rect 7840 25236 7892 25288
rect 8024 25279 8076 25288
rect 8024 25245 8033 25279
rect 8033 25245 8067 25279
rect 8067 25245 8076 25279
rect 8024 25236 8076 25245
rect 5632 25211 5684 25220
rect 5632 25177 5641 25211
rect 5641 25177 5675 25211
rect 5675 25177 5684 25211
rect 5632 25168 5684 25177
rect 8208 25168 8260 25220
rect 3516 25100 3568 25152
rect 7932 25100 7984 25152
rect 8852 25304 8904 25356
rect 9312 25304 9364 25356
rect 11336 25347 11388 25356
rect 11336 25313 11345 25347
rect 11345 25313 11379 25347
rect 11379 25313 11388 25347
rect 11336 25304 11388 25313
rect 11980 25304 12032 25356
rect 13820 25304 13872 25356
rect 9220 25236 9272 25288
rect 11244 25279 11296 25288
rect 11244 25245 11253 25279
rect 11253 25245 11287 25279
rect 11287 25245 11296 25279
rect 11244 25236 11296 25245
rect 10140 25168 10192 25220
rect 12992 25279 13044 25288
rect 12992 25245 13001 25279
rect 13001 25245 13035 25279
rect 13035 25245 13044 25279
rect 12992 25236 13044 25245
rect 14096 25236 14148 25288
rect 14464 25304 14516 25356
rect 14004 25168 14056 25220
rect 12072 25100 12124 25152
rect 12164 25143 12216 25152
rect 12164 25109 12173 25143
rect 12173 25109 12207 25143
rect 12207 25109 12216 25143
rect 12164 25100 12216 25109
rect 12256 25100 12308 25152
rect 13360 25100 13412 25152
rect 14924 25347 14976 25356
rect 14924 25313 14933 25347
rect 14933 25313 14967 25347
rect 14967 25313 14976 25347
rect 14924 25304 14976 25313
rect 15200 25211 15252 25220
rect 15200 25177 15234 25211
rect 15234 25177 15252 25211
rect 15200 25168 15252 25177
rect 15568 25100 15620 25152
rect 16212 25100 16264 25152
rect 4874 24998 4926 25050
rect 4938 24998 4990 25050
rect 5002 24998 5054 25050
rect 5066 24998 5118 25050
rect 5130 24998 5182 25050
rect 2044 24939 2096 24948
rect 2044 24905 2053 24939
rect 2053 24905 2087 24939
rect 2087 24905 2096 24939
rect 2044 24896 2096 24905
rect 4620 24896 4672 24948
rect 7656 24896 7708 24948
rect 3608 24828 3660 24880
rect 2872 24760 2924 24812
rect 3424 24760 3476 24812
rect 3516 24803 3568 24812
rect 3516 24769 3525 24803
rect 3525 24769 3559 24803
rect 3559 24769 3568 24803
rect 3516 24760 3568 24769
rect 3976 24803 4028 24812
rect 3976 24769 3985 24803
rect 3985 24769 4019 24803
rect 4019 24769 4028 24803
rect 3976 24760 4028 24769
rect 4712 24828 4764 24880
rect 1860 24735 1912 24744
rect 1860 24701 1878 24735
rect 1878 24701 1912 24735
rect 1860 24692 1912 24701
rect 2596 24692 2648 24744
rect 3884 24735 3936 24744
rect 3884 24701 3893 24735
rect 3893 24701 3927 24735
rect 3927 24701 3936 24735
rect 3884 24692 3936 24701
rect 3792 24624 3844 24676
rect 4896 24692 4948 24744
rect 4620 24624 4672 24676
rect 5632 24803 5684 24812
rect 5632 24769 5641 24803
rect 5641 24769 5675 24803
rect 5675 24769 5684 24803
rect 5632 24760 5684 24769
rect 5816 24760 5868 24812
rect 7840 24828 7892 24880
rect 8116 24896 8168 24948
rect 9312 24939 9364 24948
rect 9312 24905 9321 24939
rect 9321 24905 9355 24939
rect 9355 24905 9364 24939
rect 9312 24896 9364 24905
rect 11336 24939 11388 24948
rect 11336 24905 11345 24939
rect 11345 24905 11379 24939
rect 11379 24905 11388 24939
rect 11336 24896 11388 24905
rect 12992 24896 13044 24948
rect 13360 24939 13412 24948
rect 13360 24905 13369 24939
rect 13369 24905 13403 24939
rect 13403 24905 13412 24939
rect 13360 24896 13412 24905
rect 13544 24896 13596 24948
rect 15752 24896 15804 24948
rect 7104 24803 7156 24812
rect 7104 24769 7138 24803
rect 7138 24769 7156 24803
rect 5816 24624 5868 24676
rect 6184 24624 6236 24676
rect 6276 24624 6328 24676
rect 7104 24760 7156 24769
rect 8668 24871 8720 24880
rect 8668 24837 8677 24871
rect 8677 24837 8711 24871
rect 8711 24837 8720 24871
rect 8668 24828 8720 24837
rect 9680 24760 9732 24812
rect 11244 24760 11296 24812
rect 11612 24760 11664 24812
rect 12348 24760 12400 24812
rect 8300 24692 8352 24744
rect 9312 24692 9364 24744
rect 11520 24735 11572 24744
rect 11520 24701 11529 24735
rect 11529 24701 11563 24735
rect 11563 24701 11572 24735
rect 11520 24692 11572 24701
rect 13728 24760 13780 24812
rect 12624 24692 12676 24744
rect 14280 24760 14332 24812
rect 14372 24803 14424 24812
rect 14372 24769 14381 24803
rect 14381 24769 14415 24803
rect 14415 24769 14424 24803
rect 14372 24760 14424 24769
rect 15016 24828 15068 24880
rect 14556 24803 14608 24812
rect 14556 24769 14565 24803
rect 14565 24769 14599 24803
rect 14599 24769 14608 24803
rect 14556 24760 14608 24769
rect 14924 24803 14976 24812
rect 14924 24769 14933 24803
rect 14933 24769 14967 24803
rect 14967 24769 14976 24803
rect 14924 24760 14976 24769
rect 16212 24828 16264 24880
rect 15476 24760 15528 24812
rect 1768 24556 1820 24608
rect 3424 24556 3476 24608
rect 4068 24556 4120 24608
rect 4712 24556 4764 24608
rect 5448 24599 5500 24608
rect 5448 24565 5457 24599
rect 5457 24565 5491 24599
rect 5491 24565 5500 24599
rect 5448 24556 5500 24565
rect 7748 24556 7800 24608
rect 8484 24556 8536 24608
rect 11428 24556 11480 24608
rect 12808 24556 12860 24608
rect 12992 24599 13044 24608
rect 12992 24565 13001 24599
rect 13001 24565 13035 24599
rect 13035 24565 13044 24599
rect 12992 24556 13044 24565
rect 13912 24667 13964 24676
rect 13912 24633 13921 24667
rect 13921 24633 13955 24667
rect 13955 24633 13964 24667
rect 13912 24624 13964 24633
rect 14096 24624 14148 24676
rect 14372 24624 14424 24676
rect 14740 24624 14792 24676
rect 14924 24624 14976 24676
rect 14648 24556 14700 24608
rect 15200 24556 15252 24608
rect 15292 24556 15344 24608
rect 15660 24556 15712 24608
rect 15844 24556 15896 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 1860 24352 1912 24404
rect 4252 24352 4304 24404
rect 4896 24352 4948 24404
rect 5356 24352 5408 24404
rect 3976 24284 4028 24336
rect 6184 24352 6236 24404
rect 7104 24352 7156 24404
rect 8852 24352 8904 24404
rect 10140 24395 10192 24404
rect 10140 24361 10149 24395
rect 10149 24361 10183 24395
rect 10183 24361 10192 24395
rect 10140 24352 10192 24361
rect 10232 24352 10284 24404
rect 10692 24352 10744 24404
rect 12256 24352 12308 24404
rect 13176 24352 13228 24404
rect 1400 24148 1452 24200
rect 1768 24191 1820 24200
rect 1768 24157 1802 24191
rect 1802 24157 1820 24191
rect 1768 24148 1820 24157
rect 2044 24148 2096 24200
rect 3056 24216 3108 24268
rect 2964 24191 3016 24200
rect 2964 24157 2973 24191
rect 2973 24157 3007 24191
rect 3007 24157 3016 24191
rect 2964 24148 3016 24157
rect 3148 24191 3200 24200
rect 3148 24157 3157 24191
rect 3157 24157 3191 24191
rect 3191 24157 3200 24191
rect 3148 24148 3200 24157
rect 3424 24191 3476 24200
rect 3424 24157 3463 24191
rect 3463 24157 3476 24191
rect 3424 24148 3476 24157
rect 3608 24191 3660 24200
rect 3608 24157 3617 24191
rect 3617 24157 3651 24191
rect 3651 24157 3660 24191
rect 3608 24148 3660 24157
rect 2596 24080 2648 24132
rect 3332 24080 3384 24132
rect 3056 24012 3108 24064
rect 3148 24012 3200 24064
rect 4068 24148 4120 24200
rect 4988 24259 5040 24268
rect 4988 24225 4997 24259
rect 4997 24225 5031 24259
rect 5031 24225 5040 24259
rect 4988 24216 5040 24225
rect 5448 24216 5500 24268
rect 5908 24216 5960 24268
rect 7380 24216 7432 24268
rect 5172 24080 5224 24132
rect 7564 24148 7616 24200
rect 8484 24191 8536 24200
rect 8484 24157 8502 24191
rect 8502 24157 8536 24191
rect 8484 24148 8536 24157
rect 9220 24148 9272 24200
rect 11060 24284 11112 24336
rect 11980 24327 12032 24336
rect 11980 24293 11989 24327
rect 11989 24293 12023 24327
rect 12023 24293 12032 24327
rect 11980 24284 12032 24293
rect 10600 24259 10652 24268
rect 10600 24225 10609 24259
rect 10609 24225 10643 24259
rect 10643 24225 10652 24259
rect 10600 24216 10652 24225
rect 10692 24259 10744 24268
rect 10692 24225 10701 24259
rect 10701 24225 10735 24259
rect 10735 24225 10744 24259
rect 10692 24216 10744 24225
rect 9864 24191 9916 24200
rect 9864 24157 9873 24191
rect 9873 24157 9907 24191
rect 9907 24157 9916 24191
rect 9864 24148 9916 24157
rect 11428 24216 11480 24268
rect 11336 24191 11388 24200
rect 11336 24157 11345 24191
rect 11345 24157 11379 24191
rect 11379 24157 11388 24191
rect 11336 24148 11388 24157
rect 12164 24216 12216 24268
rect 14280 24352 14332 24404
rect 14924 24352 14976 24404
rect 15476 24395 15528 24404
rect 15476 24361 15485 24395
rect 15485 24361 15519 24395
rect 15519 24361 15528 24395
rect 15476 24352 15528 24361
rect 15568 24395 15620 24404
rect 15568 24361 15577 24395
rect 15577 24361 15611 24395
rect 15611 24361 15620 24395
rect 15568 24352 15620 24361
rect 13636 24284 13688 24336
rect 14004 24284 14056 24336
rect 14556 24284 14608 24336
rect 15108 24284 15160 24336
rect 11704 24148 11756 24200
rect 12256 24148 12308 24200
rect 13636 24148 13688 24200
rect 13820 24216 13872 24268
rect 13912 24216 13964 24268
rect 14464 24191 14516 24200
rect 14464 24157 14473 24191
rect 14473 24157 14507 24191
rect 14507 24157 14516 24191
rect 14464 24148 14516 24157
rect 14924 24148 14976 24200
rect 15016 24191 15068 24200
rect 15016 24157 15025 24191
rect 15025 24157 15059 24191
rect 15059 24157 15068 24191
rect 15016 24148 15068 24157
rect 5540 24080 5592 24132
rect 6092 24123 6144 24132
rect 6092 24089 6101 24123
rect 6101 24089 6135 24123
rect 6135 24089 6144 24123
rect 6092 24080 6144 24089
rect 12532 24080 12584 24132
rect 12992 24080 13044 24132
rect 15568 24148 15620 24200
rect 16212 24148 16264 24200
rect 15384 24080 15436 24132
rect 15844 24123 15896 24132
rect 15844 24089 15853 24123
rect 15853 24089 15887 24123
rect 15887 24089 15896 24123
rect 15844 24080 15896 24089
rect 15936 24123 15988 24132
rect 15936 24089 15945 24123
rect 15945 24089 15979 24123
rect 15979 24089 15988 24123
rect 15936 24080 15988 24089
rect 16396 24080 16448 24132
rect 4068 24012 4120 24064
rect 5356 24012 5408 24064
rect 5448 24012 5500 24064
rect 6184 24012 6236 24064
rect 6276 24055 6328 24064
rect 6276 24021 6285 24055
rect 6285 24021 6319 24055
rect 6319 24021 6328 24055
rect 6276 24012 6328 24021
rect 9680 24055 9732 24064
rect 9680 24021 9689 24055
rect 9689 24021 9723 24055
rect 9723 24021 9732 24055
rect 9680 24012 9732 24021
rect 10968 24012 11020 24064
rect 11152 24012 11204 24064
rect 11336 24012 11388 24064
rect 11428 24055 11480 24064
rect 11428 24021 11437 24055
rect 11437 24021 11471 24055
rect 11471 24021 11480 24055
rect 11428 24012 11480 24021
rect 11704 24055 11756 24064
rect 11704 24021 11713 24055
rect 11713 24021 11747 24055
rect 11747 24021 11756 24055
rect 11704 24012 11756 24021
rect 14096 24055 14148 24064
rect 14096 24021 14105 24055
rect 14105 24021 14139 24055
rect 14139 24021 14148 24055
rect 14096 24012 14148 24021
rect 14188 24012 14240 24064
rect 4874 23910 4926 23962
rect 4938 23910 4990 23962
rect 5002 23910 5054 23962
rect 5066 23910 5118 23962
rect 5130 23910 5182 23962
rect 2964 23851 3016 23860
rect 2964 23817 2973 23851
rect 2973 23817 3007 23851
rect 3007 23817 3016 23851
rect 2964 23808 3016 23817
rect 10600 23851 10652 23860
rect 10600 23817 10609 23851
rect 10609 23817 10643 23851
rect 10643 23817 10652 23851
rect 10600 23808 10652 23817
rect 1400 23715 1452 23724
rect 1400 23681 1409 23715
rect 1409 23681 1443 23715
rect 1443 23681 1452 23715
rect 1400 23672 1452 23681
rect 1676 23715 1728 23724
rect 1676 23681 1710 23715
rect 1710 23681 1728 23715
rect 1676 23672 1728 23681
rect 2872 23715 2924 23724
rect 2872 23681 2881 23715
rect 2881 23681 2915 23715
rect 2915 23681 2924 23715
rect 2872 23672 2924 23681
rect 3056 23715 3108 23724
rect 3056 23681 3065 23715
rect 3065 23681 3099 23715
rect 3099 23681 3108 23715
rect 3056 23672 3108 23681
rect 3148 23715 3200 23724
rect 3148 23681 3157 23715
rect 3157 23681 3191 23715
rect 3191 23681 3200 23715
rect 3148 23672 3200 23681
rect 3332 23715 3384 23724
rect 3332 23681 3341 23715
rect 3341 23681 3375 23715
rect 3375 23681 3384 23715
rect 3332 23672 3384 23681
rect 3424 23715 3476 23724
rect 3424 23681 3433 23715
rect 3433 23681 3467 23715
rect 3467 23681 3476 23715
rect 3424 23672 3476 23681
rect 3700 23672 3752 23724
rect 4252 23715 4304 23724
rect 4252 23681 4261 23715
rect 4261 23681 4295 23715
rect 4295 23681 4304 23715
rect 4252 23672 4304 23681
rect 5632 23740 5684 23792
rect 9220 23740 9272 23792
rect 11520 23740 11572 23792
rect 11980 23740 12032 23792
rect 3608 23604 3660 23656
rect 4068 23604 4120 23656
rect 5356 23672 5408 23724
rect 10508 23672 10560 23724
rect 10600 23672 10652 23724
rect 11428 23672 11480 23724
rect 9220 23647 9272 23656
rect 9220 23613 9229 23647
rect 9229 23613 9263 23647
rect 9263 23613 9272 23647
rect 9220 23604 9272 23613
rect 10968 23604 11020 23656
rect 4804 23536 4856 23588
rect 11244 23536 11296 23588
rect 2964 23468 3016 23520
rect 3792 23511 3844 23520
rect 3792 23477 3801 23511
rect 3801 23477 3835 23511
rect 3835 23477 3844 23511
rect 3792 23468 3844 23477
rect 4068 23468 4120 23520
rect 5908 23468 5960 23520
rect 6276 23468 6328 23520
rect 9864 23468 9916 23520
rect 11060 23468 11112 23520
rect 11888 23715 11940 23724
rect 11888 23681 11897 23715
rect 11897 23681 11931 23715
rect 11931 23681 11940 23715
rect 11888 23672 11940 23681
rect 12072 23715 12124 23724
rect 12072 23681 12081 23715
rect 12081 23681 12115 23715
rect 12115 23681 12124 23715
rect 12072 23672 12124 23681
rect 12808 23808 12860 23860
rect 12992 23808 13044 23860
rect 13084 23851 13136 23860
rect 13084 23817 13093 23851
rect 13093 23817 13127 23851
rect 13127 23817 13136 23851
rect 13084 23808 13136 23817
rect 13820 23808 13872 23860
rect 15016 23851 15068 23860
rect 15016 23817 15025 23851
rect 15025 23817 15059 23851
rect 15059 23817 15068 23851
rect 15016 23808 15068 23817
rect 14096 23740 14148 23792
rect 14188 23740 14240 23792
rect 12532 23715 12584 23724
rect 12532 23681 12541 23715
rect 12541 23681 12575 23715
rect 12575 23681 12584 23715
rect 12532 23672 12584 23681
rect 12716 23715 12768 23724
rect 12716 23681 12725 23715
rect 12725 23681 12759 23715
rect 12759 23681 12768 23715
rect 12716 23672 12768 23681
rect 12808 23715 12860 23724
rect 12808 23681 12817 23715
rect 12817 23681 12851 23715
rect 12851 23681 12860 23715
rect 12808 23672 12860 23681
rect 13084 23672 13136 23724
rect 16488 23740 16540 23792
rect 15108 23715 15160 23724
rect 15108 23681 15117 23715
rect 15117 23681 15151 23715
rect 15151 23681 15160 23715
rect 15108 23672 15160 23681
rect 13176 23647 13228 23656
rect 13176 23613 13185 23647
rect 13185 23613 13219 23647
rect 13219 23613 13228 23647
rect 13176 23604 13228 23613
rect 12072 23536 12124 23588
rect 15200 23604 15252 23656
rect 15384 23715 15436 23724
rect 15384 23681 15393 23715
rect 15393 23681 15427 23715
rect 15427 23681 15436 23715
rect 15384 23672 15436 23681
rect 15568 23672 15620 23724
rect 15660 23604 15712 23656
rect 15936 23604 15988 23656
rect 16120 23604 16172 23656
rect 14280 23536 14332 23588
rect 15292 23468 15344 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 1676 23264 1728 23316
rect 2596 23307 2648 23316
rect 2596 23273 2605 23307
rect 2605 23273 2639 23307
rect 2639 23273 2648 23307
rect 2596 23264 2648 23273
rect 2964 23264 3016 23316
rect 8024 23307 8076 23316
rect 8024 23273 8033 23307
rect 8033 23273 8067 23307
rect 8067 23273 8076 23307
rect 8024 23264 8076 23273
rect 8668 23264 8720 23316
rect 2688 23196 2740 23248
rect 3056 23196 3108 23248
rect 2044 23128 2096 23180
rect 3332 23171 3384 23180
rect 3332 23137 3341 23171
rect 3341 23137 3375 23171
rect 3375 23137 3384 23171
rect 3332 23128 3384 23137
rect 8300 23128 8352 23180
rect 9496 23128 9548 23180
rect 10232 23264 10284 23316
rect 10508 23264 10560 23316
rect 11060 23264 11112 23316
rect 11244 23264 11296 23316
rect 11612 23264 11664 23316
rect 11888 23264 11940 23316
rect 12072 23264 12124 23316
rect 13452 23264 13504 23316
rect 13636 23264 13688 23316
rect 10140 23128 10192 23180
rect 2136 23060 2188 23112
rect 2320 23103 2372 23112
rect 2320 23069 2329 23103
rect 2329 23069 2363 23103
rect 2363 23069 2372 23103
rect 2320 23060 2372 23069
rect 2872 23060 2924 23112
rect 2964 23103 3016 23112
rect 2964 23069 2973 23103
rect 2973 23069 3007 23103
rect 3007 23069 3016 23103
rect 2964 23060 3016 23069
rect 3240 23103 3292 23112
rect 3240 23069 3249 23103
rect 3249 23069 3283 23103
rect 3283 23069 3292 23103
rect 3240 23060 3292 23069
rect 3792 23103 3844 23112
rect 3792 23069 3801 23103
rect 3801 23069 3835 23103
rect 3835 23069 3844 23103
rect 3792 23060 3844 23069
rect 2504 22924 2556 22976
rect 3056 22992 3108 23044
rect 4160 23103 4212 23112
rect 4160 23069 4169 23103
rect 4169 23069 4203 23103
rect 4203 23069 4212 23103
rect 4160 23060 4212 23069
rect 6184 23103 6236 23112
rect 6184 23069 6202 23103
rect 6202 23069 6236 23103
rect 6184 23060 6236 23069
rect 6368 23060 6420 23112
rect 4252 22992 4304 23044
rect 8576 23060 8628 23112
rect 9772 23060 9824 23112
rect 10692 23060 10744 23112
rect 10968 23103 11020 23112
rect 10968 23069 10977 23103
rect 10977 23069 11011 23103
rect 11011 23069 11020 23103
rect 10968 23060 11020 23069
rect 11612 23179 11664 23188
rect 11612 23145 11621 23179
rect 11621 23145 11655 23179
rect 11655 23145 11664 23179
rect 11612 23136 11664 23145
rect 11796 23128 11848 23180
rect 12072 23128 12124 23180
rect 13912 23196 13964 23248
rect 11244 23103 11296 23112
rect 11244 23069 11253 23103
rect 11253 23069 11287 23103
rect 11287 23069 11296 23103
rect 11244 23060 11296 23069
rect 11336 23103 11388 23112
rect 11336 23069 11345 23103
rect 11345 23069 11379 23103
rect 11379 23069 11388 23103
rect 11336 23060 11388 23069
rect 11980 23103 12032 23112
rect 11980 23069 11989 23103
rect 11989 23069 12023 23103
rect 12023 23069 12032 23103
rect 11980 23060 12032 23069
rect 12256 23103 12308 23112
rect 12256 23069 12265 23103
rect 12265 23069 12299 23103
rect 12299 23069 12308 23103
rect 12256 23060 12308 23069
rect 12440 23128 12492 23180
rect 12992 23128 13044 23180
rect 13452 23128 13504 23180
rect 12808 23060 12860 23112
rect 14096 23103 14148 23112
rect 14096 23069 14105 23103
rect 14105 23069 14139 23103
rect 14139 23069 14148 23103
rect 14096 23060 14148 23069
rect 14280 23103 14332 23112
rect 14280 23069 14289 23103
rect 14289 23069 14323 23103
rect 14323 23069 14332 23103
rect 14280 23060 14332 23069
rect 15476 23264 15528 23316
rect 14464 23103 14516 23112
rect 14464 23069 14473 23103
rect 14473 23069 14507 23103
rect 14507 23069 14516 23103
rect 14464 23060 14516 23069
rect 4620 22924 4672 22976
rect 4712 22924 4764 22976
rect 4804 22924 4856 22976
rect 5356 22924 5408 22976
rect 6920 22924 6972 22976
rect 8392 22992 8444 23044
rect 12164 22992 12216 23044
rect 12716 22992 12768 23044
rect 13912 22992 13964 23044
rect 9496 22967 9548 22976
rect 9496 22933 9505 22967
rect 9505 22933 9539 22967
rect 9539 22933 9548 22967
rect 9496 22924 9548 22933
rect 10600 22967 10652 22976
rect 10600 22933 10609 22967
rect 10609 22933 10643 22967
rect 10643 22933 10652 22967
rect 10600 22924 10652 22933
rect 11152 22924 11204 22976
rect 11980 22924 12032 22976
rect 13176 22924 13228 22976
rect 13360 22967 13412 22976
rect 13360 22933 13369 22967
rect 13369 22933 13403 22967
rect 13403 22933 13412 22967
rect 13360 22924 13412 22933
rect 14096 22924 14148 22976
rect 14832 22924 14884 22976
rect 15384 22924 15436 22976
rect 4874 22822 4926 22874
rect 4938 22822 4990 22874
rect 5002 22822 5054 22874
rect 5066 22822 5118 22874
rect 5130 22822 5182 22874
rect 2228 22720 2280 22772
rect 2504 22763 2556 22772
rect 2504 22729 2529 22763
rect 2529 22729 2556 22763
rect 2504 22720 2556 22729
rect 2872 22720 2924 22772
rect 3516 22720 3568 22772
rect 3792 22720 3844 22772
rect 5448 22652 5500 22704
rect 9772 22763 9824 22772
rect 9772 22729 9781 22763
rect 9781 22729 9815 22763
rect 9815 22729 9824 22763
rect 9772 22720 9824 22729
rect 3056 22627 3108 22636
rect 3056 22593 3065 22627
rect 3065 22593 3099 22627
rect 3099 22593 3108 22627
rect 3056 22584 3108 22593
rect 4068 22584 4120 22636
rect 4436 22584 4488 22636
rect 2412 22516 2464 22568
rect 3240 22516 3292 22568
rect 4712 22627 4764 22636
rect 4712 22593 4721 22627
rect 4721 22593 4755 22627
rect 4755 22593 4764 22627
rect 4712 22584 4764 22593
rect 5816 22627 5868 22636
rect 2320 22448 2372 22500
rect 4988 22516 5040 22568
rect 3148 22380 3200 22432
rect 4252 22448 4304 22500
rect 4712 22448 4764 22500
rect 5080 22448 5132 22500
rect 5816 22593 5825 22627
rect 5825 22593 5859 22627
rect 5859 22593 5868 22627
rect 5816 22584 5868 22593
rect 6460 22584 6512 22636
rect 8300 22652 8352 22704
rect 12164 22720 12216 22772
rect 11060 22652 11112 22704
rect 8484 22584 8536 22636
rect 10416 22627 10468 22636
rect 10416 22593 10425 22627
rect 10425 22593 10459 22627
rect 10459 22593 10468 22627
rect 10416 22584 10468 22593
rect 10600 22627 10652 22636
rect 10600 22593 10609 22627
rect 10609 22593 10643 22627
rect 10643 22593 10652 22627
rect 10600 22584 10652 22593
rect 10784 22627 10836 22636
rect 10784 22593 10793 22627
rect 10793 22593 10827 22627
rect 10827 22593 10836 22627
rect 10784 22584 10836 22593
rect 5540 22559 5592 22568
rect 5540 22525 5549 22559
rect 5549 22525 5583 22559
rect 5583 22525 5592 22559
rect 5540 22516 5592 22525
rect 5356 22448 5408 22500
rect 6276 22516 6328 22568
rect 8300 22516 8352 22568
rect 6184 22448 6236 22500
rect 4896 22423 4948 22432
rect 4896 22389 4905 22423
rect 4905 22389 4939 22423
rect 4939 22389 4948 22423
rect 4896 22380 4948 22389
rect 5632 22423 5684 22432
rect 5632 22389 5641 22423
rect 5641 22389 5675 22423
rect 5675 22389 5684 22423
rect 5632 22380 5684 22389
rect 10508 22516 10560 22568
rect 10968 22627 11020 22636
rect 10968 22593 10977 22627
rect 10977 22593 11011 22627
rect 11011 22593 11020 22627
rect 10968 22584 11020 22593
rect 11520 22627 11572 22636
rect 11520 22593 11529 22627
rect 11529 22593 11563 22627
rect 11563 22593 11572 22627
rect 11520 22584 11572 22593
rect 12992 22584 13044 22636
rect 15108 22720 15160 22772
rect 16028 22720 16080 22772
rect 15752 22695 15804 22704
rect 15752 22661 15761 22695
rect 15761 22661 15795 22695
rect 15795 22661 15804 22695
rect 15752 22652 15804 22661
rect 16488 22652 16540 22704
rect 9496 22448 9548 22500
rect 12440 22448 12492 22500
rect 9864 22423 9916 22432
rect 9864 22389 9873 22423
rect 9873 22389 9907 22423
rect 9907 22389 9916 22423
rect 9864 22380 9916 22389
rect 10048 22380 10100 22432
rect 11796 22380 11848 22432
rect 14556 22584 14608 22636
rect 16304 22584 16356 22636
rect 13912 22559 13964 22568
rect 13912 22525 13921 22559
rect 13921 22525 13955 22559
rect 13955 22525 13964 22559
rect 13912 22516 13964 22525
rect 13820 22448 13872 22500
rect 15016 22448 15068 22500
rect 14096 22380 14148 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 3332 22176 3384 22228
rect 4436 22176 4488 22228
rect 4988 22176 5040 22228
rect 8392 22176 8444 22228
rect 8484 22176 8536 22228
rect 10784 22176 10836 22228
rect 11612 22176 11664 22228
rect 13452 22176 13504 22228
rect 13636 22176 13688 22228
rect 14372 22176 14424 22228
rect 14924 22176 14976 22228
rect 4344 22108 4396 22160
rect 5080 22108 5132 22160
rect 6368 22108 6420 22160
rect 3332 22083 3384 22092
rect 3332 22049 3341 22083
rect 3341 22049 3375 22083
rect 3375 22049 3384 22083
rect 3332 22040 3384 22049
rect 3976 22015 4028 22024
rect 3976 21981 3985 22015
rect 3985 21981 4019 22015
rect 4019 21981 4028 22015
rect 3976 21972 4028 21981
rect 4620 22040 4672 22092
rect 5816 22040 5868 22092
rect 10600 22108 10652 22160
rect 11888 22108 11940 22160
rect 4804 21972 4856 22024
rect 5448 22015 5500 22024
rect 5448 21981 5457 22015
rect 5457 21981 5491 22015
rect 5491 21981 5500 22015
rect 6368 22015 6420 22024
rect 5448 21972 5500 21981
rect 6368 21981 6377 22015
rect 6377 21981 6411 22015
rect 6411 21981 6420 22015
rect 6368 21972 6420 21981
rect 9404 22040 9456 22092
rect 10416 22040 10468 22092
rect 6828 22015 6880 22024
rect 6828 21981 6837 22015
rect 6837 21981 6871 22015
rect 6871 21981 6880 22015
rect 6828 21972 6880 21981
rect 3884 21904 3936 21956
rect 4712 21904 4764 21956
rect 7012 21904 7064 21956
rect 7564 21904 7616 21956
rect 9312 21972 9364 22024
rect 7840 21904 7892 21956
rect 9496 21904 9548 21956
rect 9956 21972 10008 22024
rect 10324 21972 10376 22024
rect 12072 22040 12124 22092
rect 12440 22083 12492 22092
rect 12440 22049 12449 22083
rect 12449 22049 12483 22083
rect 12483 22049 12492 22083
rect 12440 22040 12492 22049
rect 12992 22108 13044 22160
rect 14188 22040 14240 22092
rect 14280 22040 14332 22092
rect 14740 22040 14792 22092
rect 11704 21972 11756 22024
rect 12256 22015 12308 22024
rect 12256 21981 12265 22015
rect 12265 21981 12299 22015
rect 12299 21981 12308 22015
rect 12256 21972 12308 21981
rect 13360 21972 13412 22024
rect 15108 21972 15160 22024
rect 15384 22015 15436 22024
rect 15384 21981 15393 22015
rect 15393 21981 15427 22015
rect 15427 21981 15436 22015
rect 15384 21972 15436 21981
rect 15936 21972 15988 22024
rect 16028 22015 16080 22024
rect 16028 21981 16037 22015
rect 16037 21981 16071 22015
rect 16071 21981 16080 22015
rect 16028 21972 16080 21981
rect 10232 21904 10284 21956
rect 4620 21879 4672 21888
rect 4620 21845 4629 21879
rect 4629 21845 4663 21879
rect 4663 21845 4672 21879
rect 4620 21836 4672 21845
rect 6736 21879 6788 21888
rect 6736 21845 6745 21879
rect 6745 21845 6779 21879
rect 6779 21845 6788 21879
rect 6736 21836 6788 21845
rect 9128 21836 9180 21888
rect 9864 21836 9916 21888
rect 10784 21836 10836 21888
rect 11520 21904 11572 21956
rect 11980 21904 12032 21956
rect 13268 21904 13320 21956
rect 14464 21904 14516 21956
rect 15292 21904 15344 21956
rect 15200 21879 15252 21888
rect 15200 21845 15209 21879
rect 15209 21845 15243 21879
rect 15243 21845 15252 21879
rect 15200 21836 15252 21845
rect 15844 21879 15896 21888
rect 15844 21845 15853 21879
rect 15853 21845 15887 21879
rect 15887 21845 15896 21879
rect 15844 21836 15896 21845
rect 16212 21879 16264 21888
rect 16212 21845 16221 21879
rect 16221 21845 16255 21879
rect 16255 21845 16264 21879
rect 16212 21836 16264 21845
rect 4874 21734 4926 21786
rect 4938 21734 4990 21786
rect 5002 21734 5054 21786
rect 5066 21734 5118 21786
rect 5130 21734 5182 21786
rect 848 21496 900 21548
rect 3608 21632 3660 21684
rect 3884 21675 3936 21684
rect 3884 21641 3893 21675
rect 3893 21641 3927 21675
rect 3927 21641 3936 21675
rect 3884 21632 3936 21641
rect 5264 21675 5316 21684
rect 5264 21641 5273 21675
rect 5273 21641 5307 21675
rect 5307 21641 5316 21675
rect 5264 21632 5316 21641
rect 5356 21675 5408 21684
rect 5356 21641 5365 21675
rect 5365 21641 5399 21675
rect 5399 21641 5408 21675
rect 5356 21632 5408 21641
rect 7564 21675 7616 21684
rect 7564 21641 7573 21675
rect 7573 21641 7607 21675
rect 7607 21641 7616 21675
rect 7564 21632 7616 21641
rect 10876 21675 10928 21684
rect 10876 21641 10885 21675
rect 10885 21641 10919 21675
rect 10919 21641 10928 21675
rect 10876 21632 10928 21641
rect 12072 21632 12124 21684
rect 12348 21632 12400 21684
rect 14096 21632 14148 21684
rect 14464 21632 14516 21684
rect 14556 21675 14608 21684
rect 14556 21641 14565 21675
rect 14565 21641 14599 21675
rect 14599 21641 14608 21675
rect 14556 21632 14608 21641
rect 16028 21632 16080 21684
rect 4988 21564 5040 21616
rect 5632 21564 5684 21616
rect 5816 21564 5868 21616
rect 6184 21564 6236 21616
rect 6828 21564 6880 21616
rect 7012 21564 7064 21616
rect 8208 21607 8260 21616
rect 8208 21573 8217 21607
rect 8217 21573 8251 21607
rect 8251 21573 8260 21607
rect 8208 21564 8260 21573
rect 10232 21564 10284 21616
rect 10416 21564 10468 21616
rect 11244 21564 11296 21616
rect 3148 21496 3200 21548
rect 3332 21496 3384 21548
rect 3884 21496 3936 21548
rect 4344 21539 4396 21548
rect 4344 21505 4353 21539
rect 4353 21505 4387 21539
rect 4387 21505 4396 21539
rect 4344 21496 4396 21505
rect 4436 21539 4488 21548
rect 4436 21505 4445 21539
rect 4445 21505 4479 21539
rect 4479 21505 4488 21539
rect 4436 21496 4488 21505
rect 4896 21539 4948 21548
rect 4896 21505 4905 21539
rect 4905 21505 4939 21539
rect 4939 21505 4948 21539
rect 4896 21496 4948 21505
rect 5080 21428 5132 21480
rect 5908 21539 5960 21548
rect 5908 21505 5917 21539
rect 5917 21505 5951 21539
rect 5951 21505 5960 21539
rect 5908 21496 5960 21505
rect 6644 21496 6696 21548
rect 6920 21539 6972 21548
rect 6920 21505 6929 21539
rect 6929 21505 6963 21539
rect 6963 21505 6972 21539
rect 6920 21496 6972 21505
rect 7840 21539 7892 21548
rect 7840 21505 7849 21539
rect 7849 21505 7883 21539
rect 7883 21505 7892 21539
rect 7840 21496 7892 21505
rect 9220 21496 9272 21548
rect 9772 21539 9824 21548
rect 9772 21505 9806 21539
rect 9806 21505 9824 21539
rect 9772 21496 9824 21505
rect 10784 21496 10836 21548
rect 11428 21496 11480 21548
rect 11520 21539 11572 21548
rect 11520 21505 11529 21539
rect 11529 21505 11563 21539
rect 11563 21505 11572 21539
rect 11520 21496 11572 21505
rect 11704 21539 11756 21548
rect 11704 21505 11713 21539
rect 11713 21505 11747 21539
rect 11747 21505 11756 21539
rect 11704 21496 11756 21505
rect 12256 21564 12308 21616
rect 14372 21564 14424 21616
rect 14740 21564 14792 21616
rect 12348 21506 12400 21558
rect 12624 21539 12676 21548
rect 12624 21505 12658 21539
rect 12658 21505 12676 21539
rect 12624 21496 12676 21505
rect 14924 21539 14976 21548
rect 14924 21505 14933 21539
rect 14933 21505 14967 21539
rect 14967 21505 14976 21539
rect 14924 21496 14976 21505
rect 15016 21539 15068 21548
rect 15016 21505 15025 21539
rect 15025 21505 15059 21539
rect 15059 21505 15068 21539
rect 15016 21496 15068 21505
rect 15568 21564 15620 21616
rect 8944 21471 8996 21480
rect 8944 21437 8953 21471
rect 8953 21437 8987 21471
rect 8987 21437 8996 21471
rect 8944 21428 8996 21437
rect 11152 21428 11204 21480
rect 11336 21428 11388 21480
rect 5264 21360 5316 21412
rect 11888 21471 11940 21480
rect 11888 21437 11897 21471
rect 11897 21437 11931 21471
rect 11931 21437 11940 21471
rect 11888 21428 11940 21437
rect 11980 21428 12032 21480
rect 15844 21496 15896 21548
rect 16028 21539 16080 21548
rect 16028 21505 16037 21539
rect 16037 21505 16071 21539
rect 16071 21505 16080 21539
rect 16028 21496 16080 21505
rect 3424 21292 3476 21344
rect 3884 21292 3936 21344
rect 4712 21292 4764 21344
rect 5632 21335 5684 21344
rect 5632 21301 5641 21335
rect 5641 21301 5675 21335
rect 5675 21301 5684 21335
rect 5632 21292 5684 21301
rect 5816 21292 5868 21344
rect 6552 21292 6604 21344
rect 8668 21292 8720 21344
rect 9496 21292 9548 21344
rect 16488 21428 16540 21480
rect 15384 21360 15436 21412
rect 15844 21360 15896 21412
rect 11888 21292 11940 21344
rect 13268 21292 13320 21344
rect 13820 21335 13872 21344
rect 13820 21301 13829 21335
rect 13829 21301 13863 21335
rect 13863 21301 13872 21335
rect 13820 21292 13872 21301
rect 14280 21292 14332 21344
rect 14924 21292 14976 21344
rect 16304 21292 16356 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 3332 21131 3384 21140
rect 3332 21097 3341 21131
rect 3341 21097 3375 21131
rect 3375 21097 3384 21131
rect 3332 21088 3384 21097
rect 3792 21131 3844 21140
rect 3792 21097 3801 21131
rect 3801 21097 3835 21131
rect 3835 21097 3844 21131
rect 3792 21088 3844 21097
rect 2044 21020 2096 21072
rect 2136 20952 2188 21004
rect 2780 20995 2832 21004
rect 2780 20961 2789 20995
rect 2789 20961 2823 20995
rect 2823 20961 2832 20995
rect 2780 20952 2832 20961
rect 2412 20884 2464 20936
rect 2228 20859 2280 20868
rect 2228 20825 2237 20859
rect 2237 20825 2271 20859
rect 2271 20825 2280 20859
rect 2228 20816 2280 20825
rect 2872 20884 2924 20936
rect 3424 20884 3476 20936
rect 2964 20816 3016 20868
rect 7288 21088 7340 21140
rect 8484 21088 8536 21140
rect 9772 21131 9824 21140
rect 9772 21097 9781 21131
rect 9781 21097 9815 21131
rect 9815 21097 9824 21131
rect 9772 21088 9824 21097
rect 11704 21088 11756 21140
rect 12348 21131 12400 21140
rect 12348 21097 12357 21131
rect 12357 21097 12391 21131
rect 12391 21097 12400 21131
rect 12348 21088 12400 21097
rect 12624 21088 12676 21140
rect 13728 21088 13780 21140
rect 15108 21088 15160 21140
rect 4804 21020 4856 21072
rect 4988 21020 5040 21072
rect 6276 21020 6328 21072
rect 6368 21020 6420 21072
rect 4344 20927 4396 20936
rect 4344 20893 4353 20927
rect 4353 20893 4387 20927
rect 4387 20893 4396 20927
rect 4344 20884 4396 20893
rect 4528 20927 4580 20936
rect 4528 20893 4537 20927
rect 4537 20893 4571 20927
rect 4571 20893 4580 20927
rect 4528 20884 4580 20893
rect 5080 20952 5132 21004
rect 6736 20995 6788 21004
rect 6736 20961 6745 20995
rect 6745 20961 6779 20995
rect 6779 20961 6788 20995
rect 6736 20952 6788 20961
rect 10140 21063 10192 21072
rect 10140 21029 10149 21063
rect 10149 21029 10183 21063
rect 10183 21029 10192 21063
rect 10140 21020 10192 21029
rect 10324 21020 10376 21072
rect 9312 20952 9364 21004
rect 4896 20884 4948 20936
rect 5264 20884 5316 20936
rect 6460 20884 6512 20936
rect 8300 20884 8352 20936
rect 8944 20927 8996 20936
rect 8944 20893 8953 20927
rect 8953 20893 8987 20927
rect 8987 20893 8996 20927
rect 8944 20884 8996 20893
rect 9956 20927 10008 20936
rect 9956 20893 9965 20927
rect 9965 20893 9999 20927
rect 9999 20893 10008 20927
rect 9956 20884 10008 20893
rect 10324 20884 10376 20936
rect 10600 20927 10652 20936
rect 10600 20893 10609 20927
rect 10609 20893 10643 20927
rect 10643 20893 10652 20927
rect 10600 20884 10652 20893
rect 10876 21020 10928 21072
rect 11612 21020 11664 21072
rect 10784 20884 10836 20936
rect 11704 20927 11756 20936
rect 11704 20893 11713 20927
rect 11713 20893 11747 20927
rect 11747 20893 11756 20927
rect 11704 20884 11756 20893
rect 11888 20927 11940 20936
rect 11888 20893 11897 20927
rect 11897 20893 11931 20927
rect 11931 20893 11940 20927
rect 11888 20884 11940 20893
rect 12164 20952 12216 21004
rect 12256 20884 12308 20936
rect 12808 21020 12860 21072
rect 12992 21020 13044 21072
rect 14372 21020 14424 21072
rect 13176 20995 13228 21004
rect 13176 20961 13185 20995
rect 13185 20961 13219 20995
rect 13219 20961 13228 20995
rect 13176 20952 13228 20961
rect 13268 20995 13320 21004
rect 13268 20961 13277 20995
rect 13277 20961 13311 20995
rect 13311 20961 13320 20995
rect 13268 20952 13320 20961
rect 12624 20927 12676 20936
rect 12624 20893 12633 20927
rect 12633 20893 12667 20927
rect 12667 20893 12676 20927
rect 12624 20884 12676 20893
rect 12900 20884 12952 20936
rect 13820 20884 13872 20936
rect 14188 20884 14240 20936
rect 14464 20884 14516 20936
rect 5356 20816 5408 20868
rect 1492 20791 1544 20800
rect 1492 20757 1501 20791
rect 1501 20757 1535 20791
rect 1535 20757 1544 20791
rect 1492 20748 1544 20757
rect 2412 20791 2464 20800
rect 2412 20757 2421 20791
rect 2421 20757 2455 20791
rect 2455 20757 2464 20791
rect 2412 20748 2464 20757
rect 4804 20748 4856 20800
rect 8852 20816 8904 20868
rect 10968 20816 11020 20868
rect 14004 20816 14056 20868
rect 11060 20748 11112 20800
rect 12440 20748 12492 20800
rect 12900 20748 12952 20800
rect 14372 20859 14424 20868
rect 14372 20825 14381 20859
rect 14381 20825 14415 20859
rect 14415 20825 14424 20859
rect 14372 20816 14424 20825
rect 15016 20816 15068 20868
rect 15936 20748 15988 20800
rect 4874 20646 4926 20698
rect 4938 20646 4990 20698
rect 5002 20646 5054 20698
rect 5066 20646 5118 20698
rect 5130 20646 5182 20698
rect 3148 20544 3200 20596
rect 4344 20544 4396 20596
rect 6460 20544 6512 20596
rect 8852 20587 8904 20596
rect 8852 20553 8861 20587
rect 8861 20553 8895 20587
rect 8895 20553 8904 20587
rect 8852 20544 8904 20553
rect 10324 20544 10376 20596
rect 11244 20544 11296 20596
rect 2412 20476 2464 20528
rect 3976 20476 4028 20528
rect 2872 20408 2924 20460
rect 1400 20340 1452 20392
rect 2964 20383 3016 20392
rect 2964 20349 2973 20383
rect 2973 20349 3007 20383
rect 3007 20349 3016 20383
rect 2964 20340 3016 20349
rect 3148 20408 3200 20460
rect 3608 20408 3660 20460
rect 4160 20451 4212 20460
rect 4160 20417 4169 20451
rect 4169 20417 4203 20451
rect 4203 20417 4212 20451
rect 4160 20408 4212 20417
rect 7288 20476 7340 20528
rect 9956 20476 10008 20528
rect 10508 20476 10560 20528
rect 4620 20408 4672 20460
rect 4068 20340 4120 20392
rect 8484 20408 8536 20460
rect 10416 20408 10468 20460
rect 5264 20383 5316 20392
rect 5264 20349 5273 20383
rect 5273 20349 5307 20383
rect 5307 20349 5316 20383
rect 5264 20340 5316 20349
rect 4896 20272 4948 20324
rect 6092 20340 6144 20392
rect 8300 20340 8352 20392
rect 8392 20340 8444 20392
rect 6644 20272 6696 20324
rect 10876 20383 10928 20392
rect 10876 20349 10885 20383
rect 10885 20349 10919 20383
rect 10919 20349 10928 20383
rect 10876 20340 10928 20349
rect 11060 20451 11112 20460
rect 11060 20417 11069 20451
rect 11069 20417 11103 20451
rect 11103 20417 11112 20451
rect 11060 20408 11112 20417
rect 11336 20476 11388 20528
rect 12164 20476 12216 20528
rect 12900 20451 12952 20460
rect 12900 20417 12909 20451
rect 12909 20417 12943 20451
rect 12943 20417 12952 20451
rect 12900 20408 12952 20417
rect 13176 20476 13228 20528
rect 14372 20544 14424 20596
rect 14832 20587 14884 20596
rect 14832 20553 14841 20587
rect 14841 20553 14875 20587
rect 14875 20553 14884 20587
rect 14832 20544 14884 20553
rect 15016 20544 15068 20596
rect 15108 20544 15160 20596
rect 14648 20476 14700 20528
rect 14740 20476 14792 20528
rect 12164 20340 12216 20392
rect 15384 20451 15436 20460
rect 15384 20417 15393 20451
rect 15393 20417 15427 20451
rect 15427 20417 15436 20451
rect 15384 20408 15436 20417
rect 15568 20451 15620 20460
rect 15568 20417 15577 20451
rect 15577 20417 15611 20451
rect 15611 20417 15620 20451
rect 15568 20408 15620 20417
rect 11060 20272 11112 20324
rect 3884 20247 3936 20256
rect 3884 20213 3893 20247
rect 3893 20213 3927 20247
rect 3927 20213 3936 20247
rect 3884 20204 3936 20213
rect 7932 20204 7984 20256
rect 10968 20204 11020 20256
rect 15476 20340 15528 20392
rect 15384 20272 15436 20324
rect 16028 20408 16080 20460
rect 16120 20451 16172 20460
rect 16120 20417 16129 20451
rect 16129 20417 16163 20451
rect 16163 20417 16172 20451
rect 16120 20408 16172 20417
rect 16304 20340 16356 20392
rect 14188 20204 14240 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 1400 20000 1452 20052
rect 2872 19932 2924 19984
rect 3608 20043 3660 20052
rect 3608 20009 3617 20043
rect 3617 20009 3651 20043
rect 3651 20009 3660 20043
rect 3608 20000 3660 20009
rect 4160 20043 4212 20052
rect 4160 20009 4169 20043
rect 4169 20009 4203 20043
rect 4203 20009 4212 20043
rect 4160 20000 4212 20009
rect 4344 20043 4396 20052
rect 4344 20009 4353 20043
rect 4353 20009 4387 20043
rect 4387 20009 4396 20043
rect 4344 20000 4396 20009
rect 4528 20000 4580 20052
rect 4804 20000 4856 20052
rect 6276 20000 6328 20052
rect 8208 20000 8260 20052
rect 10784 20000 10836 20052
rect 1400 19907 1452 19916
rect 1400 19873 1409 19907
rect 1409 19873 1443 19907
rect 1443 19873 1452 19907
rect 1400 19864 1452 19873
rect 1492 19796 1544 19848
rect 4712 19864 4764 19916
rect 5172 19864 5224 19916
rect 4252 19796 4304 19848
rect 4436 19839 4488 19848
rect 4436 19805 4445 19839
rect 4445 19805 4479 19839
rect 4479 19805 4488 19839
rect 4436 19796 4488 19805
rect 4896 19839 4948 19848
rect 4896 19805 4905 19839
rect 4905 19805 4939 19839
rect 4939 19805 4948 19839
rect 4896 19796 4948 19805
rect 8392 19864 8444 19916
rect 8760 19932 8812 19984
rect 9312 19932 9364 19984
rect 11520 20000 11572 20052
rect 9404 19864 9456 19916
rect 11244 19864 11296 19916
rect 12348 20000 12400 20052
rect 5448 19796 5500 19848
rect 5632 19839 5684 19848
rect 5632 19805 5666 19839
rect 5666 19805 5684 19839
rect 5632 19796 5684 19805
rect 4160 19728 4212 19780
rect 5816 19728 5868 19780
rect 3424 19660 3476 19712
rect 4344 19660 4396 19712
rect 5908 19660 5960 19712
rect 7840 19839 7892 19848
rect 7840 19805 7849 19839
rect 7849 19805 7883 19839
rect 7883 19805 7892 19839
rect 7840 19796 7892 19805
rect 7932 19839 7984 19848
rect 7932 19805 7941 19839
rect 7941 19805 7975 19839
rect 7975 19805 7984 19839
rect 7932 19796 7984 19805
rect 8668 19839 8720 19848
rect 8668 19805 8677 19839
rect 8677 19805 8711 19839
rect 8711 19805 8720 19839
rect 8668 19796 8720 19805
rect 8944 19839 8996 19848
rect 8944 19805 8953 19839
rect 8953 19805 8987 19839
rect 8987 19805 8996 19839
rect 8944 19796 8996 19805
rect 9864 19796 9916 19848
rect 8116 19728 8168 19780
rect 8852 19728 8904 19780
rect 9220 19771 9272 19780
rect 9220 19737 9229 19771
rect 9229 19737 9263 19771
rect 9263 19737 9272 19771
rect 9220 19728 9272 19737
rect 10048 19839 10100 19848
rect 10048 19805 10057 19839
rect 10057 19805 10091 19839
rect 10091 19805 10100 19839
rect 10048 19796 10100 19805
rect 10784 19796 10836 19848
rect 11060 19839 11112 19848
rect 11060 19805 11069 19839
rect 11069 19805 11103 19839
rect 11103 19805 11112 19839
rect 11060 19796 11112 19805
rect 11428 19839 11480 19848
rect 11428 19805 11437 19839
rect 11437 19805 11471 19839
rect 11471 19805 11480 19839
rect 11428 19796 11480 19805
rect 12256 19932 12308 19984
rect 12900 19932 12952 19984
rect 13084 19932 13136 19984
rect 14740 20000 14792 20052
rect 16120 20000 16172 20052
rect 10692 19728 10744 19780
rect 11704 19728 11756 19780
rect 14188 19796 14240 19848
rect 16304 19864 16356 19916
rect 13544 19728 13596 19780
rect 15660 19839 15712 19848
rect 15660 19805 15669 19839
rect 15669 19805 15703 19839
rect 15703 19805 15712 19839
rect 15660 19796 15712 19805
rect 15936 19839 15988 19848
rect 15936 19805 15945 19839
rect 15945 19805 15979 19839
rect 15979 19805 15988 19839
rect 15936 19796 15988 19805
rect 16212 19796 16264 19848
rect 14372 19771 14424 19780
rect 14372 19737 14406 19771
rect 14406 19737 14424 19771
rect 14372 19728 14424 19737
rect 8392 19660 8444 19712
rect 9496 19703 9548 19712
rect 9496 19669 9505 19703
rect 9505 19669 9539 19703
rect 9539 19669 9548 19703
rect 9496 19660 9548 19669
rect 10508 19660 10560 19712
rect 11060 19660 11112 19712
rect 11428 19660 11480 19712
rect 11612 19660 11664 19712
rect 13084 19660 13136 19712
rect 15200 19660 15252 19712
rect 16028 19660 16080 19712
rect 4874 19558 4926 19610
rect 4938 19558 4990 19610
rect 5002 19558 5054 19610
rect 5066 19558 5118 19610
rect 5130 19558 5182 19610
rect 3424 19456 3476 19508
rect 4160 19456 4212 19508
rect 4804 19456 4856 19508
rect 5264 19456 5316 19508
rect 3700 19388 3752 19440
rect 3976 19388 4028 19440
rect 6460 19456 6512 19508
rect 8392 19456 8444 19508
rect 10692 19499 10744 19508
rect 10692 19465 10701 19499
rect 10701 19465 10735 19499
rect 10735 19465 10744 19499
rect 10692 19456 10744 19465
rect 10876 19499 10928 19508
rect 10876 19465 10885 19499
rect 10885 19465 10919 19499
rect 10919 19465 10928 19499
rect 10876 19456 10928 19465
rect 11060 19456 11112 19508
rect 11612 19499 11664 19508
rect 11612 19465 11621 19499
rect 11621 19465 11655 19499
rect 11655 19465 11664 19499
rect 11612 19456 11664 19465
rect 14372 19456 14424 19508
rect 4068 19320 4120 19372
rect 4252 19363 4304 19372
rect 4252 19329 4261 19363
rect 4261 19329 4295 19363
rect 4295 19329 4304 19363
rect 4252 19320 4304 19329
rect 4712 19320 4764 19372
rect 5172 19363 5224 19372
rect 5172 19329 5181 19363
rect 5181 19329 5215 19363
rect 5215 19329 5224 19363
rect 5172 19320 5224 19329
rect 5908 19431 5960 19440
rect 5908 19397 5917 19431
rect 5917 19397 5951 19431
rect 5951 19397 5960 19431
rect 5908 19388 5960 19397
rect 4436 19252 4488 19304
rect 5816 19320 5868 19372
rect 7564 19320 7616 19372
rect 8668 19388 8720 19440
rect 9496 19388 9548 19440
rect 10692 19320 10744 19372
rect 12348 19388 12400 19440
rect 13176 19388 13228 19440
rect 13728 19388 13780 19440
rect 14556 19456 14608 19508
rect 11152 19320 11204 19372
rect 11336 19363 11388 19372
rect 11336 19329 11345 19363
rect 11345 19329 11379 19363
rect 11379 19329 11388 19363
rect 11336 19320 11388 19329
rect 6920 19295 6972 19304
rect 6920 19261 6929 19295
rect 6929 19261 6963 19295
rect 6963 19261 6972 19295
rect 6920 19252 6972 19261
rect 8300 19252 8352 19304
rect 10324 19252 10376 19304
rect 3976 19227 4028 19236
rect 3976 19193 3985 19227
rect 3985 19193 4019 19227
rect 4019 19193 4028 19227
rect 3976 19184 4028 19193
rect 4528 19184 4580 19236
rect 10048 19184 10100 19236
rect 10600 19184 10652 19236
rect 11704 19363 11756 19372
rect 11704 19329 11713 19363
rect 11713 19329 11747 19363
rect 11747 19329 11756 19363
rect 11704 19320 11756 19329
rect 11888 19363 11940 19372
rect 11888 19329 11897 19363
rect 11897 19329 11931 19363
rect 11931 19329 11940 19363
rect 11888 19320 11940 19329
rect 12164 19363 12216 19372
rect 12164 19329 12173 19363
rect 12173 19329 12207 19363
rect 12207 19329 12216 19363
rect 12164 19320 12216 19329
rect 12256 19363 12308 19372
rect 12256 19329 12265 19363
rect 12265 19329 12299 19363
rect 12299 19329 12308 19363
rect 12256 19320 12308 19329
rect 12716 19320 12768 19372
rect 13084 19295 13136 19304
rect 13084 19261 13093 19295
rect 13093 19261 13127 19295
rect 13127 19261 13136 19295
rect 13084 19252 13136 19261
rect 13912 19295 13964 19304
rect 13912 19261 13921 19295
rect 13921 19261 13955 19295
rect 13955 19261 13964 19295
rect 13912 19252 13964 19261
rect 14556 19363 14608 19372
rect 14556 19329 14565 19363
rect 14565 19329 14599 19363
rect 14599 19329 14608 19363
rect 14556 19320 14608 19329
rect 14924 19388 14976 19440
rect 15568 19388 15620 19440
rect 15016 19320 15068 19372
rect 14280 19252 14332 19304
rect 2320 19159 2372 19168
rect 2320 19125 2329 19159
rect 2329 19125 2363 19159
rect 2363 19125 2372 19159
rect 2320 19116 2372 19125
rect 2688 19116 2740 19168
rect 3148 19116 3200 19168
rect 4344 19116 4396 19168
rect 4712 19116 4764 19168
rect 6552 19116 6604 19168
rect 6644 19116 6696 19168
rect 8116 19116 8168 19168
rect 8760 19159 8812 19168
rect 8760 19125 8769 19159
rect 8769 19125 8803 19159
rect 8803 19125 8812 19159
rect 8760 19116 8812 19125
rect 9404 19116 9456 19168
rect 9956 19116 10008 19168
rect 12532 19159 12584 19168
rect 12532 19125 12541 19159
rect 12541 19125 12575 19159
rect 12575 19125 12584 19159
rect 12532 19116 12584 19125
rect 15108 19116 15160 19168
rect 15936 19116 15988 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 8852 18912 8904 18964
rect 9036 18912 9088 18964
rect 10048 18912 10100 18964
rect 10324 18912 10376 18964
rect 11704 18912 11756 18964
rect 11888 18955 11940 18964
rect 11888 18921 11897 18955
rect 11897 18921 11931 18955
rect 11931 18921 11940 18955
rect 11888 18912 11940 18921
rect 8576 18844 8628 18896
rect 9772 18844 9824 18896
rect 9956 18887 10008 18896
rect 9956 18853 9965 18887
rect 9965 18853 9999 18887
rect 9999 18853 10008 18887
rect 9956 18844 10008 18853
rect 9680 18819 9732 18828
rect 9680 18785 9689 18819
rect 9689 18785 9723 18819
rect 9723 18785 9732 18819
rect 9680 18776 9732 18785
rect 6920 18708 6972 18760
rect 8300 18751 8352 18760
rect 8300 18717 8309 18751
rect 8309 18717 8343 18751
rect 8343 18717 8352 18751
rect 8300 18708 8352 18717
rect 8484 18751 8536 18760
rect 8484 18717 8493 18751
rect 8493 18717 8527 18751
rect 8527 18717 8536 18751
rect 8484 18708 8536 18717
rect 9496 18708 9548 18760
rect 9588 18751 9640 18760
rect 9588 18717 9597 18751
rect 9597 18717 9631 18751
rect 9631 18717 9640 18751
rect 9588 18708 9640 18717
rect 10416 18708 10468 18760
rect 11152 18844 11204 18896
rect 10876 18776 10928 18828
rect 6000 18615 6052 18624
rect 6000 18581 6009 18615
rect 6009 18581 6043 18615
rect 6043 18581 6052 18615
rect 6000 18572 6052 18581
rect 7012 18640 7064 18692
rect 8208 18640 8260 18692
rect 9128 18683 9180 18692
rect 9128 18649 9146 18683
rect 9146 18649 9180 18683
rect 9128 18640 9180 18649
rect 9312 18640 9364 18692
rect 9956 18640 10008 18692
rect 10600 18640 10652 18692
rect 11060 18708 11112 18760
rect 11244 18751 11296 18760
rect 11244 18717 11253 18751
rect 11253 18717 11287 18751
rect 11287 18717 11296 18751
rect 11244 18708 11296 18717
rect 11428 18640 11480 18692
rect 7104 18572 7156 18624
rect 7840 18572 7892 18624
rect 8300 18572 8352 18624
rect 8668 18572 8720 18624
rect 9772 18572 9824 18624
rect 10692 18572 10744 18624
rect 10876 18572 10928 18624
rect 11612 18708 11664 18760
rect 12624 18912 12676 18964
rect 14096 18912 14148 18964
rect 15016 18912 15068 18964
rect 13912 18844 13964 18896
rect 15384 18912 15436 18964
rect 15200 18844 15252 18896
rect 12256 18751 12308 18760
rect 12256 18717 12265 18751
rect 12265 18717 12299 18751
rect 12299 18717 12308 18751
rect 12256 18708 12308 18717
rect 12532 18751 12584 18760
rect 12532 18717 12566 18751
rect 12566 18717 12584 18751
rect 12532 18708 12584 18717
rect 13912 18751 13964 18760
rect 13912 18717 13921 18751
rect 13921 18717 13955 18751
rect 13955 18717 13964 18751
rect 13912 18708 13964 18717
rect 14648 18708 14700 18760
rect 14740 18751 14792 18760
rect 14740 18717 14749 18751
rect 14749 18717 14783 18751
rect 14783 18717 14792 18751
rect 14740 18708 14792 18717
rect 15108 18708 15160 18760
rect 15476 18776 15528 18828
rect 15384 18751 15436 18760
rect 15384 18717 15393 18751
rect 15393 18717 15427 18751
rect 15427 18717 15436 18751
rect 15384 18708 15436 18717
rect 15568 18751 15620 18760
rect 15568 18717 15577 18751
rect 15577 18717 15611 18751
rect 15611 18717 15620 18751
rect 15568 18708 15620 18717
rect 16120 18708 16172 18760
rect 16304 18708 16356 18760
rect 11704 18615 11756 18624
rect 11704 18581 11713 18615
rect 11713 18581 11747 18615
rect 11747 18581 11756 18615
rect 11704 18572 11756 18581
rect 13268 18572 13320 18624
rect 15752 18640 15804 18692
rect 15936 18683 15988 18692
rect 15936 18649 15945 18683
rect 15945 18649 15979 18683
rect 15979 18649 15988 18683
rect 15936 18640 15988 18649
rect 16028 18683 16080 18692
rect 16028 18649 16037 18683
rect 16037 18649 16071 18683
rect 16071 18649 16080 18683
rect 16028 18640 16080 18649
rect 4874 18470 4926 18522
rect 4938 18470 4990 18522
rect 5002 18470 5054 18522
rect 5066 18470 5118 18522
rect 5130 18470 5182 18522
rect 3976 18368 4028 18420
rect 3240 18300 3292 18352
rect 3792 18300 3844 18352
rect 4160 18300 4212 18352
rect 2412 18232 2464 18284
rect 3056 18232 3108 18284
rect 7932 18368 7984 18420
rect 8484 18411 8536 18420
rect 8484 18377 8493 18411
rect 8493 18377 8527 18411
rect 8527 18377 8536 18411
rect 8484 18368 8536 18377
rect 9128 18368 9180 18420
rect 4988 18232 5040 18284
rect 5172 18232 5224 18284
rect 6000 18232 6052 18284
rect 6644 18232 6696 18284
rect 7012 18300 7064 18352
rect 7380 18343 7432 18352
rect 7380 18309 7414 18343
rect 7414 18309 7432 18343
rect 7380 18300 7432 18309
rect 8392 18300 8444 18352
rect 9588 18300 9640 18352
rect 10140 18411 10192 18420
rect 10140 18377 10149 18411
rect 10149 18377 10183 18411
rect 10183 18377 10192 18411
rect 10140 18368 10192 18377
rect 10508 18368 10560 18420
rect 13912 18368 13964 18420
rect 14188 18411 14240 18420
rect 14188 18377 14197 18411
rect 14197 18377 14231 18411
rect 14231 18377 14240 18411
rect 14188 18368 14240 18377
rect 15384 18368 15436 18420
rect 10324 18300 10376 18352
rect 6920 18232 6972 18284
rect 7748 18232 7800 18284
rect 2136 18028 2188 18080
rect 8760 18096 8812 18148
rect 9680 18232 9732 18284
rect 9864 18232 9916 18284
rect 9864 18096 9916 18148
rect 9404 18071 9456 18080
rect 9404 18037 9413 18071
rect 9413 18037 9447 18071
rect 9447 18037 9456 18071
rect 9404 18028 9456 18037
rect 9588 18028 9640 18080
rect 10600 18275 10652 18284
rect 10600 18241 10609 18275
rect 10609 18241 10643 18275
rect 10643 18241 10652 18275
rect 10600 18232 10652 18241
rect 11520 18232 11572 18284
rect 12256 18300 12308 18352
rect 12164 18275 12216 18284
rect 12164 18241 12198 18275
rect 12198 18241 12216 18275
rect 12164 18232 12216 18241
rect 14280 18232 14332 18284
rect 15752 18300 15804 18352
rect 14556 18232 14608 18284
rect 15660 18232 15712 18284
rect 15844 18232 15896 18284
rect 10692 18164 10744 18216
rect 14096 18096 14148 18148
rect 10600 18028 10652 18080
rect 10968 18028 11020 18080
rect 13360 18071 13412 18080
rect 13360 18037 13369 18071
rect 13369 18037 13403 18071
rect 13403 18037 13412 18071
rect 13360 18028 13412 18037
rect 15384 18028 15436 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 1952 17824 2004 17876
rect 2872 17824 2924 17876
rect 3332 17824 3384 17876
rect 4620 17824 4672 17876
rect 5356 17867 5408 17876
rect 5356 17833 5365 17867
rect 5365 17833 5399 17867
rect 5399 17833 5408 17867
rect 5356 17824 5408 17833
rect 7380 17824 7432 17876
rect 7564 17867 7616 17876
rect 7564 17833 7573 17867
rect 7573 17833 7607 17867
rect 7607 17833 7616 17867
rect 7564 17824 7616 17833
rect 10232 17867 10284 17876
rect 10232 17833 10241 17867
rect 10241 17833 10275 17867
rect 10275 17833 10284 17867
rect 10232 17824 10284 17833
rect 12164 17824 12216 17876
rect 12348 17824 12400 17876
rect 2964 17756 3016 17808
rect 3792 17756 3844 17808
rect 8760 17756 8812 17808
rect 14556 17824 14608 17876
rect 112 17688 164 17740
rect 2412 17663 2464 17672
rect 2412 17629 2421 17663
rect 2421 17629 2455 17663
rect 2455 17629 2464 17663
rect 2412 17620 2464 17629
rect 1768 17595 1820 17604
rect 1768 17561 1777 17595
rect 1777 17561 1811 17595
rect 1811 17561 1820 17595
rect 1768 17552 1820 17561
rect 2320 17552 2372 17604
rect 2688 17663 2740 17672
rect 2688 17629 2697 17663
rect 2697 17629 2731 17663
rect 2731 17629 2740 17663
rect 2688 17620 2740 17629
rect 3056 17620 3108 17672
rect 3332 17620 3384 17672
rect 3424 17663 3476 17672
rect 3424 17629 3433 17663
rect 3433 17629 3467 17663
rect 3467 17629 3476 17663
rect 3424 17620 3476 17629
rect 3516 17552 3568 17604
rect 3792 17663 3844 17672
rect 3792 17629 3801 17663
rect 3801 17629 3835 17663
rect 3835 17629 3844 17663
rect 3792 17620 3844 17629
rect 3884 17663 3936 17672
rect 3884 17629 3893 17663
rect 3893 17629 3927 17663
rect 3927 17629 3936 17663
rect 3884 17620 3936 17629
rect 4988 17620 5040 17672
rect 5172 17663 5224 17672
rect 5172 17629 5181 17663
rect 5181 17629 5215 17663
rect 5215 17629 5224 17663
rect 5172 17620 5224 17629
rect 4068 17552 4120 17604
rect 1400 17527 1452 17536
rect 1400 17493 1409 17527
rect 1409 17493 1443 17527
rect 1443 17493 1452 17527
rect 1400 17484 1452 17493
rect 1584 17527 1636 17536
rect 1584 17493 1611 17527
rect 1611 17493 1636 17527
rect 1584 17484 1636 17493
rect 1860 17527 1912 17536
rect 1860 17493 1869 17527
rect 1869 17493 1903 17527
rect 1903 17493 1912 17527
rect 1860 17484 1912 17493
rect 2412 17484 2464 17536
rect 2504 17527 2556 17536
rect 2504 17493 2513 17527
rect 2513 17493 2547 17527
rect 2547 17493 2556 17527
rect 2504 17484 2556 17493
rect 3148 17527 3200 17536
rect 3148 17493 3157 17527
rect 3157 17493 3191 17527
rect 3191 17493 3200 17527
rect 3148 17484 3200 17493
rect 3424 17484 3476 17536
rect 5172 17484 5224 17536
rect 6092 17484 6144 17536
rect 7840 17663 7892 17672
rect 7840 17629 7849 17663
rect 7849 17629 7883 17663
rect 7883 17629 7892 17663
rect 7840 17620 7892 17629
rect 7932 17663 7984 17672
rect 7932 17629 7941 17663
rect 7941 17629 7975 17663
rect 7975 17629 7984 17663
rect 7932 17620 7984 17629
rect 8300 17620 8352 17672
rect 8392 17663 8444 17672
rect 8392 17629 8401 17663
rect 8401 17629 8435 17663
rect 8435 17629 8444 17663
rect 8392 17620 8444 17629
rect 8668 17663 8720 17672
rect 8668 17629 8677 17663
rect 8677 17629 8711 17663
rect 8711 17629 8720 17663
rect 8668 17620 8720 17629
rect 11704 17688 11756 17740
rect 13360 17620 13412 17672
rect 8852 17552 8904 17604
rect 12900 17552 12952 17604
rect 13636 17663 13688 17672
rect 13636 17629 13645 17663
rect 13645 17629 13679 17663
rect 13679 17629 13688 17663
rect 13636 17620 13688 17629
rect 13912 17663 13964 17672
rect 13912 17629 13921 17663
rect 13921 17629 13955 17663
rect 13955 17629 13964 17663
rect 13912 17620 13964 17629
rect 14096 17663 14148 17672
rect 14096 17629 14105 17663
rect 14105 17629 14139 17663
rect 14139 17629 14148 17663
rect 14096 17620 14148 17629
rect 14280 17620 14332 17672
rect 15108 17824 15160 17876
rect 14832 17756 14884 17808
rect 14924 17620 14976 17672
rect 15568 17688 15620 17740
rect 16212 17688 16264 17740
rect 16304 17663 16356 17672
rect 16304 17629 16313 17663
rect 16313 17629 16347 17663
rect 16347 17629 16356 17663
rect 16304 17620 16356 17629
rect 15292 17595 15344 17604
rect 15292 17561 15301 17595
rect 15301 17561 15335 17595
rect 15335 17561 15344 17595
rect 15292 17552 15344 17561
rect 15660 17552 15712 17604
rect 15844 17552 15896 17604
rect 15016 17484 15068 17536
rect 16028 17484 16080 17536
rect 16304 17484 16356 17536
rect 4874 17382 4926 17434
rect 4938 17382 4990 17434
rect 5002 17382 5054 17434
rect 5066 17382 5118 17434
rect 5130 17382 5182 17434
rect 2964 17323 3016 17332
rect 2964 17289 2973 17323
rect 2973 17289 3007 17323
rect 3007 17289 3016 17323
rect 2964 17280 3016 17289
rect 8392 17280 8444 17332
rect 1400 17144 1452 17196
rect 1860 17187 1912 17196
rect 1860 17153 1894 17187
rect 1894 17153 1912 17187
rect 1860 17144 1912 17153
rect 3148 17187 3200 17196
rect 3148 17153 3157 17187
rect 3157 17153 3191 17187
rect 3191 17153 3200 17187
rect 3148 17144 3200 17153
rect 5080 17212 5132 17264
rect 3516 17144 3568 17196
rect 3700 17187 3752 17196
rect 3700 17153 3734 17187
rect 3734 17153 3752 17187
rect 3700 17144 3752 17153
rect 5356 17255 5408 17264
rect 5356 17221 5381 17255
rect 5381 17221 5408 17255
rect 5356 17212 5408 17221
rect 6276 17212 6328 17264
rect 5632 17187 5684 17196
rect 5632 17153 5641 17187
rect 5641 17153 5675 17187
rect 5675 17153 5684 17187
rect 5632 17144 5684 17153
rect 5908 17187 5960 17196
rect 5908 17153 5917 17187
rect 5917 17153 5951 17187
rect 5951 17153 5960 17187
rect 5908 17144 5960 17153
rect 8944 17280 8996 17332
rect 9312 17280 9364 17332
rect 10784 17280 10836 17332
rect 11428 17280 11480 17332
rect 13084 17323 13136 17332
rect 13084 17289 13093 17323
rect 13093 17289 13127 17323
rect 13127 17289 13136 17323
rect 13084 17280 13136 17289
rect 13820 17323 13872 17332
rect 13820 17289 13829 17323
rect 13829 17289 13863 17323
rect 13863 17289 13872 17323
rect 13820 17280 13872 17289
rect 14464 17323 14516 17332
rect 14464 17289 14473 17323
rect 14473 17289 14507 17323
rect 14507 17289 14516 17323
rect 14464 17280 14516 17289
rect 14740 17280 14792 17332
rect 8760 17212 8812 17264
rect 9128 17187 9180 17196
rect 9128 17153 9137 17187
rect 9137 17153 9171 17187
rect 9171 17153 9180 17187
rect 9128 17144 9180 17153
rect 9404 17187 9456 17196
rect 9404 17153 9443 17187
rect 9443 17153 9456 17187
rect 9404 17144 9456 17153
rect 9864 17212 9916 17264
rect 10324 17212 10376 17264
rect 5724 17076 5776 17128
rect 8668 17076 8720 17128
rect 9680 17076 9732 17128
rect 10692 17076 10744 17128
rect 12256 17144 12308 17196
rect 12900 17144 12952 17196
rect 13268 17187 13320 17196
rect 13268 17153 13277 17187
rect 13277 17153 13311 17187
rect 13311 17153 13320 17187
rect 13268 17144 13320 17153
rect 13912 17144 13964 17196
rect 15292 17212 15344 17264
rect 14096 17187 14148 17196
rect 14096 17153 14105 17187
rect 14105 17153 14139 17187
rect 14139 17153 14148 17187
rect 14096 17144 14148 17153
rect 14556 17144 14608 17196
rect 11612 17076 11664 17128
rect 12348 17076 12400 17128
rect 14832 17187 14884 17196
rect 14832 17153 14841 17187
rect 14841 17153 14875 17187
rect 14875 17153 14884 17187
rect 14832 17144 14884 17153
rect 15016 17187 15068 17196
rect 15016 17153 15025 17187
rect 15025 17153 15059 17187
rect 15059 17153 15068 17187
rect 15016 17144 15068 17153
rect 15384 17144 15436 17196
rect 15752 17187 15804 17196
rect 15752 17153 15761 17187
rect 15761 17153 15795 17187
rect 15795 17153 15804 17187
rect 15752 17144 15804 17153
rect 14740 17076 14792 17128
rect 15568 17076 15620 17128
rect 16396 17076 16448 17128
rect 11152 17008 11204 17060
rect 11796 17008 11848 17060
rect 15016 17008 15068 17060
rect 15200 17051 15252 17060
rect 15200 17017 15209 17051
rect 15209 17017 15243 17051
rect 15243 17017 15252 17051
rect 15200 17008 15252 17017
rect 3792 16940 3844 16992
rect 4068 16940 4120 16992
rect 5264 16940 5316 16992
rect 5540 16983 5592 16992
rect 5540 16949 5549 16983
rect 5549 16949 5583 16983
rect 5583 16949 5592 16983
rect 5540 16940 5592 16949
rect 5816 16940 5868 16992
rect 7104 16940 7156 16992
rect 12624 16940 12676 16992
rect 14280 16940 14332 16992
rect 15476 16940 15528 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 2320 16736 2372 16788
rect 3700 16736 3752 16788
rect 5264 16736 5316 16788
rect 5908 16736 5960 16788
rect 8944 16736 8996 16788
rect 9312 16736 9364 16788
rect 9772 16779 9824 16788
rect 9772 16745 9781 16779
rect 9781 16745 9815 16779
rect 9815 16745 9824 16779
rect 9772 16736 9824 16745
rect 10876 16736 10928 16788
rect 12992 16736 13044 16788
rect 15384 16736 15436 16788
rect 1400 16643 1452 16652
rect 1400 16609 1409 16643
rect 1409 16609 1443 16643
rect 1443 16609 1452 16643
rect 1400 16600 1452 16609
rect 1492 16532 1544 16584
rect 3792 16575 3844 16584
rect 3792 16541 3801 16575
rect 3801 16541 3835 16575
rect 3835 16541 3844 16575
rect 3792 16532 3844 16541
rect 4068 16575 4120 16584
rect 4068 16541 4077 16575
rect 4077 16541 4111 16575
rect 4111 16541 4120 16575
rect 4068 16532 4120 16541
rect 2872 16464 2924 16516
rect 3976 16507 4028 16516
rect 3976 16473 3985 16507
rect 3985 16473 4019 16507
rect 4019 16473 4028 16507
rect 3976 16464 4028 16473
rect 4252 16532 4304 16584
rect 4712 16600 4764 16652
rect 5080 16600 5132 16652
rect 5264 16643 5316 16652
rect 5264 16609 5273 16643
rect 5273 16609 5307 16643
rect 5307 16609 5316 16643
rect 5264 16600 5316 16609
rect 4620 16532 4672 16584
rect 5540 16575 5592 16584
rect 5540 16541 5574 16575
rect 5574 16541 5592 16575
rect 4712 16464 4764 16516
rect 3056 16396 3108 16448
rect 3332 16439 3384 16448
rect 3332 16405 3341 16439
rect 3341 16405 3375 16439
rect 3375 16405 3384 16439
rect 3332 16396 3384 16405
rect 3516 16396 3568 16448
rect 4160 16396 4212 16448
rect 4528 16439 4580 16448
rect 4528 16405 4537 16439
rect 4537 16405 4571 16439
rect 4571 16405 4580 16439
rect 4528 16396 4580 16405
rect 5540 16532 5592 16541
rect 8116 16575 8168 16584
rect 8116 16541 8125 16575
rect 8125 16541 8159 16575
rect 8159 16541 8168 16575
rect 8116 16532 8168 16541
rect 9404 16532 9456 16584
rect 9772 16600 9824 16652
rect 10508 16668 10560 16720
rect 11704 16668 11756 16720
rect 10140 16600 10192 16652
rect 6000 16464 6052 16516
rect 9036 16464 9088 16516
rect 9956 16532 10008 16584
rect 10416 16575 10468 16584
rect 10416 16541 10425 16575
rect 10425 16541 10459 16575
rect 10459 16541 10468 16575
rect 10416 16532 10468 16541
rect 11336 16600 11388 16652
rect 6276 16396 6328 16448
rect 9312 16396 9364 16448
rect 9496 16396 9548 16448
rect 10048 16464 10100 16516
rect 10784 16532 10836 16584
rect 12440 16532 12492 16584
rect 13084 16532 13136 16584
rect 13820 16668 13872 16720
rect 15476 16600 15528 16652
rect 13268 16575 13320 16584
rect 13268 16541 13277 16575
rect 13277 16541 13311 16575
rect 13311 16541 13320 16575
rect 13268 16532 13320 16541
rect 13452 16575 13504 16584
rect 13452 16541 13461 16575
rect 13461 16541 13495 16575
rect 13495 16541 13504 16575
rect 13452 16532 13504 16541
rect 9956 16439 10008 16448
rect 9956 16405 9965 16439
rect 9965 16405 9999 16439
rect 9999 16405 10008 16439
rect 9956 16396 10008 16405
rect 10416 16396 10468 16448
rect 10600 16396 10652 16448
rect 11152 16507 11204 16516
rect 11152 16473 11161 16507
rect 11161 16473 11195 16507
rect 11195 16473 11204 16507
rect 11152 16464 11204 16473
rect 14004 16532 14056 16584
rect 14740 16532 14792 16584
rect 16028 16575 16080 16584
rect 16028 16541 16037 16575
rect 16037 16541 16071 16575
rect 16071 16541 16080 16575
rect 16028 16532 16080 16541
rect 13728 16464 13780 16516
rect 14556 16464 14608 16516
rect 14832 16464 14884 16516
rect 15108 16464 15160 16516
rect 15752 16464 15804 16516
rect 16304 16532 16356 16584
rect 11888 16396 11940 16448
rect 12532 16396 12584 16448
rect 12900 16396 12952 16448
rect 13360 16396 13412 16448
rect 14004 16396 14056 16448
rect 15016 16396 15068 16448
rect 15568 16439 15620 16448
rect 15568 16405 15577 16439
rect 15577 16405 15611 16439
rect 15611 16405 15620 16439
rect 15568 16396 15620 16405
rect 4874 16294 4926 16346
rect 4938 16294 4990 16346
rect 5002 16294 5054 16346
rect 5066 16294 5118 16346
rect 5130 16294 5182 16346
rect 2964 16192 3016 16244
rect 3516 16235 3568 16244
rect 3516 16201 3525 16235
rect 3525 16201 3559 16235
rect 3559 16201 3568 16235
rect 3516 16192 3568 16201
rect 3976 16235 4028 16244
rect 3976 16201 3985 16235
rect 3985 16201 4019 16235
rect 4019 16201 4028 16235
rect 3976 16192 4028 16201
rect 4620 16192 4672 16244
rect 3332 16124 3384 16176
rect 5908 16192 5960 16244
rect 6000 16235 6052 16244
rect 6000 16201 6009 16235
rect 6009 16201 6043 16235
rect 6043 16201 6052 16235
rect 6000 16192 6052 16201
rect 9036 16192 9088 16244
rect 9404 16235 9456 16244
rect 9404 16201 9413 16235
rect 9413 16201 9447 16235
rect 9447 16201 9456 16235
rect 9404 16192 9456 16201
rect 9588 16192 9640 16244
rect 9772 16192 9824 16244
rect 11060 16192 11112 16244
rect 11520 16235 11572 16244
rect 11520 16201 11529 16235
rect 11529 16201 11563 16235
rect 11563 16201 11572 16235
rect 11520 16192 11572 16201
rect 15292 16192 15344 16244
rect 1400 16099 1452 16108
rect 1400 16065 1409 16099
rect 1409 16065 1443 16099
rect 1443 16065 1452 16099
rect 1400 16056 1452 16065
rect 1676 16099 1728 16108
rect 1676 16065 1710 16099
rect 1710 16065 1728 16099
rect 1676 16056 1728 16065
rect 2044 16056 2096 16108
rect 3148 16056 3200 16108
rect 3608 16056 3660 16108
rect 4068 16056 4120 16108
rect 4252 16099 4304 16108
rect 4252 16065 4260 16099
rect 4260 16065 4294 16099
rect 4294 16065 4304 16099
rect 4252 16056 4304 16065
rect 4344 16099 4396 16108
rect 4344 16065 4353 16099
rect 4353 16065 4387 16099
rect 4387 16065 4396 16099
rect 4344 16056 4396 16065
rect 5080 16124 5132 16176
rect 5632 16124 5684 16176
rect 5724 16124 5776 16176
rect 6460 16124 6512 16176
rect 4712 16056 4764 16108
rect 3976 15988 4028 16040
rect 2780 15963 2832 15972
rect 2780 15929 2789 15963
rect 2789 15929 2823 15963
rect 2823 15929 2832 15963
rect 2780 15920 2832 15929
rect 3608 15920 3660 15972
rect 4344 15920 4396 15972
rect 2964 15852 3016 15904
rect 4988 15920 5040 15972
rect 7380 16056 7432 16108
rect 8760 16099 8812 16108
rect 8760 16065 8769 16099
rect 8769 16065 8803 16099
rect 8803 16065 8812 16099
rect 8760 16056 8812 16065
rect 8944 16099 8996 16108
rect 8944 16065 8953 16099
rect 8953 16065 8987 16099
rect 8987 16065 8996 16099
rect 8944 16056 8996 16065
rect 9128 16056 9180 16108
rect 9588 16099 9640 16108
rect 9588 16065 9597 16099
rect 9597 16065 9631 16099
rect 9631 16065 9640 16099
rect 9588 16056 9640 16065
rect 9680 16099 9732 16108
rect 9680 16065 9689 16099
rect 9689 16065 9723 16099
rect 9723 16065 9732 16099
rect 9680 16056 9732 16065
rect 10140 16124 10192 16176
rect 5540 15920 5592 15972
rect 5724 15920 5776 15972
rect 4528 15852 4580 15904
rect 4896 15852 4948 15904
rect 5632 15852 5684 15904
rect 5816 15895 5868 15904
rect 5816 15861 5825 15895
rect 5825 15861 5859 15895
rect 5859 15861 5868 15895
rect 5816 15852 5868 15861
rect 10692 16056 10744 16108
rect 11428 16124 11480 16176
rect 11888 16167 11940 16176
rect 11888 16133 11897 16167
rect 11897 16133 11931 16167
rect 11931 16133 11940 16167
rect 11888 16124 11940 16133
rect 12256 16099 12308 16108
rect 12256 16065 12265 16099
rect 12265 16065 12299 16099
rect 12299 16065 12308 16099
rect 12256 16056 12308 16065
rect 9956 15988 10008 16040
rect 10140 15988 10192 16040
rect 10600 16031 10652 16040
rect 10600 15997 10609 16031
rect 10609 15997 10643 16031
rect 10643 15997 10652 16031
rect 10600 15988 10652 15997
rect 10876 15988 10928 16040
rect 11520 15988 11572 16040
rect 7196 15895 7248 15904
rect 7196 15861 7205 15895
rect 7205 15861 7239 15895
rect 7239 15861 7248 15895
rect 7196 15852 7248 15861
rect 8944 15895 8996 15904
rect 8944 15861 8953 15895
rect 8953 15861 8987 15895
rect 8987 15861 8996 15895
rect 8944 15852 8996 15861
rect 9956 15852 10008 15904
rect 10048 15895 10100 15904
rect 10048 15861 10057 15895
rect 10057 15861 10091 15895
rect 10091 15861 10100 15895
rect 10048 15852 10100 15861
rect 10324 15895 10376 15904
rect 10324 15861 10333 15895
rect 10333 15861 10367 15895
rect 10367 15861 10376 15895
rect 10324 15852 10376 15861
rect 11336 15920 11388 15972
rect 12532 15988 12584 16040
rect 13268 16056 13320 16108
rect 13452 16124 13504 16176
rect 14096 16124 14148 16176
rect 13452 15988 13504 16040
rect 13912 16056 13964 16108
rect 14648 16099 14700 16108
rect 14648 16065 14657 16099
rect 14657 16065 14691 16099
rect 14691 16065 14700 16099
rect 14648 16056 14700 16065
rect 14924 16124 14976 16176
rect 15568 16124 15620 16176
rect 15660 16056 15712 16108
rect 10784 15852 10836 15904
rect 11704 15895 11756 15904
rect 11704 15861 11713 15895
rect 11713 15861 11747 15895
rect 11747 15861 11756 15895
rect 11704 15852 11756 15861
rect 13176 15895 13228 15904
rect 13176 15861 13185 15895
rect 13185 15861 13219 15895
rect 13219 15861 13228 15895
rect 13176 15852 13228 15861
rect 14096 15920 14148 15972
rect 14556 15920 14608 15972
rect 15844 15852 15896 15904
rect 16028 15852 16080 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 1676 15648 1728 15700
rect 1768 15691 1820 15700
rect 1768 15657 1777 15691
rect 1777 15657 1811 15691
rect 1811 15657 1820 15691
rect 1768 15648 1820 15657
rect 2688 15648 2740 15700
rect 3884 15648 3936 15700
rect 4620 15648 4672 15700
rect 4804 15648 4856 15700
rect 5356 15648 5408 15700
rect 5632 15648 5684 15700
rect 6276 15648 6328 15700
rect 6920 15648 6972 15700
rect 7380 15648 7432 15700
rect 8208 15648 8260 15700
rect 8576 15648 8628 15700
rect 2780 15512 2832 15564
rect 3056 15623 3108 15632
rect 3056 15589 3065 15623
rect 3065 15589 3099 15623
rect 3099 15589 3108 15623
rect 3056 15580 3108 15589
rect 3608 15580 3660 15632
rect 3332 15512 3384 15564
rect 1952 15376 2004 15428
rect 2872 15444 2924 15496
rect 3424 15444 3476 15496
rect 3884 15444 3936 15496
rect 4804 15555 4856 15564
rect 4804 15521 4813 15555
rect 4813 15521 4847 15555
rect 4847 15521 4856 15555
rect 4804 15512 4856 15521
rect 4068 15487 4120 15496
rect 4068 15453 4077 15487
rect 4077 15453 4111 15487
rect 4111 15453 4120 15487
rect 4068 15444 4120 15453
rect 3700 15376 3752 15428
rect 4896 15487 4948 15496
rect 4896 15453 4905 15487
rect 4905 15453 4939 15487
rect 4939 15453 4948 15487
rect 4896 15444 4948 15453
rect 4988 15487 5040 15496
rect 4988 15453 4997 15487
rect 4997 15453 5031 15487
rect 5031 15453 5040 15487
rect 4988 15444 5040 15453
rect 5172 15487 5224 15496
rect 5172 15453 5181 15487
rect 5181 15453 5215 15487
rect 5215 15453 5224 15487
rect 5172 15444 5224 15453
rect 5448 15512 5500 15564
rect 5632 15487 5684 15496
rect 5632 15453 5641 15487
rect 5641 15453 5675 15487
rect 5675 15453 5684 15487
rect 5632 15444 5684 15453
rect 5908 15487 5960 15496
rect 5908 15453 5917 15487
rect 5917 15453 5951 15487
rect 5951 15453 5960 15487
rect 5908 15444 5960 15453
rect 6276 15487 6328 15496
rect 6276 15453 6285 15487
rect 6285 15453 6319 15487
rect 6319 15453 6328 15487
rect 6276 15444 6328 15453
rect 8116 15512 8168 15564
rect 7196 15444 7248 15496
rect 8392 15444 8444 15496
rect 9680 15648 9732 15700
rect 9772 15691 9824 15700
rect 9772 15657 9781 15691
rect 9781 15657 9815 15691
rect 9815 15657 9824 15691
rect 9772 15648 9824 15657
rect 9956 15648 10008 15700
rect 10508 15648 10560 15700
rect 10600 15580 10652 15632
rect 10876 15580 10928 15632
rect 8852 15512 8904 15564
rect 10784 15512 10836 15564
rect 9496 15487 9548 15496
rect 9496 15453 9506 15487
rect 9506 15453 9540 15487
rect 9540 15453 9548 15487
rect 9496 15444 9548 15453
rect 5816 15419 5868 15428
rect 5816 15385 5825 15419
rect 5825 15385 5859 15419
rect 5859 15385 5868 15419
rect 5816 15376 5868 15385
rect 6184 15419 6236 15428
rect 6184 15385 6193 15419
rect 6193 15385 6227 15419
rect 6227 15385 6236 15419
rect 6184 15376 6236 15385
rect 9772 15444 9824 15496
rect 9956 15487 10008 15496
rect 9956 15453 9965 15487
rect 9965 15453 9999 15487
rect 9999 15453 10008 15487
rect 9956 15444 10008 15453
rect 10140 15444 10192 15496
rect 10324 15444 10376 15496
rect 10416 15487 10468 15496
rect 10416 15453 10425 15487
rect 10425 15453 10459 15487
rect 10459 15453 10468 15487
rect 10416 15444 10468 15453
rect 10508 15487 10560 15496
rect 10508 15453 10517 15487
rect 10517 15453 10551 15487
rect 10551 15453 10560 15487
rect 10508 15444 10560 15453
rect 10600 15487 10652 15496
rect 10600 15453 10609 15487
rect 10609 15453 10643 15487
rect 10643 15453 10652 15487
rect 10600 15444 10652 15453
rect 10968 15444 11020 15496
rect 11704 15580 11756 15632
rect 11888 15512 11940 15564
rect 3148 15308 3200 15360
rect 3884 15308 3936 15360
rect 3976 15308 4028 15360
rect 6368 15308 6420 15360
rect 6552 15351 6604 15360
rect 6552 15317 6561 15351
rect 6561 15317 6595 15351
rect 6595 15317 6604 15351
rect 6552 15308 6604 15317
rect 8300 15351 8352 15360
rect 8300 15317 8309 15351
rect 8309 15317 8343 15351
rect 8343 15317 8352 15351
rect 8300 15308 8352 15317
rect 9312 15351 9364 15360
rect 9312 15317 9321 15351
rect 9321 15317 9355 15351
rect 9355 15317 9364 15351
rect 9312 15308 9364 15317
rect 9772 15308 9824 15360
rect 10324 15308 10376 15360
rect 10968 15308 11020 15360
rect 11336 15308 11388 15360
rect 11796 15444 11848 15496
rect 14004 15648 14056 15700
rect 14648 15648 14700 15700
rect 14832 15648 14884 15700
rect 13728 15580 13780 15632
rect 15016 15512 15068 15564
rect 12348 15487 12400 15496
rect 12348 15453 12357 15487
rect 12357 15453 12391 15487
rect 12391 15453 12400 15487
rect 12348 15444 12400 15453
rect 12532 15444 12584 15496
rect 11612 15376 11664 15428
rect 12900 15376 12952 15428
rect 13268 15419 13320 15428
rect 13268 15385 13277 15419
rect 13277 15385 13311 15419
rect 13311 15385 13320 15419
rect 13268 15376 13320 15385
rect 13360 15376 13412 15428
rect 14188 15444 14240 15496
rect 14924 15487 14976 15496
rect 14924 15453 14933 15487
rect 14933 15453 14967 15487
rect 14967 15453 14976 15487
rect 14924 15444 14976 15453
rect 15292 15487 15344 15496
rect 15292 15453 15301 15487
rect 15301 15453 15335 15487
rect 15335 15453 15344 15487
rect 15292 15444 15344 15453
rect 15568 15487 15620 15496
rect 15568 15453 15577 15487
rect 15577 15453 15611 15487
rect 15611 15453 15620 15487
rect 15568 15444 15620 15453
rect 16028 15487 16080 15496
rect 16028 15453 16037 15487
rect 16037 15453 16071 15487
rect 16071 15453 16080 15487
rect 16028 15444 16080 15453
rect 16120 15487 16172 15496
rect 16120 15453 16129 15487
rect 16129 15453 16163 15487
rect 16163 15453 16172 15487
rect 16120 15444 16172 15453
rect 16396 15444 16448 15496
rect 11520 15308 11572 15360
rect 12072 15308 12124 15360
rect 12532 15351 12584 15360
rect 12532 15317 12541 15351
rect 12541 15317 12575 15351
rect 12575 15317 12584 15351
rect 12532 15308 12584 15317
rect 12624 15308 12676 15360
rect 12992 15308 13044 15360
rect 13820 15308 13872 15360
rect 14372 15308 14424 15360
rect 14648 15308 14700 15360
rect 4874 15206 4926 15258
rect 4938 15206 4990 15258
rect 5002 15206 5054 15258
rect 5066 15206 5118 15258
rect 5130 15206 5182 15258
rect 1584 15104 1636 15156
rect 2412 15104 2464 15156
rect 3700 15104 3752 15156
rect 4896 15104 4948 15156
rect 5724 15147 5776 15156
rect 5724 15113 5733 15147
rect 5733 15113 5767 15147
rect 5767 15113 5776 15147
rect 5724 15104 5776 15113
rect 6184 15147 6236 15156
rect 6184 15113 6193 15147
rect 6193 15113 6227 15147
rect 6227 15113 6236 15147
rect 6184 15104 6236 15113
rect 5448 15036 5500 15088
rect 6920 15104 6972 15156
rect 8300 15104 8352 15156
rect 9864 15104 9916 15156
rect 2044 14968 2096 15020
rect 2136 15011 2188 15020
rect 2136 14977 2145 15011
rect 2145 14977 2179 15011
rect 2179 14977 2188 15011
rect 2136 14968 2188 14977
rect 2504 15011 2556 15020
rect 2504 14977 2513 15011
rect 2513 14977 2547 15011
rect 2547 14977 2556 15011
rect 2504 14968 2556 14977
rect 4712 14968 4764 15020
rect 5172 14968 5224 15020
rect 5540 15011 5592 15020
rect 5540 14977 5549 15011
rect 5549 14977 5583 15011
rect 5583 14977 5592 15011
rect 5540 14968 5592 14977
rect 6000 15011 6052 15020
rect 6000 14977 6009 15011
rect 6009 14977 6043 15011
rect 6043 14977 6052 15011
rect 6000 14968 6052 14977
rect 8944 15036 8996 15088
rect 10692 15104 10744 15156
rect 10784 15104 10836 15156
rect 10876 15104 10928 15156
rect 11060 15104 11112 15156
rect 11796 15104 11848 15156
rect 6368 14900 6420 14952
rect 8116 14968 8168 15020
rect 10508 15036 10560 15088
rect 9220 14900 9272 14952
rect 10600 15011 10652 15020
rect 10600 14977 10609 15011
rect 10609 14977 10643 15011
rect 10643 14977 10652 15011
rect 10600 14968 10652 14977
rect 10784 14968 10836 15020
rect 9864 14832 9916 14884
rect 10140 14832 10192 14884
rect 10416 14832 10468 14884
rect 10876 14832 10928 14884
rect 11060 15011 11112 15020
rect 11060 14977 11069 15011
rect 11069 14977 11103 15011
rect 11103 14977 11112 15011
rect 11060 14968 11112 14977
rect 11428 15036 11480 15088
rect 11704 15011 11756 15020
rect 11704 14977 11713 15011
rect 11713 14977 11747 15011
rect 11747 14977 11756 15011
rect 11704 14968 11756 14977
rect 11796 15011 11848 15020
rect 11796 14977 11805 15011
rect 11805 14977 11839 15011
rect 11839 14977 11848 15011
rect 11796 14968 11848 14977
rect 11612 14900 11664 14952
rect 12348 14968 12400 15020
rect 14096 14968 14148 15020
rect 14464 14968 14516 15020
rect 12072 14900 12124 14952
rect 12440 14832 12492 14884
rect 13268 14900 13320 14952
rect 13820 14943 13872 14952
rect 13820 14909 13829 14943
rect 13829 14909 13863 14943
rect 13863 14909 13872 14943
rect 13820 14900 13872 14909
rect 14740 15011 14792 15020
rect 14740 14977 14749 15011
rect 14749 14977 14783 15011
rect 14783 14977 14792 15011
rect 14740 14968 14792 14977
rect 15016 15011 15068 15020
rect 15016 14977 15025 15011
rect 15025 14977 15059 15011
rect 15059 14977 15068 15011
rect 15016 14968 15068 14977
rect 15384 15011 15436 15020
rect 15384 14977 15393 15011
rect 15393 14977 15427 15011
rect 15427 14977 15436 15011
rect 15384 14968 15436 14977
rect 16212 15079 16264 15088
rect 16212 15045 16221 15079
rect 16221 15045 16255 15079
rect 16255 15045 16264 15079
rect 16212 15036 16264 15045
rect 15660 14968 15712 15020
rect 15936 14968 15988 15020
rect 16028 15011 16080 15020
rect 16028 14977 16037 15011
rect 16037 14977 16071 15011
rect 16071 14977 16080 15011
rect 16028 14968 16080 14977
rect 14832 14832 14884 14884
rect 15016 14832 15068 14884
rect 15936 14832 15988 14884
rect 4712 14764 4764 14816
rect 9496 14764 9548 14816
rect 10600 14764 10652 14816
rect 12164 14807 12216 14816
rect 12164 14773 12173 14807
rect 12173 14773 12207 14807
rect 12207 14773 12216 14807
rect 12164 14764 12216 14773
rect 12348 14764 12400 14816
rect 13728 14764 13780 14816
rect 14740 14764 14792 14816
rect 15108 14807 15160 14816
rect 15108 14773 15117 14807
rect 15117 14773 15151 14807
rect 15151 14773 15160 14807
rect 15108 14764 15160 14773
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 5632 14603 5684 14612
rect 5632 14569 5641 14603
rect 5641 14569 5675 14603
rect 5675 14569 5684 14603
rect 5632 14560 5684 14569
rect 10508 14560 10560 14612
rect 6276 14492 6328 14544
rect 8760 14535 8812 14544
rect 8760 14501 8769 14535
rect 8769 14501 8803 14535
rect 8803 14501 8812 14535
rect 8760 14492 8812 14501
rect 9036 14492 9088 14544
rect 9496 14492 9548 14544
rect 4068 14424 4120 14476
rect 4896 14424 4948 14476
rect 3332 14399 3384 14408
rect 3332 14365 3341 14399
rect 3341 14365 3375 14399
rect 3375 14365 3384 14399
rect 3332 14356 3384 14365
rect 4344 14356 4396 14408
rect 4620 14356 4672 14408
rect 5264 14356 5316 14408
rect 5448 14399 5500 14408
rect 5448 14365 5457 14399
rect 5457 14365 5491 14399
rect 5491 14365 5500 14399
rect 5448 14356 5500 14365
rect 6092 14356 6144 14408
rect 6184 14399 6236 14408
rect 6184 14365 6193 14399
rect 6193 14365 6227 14399
rect 6227 14365 6236 14399
rect 6184 14356 6236 14365
rect 6368 14356 6420 14408
rect 6920 14424 6972 14476
rect 7196 14424 7248 14476
rect 9220 14424 9272 14476
rect 9680 14492 9732 14544
rect 10600 14535 10652 14544
rect 10600 14501 10609 14535
rect 10609 14501 10643 14535
rect 10643 14501 10652 14535
rect 10600 14492 10652 14501
rect 10784 14560 10836 14612
rect 9956 14424 10008 14476
rect 11060 14424 11112 14476
rect 4804 14288 4856 14340
rect 8024 14356 8076 14408
rect 7288 14288 7340 14340
rect 8300 14399 8352 14408
rect 8300 14365 8309 14399
rect 8309 14365 8343 14399
rect 8343 14365 8352 14399
rect 8300 14356 8352 14365
rect 8576 14399 8628 14408
rect 8576 14365 8585 14399
rect 8585 14365 8619 14399
rect 8619 14365 8628 14399
rect 8576 14356 8628 14365
rect 8944 14356 8996 14408
rect 15200 14560 15252 14612
rect 8392 14288 8444 14340
rect 11336 14492 11388 14544
rect 14004 14492 14056 14544
rect 15660 14560 15712 14612
rect 16120 14492 16172 14544
rect 11704 14424 11756 14476
rect 13360 14424 13412 14476
rect 11428 14399 11480 14408
rect 11428 14365 11437 14399
rect 11437 14365 11471 14399
rect 11471 14365 11480 14399
rect 11428 14356 11480 14365
rect 11612 14356 11664 14408
rect 11888 14356 11940 14408
rect 3424 14263 3476 14272
rect 3424 14229 3433 14263
rect 3433 14229 3467 14263
rect 3467 14229 3476 14263
rect 3424 14220 3476 14229
rect 4252 14220 4304 14272
rect 4620 14220 4672 14272
rect 5172 14220 5224 14272
rect 5540 14220 5592 14272
rect 5632 14220 5684 14272
rect 6000 14220 6052 14272
rect 6920 14263 6972 14272
rect 6920 14229 6929 14263
rect 6929 14229 6963 14263
rect 6963 14229 6972 14263
rect 6920 14220 6972 14229
rect 8300 14220 8352 14272
rect 10692 14220 10744 14272
rect 11060 14220 11112 14272
rect 12164 14288 12216 14340
rect 12900 14288 12952 14340
rect 12808 14220 12860 14272
rect 13268 14220 13320 14272
rect 13360 14220 13412 14272
rect 13912 14424 13964 14476
rect 14556 14356 14608 14408
rect 14740 14399 14792 14408
rect 14740 14365 14774 14399
rect 14774 14365 14792 14399
rect 14740 14356 14792 14365
rect 15660 14356 15712 14408
rect 15292 14288 15344 14340
rect 16212 14288 16264 14340
rect 13820 14263 13872 14272
rect 13820 14229 13829 14263
rect 13829 14229 13863 14263
rect 13863 14229 13872 14263
rect 13820 14220 13872 14229
rect 14924 14220 14976 14272
rect 16028 14220 16080 14272
rect 4874 14118 4926 14170
rect 4938 14118 4990 14170
rect 5002 14118 5054 14170
rect 5066 14118 5118 14170
rect 5130 14118 5182 14170
rect 2872 14016 2924 14068
rect 3148 14016 3200 14068
rect 3792 13948 3844 14000
rect 2044 13923 2096 13932
rect 2044 13889 2053 13923
rect 2053 13889 2087 13923
rect 2087 13889 2096 13923
rect 2044 13880 2096 13889
rect 2412 13812 2464 13864
rect 3608 13923 3660 13932
rect 3608 13889 3617 13923
rect 3617 13889 3651 13923
rect 3651 13889 3660 13923
rect 3608 13880 3660 13889
rect 4252 13880 4304 13932
rect 5172 14016 5224 14068
rect 5448 14016 5500 14068
rect 7104 14016 7156 14068
rect 9128 14016 9180 14068
rect 10508 14016 10560 14068
rect 11060 14016 11112 14068
rect 12808 14059 12860 14068
rect 12808 14025 12817 14059
rect 12817 14025 12851 14059
rect 12851 14025 12860 14059
rect 12808 14016 12860 14025
rect 14188 14059 14240 14068
rect 14188 14025 14197 14059
rect 14197 14025 14231 14059
rect 14231 14025 14240 14059
rect 14188 14016 14240 14025
rect 15200 14016 15252 14068
rect 16212 14059 16264 14068
rect 16212 14025 16221 14059
rect 16221 14025 16255 14059
rect 16255 14025 16264 14059
rect 16212 14016 16264 14025
rect 4436 13880 4488 13932
rect 4068 13812 4120 13864
rect 5172 13880 5224 13932
rect 5724 13923 5776 13932
rect 5724 13889 5742 13923
rect 5742 13889 5776 13923
rect 5724 13880 5776 13889
rect 6828 13880 6880 13932
rect 6920 13923 6972 13932
rect 6920 13889 6929 13923
rect 6929 13889 6963 13923
rect 6963 13889 6972 13923
rect 6920 13880 6972 13889
rect 7012 13923 7064 13932
rect 7012 13889 7021 13923
rect 7021 13889 7055 13923
rect 7055 13889 7064 13923
rect 7012 13880 7064 13889
rect 8116 13948 8168 14000
rect 10232 13948 10284 14000
rect 13268 13948 13320 14000
rect 8024 13923 8076 13932
rect 8024 13889 8033 13923
rect 8033 13889 8067 13923
rect 8067 13889 8076 13923
rect 8024 13880 8076 13889
rect 8300 13923 8352 13932
rect 8300 13889 8334 13923
rect 8334 13889 8352 13923
rect 8300 13880 8352 13889
rect 9496 13880 9548 13932
rect 10140 13923 10192 13932
rect 10140 13889 10149 13923
rect 10149 13889 10183 13923
rect 10183 13889 10192 13923
rect 10140 13880 10192 13889
rect 10600 13923 10652 13932
rect 10600 13889 10609 13923
rect 10609 13889 10643 13923
rect 10643 13889 10652 13923
rect 10600 13880 10652 13889
rect 3608 13744 3660 13796
rect 4344 13744 4396 13796
rect 4896 13744 4948 13796
rect 6644 13787 6696 13796
rect 6644 13753 6653 13787
rect 6653 13753 6687 13787
rect 6687 13753 6696 13787
rect 6644 13744 6696 13753
rect 10508 13812 10560 13864
rect 11244 13880 11296 13932
rect 12072 13880 12124 13932
rect 13912 13923 13964 13932
rect 13912 13889 13921 13923
rect 13921 13889 13955 13923
rect 13955 13889 13964 13923
rect 13912 13880 13964 13889
rect 15108 13948 15160 14000
rect 10784 13812 10836 13864
rect 12440 13812 12492 13864
rect 13820 13855 13872 13864
rect 13820 13821 13829 13855
rect 13829 13821 13863 13855
rect 13863 13821 13872 13855
rect 13820 13812 13872 13821
rect 16028 13923 16080 13932
rect 16028 13889 16037 13923
rect 16037 13889 16071 13923
rect 16071 13889 16080 13923
rect 16028 13880 16080 13889
rect 14372 13812 14424 13864
rect 14556 13855 14608 13864
rect 14556 13821 14565 13855
rect 14565 13821 14599 13855
rect 14599 13821 14608 13855
rect 14556 13812 14608 13821
rect 14004 13744 14056 13796
rect 1952 13719 2004 13728
rect 1952 13685 1961 13719
rect 1961 13685 1995 13719
rect 1995 13685 2004 13719
rect 1952 13676 2004 13685
rect 3700 13676 3752 13728
rect 3976 13676 4028 13728
rect 4068 13719 4120 13728
rect 4068 13685 4077 13719
rect 4077 13685 4111 13719
rect 4111 13685 4120 13719
rect 4068 13676 4120 13685
rect 4436 13676 4488 13728
rect 5356 13676 5408 13728
rect 5816 13676 5868 13728
rect 12164 13719 12216 13728
rect 12164 13685 12173 13719
rect 12173 13685 12207 13719
rect 12207 13685 12216 13719
rect 12164 13676 12216 13685
rect 12256 13676 12308 13728
rect 15660 13676 15712 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 4804 13472 4856 13524
rect 5264 13472 5316 13524
rect 7196 13515 7248 13524
rect 7196 13481 7205 13515
rect 7205 13481 7239 13515
rect 7239 13481 7248 13515
rect 7196 13472 7248 13481
rect 12992 13472 13044 13524
rect 13912 13472 13964 13524
rect 15108 13472 15160 13524
rect 2412 13404 2464 13456
rect 3148 13404 3200 13456
rect 2872 13268 2924 13320
rect 3056 13268 3108 13320
rect 3608 13311 3660 13320
rect 3608 13277 3617 13311
rect 3617 13277 3651 13311
rect 3651 13277 3660 13311
rect 3608 13268 3660 13277
rect 4252 13404 4304 13456
rect 4896 13336 4948 13388
rect 5264 13336 5316 13388
rect 6000 13336 6052 13388
rect 7288 13404 7340 13456
rect 1676 13243 1728 13252
rect 1676 13209 1710 13243
rect 1710 13209 1728 13243
rect 1676 13200 1728 13209
rect 3240 13243 3292 13252
rect 3240 13209 3249 13243
rect 3249 13209 3283 13243
rect 3283 13209 3292 13243
rect 3240 13200 3292 13209
rect 3424 13200 3476 13252
rect 2872 13132 2924 13184
rect 3516 13132 3568 13184
rect 4252 13311 4304 13320
rect 4252 13277 4261 13311
rect 4261 13277 4295 13311
rect 4295 13277 4304 13311
rect 4252 13268 4304 13277
rect 7012 13268 7064 13320
rect 7288 13311 7340 13320
rect 7288 13277 7297 13311
rect 7297 13277 7331 13311
rect 7331 13277 7340 13311
rect 7288 13268 7340 13277
rect 7472 13268 7524 13320
rect 8208 13268 8260 13320
rect 8300 13268 8352 13320
rect 9680 13268 9732 13320
rect 9864 13311 9916 13320
rect 9864 13277 9873 13311
rect 9873 13277 9907 13311
rect 9907 13277 9916 13311
rect 9864 13268 9916 13277
rect 9956 13268 10008 13320
rect 10600 13268 10652 13320
rect 10692 13311 10744 13320
rect 10692 13277 10701 13311
rect 10701 13277 10735 13311
rect 10735 13277 10744 13311
rect 10692 13268 10744 13277
rect 6828 13243 6880 13252
rect 6828 13209 6837 13243
rect 6837 13209 6871 13243
rect 6871 13209 6880 13243
rect 6828 13200 6880 13209
rect 11520 13404 11572 13456
rect 11060 13336 11112 13388
rect 13820 13404 13872 13456
rect 14188 13404 14240 13456
rect 15384 13515 15436 13524
rect 15384 13481 15393 13515
rect 15393 13481 15427 13515
rect 15427 13481 15436 13515
rect 15384 13472 15436 13481
rect 15568 13515 15620 13524
rect 15568 13481 15577 13515
rect 15577 13481 15611 13515
rect 15611 13481 15620 13515
rect 15568 13472 15620 13481
rect 14372 13336 14424 13388
rect 11980 13311 12032 13320
rect 11980 13277 11989 13311
rect 11989 13277 12023 13311
rect 12023 13277 12032 13311
rect 11980 13268 12032 13277
rect 12256 13311 12308 13320
rect 12256 13277 12290 13311
rect 12290 13277 12308 13311
rect 12256 13268 12308 13277
rect 14096 13268 14148 13320
rect 15292 13336 15344 13388
rect 15200 13311 15252 13320
rect 15200 13277 15209 13311
rect 15209 13277 15243 13311
rect 15243 13277 15252 13311
rect 15200 13268 15252 13277
rect 16120 13311 16172 13320
rect 16120 13277 16129 13311
rect 16129 13277 16163 13311
rect 16163 13277 16172 13311
rect 16120 13268 16172 13277
rect 4160 13132 4212 13184
rect 6552 13132 6604 13184
rect 7380 13132 7432 13184
rect 7748 13132 7800 13184
rect 9772 13132 9824 13184
rect 11796 13132 11848 13184
rect 14740 13200 14792 13252
rect 15292 13200 15344 13252
rect 14096 13175 14148 13184
rect 14096 13141 14105 13175
rect 14105 13141 14139 13175
rect 14139 13141 14148 13175
rect 14096 13132 14148 13141
rect 14648 13132 14700 13184
rect 15752 13132 15804 13184
rect 4874 13030 4926 13082
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 1676 12928 1728 12980
rect 1952 12928 2004 12980
rect 3792 12928 3844 12980
rect 2412 12903 2464 12912
rect 2412 12869 2421 12903
rect 2421 12869 2455 12903
rect 2455 12869 2464 12903
rect 2412 12860 2464 12869
rect 2872 12860 2924 12912
rect 5724 12928 5776 12980
rect 5816 12971 5868 12980
rect 5816 12937 5825 12971
rect 5825 12937 5859 12971
rect 5859 12937 5868 12971
rect 5816 12928 5868 12937
rect 7288 12928 7340 12980
rect 8300 12971 8352 12980
rect 8300 12937 8309 12971
rect 8309 12937 8343 12971
rect 8343 12937 8352 12971
rect 8300 12928 8352 12937
rect 1860 12792 1912 12844
rect 2044 12792 2096 12844
rect 2320 12724 2372 12776
rect 2504 12724 2556 12776
rect 2780 12724 2832 12776
rect 3148 12792 3200 12844
rect 2596 12656 2648 12708
rect 3700 12835 3752 12844
rect 3700 12801 3709 12835
rect 3709 12801 3743 12835
rect 3743 12801 3752 12835
rect 3700 12792 3752 12801
rect 3976 12792 4028 12844
rect 3884 12724 3936 12776
rect 4160 12835 4212 12844
rect 4160 12801 4169 12835
rect 4169 12801 4203 12835
rect 4203 12801 4212 12835
rect 4160 12792 4212 12801
rect 4988 12792 5040 12844
rect 5540 12792 5592 12844
rect 5632 12835 5684 12844
rect 5632 12801 5641 12835
rect 5641 12801 5675 12835
rect 5675 12801 5684 12835
rect 5632 12792 5684 12801
rect 5724 12792 5776 12844
rect 5908 12792 5960 12844
rect 6828 12860 6880 12912
rect 10692 12928 10744 12980
rect 12164 12928 12216 12980
rect 6552 12835 6604 12844
rect 6552 12801 6561 12835
rect 6561 12801 6595 12835
rect 6595 12801 6604 12835
rect 6552 12792 6604 12801
rect 5356 12767 5408 12776
rect 5356 12733 5365 12767
rect 5365 12733 5399 12767
rect 5399 12733 5408 12767
rect 5356 12724 5408 12733
rect 4896 12656 4948 12708
rect 3148 12588 3200 12640
rect 3424 12588 3476 12640
rect 3608 12588 3660 12640
rect 4712 12588 4764 12640
rect 5356 12588 5408 12640
rect 6920 12724 6972 12776
rect 7748 12835 7800 12844
rect 7748 12801 7766 12835
rect 7766 12801 7800 12835
rect 7748 12792 7800 12801
rect 8024 12835 8076 12844
rect 8024 12801 8033 12835
rect 8033 12801 8067 12835
rect 8067 12801 8076 12835
rect 8024 12792 8076 12801
rect 10784 12903 10836 12912
rect 10784 12869 10793 12903
rect 10793 12869 10827 12903
rect 10827 12869 10836 12903
rect 10784 12860 10836 12869
rect 12072 12860 12124 12912
rect 14096 12928 14148 12980
rect 15108 12928 15160 12980
rect 8208 12792 8260 12844
rect 12348 12792 12400 12844
rect 14188 12860 14240 12912
rect 16028 12928 16080 12980
rect 9128 12767 9180 12776
rect 9128 12733 9137 12767
rect 9137 12733 9171 12767
rect 9171 12733 9180 12767
rect 9128 12724 9180 12733
rect 9312 12767 9364 12776
rect 9312 12733 9321 12767
rect 9321 12733 9355 12767
rect 9355 12733 9364 12767
rect 9312 12724 9364 12733
rect 9956 12724 10008 12776
rect 6000 12656 6052 12708
rect 8208 12656 8260 12708
rect 9864 12656 9916 12708
rect 12072 12767 12124 12776
rect 12072 12733 12081 12767
rect 12081 12733 12115 12767
rect 12115 12733 12124 12767
rect 12072 12724 12124 12733
rect 12624 12724 12676 12776
rect 13636 12724 13688 12776
rect 14372 12792 14424 12844
rect 14924 12835 14976 12844
rect 14924 12801 14933 12835
rect 14933 12801 14967 12835
rect 14967 12801 14976 12835
rect 14924 12792 14976 12801
rect 14648 12767 14700 12776
rect 14648 12733 14657 12767
rect 14657 12733 14691 12767
rect 14691 12733 14700 12767
rect 14648 12724 14700 12733
rect 14740 12724 14792 12776
rect 15200 12724 15252 12776
rect 15660 12792 15712 12844
rect 15752 12835 15804 12844
rect 15752 12801 15761 12835
rect 15761 12801 15795 12835
rect 15795 12801 15804 12835
rect 15752 12792 15804 12801
rect 15844 12835 15896 12844
rect 15844 12801 15853 12835
rect 15853 12801 15887 12835
rect 15887 12801 15896 12835
rect 15844 12792 15896 12801
rect 12348 12656 12400 12708
rect 13544 12656 13596 12708
rect 5540 12588 5592 12640
rect 7012 12588 7064 12640
rect 8116 12588 8168 12640
rect 8300 12588 8352 12640
rect 11520 12631 11572 12640
rect 11520 12597 11529 12631
rect 11529 12597 11563 12631
rect 11563 12597 11572 12631
rect 11520 12588 11572 12597
rect 12256 12588 12308 12640
rect 14188 12588 14240 12640
rect 14832 12588 14884 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 3240 12384 3292 12436
rect 3056 12316 3108 12368
rect 5172 12384 5224 12436
rect 5724 12384 5776 12436
rect 6828 12384 6880 12436
rect 2504 12223 2556 12232
rect 1492 12155 1544 12164
rect 1492 12121 1501 12155
rect 1501 12121 1535 12155
rect 1535 12121 1544 12155
rect 2504 12189 2513 12223
rect 2513 12189 2547 12223
rect 2547 12189 2556 12223
rect 2504 12180 2556 12189
rect 2688 12248 2740 12300
rect 3424 12248 3476 12300
rect 6184 12248 6236 12300
rect 1492 12112 1544 12121
rect 1768 12044 1820 12096
rect 2780 12112 2832 12164
rect 4620 12180 4672 12232
rect 4804 12223 4856 12232
rect 4804 12189 4813 12223
rect 4813 12189 4847 12223
rect 4847 12189 4856 12223
rect 4804 12180 4856 12189
rect 3884 12112 3936 12164
rect 2228 12087 2280 12096
rect 2228 12053 2237 12087
rect 2237 12053 2271 12087
rect 2271 12053 2280 12087
rect 2228 12044 2280 12053
rect 2320 12087 2372 12096
rect 2320 12053 2329 12087
rect 2329 12053 2363 12087
rect 2363 12053 2372 12087
rect 2320 12044 2372 12053
rect 3148 12044 3200 12096
rect 3976 12044 4028 12096
rect 4436 12087 4488 12096
rect 4436 12053 4445 12087
rect 4445 12053 4479 12087
rect 4479 12053 4488 12087
rect 4436 12044 4488 12053
rect 4896 12112 4948 12164
rect 5264 12112 5316 12164
rect 5816 12044 5868 12096
rect 6092 12180 6144 12232
rect 8024 12180 8076 12232
rect 9128 12384 9180 12436
rect 10692 12384 10744 12436
rect 15016 12384 15068 12436
rect 14004 12316 14056 12368
rect 14648 12316 14700 12368
rect 9772 12291 9824 12300
rect 9772 12257 9781 12291
rect 9781 12257 9815 12291
rect 9815 12257 9824 12291
rect 9772 12248 9824 12257
rect 9128 12223 9180 12232
rect 9128 12189 9137 12223
rect 9137 12189 9171 12223
rect 9171 12189 9180 12223
rect 9128 12180 9180 12189
rect 10048 12180 10100 12232
rect 11796 12248 11848 12300
rect 11980 12291 12032 12300
rect 11980 12257 11989 12291
rect 11989 12257 12023 12291
rect 12023 12257 12032 12291
rect 11980 12248 12032 12257
rect 13544 12248 13596 12300
rect 15292 12248 15344 12300
rect 15936 12248 15988 12300
rect 11428 12223 11480 12232
rect 11428 12189 11437 12223
rect 11437 12189 11471 12223
rect 11471 12189 11480 12223
rect 11428 12180 11480 12189
rect 11888 12223 11940 12232
rect 11888 12189 11897 12223
rect 11897 12189 11931 12223
rect 11931 12189 11940 12223
rect 11888 12180 11940 12189
rect 6000 12112 6052 12164
rect 6644 12087 6696 12096
rect 6644 12053 6653 12087
rect 6653 12053 6687 12087
rect 6687 12053 6696 12087
rect 6644 12044 6696 12053
rect 7288 12112 7340 12164
rect 12256 12155 12308 12164
rect 12256 12121 12290 12155
rect 12290 12121 12308 12155
rect 12256 12112 12308 12121
rect 13912 12180 13964 12232
rect 14188 12180 14240 12232
rect 15476 12223 15528 12232
rect 15476 12189 15485 12223
rect 15485 12189 15519 12223
rect 15519 12189 15528 12223
rect 15476 12180 15528 12189
rect 15660 12180 15712 12232
rect 15752 12223 15804 12232
rect 15752 12189 15761 12223
rect 15761 12189 15795 12223
rect 15795 12189 15804 12223
rect 15752 12180 15804 12189
rect 14556 12112 14608 12164
rect 14924 12112 14976 12164
rect 8668 12087 8720 12096
rect 8668 12053 8677 12087
rect 8677 12053 8711 12087
rect 8711 12053 8720 12087
rect 8668 12044 8720 12053
rect 9036 12087 9088 12096
rect 9036 12053 9045 12087
rect 9045 12053 9079 12087
rect 9079 12053 9088 12087
rect 9036 12044 9088 12053
rect 10692 12044 10744 12096
rect 11704 12044 11756 12096
rect 13912 12044 13964 12096
rect 14096 12044 14148 12096
rect 14740 12044 14792 12096
rect 15200 12044 15252 12096
rect 15568 12044 15620 12096
rect 16028 12155 16080 12164
rect 16028 12121 16037 12155
rect 16037 12121 16071 12155
rect 16071 12121 16080 12155
rect 16028 12112 16080 12121
rect 16396 12112 16448 12164
rect 16212 12087 16264 12096
rect 16212 12053 16221 12087
rect 16221 12053 16255 12087
rect 16255 12053 16264 12087
rect 16212 12044 16264 12053
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 1492 11840 1544 11892
rect 2228 11840 2280 11892
rect 2872 11840 2924 11892
rect 1860 11772 1912 11824
rect 3976 11840 4028 11892
rect 4436 11840 4488 11892
rect 4896 11840 4948 11892
rect 5264 11840 5316 11892
rect 6184 11840 6236 11892
rect 8668 11840 8720 11892
rect 10784 11840 10836 11892
rect 11888 11840 11940 11892
rect 13544 11840 13596 11892
rect 13728 11840 13780 11892
rect 3148 11772 3200 11824
rect 3240 11815 3292 11824
rect 3240 11781 3249 11815
rect 3249 11781 3283 11815
rect 3283 11781 3292 11815
rect 3240 11772 3292 11781
rect 4804 11772 4856 11824
rect 5080 11772 5132 11824
rect 6460 11772 6512 11824
rect 8300 11772 8352 11824
rect 9864 11815 9916 11824
rect 9864 11781 9873 11815
rect 9873 11781 9907 11815
rect 9907 11781 9916 11815
rect 9864 11772 9916 11781
rect 11520 11772 11572 11824
rect 12348 11815 12400 11824
rect 12348 11781 12382 11815
rect 12382 11781 12400 11815
rect 12348 11772 12400 11781
rect 3424 11747 3476 11756
rect 3424 11713 3433 11747
rect 3433 11713 3467 11747
rect 3467 11713 3476 11747
rect 3424 11704 3476 11713
rect 3516 11704 3568 11756
rect 3976 11704 4028 11756
rect 4160 11747 4212 11756
rect 4160 11713 4169 11747
rect 4169 11713 4203 11747
rect 4203 11713 4212 11747
rect 4160 11704 4212 11713
rect 3884 11611 3936 11620
rect 3884 11577 3893 11611
rect 3893 11577 3927 11611
rect 3927 11577 3936 11611
rect 4712 11704 4764 11756
rect 5816 11747 5868 11756
rect 5816 11713 5825 11747
rect 5825 11713 5859 11747
rect 5859 11713 5868 11747
rect 5816 11704 5868 11713
rect 5632 11636 5684 11688
rect 7104 11704 7156 11756
rect 7932 11704 7984 11756
rect 8392 11704 8444 11756
rect 9312 11747 9364 11756
rect 9312 11713 9321 11747
rect 9321 11713 9355 11747
rect 9355 11713 9364 11747
rect 9312 11704 9364 11713
rect 9496 11747 9548 11756
rect 9496 11713 9505 11747
rect 9505 11713 9539 11747
rect 9539 11713 9548 11747
rect 9496 11704 9548 11713
rect 11428 11704 11480 11756
rect 12072 11747 12124 11756
rect 12072 11713 12081 11747
rect 12081 11713 12115 11747
rect 12115 11713 12124 11747
rect 12072 11704 12124 11713
rect 15108 11840 15160 11892
rect 13912 11704 13964 11756
rect 14832 11772 14884 11824
rect 14096 11747 14148 11756
rect 14096 11713 14105 11747
rect 14105 11713 14139 11747
rect 14139 11713 14148 11747
rect 14096 11704 14148 11713
rect 14372 11747 14424 11756
rect 8852 11636 8904 11688
rect 3884 11568 3936 11577
rect 5264 11568 5316 11620
rect 7196 11568 7248 11620
rect 7288 11611 7340 11620
rect 7288 11577 7297 11611
rect 7297 11577 7331 11611
rect 7331 11577 7340 11611
rect 7288 11568 7340 11577
rect 14004 11568 14056 11620
rect 2964 11500 3016 11552
rect 3056 11543 3108 11552
rect 3056 11509 3065 11543
rect 3065 11509 3099 11543
rect 3099 11509 3108 11543
rect 3056 11500 3108 11509
rect 3424 11500 3476 11552
rect 3516 11500 3568 11552
rect 6920 11500 6972 11552
rect 9220 11543 9272 11552
rect 9220 11509 9229 11543
rect 9229 11509 9263 11543
rect 9263 11509 9272 11543
rect 9220 11500 9272 11509
rect 9956 11500 10008 11552
rect 14372 11713 14381 11747
rect 14381 11713 14415 11747
rect 14415 11713 14424 11747
rect 14372 11704 14424 11713
rect 14280 11636 14332 11688
rect 14924 11747 14976 11756
rect 14924 11713 14933 11747
rect 14933 11713 14967 11747
rect 14967 11713 14976 11747
rect 14924 11704 14976 11713
rect 14832 11636 14884 11688
rect 14372 11500 14424 11552
rect 15108 11500 15160 11552
rect 16028 11500 16080 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 1768 11296 1820 11348
rect 2780 11339 2832 11348
rect 2780 11305 2789 11339
rect 2789 11305 2823 11339
rect 2823 11305 2832 11339
rect 2780 11296 2832 11305
rect 3148 11296 3200 11348
rect 5264 11339 5316 11348
rect 5264 11305 5273 11339
rect 5273 11305 5307 11339
rect 5307 11305 5316 11339
rect 5264 11296 5316 11305
rect 5724 11296 5776 11348
rect 6184 11296 6236 11348
rect 8576 11339 8628 11348
rect 8576 11305 8585 11339
rect 8585 11305 8619 11339
rect 8619 11305 8628 11339
rect 8576 11296 8628 11305
rect 4620 11228 4672 11280
rect 2780 11092 2832 11144
rect 6552 11160 6604 11212
rect 8944 11339 8996 11348
rect 8944 11305 8953 11339
rect 8953 11305 8987 11339
rect 8987 11305 8996 11339
rect 8944 11296 8996 11305
rect 9128 11296 9180 11348
rect 10508 11296 10560 11348
rect 9680 11228 9732 11280
rect 1676 11067 1728 11076
rect 1676 11033 1710 11067
rect 1710 11033 1728 11067
rect 1676 11024 1728 11033
rect 2228 11024 2280 11076
rect 4160 11092 4212 11144
rect 4528 11135 4580 11144
rect 4528 11101 4537 11135
rect 4537 11101 4571 11135
rect 4571 11101 4580 11135
rect 4528 11092 4580 11101
rect 3148 11024 3200 11076
rect 3792 11024 3844 11076
rect 4896 11092 4948 11144
rect 5724 11092 5776 11144
rect 13268 11296 13320 11348
rect 13452 11296 13504 11348
rect 14188 11296 14240 11348
rect 14556 11296 14608 11348
rect 14832 11339 14884 11348
rect 14832 11305 14841 11339
rect 14841 11305 14875 11339
rect 14875 11305 14884 11339
rect 14832 11296 14884 11305
rect 16212 11296 16264 11348
rect 13912 11203 13964 11212
rect 9220 11092 9272 11144
rect 9496 11135 9548 11144
rect 9496 11101 9505 11135
rect 9505 11101 9539 11135
rect 9539 11101 9548 11135
rect 9496 11092 9548 11101
rect 10232 11092 10284 11144
rect 11704 11135 11756 11144
rect 11704 11101 11713 11135
rect 11713 11101 11747 11135
rect 11747 11101 11756 11135
rect 11704 11092 11756 11101
rect 13912 11169 13921 11203
rect 13921 11169 13955 11203
rect 13955 11169 13964 11203
rect 13912 11160 13964 11169
rect 13820 11092 13872 11144
rect 15936 11228 15988 11280
rect 14924 11203 14976 11212
rect 14924 11169 14933 11203
rect 14933 11169 14967 11203
rect 14967 11169 14976 11203
rect 14924 11160 14976 11169
rect 4712 11024 4764 11076
rect 5540 11024 5592 11076
rect 5816 11024 5868 11076
rect 8852 11024 8904 11076
rect 9036 11024 9088 11076
rect 2044 10956 2096 11008
rect 2596 10956 2648 11008
rect 4804 10956 4856 11008
rect 5080 10956 5132 11008
rect 8116 10956 8168 11008
rect 8760 10956 8812 11008
rect 9128 10956 9180 11008
rect 12072 11024 12124 11076
rect 13912 11024 13964 11076
rect 12716 10956 12768 11008
rect 14096 10956 14148 11008
rect 14464 11135 14516 11144
rect 14464 11101 14473 11135
rect 14473 11101 14507 11135
rect 14507 11101 14516 11135
rect 14464 11092 14516 11101
rect 14556 11135 14608 11144
rect 14556 11101 14565 11135
rect 14565 11101 14599 11135
rect 14599 11101 14608 11135
rect 14556 11092 14608 11101
rect 15200 11135 15252 11144
rect 15200 11101 15234 11135
rect 15234 11101 15252 11135
rect 15200 11092 15252 11101
rect 14280 11024 14332 11076
rect 15292 11024 15344 11076
rect 15752 10956 15804 11008
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 1676 10795 1728 10804
rect 1676 10761 1685 10795
rect 1685 10761 1719 10795
rect 1719 10761 1728 10795
rect 1676 10752 1728 10761
rect 2044 10727 2096 10736
rect 2044 10693 2053 10727
rect 2053 10693 2087 10727
rect 2087 10693 2096 10727
rect 2044 10684 2096 10693
rect 3240 10752 3292 10804
rect 7196 10752 7248 10804
rect 13636 10795 13688 10804
rect 13636 10761 13645 10795
rect 13645 10761 13679 10795
rect 13679 10761 13688 10795
rect 13636 10752 13688 10761
rect 2596 10684 2648 10736
rect 5724 10727 5776 10736
rect 5724 10693 5733 10727
rect 5733 10693 5767 10727
rect 5767 10693 5776 10727
rect 5724 10684 5776 10693
rect 8668 10684 8720 10736
rect 2320 10616 2372 10668
rect 3516 10616 3568 10668
rect 4068 10659 4120 10668
rect 4068 10625 4077 10659
rect 4077 10625 4111 10659
rect 4111 10625 4120 10659
rect 4068 10616 4120 10625
rect 4712 10659 4764 10668
rect 4712 10625 4721 10659
rect 4721 10625 4755 10659
rect 4755 10625 4764 10659
rect 4712 10616 4764 10625
rect 4988 10659 5040 10668
rect 4988 10625 4997 10659
rect 4997 10625 5031 10659
rect 5031 10625 5040 10659
rect 4988 10616 5040 10625
rect 5264 10548 5316 10600
rect 3424 10480 3476 10532
rect 4528 10480 4580 10532
rect 4804 10480 4856 10532
rect 5632 10616 5684 10668
rect 7380 10659 7432 10668
rect 7380 10625 7389 10659
rect 7389 10625 7423 10659
rect 7423 10625 7432 10659
rect 7380 10616 7432 10625
rect 9036 10616 9088 10668
rect 8576 10548 8628 10600
rect 8852 10548 8904 10600
rect 9772 10616 9824 10668
rect 12072 10659 12124 10668
rect 12072 10625 12081 10659
rect 12081 10625 12115 10659
rect 12115 10625 12124 10659
rect 12072 10616 12124 10625
rect 15016 10752 15068 10804
rect 15292 10752 15344 10804
rect 15844 10752 15896 10804
rect 10508 10548 10560 10600
rect 14096 10659 14148 10668
rect 14096 10625 14105 10659
rect 14105 10625 14139 10659
rect 14139 10625 14148 10659
rect 14096 10616 14148 10625
rect 14372 10659 14424 10668
rect 14372 10625 14381 10659
rect 14381 10625 14415 10659
rect 14415 10625 14424 10659
rect 14372 10616 14424 10625
rect 14464 10659 14516 10668
rect 14464 10625 14473 10659
rect 14473 10625 14507 10659
rect 14507 10625 14516 10659
rect 14464 10616 14516 10625
rect 15476 10616 15528 10668
rect 14832 10548 14884 10600
rect 14924 10591 14976 10600
rect 14924 10557 14933 10591
rect 14933 10557 14967 10591
rect 14967 10557 14976 10591
rect 14924 10548 14976 10557
rect 8208 10480 8260 10532
rect 1860 10455 1912 10464
rect 1860 10421 1869 10455
rect 1869 10421 1903 10455
rect 1903 10421 1912 10455
rect 1860 10412 1912 10421
rect 5908 10455 5960 10464
rect 5908 10421 5917 10455
rect 5917 10421 5951 10455
rect 5951 10421 5960 10455
rect 5908 10412 5960 10421
rect 7656 10455 7708 10464
rect 7656 10421 7665 10455
rect 7665 10421 7699 10455
rect 7699 10421 7708 10455
rect 7656 10412 7708 10421
rect 8484 10455 8536 10464
rect 8484 10421 8493 10455
rect 8493 10421 8527 10455
rect 8527 10421 8536 10455
rect 8484 10412 8536 10421
rect 9128 10412 9180 10464
rect 10968 10412 11020 10464
rect 14004 10412 14056 10464
rect 15200 10412 15252 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 3240 10208 3292 10260
rect 5724 10208 5776 10260
rect 7196 10208 7248 10260
rect 7932 10208 7984 10260
rect 8668 10208 8720 10260
rect 8760 10251 8812 10260
rect 8760 10217 8769 10251
rect 8769 10217 8803 10251
rect 8803 10217 8812 10251
rect 8760 10208 8812 10217
rect 15292 10208 15344 10260
rect 16304 10208 16356 10260
rect 8116 10183 8168 10192
rect 8116 10149 8125 10183
rect 8125 10149 8159 10183
rect 8159 10149 8168 10183
rect 8116 10140 8168 10149
rect 2780 10072 2832 10124
rect 3976 10072 4028 10124
rect 3332 10047 3384 10056
rect 3332 10013 3341 10047
rect 3341 10013 3375 10047
rect 3375 10013 3384 10047
rect 3332 10004 3384 10013
rect 3608 10047 3660 10056
rect 3608 10013 3617 10047
rect 3617 10013 3651 10047
rect 3651 10013 3660 10047
rect 3608 10004 3660 10013
rect 4712 10004 4764 10056
rect 5448 10004 5500 10056
rect 6644 10047 6696 10056
rect 6644 10013 6653 10047
rect 6653 10013 6687 10047
rect 6687 10013 6696 10047
rect 6644 10004 6696 10013
rect 6920 10004 6972 10056
rect 8300 10004 8352 10056
rect 8484 10072 8536 10124
rect 12900 10072 12952 10124
rect 8576 10047 8628 10056
rect 8576 10013 8585 10047
rect 8585 10013 8619 10047
rect 8619 10013 8628 10047
rect 8576 10004 8628 10013
rect 4896 9936 4948 9988
rect 6368 9979 6420 9988
rect 6368 9945 6386 9979
rect 6386 9945 6420 9979
rect 6368 9936 6420 9945
rect 4528 9868 4580 9920
rect 6460 9868 6512 9920
rect 7380 9868 7432 9920
rect 9128 10004 9180 10056
rect 10508 10047 10560 10056
rect 10508 10013 10517 10047
rect 10517 10013 10551 10047
rect 10551 10013 10560 10047
rect 10508 10004 10560 10013
rect 13176 10047 13228 10056
rect 13176 10013 13185 10047
rect 13185 10013 13219 10047
rect 13219 10013 13228 10047
rect 13176 10004 13228 10013
rect 14096 10140 14148 10192
rect 14004 10004 14056 10056
rect 11428 9979 11480 9988
rect 11428 9945 11462 9979
rect 11462 9945 11480 9979
rect 11428 9936 11480 9945
rect 11520 9936 11572 9988
rect 12072 9936 12124 9988
rect 13084 9936 13136 9988
rect 16120 10004 16172 10056
rect 8760 9868 8812 9920
rect 12440 9868 12492 9920
rect 14832 9868 14884 9920
rect 15568 9868 15620 9920
rect 16120 9868 16172 9920
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 3332 9664 3384 9716
rect 4712 9664 4764 9716
rect 6368 9707 6420 9716
rect 6368 9673 6377 9707
rect 6377 9673 6411 9707
rect 6411 9673 6420 9707
rect 6368 9664 6420 9673
rect 6920 9707 6972 9716
rect 6920 9673 6929 9707
rect 6929 9673 6963 9707
rect 6963 9673 6972 9707
rect 6920 9664 6972 9673
rect 8576 9664 8628 9716
rect 9036 9707 9088 9716
rect 9036 9673 9045 9707
rect 9045 9673 9079 9707
rect 9079 9673 9088 9707
rect 9036 9664 9088 9673
rect 12900 9707 12952 9716
rect 12900 9673 12909 9707
rect 12909 9673 12943 9707
rect 12943 9673 12952 9707
rect 12900 9664 12952 9673
rect 3884 9596 3936 9648
rect 4620 9596 4672 9648
rect 5908 9596 5960 9648
rect 3332 9571 3384 9580
rect 3332 9537 3341 9571
rect 3341 9537 3375 9571
rect 3375 9537 3384 9571
rect 3332 9528 3384 9537
rect 2964 9460 3016 9512
rect 3608 9460 3660 9512
rect 3976 9528 4028 9580
rect 6276 9528 6328 9580
rect 5448 9460 5500 9512
rect 6460 9460 6512 9512
rect 8668 9528 8720 9580
rect 12440 9596 12492 9648
rect 14556 9664 14608 9716
rect 13820 9596 13872 9648
rect 14188 9596 14240 9648
rect 14832 9639 14884 9648
rect 14832 9605 14841 9639
rect 14841 9605 14875 9639
rect 14875 9605 14884 9639
rect 14832 9596 14884 9605
rect 9864 9528 9916 9580
rect 10416 9528 10468 9580
rect 11520 9571 11572 9580
rect 11520 9537 11529 9571
rect 11529 9537 11563 9571
rect 11563 9537 11572 9571
rect 11520 9528 11572 9537
rect 12624 9528 12676 9580
rect 13084 9571 13136 9580
rect 13084 9537 13093 9571
rect 13093 9537 13127 9571
rect 13127 9537 13136 9571
rect 13084 9528 13136 9537
rect 13360 9571 13412 9580
rect 13360 9537 13394 9571
rect 13394 9537 13412 9571
rect 13360 9528 13412 9537
rect 14740 9571 14792 9580
rect 14740 9537 14749 9571
rect 14749 9537 14783 9571
rect 14783 9537 14792 9571
rect 14740 9528 14792 9537
rect 15660 9596 15712 9648
rect 16120 9596 16172 9648
rect 15016 9528 15068 9580
rect 6736 9392 6788 9444
rect 8392 9503 8444 9512
rect 8392 9469 8401 9503
rect 8401 9469 8435 9503
rect 8435 9469 8444 9503
rect 8392 9460 8444 9469
rect 9588 9503 9640 9512
rect 9588 9469 9597 9503
rect 9597 9469 9631 9503
rect 9631 9469 9640 9503
rect 9588 9460 9640 9469
rect 16028 9571 16080 9580
rect 16028 9537 16037 9571
rect 16037 9537 16071 9571
rect 16071 9537 16080 9571
rect 16028 9528 16080 9537
rect 15936 9460 15988 9512
rect 14556 9435 14608 9444
rect 14556 9401 14565 9435
rect 14565 9401 14599 9435
rect 14599 9401 14608 9435
rect 14556 9392 14608 9401
rect 4068 9324 4120 9376
rect 6552 9367 6604 9376
rect 6552 9333 6561 9367
rect 6561 9333 6595 9367
rect 6595 9333 6604 9367
rect 6552 9324 6604 9333
rect 9220 9324 9272 9376
rect 10784 9324 10836 9376
rect 12256 9324 12308 9376
rect 13268 9324 13320 9376
rect 14464 9367 14516 9376
rect 14464 9333 14473 9367
rect 14473 9333 14507 9367
rect 14507 9333 14516 9367
rect 14464 9324 14516 9333
rect 14648 9324 14700 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 1860 9120 1912 9172
rect 3608 9163 3660 9172
rect 3608 9129 3617 9163
rect 3617 9129 3651 9163
rect 3651 9129 3660 9163
rect 3608 9120 3660 9129
rect 1584 9052 1636 9104
rect 2320 8984 2372 9036
rect 1492 8848 1544 8900
rect 2044 8848 2096 8900
rect 3148 8916 3200 8968
rect 3516 8916 3568 8968
rect 4068 9120 4120 9172
rect 4804 9120 4856 9172
rect 8392 9120 8444 9172
rect 8576 9163 8628 9172
rect 8576 9129 8585 9163
rect 8585 9129 8619 9163
rect 8619 9129 8628 9163
rect 8576 9120 8628 9129
rect 11428 9163 11480 9172
rect 11428 9129 11437 9163
rect 11437 9129 11471 9163
rect 11471 9129 11480 9163
rect 11428 9120 11480 9129
rect 13452 9163 13504 9172
rect 13452 9129 13461 9163
rect 13461 9129 13495 9163
rect 13495 9129 13504 9163
rect 13452 9120 13504 9129
rect 16212 9163 16264 9172
rect 16212 9129 16221 9163
rect 16221 9129 16255 9163
rect 16255 9129 16264 9163
rect 16212 9120 16264 9129
rect 6276 9052 6328 9104
rect 3700 8984 3752 9036
rect 3976 9027 4028 9036
rect 3976 8993 3985 9027
rect 3985 8993 4019 9027
rect 4019 8993 4028 9027
rect 3976 8984 4028 8993
rect 1768 8823 1820 8832
rect 1768 8789 1777 8823
rect 1777 8789 1811 8823
rect 1811 8789 1820 8823
rect 1768 8780 1820 8789
rect 2320 8823 2372 8832
rect 2320 8789 2329 8823
rect 2329 8789 2363 8823
rect 2363 8789 2372 8823
rect 2320 8780 2372 8789
rect 2964 8848 3016 8900
rect 3424 8891 3476 8900
rect 3424 8857 3433 8891
rect 3433 8857 3467 8891
rect 3467 8857 3476 8891
rect 3424 8848 3476 8857
rect 2872 8780 2924 8832
rect 3332 8780 3384 8832
rect 8300 8984 8352 9036
rect 12256 9052 12308 9104
rect 5264 8916 5316 8968
rect 5540 8916 5592 8968
rect 6368 8848 6420 8900
rect 6644 8848 6696 8900
rect 7656 8916 7708 8968
rect 8392 8891 8444 8900
rect 8392 8857 8401 8891
rect 8401 8857 8435 8891
rect 8435 8857 8444 8891
rect 8392 8848 8444 8857
rect 11980 9027 12032 9036
rect 11980 8993 11989 9027
rect 11989 8993 12023 9027
rect 12023 8993 12032 9027
rect 11980 8984 12032 8993
rect 12164 8984 12216 9036
rect 11704 8916 11756 8968
rect 13544 8959 13596 8968
rect 13544 8925 13553 8959
rect 13553 8925 13587 8959
rect 13587 8925 13596 8959
rect 13544 8916 13596 8925
rect 13820 8916 13872 8968
rect 14464 9052 14516 9104
rect 14924 8916 14976 8968
rect 15200 8959 15252 8968
rect 15200 8925 15209 8959
rect 15209 8925 15243 8959
rect 15243 8925 15252 8959
rect 15200 8916 15252 8925
rect 9864 8848 9916 8900
rect 12440 8848 12492 8900
rect 12532 8891 12584 8900
rect 12532 8857 12541 8891
rect 12541 8857 12575 8891
rect 12575 8857 12584 8891
rect 12532 8848 12584 8857
rect 15016 8848 15068 8900
rect 15384 8916 15436 8968
rect 15752 8959 15804 8968
rect 15752 8925 15761 8959
rect 15761 8925 15795 8959
rect 15795 8925 15804 8959
rect 15752 8916 15804 8925
rect 15844 8916 15896 8968
rect 15936 8891 15988 8900
rect 15936 8857 15945 8891
rect 15945 8857 15979 8891
rect 15979 8857 15988 8891
rect 15936 8848 15988 8857
rect 16120 8848 16172 8900
rect 8300 8780 8352 8832
rect 9036 8780 9088 8832
rect 11152 8780 11204 8832
rect 11888 8823 11940 8832
rect 11888 8789 11897 8823
rect 11897 8789 11931 8823
rect 11931 8789 11940 8823
rect 11888 8780 11940 8789
rect 12348 8780 12400 8832
rect 13912 8780 13964 8832
rect 14832 8823 14884 8832
rect 14832 8789 14841 8823
rect 14841 8789 14875 8823
rect 14875 8789 14884 8823
rect 14832 8780 14884 8789
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 2320 8576 2372 8628
rect 3884 8576 3936 8628
rect 4712 8576 4764 8628
rect 5356 8576 5408 8628
rect 8484 8576 8536 8628
rect 9772 8619 9824 8628
rect 9772 8585 9781 8619
rect 9781 8585 9815 8619
rect 9815 8585 9824 8619
rect 9772 8576 9824 8585
rect 10416 8619 10468 8628
rect 10416 8585 10425 8619
rect 10425 8585 10459 8619
rect 10459 8585 10468 8619
rect 10416 8576 10468 8585
rect 10784 8619 10836 8628
rect 10784 8585 10793 8619
rect 10793 8585 10827 8619
rect 10827 8585 10836 8619
rect 10784 8576 10836 8585
rect 12624 8576 12676 8628
rect 12900 8576 12952 8628
rect 2412 8508 2464 8560
rect 2504 8483 2556 8492
rect 2504 8449 2522 8483
rect 2522 8449 2556 8483
rect 2504 8440 2556 8449
rect 2872 8551 2924 8560
rect 2872 8517 2881 8551
rect 2881 8517 2915 8551
rect 2915 8517 2924 8551
rect 2872 8508 2924 8517
rect 2780 8483 2832 8492
rect 2780 8449 2789 8483
rect 2789 8449 2823 8483
rect 2823 8449 2832 8483
rect 2780 8440 2832 8449
rect 3976 8508 4028 8560
rect 5540 8508 5592 8560
rect 2964 8304 3016 8356
rect 3516 8483 3568 8492
rect 3516 8449 3525 8483
rect 3525 8449 3559 8483
rect 3559 8449 3568 8483
rect 3516 8440 3568 8449
rect 5448 8483 5500 8492
rect 5448 8449 5457 8483
rect 5457 8449 5491 8483
rect 5491 8449 5500 8483
rect 5448 8440 5500 8449
rect 8116 8508 8168 8560
rect 5724 8483 5776 8492
rect 5724 8449 5733 8483
rect 5733 8449 5767 8483
rect 5767 8449 5776 8483
rect 5724 8440 5776 8449
rect 6276 8440 6328 8492
rect 12808 8508 12860 8560
rect 8484 8440 8536 8492
rect 9864 8483 9916 8492
rect 9864 8449 9873 8483
rect 9873 8449 9907 8483
rect 9907 8449 9916 8483
rect 9864 8440 9916 8449
rect 4804 8372 4856 8424
rect 4068 8304 4120 8356
rect 5908 8372 5960 8424
rect 6736 8415 6788 8424
rect 6736 8381 6745 8415
rect 6745 8381 6779 8415
rect 6779 8381 6788 8415
rect 6736 8372 6788 8381
rect 5540 8347 5592 8356
rect 5540 8313 5549 8347
rect 5549 8313 5583 8347
rect 5583 8313 5592 8347
rect 5540 8304 5592 8313
rect 6368 8304 6420 8356
rect 9588 8372 9640 8424
rect 11888 8440 11940 8492
rect 13360 8619 13412 8628
rect 13360 8585 13369 8619
rect 13369 8585 13403 8619
rect 13403 8585 13412 8619
rect 13360 8576 13412 8585
rect 13728 8576 13780 8628
rect 13728 8483 13780 8492
rect 13728 8449 13737 8483
rect 13737 8449 13771 8483
rect 13771 8449 13780 8483
rect 13728 8440 13780 8449
rect 13912 8440 13964 8492
rect 14004 8483 14056 8492
rect 14004 8449 14013 8483
rect 14013 8449 14047 8483
rect 14047 8449 14056 8483
rect 14648 8508 14700 8560
rect 14004 8440 14056 8449
rect 15752 8576 15804 8628
rect 14832 8508 14884 8560
rect 10968 8415 11020 8424
rect 10968 8381 10977 8415
rect 10977 8381 11011 8415
rect 11011 8381 11020 8415
rect 10968 8372 11020 8381
rect 12348 8415 12400 8424
rect 12348 8381 12357 8415
rect 12357 8381 12391 8415
rect 12391 8381 12400 8415
rect 12348 8372 12400 8381
rect 13084 8415 13136 8424
rect 13084 8381 13093 8415
rect 13093 8381 13127 8415
rect 13127 8381 13136 8415
rect 13084 8372 13136 8381
rect 13360 8372 13412 8424
rect 14372 8304 14424 8356
rect 3148 8236 3200 8288
rect 4620 8236 4672 8288
rect 5356 8236 5408 8288
rect 9772 8236 9824 8288
rect 10692 8236 10744 8288
rect 11244 8236 11296 8288
rect 11796 8236 11848 8288
rect 12992 8236 13044 8288
rect 15752 8440 15804 8492
rect 14924 8415 14976 8424
rect 14924 8381 14933 8415
rect 14933 8381 14967 8415
rect 14967 8381 14976 8415
rect 14924 8372 14976 8381
rect 15200 8236 15252 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 2780 8032 2832 8084
rect 2872 8032 2924 8084
rect 2596 7964 2648 8016
rect 8392 8032 8444 8084
rect 8944 8075 8996 8084
rect 8944 8041 8953 8075
rect 8953 8041 8987 8075
rect 8987 8041 8996 8075
rect 8944 8032 8996 8041
rect 11060 8075 11112 8084
rect 5448 7964 5500 8016
rect 5632 7964 5684 8016
rect 6276 7964 6328 8016
rect 11060 8041 11069 8075
rect 11069 8041 11103 8075
rect 11103 8041 11112 8075
rect 11060 8032 11112 8041
rect 11704 8032 11756 8084
rect 12164 8032 12216 8084
rect 12716 8032 12768 8084
rect 13452 8032 13504 8084
rect 16028 8032 16080 8084
rect 1676 7828 1728 7880
rect 1860 7871 1912 7880
rect 1860 7837 1894 7871
rect 1894 7837 1912 7871
rect 1860 7828 1912 7837
rect 3056 7828 3108 7880
rect 3516 7828 3568 7880
rect 3976 7828 4028 7880
rect 4160 7871 4212 7880
rect 4160 7837 4169 7871
rect 4169 7837 4203 7871
rect 4203 7837 4212 7871
rect 4160 7828 4212 7837
rect 5724 7828 5776 7880
rect 6092 7828 6144 7880
rect 6276 7828 6328 7880
rect 6736 7871 6788 7880
rect 6736 7837 6745 7871
rect 6745 7837 6779 7871
rect 6779 7837 6788 7871
rect 6736 7828 6788 7837
rect 9772 7964 9824 8016
rect 12808 7964 12860 8016
rect 14832 7964 14884 8016
rect 8576 7896 8628 7948
rect 2412 7760 2464 7812
rect 4804 7760 4856 7812
rect 6920 7760 6972 7812
rect 9128 7760 9180 7812
rect 9864 7828 9916 7880
rect 12532 7896 12584 7948
rect 14924 7939 14976 7948
rect 14924 7905 14933 7939
rect 14933 7905 14967 7939
rect 14967 7905 14976 7939
rect 14924 7896 14976 7905
rect 10416 7760 10468 7812
rect 10600 7803 10652 7812
rect 10600 7769 10618 7803
rect 10618 7769 10652 7803
rect 10600 7760 10652 7769
rect 2872 7692 2924 7744
rect 3148 7692 3200 7744
rect 3424 7692 3476 7744
rect 4252 7735 4304 7744
rect 4252 7701 4261 7735
rect 4261 7701 4295 7735
rect 4295 7701 4304 7735
rect 4252 7692 4304 7701
rect 5264 7692 5316 7744
rect 5356 7735 5408 7744
rect 5356 7701 5365 7735
rect 5365 7701 5399 7735
rect 5399 7701 5408 7735
rect 5356 7692 5408 7701
rect 5724 7692 5776 7744
rect 6000 7735 6052 7744
rect 6000 7701 6009 7735
rect 6009 7701 6043 7735
rect 6043 7701 6052 7735
rect 6000 7692 6052 7701
rect 6092 7735 6144 7744
rect 6092 7701 6101 7735
rect 6101 7701 6135 7735
rect 6135 7701 6144 7735
rect 6092 7692 6144 7701
rect 6736 7692 6788 7744
rect 7104 7735 7156 7744
rect 7104 7701 7113 7735
rect 7113 7701 7147 7735
rect 7147 7701 7156 7735
rect 7104 7692 7156 7701
rect 9956 7692 10008 7744
rect 11244 7828 11296 7880
rect 11796 7871 11848 7880
rect 11796 7837 11830 7871
rect 11830 7837 11848 7871
rect 11796 7828 11848 7837
rect 12900 7828 12952 7880
rect 13544 7828 13596 7880
rect 13636 7871 13688 7880
rect 13636 7837 13645 7871
rect 13645 7837 13679 7871
rect 13679 7837 13688 7871
rect 13636 7828 13688 7837
rect 13728 7828 13780 7880
rect 14004 7828 14056 7880
rect 14280 7871 14332 7880
rect 14280 7837 14289 7871
rect 14289 7837 14323 7871
rect 14323 7837 14332 7871
rect 14280 7828 14332 7837
rect 14372 7871 14424 7880
rect 14372 7837 14381 7871
rect 14381 7837 14415 7871
rect 14415 7837 14424 7871
rect 14372 7828 14424 7837
rect 14464 7871 14516 7880
rect 14464 7837 14473 7871
rect 14473 7837 14507 7871
rect 14507 7837 14516 7871
rect 14464 7828 14516 7837
rect 15200 7871 15252 7880
rect 15200 7837 15234 7871
rect 15234 7837 15252 7871
rect 15200 7828 15252 7837
rect 12164 7760 12216 7812
rect 15108 7760 15160 7812
rect 14740 7735 14792 7744
rect 14740 7701 14749 7735
rect 14749 7701 14783 7735
rect 14783 7701 14792 7735
rect 14740 7692 14792 7701
rect 14832 7692 14884 7744
rect 15016 7692 15068 7744
rect 16304 7692 16356 7744
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 2964 7488 3016 7540
rect 3056 7531 3108 7540
rect 3056 7497 3065 7531
rect 3065 7497 3099 7531
rect 3099 7497 3108 7531
rect 3056 7488 3108 7497
rect 1492 7463 1544 7472
rect 1492 7429 1501 7463
rect 1501 7429 1535 7463
rect 1535 7429 1544 7463
rect 1492 7420 1544 7429
rect 4252 7488 4304 7540
rect 4712 7531 4764 7540
rect 4712 7497 4721 7531
rect 4721 7497 4755 7531
rect 4755 7497 4764 7531
rect 4712 7488 4764 7497
rect 6092 7488 6144 7540
rect 6184 7531 6236 7540
rect 6184 7497 6193 7531
rect 6193 7497 6227 7531
rect 6227 7497 6236 7531
rect 6184 7488 6236 7497
rect 8484 7488 8536 7540
rect 9588 7488 9640 7540
rect 11336 7488 11388 7540
rect 13636 7488 13688 7540
rect 16212 7531 16264 7540
rect 16212 7497 16221 7531
rect 16221 7497 16255 7531
rect 16255 7497 16264 7531
rect 16212 7488 16264 7497
rect 1584 7395 1636 7404
rect 1584 7361 1593 7395
rect 1593 7361 1627 7395
rect 1627 7361 1636 7395
rect 1584 7352 1636 7361
rect 1676 7395 1728 7404
rect 1676 7361 1685 7395
rect 1685 7361 1719 7395
rect 1719 7361 1728 7395
rect 1676 7352 1728 7361
rect 2228 7352 2280 7404
rect 3976 7395 4028 7404
rect 3976 7361 3985 7395
rect 3985 7361 4019 7395
rect 4019 7361 4028 7395
rect 3976 7352 4028 7361
rect 4068 7395 4120 7404
rect 4068 7361 4077 7395
rect 4077 7361 4111 7395
rect 4111 7361 4120 7395
rect 4068 7352 4120 7361
rect 4712 7395 4764 7404
rect 4712 7361 4721 7395
rect 4721 7361 4755 7395
rect 4755 7361 4764 7395
rect 4712 7352 4764 7361
rect 5356 7352 5408 7404
rect 5632 7352 5684 7404
rect 6368 7395 6420 7404
rect 6368 7361 6377 7395
rect 6377 7361 6411 7395
rect 6411 7361 6420 7395
rect 6368 7352 6420 7361
rect 7012 7352 7064 7404
rect 8300 7352 8352 7404
rect 8760 7352 8812 7404
rect 9864 7420 9916 7472
rect 1952 7148 2004 7200
rect 2320 7148 2372 7200
rect 4620 7216 4672 7268
rect 8208 7284 8260 7336
rect 8668 7284 8720 7336
rect 9680 7352 9732 7404
rect 11152 7395 11204 7404
rect 11152 7361 11161 7395
rect 11161 7361 11195 7395
rect 11195 7361 11204 7395
rect 11152 7352 11204 7361
rect 12532 7420 12584 7472
rect 11612 7352 11664 7404
rect 14924 7420 14976 7472
rect 13176 7352 13228 7404
rect 14740 7352 14792 7404
rect 16028 7395 16080 7404
rect 16028 7361 16037 7395
rect 16037 7361 16071 7395
rect 16071 7361 16080 7395
rect 16028 7352 16080 7361
rect 12992 7216 13044 7268
rect 6000 7148 6052 7200
rect 6644 7148 6696 7200
rect 8024 7148 8076 7200
rect 10416 7191 10468 7200
rect 10416 7157 10425 7191
rect 10425 7157 10459 7191
rect 10459 7157 10468 7191
rect 10416 7148 10468 7157
rect 10784 7148 10836 7200
rect 14004 7148 14056 7200
rect 14556 7191 14608 7200
rect 14556 7157 14565 7191
rect 14565 7157 14599 7191
rect 14599 7157 14608 7191
rect 14556 7148 14608 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 2320 6987 2372 6996
rect 2320 6953 2329 6987
rect 2329 6953 2363 6987
rect 2363 6953 2372 6987
rect 2320 6944 2372 6953
rect 2412 6876 2464 6928
rect 3148 6987 3200 6996
rect 3148 6953 3157 6987
rect 3157 6953 3191 6987
rect 3191 6953 3200 6987
rect 3148 6944 3200 6953
rect 3424 6987 3476 6996
rect 3424 6953 3433 6987
rect 3433 6953 3467 6987
rect 3467 6953 3476 6987
rect 3424 6944 3476 6953
rect 4804 6944 4856 6996
rect 5172 6987 5224 6996
rect 5172 6953 5181 6987
rect 5181 6953 5215 6987
rect 5215 6953 5224 6987
rect 5172 6944 5224 6953
rect 5724 6944 5776 6996
rect 6184 6944 6236 6996
rect 6736 6944 6788 6996
rect 7012 6987 7064 6996
rect 7012 6953 7021 6987
rect 7021 6953 7055 6987
rect 7055 6953 7064 6987
rect 7012 6944 7064 6953
rect 11336 6987 11388 6996
rect 11336 6953 11345 6987
rect 11345 6953 11379 6987
rect 11379 6953 11388 6987
rect 11336 6944 11388 6953
rect 11612 6944 11664 6996
rect 13176 6944 13228 6996
rect 14464 6944 14516 6996
rect 2320 6808 2372 6860
rect 2780 6808 2832 6860
rect 3240 6808 3292 6860
rect 9128 6808 9180 6860
rect 11060 6808 11112 6860
rect 12164 6851 12216 6860
rect 12164 6817 12173 6851
rect 12173 6817 12207 6851
rect 12207 6817 12216 6851
rect 12164 6808 12216 6817
rect 14924 6851 14976 6860
rect 14924 6817 14933 6851
rect 14933 6817 14967 6851
rect 14967 6817 14976 6851
rect 14924 6808 14976 6817
rect 2872 6740 2924 6792
rect 2228 6672 2280 6724
rect 2320 6715 2372 6724
rect 2320 6681 2345 6715
rect 2345 6681 2372 6715
rect 2320 6672 2372 6681
rect 2688 6672 2740 6724
rect 2964 6715 3016 6724
rect 3884 6740 3936 6792
rect 4620 6740 4672 6792
rect 2964 6681 2989 6715
rect 2989 6681 3016 6715
rect 2964 6672 3016 6681
rect 2504 6647 2556 6656
rect 2504 6613 2513 6647
rect 2513 6613 2547 6647
rect 2547 6613 2556 6647
rect 2504 6604 2556 6613
rect 2596 6604 2648 6656
rect 2872 6604 2924 6656
rect 3976 6604 4028 6656
rect 5448 6783 5500 6792
rect 5448 6749 5457 6783
rect 5457 6749 5491 6783
rect 5491 6749 5500 6783
rect 5448 6740 5500 6749
rect 5632 6740 5684 6792
rect 6920 6740 6972 6792
rect 8024 6783 8076 6792
rect 8024 6749 8033 6783
rect 8033 6749 8067 6783
rect 8067 6749 8076 6783
rect 8024 6740 8076 6749
rect 5356 6715 5408 6724
rect 5356 6681 5365 6715
rect 5365 6681 5399 6715
rect 5399 6681 5408 6715
rect 5356 6672 5408 6681
rect 5908 6672 5960 6724
rect 7104 6672 7156 6724
rect 10692 6783 10744 6792
rect 10692 6749 10701 6783
rect 10701 6749 10735 6783
rect 10735 6749 10744 6783
rect 10692 6740 10744 6749
rect 10784 6740 10836 6792
rect 12624 6740 12676 6792
rect 13268 6783 13320 6792
rect 13268 6749 13277 6783
rect 13277 6749 13311 6783
rect 13311 6749 13320 6783
rect 13268 6740 13320 6749
rect 13360 6783 13412 6792
rect 13360 6749 13369 6783
rect 13369 6749 13403 6783
rect 13403 6749 13412 6783
rect 13360 6740 13412 6749
rect 13544 6740 13596 6792
rect 13728 6740 13780 6792
rect 14004 6740 14056 6792
rect 14188 6740 14240 6792
rect 14648 6740 14700 6792
rect 11152 6672 11204 6724
rect 12992 6672 13044 6724
rect 14372 6715 14424 6724
rect 14372 6681 14381 6715
rect 14381 6681 14415 6715
rect 14415 6681 14424 6715
rect 14372 6672 14424 6681
rect 14556 6672 14608 6724
rect 15568 6672 15620 6724
rect 10048 6604 10100 6656
rect 11888 6647 11940 6656
rect 11888 6613 11897 6647
rect 11897 6613 11931 6647
rect 11931 6613 11940 6647
rect 11888 6604 11940 6613
rect 13176 6604 13228 6656
rect 13636 6604 13688 6656
rect 14464 6604 14516 6656
rect 15936 6604 15988 6656
rect 16212 6604 16264 6656
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 3884 6400 3936 6452
rect 5540 6400 5592 6452
rect 3148 6332 3200 6384
rect 3240 6307 3292 6316
rect 3240 6273 3249 6307
rect 3249 6273 3283 6307
rect 3283 6273 3292 6307
rect 3240 6264 3292 6273
rect 6920 6400 6972 6452
rect 8852 6400 8904 6452
rect 10968 6400 11020 6452
rect 11244 6400 11296 6452
rect 11980 6400 12032 6452
rect 13084 6400 13136 6452
rect 13544 6443 13596 6452
rect 13544 6409 13553 6443
rect 13553 6409 13587 6443
rect 13587 6409 13596 6443
rect 13544 6400 13596 6409
rect 14280 6400 14332 6452
rect 15200 6400 15252 6452
rect 15568 6443 15620 6452
rect 15568 6409 15577 6443
rect 15577 6409 15611 6443
rect 15611 6409 15620 6443
rect 15568 6400 15620 6409
rect 15660 6443 15712 6452
rect 15660 6409 15669 6443
rect 15669 6409 15703 6443
rect 15703 6409 15712 6443
rect 15660 6400 15712 6409
rect 2872 6239 2924 6248
rect 2872 6205 2881 6239
rect 2881 6205 2915 6239
rect 2915 6205 2924 6239
rect 2872 6196 2924 6205
rect 4068 6264 4120 6316
rect 6736 6264 6788 6316
rect 6644 6196 6696 6248
rect 9680 6307 9732 6316
rect 9680 6273 9689 6307
rect 9689 6273 9723 6307
rect 9723 6273 9732 6307
rect 9680 6264 9732 6273
rect 9772 6307 9824 6316
rect 9772 6273 9781 6307
rect 9781 6273 9815 6307
rect 9815 6273 9824 6307
rect 9772 6264 9824 6273
rect 9956 6264 10008 6316
rect 10048 6239 10100 6248
rect 10048 6205 10057 6239
rect 10057 6205 10091 6239
rect 10091 6205 10100 6239
rect 10048 6196 10100 6205
rect 11152 6264 11204 6316
rect 12900 6332 12952 6384
rect 11060 6196 11112 6248
rect 11244 6196 11296 6248
rect 13544 6264 13596 6316
rect 6184 6128 6236 6180
rect 13636 6196 13688 6248
rect 13912 6307 13964 6316
rect 13912 6273 13921 6307
rect 13921 6273 13955 6307
rect 13955 6273 13964 6307
rect 13912 6264 13964 6273
rect 14464 6375 14516 6384
rect 14464 6341 14473 6375
rect 14473 6341 14507 6375
rect 14507 6341 14516 6375
rect 14464 6332 14516 6341
rect 14648 6332 14700 6384
rect 16028 6400 16080 6452
rect 14372 6264 14424 6316
rect 14556 6307 14608 6316
rect 14556 6273 14565 6307
rect 14565 6273 14599 6307
rect 14599 6273 14608 6307
rect 14556 6264 14608 6273
rect 15016 6262 15068 6314
rect 14004 6196 14056 6248
rect 14096 6196 14148 6248
rect 15209 6307 15261 6316
rect 15209 6273 15212 6307
rect 15212 6273 15246 6307
rect 15246 6273 15261 6307
rect 15209 6264 15261 6273
rect 15752 6264 15804 6316
rect 16028 6307 16080 6316
rect 16028 6273 16037 6307
rect 16037 6273 16071 6307
rect 16071 6273 16080 6307
rect 16028 6264 16080 6273
rect 16212 6307 16264 6316
rect 16212 6273 16221 6307
rect 16221 6273 16255 6307
rect 16255 6273 16264 6307
rect 16212 6264 16264 6273
rect 3424 6060 3476 6112
rect 4712 6103 4764 6112
rect 4712 6069 4721 6103
rect 4721 6069 4755 6103
rect 4755 6069 4764 6103
rect 4712 6060 4764 6069
rect 4804 6060 4856 6112
rect 5448 6103 5500 6112
rect 5448 6069 5457 6103
rect 5457 6069 5491 6103
rect 5491 6069 5500 6103
rect 5448 6060 5500 6069
rect 9956 6103 10008 6112
rect 9956 6069 9965 6103
rect 9965 6069 9999 6103
rect 9999 6069 10008 6103
rect 9956 6060 10008 6069
rect 10876 6060 10928 6112
rect 11704 6103 11756 6112
rect 11704 6069 11713 6103
rect 11713 6069 11747 6103
rect 11747 6069 11756 6103
rect 11704 6060 11756 6069
rect 15200 6128 15252 6180
rect 12716 6060 12768 6112
rect 12808 6103 12860 6112
rect 12808 6069 12817 6103
rect 12817 6069 12851 6103
rect 12851 6069 12860 6103
rect 12808 6060 12860 6069
rect 13728 6060 13780 6112
rect 13820 6060 13872 6112
rect 15016 6060 15068 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 3884 5856 3936 5908
rect 6920 5856 6972 5908
rect 10600 5899 10652 5908
rect 10600 5865 10609 5899
rect 10609 5865 10643 5899
rect 10643 5865 10652 5899
rect 10600 5856 10652 5865
rect 12072 5856 12124 5908
rect 14096 5856 14148 5908
rect 2688 5788 2740 5840
rect 4068 5788 4120 5840
rect 14188 5788 14240 5840
rect 14740 5831 14792 5840
rect 14740 5797 14749 5831
rect 14749 5797 14783 5831
rect 14783 5797 14792 5831
rect 14740 5788 14792 5797
rect 4712 5584 4764 5636
rect 5448 5584 5500 5636
rect 9956 5652 10008 5704
rect 10784 5695 10836 5704
rect 10784 5661 10793 5695
rect 10793 5661 10827 5695
rect 10827 5661 10836 5695
rect 10784 5652 10836 5661
rect 10876 5652 10928 5704
rect 11704 5652 11756 5704
rect 12256 5652 12308 5704
rect 12808 5695 12860 5704
rect 12808 5661 12817 5695
rect 12817 5661 12851 5695
rect 12851 5661 12860 5695
rect 12808 5652 12860 5661
rect 13912 5720 13964 5772
rect 16028 5856 16080 5908
rect 15292 5788 15344 5840
rect 14188 5652 14240 5704
rect 13084 5627 13136 5636
rect 13084 5593 13093 5627
rect 13093 5593 13127 5627
rect 13127 5593 13136 5627
rect 13084 5584 13136 5593
rect 13544 5627 13596 5636
rect 13544 5593 13553 5627
rect 13553 5593 13587 5627
rect 13587 5593 13596 5627
rect 13544 5584 13596 5593
rect 5540 5516 5592 5568
rect 10968 5516 11020 5568
rect 11520 5516 11572 5568
rect 12348 5559 12400 5568
rect 12348 5525 12357 5559
rect 12357 5525 12391 5559
rect 12391 5525 12400 5559
rect 12348 5516 12400 5525
rect 13636 5516 13688 5568
rect 13820 5584 13872 5636
rect 14648 5652 14700 5704
rect 14188 5516 14240 5568
rect 14372 5516 14424 5568
rect 14556 5584 14608 5636
rect 14740 5584 14792 5636
rect 15016 5627 15068 5636
rect 15016 5593 15025 5627
rect 15025 5593 15059 5627
rect 15059 5593 15068 5627
rect 15016 5584 15068 5593
rect 15660 5652 15712 5704
rect 15844 5695 15896 5704
rect 15844 5661 15853 5695
rect 15853 5661 15887 5695
rect 15887 5661 15896 5695
rect 15844 5652 15896 5661
rect 15936 5695 15988 5704
rect 15936 5661 15945 5695
rect 15945 5661 15979 5695
rect 15979 5661 15988 5695
rect 15936 5652 15988 5661
rect 16120 5695 16172 5704
rect 16120 5661 16129 5695
rect 16129 5661 16163 5695
rect 16163 5661 16172 5695
rect 16120 5652 16172 5661
rect 14832 5516 14884 5568
rect 15292 5516 15344 5568
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 9404 5312 9456 5364
rect 10784 5312 10836 5364
rect 11980 5355 12032 5364
rect 11980 5321 11989 5355
rect 11989 5321 12023 5355
rect 12023 5321 12032 5355
rect 11980 5312 12032 5321
rect 12716 5312 12768 5364
rect 15384 5312 15436 5364
rect 9220 5244 9272 5296
rect 9496 5244 9548 5296
rect 11060 5244 11112 5296
rect 10876 5176 10928 5228
rect 11704 5176 11756 5228
rect 12900 5219 12952 5228
rect 12900 5185 12909 5219
rect 12909 5185 12943 5219
rect 12943 5185 12952 5219
rect 12900 5176 12952 5185
rect 13360 5244 13412 5296
rect 13820 5244 13872 5296
rect 9496 5040 9548 5092
rect 12072 5151 12124 5160
rect 12072 5117 12081 5151
rect 12081 5117 12115 5151
rect 12115 5117 12124 5151
rect 12072 5108 12124 5117
rect 12164 5151 12216 5160
rect 12164 5117 12173 5151
rect 12173 5117 12207 5151
rect 12207 5117 12216 5151
rect 12164 5108 12216 5117
rect 12992 5151 13044 5160
rect 12992 5117 13001 5151
rect 13001 5117 13035 5151
rect 13035 5117 13044 5151
rect 12992 5108 13044 5117
rect 12900 5040 12952 5092
rect 11152 5015 11204 5024
rect 11152 4981 11161 5015
rect 11161 4981 11195 5015
rect 11195 4981 11204 5015
rect 11152 4972 11204 4981
rect 11704 4972 11756 5024
rect 12440 5015 12492 5024
rect 12440 4981 12449 5015
rect 12449 4981 12483 5015
rect 12483 4981 12492 5015
rect 12440 4972 12492 4981
rect 13360 4972 13412 5024
rect 13636 5040 13688 5092
rect 13912 5219 13964 5228
rect 13912 5185 13921 5219
rect 13921 5185 13955 5219
rect 13955 5185 13964 5219
rect 13912 5176 13964 5185
rect 14372 5176 14424 5228
rect 15108 5219 15160 5228
rect 15108 5185 15117 5219
rect 15117 5185 15151 5219
rect 15151 5185 15160 5219
rect 15108 5176 15160 5185
rect 15200 5219 15252 5228
rect 15200 5185 15209 5219
rect 15209 5185 15243 5219
rect 15243 5185 15252 5219
rect 15200 5176 15252 5185
rect 15384 5219 15436 5228
rect 15384 5185 15393 5219
rect 15393 5185 15427 5219
rect 15427 5185 15436 5219
rect 15384 5176 15436 5185
rect 16120 5219 16172 5228
rect 14188 5108 14240 5160
rect 14648 5108 14700 5160
rect 13912 5040 13964 5092
rect 14372 4972 14424 5024
rect 14740 5015 14792 5024
rect 14740 4981 14749 5015
rect 14749 4981 14783 5015
rect 14783 4981 14792 5015
rect 14740 4972 14792 4981
rect 15108 5040 15160 5092
rect 16120 5185 16129 5219
rect 16129 5185 16163 5219
rect 16163 5185 16172 5219
rect 16120 5176 16172 5185
rect 15384 4972 15436 5024
rect 15476 5015 15528 5024
rect 15476 4981 15485 5015
rect 15485 4981 15519 5015
rect 15519 4981 15528 5015
rect 15476 4972 15528 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 8944 4768 8996 4820
rect 11152 4811 11204 4820
rect 11152 4777 11161 4811
rect 11161 4777 11195 4811
rect 11195 4777 11204 4811
rect 11152 4768 11204 4777
rect 12716 4768 12768 4820
rect 14280 4768 14332 4820
rect 15844 4700 15896 4752
rect 9128 4632 9180 4684
rect 12900 4632 12952 4684
rect 8852 4564 8904 4616
rect 9312 4564 9364 4616
rect 9404 4607 9456 4616
rect 9404 4573 9413 4607
rect 9413 4573 9447 4607
rect 9447 4573 9456 4607
rect 9404 4564 9456 4573
rect 9496 4607 9548 4616
rect 9496 4573 9505 4607
rect 9505 4573 9539 4607
rect 9539 4573 9548 4607
rect 9496 4564 9548 4573
rect 9864 4564 9916 4616
rect 11428 4607 11480 4616
rect 11428 4573 11437 4607
rect 11437 4573 11471 4607
rect 11471 4573 11480 4607
rect 11428 4564 11480 4573
rect 11704 4607 11756 4616
rect 11704 4573 11738 4607
rect 11738 4573 11756 4607
rect 11704 4564 11756 4573
rect 11612 4496 11664 4548
rect 14372 4564 14424 4616
rect 14648 4564 14700 4616
rect 14924 4564 14976 4616
rect 9588 4428 9640 4480
rect 10784 4428 10836 4480
rect 12072 4428 12124 4480
rect 14740 4496 14792 4548
rect 16028 4607 16080 4616
rect 16028 4573 16037 4607
rect 16037 4573 16071 4607
rect 16071 4573 16080 4607
rect 16028 4564 16080 4573
rect 16120 4564 16172 4616
rect 16304 4496 16356 4548
rect 12900 4428 12952 4480
rect 15568 4471 15620 4480
rect 15568 4437 15577 4471
rect 15577 4437 15611 4471
rect 15611 4437 15620 4471
rect 15568 4428 15620 4437
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 10968 4224 11020 4276
rect 11612 4267 11664 4276
rect 11612 4233 11621 4267
rect 11621 4233 11655 4267
rect 11655 4233 11664 4267
rect 11612 4224 11664 4233
rect 8852 4156 8904 4208
rect 9312 4199 9364 4208
rect 9312 4165 9321 4199
rect 9321 4165 9355 4199
rect 9355 4165 9364 4199
rect 9312 4156 9364 4165
rect 9772 4156 9824 4208
rect 12900 4156 12952 4208
rect 9128 4131 9180 4140
rect 9128 4097 9137 4131
rect 9137 4097 9171 4131
rect 9171 4097 9180 4131
rect 9128 4088 9180 4097
rect 9588 4131 9640 4140
rect 9588 4097 9597 4131
rect 9597 4097 9631 4131
rect 9631 4097 9640 4131
rect 9588 4088 9640 4097
rect 10416 4088 10468 4140
rect 13820 4156 13872 4208
rect 14924 4156 14976 4208
rect 13360 4131 13412 4140
rect 13360 4097 13394 4131
rect 13394 4097 13412 4131
rect 13360 4088 13412 4097
rect 15476 4088 15528 4140
rect 9404 4020 9456 4072
rect 9864 4063 9916 4072
rect 9864 4029 9873 4063
rect 9873 4029 9907 4063
rect 9907 4029 9916 4063
rect 9864 4020 9916 4029
rect 8024 3927 8076 3936
rect 8024 3893 8033 3927
rect 8033 3893 8067 3927
rect 8067 3893 8076 3927
rect 8024 3884 8076 3893
rect 8944 3927 8996 3936
rect 8944 3893 8953 3927
rect 8953 3893 8987 3927
rect 8987 3893 8996 3927
rect 8944 3884 8996 3893
rect 11244 3995 11296 4004
rect 11244 3961 11253 3995
rect 11253 3961 11287 3995
rect 11287 3961 11296 3995
rect 11244 3952 11296 3961
rect 15016 3952 15068 4004
rect 10876 3884 10928 3936
rect 14464 3927 14516 3936
rect 14464 3893 14473 3927
rect 14473 3893 14507 3927
rect 14507 3893 14516 3927
rect 14464 3884 14516 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 9772 3723 9824 3732
rect 9772 3689 9781 3723
rect 9781 3689 9815 3723
rect 9815 3689 9824 3723
rect 9772 3680 9824 3689
rect 10876 3680 10928 3732
rect 12164 3680 12216 3732
rect 14188 3680 14240 3732
rect 8024 3544 8076 3596
rect 8760 3519 8812 3528
rect 8760 3485 8769 3519
rect 8769 3485 8803 3519
rect 8803 3485 8812 3519
rect 8760 3476 8812 3485
rect 9220 3519 9272 3528
rect 9220 3485 9229 3519
rect 9229 3485 9263 3519
rect 9263 3485 9272 3519
rect 9220 3476 9272 3485
rect 9864 3587 9916 3596
rect 9864 3553 9873 3587
rect 9873 3553 9907 3587
rect 9907 3553 9916 3587
rect 9864 3544 9916 3553
rect 11428 3544 11480 3596
rect 11980 3587 12032 3596
rect 11980 3553 11989 3587
rect 11989 3553 12023 3587
rect 12023 3553 12032 3587
rect 11980 3544 12032 3553
rect 13912 3612 13964 3664
rect 9128 3408 9180 3460
rect 13084 3476 13136 3528
rect 14280 3476 14332 3528
rect 14372 3519 14424 3528
rect 14372 3485 14381 3519
rect 14381 3485 14415 3519
rect 14415 3485 14424 3519
rect 14372 3476 14424 3485
rect 15660 3680 15712 3732
rect 14924 3587 14976 3596
rect 14924 3553 14933 3587
rect 14933 3553 14967 3587
rect 14967 3553 14976 3587
rect 14924 3544 14976 3553
rect 11152 3408 11204 3460
rect 11520 3451 11572 3460
rect 11520 3417 11545 3451
rect 11545 3417 11572 3451
rect 11520 3408 11572 3417
rect 12440 3408 12492 3460
rect 13912 3408 13964 3460
rect 15568 3476 15620 3528
rect 15844 3408 15896 3460
rect 8760 3340 8812 3392
rect 14096 3383 14148 3392
rect 14096 3349 14105 3383
rect 14105 3349 14139 3383
rect 14139 3349 14148 3383
rect 14096 3340 14148 3349
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 9220 3136 9272 3188
rect 10416 3179 10468 3188
rect 10416 3145 10425 3179
rect 10425 3145 10459 3179
rect 10459 3145 10468 3179
rect 10416 3136 10468 3145
rect 11244 3136 11296 3188
rect 13912 3136 13964 3188
rect 14556 3136 14608 3188
rect 15936 3136 15988 3188
rect 8944 3068 8996 3120
rect 11980 3068 12032 3120
rect 5540 3000 5592 3052
rect 13820 3068 13872 3120
rect 14740 3068 14792 3120
rect 15292 3068 15344 3120
rect 14096 3000 14148 3052
rect 14188 3043 14240 3052
rect 14188 3009 14197 3043
rect 14197 3009 14231 3043
rect 14231 3009 14240 3043
rect 14188 3000 14240 3009
rect 14280 3000 14332 3052
rect 14556 3000 14608 3052
rect 14924 3043 14976 3052
rect 14924 3009 14933 3043
rect 14933 3009 14967 3043
rect 14967 3009 14976 3043
rect 14924 3000 14976 3009
rect 10876 2975 10928 2984
rect 10876 2941 10885 2975
rect 10885 2941 10919 2975
rect 10919 2941 10928 2975
rect 10876 2932 10928 2941
rect 10968 2975 11020 2984
rect 10968 2941 10977 2975
rect 10977 2941 11011 2975
rect 11011 2941 11020 2975
rect 10968 2932 11020 2941
rect 13820 2864 13872 2916
rect 14464 2864 14516 2916
rect 14648 2796 14700 2848
rect 14740 2796 14792 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 14832 2635 14884 2644
rect 14832 2601 14841 2635
rect 14841 2601 14875 2635
rect 14875 2601 14884 2635
rect 14832 2592 14884 2601
rect 15200 2635 15252 2644
rect 15200 2601 15209 2635
rect 15209 2601 15243 2635
rect 15243 2601 15252 2635
rect 15200 2592 15252 2601
rect 16028 2592 16080 2644
rect 16212 2635 16264 2644
rect 16212 2601 16221 2635
rect 16221 2601 16255 2635
rect 16255 2601 16264 2635
rect 16212 2592 16264 2601
rect 8852 2524 8904 2576
rect 10876 2524 10928 2576
rect 14556 2524 14608 2576
rect 9312 2456 9364 2508
rect 7104 2388 7156 2440
rect 8760 2431 8812 2440
rect 8760 2397 8769 2431
rect 8769 2397 8803 2431
rect 8803 2397 8812 2431
rect 8760 2388 8812 2397
rect 9220 2388 9272 2440
rect 13820 2388 13872 2440
rect 13912 2431 13964 2440
rect 13912 2397 13921 2431
rect 13921 2397 13955 2431
rect 13955 2397 13964 2431
rect 13912 2388 13964 2397
rect 14004 2388 14056 2440
rect 14648 2431 14700 2440
rect 14648 2397 14657 2431
rect 14657 2397 14691 2431
rect 14691 2397 14700 2431
rect 14648 2388 14700 2397
rect 14740 2388 14792 2440
rect 15660 2388 15712 2440
rect 7748 2320 7800 2372
rect 9680 2320 9732 2372
rect 8392 2252 8444 2304
rect 9036 2252 9088 2304
rect 12900 2252 12952 2304
rect 13544 2252 13596 2304
rect 14188 2252 14240 2304
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
<< metal2 >>
rect 7746 34714 7802 35514
rect 12898 34714 12954 35514
rect 13542 34714 13598 35514
rect 14830 34714 14886 35514
rect 15474 34714 15530 35514
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 7760 33114 7788 34714
rect 12912 33114 12940 34714
rect 7748 33108 7800 33114
rect 7748 33050 7800 33056
rect 12900 33108 12952 33114
rect 12900 33050 12952 33056
rect 12992 33108 13044 33114
rect 12992 33050 13044 33056
rect 8116 32904 8168 32910
rect 8116 32846 8168 32852
rect 10600 32904 10652 32910
rect 10600 32846 10652 32852
rect 10876 32904 10928 32910
rect 10876 32846 10928 32852
rect 11336 32904 11388 32910
rect 11336 32846 11388 32852
rect 11520 32904 11572 32910
rect 11520 32846 11572 32852
rect 12806 32872 12862 32881
rect 4874 32668 5182 32677
rect 4874 32666 4880 32668
rect 4936 32666 4960 32668
rect 5016 32666 5040 32668
rect 5096 32666 5120 32668
rect 5176 32666 5182 32668
rect 4936 32614 4938 32666
rect 5118 32614 5120 32666
rect 4874 32612 4880 32614
rect 4936 32612 4960 32614
rect 5016 32612 5040 32614
rect 5096 32612 5120 32614
rect 5176 32612 5182 32614
rect 4874 32603 5182 32612
rect 7196 32428 7248 32434
rect 7196 32370 7248 32376
rect 7380 32428 7432 32434
rect 7380 32370 7432 32376
rect 7472 32428 7524 32434
rect 7472 32370 7524 32376
rect 7012 32292 7064 32298
rect 7012 32234 7064 32240
rect 7104 32292 7156 32298
rect 7104 32234 7156 32240
rect 6736 32224 6788 32230
rect 6736 32166 6788 32172
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 6748 31754 6776 32166
rect 7024 31929 7052 32234
rect 7010 31920 7066 31929
rect 7010 31855 7066 31864
rect 6736 31748 6788 31754
rect 6736 31690 6788 31696
rect 6920 31748 6972 31754
rect 6920 31690 6972 31696
rect 4874 31580 5182 31589
rect 4874 31578 4880 31580
rect 4936 31578 4960 31580
rect 5016 31578 5040 31580
rect 5096 31578 5120 31580
rect 5176 31578 5182 31580
rect 4936 31526 4938 31578
rect 5118 31526 5120 31578
rect 4874 31524 4880 31526
rect 4936 31524 4960 31526
rect 5016 31524 5040 31526
rect 5096 31524 5120 31526
rect 5176 31524 5182 31526
rect 4874 31515 5182 31524
rect 6092 31272 6144 31278
rect 6092 31214 6144 31220
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 6104 30938 6132 31214
rect 6932 31210 6960 31690
rect 7116 31346 7144 32234
rect 7208 31793 7236 32370
rect 7194 31784 7250 31793
rect 7194 31719 7250 31728
rect 7392 31482 7420 32370
rect 7380 31476 7432 31482
rect 7380 31418 7432 31424
rect 7104 31340 7156 31346
rect 7104 31282 7156 31288
rect 6920 31204 6972 31210
rect 6920 31146 6972 31152
rect 6736 31136 6788 31142
rect 6736 31078 6788 31084
rect 6092 30932 6144 30938
rect 6092 30874 6144 30880
rect 4874 30492 5182 30501
rect 4874 30490 4880 30492
rect 4936 30490 4960 30492
rect 5016 30490 5040 30492
rect 5096 30490 5120 30492
rect 5176 30490 5182 30492
rect 4936 30438 4938 30490
rect 5118 30438 5120 30490
rect 4874 30436 4880 30438
rect 4936 30436 4960 30438
rect 5016 30436 5040 30438
rect 5096 30436 5120 30438
rect 5176 30436 5182 30438
rect 4874 30427 5182 30436
rect 5908 30252 5960 30258
rect 5908 30194 5960 30200
rect 110 30152 166 30161
rect 110 30087 166 30096
rect 124 17746 152 30087
rect 5540 30048 5592 30054
rect 5540 29990 5592 29996
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4874 29404 5182 29413
rect 4874 29402 4880 29404
rect 4936 29402 4960 29404
rect 5016 29402 5040 29404
rect 5096 29402 5120 29404
rect 5176 29402 5182 29404
rect 4936 29350 4938 29402
rect 5118 29350 5120 29402
rect 4874 29348 4880 29350
rect 4936 29348 4960 29350
rect 5016 29348 5040 29350
rect 5096 29348 5120 29350
rect 5176 29348 5182 29350
rect 4874 29339 5182 29348
rect 5552 29170 5580 29990
rect 5724 29504 5776 29510
rect 5724 29446 5776 29452
rect 5540 29164 5592 29170
rect 5540 29106 5592 29112
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 5736 28558 5764 29446
rect 5920 29238 5948 30194
rect 6104 30190 6132 30874
rect 6460 30728 6512 30734
rect 6460 30670 6512 30676
rect 6472 30326 6500 30670
rect 6748 30394 6776 31078
rect 6932 30734 6960 31146
rect 7484 30818 7512 32370
rect 7656 32360 7708 32366
rect 7656 32302 7708 32308
rect 7564 31340 7616 31346
rect 7564 31282 7616 31288
rect 7392 30790 7512 30818
rect 6920 30728 6972 30734
rect 6920 30670 6972 30676
rect 7012 30660 7064 30666
rect 7012 30602 7064 30608
rect 6736 30388 6788 30394
rect 6736 30330 6788 30336
rect 6828 30388 6880 30394
rect 6828 30330 6880 30336
rect 6460 30320 6512 30326
rect 6460 30262 6512 30268
rect 6184 30252 6236 30258
rect 6184 30194 6236 30200
rect 6092 30184 6144 30190
rect 6092 30126 6144 30132
rect 6104 29850 6132 30126
rect 6092 29844 6144 29850
rect 6092 29786 6144 29792
rect 6104 29510 6132 29786
rect 6196 29646 6224 30194
rect 6184 29640 6236 29646
rect 6840 29594 6868 30330
rect 7024 30054 7052 30602
rect 7012 30048 7064 30054
rect 7012 29990 7064 29996
rect 7392 29850 7420 30790
rect 7472 30728 7524 30734
rect 7472 30670 7524 30676
rect 7484 30258 7512 30670
rect 7472 30252 7524 30258
rect 7472 30194 7524 30200
rect 7576 30138 7604 31282
rect 7668 31278 7696 32302
rect 8128 32026 8156 32846
rect 10416 32768 10468 32774
rect 10416 32710 10468 32716
rect 9128 32428 9180 32434
rect 9128 32370 9180 32376
rect 8392 32224 8444 32230
rect 8392 32166 8444 32172
rect 8116 32020 8168 32026
rect 8116 31962 8168 31968
rect 8128 31822 8156 31962
rect 8404 31890 8432 32166
rect 9140 32026 9168 32370
rect 9128 32020 9180 32026
rect 9128 31962 9180 31968
rect 8392 31884 8444 31890
rect 8392 31826 8444 31832
rect 8116 31816 8168 31822
rect 8484 31816 8536 31822
rect 8116 31758 8168 31764
rect 8404 31764 8484 31770
rect 8404 31758 8536 31764
rect 9404 31816 9456 31822
rect 9404 31758 9456 31764
rect 9680 31816 9732 31822
rect 9680 31758 9732 31764
rect 8404 31742 8524 31758
rect 8852 31748 8904 31754
rect 7932 31680 7984 31686
rect 7932 31622 7984 31628
rect 7944 31414 7972 31622
rect 7932 31408 7984 31414
rect 7932 31350 7984 31356
rect 7656 31272 7708 31278
rect 7656 31214 7708 31220
rect 8024 31272 8076 31278
rect 8024 31214 8076 31220
rect 7484 30110 7604 30138
rect 7104 29844 7156 29850
rect 7104 29786 7156 29792
rect 7380 29844 7432 29850
rect 7380 29786 7432 29792
rect 6918 29744 6974 29753
rect 6918 29679 6974 29688
rect 6932 29646 6960 29679
rect 6184 29582 6236 29588
rect 6656 29566 6868 29594
rect 6920 29640 6972 29646
rect 6920 29582 6972 29588
rect 7116 29578 7144 29786
rect 7196 29776 7248 29782
rect 7196 29718 7248 29724
rect 7286 29744 7342 29753
rect 7104 29572 7156 29578
rect 6092 29504 6144 29510
rect 6092 29446 6144 29452
rect 6656 29306 6684 29566
rect 7104 29514 7156 29520
rect 6736 29504 6788 29510
rect 6736 29446 6788 29452
rect 6920 29504 6972 29510
rect 6920 29446 6972 29452
rect 6748 29306 6776 29446
rect 6644 29300 6696 29306
rect 6644 29242 6696 29248
rect 6736 29300 6788 29306
rect 6736 29242 6788 29248
rect 5908 29232 5960 29238
rect 5908 29174 5960 29180
rect 6828 29232 6880 29238
rect 6828 29174 6880 29180
rect 6644 29164 6696 29170
rect 6644 29106 6696 29112
rect 6656 28642 6684 29106
rect 6840 28762 6868 29174
rect 6932 29170 6960 29446
rect 6920 29164 6972 29170
rect 6920 29106 6972 29112
rect 7208 29034 7236 29718
rect 7286 29679 7342 29688
rect 7300 29034 7328 29679
rect 7196 29028 7248 29034
rect 7196 28970 7248 28976
rect 7288 29028 7340 29034
rect 7288 28970 7340 28976
rect 6828 28756 6880 28762
rect 6828 28698 6880 28704
rect 6656 28614 6868 28642
rect 6840 28558 6868 28614
rect 7208 28558 7236 28970
rect 5724 28552 5776 28558
rect 5724 28494 5776 28500
rect 6828 28552 6880 28558
rect 6828 28494 6880 28500
rect 7196 28552 7248 28558
rect 7196 28494 7248 28500
rect 2964 28484 3016 28490
rect 2964 28426 3016 28432
rect 2596 28076 2648 28082
rect 2596 28018 2648 28024
rect 2412 27396 2464 27402
rect 2412 27338 2464 27344
rect 2136 27124 2188 27130
rect 2136 27066 2188 27072
rect 1676 26988 1728 26994
rect 1676 26930 1728 26936
rect 1688 26518 1716 26930
rect 2044 26920 2096 26926
rect 2044 26862 2096 26868
rect 1676 26512 1728 26518
rect 1676 26454 1728 26460
rect 846 25392 902 25401
rect 846 25327 902 25336
rect 860 25294 888 25327
rect 848 25288 900 25294
rect 848 25230 900 25236
rect 2056 24954 2084 26862
rect 2044 24948 2096 24954
rect 2044 24890 2096 24896
rect 1860 24744 1912 24750
rect 1860 24686 1912 24692
rect 1768 24608 1820 24614
rect 1768 24550 1820 24556
rect 1780 24206 1808 24550
rect 1872 24410 1900 24686
rect 1860 24404 1912 24410
rect 1860 24346 1912 24352
rect 1400 24200 1452 24206
rect 1400 24142 1452 24148
rect 1768 24200 1820 24206
rect 1768 24142 1820 24148
rect 2044 24200 2096 24206
rect 2044 24142 2096 24148
rect 1412 23730 1440 24142
rect 1400 23724 1452 23730
rect 1400 23666 1452 23672
rect 1676 23724 1728 23730
rect 1676 23666 1728 23672
rect 1688 23322 1716 23666
rect 1676 23316 1728 23322
rect 1676 23258 1728 23264
rect 2056 23186 2084 24142
rect 2044 23180 2096 23186
rect 2044 23122 2096 23128
rect 848 21548 900 21554
rect 848 21490 900 21496
rect 860 21321 888 21490
rect 846 21312 902 21321
rect 846 21247 902 21256
rect 2056 21078 2084 23122
rect 2148 23118 2176 27066
rect 2320 27056 2372 27062
rect 2320 26998 2372 27004
rect 2228 26920 2280 26926
rect 2228 26862 2280 26868
rect 2240 26586 2268 26862
rect 2228 26580 2280 26586
rect 2332 26568 2360 26998
rect 2424 26858 2452 27338
rect 2412 26852 2464 26858
rect 2412 26794 2464 26800
rect 2608 26586 2636 28018
rect 2780 28008 2832 28014
rect 2780 27950 2832 27956
rect 2792 27470 2820 27950
rect 2780 27464 2832 27470
rect 2780 27406 2832 27412
rect 2872 27124 2924 27130
rect 2872 27066 2924 27072
rect 2780 27056 2832 27062
rect 2778 27024 2780 27033
rect 2832 27024 2834 27033
rect 2700 26982 2778 27010
rect 2596 26580 2648 26586
rect 2332 26540 2544 26568
rect 2228 26522 2280 26528
rect 2516 26450 2544 26540
rect 2596 26522 2648 26528
rect 2594 26480 2650 26489
rect 2412 26444 2464 26450
rect 2412 26386 2464 26392
rect 2504 26444 2556 26450
rect 2594 26415 2650 26424
rect 2504 26386 2556 26392
rect 2424 25974 2452 26386
rect 2412 25968 2464 25974
rect 2412 25910 2464 25916
rect 2608 24750 2636 26415
rect 2596 24744 2648 24750
rect 2596 24686 2648 24692
rect 2596 24132 2648 24138
rect 2596 24074 2648 24080
rect 2608 23322 2636 24074
rect 2596 23316 2648 23322
rect 2596 23258 2648 23264
rect 2700 23254 2728 26982
rect 2778 26959 2834 26968
rect 2884 26897 2912 27066
rect 2976 26926 3004 28426
rect 4874 28316 5182 28325
rect 4874 28314 4880 28316
rect 4936 28314 4960 28316
rect 5016 28314 5040 28316
rect 5096 28314 5120 28316
rect 5176 28314 5182 28316
rect 4936 28262 4938 28314
rect 5118 28262 5120 28314
rect 4874 28260 4880 28262
rect 4936 28260 4960 28262
rect 5016 28260 5040 28262
rect 5096 28260 5120 28262
rect 5176 28260 5182 28262
rect 4874 28251 5182 28260
rect 3424 28076 3476 28082
rect 3424 28018 3476 28024
rect 4712 28076 4764 28082
rect 4712 28018 4764 28024
rect 6736 28076 6788 28082
rect 6736 28018 6788 28024
rect 3332 27328 3384 27334
rect 3332 27270 3384 27276
rect 2964 26920 3016 26926
rect 2870 26888 2926 26897
rect 3344 26908 3372 27270
rect 2964 26862 3016 26868
rect 3252 26880 3372 26908
rect 2870 26823 2926 26832
rect 2780 26580 2832 26586
rect 2780 26522 2832 26528
rect 2792 26489 2820 26522
rect 2778 26480 2834 26489
rect 2778 26415 2834 26424
rect 2976 26364 3004 26862
rect 3056 26852 3108 26858
rect 3056 26794 3108 26800
rect 3068 26761 3096 26794
rect 3054 26752 3110 26761
rect 3054 26687 3110 26696
rect 3148 26376 3200 26382
rect 2976 26336 3148 26364
rect 2872 26240 2924 26246
rect 2872 26182 2924 26188
rect 2884 24818 2912 26182
rect 2872 24812 2924 24818
rect 2872 24754 2924 24760
rect 3068 24274 3096 26336
rect 3148 26318 3200 26324
rect 3252 26246 3280 26880
rect 3436 26790 3464 28018
rect 3792 27940 3844 27946
rect 3792 27882 3844 27888
rect 3804 27470 3832 27882
rect 3976 27872 4028 27878
rect 3976 27814 4028 27820
rect 3792 27464 3844 27470
rect 3792 27406 3844 27412
rect 3884 27328 3936 27334
rect 3884 27270 3936 27276
rect 3896 27130 3924 27270
rect 3884 27124 3936 27130
rect 3884 27066 3936 27072
rect 3516 26988 3568 26994
rect 3516 26930 3568 26936
rect 3424 26784 3476 26790
rect 3528 26761 3556 26930
rect 3424 26726 3476 26732
rect 3514 26752 3570 26761
rect 3332 26376 3384 26382
rect 3332 26318 3384 26324
rect 3240 26240 3292 26246
rect 3240 26182 3292 26188
rect 3148 25968 3200 25974
rect 3148 25910 3200 25916
rect 3056 24268 3108 24274
rect 3056 24210 3108 24216
rect 3160 24206 3188 25910
rect 3252 25702 3280 26182
rect 3344 25974 3372 26318
rect 3332 25968 3384 25974
rect 3332 25910 3384 25916
rect 3436 25770 3464 26726
rect 3514 26687 3570 26696
rect 3792 26580 3844 26586
rect 3792 26522 3844 26528
rect 3804 26314 3832 26522
rect 3884 26376 3936 26382
rect 3988 26364 4016 27814
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4160 27464 4212 27470
rect 4160 27406 4212 27412
rect 4068 27396 4120 27402
rect 4068 27338 4120 27344
rect 3936 26336 4016 26364
rect 3884 26318 3936 26324
rect 3516 26308 3568 26314
rect 3516 26250 3568 26256
rect 3792 26308 3844 26314
rect 3792 26250 3844 26256
rect 3424 25764 3476 25770
rect 3424 25706 3476 25712
rect 3240 25696 3292 25702
rect 3528 25650 3556 26250
rect 3988 26042 4016 26336
rect 3976 26036 4028 26042
rect 3976 25978 4028 25984
rect 3240 25638 3292 25644
rect 2964 24200 3016 24206
rect 2964 24142 3016 24148
rect 3148 24200 3200 24206
rect 3148 24142 3200 24148
rect 2976 23866 3004 24142
rect 3056 24064 3108 24070
rect 3056 24006 3108 24012
rect 3148 24064 3200 24070
rect 3252 24052 3280 25638
rect 3436 25622 3556 25650
rect 3436 24818 3464 25622
rect 3516 25152 3568 25158
rect 3516 25094 3568 25100
rect 3528 24818 3556 25094
rect 3608 24880 3660 24886
rect 3608 24822 3660 24828
rect 3424 24812 3476 24818
rect 3424 24754 3476 24760
rect 3516 24812 3568 24818
rect 3516 24754 3568 24760
rect 3436 24698 3464 24754
rect 3436 24670 3556 24698
rect 3424 24608 3476 24614
rect 3424 24550 3476 24556
rect 3436 24206 3464 24550
rect 3424 24200 3476 24206
rect 3422 24168 3424 24177
rect 3476 24168 3478 24177
rect 3332 24132 3384 24138
rect 3422 24103 3478 24112
rect 3332 24074 3384 24080
rect 3200 24024 3280 24052
rect 3148 24006 3200 24012
rect 2964 23860 3016 23866
rect 2964 23802 3016 23808
rect 3068 23730 3096 24006
rect 3160 23730 3188 24006
rect 3344 23730 3372 24074
rect 2872 23724 2924 23730
rect 2872 23666 2924 23672
rect 3056 23724 3108 23730
rect 3056 23666 3108 23672
rect 3148 23724 3200 23730
rect 3148 23666 3200 23672
rect 3332 23724 3384 23730
rect 3332 23666 3384 23672
rect 3424 23724 3476 23730
rect 3424 23666 3476 23672
rect 2688 23248 2740 23254
rect 2740 23208 2820 23236
rect 2688 23190 2740 23196
rect 2136 23112 2188 23118
rect 2136 23054 2188 23060
rect 2320 23112 2372 23118
rect 2320 23054 2372 23060
rect 2044 21072 2096 21078
rect 2044 21014 2096 21020
rect 2148 21010 2176 23054
rect 2228 22772 2280 22778
rect 2228 22714 2280 22720
rect 2136 21004 2188 21010
rect 2136 20946 2188 20952
rect 2240 20913 2268 22714
rect 2332 22506 2360 23054
rect 2504 22976 2556 22982
rect 2504 22918 2556 22924
rect 2516 22778 2544 22918
rect 2504 22772 2556 22778
rect 2504 22714 2556 22720
rect 2412 22568 2464 22574
rect 2412 22510 2464 22516
rect 2320 22500 2372 22506
rect 2320 22442 2372 22448
rect 2424 22094 2452 22510
rect 2332 22066 2452 22094
rect 2226 20904 2282 20913
rect 2226 20839 2228 20848
rect 2280 20839 2282 20848
rect 2228 20810 2280 20816
rect 1492 20800 1544 20806
rect 1492 20742 1544 20748
rect 1400 20392 1452 20398
rect 1400 20334 1452 20340
rect 1412 20058 1440 20334
rect 1400 20052 1452 20058
rect 1400 19994 1452 20000
rect 1412 19922 1440 19994
rect 1400 19916 1452 19922
rect 1400 19858 1452 19864
rect 1504 19854 1532 20742
rect 1492 19848 1544 19854
rect 1492 19790 1544 19796
rect 2332 19174 2360 22066
rect 2792 21010 2820 23208
rect 2884 23118 2912 23666
rect 2964 23520 3016 23526
rect 2964 23462 3016 23468
rect 2976 23322 3004 23462
rect 2964 23316 3016 23322
rect 2964 23258 3016 23264
rect 2976 23118 3004 23258
rect 3068 23254 3096 23666
rect 3056 23248 3108 23254
rect 3056 23190 3108 23196
rect 3332 23180 3384 23186
rect 3332 23122 3384 23128
rect 2872 23112 2924 23118
rect 2872 23054 2924 23060
rect 2964 23112 3016 23118
rect 2964 23054 3016 23060
rect 3240 23112 3292 23118
rect 3240 23054 3292 23060
rect 2884 22778 2912 23054
rect 2976 22930 3004 23054
rect 3056 23044 3108 23050
rect 3108 23004 3188 23032
rect 3056 22986 3108 22992
rect 2976 22902 3096 22930
rect 2872 22772 2924 22778
rect 2872 22714 2924 22720
rect 3068 22642 3096 22902
rect 3056 22636 3108 22642
rect 3056 22578 3108 22584
rect 3160 22438 3188 23004
rect 3252 22574 3280 23054
rect 3240 22568 3292 22574
rect 3240 22510 3292 22516
rect 3148 22432 3200 22438
rect 3148 22374 3200 22380
rect 3160 21554 3188 22374
rect 3344 22234 3372 23122
rect 3332 22228 3384 22234
rect 3332 22170 3384 22176
rect 3332 22094 3384 22098
rect 3436 22094 3464 23666
rect 3528 22778 3556 24670
rect 3620 24206 3648 24822
rect 3988 24818 4016 25978
rect 4080 25770 4108 27338
rect 4172 27062 4200 27406
rect 4620 27396 4672 27402
rect 4620 27338 4672 27344
rect 4160 27056 4212 27062
rect 4160 26998 4212 27004
rect 4172 26790 4200 26998
rect 4160 26784 4212 26790
rect 4160 26726 4212 26732
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4632 26518 4660 27338
rect 4724 27130 4752 28018
rect 5816 27940 5868 27946
rect 5816 27882 5868 27888
rect 5632 27464 5684 27470
rect 5632 27406 5684 27412
rect 5264 27328 5316 27334
rect 5264 27270 5316 27276
rect 4874 27228 5182 27237
rect 4874 27226 4880 27228
rect 4936 27226 4960 27228
rect 5016 27226 5040 27228
rect 5096 27226 5120 27228
rect 5176 27226 5182 27228
rect 4936 27174 4938 27226
rect 5118 27174 5120 27226
rect 4874 27172 4880 27174
rect 4936 27172 4960 27174
rect 5016 27172 5040 27174
rect 5096 27172 5120 27174
rect 5176 27172 5182 27174
rect 4874 27163 5182 27172
rect 4712 27124 4764 27130
rect 4712 27066 4764 27072
rect 4620 26512 4672 26518
rect 4620 26454 4672 26460
rect 4252 26444 4304 26450
rect 4252 26386 4304 26392
rect 4264 26246 4292 26386
rect 4436 26308 4488 26314
rect 4436 26250 4488 26256
rect 4252 26240 4304 26246
rect 4252 26182 4304 26188
rect 4448 25838 4476 26250
rect 4620 26240 4672 26246
rect 4620 26182 4672 26188
rect 4436 25832 4488 25838
rect 4436 25774 4488 25780
rect 4068 25764 4120 25770
rect 4068 25706 4120 25712
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4632 25362 4660 26182
rect 4724 25974 4752 27066
rect 4802 27024 4858 27033
rect 4802 26959 4858 26968
rect 4988 26988 5040 26994
rect 4816 26450 4844 26959
rect 4988 26930 5040 26936
rect 4804 26444 4856 26450
rect 4804 26386 4856 26392
rect 4804 26308 4856 26314
rect 4804 26250 4856 26256
rect 4712 25968 4764 25974
rect 4712 25910 4764 25916
rect 4620 25356 4672 25362
rect 4620 25298 4672 25304
rect 4632 24954 4660 25298
rect 4620 24948 4672 24954
rect 4620 24890 4672 24896
rect 4724 24886 4752 25910
rect 4816 25906 4844 26250
rect 5000 26246 5028 26930
rect 5078 26888 5134 26897
rect 5078 26823 5134 26832
rect 5092 26450 5120 26823
rect 5080 26444 5132 26450
rect 5080 26386 5132 26392
rect 4988 26240 5040 26246
rect 5092 26228 5120 26386
rect 5276 26314 5304 27270
rect 5644 26790 5672 27406
rect 5632 26784 5684 26790
rect 5632 26726 5684 26732
rect 5540 26444 5592 26450
rect 5540 26386 5592 26392
rect 5356 26376 5408 26382
rect 5356 26318 5408 26324
rect 5264 26308 5316 26314
rect 5264 26250 5316 26256
rect 5092 26200 5237 26228
rect 4988 26182 5040 26188
rect 5209 26194 5237 26200
rect 5209 26166 5304 26194
rect 4874 26140 5182 26149
rect 4874 26138 4880 26140
rect 4936 26138 4960 26140
rect 5016 26138 5040 26140
rect 5096 26138 5120 26140
rect 5176 26138 5182 26140
rect 4936 26086 4938 26138
rect 5118 26086 5120 26138
rect 4874 26084 4880 26086
rect 4936 26084 4960 26086
rect 5016 26084 5040 26086
rect 5096 26084 5120 26086
rect 5176 26084 5182 26086
rect 4874 26075 5182 26084
rect 4804 25900 4856 25906
rect 4804 25842 4856 25848
rect 4816 25702 4844 25842
rect 4804 25696 4856 25702
rect 4804 25638 4856 25644
rect 4816 24936 4844 25638
rect 4874 25052 5182 25061
rect 4874 25050 4880 25052
rect 4936 25050 4960 25052
rect 5016 25050 5040 25052
rect 5096 25050 5120 25052
rect 5176 25050 5182 25052
rect 4936 24998 4938 25050
rect 5118 24998 5120 25050
rect 4874 24996 4880 24998
rect 4936 24996 4960 24998
rect 5016 24996 5040 24998
rect 5096 24996 5120 24998
rect 5176 24996 5182 24998
rect 4874 24987 5182 24996
rect 4816 24908 4936 24936
rect 4712 24880 4764 24886
rect 4712 24822 4764 24828
rect 3976 24812 4028 24818
rect 3976 24754 4028 24760
rect 3884 24744 3936 24750
rect 3884 24686 3936 24692
rect 4724 24698 4752 24822
rect 4908 24750 4936 24908
rect 4896 24744 4948 24750
rect 3792 24676 3844 24682
rect 3792 24618 3844 24624
rect 3608 24200 3660 24206
rect 3608 24142 3660 24148
rect 3700 23724 3752 23730
rect 3804 23712 3832 24618
rect 3896 24154 3924 24686
rect 4620 24676 4672 24682
rect 4724 24670 4844 24698
rect 4896 24686 4948 24692
rect 4620 24618 4672 24624
rect 4068 24608 4120 24614
rect 4068 24550 4120 24556
rect 3976 24336 4028 24342
rect 3974 24304 3976 24313
rect 4028 24304 4030 24313
rect 3974 24239 4030 24248
rect 4080 24206 4108 24550
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4252 24404 4304 24410
rect 4252 24346 4304 24352
rect 4068 24200 4120 24206
rect 3896 24126 4016 24154
rect 4068 24142 4120 24148
rect 3988 24018 4016 24126
rect 4068 24064 4120 24070
rect 3988 24012 4068 24018
rect 3988 24006 4120 24012
rect 3988 23990 4108 24006
rect 3752 23684 3832 23712
rect 3700 23666 3752 23672
rect 3608 23656 3660 23662
rect 3608 23598 3660 23604
rect 3516 22772 3568 22778
rect 3516 22714 3568 22720
rect 3332 22092 3464 22094
rect 3252 22052 3332 22080
rect 3148 21548 3200 21554
rect 3148 21490 3200 21496
rect 2780 21004 2832 21010
rect 2608 20964 2780 20992
rect 2412 20936 2464 20942
rect 2608 20924 2636 20964
rect 2780 20946 2832 20952
rect 2464 20896 2636 20924
rect 2872 20936 2924 20942
rect 2870 20904 2872 20913
rect 2924 20904 2926 20913
rect 2412 20878 2464 20884
rect 2870 20839 2926 20848
rect 2964 20868 3016 20874
rect 2412 20800 2464 20806
rect 2412 20742 2464 20748
rect 2424 20534 2452 20742
rect 2412 20528 2464 20534
rect 2412 20470 2464 20476
rect 2884 20466 2912 20839
rect 2964 20810 3016 20816
rect 2872 20460 2924 20466
rect 2872 20402 2924 20408
rect 2884 19990 2912 20402
rect 2976 20398 3004 20810
rect 3160 20602 3188 21490
rect 3148 20596 3200 20602
rect 3148 20538 3200 20544
rect 3160 20466 3188 20538
rect 3148 20460 3200 20466
rect 3148 20402 3200 20408
rect 2964 20392 3016 20398
rect 2964 20334 3016 20340
rect 2872 19984 2924 19990
rect 2872 19926 2924 19932
rect 2320 19168 2372 19174
rect 2320 19110 2372 19116
rect 2688 19168 2740 19174
rect 2688 19110 2740 19116
rect 3148 19168 3200 19174
rect 3252 19156 3280 22052
rect 3384 22066 3464 22092
rect 3332 22034 3384 22040
rect 3620 21690 3648 23598
rect 3608 21684 3660 21690
rect 3608 21626 3660 21632
rect 3332 21548 3384 21554
rect 3332 21490 3384 21496
rect 3344 21146 3372 21490
rect 3424 21344 3476 21350
rect 3424 21286 3476 21292
rect 3332 21140 3384 21146
rect 3332 21082 3384 21088
rect 3436 20942 3464 21286
rect 3424 20936 3476 20942
rect 3424 20878 3476 20884
rect 3436 19718 3464 20878
rect 3620 20618 3648 21626
rect 3712 20754 3740 23666
rect 4080 23662 4108 23990
rect 4264 23730 4292 24346
rect 4252 23724 4304 23730
rect 4252 23666 4304 23672
rect 4068 23656 4120 23662
rect 4068 23598 4120 23604
rect 3792 23520 3844 23526
rect 3792 23462 3844 23468
rect 4068 23520 4120 23526
rect 4068 23462 4120 23468
rect 3804 23118 3832 23462
rect 3792 23112 3844 23118
rect 3792 23054 3844 23060
rect 4080 23100 4108 23462
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4160 23112 4212 23118
rect 4080 23072 4160 23100
rect 3792 22772 3844 22778
rect 3792 22714 3844 22720
rect 3804 21146 3832 22714
rect 4080 22642 4108 23072
rect 4632 23066 4660 24618
rect 4712 24608 4764 24614
rect 4712 24550 4764 24556
rect 4160 23054 4212 23060
rect 4252 23044 4304 23050
rect 4252 22986 4304 22992
rect 4448 23038 4660 23066
rect 4068 22636 4120 22642
rect 4068 22578 4120 22584
rect 4264 22506 4292 22986
rect 4448 22642 4476 23038
rect 4724 22982 4752 24550
rect 4816 23594 4844 24670
rect 4908 24410 4936 24686
rect 4896 24404 4948 24410
rect 4896 24346 4948 24352
rect 4988 24268 5040 24274
rect 5276 24256 5304 26166
rect 5368 26042 5396 26318
rect 5552 26042 5580 26386
rect 5356 26036 5408 26042
rect 5356 25978 5408 25984
rect 5540 26036 5592 26042
rect 5540 25978 5592 25984
rect 5368 25838 5396 25978
rect 5356 25832 5408 25838
rect 5356 25774 5408 25780
rect 5368 24410 5396 25774
rect 5644 25226 5672 26726
rect 5828 26314 5856 27882
rect 6000 27396 6052 27402
rect 6000 27338 6052 27344
rect 5906 27024 5962 27033
rect 5906 26959 5962 26968
rect 5816 26308 5868 26314
rect 5816 26250 5868 26256
rect 5920 26246 5948 26959
rect 6012 26518 6040 27338
rect 6748 27334 6776 28018
rect 6276 27328 6328 27334
rect 6276 27270 6328 27276
rect 6736 27328 6788 27334
rect 6736 27270 6788 27276
rect 6092 26784 6144 26790
rect 6092 26726 6144 26732
rect 6000 26512 6052 26518
rect 6000 26454 6052 26460
rect 6000 26376 6052 26382
rect 6104 26364 6132 26726
rect 6288 26382 6316 27270
rect 6052 26336 6132 26364
rect 6000 26318 6052 26324
rect 5724 26240 5776 26246
rect 5724 26182 5776 26188
rect 5908 26240 5960 26246
rect 5908 26182 5960 26188
rect 5736 25906 5764 26182
rect 5724 25900 5776 25906
rect 5724 25842 5776 25848
rect 5816 25900 5868 25906
rect 5816 25842 5868 25848
rect 5828 25702 5856 25842
rect 5816 25696 5868 25702
rect 5816 25638 5868 25644
rect 5632 25220 5684 25226
rect 5632 25162 5684 25168
rect 5644 24818 5672 25162
rect 5828 24818 5856 25638
rect 5632 24812 5684 24818
rect 5632 24754 5684 24760
rect 5816 24812 5868 24818
rect 5816 24754 5868 24760
rect 5448 24608 5500 24614
rect 5448 24550 5500 24556
rect 5356 24404 5408 24410
rect 5356 24346 5408 24352
rect 5460 24274 5488 24550
rect 5448 24268 5500 24274
rect 5040 24228 5396 24256
rect 4988 24210 5040 24216
rect 5368 24154 5396 24228
rect 5448 24210 5500 24216
rect 5172 24132 5224 24138
rect 5368 24126 5488 24154
rect 5224 24092 5304 24120
rect 5172 24074 5224 24080
rect 4874 23964 5182 23973
rect 4874 23962 4880 23964
rect 4936 23962 4960 23964
rect 5016 23962 5040 23964
rect 5096 23962 5120 23964
rect 5176 23962 5182 23964
rect 4936 23910 4938 23962
rect 5118 23910 5120 23962
rect 4874 23908 4880 23910
rect 4936 23908 4960 23910
rect 5016 23908 5040 23910
rect 5096 23908 5120 23910
rect 5176 23908 5182 23910
rect 4874 23899 5182 23908
rect 4804 23588 4856 23594
rect 4804 23530 4856 23536
rect 4620 22976 4672 22982
rect 4620 22918 4672 22924
rect 4712 22976 4764 22982
rect 4712 22918 4764 22924
rect 4804 22976 4856 22982
rect 4804 22918 4856 22924
rect 4436 22636 4488 22642
rect 4436 22578 4488 22584
rect 4252 22500 4304 22506
rect 4252 22442 4304 22448
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4436 22228 4488 22234
rect 4436 22170 4488 22176
rect 4344 22160 4396 22166
rect 4344 22102 4396 22108
rect 3976 22024 4028 22030
rect 3976 21966 4028 21972
rect 3884 21956 3936 21962
rect 3884 21898 3936 21904
rect 3896 21690 3924 21898
rect 3884 21684 3936 21690
rect 3884 21626 3936 21632
rect 3884 21548 3936 21554
rect 3884 21490 3936 21496
rect 3896 21350 3924 21490
rect 3884 21344 3936 21350
rect 3884 21286 3936 21292
rect 3792 21140 3844 21146
rect 3792 21082 3844 21088
rect 3712 20726 3832 20754
rect 3620 20590 3740 20618
rect 3608 20460 3660 20466
rect 3608 20402 3660 20408
rect 3620 20058 3648 20402
rect 3608 20052 3660 20058
rect 3608 19994 3660 20000
rect 3424 19712 3476 19718
rect 3424 19654 3476 19660
rect 3436 19514 3464 19654
rect 3424 19508 3476 19514
rect 3424 19450 3476 19456
rect 3712 19446 3740 20590
rect 3700 19440 3752 19446
rect 3700 19382 3752 19388
rect 3200 19128 3280 19156
rect 3148 19110 3200 19116
rect 2412 18284 2464 18290
rect 2464 18244 2544 18272
rect 2412 18226 2464 18232
rect 2136 18080 2188 18086
rect 2136 18022 2188 18028
rect 1952 17876 2004 17882
rect 1952 17818 2004 17824
rect 112 17740 164 17746
rect 112 17682 164 17688
rect 1768 17604 1820 17610
rect 1768 17546 1820 17552
rect 1400 17536 1452 17542
rect 1584 17536 1636 17542
rect 1452 17496 1532 17524
rect 1400 17478 1452 17484
rect 1400 17196 1452 17202
rect 1400 17138 1452 17144
rect 1412 16658 1440 17138
rect 1400 16652 1452 16658
rect 1400 16594 1452 16600
rect 1412 16114 1440 16594
rect 1504 16590 1532 17496
rect 1584 17478 1636 17484
rect 1492 16584 1544 16590
rect 1492 16526 1544 16532
rect 1400 16108 1452 16114
rect 1400 16050 1452 16056
rect 1596 15162 1624 17478
rect 1676 16108 1728 16114
rect 1676 16050 1728 16056
rect 1688 15706 1716 16050
rect 1780 15706 1808 17546
rect 1860 17536 1912 17542
rect 1860 17478 1912 17484
rect 1872 17202 1900 17478
rect 1860 17196 1912 17202
rect 1860 17138 1912 17144
rect 1676 15700 1728 15706
rect 1676 15642 1728 15648
rect 1768 15700 1820 15706
rect 1768 15642 1820 15648
rect 1964 15434 1992 17818
rect 2044 16108 2096 16114
rect 2044 16050 2096 16056
rect 1952 15428 2004 15434
rect 1872 15388 1952 15416
rect 1584 15156 1636 15162
rect 1584 15098 1636 15104
rect 1676 13252 1728 13258
rect 1676 13194 1728 13200
rect 1688 12986 1716 13194
rect 1676 12980 1728 12986
rect 1676 12922 1728 12928
rect 1872 12850 1900 15388
rect 1952 15370 2004 15376
rect 2056 15026 2084 16050
rect 2148 15026 2176 18022
rect 2412 17672 2464 17678
rect 2410 17640 2412 17649
rect 2464 17640 2466 17649
rect 2320 17604 2372 17610
rect 2410 17575 2466 17584
rect 2320 17546 2372 17552
rect 2332 16794 2360 17546
rect 2516 17542 2544 18244
rect 2700 17678 2728 19110
rect 3056 18284 3108 18290
rect 3056 18226 3108 18232
rect 2792 17882 2912 17898
rect 2792 17876 2924 17882
rect 2792 17870 2872 17876
rect 2688 17672 2740 17678
rect 2688 17614 2740 17620
rect 2412 17536 2464 17542
rect 2412 17478 2464 17484
rect 2504 17536 2556 17542
rect 2504 17478 2556 17484
rect 2320 16788 2372 16794
rect 2320 16730 2372 16736
rect 2044 15020 2096 15026
rect 2044 14962 2096 14968
rect 2136 15020 2188 15026
rect 2136 14962 2188 14968
rect 2056 13938 2084 14962
rect 2044 13932 2096 13938
rect 2044 13874 2096 13880
rect 1952 13728 2004 13734
rect 1952 13670 2004 13676
rect 1964 12986 1992 13670
rect 1952 12980 2004 12986
rect 1952 12922 2004 12928
rect 2056 12850 2084 13874
rect 1860 12844 1912 12850
rect 1860 12786 1912 12792
rect 2044 12844 2096 12850
rect 2044 12786 2096 12792
rect 1492 12164 1544 12170
rect 1492 12106 1544 12112
rect 1504 11898 1532 12106
rect 1768 12096 1820 12102
rect 1768 12038 1820 12044
rect 1492 11892 1544 11898
rect 1492 11834 1544 11840
rect 1780 11354 1808 12038
rect 1872 11830 1900 12786
rect 2332 12782 2360 16730
rect 2424 15162 2452 17478
rect 2412 15156 2464 15162
rect 2412 15098 2464 15104
rect 2516 15026 2544 17478
rect 2792 17082 2820 17870
rect 2872 17818 2924 17824
rect 2964 17808 3016 17814
rect 2964 17750 3016 17756
rect 2976 17338 3004 17750
rect 3068 17678 3096 18226
rect 3056 17672 3108 17678
rect 3056 17614 3108 17620
rect 2964 17332 3016 17338
rect 2964 17274 3016 17280
rect 2792 17054 2912 17082
rect 2884 16522 2912 17054
rect 2872 16516 2924 16522
rect 2872 16458 2924 16464
rect 2884 16130 2912 16458
rect 2976 16250 3004 17274
rect 3068 16454 3096 17614
rect 3160 17542 3188 19110
rect 3804 18358 3832 20726
rect 3896 20262 3924 21286
rect 3988 20534 4016 21966
rect 4356 21554 4384 22102
rect 4448 21554 4476 22170
rect 4632 22098 4660 22918
rect 4712 22636 4764 22642
rect 4712 22578 4764 22584
rect 4724 22506 4752 22578
rect 4712 22500 4764 22506
rect 4712 22442 4764 22448
rect 4620 22092 4672 22098
rect 4620 22034 4672 22040
rect 4724 21962 4752 22442
rect 4816 22030 4844 22918
rect 4874 22876 5182 22885
rect 4874 22874 4880 22876
rect 4936 22874 4960 22876
rect 5016 22874 5040 22876
rect 5096 22874 5120 22876
rect 5176 22874 5182 22876
rect 4936 22822 4938 22874
rect 5118 22822 5120 22874
rect 4874 22820 4880 22822
rect 4936 22820 4960 22822
rect 5016 22820 5040 22822
rect 5096 22820 5120 22822
rect 5176 22820 5182 22822
rect 4874 22811 5182 22820
rect 4988 22568 5040 22574
rect 4988 22510 5040 22516
rect 4896 22432 4948 22438
rect 4896 22374 4948 22380
rect 4804 22024 4856 22030
rect 4804 21966 4856 21972
rect 4712 21956 4764 21962
rect 4712 21898 4764 21904
rect 4620 21888 4672 21894
rect 4908 21876 4936 22374
rect 5000 22234 5028 22510
rect 5080 22500 5132 22506
rect 5080 22442 5132 22448
rect 4988 22228 5040 22234
rect 4988 22170 5040 22176
rect 5092 22166 5120 22442
rect 5080 22160 5132 22166
rect 5080 22102 5132 22108
rect 4620 21830 4672 21836
rect 4816 21848 4936 21876
rect 4344 21548 4396 21554
rect 4344 21490 4396 21496
rect 4436 21548 4488 21554
rect 4436 21490 4488 21496
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4344 20936 4396 20942
rect 4344 20878 4396 20884
rect 4528 20936 4580 20942
rect 4528 20878 4580 20884
rect 4158 20632 4214 20641
rect 4356 20602 4384 20878
rect 4158 20567 4214 20576
rect 4344 20596 4396 20602
rect 3976 20528 4028 20534
rect 3976 20470 4028 20476
rect 3884 20256 3936 20262
rect 3884 20198 3936 20204
rect 3988 19446 4016 20470
rect 4172 20466 4200 20567
rect 4344 20538 4396 20544
rect 4160 20460 4212 20466
rect 4160 20402 4212 20408
rect 4068 20392 4120 20398
rect 4068 20334 4120 20340
rect 4540 20346 4568 20878
rect 4632 20466 4660 21830
rect 4712 21344 4764 21350
rect 4712 21286 4764 21292
rect 4620 20460 4672 20466
rect 4620 20402 4672 20408
rect 4080 20040 4108 20334
rect 4540 20318 4660 20346
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4160 20052 4212 20058
rect 4080 20012 4160 20040
rect 4160 19994 4212 20000
rect 4344 20052 4396 20058
rect 4344 19994 4396 20000
rect 4528 20052 4580 20058
rect 4528 19994 4580 20000
rect 4252 19848 4304 19854
rect 4252 19790 4304 19796
rect 4160 19780 4212 19786
rect 4160 19722 4212 19728
rect 4172 19514 4200 19722
rect 4160 19508 4212 19514
rect 4160 19450 4212 19456
rect 3976 19440 4028 19446
rect 3976 19382 4028 19388
rect 4264 19378 4292 19790
rect 4356 19718 4384 19994
rect 4436 19848 4488 19854
rect 4436 19790 4488 19796
rect 4344 19712 4396 19718
rect 4344 19654 4396 19660
rect 4068 19372 4120 19378
rect 4068 19314 4120 19320
rect 4252 19372 4304 19378
rect 4252 19314 4304 19320
rect 3976 19236 4028 19242
rect 3976 19178 4028 19184
rect 3988 18426 4016 19178
rect 4080 18952 4108 19314
rect 4264 19281 4292 19314
rect 4250 19272 4306 19281
rect 4250 19207 4306 19216
rect 4356 19174 4384 19654
rect 4448 19310 4476 19790
rect 4436 19304 4488 19310
rect 4436 19246 4488 19252
rect 4540 19242 4568 19994
rect 4528 19236 4580 19242
rect 4528 19178 4580 19184
rect 4344 19168 4396 19174
rect 4344 19110 4396 19116
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4080 18924 4200 18952
rect 3976 18420 4028 18426
rect 3976 18362 4028 18368
rect 4172 18358 4200 18924
rect 3240 18352 3292 18358
rect 3240 18294 3292 18300
rect 3792 18352 3844 18358
rect 3792 18294 3844 18300
rect 4160 18352 4212 18358
rect 4160 18294 4212 18300
rect 3148 17536 3200 17542
rect 3148 17478 3200 17484
rect 3146 17232 3202 17241
rect 3146 17167 3148 17176
rect 3200 17167 3202 17176
rect 3148 17138 3200 17144
rect 3056 16448 3108 16454
rect 3056 16390 3108 16396
rect 2964 16244 3016 16250
rect 2964 16186 3016 16192
rect 2884 16102 3004 16130
rect 2780 15972 2832 15978
rect 2780 15914 2832 15920
rect 2688 15700 2740 15706
rect 2688 15642 2740 15648
rect 2700 15609 2728 15642
rect 2686 15600 2742 15609
rect 2792 15570 2820 15914
rect 2976 15910 3004 16102
rect 3068 16096 3096 16390
rect 3148 16108 3200 16114
rect 3068 16068 3148 16096
rect 2964 15904 3016 15910
rect 2964 15846 3016 15852
rect 2870 15736 2926 15745
rect 2870 15671 2926 15680
rect 2686 15535 2742 15544
rect 2780 15564 2832 15570
rect 2780 15506 2832 15512
rect 2884 15502 2912 15671
rect 2872 15496 2924 15502
rect 2872 15438 2924 15444
rect 2504 15020 2556 15026
rect 2504 14962 2556 14968
rect 2872 14068 2924 14074
rect 2872 14010 2924 14016
rect 2412 13864 2464 13870
rect 2412 13806 2464 13812
rect 2424 13462 2452 13806
rect 2412 13456 2464 13462
rect 2412 13398 2464 13404
rect 2424 12918 2452 13398
rect 2884 13326 2912 14010
rect 2872 13320 2924 13326
rect 2792 13280 2872 13308
rect 2412 12912 2464 12918
rect 2464 12860 2728 12866
rect 2412 12854 2728 12860
rect 2424 12838 2728 12854
rect 2320 12776 2372 12782
rect 2320 12718 2372 12724
rect 2504 12776 2556 12782
rect 2504 12718 2556 12724
rect 2516 12238 2544 12718
rect 2596 12708 2648 12714
rect 2596 12650 2648 12656
rect 2504 12232 2556 12238
rect 2504 12174 2556 12180
rect 2228 12096 2280 12102
rect 2228 12038 2280 12044
rect 2320 12096 2372 12102
rect 2320 12038 2372 12044
rect 2240 11898 2268 12038
rect 2228 11892 2280 11898
rect 2228 11834 2280 11840
rect 1860 11824 1912 11830
rect 1860 11766 1912 11772
rect 1768 11348 1820 11354
rect 1768 11290 1820 11296
rect 1676 11076 1728 11082
rect 1676 11018 1728 11024
rect 1688 10810 1716 11018
rect 1676 10804 1728 10810
rect 1676 10746 1728 10752
rect 1872 10470 1900 11766
rect 2240 11082 2268 11834
rect 2228 11076 2280 11082
rect 2228 11018 2280 11024
rect 2044 11008 2096 11014
rect 2044 10950 2096 10956
rect 2056 10742 2084 10950
rect 2044 10736 2096 10742
rect 2044 10678 2096 10684
rect 1860 10464 1912 10470
rect 1860 10406 1912 10412
rect 1872 9178 1900 10406
rect 1860 9172 1912 9178
rect 1860 9114 1912 9120
rect 1584 9104 1636 9110
rect 1584 9046 1636 9052
rect 1492 8900 1544 8906
rect 1492 8842 1544 8848
rect 1504 7478 1532 8842
rect 1492 7472 1544 7478
rect 1492 7414 1544 7420
rect 1596 7410 1624 9046
rect 1768 8832 1820 8838
rect 1768 8774 1820 8780
rect 1676 7880 1728 7886
rect 1780 7868 1808 8774
rect 1872 7970 1900 9114
rect 2056 8906 2084 10678
rect 2332 10674 2360 12038
rect 2608 11014 2636 12650
rect 2700 12306 2728 12838
rect 2792 12782 2820 13280
rect 2872 13262 2924 13268
rect 2872 13184 2924 13190
rect 2872 13126 2924 13132
rect 2884 12918 2912 13126
rect 2872 12912 2924 12918
rect 2872 12854 2924 12860
rect 2780 12776 2832 12782
rect 2832 12736 2912 12764
rect 2780 12718 2832 12724
rect 2688 12300 2740 12306
rect 2688 12242 2740 12248
rect 2780 12164 2832 12170
rect 2780 12106 2832 12112
rect 2792 11354 2820 12106
rect 2884 12073 2912 12736
rect 2870 12064 2926 12073
rect 2870 11999 2926 12008
rect 2872 11892 2924 11898
rect 2872 11834 2924 11840
rect 2884 11506 2912 11834
rect 2976 11642 3004 15846
rect 3068 15638 3096 16068
rect 3148 16050 3200 16056
rect 3252 15688 3280 18294
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4632 17882 4660 20318
rect 4724 19922 4752 21286
rect 4816 21078 4844 21848
rect 4874 21788 5182 21797
rect 4874 21786 4880 21788
rect 4936 21786 4960 21788
rect 5016 21786 5040 21788
rect 5096 21786 5120 21788
rect 5176 21786 5182 21788
rect 4936 21734 4938 21786
rect 5118 21734 5120 21786
rect 4874 21732 4880 21734
rect 4936 21732 4960 21734
rect 5016 21732 5040 21734
rect 5096 21732 5120 21734
rect 5176 21732 5182 21734
rect 4874 21723 5182 21732
rect 5276 21690 5304 24092
rect 5460 24070 5488 24126
rect 5540 24132 5592 24138
rect 5540 24074 5592 24080
rect 5356 24064 5408 24070
rect 5356 24006 5408 24012
rect 5448 24064 5500 24070
rect 5448 24006 5500 24012
rect 5368 23730 5396 24006
rect 5356 23724 5408 23730
rect 5356 23666 5408 23672
rect 5356 22976 5408 22982
rect 5356 22918 5408 22924
rect 5368 22506 5396 22918
rect 5460 22710 5488 24006
rect 5448 22704 5500 22710
rect 5448 22646 5500 22652
rect 5356 22500 5408 22506
rect 5356 22442 5408 22448
rect 5460 22386 5488 22646
rect 5552 22574 5580 24074
rect 5644 23798 5672 24754
rect 5816 24676 5868 24682
rect 5816 24618 5868 24624
rect 5632 23792 5684 23798
rect 5632 23734 5684 23740
rect 5828 22642 5856 24618
rect 5920 24274 5948 26182
rect 6104 25974 6132 26336
rect 6276 26376 6328 26382
rect 6276 26318 6328 26324
rect 6092 25968 6144 25974
rect 6092 25910 6144 25916
rect 5908 24268 5960 24274
rect 5908 24210 5960 24216
rect 6104 24138 6132 25910
rect 6552 25832 6604 25838
rect 6552 25774 6604 25780
rect 6564 25498 6592 25774
rect 6552 25492 6604 25498
rect 6552 25434 6604 25440
rect 6840 25430 6868 28494
rect 7012 28144 7064 28150
rect 7484 28098 7512 30110
rect 7668 28626 7696 31214
rect 8036 30938 8064 31214
rect 8024 30932 8076 30938
rect 8024 30874 8076 30880
rect 8404 30734 8432 31742
rect 8852 31690 8904 31696
rect 8484 31680 8536 31686
rect 8484 31622 8536 31628
rect 8496 31346 8524 31622
rect 8484 31340 8536 31346
rect 8484 31282 8536 31288
rect 8484 30864 8536 30870
rect 8484 30806 8536 30812
rect 8496 30734 8524 30806
rect 8864 30734 8892 31690
rect 9416 31142 9444 31758
rect 9692 31346 9720 31758
rect 10428 31754 10456 32710
rect 10428 31726 10548 31754
rect 9680 31340 9732 31346
rect 9680 31282 9732 31288
rect 9956 31340 10008 31346
rect 9956 31282 10008 31288
rect 9404 31136 9456 31142
rect 9404 31078 9456 31084
rect 8392 30728 8444 30734
rect 8392 30670 8444 30676
rect 8484 30728 8536 30734
rect 8484 30670 8536 30676
rect 8852 30728 8904 30734
rect 8852 30670 8904 30676
rect 9128 30728 9180 30734
rect 9128 30670 9180 30676
rect 9220 30728 9272 30734
rect 9220 30670 9272 30676
rect 8024 30592 8076 30598
rect 8024 30534 8076 30540
rect 8036 30326 8064 30534
rect 8024 30320 8076 30326
rect 8024 30262 8076 30268
rect 7932 30252 7984 30258
rect 7932 30194 7984 30200
rect 7748 30048 7800 30054
rect 7748 29990 7800 29996
rect 7760 29714 7788 29990
rect 7840 29844 7892 29850
rect 7840 29786 7892 29792
rect 7748 29708 7800 29714
rect 7748 29650 7800 29656
rect 7656 28620 7708 28626
rect 7656 28562 7708 28568
rect 7564 28416 7616 28422
rect 7564 28358 7616 28364
rect 7012 28086 7064 28092
rect 6920 27872 6972 27878
rect 6920 27814 6972 27820
rect 6932 26994 6960 27814
rect 7024 27674 7052 28086
rect 7104 28076 7156 28082
rect 7104 28018 7156 28024
rect 7288 28076 7340 28082
rect 7288 28018 7340 28024
rect 7392 28070 7512 28098
rect 7012 27668 7064 27674
rect 7012 27610 7064 27616
rect 7116 27606 7144 28018
rect 7196 28008 7248 28014
rect 7196 27950 7248 27956
rect 7104 27600 7156 27606
rect 7104 27542 7156 27548
rect 7012 27328 7064 27334
rect 7012 27270 7064 27276
rect 6920 26988 6972 26994
rect 6920 26930 6972 26936
rect 6920 26308 6972 26314
rect 6920 26250 6972 26256
rect 6932 26042 6960 26250
rect 6920 26036 6972 26042
rect 6920 25978 6972 25984
rect 7024 25498 7052 27270
rect 7104 27056 7156 27062
rect 7104 26998 7156 27004
rect 7116 26382 7144 26998
rect 7104 26376 7156 26382
rect 7104 26318 7156 26324
rect 7208 25770 7236 27950
rect 7300 27402 7328 28018
rect 7392 27674 7420 28070
rect 7380 27668 7432 27674
rect 7380 27610 7432 27616
rect 7288 27396 7340 27402
rect 7288 27338 7340 27344
rect 7300 26586 7328 27338
rect 7288 26580 7340 26586
rect 7288 26522 7340 26528
rect 7196 25764 7248 25770
rect 7196 25706 7248 25712
rect 7012 25492 7064 25498
rect 7012 25434 7064 25440
rect 6828 25424 6880 25430
rect 6828 25366 6880 25372
rect 6644 25356 6696 25362
rect 6644 25298 6696 25304
rect 6184 24676 6236 24682
rect 6184 24618 6236 24624
rect 6276 24676 6328 24682
rect 6276 24618 6328 24624
rect 6196 24410 6224 24618
rect 6184 24404 6236 24410
rect 6184 24346 6236 24352
rect 6092 24132 6144 24138
rect 6092 24074 6144 24080
rect 5908 23520 5960 23526
rect 5908 23462 5960 23468
rect 5816 22636 5868 22642
rect 5816 22578 5868 22584
rect 5540 22568 5592 22574
rect 5540 22510 5592 22516
rect 5368 22358 5488 22386
rect 5632 22432 5684 22438
rect 5632 22374 5684 22380
rect 5368 21690 5396 22358
rect 5448 22024 5500 22030
rect 5448 21966 5500 21972
rect 5264 21684 5316 21690
rect 5264 21626 5316 21632
rect 5356 21684 5408 21690
rect 5356 21626 5408 21632
rect 4988 21616 5040 21622
rect 4988 21558 5040 21564
rect 4896 21548 4948 21554
rect 4896 21490 4948 21496
rect 4804 21072 4856 21078
rect 4804 21014 4856 21020
rect 4908 20942 4936 21490
rect 5000 21078 5028 21558
rect 5080 21480 5132 21486
rect 5080 21422 5132 21428
rect 4988 21072 5040 21078
rect 4988 21014 5040 21020
rect 5092 21010 5120 21422
rect 5276 21418 5304 21626
rect 5264 21412 5316 21418
rect 5264 21354 5316 21360
rect 5080 21004 5132 21010
rect 5080 20946 5132 20952
rect 5276 20942 5304 21354
rect 4896 20936 4948 20942
rect 4896 20878 4948 20884
rect 5264 20936 5316 20942
rect 5264 20878 5316 20884
rect 5368 20874 5396 21626
rect 5356 20868 5408 20874
rect 5356 20810 5408 20816
rect 4804 20800 4856 20806
rect 4804 20742 4856 20748
rect 4816 20058 4844 20742
rect 4874 20700 5182 20709
rect 4874 20698 4880 20700
rect 4936 20698 4960 20700
rect 5016 20698 5040 20700
rect 5096 20698 5120 20700
rect 5176 20698 5182 20700
rect 4936 20646 4938 20698
rect 5118 20646 5120 20698
rect 4874 20644 4880 20646
rect 4936 20644 4960 20646
rect 5016 20644 5040 20646
rect 5096 20644 5120 20646
rect 5176 20644 5182 20646
rect 4874 20635 5182 20644
rect 5264 20392 5316 20398
rect 5264 20334 5316 20340
rect 4896 20324 4948 20330
rect 4896 20266 4948 20272
rect 4804 20052 4856 20058
rect 4804 19994 4856 20000
rect 4712 19916 4764 19922
rect 4712 19858 4764 19864
rect 4724 19378 4752 19858
rect 4908 19854 4936 20266
rect 5172 19916 5224 19922
rect 5172 19858 5224 19864
rect 4896 19848 4948 19854
rect 5184 19825 5212 19858
rect 4896 19790 4948 19796
rect 5170 19816 5226 19825
rect 5170 19751 5226 19760
rect 4874 19612 5182 19621
rect 4874 19610 4880 19612
rect 4936 19610 4960 19612
rect 5016 19610 5040 19612
rect 5096 19610 5120 19612
rect 5176 19610 5182 19612
rect 4936 19558 4938 19610
rect 5118 19558 5120 19610
rect 4874 19556 4880 19558
rect 4936 19556 4960 19558
rect 5016 19556 5040 19558
rect 5096 19556 5120 19558
rect 5176 19556 5182 19558
rect 4874 19547 5182 19556
rect 5276 19514 5304 20334
rect 5460 19854 5488 21966
rect 5644 21622 5672 22374
rect 5828 22098 5856 22578
rect 5816 22092 5868 22098
rect 5816 22034 5868 22040
rect 5632 21616 5684 21622
rect 5632 21558 5684 21564
rect 5816 21616 5868 21622
rect 5816 21558 5868 21564
rect 5828 21434 5856 21558
rect 5920 21554 5948 23462
rect 5908 21548 5960 21554
rect 5908 21490 5960 21496
rect 5828 21406 5948 21434
rect 5632 21344 5684 21350
rect 5632 21286 5684 21292
rect 5816 21344 5868 21350
rect 5816 21286 5868 21292
rect 5644 19854 5672 21286
rect 5448 19848 5500 19854
rect 5354 19816 5410 19825
rect 5448 19790 5500 19796
rect 5632 19848 5684 19854
rect 5632 19790 5684 19796
rect 5828 19786 5856 21286
rect 5920 21162 5948 21406
rect 5920 21134 6040 21162
rect 5354 19751 5410 19760
rect 5816 19780 5868 19786
rect 4804 19508 4856 19514
rect 4804 19450 4856 19456
rect 5264 19508 5316 19514
rect 5264 19450 5316 19456
rect 4712 19372 4764 19378
rect 4712 19314 4764 19320
rect 4712 19168 4764 19174
rect 4712 19110 4764 19116
rect 3332 17876 3384 17882
rect 3332 17818 3384 17824
rect 4620 17876 4672 17882
rect 4620 17818 4672 17824
rect 3344 17678 3372 17818
rect 3792 17808 3844 17814
rect 3436 17734 3648 17762
rect 3792 17750 3844 17756
rect 3436 17678 3464 17734
rect 3332 17672 3384 17678
rect 3332 17614 3384 17620
rect 3424 17672 3476 17678
rect 3424 17614 3476 17620
rect 3344 16454 3372 17614
rect 3516 17604 3568 17610
rect 3516 17546 3568 17552
rect 3424 17536 3476 17542
rect 3424 17478 3476 17484
rect 3332 16448 3384 16454
rect 3332 16390 3384 16396
rect 3344 16182 3372 16390
rect 3332 16176 3384 16182
rect 3332 16118 3384 16124
rect 3160 15660 3280 15688
rect 3056 15632 3108 15638
rect 3056 15574 3108 15580
rect 3160 15473 3188 15660
rect 3238 15600 3294 15609
rect 3238 15535 3294 15544
rect 3332 15564 3384 15570
rect 3146 15464 3202 15473
rect 3146 15399 3202 15408
rect 3160 15366 3188 15399
rect 3148 15360 3200 15366
rect 3148 15302 3200 15308
rect 3160 14074 3188 15302
rect 3252 14260 3280 15535
rect 3332 15506 3384 15512
rect 3344 14414 3372 15506
rect 3436 15502 3464 17478
rect 3528 17202 3556 17546
rect 3516 17196 3568 17202
rect 3516 17138 3568 17144
rect 3516 16448 3568 16454
rect 3516 16390 3568 16396
rect 3528 16250 3556 16390
rect 3516 16244 3568 16250
rect 3516 16186 3568 16192
rect 3620 16114 3648 17734
rect 3804 17678 3832 17750
rect 3792 17672 3844 17678
rect 3884 17672 3936 17678
rect 3792 17614 3844 17620
rect 3882 17640 3884 17649
rect 3936 17640 3938 17649
rect 3882 17575 3938 17584
rect 4068 17604 4120 17610
rect 3700 17196 3752 17202
rect 3700 17138 3752 17144
rect 3712 16794 3740 17138
rect 3792 16992 3844 16998
rect 3792 16934 3844 16940
rect 3700 16788 3752 16794
rect 3700 16730 3752 16736
rect 3804 16590 3832 16934
rect 3792 16584 3844 16590
rect 3792 16526 3844 16532
rect 3608 16108 3660 16114
rect 3608 16050 3660 16056
rect 3620 15978 3648 16050
rect 3896 16028 3924 17575
rect 4068 17546 4120 17552
rect 4080 16998 4108 17546
rect 4068 16992 4120 16998
rect 4068 16934 4120 16940
rect 4080 16590 4108 16934
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4632 16590 4660 17818
rect 4724 16658 4752 19110
rect 4712 16652 4764 16658
rect 4712 16594 4764 16600
rect 4068 16584 4120 16590
rect 4068 16526 4120 16532
rect 4252 16584 4304 16590
rect 4252 16526 4304 16532
rect 4620 16584 4672 16590
rect 4620 16526 4672 16532
rect 3976 16516 4028 16522
rect 3976 16458 4028 16464
rect 3988 16250 4016 16458
rect 3976 16244 4028 16250
rect 3976 16186 4028 16192
rect 4080 16114 4108 16526
rect 4160 16448 4212 16454
rect 4160 16390 4212 16396
rect 4068 16108 4120 16114
rect 4068 16050 4120 16056
rect 3976 16040 4028 16046
rect 3896 16000 3976 16028
rect 3608 15972 3660 15978
rect 3608 15914 3660 15920
rect 3620 15638 3648 15914
rect 3896 15706 3924 16000
rect 4172 15994 4200 16390
rect 4264 16114 4292 16526
rect 4712 16516 4764 16522
rect 4712 16458 4764 16464
rect 4528 16448 4580 16454
rect 4528 16390 4580 16396
rect 4252 16108 4304 16114
rect 4252 16050 4304 16056
rect 4344 16108 4396 16114
rect 4344 16050 4396 16056
rect 3976 15982 4028 15988
rect 4080 15966 4200 15994
rect 4356 15978 4384 16050
rect 4344 15972 4396 15978
rect 3884 15700 3936 15706
rect 4080 15688 4108 15966
rect 4344 15914 4396 15920
rect 4540 15910 4568 16390
rect 4620 16244 4672 16250
rect 4620 16186 4672 16192
rect 4528 15904 4580 15910
rect 4528 15846 4580 15852
rect 4632 15858 4660 16186
rect 4724 16114 4752 16458
rect 4712 16108 4764 16114
rect 4712 16050 4764 16056
rect 4632 15830 4752 15858
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4620 15700 4672 15706
rect 4080 15660 4200 15688
rect 3884 15642 3936 15648
rect 3608 15632 3660 15638
rect 3608 15574 3660 15580
rect 3896 15502 3924 15642
rect 3424 15496 3476 15502
rect 3424 15438 3476 15444
rect 3884 15496 3936 15502
rect 4068 15496 4120 15502
rect 3884 15438 3936 15444
rect 4066 15464 4068 15473
rect 4120 15464 4122 15473
rect 3700 15428 3752 15434
rect 4066 15399 4122 15408
rect 3700 15370 3752 15376
rect 3712 15162 3740 15370
rect 3884 15360 3936 15366
rect 3884 15302 3936 15308
rect 3976 15360 4028 15366
rect 3976 15302 4028 15308
rect 3700 15156 3752 15162
rect 3700 15098 3752 15104
rect 3332 14408 3384 14414
rect 3332 14350 3384 14356
rect 3424 14272 3476 14278
rect 3252 14232 3372 14260
rect 3148 14068 3200 14074
rect 3148 14010 3200 14016
rect 3148 13456 3200 13462
rect 3148 13398 3200 13404
rect 3056 13320 3108 13326
rect 3056 13262 3108 13268
rect 3068 12374 3096 13262
rect 3160 12850 3188 13398
rect 3240 13252 3292 13258
rect 3240 13194 3292 13200
rect 3148 12844 3200 12850
rect 3148 12786 3200 12792
rect 3148 12640 3200 12646
rect 3148 12582 3200 12588
rect 3056 12368 3108 12374
rect 3056 12310 3108 12316
rect 3160 12102 3188 12582
rect 3252 12442 3280 13194
rect 3240 12436 3292 12442
rect 3240 12378 3292 12384
rect 3148 12096 3200 12102
rect 3148 12038 3200 12044
rect 3344 11914 3372 14232
rect 3424 14214 3476 14220
rect 3436 13433 3464 14214
rect 3792 14000 3844 14006
rect 3606 13968 3662 13977
rect 3792 13942 3844 13948
rect 3606 13903 3608 13912
rect 3660 13903 3662 13912
rect 3608 13874 3660 13880
rect 3608 13796 3660 13802
rect 3528 13756 3608 13784
rect 3422 13424 3478 13433
rect 3422 13359 3478 13368
rect 3528 13274 3556 13756
rect 3608 13738 3660 13744
rect 3700 13728 3752 13734
rect 3606 13696 3662 13705
rect 3700 13670 3752 13676
rect 3606 13631 3662 13640
rect 3620 13326 3648 13631
rect 3436 13258 3556 13274
rect 3608 13320 3660 13326
rect 3608 13262 3660 13268
rect 3424 13252 3556 13258
rect 3476 13246 3556 13252
rect 3424 13194 3476 13200
rect 3516 13184 3568 13190
rect 3516 13126 3568 13132
rect 3424 12640 3476 12646
rect 3528 12628 3556 13126
rect 3620 12730 3648 13262
rect 3712 12850 3740 13670
rect 3804 12986 3832 13942
rect 3896 13433 3924 15302
rect 3988 13734 4016 15302
rect 4172 14872 4200 15660
rect 4620 15642 4672 15648
rect 4080 14844 4200 14872
rect 4080 14482 4108 14844
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4068 14476 4120 14482
rect 4068 14418 4120 14424
rect 4080 13870 4108 14418
rect 4632 14414 4660 15642
rect 4724 15026 4752 15830
rect 4816 15706 4844 19450
rect 5170 19408 5226 19417
rect 5170 19343 5172 19352
rect 5224 19343 5226 19352
rect 5172 19314 5224 19320
rect 4874 18524 5182 18533
rect 4874 18522 4880 18524
rect 4936 18522 4960 18524
rect 5016 18522 5040 18524
rect 5096 18522 5120 18524
rect 5176 18522 5182 18524
rect 4936 18470 4938 18522
rect 5118 18470 5120 18522
rect 4874 18468 4880 18470
rect 4936 18468 4960 18470
rect 5016 18468 5040 18470
rect 5096 18468 5120 18470
rect 5176 18468 5182 18470
rect 4874 18459 5182 18468
rect 4988 18284 5040 18290
rect 4988 18226 5040 18232
rect 5172 18284 5224 18290
rect 5172 18226 5224 18232
rect 5000 17678 5028 18226
rect 5184 17678 5212 18226
rect 5368 17882 5396 19751
rect 5816 19722 5868 19728
rect 5828 19378 5856 19722
rect 5908 19712 5960 19718
rect 5908 19654 5960 19660
rect 5920 19446 5948 19654
rect 5908 19440 5960 19446
rect 6012 19417 6040 21134
rect 6104 20398 6132 24074
rect 6288 24070 6316 24618
rect 6184 24064 6236 24070
rect 6184 24006 6236 24012
rect 6276 24064 6328 24070
rect 6276 24006 6328 24012
rect 6196 23118 6224 24006
rect 6288 23526 6316 24006
rect 6276 23520 6328 23526
rect 6276 23462 6328 23468
rect 6184 23112 6236 23118
rect 6184 23054 6236 23060
rect 6368 23112 6420 23118
rect 6368 23054 6420 23060
rect 6276 22568 6328 22574
rect 6276 22510 6328 22516
rect 6184 22500 6236 22506
rect 6184 22442 6236 22448
rect 6196 21622 6224 22442
rect 6184 21616 6236 21622
rect 6184 21558 6236 21564
rect 6288 21078 6316 22510
rect 6380 22166 6408 23054
rect 6460 22636 6512 22642
rect 6460 22578 6512 22584
rect 6368 22160 6420 22166
rect 6368 22102 6420 22108
rect 6380 22030 6408 22102
rect 6368 22024 6420 22030
rect 6368 21966 6420 21972
rect 6380 21078 6408 21966
rect 6276 21072 6328 21078
rect 6276 21014 6328 21020
rect 6368 21072 6420 21078
rect 6368 21014 6420 21020
rect 6092 20392 6144 20398
rect 6092 20334 6144 20340
rect 6288 20058 6316 21014
rect 6472 20942 6500 22578
rect 6656 21554 6684 25298
rect 7208 25294 7236 25706
rect 7196 25288 7248 25294
rect 7196 25230 7248 25236
rect 7104 24812 7156 24818
rect 7104 24754 7156 24760
rect 7116 24410 7144 24754
rect 7104 24404 7156 24410
rect 7104 24346 7156 24352
rect 7392 24274 7420 27610
rect 7472 26784 7524 26790
rect 7472 26726 7524 26732
rect 7380 24268 7432 24274
rect 7380 24210 7432 24216
rect 6920 22976 6972 22982
rect 6920 22918 6972 22924
rect 6828 22024 6880 22030
rect 6828 21966 6880 21972
rect 6736 21888 6788 21894
rect 6736 21830 6788 21836
rect 6644 21548 6696 21554
rect 6644 21490 6696 21496
rect 6552 21344 6604 21350
rect 6552 21286 6604 21292
rect 6460 20936 6512 20942
rect 6460 20878 6512 20884
rect 6472 20602 6500 20878
rect 6460 20596 6512 20602
rect 6460 20538 6512 20544
rect 6276 20052 6328 20058
rect 6276 19994 6328 20000
rect 6472 19514 6500 20538
rect 6460 19508 6512 19514
rect 6460 19450 6512 19456
rect 5908 19382 5960 19388
rect 5998 19408 6054 19417
rect 5816 19372 5868 19378
rect 5998 19343 6054 19352
rect 5816 19314 5868 19320
rect 6564 19174 6592 21286
rect 6656 20330 6684 21490
rect 6748 21010 6776 21830
rect 6840 21622 6868 21966
rect 6828 21616 6880 21622
rect 6828 21558 6880 21564
rect 6932 21554 6960 22918
rect 7012 21956 7064 21962
rect 7012 21898 7064 21904
rect 7024 21622 7052 21898
rect 7012 21616 7064 21622
rect 7012 21558 7064 21564
rect 6920 21548 6972 21554
rect 6920 21490 6972 21496
rect 7288 21140 7340 21146
rect 7288 21082 7340 21088
rect 6736 21004 6788 21010
rect 6736 20946 6788 20952
rect 7300 20534 7328 21082
rect 7288 20528 7340 20534
rect 7288 20470 7340 20476
rect 6644 20324 6696 20330
rect 6644 20266 6696 20272
rect 6920 19304 6972 19310
rect 6920 19246 6972 19252
rect 6552 19168 6604 19174
rect 6552 19110 6604 19116
rect 6644 19168 6696 19174
rect 6644 19110 6696 19116
rect 6000 18624 6052 18630
rect 6000 18566 6052 18572
rect 6012 18290 6040 18566
rect 6656 18290 6684 19110
rect 6932 18766 6960 19246
rect 6920 18760 6972 18766
rect 6920 18702 6972 18708
rect 6932 18290 6960 18702
rect 7012 18692 7064 18698
rect 7012 18634 7064 18640
rect 7024 18358 7052 18634
rect 7104 18624 7156 18630
rect 7104 18566 7156 18572
rect 7012 18352 7064 18358
rect 7012 18294 7064 18300
rect 6000 18284 6052 18290
rect 6000 18226 6052 18232
rect 6644 18284 6696 18290
rect 6644 18226 6696 18232
rect 6920 18284 6972 18290
rect 6920 18226 6972 18232
rect 5356 17876 5408 17882
rect 5356 17818 5408 17824
rect 4988 17672 5040 17678
rect 4988 17614 5040 17620
rect 5172 17672 5224 17678
rect 5172 17614 5224 17620
rect 5184 17542 5212 17614
rect 5172 17536 5224 17542
rect 5172 17478 5224 17484
rect 4874 17436 5182 17445
rect 4874 17434 4880 17436
rect 4936 17434 4960 17436
rect 5016 17434 5040 17436
rect 5096 17434 5120 17436
rect 5176 17434 5182 17436
rect 4936 17382 4938 17434
rect 5118 17382 5120 17434
rect 4874 17380 4880 17382
rect 4936 17380 4960 17382
rect 5016 17380 5040 17382
rect 5096 17380 5120 17382
rect 5176 17380 5182 17382
rect 4874 17371 5182 17380
rect 5368 17354 5396 17818
rect 6092 17536 6144 17542
rect 6092 17478 6144 17484
rect 5368 17326 5488 17354
rect 5080 17264 5132 17270
rect 5080 17206 5132 17212
rect 5356 17264 5408 17270
rect 5356 17206 5408 17212
rect 5092 16658 5120 17206
rect 5264 16992 5316 16998
rect 5264 16934 5316 16940
rect 5276 16794 5304 16934
rect 5264 16788 5316 16794
rect 5264 16730 5316 16736
rect 5080 16652 5132 16658
rect 5080 16594 5132 16600
rect 5264 16652 5316 16658
rect 5264 16594 5316 16600
rect 4874 16348 5182 16357
rect 4874 16346 4880 16348
rect 4936 16346 4960 16348
rect 5016 16346 5040 16348
rect 5096 16346 5120 16348
rect 5176 16346 5182 16348
rect 4936 16294 4938 16346
rect 5118 16294 5120 16346
rect 4874 16292 4880 16294
rect 4936 16292 4960 16294
rect 5016 16292 5040 16294
rect 5096 16292 5120 16294
rect 5176 16292 5182 16294
rect 4874 16283 5182 16292
rect 5080 16176 5132 16182
rect 5080 16118 5132 16124
rect 4988 15972 5040 15978
rect 4988 15914 5040 15920
rect 4896 15904 4948 15910
rect 4896 15846 4948 15852
rect 4804 15700 4856 15706
rect 4804 15642 4856 15648
rect 4908 15586 4936 15846
rect 4816 15570 4936 15586
rect 4804 15564 4936 15570
rect 4856 15558 4936 15564
rect 4804 15506 4856 15512
rect 4712 15020 4764 15026
rect 4712 14962 4764 14968
rect 4712 14816 4764 14822
rect 4712 14758 4764 14764
rect 4344 14408 4396 14414
rect 4344 14350 4396 14356
rect 4620 14408 4672 14414
rect 4620 14350 4672 14356
rect 4252 14272 4304 14278
rect 4252 14214 4304 14220
rect 4264 13938 4292 14214
rect 4252 13932 4304 13938
rect 4252 13874 4304 13880
rect 4068 13864 4120 13870
rect 4068 13806 4120 13812
rect 4356 13802 4384 14350
rect 4620 14272 4672 14278
rect 4620 14214 4672 14220
rect 4436 13932 4488 13938
rect 4436 13874 4488 13880
rect 4344 13796 4396 13802
rect 4344 13738 4396 13744
rect 4448 13734 4476 13874
rect 3976 13728 4028 13734
rect 3976 13670 4028 13676
rect 4068 13728 4120 13734
rect 4068 13670 4120 13676
rect 4436 13728 4488 13734
rect 4436 13670 4488 13676
rect 3882 13424 3938 13433
rect 3882 13359 3938 13368
rect 3792 12980 3844 12986
rect 3792 12922 3844 12928
rect 3988 12850 4016 13670
rect 3700 12844 3752 12850
rect 3700 12786 3752 12792
rect 3976 12844 4028 12850
rect 3976 12786 4028 12792
rect 3884 12776 3936 12782
rect 3620 12702 3740 12730
rect 3884 12718 3936 12724
rect 3476 12600 3556 12628
rect 3608 12640 3660 12646
rect 3424 12582 3476 12588
rect 3608 12582 3660 12588
rect 3422 12336 3478 12345
rect 3478 12280 3556 12288
rect 3422 12271 3424 12280
rect 3476 12260 3556 12280
rect 3424 12242 3476 12248
rect 3252 11886 3372 11914
rect 3252 11830 3280 11886
rect 3148 11824 3200 11830
rect 3148 11766 3200 11772
rect 3240 11824 3292 11830
rect 3240 11766 3292 11772
rect 2976 11614 3096 11642
rect 3068 11558 3096 11614
rect 2964 11552 3016 11558
rect 2884 11500 2964 11506
rect 2884 11494 3016 11500
rect 3056 11552 3108 11558
rect 3056 11494 3108 11500
rect 2884 11478 3004 11494
rect 3160 11354 3188 11766
rect 2780 11348 2832 11354
rect 2780 11290 2832 11296
rect 3148 11348 3200 11354
rect 3148 11290 3200 11296
rect 2780 11144 2832 11150
rect 2780 11086 2832 11092
rect 2596 11008 2648 11014
rect 2596 10950 2648 10956
rect 2608 10742 2636 10950
rect 2596 10736 2648 10742
rect 2596 10678 2648 10684
rect 2320 10668 2372 10674
rect 2320 10610 2372 10616
rect 2332 9042 2360 10610
rect 2792 10130 2820 11086
rect 3148 11076 3200 11082
rect 3148 11018 3200 11024
rect 2780 10124 2832 10130
rect 2780 10066 2832 10072
rect 2320 9036 2372 9042
rect 2320 8978 2372 8984
rect 2332 8922 2360 8978
rect 2044 8900 2096 8906
rect 2332 8894 2452 8922
rect 2096 8860 2268 8888
rect 2044 8842 2096 8848
rect 1872 7942 1992 7970
rect 1860 7880 1912 7886
rect 1780 7840 1860 7868
rect 1676 7822 1728 7828
rect 1860 7822 1912 7828
rect 1688 7410 1716 7822
rect 1584 7404 1636 7410
rect 1584 7346 1636 7352
rect 1676 7404 1728 7410
rect 1676 7346 1728 7352
rect 1964 7206 1992 7942
rect 2240 7410 2268 8860
rect 2320 8832 2372 8838
rect 2320 8774 2372 8780
rect 2332 8634 2360 8774
rect 2320 8628 2372 8634
rect 2320 8570 2372 8576
rect 2424 8566 2452 8894
rect 2412 8560 2464 8566
rect 2412 8502 2464 8508
rect 2424 7818 2452 8502
rect 2792 8498 2820 10066
rect 2964 9512 3016 9518
rect 2964 9454 3016 9460
rect 2976 8906 3004 9454
rect 3160 8974 3188 11018
rect 3252 10810 3280 11766
rect 3528 11762 3556 12260
rect 3424 11756 3476 11762
rect 3424 11698 3476 11704
rect 3516 11756 3568 11762
rect 3516 11698 3568 11704
rect 3436 11558 3464 11698
rect 3424 11552 3476 11558
rect 3424 11494 3476 11500
rect 3516 11552 3568 11558
rect 3516 11494 3568 11500
rect 3240 10804 3292 10810
rect 3240 10746 3292 10752
rect 3252 10266 3280 10746
rect 3436 10538 3464 11494
rect 3528 10674 3556 11494
rect 3516 10668 3568 10674
rect 3516 10610 3568 10616
rect 3424 10532 3476 10538
rect 3424 10474 3476 10480
rect 3240 10260 3292 10266
rect 3240 10202 3292 10208
rect 3620 10062 3648 12582
rect 3332 10056 3384 10062
rect 3332 9998 3384 10004
rect 3608 10056 3660 10062
rect 3608 9998 3660 10004
rect 3344 9722 3372 9998
rect 3332 9716 3384 9722
rect 3332 9658 3384 9664
rect 3332 9580 3384 9586
rect 3332 9522 3384 9528
rect 3148 8968 3200 8974
rect 3148 8910 3200 8916
rect 2964 8900 3016 8906
rect 2964 8842 3016 8848
rect 2872 8832 2924 8838
rect 2872 8774 2924 8780
rect 2884 8566 2912 8774
rect 2872 8560 2924 8566
rect 2872 8502 2924 8508
rect 2504 8492 2556 8498
rect 2504 8434 2556 8440
rect 2780 8492 2832 8498
rect 2780 8434 2832 8440
rect 2412 7812 2464 7818
rect 2412 7754 2464 7760
rect 2228 7404 2280 7410
rect 2228 7346 2280 7352
rect 1952 7200 2004 7206
rect 1952 7142 2004 7148
rect 2240 6730 2268 7346
rect 2320 7200 2372 7206
rect 2320 7142 2372 7148
rect 2332 7002 2360 7142
rect 2320 6996 2372 7002
rect 2320 6938 2372 6944
rect 2424 6934 2452 7754
rect 2412 6928 2464 6934
rect 2412 6870 2464 6876
rect 2320 6860 2372 6866
rect 2320 6802 2372 6808
rect 2332 6730 2360 6802
rect 2228 6724 2280 6730
rect 2228 6666 2280 6672
rect 2320 6724 2372 6730
rect 2320 6666 2372 6672
rect 2516 6662 2544 8434
rect 2792 8090 2820 8434
rect 2884 8090 2912 8502
rect 2964 8356 3016 8362
rect 2964 8298 3016 8304
rect 2780 8084 2832 8090
rect 2780 8026 2832 8032
rect 2872 8084 2924 8090
rect 2872 8026 2924 8032
rect 2596 8016 2648 8022
rect 2596 7958 2648 7964
rect 2608 6662 2636 7958
rect 2792 6866 2820 8026
rect 2872 7744 2924 7750
rect 2872 7686 2924 7692
rect 2780 6860 2832 6866
rect 2780 6802 2832 6808
rect 2884 6798 2912 7686
rect 2976 7546 3004 8298
rect 3160 8294 3188 8910
rect 3344 8838 3372 9522
rect 3608 9512 3660 9518
rect 3608 9454 3660 9460
rect 3620 9178 3648 9454
rect 3608 9172 3660 9178
rect 3608 9114 3660 9120
rect 3712 9042 3740 12702
rect 3896 12434 3924 12718
rect 3804 12406 3924 12434
rect 3804 11506 3832 12406
rect 3884 12164 3936 12170
rect 3884 12106 3936 12112
rect 3896 11626 3924 12106
rect 3976 12096 4028 12102
rect 3976 12038 4028 12044
rect 3988 11898 4016 12038
rect 3976 11892 4028 11898
rect 3976 11834 4028 11840
rect 3976 11756 4028 11762
rect 3976 11698 4028 11704
rect 3884 11620 3936 11626
rect 3884 11562 3936 11568
rect 3988 11506 4016 11698
rect 3804 11478 4016 11506
rect 3804 11082 3832 11478
rect 3792 11076 3844 11082
rect 3792 11018 3844 11024
rect 4080 10674 4108 13670
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4252 13456 4304 13462
rect 4250 13424 4252 13433
rect 4304 13424 4306 13433
rect 4250 13359 4306 13368
rect 4252 13320 4304 13326
rect 4250 13288 4252 13297
rect 4304 13288 4306 13297
rect 4250 13223 4306 13232
rect 4160 13184 4212 13190
rect 4160 13126 4212 13132
rect 4172 12850 4200 13126
rect 4160 12844 4212 12850
rect 4160 12786 4212 12792
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4632 12434 4660 14214
rect 4724 12646 4752 14758
rect 4816 14346 4844 15506
rect 5000 15502 5028 15914
rect 4896 15496 4948 15502
rect 4894 15464 4896 15473
rect 4988 15496 5040 15502
rect 4948 15464 4950 15473
rect 5092 15473 5120 16118
rect 5170 15600 5226 15609
rect 5170 15535 5226 15544
rect 5184 15502 5212 15535
rect 5172 15496 5224 15502
rect 4988 15438 5040 15444
rect 5078 15464 5134 15473
rect 4894 15399 4950 15408
rect 5172 15438 5224 15444
rect 5078 15399 5134 15408
rect 4874 15260 5182 15269
rect 4874 15258 4880 15260
rect 4936 15258 4960 15260
rect 5016 15258 5040 15260
rect 5096 15258 5120 15260
rect 5176 15258 5182 15260
rect 4936 15206 4938 15258
rect 5118 15206 5120 15258
rect 4874 15204 4880 15206
rect 4936 15204 4960 15206
rect 5016 15204 5040 15206
rect 5096 15204 5120 15206
rect 5176 15204 5182 15206
rect 4874 15195 5182 15204
rect 4896 15156 4948 15162
rect 4896 15098 4948 15104
rect 4908 14482 4936 15098
rect 5172 15020 5224 15026
rect 5172 14962 5224 14968
rect 4896 14476 4948 14482
rect 4896 14418 4948 14424
rect 4804 14340 4856 14346
rect 4804 14282 4856 14288
rect 4816 13977 4844 14282
rect 5184 14278 5212 14962
rect 5276 14414 5304 16594
rect 5368 15706 5396 17206
rect 5356 15700 5408 15706
rect 5356 15642 5408 15648
rect 5460 15570 5488 17326
rect 5632 17196 5684 17202
rect 5632 17138 5684 17144
rect 5908 17196 5960 17202
rect 5908 17138 5960 17144
rect 5540 16992 5592 16998
rect 5540 16934 5592 16940
rect 5552 16590 5580 16934
rect 5540 16584 5592 16590
rect 5540 16526 5592 16532
rect 5644 16182 5672 17138
rect 5724 17128 5776 17134
rect 5724 17070 5776 17076
rect 5736 16182 5764 17070
rect 5816 16992 5868 16998
rect 5816 16934 5868 16940
rect 5632 16176 5684 16182
rect 5632 16118 5684 16124
rect 5724 16176 5776 16182
rect 5724 16118 5776 16124
rect 5540 15972 5592 15978
rect 5540 15914 5592 15920
rect 5724 15972 5776 15978
rect 5724 15914 5776 15920
rect 5448 15564 5500 15570
rect 5448 15506 5500 15512
rect 5448 15088 5500 15094
rect 5448 15030 5500 15036
rect 5460 14414 5488 15030
rect 5552 15026 5580 15914
rect 5632 15904 5684 15910
rect 5632 15846 5684 15852
rect 5644 15706 5672 15846
rect 5632 15700 5684 15706
rect 5632 15642 5684 15648
rect 5644 15502 5672 15642
rect 5632 15496 5684 15502
rect 5632 15438 5684 15444
rect 5540 15020 5592 15026
rect 5540 14962 5592 14968
rect 5644 14618 5672 15438
rect 5736 15162 5764 15914
rect 5828 15910 5856 16934
rect 5920 16794 5948 17138
rect 5908 16788 5960 16794
rect 5908 16730 5960 16736
rect 5920 16250 5948 16730
rect 6000 16516 6052 16522
rect 6000 16458 6052 16464
rect 6012 16250 6040 16458
rect 5908 16244 5960 16250
rect 5908 16186 5960 16192
rect 6000 16244 6052 16250
rect 6000 16186 6052 16192
rect 5816 15904 5868 15910
rect 5816 15846 5868 15852
rect 5920 15502 5948 16186
rect 5908 15496 5960 15502
rect 5908 15438 5960 15444
rect 5816 15428 5868 15434
rect 5816 15370 5868 15376
rect 5828 15337 5856 15370
rect 5814 15328 5870 15337
rect 5814 15263 5870 15272
rect 5724 15156 5776 15162
rect 5776 15116 5948 15144
rect 5724 15098 5776 15104
rect 5632 14612 5684 14618
rect 5632 14554 5684 14560
rect 5264 14408 5316 14414
rect 5264 14350 5316 14356
rect 5448 14408 5500 14414
rect 5448 14350 5500 14356
rect 5172 14272 5224 14278
rect 5172 14214 5224 14220
rect 4874 14172 5182 14181
rect 4874 14170 4880 14172
rect 4936 14170 4960 14172
rect 5016 14170 5040 14172
rect 5096 14170 5120 14172
rect 5176 14170 5182 14172
rect 4936 14118 4938 14170
rect 5118 14118 5120 14170
rect 4874 14116 4880 14118
rect 4936 14116 4960 14118
rect 5016 14116 5040 14118
rect 5096 14116 5120 14118
rect 5176 14116 5182 14118
rect 4874 14107 5182 14116
rect 5172 14068 5224 14074
rect 5172 14010 5224 14016
rect 4802 13968 4858 13977
rect 5184 13938 5212 14010
rect 4802 13903 4858 13912
rect 5172 13932 5224 13938
rect 5172 13874 5224 13880
rect 4896 13796 4948 13802
rect 4896 13738 4948 13744
rect 4804 13524 4856 13530
rect 4804 13466 4856 13472
rect 4712 12640 4764 12646
rect 4712 12582 4764 12588
rect 4632 12406 4752 12434
rect 4620 12232 4672 12238
rect 4620 12174 4672 12180
rect 4436 12096 4488 12102
rect 4158 12064 4214 12073
rect 4436 12038 4488 12044
rect 4158 11999 4214 12008
rect 4172 11762 4200 11999
rect 4448 11898 4476 12038
rect 4436 11892 4488 11898
rect 4436 11834 4488 11840
rect 4160 11756 4212 11762
rect 4160 11698 4212 11704
rect 4632 11642 4660 12174
rect 4724 11762 4752 12406
rect 4816 12238 4844 13466
rect 4908 13394 4936 13738
rect 4896 13388 4948 13394
rect 4896 13330 4948 13336
rect 5184 13274 5212 13874
rect 5276 13530 5304 14350
rect 5460 14074 5488 14350
rect 5540 14272 5592 14278
rect 5540 14214 5592 14220
rect 5632 14272 5684 14278
rect 5632 14214 5684 14220
rect 5448 14068 5500 14074
rect 5448 14010 5500 14016
rect 5356 13728 5408 13734
rect 5356 13670 5408 13676
rect 5264 13524 5316 13530
rect 5264 13466 5316 13472
rect 5276 13394 5304 13466
rect 5264 13388 5316 13394
rect 5264 13330 5316 13336
rect 5184 13246 5304 13274
rect 4874 13084 5182 13093
rect 4874 13082 4880 13084
rect 4936 13082 4960 13084
rect 5016 13082 5040 13084
rect 5096 13082 5120 13084
rect 5176 13082 5182 13084
rect 4936 13030 4938 13082
rect 5118 13030 5120 13082
rect 4874 13028 4880 13030
rect 4936 13028 4960 13030
rect 5016 13028 5040 13030
rect 5096 13028 5120 13030
rect 5176 13028 5182 13030
rect 4874 13019 5182 13028
rect 4894 12880 4950 12889
rect 4894 12815 4950 12824
rect 4988 12844 5040 12850
rect 4908 12714 4936 12815
rect 4988 12786 5040 12792
rect 4896 12708 4948 12714
rect 4896 12650 4948 12656
rect 4804 12232 4856 12238
rect 4804 12174 4856 12180
rect 4816 11830 4844 12174
rect 4908 12170 4936 12650
rect 5000 12481 5028 12786
rect 4986 12472 5042 12481
rect 4986 12407 5042 12416
rect 5172 12436 5224 12442
rect 5276 12424 5304 13246
rect 5368 12782 5396 13670
rect 5552 12850 5580 14214
rect 5644 12850 5672 14214
rect 5724 13932 5776 13938
rect 5724 13874 5776 13880
rect 5736 12986 5764 13874
rect 5816 13728 5868 13734
rect 5816 13670 5868 13676
rect 5828 12986 5856 13670
rect 5724 12980 5776 12986
rect 5724 12922 5776 12928
rect 5816 12980 5868 12986
rect 5816 12922 5868 12928
rect 5920 12850 5948 15116
rect 6104 15042 6132 17478
rect 6276 17264 6328 17270
rect 6276 17206 6328 17212
rect 6288 16454 6316 17206
rect 7116 16998 7144 18566
rect 7380 18352 7432 18358
rect 7380 18294 7432 18300
rect 7392 17882 7420 18294
rect 7380 17876 7432 17882
rect 7380 17818 7432 17824
rect 7104 16992 7156 16998
rect 7104 16934 7156 16940
rect 6276 16448 6328 16454
rect 6276 16390 6328 16396
rect 6288 15706 6316 16390
rect 6460 16176 6512 16182
rect 6460 16118 6512 16124
rect 6276 15700 6328 15706
rect 6276 15642 6328 15648
rect 6288 15502 6316 15642
rect 6276 15496 6328 15502
rect 6276 15438 6328 15444
rect 6184 15428 6236 15434
rect 6184 15370 6236 15376
rect 6196 15162 6224 15370
rect 6368 15360 6420 15366
rect 6368 15302 6420 15308
rect 6184 15156 6236 15162
rect 6184 15098 6236 15104
rect 6000 15020 6052 15026
rect 6104 15014 6316 15042
rect 6000 14962 6052 14968
rect 6012 14278 6040 14962
rect 6288 14550 6316 15014
rect 6380 14958 6408 15302
rect 6368 14952 6420 14958
rect 6368 14894 6420 14900
rect 6276 14544 6328 14550
rect 6276 14486 6328 14492
rect 6092 14408 6144 14414
rect 6092 14350 6144 14356
rect 6184 14408 6236 14414
rect 6184 14350 6236 14356
rect 6000 14272 6052 14278
rect 6000 14214 6052 14220
rect 6012 13394 6040 14214
rect 6000 13388 6052 13394
rect 6000 13330 6052 13336
rect 5540 12844 5592 12850
rect 5540 12786 5592 12792
rect 5632 12844 5684 12850
rect 5632 12786 5684 12792
rect 5724 12844 5776 12850
rect 5724 12786 5776 12792
rect 5908 12844 5960 12850
rect 5908 12786 5960 12792
rect 5356 12776 5408 12782
rect 5356 12718 5408 12724
rect 5356 12640 5408 12646
rect 5540 12640 5592 12646
rect 5356 12582 5408 12588
rect 5460 12588 5540 12594
rect 5460 12582 5592 12588
rect 5224 12396 5304 12424
rect 5172 12378 5224 12384
rect 4896 12164 4948 12170
rect 4896 12106 4948 12112
rect 5264 12164 5316 12170
rect 5264 12106 5316 12112
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 5276 11898 5304 12106
rect 4896 11892 4948 11898
rect 4896 11834 4948 11840
rect 5264 11892 5316 11898
rect 5264 11834 5316 11840
rect 4804 11824 4856 11830
rect 4804 11766 4856 11772
rect 4712 11756 4764 11762
rect 4712 11698 4764 11704
rect 4632 11614 4752 11642
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4620 11280 4672 11286
rect 4526 11248 4582 11257
rect 4620 11222 4672 11228
rect 4526 11183 4582 11192
rect 4540 11150 4568 11183
rect 4160 11144 4212 11150
rect 4160 11086 4212 11092
rect 4528 11144 4580 11150
rect 4528 11086 4580 11092
rect 4068 10668 4120 10674
rect 4068 10610 4120 10616
rect 4172 10554 4200 11086
rect 4080 10526 4200 10554
rect 4540 10538 4568 11086
rect 4528 10532 4580 10538
rect 3976 10124 4028 10130
rect 3976 10066 4028 10072
rect 3884 9648 3936 9654
rect 3884 9590 3936 9596
rect 3700 9036 3752 9042
rect 3700 8978 3752 8984
rect 3516 8968 3568 8974
rect 3516 8910 3568 8916
rect 3424 8900 3476 8906
rect 3424 8842 3476 8848
rect 3332 8832 3384 8838
rect 3332 8774 3384 8780
rect 3148 8288 3200 8294
rect 3148 8230 3200 8236
rect 3056 7880 3108 7886
rect 3056 7822 3108 7828
rect 3068 7546 3096 7822
rect 3160 7750 3188 8230
rect 3436 7750 3464 8842
rect 3528 8498 3556 8910
rect 3896 8634 3924 9590
rect 3988 9586 4016 10066
rect 3976 9580 4028 9586
rect 3976 9522 4028 9528
rect 4080 9466 4108 10526
rect 4528 10474 4580 10480
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4528 9920 4580 9926
rect 4528 9862 4580 9868
rect 3988 9438 4108 9466
rect 4540 9466 4568 9862
rect 4632 9654 4660 11222
rect 4724 11082 4752 11614
rect 4908 11150 4936 11834
rect 5080 11824 5132 11830
rect 5080 11766 5132 11772
rect 4896 11144 4948 11150
rect 4896 11086 4948 11092
rect 4712 11076 4764 11082
rect 4712 11018 4764 11024
rect 5092 11014 5120 11766
rect 5264 11620 5316 11626
rect 5264 11562 5316 11568
rect 5276 11354 5304 11562
rect 5264 11348 5316 11354
rect 5264 11290 5316 11296
rect 4804 11008 4856 11014
rect 4804 10950 4856 10956
rect 5080 11008 5132 11014
rect 5080 10950 5132 10956
rect 4816 10690 4844 10950
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 4986 10704 5042 10713
rect 4712 10668 4764 10674
rect 4816 10662 4936 10690
rect 4712 10610 4764 10616
rect 4724 10062 4752 10610
rect 4804 10532 4856 10538
rect 4804 10474 4856 10480
rect 4712 10056 4764 10062
rect 4712 9998 4764 10004
rect 4724 9722 4752 9998
rect 4712 9716 4764 9722
rect 4712 9658 4764 9664
rect 4620 9648 4672 9654
rect 4620 9590 4672 9596
rect 4540 9438 4660 9466
rect 3988 9042 4016 9438
rect 4068 9376 4120 9382
rect 4068 9318 4120 9324
rect 4080 9178 4108 9318
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4068 9172 4120 9178
rect 4068 9114 4120 9120
rect 3976 9036 4028 9042
rect 3976 8978 4028 8984
rect 3884 8628 3936 8634
rect 3884 8570 3936 8576
rect 3988 8566 4016 8978
rect 3976 8560 4028 8566
rect 3976 8502 4028 8508
rect 3516 8492 3568 8498
rect 3516 8434 3568 8440
rect 3528 7886 3556 8434
rect 3988 7886 4016 8502
rect 4068 8356 4120 8362
rect 4068 8298 4120 8304
rect 4080 8072 4108 8298
rect 4632 8294 4660 9438
rect 4816 9178 4844 10474
rect 4908 9994 4936 10662
rect 4986 10639 4988 10648
rect 5040 10639 5042 10648
rect 4988 10610 5040 10616
rect 5264 10600 5316 10606
rect 5264 10542 5316 10548
rect 4896 9988 4948 9994
rect 4896 9930 4948 9936
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 4804 9172 4856 9178
rect 4804 9114 4856 9120
rect 4712 8628 4764 8634
rect 4712 8570 4764 8576
rect 4620 8288 4672 8294
rect 4620 8230 4672 8236
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4080 8044 4200 8072
rect 4172 7886 4200 8044
rect 3516 7880 3568 7886
rect 3976 7880 4028 7886
rect 3516 7822 3568 7828
rect 3896 7840 3976 7868
rect 3148 7744 3200 7750
rect 3148 7686 3200 7692
rect 3424 7744 3476 7750
rect 3424 7686 3476 7692
rect 2964 7540 3016 7546
rect 2964 7482 3016 7488
rect 3056 7540 3108 7546
rect 3056 7482 3108 7488
rect 3436 7002 3464 7686
rect 3148 6996 3200 7002
rect 3148 6938 3200 6944
rect 3424 6996 3476 7002
rect 3424 6938 3476 6944
rect 2872 6792 2924 6798
rect 2872 6734 2924 6740
rect 2962 6760 3018 6769
rect 2688 6724 2740 6730
rect 2962 6695 2964 6704
rect 2688 6666 2740 6672
rect 3016 6695 3018 6704
rect 2964 6666 3016 6672
rect 2504 6656 2556 6662
rect 2504 6598 2556 6604
rect 2596 6656 2648 6662
rect 2596 6598 2648 6604
rect 2700 5846 2728 6666
rect 2872 6656 2924 6662
rect 2872 6598 2924 6604
rect 2884 6254 2912 6598
rect 3160 6390 3188 6938
rect 3240 6860 3292 6866
rect 3240 6802 3292 6808
rect 3148 6384 3200 6390
rect 3148 6326 3200 6332
rect 3252 6322 3280 6802
rect 3240 6316 3292 6322
rect 3240 6258 3292 6264
rect 2872 6248 2924 6254
rect 2872 6190 2924 6196
rect 3436 6118 3464 6938
rect 3896 6798 3924 7840
rect 3976 7822 4028 7828
rect 4160 7880 4212 7886
rect 4160 7822 4212 7828
rect 4252 7744 4304 7750
rect 4252 7686 4304 7692
rect 4264 7546 4292 7686
rect 4724 7546 4752 8570
rect 4816 8430 4844 9114
rect 5276 8974 5304 10542
rect 5264 8968 5316 8974
rect 5264 8910 5316 8916
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 4804 8424 4856 8430
rect 4804 8366 4856 8372
rect 5276 7857 5304 8910
rect 5368 8634 5396 12582
rect 5460 12566 5580 12582
rect 5460 10062 5488 12566
rect 5736 12442 5764 12786
rect 5920 12594 5948 12786
rect 6012 12714 6040 13330
rect 6000 12708 6052 12714
rect 6000 12650 6052 12656
rect 5920 12566 6040 12594
rect 5724 12436 5776 12442
rect 5724 12378 5776 12384
rect 6012 12170 6040 12566
rect 6104 12238 6132 14350
rect 6196 12306 6224 14350
rect 6184 12300 6236 12306
rect 6184 12242 6236 12248
rect 6092 12232 6144 12238
rect 6092 12174 6144 12180
rect 6000 12164 6052 12170
rect 6000 12106 6052 12112
rect 5816 12096 5868 12102
rect 5816 12038 5868 12044
rect 5828 11762 5856 12038
rect 6196 11898 6224 12242
rect 6184 11892 6236 11898
rect 6184 11834 6236 11840
rect 5816 11756 5868 11762
rect 5816 11698 5868 11704
rect 5632 11688 5684 11694
rect 5632 11630 5684 11636
rect 5540 11076 5592 11082
rect 5644 11064 5672 11630
rect 5724 11348 5776 11354
rect 5724 11290 5776 11296
rect 5736 11150 5764 11290
rect 5724 11144 5776 11150
rect 5724 11086 5776 11092
rect 5592 11036 5672 11064
rect 5540 11018 5592 11024
rect 5644 10674 5672 11036
rect 5736 10742 5764 11086
rect 5828 11082 5856 11698
rect 6196 11354 6224 11834
rect 6184 11348 6236 11354
rect 6184 11290 6236 11296
rect 5816 11076 5868 11082
rect 5816 11018 5868 11024
rect 5724 10736 5776 10742
rect 5724 10678 5776 10684
rect 5632 10668 5684 10674
rect 5632 10610 5684 10616
rect 5448 10056 5500 10062
rect 5448 9998 5500 10004
rect 5460 9738 5488 9998
rect 5460 9710 5580 9738
rect 5448 9512 5500 9518
rect 5448 9454 5500 9460
rect 5356 8628 5408 8634
rect 5356 8570 5408 8576
rect 5460 8498 5488 9454
rect 5552 8974 5580 9710
rect 5540 8968 5592 8974
rect 5540 8910 5592 8916
rect 5540 8560 5592 8566
rect 5540 8502 5592 8508
rect 5448 8492 5500 8498
rect 5448 8434 5500 8440
rect 5552 8362 5580 8502
rect 5540 8356 5592 8362
rect 5540 8298 5592 8304
rect 5356 8288 5408 8294
rect 5356 8230 5408 8236
rect 5262 7848 5318 7857
rect 4804 7812 4856 7818
rect 5262 7783 5318 7792
rect 4804 7754 4856 7760
rect 4252 7540 4304 7546
rect 4252 7482 4304 7488
rect 4712 7540 4764 7546
rect 4712 7482 4764 7488
rect 4066 7440 4122 7449
rect 3976 7404 4028 7410
rect 4816 7426 4844 7754
rect 5368 7750 5396 8230
rect 5448 8016 5500 8022
rect 5448 7958 5500 7964
rect 5264 7744 5316 7750
rect 5264 7686 5316 7692
rect 5356 7744 5408 7750
rect 5356 7686 5408 7692
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 4724 7410 4844 7426
rect 4066 7375 4068 7384
rect 3976 7346 4028 7352
rect 4120 7375 4122 7384
rect 4712 7404 4844 7410
rect 4068 7346 4120 7352
rect 4764 7398 4844 7404
rect 5170 7440 5226 7449
rect 5276 7426 5304 7686
rect 5276 7410 5396 7426
rect 5276 7404 5408 7410
rect 5276 7398 5356 7404
rect 5170 7375 5226 7384
rect 4712 7346 4764 7352
rect 3884 6792 3936 6798
rect 3884 6734 3936 6740
rect 3896 6458 3924 6734
rect 3988 6662 4016 7346
rect 4620 7268 4672 7274
rect 4620 7210 4672 7216
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4632 6798 4660 7210
rect 5184 7002 5212 7375
rect 5356 7346 5408 7352
rect 4804 6996 4856 7002
rect 4804 6938 4856 6944
rect 5172 6996 5224 7002
rect 5172 6938 5224 6944
rect 4620 6792 4672 6798
rect 4620 6734 4672 6740
rect 3976 6656 4028 6662
rect 3976 6598 4028 6604
rect 3884 6452 3936 6458
rect 3884 6394 3936 6400
rect 3424 6112 3476 6118
rect 3424 6054 3476 6060
rect 3896 5914 3924 6394
rect 4068 6316 4120 6322
rect 4068 6258 4120 6264
rect 3884 5908 3936 5914
rect 3884 5850 3936 5856
rect 4080 5846 4108 6258
rect 4816 6118 4844 6938
rect 5460 6798 5488 7958
rect 5448 6792 5500 6798
rect 5354 6760 5410 6769
rect 5448 6734 5500 6740
rect 5354 6695 5356 6704
rect 5408 6695 5410 6704
rect 5356 6666 5408 6672
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 5552 6458 5580 8298
rect 5644 8022 5672 10610
rect 5736 10266 5764 10678
rect 5908 10464 5960 10470
rect 5908 10406 5960 10412
rect 5724 10260 5776 10266
rect 5724 10202 5776 10208
rect 5920 9654 5948 10406
rect 5908 9648 5960 9654
rect 5908 9590 5960 9596
rect 6288 9586 6316 14486
rect 6368 14408 6420 14414
rect 6366 14376 6368 14385
rect 6420 14376 6422 14385
rect 6366 14311 6422 14320
rect 6472 12481 6500 16118
rect 7380 16108 7432 16114
rect 7380 16050 7432 16056
rect 7196 15904 7248 15910
rect 7196 15846 7248 15852
rect 6920 15700 6972 15706
rect 6920 15642 6972 15648
rect 6552 15360 6604 15366
rect 6552 15302 6604 15308
rect 6564 13818 6592 15302
rect 6932 15162 6960 15642
rect 7208 15502 7236 15846
rect 7392 15706 7420 16050
rect 7380 15700 7432 15706
rect 7380 15642 7432 15648
rect 7196 15496 7248 15502
rect 7196 15438 7248 15444
rect 6920 15156 6972 15162
rect 6920 15098 6972 15104
rect 6932 14482 6960 15098
rect 6920 14476 6972 14482
rect 6920 14418 6972 14424
rect 7196 14476 7248 14482
rect 7196 14418 7248 14424
rect 6734 14376 6790 14385
rect 6734 14311 6790 14320
rect 6564 13802 6684 13818
rect 6564 13796 6696 13802
rect 6564 13790 6644 13796
rect 6644 13738 6696 13744
rect 6552 13184 6604 13190
rect 6552 13126 6604 13132
rect 6564 12850 6592 13126
rect 6552 12844 6604 12850
rect 6552 12786 6604 12792
rect 6458 12472 6514 12481
rect 6458 12407 6514 12416
rect 6472 11830 6500 12407
rect 6644 12096 6696 12102
rect 6748 12084 6776 14311
rect 6920 14272 6972 14278
rect 6920 14214 6972 14220
rect 6932 13938 6960 14214
rect 7104 14068 7156 14074
rect 7104 14010 7156 14016
rect 6828 13932 6880 13938
rect 6828 13874 6880 13880
rect 6920 13932 6972 13938
rect 6920 13874 6972 13880
rect 7012 13932 7064 13938
rect 7012 13874 7064 13880
rect 6840 13258 6868 13874
rect 7024 13326 7052 13874
rect 7012 13320 7064 13326
rect 7012 13262 7064 13268
rect 6828 13252 6880 13258
rect 6828 13194 6880 13200
rect 6840 12918 6868 13194
rect 6828 12912 6880 12918
rect 6828 12854 6880 12860
rect 6840 12442 6868 12854
rect 6920 12776 6972 12782
rect 6920 12718 6972 12724
rect 6828 12436 6880 12442
rect 6828 12378 6880 12384
rect 6696 12056 6776 12084
rect 6644 12038 6696 12044
rect 6460 11824 6512 11830
rect 6460 11766 6512 11772
rect 6368 9988 6420 9994
rect 6368 9930 6420 9936
rect 6380 9722 6408 9930
rect 6472 9926 6500 11766
rect 6552 11212 6604 11218
rect 6552 11154 6604 11160
rect 6460 9920 6512 9926
rect 6460 9862 6512 9868
rect 6368 9716 6420 9722
rect 6368 9658 6420 9664
rect 6276 9580 6328 9586
rect 6276 9522 6328 9528
rect 6288 9110 6316 9522
rect 6472 9518 6500 9862
rect 6460 9512 6512 9518
rect 6460 9454 6512 9460
rect 6564 9382 6592 11154
rect 6644 10056 6696 10062
rect 6644 9998 6696 10004
rect 6552 9376 6604 9382
rect 6552 9318 6604 9324
rect 6276 9104 6328 9110
rect 6276 9046 6328 9052
rect 6656 8906 6684 9998
rect 6748 9450 6776 12056
rect 6932 11558 6960 12718
rect 7024 12646 7052 13262
rect 7012 12640 7064 12646
rect 7012 12582 7064 12588
rect 7116 11762 7144 14010
rect 7208 13530 7236 14418
rect 7288 14340 7340 14346
rect 7288 14282 7340 14288
rect 7196 13524 7248 13530
rect 7196 13466 7248 13472
rect 7300 13462 7328 14282
rect 7288 13456 7340 13462
rect 7288 13398 7340 13404
rect 7484 13326 7512 26726
rect 7576 24206 7604 28358
rect 7668 26246 7696 28562
rect 7852 28218 7880 29786
rect 7944 29238 7972 30194
rect 8114 29744 8170 29753
rect 8114 29679 8116 29688
rect 8168 29679 8170 29688
rect 8116 29650 8168 29656
rect 8404 29306 8432 30670
rect 8496 30394 8524 30670
rect 8484 30388 8536 30394
rect 8484 30330 8536 30336
rect 8864 30054 8892 30670
rect 8852 30048 8904 30054
rect 8852 29990 8904 29996
rect 8864 29646 8892 29990
rect 8852 29640 8904 29646
rect 8852 29582 8904 29588
rect 8668 29504 8720 29510
rect 8668 29446 8720 29452
rect 8680 29306 8708 29446
rect 8392 29300 8444 29306
rect 8392 29242 8444 29248
rect 8668 29300 8720 29306
rect 8668 29242 8720 29248
rect 7932 29232 7984 29238
rect 7932 29174 7984 29180
rect 7840 28212 7892 28218
rect 7840 28154 7892 28160
rect 7840 28076 7892 28082
rect 7840 28018 7892 28024
rect 7852 27606 7880 28018
rect 7840 27600 7892 27606
rect 7840 27542 7892 27548
rect 7852 26246 7880 27542
rect 7944 27062 7972 29174
rect 8864 28642 8892 29582
rect 9036 29504 9088 29510
rect 9036 29446 9088 29452
rect 9048 29238 9076 29446
rect 9036 29232 9088 29238
rect 9036 29174 9088 29180
rect 8944 29164 8996 29170
rect 8944 29106 8996 29112
rect 8956 28762 8984 29106
rect 9036 28960 9088 28966
rect 9036 28902 9088 28908
rect 9048 28762 9076 28902
rect 8944 28756 8996 28762
rect 8944 28698 8996 28704
rect 9036 28756 9088 28762
rect 9036 28698 9088 28704
rect 8864 28614 8984 28642
rect 8208 28484 8260 28490
rect 8208 28426 8260 28432
rect 8220 28082 8248 28426
rect 8852 28416 8904 28422
rect 8852 28358 8904 28364
rect 8208 28076 8260 28082
rect 8208 28018 8260 28024
rect 8760 28076 8812 28082
rect 8760 28018 8812 28024
rect 8220 27130 8248 28018
rect 8772 27470 8800 28018
rect 8760 27464 8812 27470
rect 8760 27406 8812 27412
rect 8484 27328 8536 27334
rect 8484 27270 8536 27276
rect 8208 27124 8260 27130
rect 8208 27066 8260 27072
rect 7932 27056 7984 27062
rect 7932 26998 7984 27004
rect 8116 26988 8168 26994
rect 8116 26930 8168 26936
rect 8128 26586 8156 26930
rect 8116 26580 8168 26586
rect 8116 26522 8168 26528
rect 8496 26450 8524 27270
rect 8772 27130 8800 27406
rect 8760 27124 8812 27130
rect 8760 27066 8812 27072
rect 8484 26444 8536 26450
rect 8484 26386 8536 26392
rect 7932 26376 7984 26382
rect 7932 26318 7984 26324
rect 7656 26240 7708 26246
rect 7656 26182 7708 26188
rect 7840 26240 7892 26246
rect 7840 26182 7892 26188
rect 7668 25650 7696 26182
rect 7852 25906 7880 26182
rect 7944 25906 7972 26318
rect 8208 25968 8260 25974
rect 8208 25910 8260 25916
rect 7840 25900 7892 25906
rect 7840 25842 7892 25848
rect 7932 25900 7984 25906
rect 7932 25842 7984 25848
rect 7668 25622 7788 25650
rect 7654 25528 7710 25537
rect 7654 25463 7656 25472
rect 7708 25463 7710 25472
rect 7656 25434 7708 25440
rect 7668 24954 7696 25434
rect 7760 25362 7788 25622
rect 7852 25498 7880 25842
rect 7840 25492 7892 25498
rect 7840 25434 7892 25440
rect 7944 25378 7972 25842
rect 8114 25528 8170 25537
rect 8114 25463 8116 25472
rect 8168 25463 8170 25472
rect 8116 25434 8168 25440
rect 7748 25356 7800 25362
rect 7748 25298 7800 25304
rect 7852 25350 7972 25378
rect 7656 24948 7708 24954
rect 7656 24890 7708 24896
rect 7760 24614 7788 25298
rect 7852 25294 7880 25350
rect 7840 25288 7892 25294
rect 7840 25230 7892 25236
rect 8024 25288 8076 25294
rect 8024 25230 8076 25236
rect 7852 24886 7880 25230
rect 7932 25152 7984 25158
rect 7932 25094 7984 25100
rect 7840 24880 7892 24886
rect 7840 24822 7892 24828
rect 7748 24608 7800 24614
rect 7748 24550 7800 24556
rect 7564 24200 7616 24206
rect 7564 24142 7616 24148
rect 7944 22094 7972 25094
rect 8036 23322 8064 25230
rect 8128 24954 8156 25434
rect 8220 25226 8248 25910
rect 8300 25424 8352 25430
rect 8300 25366 8352 25372
rect 8208 25220 8260 25226
rect 8208 25162 8260 25168
rect 8116 24948 8168 24954
rect 8116 24890 8168 24896
rect 8024 23316 8076 23322
rect 8024 23258 8076 23264
rect 7668 22066 7972 22094
rect 7564 21956 7616 21962
rect 7564 21898 7616 21904
rect 7576 21690 7604 21898
rect 7564 21684 7616 21690
rect 7564 21626 7616 21632
rect 7564 19372 7616 19378
rect 7564 19314 7616 19320
rect 7576 17882 7604 19314
rect 7564 17876 7616 17882
rect 7564 17818 7616 17824
rect 7288 13320 7340 13326
rect 7288 13262 7340 13268
rect 7472 13320 7524 13326
rect 7472 13262 7524 13268
rect 7300 12986 7328 13262
rect 7380 13184 7432 13190
rect 7380 13126 7432 13132
rect 7288 12980 7340 12986
rect 7288 12922 7340 12928
rect 7288 12164 7340 12170
rect 7288 12106 7340 12112
rect 7104 11756 7156 11762
rect 7104 11698 7156 11704
rect 7300 11626 7328 12106
rect 7196 11620 7248 11626
rect 7196 11562 7248 11568
rect 7288 11620 7340 11626
rect 7288 11562 7340 11568
rect 6920 11552 6972 11558
rect 6920 11494 6972 11500
rect 7208 10810 7236 11562
rect 7196 10804 7248 10810
rect 7196 10746 7248 10752
rect 7208 10266 7236 10746
rect 7392 10674 7420 13126
rect 7668 12434 7696 22066
rect 7840 21956 7892 21962
rect 7840 21898 7892 21904
rect 7852 21554 7880 21898
rect 8220 21622 8248 25162
rect 8312 24750 8340 25366
rect 8864 25362 8892 28358
rect 8956 27606 8984 28614
rect 9048 28558 9076 28698
rect 9036 28552 9088 28558
rect 9036 28494 9088 28500
rect 9140 28218 9168 30670
rect 9232 29646 9260 30670
rect 9416 30598 9444 31078
rect 9692 30870 9720 31282
rect 9968 30938 9996 31282
rect 9864 30932 9916 30938
rect 9864 30874 9916 30880
rect 9956 30932 10008 30938
rect 9956 30874 10008 30880
rect 9680 30864 9732 30870
rect 9680 30806 9732 30812
rect 9496 30728 9548 30734
rect 9496 30670 9548 30676
rect 9404 30592 9456 30598
rect 9404 30534 9456 30540
rect 9416 29646 9444 30534
rect 9508 29850 9536 30670
rect 9588 30388 9640 30394
rect 9588 30330 9640 30336
rect 9496 29844 9548 29850
rect 9496 29786 9548 29792
rect 9600 29782 9628 30330
rect 9588 29776 9640 29782
rect 9588 29718 9640 29724
rect 9600 29646 9628 29718
rect 9220 29640 9272 29646
rect 9220 29582 9272 29588
rect 9404 29640 9456 29646
rect 9404 29582 9456 29588
rect 9588 29640 9640 29646
rect 9588 29582 9640 29588
rect 9232 28694 9260 29582
rect 9220 28688 9272 28694
rect 9220 28630 9272 28636
rect 9416 28490 9444 29582
rect 9600 29322 9628 29582
rect 9508 29294 9628 29322
rect 9508 28966 9536 29294
rect 9692 29186 9720 30806
rect 9772 30592 9824 30598
rect 9772 30534 9824 30540
rect 9784 29646 9812 30534
rect 9876 30394 9904 30874
rect 9956 30796 10008 30802
rect 9956 30738 10008 30744
rect 10232 30796 10284 30802
rect 10232 30738 10284 30744
rect 9864 30388 9916 30394
rect 9864 30330 9916 30336
rect 9864 30048 9916 30054
rect 9864 29990 9916 29996
rect 9876 29646 9904 29990
rect 9968 29850 9996 30738
rect 10140 30728 10192 30734
rect 10140 30670 10192 30676
rect 10152 30326 10180 30670
rect 10140 30320 10192 30326
rect 10140 30262 10192 30268
rect 10048 30252 10100 30258
rect 10048 30194 10100 30200
rect 9956 29844 10008 29850
rect 9956 29786 10008 29792
rect 9956 29708 10008 29714
rect 9956 29650 10008 29656
rect 9772 29640 9824 29646
rect 9772 29582 9824 29588
rect 9864 29640 9916 29646
rect 9864 29582 9916 29588
rect 9600 29170 9720 29186
rect 9588 29164 9720 29170
rect 9640 29158 9720 29164
rect 9588 29106 9640 29112
rect 9496 28960 9548 28966
rect 9496 28902 9548 28908
rect 9692 28490 9720 29158
rect 9404 28484 9456 28490
rect 9404 28426 9456 28432
rect 9680 28484 9732 28490
rect 9680 28426 9732 28432
rect 9128 28212 9180 28218
rect 9128 28154 9180 28160
rect 9220 28008 9272 28014
rect 9220 27950 9272 27956
rect 8944 27600 8996 27606
rect 8944 27542 8996 27548
rect 9232 26042 9260 27950
rect 9692 27470 9720 28426
rect 9968 28014 9996 29650
rect 10060 28762 10088 30194
rect 10152 29714 10180 30262
rect 10140 29708 10192 29714
rect 10140 29650 10192 29656
rect 10140 29164 10192 29170
rect 10140 29106 10192 29112
rect 10152 28762 10180 29106
rect 10048 28756 10100 28762
rect 10048 28698 10100 28704
rect 10140 28756 10192 28762
rect 10140 28698 10192 28704
rect 10244 28626 10272 30738
rect 10520 30705 10548 31726
rect 10506 30696 10562 30705
rect 10416 30660 10468 30666
rect 10506 30631 10562 30640
rect 10416 30602 10468 30608
rect 10324 30048 10376 30054
rect 10324 29990 10376 29996
rect 10336 29850 10364 29990
rect 10428 29850 10456 30602
rect 10612 30258 10640 32846
rect 10784 32768 10836 32774
rect 10784 32710 10836 32716
rect 10796 32502 10824 32710
rect 10784 32496 10836 32502
rect 10784 32438 10836 32444
rect 10784 32360 10836 32366
rect 10784 32302 10836 32308
rect 10796 31958 10824 32302
rect 10784 31952 10836 31958
rect 10784 31894 10836 31900
rect 10888 31754 10916 32846
rect 11348 32570 11376 32846
rect 11336 32564 11388 32570
rect 11336 32506 11388 32512
rect 11060 32292 11112 32298
rect 11060 32234 11112 32240
rect 10968 31952 11020 31958
rect 10968 31894 11020 31900
rect 10692 31748 10744 31754
rect 10692 31690 10744 31696
rect 10796 31726 10916 31754
rect 10704 30802 10732 31690
rect 10692 30796 10744 30802
rect 10692 30738 10744 30744
rect 10796 30433 10824 31726
rect 10782 30424 10838 30433
rect 10782 30359 10838 30368
rect 10876 30388 10928 30394
rect 10876 30330 10928 30336
rect 10784 30320 10836 30326
rect 10784 30262 10836 30268
rect 10600 30252 10652 30258
rect 10600 30194 10652 30200
rect 10692 30116 10744 30122
rect 10692 30058 10744 30064
rect 10324 29844 10376 29850
rect 10324 29786 10376 29792
rect 10416 29844 10468 29850
rect 10416 29786 10468 29792
rect 10704 29646 10732 30058
rect 10692 29640 10744 29646
rect 10692 29582 10744 29588
rect 10324 29504 10376 29510
rect 10324 29446 10376 29452
rect 10508 29504 10560 29510
rect 10508 29446 10560 29452
rect 10232 28620 10284 28626
rect 10232 28562 10284 28568
rect 9956 28008 10008 28014
rect 9956 27950 10008 27956
rect 10244 27878 10272 28562
rect 10232 27872 10284 27878
rect 10232 27814 10284 27820
rect 9680 27464 9732 27470
rect 9680 27406 9732 27412
rect 9692 27062 9720 27406
rect 10244 27130 10272 27814
rect 10232 27124 10284 27130
rect 10232 27066 10284 27072
rect 9680 27056 9732 27062
rect 9680 26998 9732 27004
rect 9588 26784 9640 26790
rect 9588 26726 9640 26732
rect 9312 26580 9364 26586
rect 9312 26522 9364 26528
rect 9220 26036 9272 26042
rect 9220 25978 9272 25984
rect 9036 25900 9088 25906
rect 9036 25842 9088 25848
rect 9048 25498 9076 25842
rect 9036 25492 9088 25498
rect 9036 25434 9088 25440
rect 8852 25356 8904 25362
rect 8852 25298 8904 25304
rect 8668 24880 8720 24886
rect 8668 24822 8720 24828
rect 8300 24744 8352 24750
rect 8300 24686 8352 24692
rect 8484 24608 8536 24614
rect 8484 24550 8536 24556
rect 8496 24206 8524 24550
rect 8484 24200 8536 24206
rect 8484 24142 8536 24148
rect 8680 23322 8708 24822
rect 8864 24410 8892 25298
rect 9232 25294 9260 25978
rect 9324 25362 9352 26522
rect 9600 26382 9628 26726
rect 9692 26382 9720 26998
rect 10244 26926 10272 27066
rect 10336 26926 10364 29446
rect 10520 28558 10548 29446
rect 10704 29238 10732 29582
rect 10692 29232 10744 29238
rect 10692 29174 10744 29180
rect 10796 29034 10824 30262
rect 10888 29306 10916 30330
rect 10980 30122 11008 31894
rect 11072 30666 11100 32234
rect 11336 32224 11388 32230
rect 11336 32166 11388 32172
rect 11348 31890 11376 32166
rect 11532 32026 11560 32846
rect 12532 32836 12584 32842
rect 13004 32842 13032 33050
rect 13556 33046 13584 34714
rect 14844 33114 14872 34714
rect 14832 33108 14884 33114
rect 14832 33050 14884 33056
rect 15292 33108 15344 33114
rect 15292 33050 15344 33056
rect 13544 33040 13596 33046
rect 13544 32982 13596 32988
rect 13924 32966 14320 32994
rect 13924 32910 13952 32966
rect 13912 32904 13964 32910
rect 13912 32846 13964 32852
rect 14292 32842 14320 32966
rect 15304 32910 15332 33050
rect 15488 32978 15516 34714
rect 16488 33108 16540 33114
rect 16488 33050 16540 33056
rect 15476 32972 15528 32978
rect 15476 32914 15528 32920
rect 14924 32904 14976 32910
rect 15292 32904 15344 32910
rect 14924 32846 14976 32852
rect 15290 32872 15292 32881
rect 15384 32904 15436 32910
rect 15344 32872 15346 32881
rect 12806 32807 12808 32816
rect 12532 32778 12584 32784
rect 12860 32807 12862 32816
rect 12992 32836 13044 32842
rect 12808 32778 12860 32784
rect 12992 32778 13044 32784
rect 13360 32836 13412 32842
rect 13360 32778 13412 32784
rect 13452 32836 13504 32842
rect 13452 32778 13504 32784
rect 14188 32836 14240 32842
rect 14188 32778 14240 32784
rect 14280 32836 14332 32842
rect 14280 32778 14332 32784
rect 14372 32836 14424 32842
rect 14372 32778 14424 32784
rect 14648 32836 14700 32842
rect 14648 32778 14700 32784
rect 12256 32768 12308 32774
rect 12544 32745 12572 32778
rect 13176 32768 13228 32774
rect 12256 32710 12308 32716
rect 12530 32736 12586 32745
rect 12072 32360 12124 32366
rect 12072 32302 12124 32308
rect 11978 32192 12034 32201
rect 11978 32127 12034 32136
rect 11520 32020 11572 32026
rect 11520 31962 11572 31968
rect 11336 31884 11388 31890
rect 11336 31826 11388 31832
rect 11532 31770 11560 31962
rect 11702 31920 11758 31929
rect 11702 31855 11758 31864
rect 11440 31742 11560 31770
rect 11244 31476 11296 31482
rect 11244 31418 11296 31424
rect 11060 30660 11112 30666
rect 11060 30602 11112 30608
rect 10968 30116 11020 30122
rect 10968 30058 11020 30064
rect 11060 30116 11112 30122
rect 11060 30058 11112 30064
rect 10876 29300 10928 29306
rect 10876 29242 10928 29248
rect 10784 29028 10836 29034
rect 10784 28970 10836 28976
rect 11072 28778 11100 30058
rect 11256 29782 11284 31418
rect 11336 30184 11388 30190
rect 11336 30126 11388 30132
rect 11244 29776 11296 29782
rect 11244 29718 11296 29724
rect 11152 29708 11204 29714
rect 11152 29650 11204 29656
rect 11164 28966 11192 29650
rect 11152 28960 11204 28966
rect 11152 28902 11204 28908
rect 11072 28750 11192 28778
rect 10508 28552 10560 28558
rect 10508 28494 10560 28500
rect 10508 28416 10560 28422
rect 10508 28358 10560 28364
rect 10520 28218 10548 28358
rect 10508 28212 10560 28218
rect 10508 28154 10560 28160
rect 11164 28014 11192 28750
rect 11242 28656 11298 28665
rect 11242 28591 11298 28600
rect 10876 28008 10928 28014
rect 10876 27950 10928 27956
rect 11152 28008 11204 28014
rect 11152 27950 11204 27956
rect 10600 27396 10652 27402
rect 10600 27338 10652 27344
rect 10232 26920 10284 26926
rect 10232 26862 10284 26868
rect 10324 26920 10376 26926
rect 10324 26862 10376 26868
rect 10244 26586 10272 26862
rect 10336 26586 10364 26862
rect 10232 26580 10284 26586
rect 10232 26522 10284 26528
rect 10324 26580 10376 26586
rect 10324 26522 10376 26528
rect 9588 26376 9640 26382
rect 9588 26318 9640 26324
rect 9680 26376 9732 26382
rect 9680 26318 9732 26324
rect 9312 25356 9364 25362
rect 9312 25298 9364 25304
rect 9220 25288 9272 25294
rect 9220 25230 9272 25236
rect 9324 24954 9352 25298
rect 9312 24948 9364 24954
rect 9312 24890 9364 24896
rect 9324 24750 9352 24890
rect 9692 24818 9720 26318
rect 9772 26308 9824 26314
rect 9772 26250 9824 26256
rect 9784 26042 9812 26250
rect 9772 26036 9824 26042
rect 9772 25978 9824 25984
rect 10416 25900 10468 25906
rect 10416 25842 10468 25848
rect 10232 25832 10284 25838
rect 10232 25774 10284 25780
rect 10140 25220 10192 25226
rect 10140 25162 10192 25168
rect 9680 24812 9732 24818
rect 9680 24754 9732 24760
rect 9312 24744 9364 24750
rect 9312 24686 9364 24692
rect 10152 24410 10180 25162
rect 10244 24410 10272 25774
rect 8852 24404 8904 24410
rect 8852 24346 8904 24352
rect 10140 24404 10192 24410
rect 10140 24346 10192 24352
rect 10232 24404 10284 24410
rect 10232 24346 10284 24352
rect 9220 24200 9272 24206
rect 9220 24142 9272 24148
rect 9864 24200 9916 24206
rect 9864 24142 9916 24148
rect 9232 23798 9260 24142
rect 9680 24064 9732 24070
rect 9680 24006 9732 24012
rect 9220 23792 9272 23798
rect 9220 23734 9272 23740
rect 9232 23662 9260 23734
rect 9220 23656 9272 23662
rect 9220 23598 9272 23604
rect 8668 23316 8720 23322
rect 8668 23258 8720 23264
rect 8300 23180 8352 23186
rect 8300 23122 8352 23128
rect 8312 22710 8340 23122
rect 8576 23112 8628 23118
rect 8576 23054 8628 23060
rect 8392 23044 8444 23050
rect 8392 22986 8444 22992
rect 8300 22704 8352 22710
rect 8300 22646 8352 22652
rect 8312 22574 8340 22646
rect 8300 22568 8352 22574
rect 8300 22510 8352 22516
rect 8208 21616 8260 21622
rect 8208 21558 8260 21564
rect 7840 21548 7892 21554
rect 7840 21490 7892 21496
rect 8312 20942 8340 22510
rect 8404 22234 8432 22986
rect 8484 22636 8536 22642
rect 8484 22578 8536 22584
rect 8496 22234 8524 22578
rect 8392 22228 8444 22234
rect 8392 22170 8444 22176
rect 8484 22228 8536 22234
rect 8484 22170 8536 22176
rect 8588 22094 8616 23054
rect 8496 22066 8616 22094
rect 8496 21146 8524 22066
rect 9128 21888 9180 21894
rect 9128 21830 9180 21836
rect 8944 21480 8996 21486
rect 8944 21422 8996 21428
rect 8668 21344 8720 21350
rect 8668 21286 8720 21292
rect 8484 21140 8536 21146
rect 8484 21082 8536 21088
rect 8300 20936 8352 20942
rect 8300 20878 8352 20884
rect 8312 20398 8340 20878
rect 8496 20466 8524 21082
rect 8484 20460 8536 20466
rect 8484 20402 8536 20408
rect 8300 20392 8352 20398
rect 8300 20334 8352 20340
rect 8392 20392 8444 20398
rect 8392 20334 8444 20340
rect 7932 20256 7984 20262
rect 7932 20198 7984 20204
rect 7944 19854 7972 20198
rect 8208 20052 8260 20058
rect 8208 19994 8260 20000
rect 7840 19848 7892 19854
rect 7840 19790 7892 19796
rect 7932 19848 7984 19854
rect 7932 19790 7984 19796
rect 7852 18714 7880 19790
rect 8116 19780 8168 19786
rect 8116 19722 8168 19728
rect 8128 19174 8156 19722
rect 8116 19168 8168 19174
rect 8116 19110 8168 19116
rect 7760 18686 7880 18714
rect 7760 18290 7788 18686
rect 7840 18624 7892 18630
rect 7840 18566 7892 18572
rect 8128 18578 8156 19110
rect 8220 18698 8248 19994
rect 8312 19310 8340 20334
rect 8404 19922 8432 20334
rect 8392 19916 8444 19922
rect 8392 19858 8444 19864
rect 8680 19854 8708 21286
rect 8956 20942 8984 21422
rect 8944 20936 8996 20942
rect 8944 20878 8996 20884
rect 8852 20868 8904 20874
rect 8852 20810 8904 20816
rect 8864 20602 8892 20810
rect 8852 20596 8904 20602
rect 8852 20538 8904 20544
rect 8760 19984 8812 19990
rect 8760 19926 8812 19932
rect 8668 19848 8720 19854
rect 8668 19790 8720 19796
rect 8392 19712 8444 19718
rect 8392 19654 8444 19660
rect 8404 19514 8432 19654
rect 8680 19530 8708 19790
rect 8392 19508 8444 19514
rect 8392 19450 8444 19456
rect 8588 19502 8708 19530
rect 8300 19304 8352 19310
rect 8300 19246 8352 19252
rect 8312 18766 8340 19246
rect 8300 18760 8352 18766
rect 8300 18702 8352 18708
rect 8208 18692 8260 18698
rect 8208 18634 8260 18640
rect 8300 18624 8352 18630
rect 8128 18572 8300 18578
rect 8128 18566 8352 18572
rect 7748 18284 7800 18290
rect 7748 18226 7800 18232
rect 7852 17678 7880 18566
rect 8128 18550 8340 18566
rect 7932 18420 7984 18426
rect 7932 18362 7984 18368
rect 7944 17678 7972 18362
rect 7840 17672 7892 17678
rect 7840 17614 7892 17620
rect 7932 17672 7984 17678
rect 7932 17614 7984 17620
rect 8116 16584 8168 16590
rect 8116 16526 8168 16532
rect 8128 15570 8156 16526
rect 8220 15706 8248 18550
rect 8404 18358 8432 19450
rect 8588 18902 8616 19502
rect 8668 19440 8720 19446
rect 8668 19382 8720 19388
rect 8576 18896 8628 18902
rect 8576 18838 8628 18844
rect 8484 18760 8536 18766
rect 8484 18702 8536 18708
rect 8496 18426 8524 18702
rect 8680 18630 8708 19382
rect 8772 19174 8800 19926
rect 8944 19848 8996 19854
rect 8944 19790 8996 19796
rect 8852 19780 8904 19786
rect 8852 19722 8904 19728
rect 8760 19168 8812 19174
rect 8760 19110 8812 19116
rect 8668 18624 8720 18630
rect 8668 18566 8720 18572
rect 8484 18420 8536 18426
rect 8484 18362 8536 18368
rect 8392 18352 8444 18358
rect 8392 18294 8444 18300
rect 8404 17762 8432 18294
rect 8772 18154 8800 19110
rect 8864 18970 8892 19722
rect 8852 18964 8904 18970
rect 8852 18906 8904 18912
rect 8760 18148 8812 18154
rect 8760 18090 8812 18096
rect 8760 17808 8812 17814
rect 8312 17734 8708 17762
rect 8760 17750 8812 17756
rect 8312 17678 8340 17734
rect 8680 17678 8708 17734
rect 8300 17672 8352 17678
rect 8300 17614 8352 17620
rect 8392 17672 8444 17678
rect 8392 17614 8444 17620
rect 8668 17672 8720 17678
rect 8668 17614 8720 17620
rect 8404 17338 8432 17614
rect 8392 17332 8444 17338
rect 8392 17274 8444 17280
rect 8680 17134 8708 17614
rect 8772 17270 8800 17750
rect 8864 17610 8892 18906
rect 8852 17604 8904 17610
rect 8852 17546 8904 17552
rect 8956 17338 8984 19790
rect 9036 18964 9088 18970
rect 9036 18906 9088 18912
rect 8944 17332 8996 17338
rect 8944 17274 8996 17280
rect 8760 17264 8812 17270
rect 8760 17206 8812 17212
rect 8668 17128 8720 17134
rect 8668 17070 8720 17076
rect 8772 16114 8800 17206
rect 9048 17082 9076 18906
rect 9140 18698 9168 21830
rect 9232 21554 9260 23598
rect 9496 23180 9548 23186
rect 9496 23122 9548 23128
rect 9508 23089 9536 23122
rect 9494 23080 9550 23089
rect 9494 23015 9550 23024
rect 9496 22976 9548 22982
rect 9496 22918 9548 22924
rect 9508 22506 9536 22918
rect 9496 22500 9548 22506
rect 9496 22442 9548 22448
rect 9692 22273 9720 24006
rect 9876 23526 9904 24142
rect 9864 23520 9916 23526
rect 9864 23462 9916 23468
rect 10244 23322 10272 24346
rect 10322 23352 10378 23361
rect 10232 23316 10284 23322
rect 10322 23287 10378 23296
rect 10232 23258 10284 23264
rect 10140 23180 10192 23186
rect 10140 23122 10192 23128
rect 9772 23112 9824 23118
rect 9772 23054 9824 23060
rect 9784 22778 9812 23054
rect 9772 22772 9824 22778
rect 9772 22714 9824 22720
rect 9864 22432 9916 22438
rect 9864 22374 9916 22380
rect 10048 22432 10100 22438
rect 10048 22374 10100 22380
rect 9678 22264 9734 22273
rect 9678 22199 9734 22208
rect 9404 22092 9456 22098
rect 9404 22034 9456 22040
rect 9312 22024 9364 22030
rect 9312 21966 9364 21972
rect 9220 21548 9272 21554
rect 9220 21490 9272 21496
rect 9324 21010 9352 21966
rect 9312 21004 9364 21010
rect 9312 20946 9364 20952
rect 9324 19990 9352 20946
rect 9416 20777 9444 22034
rect 9496 21956 9548 21962
rect 9496 21898 9548 21904
rect 9508 21350 9536 21898
rect 9876 21894 9904 22374
rect 9956 22024 10008 22030
rect 9956 21966 10008 21972
rect 9864 21888 9916 21894
rect 9864 21830 9916 21836
rect 9772 21548 9824 21554
rect 9772 21490 9824 21496
rect 9496 21344 9548 21350
rect 9496 21286 9548 21292
rect 9784 21146 9812 21490
rect 9772 21140 9824 21146
rect 9772 21082 9824 21088
rect 9968 20942 9996 21966
rect 9956 20936 10008 20942
rect 9956 20878 10008 20884
rect 9402 20768 9458 20777
rect 9402 20703 9458 20712
rect 9968 20534 9996 20878
rect 9956 20528 10008 20534
rect 9956 20470 10008 20476
rect 9312 19984 9364 19990
rect 9312 19926 9364 19932
rect 9220 19780 9272 19786
rect 9220 19722 9272 19728
rect 9128 18692 9180 18698
rect 9128 18634 9180 18640
rect 9128 18420 9180 18426
rect 9128 18362 9180 18368
rect 9140 17202 9168 18362
rect 9128 17196 9180 17202
rect 9128 17138 9180 17144
rect 9048 17054 9168 17082
rect 8944 16788 8996 16794
rect 8944 16730 8996 16736
rect 8956 16114 8984 16730
rect 9036 16516 9088 16522
rect 9036 16458 9088 16464
rect 9048 16250 9076 16458
rect 9036 16244 9088 16250
rect 9036 16186 9088 16192
rect 8760 16108 8812 16114
rect 8760 16050 8812 16056
rect 8944 16108 8996 16114
rect 8944 16050 8996 16056
rect 8208 15700 8260 15706
rect 8208 15642 8260 15648
rect 8576 15700 8628 15706
rect 8576 15642 8628 15648
rect 8116 15564 8168 15570
rect 8116 15506 8168 15512
rect 8128 15026 8156 15506
rect 8392 15496 8444 15502
rect 8392 15438 8444 15444
rect 8300 15360 8352 15366
rect 8300 15302 8352 15308
rect 8312 15162 8340 15302
rect 8300 15156 8352 15162
rect 8300 15098 8352 15104
rect 8116 15020 8168 15026
rect 8116 14962 8168 14968
rect 8024 14408 8076 14414
rect 8128 14396 8156 14962
rect 8312 14414 8340 15098
rect 8076 14368 8156 14396
rect 8300 14408 8352 14414
rect 8024 14350 8076 14356
rect 8300 14350 8352 14356
rect 8036 13938 8064 14350
rect 8404 14346 8432 15438
rect 8588 14414 8616 15642
rect 8772 15337 8800 16050
rect 8944 15904 8996 15910
rect 8944 15846 8996 15852
rect 8850 15600 8906 15609
rect 8850 15535 8852 15544
rect 8904 15535 8906 15544
rect 8852 15506 8904 15512
rect 8758 15328 8814 15337
rect 8758 15263 8814 15272
rect 8772 14550 8800 15263
rect 8956 15094 8984 15846
rect 8944 15088 8996 15094
rect 8944 15030 8996 15036
rect 8760 14544 8812 14550
rect 8760 14486 8812 14492
rect 8956 14414 8984 15030
rect 9048 14550 9076 16186
rect 9140 16114 9168 17054
rect 9128 16108 9180 16114
rect 9128 16050 9180 16056
rect 9036 14544 9088 14550
rect 9036 14486 9088 14492
rect 8576 14408 8628 14414
rect 8576 14350 8628 14356
rect 8944 14408 8996 14414
rect 8944 14350 8996 14356
rect 8392 14340 8444 14346
rect 8392 14282 8444 14288
rect 8300 14272 8352 14278
rect 8300 14214 8352 14220
rect 8116 14000 8168 14006
rect 8116 13942 8168 13948
rect 8024 13932 8076 13938
rect 8024 13874 8076 13880
rect 7748 13184 7800 13190
rect 7748 13126 7800 13132
rect 7760 12850 7788 13126
rect 8036 12850 8064 13874
rect 7748 12844 7800 12850
rect 7748 12786 7800 12792
rect 8024 12844 8076 12850
rect 8024 12786 8076 12792
rect 7668 12406 7788 12434
rect 7380 10668 7432 10674
rect 7380 10610 7432 10616
rect 7196 10260 7248 10266
rect 7196 10202 7248 10208
rect 6920 10056 6972 10062
rect 6920 9998 6972 10004
rect 6932 9722 6960 9998
rect 7392 9926 7420 10610
rect 7656 10464 7708 10470
rect 7656 10406 7708 10412
rect 7380 9920 7432 9926
rect 7380 9862 7432 9868
rect 6920 9716 6972 9722
rect 6920 9658 6972 9664
rect 6736 9444 6788 9450
rect 6736 9386 6788 9392
rect 6368 8900 6420 8906
rect 6368 8842 6420 8848
rect 6644 8900 6696 8906
rect 6644 8842 6696 8848
rect 5724 8492 5776 8498
rect 5724 8434 5776 8440
rect 6276 8492 6328 8498
rect 6276 8434 6328 8440
rect 5632 8016 5684 8022
rect 5632 7958 5684 7964
rect 5736 7886 5764 8434
rect 5908 8424 5960 8430
rect 5908 8366 5960 8372
rect 5724 7880 5776 7886
rect 5724 7822 5776 7828
rect 5724 7744 5776 7750
rect 5724 7686 5776 7692
rect 5632 7404 5684 7410
rect 5632 7346 5684 7352
rect 5644 6798 5672 7346
rect 5736 7002 5764 7686
rect 5724 6996 5776 7002
rect 5724 6938 5776 6944
rect 5632 6792 5684 6798
rect 5632 6734 5684 6740
rect 5540 6452 5592 6458
rect 5540 6394 5592 6400
rect 5644 6338 5672 6734
rect 5920 6730 5948 8366
rect 6288 8022 6316 8434
rect 6380 8362 6408 8842
rect 6748 8430 6776 9386
rect 7668 8974 7696 10406
rect 7656 8968 7708 8974
rect 7656 8910 7708 8916
rect 6736 8424 6788 8430
rect 6736 8366 6788 8372
rect 6368 8356 6420 8362
rect 6368 8298 6420 8304
rect 6276 8016 6328 8022
rect 6276 7958 6328 7964
rect 6288 7886 6316 7958
rect 6092 7880 6144 7886
rect 6276 7880 6328 7886
rect 6144 7840 6224 7868
rect 6092 7822 6144 7828
rect 6000 7744 6052 7750
rect 6000 7686 6052 7692
rect 6092 7744 6144 7750
rect 6092 7686 6144 7692
rect 6012 7426 6040 7686
rect 6104 7546 6132 7686
rect 6196 7546 6224 7840
rect 6276 7822 6328 7828
rect 6092 7540 6144 7546
rect 6092 7482 6144 7488
rect 6184 7540 6236 7546
rect 6184 7482 6236 7488
rect 6288 7426 6316 7822
rect 6012 7398 6316 7426
rect 6380 7410 6408 8298
rect 6736 7880 6788 7886
rect 6736 7822 6788 7828
rect 6748 7750 6776 7822
rect 6920 7812 6972 7818
rect 6920 7754 6972 7760
rect 6736 7744 6788 7750
rect 6736 7686 6788 7692
rect 6368 7404 6420 7410
rect 6012 7206 6040 7398
rect 6368 7346 6420 7352
rect 6000 7200 6052 7206
rect 6000 7142 6052 7148
rect 6644 7200 6696 7206
rect 6644 7142 6696 7148
rect 6184 6996 6236 7002
rect 6184 6938 6236 6944
rect 5908 6724 5960 6730
rect 5908 6666 5960 6672
rect 5552 6310 5672 6338
rect 4712 6112 4764 6118
rect 4712 6054 4764 6060
rect 4804 6112 4856 6118
rect 4804 6054 4856 6060
rect 5448 6112 5500 6118
rect 5448 6054 5500 6060
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 2688 5840 2740 5846
rect 2688 5782 2740 5788
rect 4068 5840 4120 5846
rect 4068 5782 4120 5788
rect 4724 5642 4752 6054
rect 5460 5642 5488 6054
rect 4712 5636 4764 5642
rect 4712 5578 4764 5584
rect 5448 5636 5500 5642
rect 5448 5578 5500 5584
rect 5552 5574 5580 6310
rect 6196 6186 6224 6938
rect 6656 6254 6684 7142
rect 6748 7002 6776 7686
rect 6736 6996 6788 7002
rect 6736 6938 6788 6944
rect 6748 6322 6776 6938
rect 6932 6798 6960 7754
rect 7104 7744 7156 7750
rect 7104 7686 7156 7692
rect 7012 7404 7064 7410
rect 7012 7346 7064 7352
rect 7024 7002 7052 7346
rect 7012 6996 7064 7002
rect 7012 6938 7064 6944
rect 6920 6792 6972 6798
rect 6920 6734 6972 6740
rect 6932 6458 6960 6734
rect 7116 6730 7144 7686
rect 7104 6724 7156 6730
rect 7104 6666 7156 6672
rect 6920 6452 6972 6458
rect 6920 6394 6972 6400
rect 6736 6316 6788 6322
rect 6736 6258 6788 6264
rect 6644 6248 6696 6254
rect 6644 6190 6696 6196
rect 6184 6180 6236 6186
rect 6184 6122 6236 6128
rect 6932 5914 6960 6394
rect 7760 6089 7788 12406
rect 8036 12238 8064 12786
rect 8128 12646 8156 13942
rect 8312 13938 8340 14214
rect 8300 13932 8352 13938
rect 8300 13874 8352 13880
rect 8208 13320 8260 13326
rect 8208 13262 8260 13268
rect 8300 13320 8352 13326
rect 8300 13262 8352 13268
rect 8220 12850 8248 13262
rect 8312 12986 8340 13262
rect 8300 12980 8352 12986
rect 8300 12922 8352 12928
rect 8208 12844 8260 12850
rect 8208 12786 8260 12792
rect 8208 12708 8260 12714
rect 8208 12650 8260 12656
rect 8116 12640 8168 12646
rect 8116 12582 8168 12588
rect 8220 12434 8248 12650
rect 8300 12640 8352 12646
rect 8300 12582 8352 12588
rect 8128 12406 8248 12434
rect 8024 12232 8076 12238
rect 8024 12174 8076 12180
rect 7932 11756 7984 11762
rect 8036 11744 8064 12174
rect 7984 11716 8064 11744
rect 7932 11698 7984 11704
rect 8128 11014 8156 12406
rect 8312 11830 8340 12582
rect 8300 11824 8352 11830
rect 8300 11766 8352 11772
rect 8404 11762 8432 14282
rect 8392 11756 8444 11762
rect 8392 11698 8444 11704
rect 8588 11354 8616 14350
rect 9140 14074 9168 16050
rect 9232 14958 9260 19722
rect 9324 18986 9352 19926
rect 9404 19916 9456 19922
rect 9404 19858 9456 19864
rect 9416 19174 9444 19858
rect 10060 19854 10088 22374
rect 10152 21078 10180 23122
rect 10336 22094 10364 23287
rect 10428 22642 10456 25842
rect 10612 25838 10640 27338
rect 10784 26580 10836 26586
rect 10784 26522 10836 26528
rect 10692 26308 10744 26314
rect 10692 26250 10744 26256
rect 10704 26042 10732 26250
rect 10796 26042 10824 26522
rect 10692 26036 10744 26042
rect 10692 25978 10744 25984
rect 10784 26036 10836 26042
rect 10784 25978 10836 25984
rect 10600 25832 10652 25838
rect 10600 25774 10652 25780
rect 10692 24404 10744 24410
rect 10692 24346 10744 24352
rect 10704 24274 10732 24346
rect 10600 24268 10652 24274
rect 10600 24210 10652 24216
rect 10692 24268 10744 24274
rect 10692 24210 10744 24216
rect 10612 23866 10640 24210
rect 10600 23860 10652 23866
rect 10600 23802 10652 23808
rect 10612 23730 10640 23802
rect 10508 23724 10560 23730
rect 10508 23666 10560 23672
rect 10600 23724 10652 23730
rect 10600 23666 10652 23672
rect 10520 23322 10548 23666
rect 10508 23316 10560 23322
rect 10508 23258 10560 23264
rect 10692 23112 10744 23118
rect 10692 23054 10744 23060
rect 10600 22976 10652 22982
rect 10600 22918 10652 22924
rect 10612 22642 10640 22918
rect 10416 22636 10468 22642
rect 10416 22578 10468 22584
rect 10600 22636 10652 22642
rect 10600 22578 10652 22584
rect 10508 22568 10560 22574
rect 10508 22510 10560 22516
rect 10520 22148 10548 22510
rect 10600 22160 10652 22166
rect 10520 22120 10600 22148
rect 10416 22094 10468 22098
rect 10336 22092 10468 22094
rect 10336 22066 10416 22092
rect 10416 22034 10468 22040
rect 10324 22024 10376 22030
rect 10324 21966 10376 21972
rect 10232 21956 10284 21962
rect 10232 21898 10284 21904
rect 10244 21622 10272 21898
rect 10232 21616 10284 21622
rect 10232 21558 10284 21564
rect 10140 21072 10192 21078
rect 10140 21014 10192 21020
rect 9864 19848 9916 19854
rect 9864 19790 9916 19796
rect 10048 19848 10100 19854
rect 10048 19790 10100 19796
rect 9496 19712 9548 19718
rect 9496 19654 9548 19660
rect 9508 19446 9536 19654
rect 9496 19440 9548 19446
rect 9496 19382 9548 19388
rect 9876 19334 9904 19790
rect 10060 19334 10088 19790
rect 9876 19306 9996 19334
rect 10060 19306 10180 19334
rect 9968 19174 9996 19306
rect 10048 19236 10100 19242
rect 10048 19178 10100 19184
rect 9404 19168 9456 19174
rect 9956 19168 10008 19174
rect 9456 19128 9536 19156
rect 9404 19110 9456 19116
rect 9324 18958 9444 18986
rect 9312 18692 9364 18698
rect 9312 18634 9364 18640
rect 9324 17338 9352 18634
rect 9416 18086 9444 18958
rect 9508 18766 9536 19128
rect 9956 19110 10008 19116
rect 9968 18902 9996 19110
rect 10060 18970 10088 19178
rect 10048 18964 10100 18970
rect 10048 18906 10100 18912
rect 9772 18896 9824 18902
rect 9772 18838 9824 18844
rect 9956 18896 10008 18902
rect 9956 18838 10008 18844
rect 9680 18828 9732 18834
rect 9680 18770 9732 18776
rect 9496 18760 9548 18766
rect 9496 18702 9548 18708
rect 9588 18760 9640 18766
rect 9588 18702 9640 18708
rect 9508 18170 9536 18702
rect 9600 18358 9628 18702
rect 9588 18352 9640 18358
rect 9588 18294 9640 18300
rect 9692 18290 9720 18770
rect 9784 18630 9812 18838
rect 9968 18698 9996 18838
rect 9956 18692 10008 18698
rect 9956 18634 10008 18640
rect 9772 18624 9824 18630
rect 9772 18566 9824 18572
rect 9680 18284 9732 18290
rect 9864 18284 9916 18290
rect 9732 18244 9812 18272
rect 9680 18226 9732 18232
rect 9508 18142 9628 18170
rect 9600 18086 9628 18142
rect 9404 18080 9456 18086
rect 9404 18022 9456 18028
rect 9588 18080 9640 18086
rect 9588 18022 9640 18028
rect 9312 17332 9364 17338
rect 9312 17274 9364 17280
rect 9324 16794 9352 17274
rect 9416 17202 9444 18022
rect 9404 17196 9456 17202
rect 9404 17138 9456 17144
rect 9312 16788 9364 16794
rect 9312 16730 9364 16736
rect 9404 16584 9456 16590
rect 9310 16552 9366 16561
rect 9404 16526 9456 16532
rect 9310 16487 9366 16496
rect 9324 16454 9352 16487
rect 9312 16448 9364 16454
rect 9312 16390 9364 16396
rect 9416 16250 9444 16526
rect 9496 16448 9548 16454
rect 9496 16390 9548 16396
rect 9404 16244 9456 16250
rect 9404 16186 9456 16192
rect 9416 15484 9444 16186
rect 9508 15994 9536 16390
rect 9600 16250 9628 18022
rect 9680 17128 9732 17134
rect 9680 17070 9732 17076
rect 9588 16244 9640 16250
rect 9588 16186 9640 16192
rect 9586 16144 9642 16153
rect 9692 16114 9720 17070
rect 9784 16794 9812 18244
rect 9968 18272 9996 18634
rect 10152 18426 10180 19306
rect 10140 18420 10192 18426
rect 10140 18362 10192 18368
rect 9916 18244 9996 18272
rect 9864 18226 9916 18232
rect 9864 18148 9916 18154
rect 9864 18090 9916 18096
rect 9876 17270 9904 18090
rect 9864 17264 9916 17270
rect 9864 17206 9916 17212
rect 9772 16788 9824 16794
rect 9824 16748 9904 16776
rect 9772 16730 9824 16736
rect 9772 16652 9824 16658
rect 9772 16594 9824 16600
rect 9784 16250 9812 16594
rect 9772 16244 9824 16250
rect 9772 16186 9824 16192
rect 9586 16079 9588 16088
rect 9640 16079 9642 16088
rect 9680 16108 9732 16114
rect 9588 16050 9640 16056
rect 9680 16050 9732 16056
rect 9508 15966 9720 15994
rect 9692 15706 9720 15966
rect 9784 15706 9812 16186
rect 9680 15700 9732 15706
rect 9680 15642 9732 15648
rect 9772 15700 9824 15706
rect 9772 15642 9824 15648
rect 9496 15496 9548 15502
rect 9416 15456 9496 15484
rect 9496 15438 9548 15444
rect 9312 15360 9364 15366
rect 9312 15302 9364 15308
rect 9220 14952 9272 14958
rect 9220 14894 9272 14900
rect 9232 14482 9260 14894
rect 9220 14476 9272 14482
rect 9220 14418 9272 14424
rect 9128 14068 9180 14074
rect 9128 14010 9180 14016
rect 9324 12782 9352 15302
rect 9496 14816 9548 14822
rect 9496 14758 9548 14764
rect 9508 14550 9536 14758
rect 9692 14550 9720 15642
rect 9772 15496 9824 15502
rect 9770 15464 9772 15473
rect 9824 15464 9826 15473
rect 9770 15399 9826 15408
rect 9772 15360 9824 15366
rect 9772 15302 9824 15308
rect 9496 14544 9548 14550
rect 9496 14486 9548 14492
rect 9680 14544 9732 14550
rect 9680 14486 9732 14492
rect 9508 13938 9536 14486
rect 9784 14385 9812 15302
rect 9876 15162 9904 16748
rect 9968 16590 9996 18244
rect 10244 17882 10272 21558
rect 10336 21078 10364 21966
rect 10428 21622 10456 22034
rect 10416 21616 10468 21622
rect 10416 21558 10468 21564
rect 10520 21468 10548 22120
rect 10600 22102 10652 22108
rect 10428 21440 10548 21468
rect 10324 21072 10376 21078
rect 10324 21014 10376 21020
rect 10324 20936 10376 20942
rect 10324 20878 10376 20884
rect 10336 20602 10364 20878
rect 10324 20596 10376 20602
rect 10324 20538 10376 20544
rect 10428 20466 10456 21440
rect 10600 20936 10652 20942
rect 10600 20878 10652 20884
rect 10508 20528 10560 20534
rect 10508 20470 10560 20476
rect 10416 20460 10468 20466
rect 10416 20402 10468 20408
rect 10520 19718 10548 20470
rect 10508 19712 10560 19718
rect 10508 19654 10560 19660
rect 10324 19304 10376 19310
rect 10324 19246 10376 19252
rect 10336 18970 10364 19246
rect 10324 18964 10376 18970
rect 10324 18906 10376 18912
rect 10336 18358 10364 18906
rect 10416 18760 10468 18766
rect 10416 18702 10468 18708
rect 10324 18352 10376 18358
rect 10324 18294 10376 18300
rect 10232 17876 10284 17882
rect 10232 17818 10284 17824
rect 10140 16652 10192 16658
rect 10140 16594 10192 16600
rect 9956 16584 10008 16590
rect 9956 16526 10008 16532
rect 10048 16516 10100 16522
rect 10048 16458 10100 16464
rect 9956 16448 10008 16454
rect 9956 16390 10008 16396
rect 9968 16046 9996 16390
rect 10060 16153 10088 16458
rect 10152 16182 10180 16594
rect 10140 16176 10192 16182
rect 10046 16144 10102 16153
rect 10140 16118 10192 16124
rect 10046 16079 10102 16088
rect 9956 16040 10008 16046
rect 9956 15982 10008 15988
rect 10140 16040 10192 16046
rect 10140 15982 10192 15988
rect 9956 15904 10008 15910
rect 9956 15846 10008 15852
rect 10048 15904 10100 15910
rect 10048 15846 10100 15852
rect 9968 15706 9996 15846
rect 9956 15700 10008 15706
rect 9956 15642 10008 15648
rect 9954 15600 10010 15609
rect 9954 15535 10010 15544
rect 9968 15502 9996 15535
rect 9956 15496 10008 15502
rect 9956 15438 10008 15444
rect 9864 15156 9916 15162
rect 9864 15098 9916 15104
rect 9876 14890 9904 15098
rect 9864 14884 9916 14890
rect 9864 14826 9916 14832
rect 9968 14482 9996 15438
rect 9956 14476 10008 14482
rect 9956 14418 10008 14424
rect 9770 14376 9826 14385
rect 9770 14311 9826 14320
rect 9496 13932 9548 13938
rect 9496 13874 9548 13880
rect 9680 13320 9732 13326
rect 9680 13262 9732 13268
rect 9128 12776 9180 12782
rect 9128 12718 9180 12724
rect 9312 12776 9364 12782
rect 9312 12718 9364 12724
rect 9140 12442 9168 12718
rect 9128 12436 9180 12442
rect 9128 12378 9180 12384
rect 9126 12336 9182 12345
rect 9126 12271 9182 12280
rect 9140 12238 9168 12271
rect 9128 12232 9180 12238
rect 9128 12174 9180 12180
rect 8668 12096 8720 12102
rect 8668 12038 8720 12044
rect 9036 12096 9088 12102
rect 9036 12038 9088 12044
rect 8680 11898 8708 12038
rect 8668 11892 8720 11898
rect 8668 11834 8720 11840
rect 8852 11688 8904 11694
rect 8852 11630 8904 11636
rect 8576 11348 8628 11354
rect 8576 11290 8628 11296
rect 8864 11082 8892 11630
rect 8944 11348 8996 11354
rect 8944 11290 8996 11296
rect 8852 11076 8904 11082
rect 8852 11018 8904 11024
rect 8116 11008 8168 11014
rect 8116 10950 8168 10956
rect 8760 11008 8812 11014
rect 8760 10950 8812 10956
rect 8128 10418 8156 10950
rect 8668 10736 8720 10742
rect 8668 10678 8720 10684
rect 8576 10600 8628 10606
rect 8576 10542 8628 10548
rect 8208 10532 8260 10538
rect 8208 10474 8260 10480
rect 7944 10390 8156 10418
rect 7944 10266 7972 10390
rect 7932 10260 7984 10266
rect 7932 10202 7984 10208
rect 8116 10192 8168 10198
rect 8116 10134 8168 10140
rect 8128 8566 8156 10134
rect 8116 8560 8168 8566
rect 8116 8502 8168 8508
rect 8220 7342 8248 10474
rect 8484 10464 8536 10470
rect 8484 10406 8536 10412
rect 8496 10130 8524 10406
rect 8484 10124 8536 10130
rect 8484 10066 8536 10072
rect 8588 10062 8616 10542
rect 8680 10266 8708 10678
rect 8772 10266 8800 10950
rect 8852 10600 8904 10606
rect 8852 10542 8904 10548
rect 8668 10260 8720 10266
rect 8668 10202 8720 10208
rect 8760 10260 8812 10266
rect 8760 10202 8812 10208
rect 8300 10056 8352 10062
rect 8300 9998 8352 10004
rect 8576 10056 8628 10062
rect 8576 9998 8628 10004
rect 8312 9042 8340 9998
rect 8588 9874 8616 9998
rect 8496 9846 8616 9874
rect 8392 9512 8444 9518
rect 8392 9454 8444 9460
rect 8404 9178 8432 9454
rect 8392 9172 8444 9178
rect 8392 9114 8444 9120
rect 8300 9036 8352 9042
rect 8300 8978 8352 8984
rect 8392 8900 8444 8906
rect 8392 8842 8444 8848
rect 8300 8832 8352 8838
rect 8300 8774 8352 8780
rect 8312 7410 8340 8774
rect 8404 8090 8432 8842
rect 8496 8634 8524 9846
rect 8576 9716 8628 9722
rect 8576 9658 8628 9664
rect 8588 9178 8616 9658
rect 8680 9586 8708 10202
rect 8760 9920 8812 9926
rect 8760 9862 8812 9868
rect 8668 9580 8720 9586
rect 8668 9522 8720 9528
rect 8576 9172 8628 9178
rect 8576 9114 8628 9120
rect 8484 8628 8536 8634
rect 8536 8588 8616 8616
rect 8484 8570 8536 8576
rect 8484 8492 8536 8498
rect 8484 8434 8536 8440
rect 8392 8084 8444 8090
rect 8392 8026 8444 8032
rect 8496 7546 8524 8434
rect 8588 7954 8616 8588
rect 8576 7948 8628 7954
rect 8576 7890 8628 7896
rect 8484 7540 8536 7546
rect 8484 7482 8536 7488
rect 8772 7410 8800 9862
rect 8300 7404 8352 7410
rect 8300 7346 8352 7352
rect 8760 7404 8812 7410
rect 8760 7346 8812 7352
rect 8208 7336 8260 7342
rect 8208 7278 8260 7284
rect 8668 7336 8720 7342
rect 8864 7290 8892 10542
rect 8956 8090 8984 11290
rect 9048 11082 9076 12038
rect 9312 11756 9364 11762
rect 9312 11698 9364 11704
rect 9496 11756 9548 11762
rect 9496 11698 9548 11704
rect 9220 11552 9272 11558
rect 9218 11520 9220 11529
rect 9272 11520 9274 11529
rect 9218 11455 9274 11464
rect 9128 11348 9180 11354
rect 9128 11290 9180 11296
rect 9036 11076 9088 11082
rect 9036 11018 9088 11024
rect 9140 11014 9168 11290
rect 9220 11144 9272 11150
rect 9324 11098 9352 11698
rect 9508 11150 9536 11698
rect 9692 11286 9720 13262
rect 9784 13190 9812 14311
rect 9862 13424 9918 13433
rect 9862 13359 9918 13368
rect 9876 13326 9904 13359
rect 9968 13326 9996 14418
rect 9864 13320 9916 13326
rect 9864 13262 9916 13268
rect 9956 13320 10008 13326
rect 9956 13262 10008 13268
rect 9772 13184 9824 13190
rect 9772 13126 9824 13132
rect 9784 12306 9812 13126
rect 9956 12776 10008 12782
rect 9956 12718 10008 12724
rect 9864 12708 9916 12714
rect 9864 12650 9916 12656
rect 9876 12345 9904 12650
rect 9862 12336 9918 12345
rect 9772 12300 9824 12306
rect 9862 12271 9918 12280
rect 9772 12242 9824 12248
rect 9876 11830 9904 12271
rect 9864 11824 9916 11830
rect 9864 11766 9916 11772
rect 9968 11558 9996 12718
rect 10060 12238 10088 15846
rect 10152 15502 10180 15982
rect 10140 15496 10192 15502
rect 10140 15438 10192 15444
rect 10140 14884 10192 14890
rect 10140 14826 10192 14832
rect 10152 13938 10180 14826
rect 10244 14006 10272 17818
rect 10324 17264 10376 17270
rect 10324 17206 10376 17212
rect 10336 15910 10364 17206
rect 10428 16590 10456 18702
rect 10520 18426 10548 19654
rect 10612 19242 10640 20878
rect 10704 19786 10732 23054
rect 10784 22636 10836 22642
rect 10784 22578 10836 22584
rect 10796 22234 10824 22578
rect 10784 22228 10836 22234
rect 10784 22170 10836 22176
rect 10784 21888 10836 21894
rect 10784 21830 10836 21836
rect 10796 21554 10824 21830
rect 10888 21690 10916 27950
rect 11164 27538 11192 27950
rect 11152 27532 11204 27538
rect 11152 27474 11204 27480
rect 11256 27334 11284 28591
rect 11244 27328 11296 27334
rect 11244 27270 11296 27276
rect 11244 26852 11296 26858
rect 11244 26794 11296 26800
rect 11058 26616 11114 26625
rect 11058 26551 11114 26560
rect 10968 25764 11020 25770
rect 10968 25706 11020 25712
rect 10980 24993 11008 25706
rect 11072 25498 11100 26551
rect 11060 25492 11112 25498
rect 11060 25434 11112 25440
rect 11256 25294 11284 26794
rect 11348 25362 11376 30126
rect 11440 29646 11468 31742
rect 11520 31680 11572 31686
rect 11520 31622 11572 31628
rect 11532 30394 11560 31622
rect 11520 30388 11572 30394
rect 11520 30330 11572 30336
rect 11716 29646 11744 31855
rect 11992 31226 12020 32127
rect 12084 31482 12112 32302
rect 12072 31476 12124 31482
rect 12072 31418 12124 31424
rect 11992 31198 12112 31226
rect 11888 31136 11940 31142
rect 11888 31078 11940 31084
rect 11980 31136 12032 31142
rect 11980 31078 12032 31084
rect 11900 30938 11928 31078
rect 11888 30932 11940 30938
rect 11888 30874 11940 30880
rect 11796 30660 11848 30666
rect 11796 30602 11848 30608
rect 11808 29782 11836 30602
rect 11900 30394 11928 30874
rect 11888 30388 11940 30394
rect 11888 30330 11940 30336
rect 11992 30274 12020 31078
rect 11900 30246 12020 30274
rect 11796 29776 11848 29782
rect 11796 29718 11848 29724
rect 11428 29640 11480 29646
rect 11428 29582 11480 29588
rect 11612 29640 11664 29646
rect 11612 29582 11664 29588
rect 11704 29640 11756 29646
rect 11704 29582 11756 29588
rect 11624 29481 11652 29582
rect 11610 29472 11666 29481
rect 11610 29407 11666 29416
rect 11612 29300 11664 29306
rect 11612 29242 11664 29248
rect 11520 28960 11572 28966
rect 11520 28902 11572 28908
rect 11532 28558 11560 28902
rect 11624 28558 11652 29242
rect 11520 28552 11572 28558
rect 11520 28494 11572 28500
rect 11612 28552 11664 28558
rect 11612 28494 11664 28500
rect 11624 27674 11652 28494
rect 11612 27668 11664 27674
rect 11612 27610 11664 27616
rect 11900 27538 11928 30246
rect 12084 29458 12112 31198
rect 12164 30048 12216 30054
rect 12164 29990 12216 29996
rect 12176 29646 12204 29990
rect 12268 29782 12296 32710
rect 13176 32710 13228 32716
rect 12530 32671 12586 32680
rect 12348 31340 12400 31346
rect 12348 31282 12400 31288
rect 12360 30394 12388 31282
rect 12440 30592 12492 30598
rect 12440 30534 12492 30540
rect 12348 30388 12400 30394
rect 12348 30330 12400 30336
rect 12348 30116 12400 30122
rect 12348 30058 12400 30064
rect 12256 29776 12308 29782
rect 12256 29718 12308 29724
rect 12360 29714 12388 30058
rect 12348 29708 12400 29714
rect 12348 29650 12400 29656
rect 12164 29640 12216 29646
rect 12164 29582 12216 29588
rect 12084 29430 12388 29458
rect 12256 29096 12308 29102
rect 12256 29038 12308 29044
rect 12268 28558 12296 29038
rect 12256 28552 12308 28558
rect 12256 28494 12308 28500
rect 11980 28212 12032 28218
rect 11980 28154 12032 28160
rect 11888 27532 11940 27538
rect 11888 27474 11940 27480
rect 11888 27328 11940 27334
rect 11888 27270 11940 27276
rect 11794 26344 11850 26353
rect 11794 26279 11850 26288
rect 11808 26246 11836 26279
rect 11796 26240 11848 26246
rect 11796 26182 11848 26188
rect 11704 25900 11756 25906
rect 11704 25842 11756 25848
rect 11336 25356 11388 25362
rect 11336 25298 11388 25304
rect 11244 25288 11296 25294
rect 11244 25230 11296 25236
rect 10966 24984 11022 24993
rect 11348 24954 11376 25298
rect 10966 24919 11022 24928
rect 11336 24948 11388 24954
rect 11336 24890 11388 24896
rect 11244 24812 11296 24818
rect 11244 24754 11296 24760
rect 11612 24812 11664 24818
rect 11612 24754 11664 24760
rect 11060 24336 11112 24342
rect 11060 24278 11112 24284
rect 10968 24064 11020 24070
rect 11072 24018 11100 24278
rect 11020 24012 11100 24018
rect 10968 24006 11100 24012
rect 11152 24064 11204 24070
rect 11152 24006 11204 24012
rect 10980 23990 11100 24006
rect 10968 23656 11020 23662
rect 10968 23598 11020 23604
rect 10980 23118 11008 23598
rect 11060 23520 11112 23526
rect 11060 23462 11112 23468
rect 11072 23322 11100 23462
rect 11060 23316 11112 23322
rect 11060 23258 11112 23264
rect 10968 23112 11020 23118
rect 10968 23054 11020 23060
rect 11072 22710 11100 23258
rect 11164 22982 11192 24006
rect 11256 23594 11284 24754
rect 11520 24744 11572 24750
rect 11520 24686 11572 24692
rect 11428 24608 11480 24614
rect 11428 24550 11480 24556
rect 11440 24274 11468 24550
rect 11428 24268 11480 24274
rect 11428 24210 11480 24216
rect 11336 24200 11388 24206
rect 11336 24142 11388 24148
rect 11348 24070 11376 24142
rect 11336 24064 11388 24070
rect 11336 24006 11388 24012
rect 11428 24064 11480 24070
rect 11428 24006 11480 24012
rect 11440 23848 11468 24006
rect 11348 23820 11468 23848
rect 11244 23588 11296 23594
rect 11244 23530 11296 23536
rect 11242 23488 11298 23497
rect 11242 23423 11298 23432
rect 11256 23322 11284 23423
rect 11244 23316 11296 23322
rect 11244 23258 11296 23264
rect 11348 23202 11376 23820
rect 11532 23798 11560 24686
rect 11520 23792 11572 23798
rect 11520 23734 11572 23740
rect 11428 23724 11480 23730
rect 11428 23666 11480 23672
rect 11256 23174 11376 23202
rect 11256 23118 11284 23174
rect 11244 23112 11296 23118
rect 11244 23054 11296 23060
rect 11336 23112 11388 23118
rect 11336 23054 11388 23060
rect 11152 22976 11204 22982
rect 11152 22918 11204 22924
rect 11060 22704 11112 22710
rect 11060 22646 11112 22652
rect 10968 22636 11020 22642
rect 10968 22578 11020 22584
rect 10876 21684 10928 21690
rect 10876 21626 10928 21632
rect 10784 21548 10836 21554
rect 10784 21490 10836 21496
rect 10888 21078 10916 21626
rect 10876 21072 10928 21078
rect 10876 21014 10928 21020
rect 10784 20936 10836 20942
rect 10784 20878 10836 20884
rect 10796 20058 10824 20878
rect 10980 20874 11008 22578
rect 11164 21486 11192 22918
rect 11244 21616 11296 21622
rect 11244 21558 11296 21564
rect 11152 21480 11204 21486
rect 11152 21422 11204 21428
rect 10968 20868 11020 20874
rect 10968 20810 11020 20816
rect 11060 20800 11112 20806
rect 11060 20742 11112 20748
rect 11072 20466 11100 20742
rect 11060 20460 11112 20466
rect 11060 20402 11112 20408
rect 10876 20392 10928 20398
rect 10876 20334 10928 20340
rect 10784 20052 10836 20058
rect 10784 19994 10836 20000
rect 10784 19848 10836 19854
rect 10784 19790 10836 19796
rect 10692 19780 10744 19786
rect 10692 19722 10744 19728
rect 10704 19514 10732 19722
rect 10692 19508 10744 19514
rect 10692 19450 10744 19456
rect 10692 19372 10744 19378
rect 10692 19314 10744 19320
rect 10600 19236 10652 19242
rect 10600 19178 10652 19184
rect 10600 18692 10652 18698
rect 10600 18634 10652 18640
rect 10508 18420 10560 18426
rect 10508 18362 10560 18368
rect 10520 16726 10548 18362
rect 10612 18290 10640 18634
rect 10704 18630 10732 19314
rect 10692 18624 10744 18630
rect 10692 18566 10744 18572
rect 10600 18284 10652 18290
rect 10600 18226 10652 18232
rect 10612 18086 10640 18226
rect 10692 18216 10744 18222
rect 10692 18158 10744 18164
rect 10600 18080 10652 18086
rect 10600 18022 10652 18028
rect 10704 17134 10732 18158
rect 10796 17338 10824 19790
rect 10888 19514 10916 20334
rect 11060 20324 11112 20330
rect 11060 20266 11112 20272
rect 10968 20256 11020 20262
rect 10968 20198 11020 20204
rect 10876 19508 10928 19514
rect 10876 19450 10928 19456
rect 10888 18834 10916 19450
rect 10876 18828 10928 18834
rect 10876 18770 10928 18776
rect 10980 18748 11008 20198
rect 11072 19854 11100 20266
rect 11060 19848 11112 19854
rect 11060 19790 11112 19796
rect 11060 19712 11112 19718
rect 11060 19654 11112 19660
rect 11072 19514 11100 19654
rect 11060 19508 11112 19514
rect 11060 19450 11112 19456
rect 11164 19378 11192 21422
rect 11256 20602 11284 21558
rect 11348 21486 11376 23054
rect 11440 21554 11468 23666
rect 11532 22642 11560 23734
rect 11624 23322 11652 24754
rect 11716 24206 11744 25842
rect 11900 25702 11928 27270
rect 11992 26518 12020 28154
rect 12268 28150 12296 28494
rect 12256 28144 12308 28150
rect 12256 28086 12308 28092
rect 12256 27668 12308 27674
rect 12256 27610 12308 27616
rect 12268 27130 12296 27610
rect 12256 27124 12308 27130
rect 12256 27066 12308 27072
rect 11980 26512 12032 26518
rect 12032 26460 12112 26466
rect 11980 26454 12112 26460
rect 11992 26438 12112 26454
rect 12084 25974 12112 26438
rect 12072 25968 12124 25974
rect 12072 25910 12124 25916
rect 11888 25696 11940 25702
rect 11888 25638 11940 25644
rect 11980 25356 12032 25362
rect 11980 25298 12032 25304
rect 11992 24342 12020 25298
rect 12072 25152 12124 25158
rect 12072 25094 12124 25100
rect 12164 25152 12216 25158
rect 12164 25094 12216 25100
rect 12256 25152 12308 25158
rect 12256 25094 12308 25100
rect 11980 24336 12032 24342
rect 11980 24278 12032 24284
rect 11704 24200 11756 24206
rect 11756 24160 11836 24188
rect 11704 24142 11756 24148
rect 11704 24064 11756 24070
rect 11704 24006 11756 24012
rect 11716 23497 11744 24006
rect 11702 23488 11758 23497
rect 11702 23423 11758 23432
rect 11612 23316 11664 23322
rect 11612 23258 11664 23264
rect 11612 23188 11664 23194
rect 11612 23130 11664 23136
rect 11520 22636 11572 22642
rect 11520 22578 11572 22584
rect 11532 21962 11560 22578
rect 11624 22234 11652 23130
rect 11612 22228 11664 22234
rect 11612 22170 11664 22176
rect 11716 22094 11744 23423
rect 11808 23361 11836 24160
rect 11978 24168 12034 24177
rect 11978 24103 12034 24112
rect 11992 23798 12020 24103
rect 11980 23792 12032 23798
rect 11980 23734 12032 23740
rect 11888 23724 11940 23730
rect 11888 23666 11940 23672
rect 11794 23352 11850 23361
rect 11900 23322 11928 23666
rect 11794 23287 11850 23296
rect 11888 23316 11940 23322
rect 11888 23258 11940 23264
rect 11992 23202 12020 23734
rect 12084 23730 12112 25094
rect 12176 24585 12204 25094
rect 12162 24576 12218 24585
rect 12162 24511 12218 24520
rect 12268 24410 12296 25094
rect 12360 24818 12388 29430
rect 12452 26353 12480 30534
rect 12544 29510 12572 32671
rect 12624 32292 12676 32298
rect 12624 32234 12676 32240
rect 12636 30734 12664 32234
rect 13084 31748 13136 31754
rect 13084 31690 13136 31696
rect 12992 31340 13044 31346
rect 12992 31282 13044 31288
rect 12716 30796 12768 30802
rect 12716 30738 12768 30744
rect 12624 30728 12676 30734
rect 12624 30670 12676 30676
rect 12728 30190 12756 30738
rect 12808 30660 12860 30666
rect 12808 30602 12860 30608
rect 12820 30326 12848 30602
rect 12808 30320 12860 30326
rect 12808 30262 12860 30268
rect 12716 30184 12768 30190
rect 12716 30126 12768 30132
rect 13004 29850 13032 31282
rect 13096 30666 13124 31690
rect 13084 30660 13136 30666
rect 13084 30602 13136 30608
rect 13188 30190 13216 32710
rect 13372 32570 13400 32778
rect 13464 32570 13492 32778
rect 13360 32564 13412 32570
rect 13360 32506 13412 32512
rect 13452 32564 13504 32570
rect 13452 32506 13504 32512
rect 13268 30592 13320 30598
rect 13268 30534 13320 30540
rect 13280 30394 13308 30534
rect 13268 30388 13320 30394
rect 13268 30330 13320 30336
rect 13084 30184 13136 30190
rect 13084 30126 13136 30132
rect 13176 30184 13228 30190
rect 13176 30126 13228 30132
rect 12992 29844 13044 29850
rect 12992 29786 13044 29792
rect 13096 29714 13124 30126
rect 12716 29708 12768 29714
rect 12716 29650 12768 29656
rect 13084 29708 13136 29714
rect 13084 29650 13136 29656
rect 13268 29708 13320 29714
rect 13268 29650 13320 29656
rect 12532 29504 12584 29510
rect 12532 29446 12584 29452
rect 12624 29504 12676 29510
rect 12624 29446 12676 29452
rect 12636 29238 12664 29446
rect 12624 29232 12676 29238
rect 12624 29174 12676 29180
rect 12624 28076 12676 28082
rect 12624 28018 12676 28024
rect 12636 27130 12664 28018
rect 12624 27124 12676 27130
rect 12624 27066 12676 27072
rect 12728 27010 12756 29650
rect 13280 29510 13308 29650
rect 12900 29504 12952 29510
rect 12900 29446 12952 29452
rect 13268 29504 13320 29510
rect 13268 29446 13320 29452
rect 12808 28416 12860 28422
rect 12808 28358 12860 28364
rect 12820 27538 12848 28358
rect 12808 27532 12860 27538
rect 12808 27474 12860 27480
rect 12636 26982 12756 27010
rect 12636 26926 12664 26982
rect 12624 26920 12676 26926
rect 12624 26862 12676 26868
rect 12438 26344 12494 26353
rect 12438 26279 12494 26288
rect 12636 25498 12664 26862
rect 12806 26480 12862 26489
rect 12806 26415 12862 26424
rect 12624 25492 12676 25498
rect 12624 25434 12676 25440
rect 12348 24812 12400 24818
rect 12348 24754 12400 24760
rect 12636 24750 12664 25434
rect 12624 24744 12676 24750
rect 12624 24686 12676 24692
rect 12256 24404 12308 24410
rect 12256 24346 12308 24352
rect 12164 24268 12216 24274
rect 12164 24210 12216 24216
rect 12176 24177 12204 24210
rect 12256 24200 12308 24206
rect 12162 24168 12218 24177
rect 12256 24142 12308 24148
rect 12162 24103 12218 24112
rect 12072 23724 12124 23730
rect 12072 23666 12124 23672
rect 12072 23588 12124 23594
rect 12072 23530 12124 23536
rect 12084 23322 12112 23530
rect 12072 23316 12124 23322
rect 12072 23258 12124 23264
rect 11796 23180 11848 23186
rect 11796 23122 11848 23128
rect 11900 23174 12020 23202
rect 12268 23202 12296 24142
rect 12532 24132 12584 24138
rect 12532 24074 12584 24080
rect 12544 23730 12572 24074
rect 12532 23724 12584 23730
rect 12532 23666 12584 23672
rect 12072 23180 12124 23186
rect 11808 22438 11836 23122
rect 11796 22432 11848 22438
rect 11796 22374 11848 22380
rect 11900 22166 11928 23174
rect 12268 23174 12388 23202
rect 12072 23122 12124 23128
rect 11980 23112 12032 23118
rect 11980 23054 12032 23060
rect 11992 22982 12020 23054
rect 11980 22976 12032 22982
rect 11980 22918 12032 22924
rect 12084 22817 12112 23122
rect 12256 23112 12308 23118
rect 12254 23080 12256 23089
rect 12308 23080 12310 23089
rect 12164 23044 12216 23050
rect 12254 23015 12310 23024
rect 12164 22986 12216 22992
rect 12176 22953 12204 22986
rect 12162 22944 12218 22953
rect 12162 22879 12218 22888
rect 12070 22808 12126 22817
rect 12070 22743 12126 22752
rect 12164 22772 12216 22778
rect 12164 22714 12216 22720
rect 11888 22160 11940 22166
rect 11888 22102 11940 22108
rect 11624 22066 11744 22094
rect 12072 22092 12124 22098
rect 11520 21956 11572 21962
rect 11520 21898 11572 21904
rect 11428 21548 11480 21554
rect 11428 21490 11480 21496
rect 11520 21548 11572 21554
rect 11520 21490 11572 21496
rect 11336 21480 11388 21486
rect 11336 21422 11388 21428
rect 11244 20596 11296 20602
rect 11244 20538 11296 20544
rect 11336 20528 11388 20534
rect 11336 20470 11388 20476
rect 11244 19916 11296 19922
rect 11244 19858 11296 19864
rect 11152 19372 11204 19378
rect 11152 19314 11204 19320
rect 11164 18902 11192 19314
rect 11152 18896 11204 18902
rect 11152 18838 11204 18844
rect 11256 18766 11284 19858
rect 11348 19378 11376 20470
rect 11440 19854 11468 21490
rect 11532 20924 11560 21490
rect 11624 21078 11652 22066
rect 12176 22080 12204 22714
rect 12124 22052 12204 22080
rect 12072 22034 12124 22040
rect 11704 22024 11756 22030
rect 11704 21966 11756 21972
rect 11716 21554 11744 21966
rect 11980 21956 12032 21962
rect 11980 21898 12032 21904
rect 11704 21548 11756 21554
rect 11704 21490 11756 21496
rect 11716 21146 11744 21490
rect 11992 21486 12020 21898
rect 12072 21684 12124 21690
rect 12072 21626 12124 21632
rect 11888 21480 11940 21486
rect 11808 21428 11888 21434
rect 11808 21422 11940 21428
rect 11980 21480 12032 21486
rect 11980 21422 12032 21428
rect 11808 21406 11928 21422
rect 11704 21140 11756 21146
rect 11704 21082 11756 21088
rect 11612 21072 11664 21078
rect 11612 21014 11664 21020
rect 11704 20936 11756 20942
rect 11532 20896 11704 20924
rect 11704 20878 11756 20884
rect 11520 20052 11572 20058
rect 11520 19994 11572 20000
rect 11428 19848 11480 19854
rect 11428 19790 11480 19796
rect 11428 19712 11480 19718
rect 11428 19654 11480 19660
rect 11336 19372 11388 19378
rect 11336 19314 11388 19320
rect 11060 18760 11112 18766
rect 10980 18720 11060 18748
rect 11244 18760 11296 18766
rect 11060 18702 11112 18708
rect 11164 18720 11244 18748
rect 10876 18624 10928 18630
rect 10876 18566 10928 18572
rect 10784 17332 10836 17338
rect 10784 17274 10836 17280
rect 10692 17128 10744 17134
rect 10692 17070 10744 17076
rect 10888 16794 10916 18566
rect 10968 18080 11020 18086
rect 10968 18022 11020 18028
rect 10876 16788 10928 16794
rect 10876 16730 10928 16736
rect 10508 16720 10560 16726
rect 10508 16662 10560 16668
rect 10416 16584 10468 16590
rect 10416 16526 10468 16532
rect 10784 16584 10836 16590
rect 10784 16526 10836 16532
rect 10416 16448 10468 16454
rect 10416 16390 10468 16396
rect 10600 16448 10652 16454
rect 10600 16390 10652 16396
rect 10324 15904 10376 15910
rect 10324 15846 10376 15852
rect 10428 15502 10456 16390
rect 10612 16046 10640 16390
rect 10692 16108 10744 16114
rect 10692 16050 10744 16056
rect 10600 16040 10652 16046
rect 10600 15982 10652 15988
rect 10508 15700 10560 15706
rect 10508 15642 10560 15648
rect 10520 15502 10548 15642
rect 10612 15638 10640 15982
rect 10600 15632 10652 15638
rect 10600 15574 10652 15580
rect 10324 15496 10376 15502
rect 10324 15438 10376 15444
rect 10416 15496 10468 15502
rect 10416 15438 10468 15444
rect 10508 15496 10560 15502
rect 10508 15438 10560 15444
rect 10600 15496 10652 15502
rect 10600 15438 10652 15444
rect 10336 15366 10364 15438
rect 10324 15360 10376 15366
rect 10612 15337 10640 15438
rect 10324 15302 10376 15308
rect 10598 15328 10654 15337
rect 10336 14872 10364 15302
rect 10598 15263 10654 15272
rect 10704 15162 10732 16050
rect 10796 15910 10824 16526
rect 10888 16046 10916 16730
rect 10876 16040 10928 16046
rect 10876 15982 10928 15988
rect 10784 15904 10836 15910
rect 10784 15846 10836 15852
rect 10796 15570 10824 15846
rect 10876 15632 10928 15638
rect 10876 15574 10928 15580
rect 10784 15564 10836 15570
rect 10784 15506 10836 15512
rect 10796 15162 10824 15506
rect 10888 15162 10916 15574
rect 10980 15502 11008 18022
rect 11072 16250 11100 18702
rect 11164 17066 11192 18720
rect 11244 18702 11296 18708
rect 11440 18698 11468 19654
rect 11428 18692 11480 18698
rect 11428 18634 11480 18640
rect 11532 18290 11560 19994
rect 11716 19786 11744 20878
rect 11704 19780 11756 19786
rect 11704 19722 11756 19728
rect 11612 19712 11664 19718
rect 11612 19654 11664 19660
rect 11624 19514 11652 19654
rect 11612 19508 11664 19514
rect 11612 19450 11664 19456
rect 11624 18766 11652 19450
rect 11704 19372 11756 19378
rect 11808 19360 11836 21406
rect 11888 21344 11940 21350
rect 11888 21286 11940 21292
rect 11900 20942 11928 21286
rect 11888 20936 11940 20942
rect 11888 20878 11940 20884
rect 11756 19332 11836 19360
rect 11888 19372 11940 19378
rect 11704 19314 11756 19320
rect 11888 19314 11940 19320
rect 11716 18970 11744 19314
rect 11900 18970 11928 19314
rect 11704 18964 11756 18970
rect 11704 18906 11756 18912
rect 11888 18964 11940 18970
rect 11888 18906 11940 18912
rect 11612 18760 11664 18766
rect 11612 18702 11664 18708
rect 11704 18624 11756 18630
rect 11704 18566 11756 18572
rect 11520 18284 11572 18290
rect 11440 18244 11520 18272
rect 11242 17912 11298 17921
rect 11242 17847 11298 17856
rect 11152 17060 11204 17066
rect 11152 17002 11204 17008
rect 11152 16516 11204 16522
rect 11152 16458 11204 16464
rect 11060 16244 11112 16250
rect 11060 16186 11112 16192
rect 10968 15496 11020 15502
rect 10968 15438 11020 15444
rect 11058 15464 11114 15473
rect 11058 15399 11114 15408
rect 10968 15360 11020 15366
rect 10968 15302 11020 15308
rect 10692 15156 10744 15162
rect 10692 15098 10744 15104
rect 10784 15156 10836 15162
rect 10784 15098 10836 15104
rect 10876 15156 10928 15162
rect 10876 15098 10928 15104
rect 10508 15088 10560 15094
rect 10508 15030 10560 15036
rect 10416 14884 10468 14890
rect 10336 14844 10416 14872
rect 10416 14826 10468 14832
rect 10520 14618 10548 15030
rect 10600 15020 10652 15026
rect 10600 14962 10652 14968
rect 10612 14822 10640 14962
rect 10600 14816 10652 14822
rect 10600 14758 10652 14764
rect 10508 14612 10560 14618
rect 10508 14554 10560 14560
rect 10520 14074 10548 14554
rect 10600 14544 10652 14550
rect 10600 14486 10652 14492
rect 10612 14090 10640 14486
rect 10704 14278 10732 15098
rect 10784 15020 10836 15026
rect 10784 14962 10836 14968
rect 10796 14618 10824 14962
rect 10876 14884 10928 14890
rect 10876 14826 10928 14832
rect 10784 14612 10836 14618
rect 10784 14554 10836 14560
rect 10692 14272 10744 14278
rect 10692 14214 10744 14220
rect 10888 14090 10916 14826
rect 10508 14068 10560 14074
rect 10508 14010 10560 14016
rect 10612 14062 10916 14090
rect 10232 14000 10284 14006
rect 10232 13942 10284 13948
rect 10140 13932 10192 13938
rect 10140 13874 10192 13880
rect 10048 12232 10100 12238
rect 10048 12174 10100 12180
rect 9956 11552 10008 11558
rect 9956 11494 10008 11500
rect 9680 11280 9732 11286
rect 9680 11222 9732 11228
rect 10244 11150 10272 13942
rect 10612 13938 10640 14062
rect 10600 13932 10652 13938
rect 10600 13874 10652 13880
rect 10508 13864 10560 13870
rect 10508 13806 10560 13812
rect 10520 11354 10548 13806
rect 10612 13326 10640 13874
rect 10784 13864 10836 13870
rect 10784 13806 10836 13812
rect 10600 13320 10652 13326
rect 10600 13262 10652 13268
rect 10692 13320 10744 13326
rect 10692 13262 10744 13268
rect 10704 12986 10732 13262
rect 10692 12980 10744 12986
rect 10692 12922 10744 12928
rect 10704 12442 10732 12922
rect 10796 12918 10824 13806
rect 10784 12912 10836 12918
rect 10784 12854 10836 12860
rect 10692 12436 10744 12442
rect 10692 12378 10744 12384
rect 10692 12096 10744 12102
rect 10692 12038 10744 12044
rect 10704 11778 10732 12038
rect 10796 11898 10824 12854
rect 10784 11892 10836 11898
rect 10784 11834 10836 11840
rect 10704 11750 10824 11778
rect 10508 11348 10560 11354
rect 10508 11290 10560 11296
rect 9272 11092 9352 11098
rect 9220 11086 9352 11092
rect 9496 11144 9548 11150
rect 9496 11086 9548 11092
rect 10232 11144 10284 11150
rect 10232 11086 10284 11092
rect 9232 11070 9352 11086
rect 9128 11008 9180 11014
rect 9128 10950 9180 10956
rect 9036 10668 9088 10674
rect 9036 10610 9088 10616
rect 9048 9722 9076 10610
rect 9128 10464 9180 10470
rect 9128 10406 9180 10412
rect 9140 10062 9168 10406
rect 9128 10056 9180 10062
rect 9128 9998 9180 10004
rect 9036 9716 9088 9722
rect 9036 9658 9088 9664
rect 9140 9330 9168 9998
rect 9220 9376 9272 9382
rect 9140 9324 9220 9330
rect 9140 9318 9272 9324
rect 9140 9302 9260 9318
rect 9036 8832 9088 8838
rect 9140 8820 9168 9302
rect 9088 8792 9168 8820
rect 9036 8774 9088 8780
rect 8944 8084 8996 8090
rect 8944 8026 8996 8032
rect 8720 7284 8892 7290
rect 8668 7278 8892 7284
rect 8680 7262 8892 7278
rect 8024 7200 8076 7206
rect 8024 7142 8076 7148
rect 8036 6798 8064 7142
rect 8024 6792 8076 6798
rect 8024 6734 8076 6740
rect 8864 6458 8892 7262
rect 8852 6452 8904 6458
rect 8852 6394 8904 6400
rect 7746 6080 7802 6089
rect 7746 6015 7802 6024
rect 6920 5908 6972 5914
rect 6920 5850 6972 5856
rect 5540 5568 5592 5574
rect 5540 5510 5592 5516
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 5552 3058 5580 5510
rect 8956 4826 8984 8026
rect 9128 7812 9180 7818
rect 9128 7754 9180 7760
rect 9140 6866 9168 7754
rect 9128 6860 9180 6866
rect 9128 6802 9180 6808
rect 9220 5296 9272 5302
rect 9220 5238 9272 5244
rect 8944 4820 8996 4826
rect 8944 4762 8996 4768
rect 9128 4684 9180 4690
rect 9128 4626 9180 4632
rect 8852 4616 8904 4622
rect 8852 4558 8904 4564
rect 8864 4214 8892 4558
rect 8852 4208 8904 4214
rect 8852 4150 8904 4156
rect 8758 4040 8814 4049
rect 8758 3975 8814 3984
rect 8024 3936 8076 3942
rect 8024 3878 8076 3884
rect 8036 3602 8064 3878
rect 8024 3596 8076 3602
rect 8024 3538 8076 3544
rect 8772 3534 8800 3975
rect 8760 3528 8812 3534
rect 8760 3470 8812 3476
rect 8760 3392 8812 3398
rect 8760 3334 8812 3340
rect 5540 3052 5592 3058
rect 5540 2994 5592 3000
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 8772 2446 8800 3334
rect 8864 2582 8892 4150
rect 9140 4146 9168 4626
rect 9232 4434 9260 5238
rect 9324 4622 9352 11070
rect 9404 5364 9456 5370
rect 9404 5306 9456 5312
rect 9416 4622 9444 5306
rect 9508 5302 9536 11086
rect 9772 10668 9824 10674
rect 9772 10610 9824 10616
rect 9588 9512 9640 9518
rect 9588 9454 9640 9460
rect 9600 8430 9628 9454
rect 9784 8634 9812 10610
rect 10508 10600 10560 10606
rect 10508 10542 10560 10548
rect 10520 10062 10548 10542
rect 10508 10056 10560 10062
rect 10508 9998 10560 10004
rect 9864 9580 9916 9586
rect 9864 9522 9916 9528
rect 10416 9580 10468 9586
rect 10416 9522 10468 9528
rect 9876 8906 9904 9522
rect 9864 8900 9916 8906
rect 9864 8842 9916 8848
rect 9772 8628 9824 8634
rect 9772 8570 9824 8576
rect 9588 8424 9640 8430
rect 9588 8366 9640 8372
rect 9600 7546 9628 8366
rect 9784 8294 9812 8570
rect 9876 8498 9904 8842
rect 10428 8634 10456 9522
rect 10416 8628 10468 8634
rect 10416 8570 10468 8576
rect 9864 8492 9916 8498
rect 9864 8434 9916 8440
rect 9772 8288 9824 8294
rect 9772 8230 9824 8236
rect 9784 8022 9812 8230
rect 9772 8016 9824 8022
rect 9772 7958 9824 7964
rect 9588 7540 9640 7546
rect 9588 7482 9640 7488
rect 9680 7404 9732 7410
rect 9680 7346 9732 7352
rect 9692 6322 9720 7346
rect 9784 6322 9812 7958
rect 9876 7886 9904 8434
rect 9864 7880 9916 7886
rect 9864 7822 9916 7828
rect 9876 7478 9904 7822
rect 10416 7812 10468 7818
rect 10520 7800 10548 9998
rect 10796 9382 10824 11750
rect 10980 10985 11008 15302
rect 11072 15162 11100 15399
rect 11060 15156 11112 15162
rect 11060 15098 11112 15104
rect 11072 15026 11100 15098
rect 11060 15020 11112 15026
rect 11060 14962 11112 14968
rect 11164 14498 11192 16458
rect 11072 14482 11192 14498
rect 11060 14476 11192 14482
rect 11112 14470 11192 14476
rect 11060 14418 11112 14424
rect 11072 14278 11100 14418
rect 11060 14272 11112 14278
rect 11060 14214 11112 14220
rect 11072 14074 11100 14214
rect 11060 14068 11112 14074
rect 11060 14010 11112 14016
rect 11072 13394 11100 14010
rect 11256 13938 11284 17847
rect 11440 17490 11468 18244
rect 11520 18226 11572 18232
rect 11716 17746 11744 18566
rect 11704 17740 11756 17746
rect 11704 17682 11756 17688
rect 11348 17462 11468 17490
rect 11348 16658 11376 17462
rect 11428 17332 11480 17338
rect 11428 17274 11480 17280
rect 11336 16652 11388 16658
rect 11336 16594 11388 16600
rect 11348 15978 11376 16594
rect 11440 16182 11468 17274
rect 11612 17128 11664 17134
rect 11612 17070 11664 17076
rect 11518 16688 11574 16697
rect 11518 16623 11574 16632
rect 11532 16250 11560 16623
rect 11520 16244 11572 16250
rect 11520 16186 11572 16192
rect 11428 16176 11480 16182
rect 11428 16118 11480 16124
rect 11336 15972 11388 15978
rect 11336 15914 11388 15920
rect 11336 15360 11388 15366
rect 11336 15302 11388 15308
rect 11348 14550 11376 15302
rect 11440 15178 11468 16118
rect 11520 16040 11572 16046
rect 11520 15982 11572 15988
rect 11532 15366 11560 15982
rect 11624 15434 11652 17070
rect 11796 17060 11848 17066
rect 11796 17002 11848 17008
rect 11704 16720 11756 16726
rect 11704 16662 11756 16668
rect 11716 15910 11744 16662
rect 11704 15904 11756 15910
rect 11704 15846 11756 15852
rect 11716 15638 11744 15846
rect 11704 15632 11756 15638
rect 11704 15574 11756 15580
rect 11808 15502 11836 17002
rect 11888 16448 11940 16454
rect 11888 16390 11940 16396
rect 11900 16182 11928 16390
rect 11888 16176 11940 16182
rect 11888 16118 11940 16124
rect 11900 15570 11928 16118
rect 11888 15564 11940 15570
rect 11888 15506 11940 15512
rect 11796 15496 11848 15502
rect 12084 15450 12112 21626
rect 12176 21010 12204 22052
rect 12256 22024 12308 22030
rect 12360 21978 12388 23174
rect 12440 23180 12492 23186
rect 12440 23122 12492 23128
rect 12452 22506 12480 23122
rect 12530 22944 12586 22953
rect 12636 22930 12664 24686
rect 12820 24614 12848 26415
rect 12808 24608 12860 24614
rect 12808 24550 12860 24556
rect 12820 23866 12848 24550
rect 12808 23860 12860 23866
rect 12808 23802 12860 23808
rect 12716 23724 12768 23730
rect 12716 23666 12768 23672
rect 12808 23724 12860 23730
rect 12912 23712 12940 29446
rect 13372 29238 13400 32506
rect 13464 29730 13492 32506
rect 14004 32496 14056 32502
rect 14004 32438 14056 32444
rect 13544 32428 13596 32434
rect 13544 32370 13596 32376
rect 13728 32428 13780 32434
rect 13728 32370 13780 32376
rect 13556 30326 13584 32370
rect 13740 32026 13768 32370
rect 13912 32360 13964 32366
rect 13912 32302 13964 32308
rect 13728 32020 13780 32026
rect 13728 31962 13780 31968
rect 13820 32020 13872 32026
rect 13820 31962 13872 31968
rect 13832 31929 13860 31962
rect 13818 31920 13874 31929
rect 13818 31855 13874 31864
rect 13924 31822 13952 32302
rect 13728 31816 13780 31822
rect 13728 31758 13780 31764
rect 13912 31816 13964 31822
rect 13912 31758 13964 31764
rect 13636 31680 13688 31686
rect 13636 31622 13688 31628
rect 13648 31521 13676 31622
rect 13634 31512 13690 31521
rect 13634 31447 13690 31456
rect 13740 31414 13768 31758
rect 13728 31408 13780 31414
rect 13728 31350 13780 31356
rect 13636 31340 13688 31346
rect 13636 31282 13688 31288
rect 13544 30320 13596 30326
rect 13544 30262 13596 30268
rect 13464 29702 13584 29730
rect 13556 29578 13584 29702
rect 13452 29572 13504 29578
rect 13452 29514 13504 29520
rect 13544 29572 13596 29578
rect 13544 29514 13596 29520
rect 13360 29232 13412 29238
rect 13360 29174 13412 29180
rect 13464 29034 13492 29514
rect 13452 29028 13504 29034
rect 13452 28970 13504 28976
rect 13556 28994 13584 29514
rect 13648 29510 13676 31282
rect 14016 30734 14044 32438
rect 14096 32224 14148 32230
rect 14096 32166 14148 32172
rect 14108 31346 14136 32166
rect 14200 31414 14228 32778
rect 14292 32450 14320 32778
rect 14384 32570 14412 32778
rect 14464 32768 14516 32774
rect 14464 32710 14516 32716
rect 14476 32570 14504 32710
rect 14372 32564 14424 32570
rect 14372 32506 14424 32512
rect 14464 32564 14516 32570
rect 14464 32506 14516 32512
rect 14292 32422 14412 32450
rect 14384 32337 14412 32422
rect 14464 32428 14516 32434
rect 14464 32370 14516 32376
rect 14370 32328 14426 32337
rect 14370 32263 14426 32272
rect 14372 32224 14424 32230
rect 14372 32166 14424 32172
rect 14278 31920 14334 31929
rect 14278 31855 14334 31864
rect 14292 31482 14320 31855
rect 14384 31754 14412 32166
rect 14476 31754 14504 32370
rect 14660 32366 14688 32778
rect 14832 32768 14884 32774
rect 14752 32728 14832 32756
rect 14648 32360 14700 32366
rect 14554 32328 14610 32337
rect 14648 32302 14700 32308
rect 14554 32263 14610 32272
rect 14568 31929 14596 32263
rect 14554 31920 14610 31929
rect 14554 31855 14610 31864
rect 14752 31754 14780 32728
rect 14832 32710 14884 32716
rect 14936 32502 14964 32846
rect 15384 32846 15436 32852
rect 16120 32904 16172 32910
rect 16120 32846 16172 32852
rect 15290 32807 15346 32816
rect 15292 32768 15344 32774
rect 15292 32710 15344 32716
rect 14924 32496 14976 32502
rect 14924 32438 14976 32444
rect 15016 32428 15068 32434
rect 15016 32370 15068 32376
rect 14832 32360 14884 32366
rect 14832 32302 14884 32308
rect 14922 32328 14978 32337
rect 14372 31748 14424 31754
rect 14372 31690 14424 31696
rect 14464 31748 14516 31754
rect 14464 31690 14516 31696
rect 14660 31726 14780 31754
rect 14280 31476 14332 31482
rect 14280 31418 14332 31424
rect 14188 31408 14240 31414
rect 14188 31350 14240 31356
rect 14096 31340 14148 31346
rect 14096 31282 14148 31288
rect 14004 30728 14056 30734
rect 14004 30670 14056 30676
rect 14096 30252 14148 30258
rect 14096 30194 14148 30200
rect 14108 30161 14136 30194
rect 14094 30152 14150 30161
rect 14094 30087 14150 30096
rect 14108 30054 14136 30087
rect 14096 30048 14148 30054
rect 14096 29990 14148 29996
rect 14096 29844 14148 29850
rect 14096 29786 14148 29792
rect 13728 29572 13780 29578
rect 13728 29514 13780 29520
rect 13636 29504 13688 29510
rect 13636 29446 13688 29452
rect 13648 29306 13676 29446
rect 13636 29300 13688 29306
rect 13636 29242 13688 29248
rect 13740 29102 13768 29514
rect 14108 29306 14136 29786
rect 14096 29300 14148 29306
rect 14096 29242 14148 29248
rect 13728 29096 13780 29102
rect 13728 29038 13780 29044
rect 13556 28966 13676 28994
rect 13360 28688 13412 28694
rect 13360 28630 13412 28636
rect 12992 28484 13044 28490
rect 12992 28426 13044 28432
rect 13004 28218 13032 28426
rect 12992 28212 13044 28218
rect 12992 28154 13044 28160
rect 12992 28076 13044 28082
rect 12992 28018 13044 28024
rect 13004 27713 13032 28018
rect 13084 28008 13136 28014
rect 13084 27950 13136 27956
rect 12990 27704 13046 27713
rect 12990 27639 13046 27648
rect 12992 27464 13044 27470
rect 12992 27406 13044 27412
rect 13004 25294 13032 27406
rect 12992 25288 13044 25294
rect 12992 25230 13044 25236
rect 13004 24954 13032 25230
rect 12992 24948 13044 24954
rect 12992 24890 13044 24896
rect 12992 24608 13044 24614
rect 12992 24550 13044 24556
rect 13004 24138 13032 24550
rect 12992 24132 13044 24138
rect 12992 24074 13044 24080
rect 13096 23866 13124 27950
rect 13176 27328 13228 27334
rect 13176 27270 13228 27276
rect 13188 26382 13216 27270
rect 13268 27056 13320 27062
rect 13268 26998 13320 27004
rect 13176 26376 13228 26382
rect 13176 26318 13228 26324
rect 13280 25906 13308 26998
rect 13372 26994 13400 28630
rect 13544 27872 13596 27878
rect 13544 27814 13596 27820
rect 13452 27532 13504 27538
rect 13452 27474 13504 27480
rect 13360 26988 13412 26994
rect 13464 26976 13492 27474
rect 13556 27470 13584 27814
rect 13544 27464 13596 27470
rect 13544 27406 13596 27412
rect 13464 26948 13584 26976
rect 13360 26930 13412 26936
rect 13450 26888 13506 26897
rect 13450 26823 13506 26832
rect 13464 26790 13492 26823
rect 13452 26784 13504 26790
rect 13452 26726 13504 26732
rect 13464 26246 13492 26726
rect 13360 26240 13412 26246
rect 13360 26182 13412 26188
rect 13452 26240 13504 26246
rect 13452 26182 13504 26188
rect 13372 25974 13400 26182
rect 13360 25968 13412 25974
rect 13360 25910 13412 25916
rect 13464 25906 13492 26182
rect 13268 25900 13320 25906
rect 13268 25842 13320 25848
rect 13452 25900 13504 25906
rect 13452 25842 13504 25848
rect 13176 24404 13228 24410
rect 13176 24346 13228 24352
rect 12992 23860 13044 23866
rect 12992 23802 13044 23808
rect 13084 23860 13136 23866
rect 13084 23802 13136 23808
rect 12860 23684 12940 23712
rect 12808 23666 12860 23672
rect 12728 23050 12756 23666
rect 12820 23633 12848 23666
rect 12806 23624 12862 23633
rect 12806 23559 12862 23568
rect 13004 23474 13032 23802
rect 13084 23724 13136 23730
rect 13084 23666 13136 23672
rect 12912 23446 13032 23474
rect 12808 23112 12860 23118
rect 12808 23054 12860 23060
rect 12716 23044 12768 23050
rect 12716 22986 12768 22992
rect 12586 22902 12664 22930
rect 12530 22879 12586 22888
rect 12440 22500 12492 22506
rect 12440 22442 12492 22448
rect 12438 22264 12494 22273
rect 12438 22199 12494 22208
rect 12452 22098 12480 22199
rect 12440 22092 12492 22098
rect 12440 22034 12492 22040
rect 12308 21972 12388 21978
rect 12256 21966 12388 21972
rect 12268 21950 12388 21966
rect 12268 21622 12296 21950
rect 12544 21876 12572 22879
rect 12360 21848 12572 21876
rect 12360 21690 12388 21848
rect 12348 21684 12400 21690
rect 12348 21626 12400 21632
rect 12256 21616 12308 21622
rect 12256 21558 12308 21564
rect 12348 21558 12400 21564
rect 12348 21500 12400 21506
rect 12624 21548 12676 21554
rect 12360 21298 12388 21500
rect 12624 21490 12676 21496
rect 12268 21270 12388 21298
rect 12164 21004 12216 21010
rect 12164 20946 12216 20952
rect 12176 20534 12204 20946
rect 12268 20942 12296 21270
rect 12346 21176 12402 21185
rect 12636 21146 12664 21490
rect 12346 21111 12348 21120
rect 12400 21111 12402 21120
rect 12624 21140 12676 21146
rect 12348 21082 12400 21088
rect 12624 21082 12676 21088
rect 12256 20936 12308 20942
rect 12624 20936 12676 20942
rect 12308 20896 12388 20924
rect 12256 20878 12308 20884
rect 12164 20528 12216 20534
rect 12164 20470 12216 20476
rect 12164 20392 12216 20398
rect 12164 20334 12216 20340
rect 12176 19417 12204 20334
rect 12360 20058 12388 20896
rect 12624 20878 12676 20884
rect 12440 20800 12492 20806
rect 12440 20742 12492 20748
rect 12348 20052 12400 20058
rect 12348 19994 12400 20000
rect 12256 19984 12308 19990
rect 12256 19926 12308 19932
rect 12162 19408 12218 19417
rect 12268 19378 12296 19926
rect 12348 19440 12400 19446
rect 12348 19382 12400 19388
rect 12162 19343 12164 19352
rect 12216 19343 12218 19352
rect 12256 19372 12308 19378
rect 12164 19314 12216 19320
rect 12256 19314 12308 19320
rect 12256 18760 12308 18766
rect 12256 18702 12308 18708
rect 12268 18358 12296 18702
rect 12256 18352 12308 18358
rect 12256 18294 12308 18300
rect 12164 18284 12216 18290
rect 12164 18226 12216 18232
rect 12176 17882 12204 18226
rect 12360 17882 12388 19382
rect 12164 17876 12216 17882
rect 12164 17818 12216 17824
rect 12348 17876 12400 17882
rect 12348 17818 12400 17824
rect 12256 17196 12308 17202
rect 12256 17138 12308 17144
rect 12268 16980 12296 17138
rect 12360 17134 12388 17818
rect 12348 17128 12400 17134
rect 12348 17070 12400 17076
rect 12268 16952 12388 16980
rect 12256 16108 12308 16114
rect 12256 16050 12308 16056
rect 12268 15609 12296 16050
rect 12254 15600 12310 15609
rect 12254 15535 12310 15544
rect 12360 15502 12388 16952
rect 12452 16590 12480 20742
rect 12532 19168 12584 19174
rect 12532 19110 12584 19116
rect 12544 18766 12572 19110
rect 12636 18970 12664 20878
rect 12728 19378 12756 22986
rect 12820 21078 12848 23054
rect 12808 21072 12860 21078
rect 12808 21014 12860 21020
rect 12912 20942 12940 23446
rect 12992 23180 13044 23186
rect 12992 23122 13044 23128
rect 13004 22642 13032 23122
rect 12992 22636 13044 22642
rect 12992 22578 13044 22584
rect 12992 22160 13044 22166
rect 12992 22102 13044 22108
rect 13004 22001 13032 22102
rect 12990 21992 13046 22001
rect 12990 21927 13046 21936
rect 12992 21072 13044 21078
rect 12992 21014 13044 21020
rect 12900 20936 12952 20942
rect 12900 20878 12952 20884
rect 12900 20800 12952 20806
rect 12900 20742 12952 20748
rect 12912 20466 12940 20742
rect 12900 20460 12952 20466
rect 12900 20402 12952 20408
rect 12900 19984 12952 19990
rect 12900 19926 12952 19932
rect 12716 19372 12768 19378
rect 12716 19314 12768 19320
rect 12624 18964 12676 18970
rect 12624 18906 12676 18912
rect 12532 18760 12584 18766
rect 12532 18702 12584 18708
rect 12912 17610 12940 19926
rect 12900 17604 12952 17610
rect 12900 17546 12952 17552
rect 12912 17202 12940 17546
rect 12900 17196 12952 17202
rect 12900 17138 12952 17144
rect 13004 17082 13032 21014
rect 13096 19990 13124 23666
rect 13188 23662 13216 24346
rect 13176 23656 13228 23662
rect 13176 23598 13228 23604
rect 13176 22976 13228 22982
rect 13176 22918 13228 22924
rect 13188 21010 13216 22918
rect 13280 21962 13308 25842
rect 13360 25152 13412 25158
rect 13556 25106 13584 26948
rect 13648 26450 13676 28966
rect 13728 28960 13780 28966
rect 13728 28902 13780 28908
rect 13740 28218 13768 28902
rect 13728 28212 13780 28218
rect 13728 28154 13780 28160
rect 13636 26444 13688 26450
rect 13636 26386 13688 26392
rect 13360 25094 13412 25100
rect 13372 24954 13400 25094
rect 13464 25078 13584 25106
rect 13360 24948 13412 24954
rect 13360 24890 13412 24896
rect 13464 23322 13492 25078
rect 13544 24948 13596 24954
rect 13544 24890 13596 24896
rect 13452 23316 13504 23322
rect 13452 23258 13504 23264
rect 13452 23180 13504 23186
rect 13452 23122 13504 23128
rect 13360 22976 13412 22982
rect 13360 22918 13412 22924
rect 13372 22030 13400 22918
rect 13464 22234 13492 23122
rect 13452 22228 13504 22234
rect 13452 22170 13504 22176
rect 13556 22094 13584 24890
rect 13648 24342 13676 26386
rect 13820 26376 13872 26382
rect 13818 26344 13820 26353
rect 13872 26344 13874 26353
rect 13818 26279 13874 26288
rect 13912 26308 13964 26314
rect 13912 26250 13964 26256
rect 13924 25702 13952 26250
rect 13912 25696 13964 25702
rect 13912 25638 13964 25644
rect 13820 25356 13872 25362
rect 13820 25298 13872 25304
rect 13728 24812 13780 24818
rect 13728 24754 13780 24760
rect 13636 24336 13688 24342
rect 13636 24278 13688 24284
rect 13648 24206 13676 24278
rect 13636 24200 13688 24206
rect 13636 24142 13688 24148
rect 13636 23316 13688 23322
rect 13636 23258 13688 23264
rect 13648 22234 13676 23258
rect 13636 22228 13688 22234
rect 13636 22170 13688 22176
rect 13556 22066 13676 22094
rect 13360 22024 13412 22030
rect 13360 21966 13412 21972
rect 13268 21956 13320 21962
rect 13268 21898 13320 21904
rect 13268 21344 13320 21350
rect 13268 21286 13320 21292
rect 13280 21010 13308 21286
rect 13176 21004 13228 21010
rect 13176 20946 13228 20952
rect 13268 21004 13320 21010
rect 13268 20946 13320 20952
rect 13176 20528 13228 20534
rect 13176 20470 13228 20476
rect 13084 19984 13136 19990
rect 13084 19926 13136 19932
rect 13084 19712 13136 19718
rect 13084 19654 13136 19660
rect 13096 19310 13124 19654
rect 13188 19446 13216 20470
rect 13544 19780 13596 19786
rect 13544 19722 13596 19728
rect 13176 19440 13228 19446
rect 13176 19382 13228 19388
rect 13084 19304 13136 19310
rect 13084 19246 13136 19252
rect 13268 18624 13320 18630
rect 13268 18566 13320 18572
rect 13082 18456 13138 18465
rect 13082 18391 13138 18400
rect 13096 17338 13124 18391
rect 13084 17332 13136 17338
rect 13084 17274 13136 17280
rect 13280 17202 13308 18566
rect 13360 18080 13412 18086
rect 13360 18022 13412 18028
rect 13372 17678 13400 18022
rect 13360 17672 13412 17678
rect 13360 17614 13412 17620
rect 13268 17196 13320 17202
rect 13268 17138 13320 17144
rect 12728 17054 13032 17082
rect 12624 16992 12676 16998
rect 12624 16934 12676 16940
rect 12440 16584 12492 16590
rect 12440 16526 12492 16532
rect 11796 15438 11848 15444
rect 11612 15428 11664 15434
rect 11612 15370 11664 15376
rect 11520 15360 11572 15366
rect 11520 15302 11572 15308
rect 11440 15150 11560 15178
rect 11428 15088 11480 15094
rect 11428 15030 11480 15036
rect 11336 14544 11388 14550
rect 11336 14486 11388 14492
rect 11440 14414 11468 15030
rect 11428 14408 11480 14414
rect 11428 14350 11480 14356
rect 11244 13932 11296 13938
rect 11244 13874 11296 13880
rect 11532 13462 11560 15150
rect 11624 15042 11652 15370
rect 11808 15162 11836 15438
rect 11992 15422 12112 15450
rect 12348 15496 12400 15502
rect 12452 15484 12480 16526
rect 12532 16448 12584 16454
rect 12532 16390 12584 16396
rect 12544 16046 12572 16390
rect 12532 16040 12584 16046
rect 12532 15982 12584 15988
rect 12532 15496 12584 15502
rect 12452 15456 12532 15484
rect 12348 15438 12400 15444
rect 12532 15438 12584 15444
rect 11796 15156 11848 15162
rect 11796 15098 11848 15104
rect 11794 15056 11850 15065
rect 11624 15026 11744 15042
rect 11624 15020 11756 15026
rect 11624 15014 11704 15020
rect 11794 14991 11796 15000
rect 11704 14962 11756 14968
rect 11848 14991 11850 15000
rect 11796 14962 11848 14968
rect 11612 14952 11664 14958
rect 11612 14894 11664 14900
rect 11624 14414 11652 14894
rect 11716 14482 11744 14962
rect 11992 14498 12020 15422
rect 12072 15360 12124 15366
rect 12072 15302 12124 15308
rect 12084 14958 12112 15302
rect 12360 15026 12388 15438
rect 12636 15366 12664 16934
rect 12532 15360 12584 15366
rect 12530 15328 12532 15337
rect 12624 15360 12676 15366
rect 12584 15328 12586 15337
rect 12624 15302 12676 15308
rect 12530 15263 12586 15272
rect 12348 15020 12400 15026
rect 12348 14962 12400 14968
rect 12072 14952 12124 14958
rect 12072 14894 12124 14900
rect 12440 14884 12492 14890
rect 12440 14826 12492 14832
rect 12164 14816 12216 14822
rect 12164 14758 12216 14764
rect 12348 14816 12400 14822
rect 12348 14758 12400 14764
rect 11704 14476 11756 14482
rect 11992 14470 12112 14498
rect 11704 14418 11756 14424
rect 11612 14408 11664 14414
rect 11610 14376 11612 14385
rect 11888 14408 11940 14414
rect 11664 14376 11666 14385
rect 11940 14356 12020 14362
rect 11888 14350 12020 14356
rect 11900 14334 12020 14350
rect 11610 14311 11666 14320
rect 11520 13456 11572 13462
rect 11520 13398 11572 13404
rect 11060 13388 11112 13394
rect 11060 13330 11112 13336
rect 11992 13326 12020 14334
rect 12084 13938 12112 14470
rect 12176 14346 12204 14758
rect 12164 14340 12216 14346
rect 12164 14282 12216 14288
rect 12072 13932 12124 13938
rect 12072 13874 12124 13880
rect 11980 13320 12032 13326
rect 11980 13262 12032 13268
rect 11796 13184 11848 13190
rect 11796 13126 11848 13132
rect 11520 12640 11572 12646
rect 11520 12582 11572 12588
rect 11428 12232 11480 12238
rect 11428 12174 11480 12180
rect 11440 11762 11468 12174
rect 11532 11830 11560 12582
rect 11808 12306 11836 13126
rect 11992 12306 12020 13262
rect 12084 12918 12112 13874
rect 12164 13728 12216 13734
rect 12164 13670 12216 13676
rect 12256 13728 12308 13734
rect 12256 13670 12308 13676
rect 12176 12986 12204 13670
rect 12268 13326 12296 13670
rect 12256 13320 12308 13326
rect 12256 13262 12308 13268
rect 12164 12980 12216 12986
rect 12164 12922 12216 12928
rect 12072 12912 12124 12918
rect 12072 12854 12124 12860
rect 12084 12782 12112 12854
rect 12360 12850 12388 14758
rect 12452 13870 12480 14826
rect 12440 13864 12492 13870
rect 12440 13806 12492 13812
rect 12348 12844 12400 12850
rect 12348 12786 12400 12792
rect 12636 12782 12664 15302
rect 12072 12776 12124 12782
rect 12072 12718 12124 12724
rect 12624 12776 12676 12782
rect 12624 12718 12676 12724
rect 12348 12708 12400 12714
rect 12348 12650 12400 12656
rect 12256 12640 12308 12646
rect 12256 12582 12308 12588
rect 11796 12300 11848 12306
rect 11796 12242 11848 12248
rect 11980 12300 12032 12306
rect 11980 12242 12032 12248
rect 11888 12232 11940 12238
rect 11888 12174 11940 12180
rect 11704 12096 11756 12102
rect 11704 12038 11756 12044
rect 11520 11824 11572 11830
rect 11520 11766 11572 11772
rect 11428 11756 11480 11762
rect 11428 11698 11480 11704
rect 11716 11150 11744 12038
rect 11900 11898 11928 12174
rect 12268 12170 12296 12582
rect 12256 12164 12308 12170
rect 12256 12106 12308 12112
rect 12254 12064 12310 12073
rect 12254 11999 12310 12008
rect 11888 11892 11940 11898
rect 11888 11834 11940 11840
rect 12072 11756 12124 11762
rect 12072 11698 12124 11704
rect 11704 11144 11756 11150
rect 11704 11086 11756 11092
rect 10966 10976 11022 10985
rect 10966 10911 11022 10920
rect 10968 10464 11020 10470
rect 10968 10406 11020 10412
rect 10784 9376 10836 9382
rect 10784 9318 10836 9324
rect 10796 8634 10824 9318
rect 10784 8628 10836 8634
rect 10784 8570 10836 8576
rect 10980 8430 11008 10406
rect 11428 9988 11480 9994
rect 11428 9930 11480 9936
rect 11520 9988 11572 9994
rect 11520 9930 11572 9936
rect 11440 9178 11468 9930
rect 11532 9586 11560 9930
rect 11520 9580 11572 9586
rect 11520 9522 11572 9528
rect 11428 9172 11480 9178
rect 11428 9114 11480 9120
rect 11716 8974 11744 11086
rect 12084 11082 12112 11698
rect 12072 11076 12124 11082
rect 12072 11018 12124 11024
rect 12084 10674 12112 11018
rect 12072 10668 12124 10674
rect 12072 10610 12124 10616
rect 12084 9994 12112 10610
rect 12072 9988 12124 9994
rect 12072 9930 12124 9936
rect 12070 9616 12126 9625
rect 12070 9551 12126 9560
rect 11980 9036 12032 9042
rect 11980 8978 12032 8984
rect 11704 8968 11756 8974
rect 11704 8910 11756 8916
rect 11152 8832 11204 8838
rect 11152 8774 11204 8780
rect 11888 8832 11940 8838
rect 11888 8774 11940 8780
rect 10968 8424 11020 8430
rect 10968 8366 11020 8372
rect 10692 8288 10744 8294
rect 10692 8230 10744 8236
rect 10468 7772 10548 7800
rect 10600 7812 10652 7818
rect 10416 7754 10468 7760
rect 10600 7754 10652 7760
rect 9956 7744 10008 7750
rect 9956 7686 10008 7692
rect 9864 7472 9916 7478
rect 9864 7414 9916 7420
rect 9680 6316 9732 6322
rect 9680 6258 9732 6264
rect 9772 6316 9824 6322
rect 9772 6258 9824 6264
rect 9496 5296 9548 5302
rect 9496 5238 9548 5244
rect 9496 5092 9548 5098
rect 9496 5034 9548 5040
rect 9508 4622 9536 5034
rect 9876 4622 9904 7414
rect 9968 6322 9996 7686
rect 10428 7206 10456 7754
rect 10416 7200 10468 7206
rect 10416 7142 10468 7148
rect 10048 6656 10100 6662
rect 10048 6598 10100 6604
rect 9956 6316 10008 6322
rect 9956 6258 10008 6264
rect 10060 6254 10088 6598
rect 10048 6248 10100 6254
rect 10048 6190 10100 6196
rect 9956 6112 10008 6118
rect 9956 6054 10008 6060
rect 9968 5710 9996 6054
rect 10612 5914 10640 7754
rect 10704 6798 10732 8230
rect 10784 7200 10836 7206
rect 10784 7142 10836 7148
rect 10796 6798 10824 7142
rect 10692 6792 10744 6798
rect 10692 6734 10744 6740
rect 10784 6792 10836 6798
rect 10784 6734 10836 6740
rect 10980 6458 11008 8366
rect 11060 8084 11112 8090
rect 11060 8026 11112 8032
rect 11072 6866 11100 8026
rect 11164 7410 11192 8774
rect 11900 8498 11928 8774
rect 11888 8492 11940 8498
rect 11888 8434 11940 8440
rect 11244 8288 11296 8294
rect 11244 8230 11296 8236
rect 11796 8288 11848 8294
rect 11796 8230 11848 8236
rect 11256 7886 11284 8230
rect 11704 8084 11756 8090
rect 11704 8026 11756 8032
rect 11244 7880 11296 7886
rect 11244 7822 11296 7828
rect 11336 7540 11388 7546
rect 11336 7482 11388 7488
rect 11152 7404 11204 7410
rect 11152 7346 11204 7352
rect 11060 6860 11112 6866
rect 11060 6802 11112 6808
rect 11164 6730 11192 7346
rect 11348 7002 11376 7482
rect 11612 7404 11664 7410
rect 11612 7346 11664 7352
rect 11624 7002 11652 7346
rect 11336 6996 11388 7002
rect 11256 6956 11336 6984
rect 11152 6724 11204 6730
rect 11152 6666 11204 6672
rect 11256 6458 11284 6956
rect 11336 6938 11388 6944
rect 11612 6996 11664 7002
rect 11612 6938 11664 6944
rect 10968 6452 11020 6458
rect 10968 6394 11020 6400
rect 11244 6452 11296 6458
rect 11244 6394 11296 6400
rect 11152 6316 11204 6322
rect 11152 6258 11204 6264
rect 11060 6248 11112 6254
rect 11060 6190 11112 6196
rect 10876 6112 10928 6118
rect 10876 6054 10928 6060
rect 10600 5908 10652 5914
rect 10600 5850 10652 5856
rect 10888 5710 10916 6054
rect 9956 5704 10008 5710
rect 9956 5646 10008 5652
rect 10784 5704 10836 5710
rect 10784 5646 10836 5652
rect 10876 5704 10928 5710
rect 10876 5646 10928 5652
rect 10796 5370 10824 5646
rect 10784 5364 10836 5370
rect 10784 5306 10836 5312
rect 10888 5234 10916 5646
rect 10968 5568 11020 5574
rect 10968 5510 11020 5516
rect 10876 5228 10928 5234
rect 10876 5170 10928 5176
rect 9312 4616 9364 4622
rect 9312 4558 9364 4564
rect 9404 4616 9456 4622
rect 9404 4558 9456 4564
rect 9496 4616 9548 4622
rect 9496 4558 9548 4564
rect 9864 4616 9916 4622
rect 9864 4558 9916 4564
rect 9232 4406 9352 4434
rect 9324 4214 9352 4406
rect 9312 4208 9364 4214
rect 9312 4150 9364 4156
rect 9128 4140 9180 4146
rect 9128 4082 9180 4088
rect 8944 3936 8996 3942
rect 8944 3878 8996 3884
rect 8956 3126 8984 3878
rect 9140 3466 9168 4082
rect 9220 3528 9272 3534
rect 9220 3470 9272 3476
rect 9128 3460 9180 3466
rect 9128 3402 9180 3408
rect 9232 3194 9260 3470
rect 9220 3188 9272 3194
rect 9220 3130 9272 3136
rect 8944 3120 8996 3126
rect 8944 3062 8996 3068
rect 8852 2576 8904 2582
rect 8852 2518 8904 2524
rect 9232 2446 9260 3130
rect 9324 2514 9352 4150
rect 9416 4078 9444 4558
rect 9588 4480 9640 4486
rect 9588 4422 9640 4428
rect 9600 4146 9628 4422
rect 9772 4208 9824 4214
rect 9772 4150 9824 4156
rect 9588 4140 9640 4146
rect 9588 4082 9640 4088
rect 9404 4072 9456 4078
rect 9404 4014 9456 4020
rect 9784 3738 9812 4150
rect 9876 4078 9904 4558
rect 10784 4480 10836 4486
rect 10784 4422 10836 4428
rect 10416 4140 10468 4146
rect 10416 4082 10468 4088
rect 9864 4072 9916 4078
rect 9864 4014 9916 4020
rect 9772 3732 9824 3738
rect 9772 3674 9824 3680
rect 9876 3602 9904 4014
rect 9864 3596 9916 3602
rect 9864 3538 9916 3544
rect 10428 3194 10456 4082
rect 10796 3618 10824 4422
rect 10888 3942 10916 5170
rect 10980 4282 11008 5510
rect 11072 5302 11100 6190
rect 11060 5296 11112 5302
rect 11060 5238 11112 5244
rect 11164 5030 11192 6258
rect 11256 6254 11284 6394
rect 11244 6248 11296 6254
rect 11244 6190 11296 6196
rect 11716 6118 11744 8026
rect 11808 7886 11836 8230
rect 11796 7880 11848 7886
rect 11796 7822 11848 7828
rect 11900 6662 11928 8434
rect 11888 6656 11940 6662
rect 11888 6598 11940 6604
rect 11704 6112 11756 6118
rect 11704 6054 11756 6060
rect 11242 5808 11298 5817
rect 11242 5743 11298 5752
rect 11152 5024 11204 5030
rect 11152 4966 11204 4972
rect 11164 4826 11192 4966
rect 11152 4820 11204 4826
rect 11152 4762 11204 4768
rect 10968 4276 11020 4282
rect 10968 4218 11020 4224
rect 10876 3936 10928 3942
rect 10876 3878 10928 3884
rect 10888 3738 10916 3878
rect 10876 3732 10928 3738
rect 10876 3674 10928 3680
rect 10796 3590 10916 3618
rect 10416 3188 10468 3194
rect 10416 3130 10468 3136
rect 10888 2990 10916 3590
rect 10980 2990 11008 4218
rect 11164 3466 11192 4762
rect 11256 4010 11284 5743
rect 11716 5710 11744 6054
rect 11900 5794 11928 6598
rect 11992 6458 12020 8978
rect 11980 6452 12032 6458
rect 11980 6394 12032 6400
rect 12084 5914 12112 9551
rect 12268 9382 12296 11999
rect 12360 11830 12388 12650
rect 12348 11824 12400 11830
rect 12348 11766 12400 11772
rect 12636 11370 12664 12718
rect 12728 12209 12756 17054
rect 12992 16788 13044 16794
rect 12992 16730 13044 16736
rect 12900 16448 12952 16454
rect 12900 16390 12952 16396
rect 12912 15434 12940 16390
rect 12900 15428 12952 15434
rect 12900 15370 12952 15376
rect 12912 14346 12940 15370
rect 13004 15366 13032 16730
rect 13084 16584 13136 16590
rect 13084 16526 13136 16532
rect 13268 16584 13320 16590
rect 13268 16526 13320 16532
rect 13452 16584 13504 16590
rect 13452 16526 13504 16532
rect 13096 15994 13124 16526
rect 13280 16289 13308 16526
rect 13360 16448 13412 16454
rect 13360 16390 13412 16396
rect 13266 16280 13322 16289
rect 13266 16215 13322 16224
rect 13268 16108 13320 16114
rect 13268 16050 13320 16056
rect 13096 15966 13216 15994
rect 13188 15910 13216 15966
rect 13176 15904 13228 15910
rect 13176 15846 13228 15852
rect 13280 15434 13308 16050
rect 13372 15434 13400 16390
rect 13464 16182 13492 16526
rect 13452 16176 13504 16182
rect 13452 16118 13504 16124
rect 13452 16040 13504 16046
rect 13452 15982 13504 15988
rect 13268 15428 13320 15434
rect 13268 15370 13320 15376
rect 13360 15428 13412 15434
rect 13360 15370 13412 15376
rect 12992 15360 13044 15366
rect 12992 15302 13044 15308
rect 12900 14340 12952 14346
rect 12900 14282 12952 14288
rect 12808 14272 12860 14278
rect 12808 14214 12860 14220
rect 12820 14074 12848 14214
rect 12808 14068 12860 14074
rect 12808 14010 12860 14016
rect 13004 13530 13032 15302
rect 13268 14952 13320 14958
rect 13268 14894 13320 14900
rect 13280 14278 13308 14894
rect 13372 14482 13400 15370
rect 13360 14476 13412 14482
rect 13360 14418 13412 14424
rect 13268 14272 13320 14278
rect 13268 14214 13320 14220
rect 13360 14272 13412 14278
rect 13464 14260 13492 15982
rect 13412 14232 13492 14260
rect 13360 14214 13412 14220
rect 13280 14006 13308 14214
rect 13268 14000 13320 14006
rect 13268 13942 13320 13948
rect 12992 13524 13044 13530
rect 12992 13466 13044 13472
rect 12714 12200 12770 12209
rect 12714 12135 12770 12144
rect 12636 11342 12848 11370
rect 12716 11008 12768 11014
rect 12716 10950 12768 10956
rect 12440 9920 12492 9926
rect 12440 9862 12492 9868
rect 12452 9654 12480 9862
rect 12440 9648 12492 9654
rect 12440 9590 12492 9596
rect 12256 9376 12308 9382
rect 12256 9318 12308 9324
rect 12256 9104 12308 9110
rect 12256 9046 12308 9052
rect 12164 9036 12216 9042
rect 12164 8978 12216 8984
rect 12176 8090 12204 8978
rect 12164 8084 12216 8090
rect 12164 8026 12216 8032
rect 12164 7812 12216 7818
rect 12164 7754 12216 7760
rect 12176 6866 12204 7754
rect 12164 6860 12216 6866
rect 12164 6802 12216 6808
rect 12072 5908 12124 5914
rect 12072 5850 12124 5856
rect 11900 5766 12112 5794
rect 11704 5704 11756 5710
rect 11704 5646 11756 5652
rect 11520 5568 11572 5574
rect 11520 5510 11572 5516
rect 11428 4616 11480 4622
rect 11428 4558 11480 4564
rect 11244 4004 11296 4010
rect 11244 3946 11296 3952
rect 11152 3460 11204 3466
rect 11152 3402 11204 3408
rect 11256 3194 11284 3946
rect 11440 3602 11468 4558
rect 11428 3596 11480 3602
rect 11428 3538 11480 3544
rect 11532 3466 11560 5510
rect 11716 5234 11744 5646
rect 11978 5400 12034 5409
rect 11978 5335 11980 5344
rect 12032 5335 12034 5344
rect 11980 5306 12032 5312
rect 11704 5228 11756 5234
rect 11704 5170 11756 5176
rect 12084 5166 12112 5766
rect 12268 5710 12296 9046
rect 12452 8906 12480 9590
rect 12624 9580 12676 9586
rect 12624 9522 12676 9528
rect 12440 8900 12492 8906
rect 12440 8842 12492 8848
rect 12532 8900 12584 8906
rect 12532 8842 12584 8848
rect 12348 8832 12400 8838
rect 12348 8774 12400 8780
rect 12360 8430 12388 8774
rect 12348 8424 12400 8430
rect 12348 8366 12400 8372
rect 12544 7954 12572 8842
rect 12636 8634 12664 9522
rect 12624 8628 12676 8634
rect 12624 8570 12676 8576
rect 12728 8514 12756 10950
rect 12820 8566 12848 11342
rect 13268 11348 13320 11354
rect 13372 11336 13400 14214
rect 13556 12714 13584 19722
rect 13648 17678 13676 22066
rect 13740 21146 13768 24754
rect 13832 24274 13860 25298
rect 14108 25294 14136 29242
rect 14200 25702 14228 31350
rect 14556 30864 14608 30870
rect 14556 30806 14608 30812
rect 14372 30728 14424 30734
rect 14372 30670 14424 30676
rect 14280 30660 14332 30666
rect 14280 30602 14332 30608
rect 14292 30258 14320 30602
rect 14280 30252 14332 30258
rect 14280 30194 14332 30200
rect 14292 29594 14320 30194
rect 14384 29714 14412 30670
rect 14568 30258 14596 30806
rect 14660 30734 14688 31726
rect 14844 30818 14872 32302
rect 14922 32263 14978 32272
rect 14936 32230 14964 32263
rect 14924 32224 14976 32230
rect 14924 32166 14976 32172
rect 14924 31816 14976 31822
rect 14924 31758 14976 31764
rect 14752 30790 14872 30818
rect 14648 30728 14700 30734
rect 14648 30670 14700 30676
rect 14556 30252 14608 30258
rect 14556 30194 14608 30200
rect 14464 30184 14516 30190
rect 14464 30126 14516 30132
rect 14372 29708 14424 29714
rect 14372 29650 14424 29656
rect 14292 29566 14412 29594
rect 14280 29504 14332 29510
rect 14280 29446 14332 29452
rect 14292 28558 14320 29446
rect 14384 28558 14412 29566
rect 14476 29170 14504 30126
rect 14568 29510 14596 30194
rect 14556 29504 14608 29510
rect 14556 29446 14608 29452
rect 14464 29164 14516 29170
rect 14464 29106 14516 29112
rect 14476 28762 14504 29106
rect 14568 29050 14596 29446
rect 14648 29300 14700 29306
rect 14648 29242 14700 29248
rect 14660 29170 14688 29242
rect 14648 29164 14700 29170
rect 14648 29106 14700 29112
rect 14568 29022 14688 29050
rect 14556 28960 14608 28966
rect 14556 28902 14608 28908
rect 14464 28756 14516 28762
rect 14464 28698 14516 28704
rect 14568 28694 14596 28902
rect 14556 28688 14608 28694
rect 14556 28630 14608 28636
rect 14660 28626 14688 29022
rect 14648 28620 14700 28626
rect 14648 28562 14700 28568
rect 14280 28552 14332 28558
rect 14280 28494 14332 28500
rect 14372 28552 14424 28558
rect 14752 28506 14780 30790
rect 14936 30734 14964 31758
rect 14924 30728 14976 30734
rect 14924 30670 14976 30676
rect 14832 30660 14884 30666
rect 14832 30602 14884 30608
rect 14844 29850 14872 30602
rect 14936 30258 14964 30670
rect 15028 30258 15056 32370
rect 15108 32292 15160 32298
rect 15108 32234 15160 32240
rect 15120 31822 15148 32234
rect 15108 31816 15160 31822
rect 15108 31758 15160 31764
rect 15200 31816 15252 31822
rect 15200 31758 15252 31764
rect 14924 30252 14976 30258
rect 14924 30194 14976 30200
rect 15016 30252 15068 30258
rect 15016 30194 15068 30200
rect 14832 29844 14884 29850
rect 14832 29786 14884 29792
rect 14832 29640 14884 29646
rect 14832 29582 14884 29588
rect 14844 29034 14872 29582
rect 14832 29028 14884 29034
rect 14832 28970 14884 28976
rect 14936 28626 14964 30194
rect 15016 29164 15068 29170
rect 15016 29106 15068 29112
rect 15028 29073 15056 29106
rect 15014 29064 15070 29073
rect 15014 28999 15070 29008
rect 14832 28620 14884 28626
rect 14832 28562 14884 28568
rect 14924 28620 14976 28626
rect 14924 28562 14976 28568
rect 14372 28494 14424 28500
rect 14280 27668 14332 27674
rect 14280 27610 14332 27616
rect 14188 25696 14240 25702
rect 14188 25638 14240 25644
rect 14096 25288 14148 25294
rect 13910 25256 13966 25265
rect 14096 25230 14148 25236
rect 13910 25191 13966 25200
rect 14004 25220 14056 25226
rect 13924 24682 13952 25191
rect 14004 25162 14056 25168
rect 13912 24676 13964 24682
rect 13912 24618 13964 24624
rect 14016 24426 14044 25162
rect 14108 24682 14136 25230
rect 14292 24818 14320 27610
rect 14384 26500 14412 28494
rect 14660 28478 14780 28506
rect 14556 27872 14608 27878
rect 14556 27814 14608 27820
rect 14568 27130 14596 27814
rect 14556 27124 14608 27130
rect 14556 27066 14608 27072
rect 14556 26512 14608 26518
rect 14384 26472 14556 26500
rect 14556 26454 14608 26460
rect 14464 25832 14516 25838
rect 14464 25774 14516 25780
rect 14372 25764 14424 25770
rect 14372 25706 14424 25712
rect 14384 24818 14412 25706
rect 14476 25362 14504 25774
rect 14464 25356 14516 25362
rect 14464 25298 14516 25304
rect 14568 25242 14596 26454
rect 14476 25214 14596 25242
rect 14280 24812 14332 24818
rect 14280 24754 14332 24760
rect 14372 24812 14424 24818
rect 14372 24754 14424 24760
rect 14096 24676 14148 24682
rect 14096 24618 14148 24624
rect 14016 24398 14228 24426
rect 14292 24410 14320 24754
rect 14372 24676 14424 24682
rect 14372 24618 14424 24624
rect 14004 24336 14056 24342
rect 14004 24278 14056 24284
rect 13820 24268 13872 24274
rect 13820 24210 13872 24216
rect 13912 24268 13964 24274
rect 13912 24210 13964 24216
rect 13832 23866 13860 24210
rect 13820 23860 13872 23866
rect 13820 23802 13872 23808
rect 13818 23352 13874 23361
rect 13818 23287 13874 23296
rect 13832 22506 13860 23287
rect 13924 23254 13952 24210
rect 13912 23248 13964 23254
rect 13912 23190 13964 23196
rect 13912 23044 13964 23050
rect 13912 22986 13964 22992
rect 13924 22574 13952 22986
rect 13912 22568 13964 22574
rect 13912 22510 13964 22516
rect 13820 22500 13872 22506
rect 13820 22442 13872 22448
rect 13820 21344 13872 21350
rect 13820 21286 13872 21292
rect 13728 21140 13780 21146
rect 13728 21082 13780 21088
rect 13832 20942 13860 21286
rect 13820 20936 13872 20942
rect 13820 20878 13872 20884
rect 14016 20874 14044 24278
rect 14200 24070 14228 24398
rect 14280 24404 14332 24410
rect 14280 24346 14332 24352
rect 14096 24064 14148 24070
rect 14096 24006 14148 24012
rect 14188 24064 14240 24070
rect 14188 24006 14240 24012
rect 14108 23798 14136 24006
rect 14200 23798 14228 24006
rect 14096 23792 14148 23798
rect 14096 23734 14148 23740
rect 14188 23792 14240 23798
rect 14188 23734 14240 23740
rect 14280 23588 14332 23594
rect 14280 23530 14332 23536
rect 14292 23118 14320 23530
rect 14096 23112 14148 23118
rect 14096 23054 14148 23060
rect 14280 23112 14332 23118
rect 14280 23054 14332 23060
rect 14108 22982 14136 23054
rect 14096 22976 14148 22982
rect 14096 22918 14148 22924
rect 14096 22432 14148 22438
rect 14096 22374 14148 22380
rect 14108 21690 14136 22374
rect 14384 22234 14412 24618
rect 14476 24206 14504 25214
rect 14556 24812 14608 24818
rect 14660 24800 14688 28478
rect 14740 28416 14792 28422
rect 14740 28358 14792 28364
rect 14752 27402 14780 28358
rect 14844 27674 14872 28562
rect 14832 27668 14884 27674
rect 14832 27610 14884 27616
rect 14936 27470 14964 28562
rect 15120 28150 15148 31758
rect 15212 31346 15240 31758
rect 15200 31340 15252 31346
rect 15200 31282 15252 31288
rect 15212 29458 15240 31282
rect 15304 29646 15332 32710
rect 15396 32026 15424 32846
rect 15660 32836 15712 32842
rect 15660 32778 15712 32784
rect 15752 32836 15804 32842
rect 15752 32778 15804 32784
rect 15844 32836 15896 32842
rect 15844 32778 15896 32784
rect 15476 32768 15528 32774
rect 15476 32710 15528 32716
rect 15384 32020 15436 32026
rect 15384 31962 15436 31968
rect 15384 31272 15436 31278
rect 15384 31214 15436 31220
rect 15396 30569 15424 31214
rect 15382 30560 15438 30569
rect 15382 30495 15438 30504
rect 15382 30016 15438 30025
rect 15382 29951 15438 29960
rect 15292 29640 15344 29646
rect 15292 29582 15344 29588
rect 15212 29430 15332 29458
rect 15304 29170 15332 29430
rect 15292 29164 15344 29170
rect 15292 29106 15344 29112
rect 15200 29028 15252 29034
rect 15200 28970 15252 28976
rect 15108 28144 15160 28150
rect 15028 28104 15108 28132
rect 14924 27464 14976 27470
rect 14924 27406 14976 27412
rect 14740 27396 14792 27402
rect 14740 27338 14792 27344
rect 14936 26994 14964 27406
rect 14740 26988 14792 26994
rect 14740 26930 14792 26936
rect 14924 26988 14976 26994
rect 14924 26930 14976 26936
rect 14752 26586 14780 26930
rect 14740 26580 14792 26586
rect 14740 26522 14792 26528
rect 14832 26240 14884 26246
rect 14832 26182 14884 26188
rect 14844 26042 14872 26182
rect 14832 26036 14884 26042
rect 14832 25978 14884 25984
rect 14936 25974 14964 26930
rect 14924 25968 14976 25974
rect 14924 25910 14976 25916
rect 14832 25832 14884 25838
rect 14832 25774 14884 25780
rect 14844 25498 14872 25774
rect 14832 25492 14884 25498
rect 14832 25434 14884 25440
rect 14936 25362 14964 25910
rect 14924 25356 14976 25362
rect 14924 25298 14976 25304
rect 14936 24818 14964 25298
rect 15028 24886 15056 28104
rect 15108 28086 15160 28092
rect 15108 27328 15160 27334
rect 15108 27270 15160 27276
rect 15120 26042 15148 27270
rect 15108 26036 15160 26042
rect 15108 25978 15160 25984
rect 15212 25906 15240 28970
rect 15304 28762 15332 29106
rect 15396 29034 15424 29951
rect 15488 29238 15516 32710
rect 15672 32502 15700 32778
rect 15660 32496 15712 32502
rect 15660 32438 15712 32444
rect 15764 32450 15792 32778
rect 15856 32745 15884 32778
rect 15842 32736 15898 32745
rect 15842 32671 15898 32680
rect 15764 32434 15976 32450
rect 15764 32428 15988 32434
rect 15764 32422 15936 32428
rect 15936 32370 15988 32376
rect 15660 32360 15712 32366
rect 15660 32302 15712 32308
rect 15844 32360 15896 32366
rect 15844 32302 15896 32308
rect 15568 32224 15620 32230
rect 15672 32201 15700 32302
rect 15568 32166 15620 32172
rect 15658 32192 15714 32201
rect 15580 32065 15608 32166
rect 15658 32127 15714 32136
rect 15566 32056 15622 32065
rect 15566 31991 15622 32000
rect 15856 31210 15884 32302
rect 15948 31890 15976 32370
rect 16132 32201 16160 32846
rect 16212 32836 16264 32842
rect 16212 32778 16264 32784
rect 16118 32192 16174 32201
rect 16118 32127 16174 32136
rect 16028 31952 16080 31958
rect 16028 31894 16080 31900
rect 15936 31884 15988 31890
rect 15936 31826 15988 31832
rect 15844 31204 15896 31210
rect 15844 31146 15896 31152
rect 15752 31136 15804 31142
rect 15752 31078 15804 31084
rect 15568 30252 15620 30258
rect 15568 30194 15620 30200
rect 15580 29850 15608 30194
rect 15568 29844 15620 29850
rect 15568 29786 15620 29792
rect 15660 29708 15712 29714
rect 15660 29650 15712 29656
rect 15476 29232 15528 29238
rect 15476 29174 15528 29180
rect 15476 29096 15528 29102
rect 15476 29038 15528 29044
rect 15384 29028 15436 29034
rect 15384 28970 15436 28976
rect 15292 28756 15344 28762
rect 15292 28698 15344 28704
rect 15292 28484 15344 28490
rect 15292 28426 15344 28432
rect 15304 28218 15332 28426
rect 15384 28416 15436 28422
rect 15384 28358 15436 28364
rect 15292 28212 15344 28218
rect 15292 28154 15344 28160
rect 15396 27985 15424 28358
rect 15382 27976 15438 27985
rect 15382 27911 15438 27920
rect 15384 27396 15436 27402
rect 15384 27338 15436 27344
rect 15292 27328 15344 27334
rect 15292 27270 15344 27276
rect 15304 26790 15332 27270
rect 15292 26784 15344 26790
rect 15292 26726 15344 26732
rect 15200 25900 15252 25906
rect 15200 25842 15252 25848
rect 15200 25220 15252 25226
rect 15200 25162 15252 25168
rect 15016 24880 15068 24886
rect 15016 24822 15068 24828
rect 14924 24812 14976 24818
rect 14660 24772 14872 24800
rect 14556 24754 14608 24760
rect 14568 24342 14596 24754
rect 14740 24676 14792 24682
rect 14740 24618 14792 24624
rect 14648 24608 14700 24614
rect 14648 24550 14700 24556
rect 14660 24449 14688 24550
rect 14646 24440 14702 24449
rect 14646 24375 14702 24384
rect 14556 24336 14608 24342
rect 14556 24278 14608 24284
rect 14464 24200 14516 24206
rect 14464 24142 14516 24148
rect 14476 23882 14504 24142
rect 14476 23854 14688 23882
rect 14462 23216 14518 23225
rect 14462 23151 14518 23160
rect 14476 23118 14504 23151
rect 14464 23112 14516 23118
rect 14464 23054 14516 23060
rect 14372 22228 14424 22234
rect 14372 22170 14424 22176
rect 14188 22092 14240 22098
rect 14188 22034 14240 22040
rect 14280 22092 14332 22098
rect 14476 22094 14504 23054
rect 14556 22636 14608 22642
rect 14556 22578 14608 22584
rect 14280 22034 14332 22040
rect 14384 22066 14504 22094
rect 14096 21684 14148 21690
rect 14096 21626 14148 21632
rect 14200 21026 14228 22034
rect 14292 21350 14320 22034
rect 14384 21622 14412 22066
rect 14464 21956 14516 21962
rect 14464 21898 14516 21904
rect 14476 21690 14504 21898
rect 14568 21690 14596 22578
rect 14464 21684 14516 21690
rect 14464 21626 14516 21632
rect 14556 21684 14608 21690
rect 14556 21626 14608 21632
rect 14372 21616 14424 21622
rect 14372 21558 14424 21564
rect 14280 21344 14332 21350
rect 14280 21286 14332 21292
rect 14384 21078 14412 21558
rect 14108 20998 14228 21026
rect 14372 21072 14424 21078
rect 14372 21014 14424 21020
rect 14004 20868 14056 20874
rect 14004 20810 14056 20816
rect 13728 19440 13780 19446
rect 13728 19382 13780 19388
rect 13636 17672 13688 17678
rect 13636 17614 13688 17620
rect 13648 12782 13676 17614
rect 13740 16522 13768 19382
rect 13912 19304 13964 19310
rect 13912 19246 13964 19252
rect 13924 18902 13952 19246
rect 13912 18896 13964 18902
rect 13912 18838 13964 18844
rect 13924 18766 13952 18838
rect 13912 18760 13964 18766
rect 13912 18702 13964 18708
rect 13912 18420 13964 18426
rect 13912 18362 13964 18368
rect 13924 17678 13952 18362
rect 13912 17672 13964 17678
rect 13818 17640 13874 17649
rect 13912 17614 13964 17620
rect 13818 17575 13874 17584
rect 13832 17338 13860 17575
rect 13820 17332 13872 17338
rect 13820 17274 13872 17280
rect 14016 17218 14044 20810
rect 14108 18970 14136 20998
rect 14476 20942 14504 21626
rect 14660 21570 14688 23854
rect 14752 22098 14780 24618
rect 14844 22982 14872 24772
rect 14924 24754 14976 24760
rect 15028 24698 15056 24822
rect 14936 24682 15056 24698
rect 14924 24676 15056 24682
rect 14976 24670 15056 24676
rect 14924 24618 14976 24624
rect 15212 24614 15240 25162
rect 15200 24608 15252 24614
rect 15200 24550 15252 24556
rect 15292 24608 15344 24614
rect 15292 24550 15344 24556
rect 15106 24440 15162 24449
rect 14924 24404 14976 24410
rect 15106 24375 15162 24384
rect 14924 24346 14976 24352
rect 14936 24206 14964 24346
rect 15120 24342 15148 24375
rect 15108 24336 15160 24342
rect 15108 24278 15160 24284
rect 14924 24200 14976 24206
rect 14924 24142 14976 24148
rect 15016 24200 15068 24206
rect 15016 24142 15068 24148
rect 15028 23866 15056 24142
rect 15198 23896 15254 23905
rect 15016 23860 15068 23866
rect 15198 23831 15254 23840
rect 15016 23802 15068 23808
rect 15108 23724 15160 23730
rect 15108 23666 15160 23672
rect 14832 22976 14884 22982
rect 14832 22918 14884 22924
rect 14740 22092 14792 22098
rect 14740 22034 14792 22040
rect 14844 21842 14872 22918
rect 15120 22778 15148 23666
rect 15212 23662 15240 23831
rect 15200 23656 15252 23662
rect 15200 23598 15252 23604
rect 15304 23526 15332 24550
rect 15396 24138 15424 27338
rect 15488 27334 15516 29038
rect 15568 28552 15620 28558
rect 15568 28494 15620 28500
rect 15580 28082 15608 28494
rect 15568 28076 15620 28082
rect 15568 28018 15620 28024
rect 15672 27402 15700 29650
rect 15764 28082 15792 31078
rect 15934 30288 15990 30297
rect 15934 30223 15990 30232
rect 15844 30048 15896 30054
rect 15844 29990 15896 29996
rect 15856 29646 15884 29990
rect 15844 29640 15896 29646
rect 15844 29582 15896 29588
rect 15948 29322 15976 30223
rect 15856 29306 15976 29322
rect 15856 29300 15988 29306
rect 15856 29294 15936 29300
rect 15856 28082 15884 29294
rect 15936 29242 15988 29248
rect 15934 29200 15990 29209
rect 16040 29170 16068 31894
rect 16132 31822 16160 32127
rect 16120 31816 16172 31822
rect 16120 31758 16172 31764
rect 16120 31680 16172 31686
rect 16120 31622 16172 31628
rect 15934 29135 15936 29144
rect 15988 29135 15990 29144
rect 16028 29164 16080 29170
rect 15936 29106 15988 29112
rect 16028 29106 16080 29112
rect 16132 28082 16160 31622
rect 16224 30394 16252 32778
rect 16396 31884 16448 31890
rect 16396 31826 16448 31832
rect 16302 31376 16358 31385
rect 16302 31311 16304 31320
rect 16356 31311 16358 31320
rect 16304 31282 16356 31288
rect 16304 31204 16356 31210
rect 16304 31146 16356 31152
rect 16316 30938 16344 31146
rect 16304 30932 16356 30938
rect 16304 30874 16356 30880
rect 16212 30388 16264 30394
rect 16212 30330 16264 30336
rect 16302 29336 16358 29345
rect 16302 29271 16358 29280
rect 16316 29170 16344 29271
rect 16304 29164 16356 29170
rect 16304 29106 16356 29112
rect 15752 28076 15804 28082
rect 15752 28018 15804 28024
rect 15844 28076 15896 28082
rect 15844 28018 15896 28024
rect 16120 28076 16172 28082
rect 16120 28018 16172 28024
rect 16304 28076 16356 28082
rect 16304 28018 16356 28024
rect 15752 27940 15804 27946
rect 15752 27882 15804 27888
rect 15764 27470 15792 27882
rect 16212 27872 16264 27878
rect 16212 27814 16264 27820
rect 15752 27464 15804 27470
rect 15752 27406 15804 27412
rect 16028 27464 16080 27470
rect 16028 27406 16080 27412
rect 16120 27464 16172 27470
rect 16120 27406 16172 27412
rect 15660 27396 15712 27402
rect 15660 27338 15712 27344
rect 15476 27328 15528 27334
rect 15476 27270 15528 27276
rect 15568 27328 15620 27334
rect 15568 27270 15620 27276
rect 15580 27062 15608 27270
rect 15568 27056 15620 27062
rect 15568 26998 15620 27004
rect 15568 25900 15620 25906
rect 15568 25842 15620 25848
rect 15660 25900 15712 25906
rect 15660 25842 15712 25848
rect 15580 25401 15608 25842
rect 15566 25392 15622 25401
rect 15566 25327 15622 25336
rect 15568 25152 15620 25158
rect 15568 25094 15620 25100
rect 15476 24812 15528 24818
rect 15476 24754 15528 24760
rect 15488 24410 15516 24754
rect 15580 24410 15608 25094
rect 15672 24614 15700 25842
rect 15764 24954 15792 27406
rect 15844 26376 15896 26382
rect 15842 26344 15844 26353
rect 15896 26344 15898 26353
rect 15842 26279 15898 26288
rect 15844 25696 15896 25702
rect 15844 25638 15896 25644
rect 15752 24948 15804 24954
rect 15752 24890 15804 24896
rect 15856 24834 15884 25638
rect 15764 24806 15884 24834
rect 15660 24608 15712 24614
rect 15660 24550 15712 24556
rect 15476 24404 15528 24410
rect 15476 24346 15528 24352
rect 15568 24404 15620 24410
rect 15568 24346 15620 24352
rect 15568 24200 15620 24206
rect 15568 24142 15620 24148
rect 15384 24132 15436 24138
rect 15436 24092 15516 24120
rect 15384 24074 15436 24080
rect 15384 23724 15436 23730
rect 15384 23666 15436 23672
rect 15292 23520 15344 23526
rect 15292 23462 15344 23468
rect 15198 23216 15254 23225
rect 15198 23151 15254 23160
rect 15108 22772 15160 22778
rect 15108 22714 15160 22720
rect 15016 22500 15068 22506
rect 15016 22442 15068 22448
rect 14924 22228 14976 22234
rect 14924 22170 14976 22176
rect 14752 21814 14872 21842
rect 14752 21622 14780 21814
rect 14936 21672 14964 22170
rect 14844 21644 14964 21672
rect 14568 21542 14688 21570
rect 14740 21616 14792 21622
rect 14740 21558 14792 21564
rect 14188 20936 14240 20942
rect 14188 20878 14240 20884
rect 14464 20936 14516 20942
rect 14464 20878 14516 20884
rect 14200 20262 14228 20878
rect 14372 20868 14424 20874
rect 14372 20810 14424 20816
rect 14384 20602 14412 20810
rect 14372 20596 14424 20602
rect 14372 20538 14424 20544
rect 14188 20256 14240 20262
rect 14188 20198 14240 20204
rect 14200 19854 14228 20198
rect 14188 19848 14240 19854
rect 14240 19808 14320 19836
rect 14188 19790 14240 19796
rect 14292 19310 14320 19808
rect 14372 19780 14424 19786
rect 14372 19722 14424 19728
rect 14384 19514 14412 19722
rect 14568 19514 14596 21542
rect 14752 20856 14780 21558
rect 14660 20828 14780 20856
rect 14660 20534 14688 20828
rect 14844 20754 14872 21644
rect 15028 21554 15056 22442
rect 15120 22030 15148 22714
rect 15108 22024 15160 22030
rect 15108 21966 15160 21972
rect 15212 21894 15240 23151
rect 15396 22982 15424 23666
rect 15488 23322 15516 24092
rect 15580 23730 15608 24142
rect 15568 23724 15620 23730
rect 15568 23666 15620 23672
rect 15660 23656 15712 23662
rect 15660 23598 15712 23604
rect 15476 23316 15528 23322
rect 15476 23258 15528 23264
rect 15384 22976 15436 22982
rect 15384 22918 15436 22924
rect 15290 22536 15346 22545
rect 15290 22471 15346 22480
rect 15304 21962 15332 22471
rect 15396 22030 15424 22918
rect 15384 22024 15436 22030
rect 15384 21966 15436 21972
rect 15292 21956 15344 21962
rect 15292 21898 15344 21904
rect 15200 21888 15252 21894
rect 15200 21830 15252 21836
rect 14924 21548 14976 21554
rect 14924 21490 14976 21496
rect 15016 21548 15068 21554
rect 15016 21490 15068 21496
rect 14936 21350 14964 21490
rect 15384 21412 15436 21418
rect 15384 21354 15436 21360
rect 14924 21344 14976 21350
rect 14924 21286 14976 21292
rect 14752 20726 14872 20754
rect 14752 20534 14780 20726
rect 14830 20632 14886 20641
rect 14830 20567 14832 20576
rect 14884 20567 14886 20576
rect 14832 20538 14884 20544
rect 14648 20528 14700 20534
rect 14648 20470 14700 20476
rect 14740 20528 14792 20534
rect 14740 20470 14792 20476
rect 14740 20052 14792 20058
rect 14660 20012 14740 20040
rect 14372 19508 14424 19514
rect 14372 19450 14424 19456
rect 14556 19508 14608 19514
rect 14556 19450 14608 19456
rect 14370 19408 14426 19417
rect 14556 19372 14608 19378
rect 14370 19343 14426 19352
rect 14280 19304 14332 19310
rect 14280 19246 14332 19252
rect 14186 19136 14242 19145
rect 14186 19071 14242 19080
rect 14096 18964 14148 18970
rect 14096 18906 14148 18912
rect 14200 18426 14228 19071
rect 14188 18420 14240 18426
rect 14188 18362 14240 18368
rect 14292 18290 14320 19246
rect 14280 18284 14332 18290
rect 14280 18226 14332 18232
rect 14096 18148 14148 18154
rect 14096 18090 14148 18096
rect 14108 17678 14136 18090
rect 14096 17672 14148 17678
rect 14096 17614 14148 17620
rect 14280 17672 14332 17678
rect 14280 17614 14332 17620
rect 14016 17202 14136 17218
rect 13912 17196 13964 17202
rect 14016 17196 14148 17202
rect 14016 17190 14096 17196
rect 13912 17138 13964 17144
rect 14096 17138 14148 17144
rect 13820 16720 13872 16726
rect 13820 16662 13872 16668
rect 13728 16516 13780 16522
rect 13728 16458 13780 16464
rect 13728 15632 13780 15638
rect 13728 15574 13780 15580
rect 13740 14822 13768 15574
rect 13832 15366 13860 16662
rect 13924 16402 13952 17138
rect 14004 16584 14056 16590
rect 14002 16552 14004 16561
rect 14056 16552 14058 16561
rect 14002 16487 14058 16496
rect 14004 16448 14056 16454
rect 13924 16396 14004 16402
rect 13924 16390 14056 16396
rect 13924 16374 14044 16390
rect 13924 16114 13952 16374
rect 14108 16182 14136 17138
rect 14292 16998 14320 17614
rect 14280 16992 14332 16998
rect 14280 16934 14332 16940
rect 14096 16176 14148 16182
rect 14384 16130 14412 19343
rect 14476 19332 14556 19360
rect 14476 17338 14504 19332
rect 14556 19314 14608 19320
rect 14660 18766 14688 20012
rect 14740 19994 14792 20000
rect 14936 19530 14964 21286
rect 15108 21140 15160 21146
rect 15108 21082 15160 21088
rect 15016 20868 15068 20874
rect 15016 20810 15068 20816
rect 15028 20602 15056 20810
rect 15120 20602 15148 21082
rect 15016 20596 15068 20602
rect 15016 20538 15068 20544
rect 15108 20596 15160 20602
rect 15108 20538 15160 20544
rect 15396 20466 15424 21354
rect 15384 20460 15436 20466
rect 15384 20402 15436 20408
rect 15488 20398 15516 23258
rect 15568 21616 15620 21622
rect 15568 21558 15620 21564
rect 15580 20466 15608 21558
rect 15568 20460 15620 20466
rect 15568 20402 15620 20408
rect 15476 20392 15528 20398
rect 15476 20334 15528 20340
rect 15384 20324 15436 20330
rect 15384 20266 15436 20272
rect 15198 19816 15254 19825
rect 15198 19751 15254 19760
rect 15212 19718 15240 19751
rect 15200 19712 15252 19718
rect 15200 19654 15252 19660
rect 14844 19502 14964 19530
rect 14648 18760 14700 18766
rect 14648 18702 14700 18708
rect 14740 18760 14792 18766
rect 14740 18702 14792 18708
rect 14556 18284 14608 18290
rect 14556 18226 14608 18232
rect 14568 17882 14596 18226
rect 14556 17876 14608 17882
rect 14556 17818 14608 17824
rect 14464 17332 14516 17338
rect 14464 17274 14516 17280
rect 14660 17218 14688 18702
rect 14752 17338 14780 18702
rect 14844 17814 14872 19502
rect 14924 19440 14976 19446
rect 14924 19382 14976 19388
rect 14832 17808 14884 17814
rect 14832 17750 14884 17756
rect 14844 17490 14872 17750
rect 14936 17678 14964 19382
rect 15016 19372 15068 19378
rect 15016 19314 15068 19320
rect 15028 18970 15056 19314
rect 15108 19168 15160 19174
rect 15108 19110 15160 19116
rect 15016 18964 15068 18970
rect 15016 18906 15068 18912
rect 15120 18766 15148 19110
rect 15396 18970 15424 20266
rect 15384 18964 15436 18970
rect 15384 18906 15436 18912
rect 15200 18896 15252 18902
rect 15396 18873 15424 18906
rect 15200 18838 15252 18844
rect 15382 18864 15438 18873
rect 15108 18760 15160 18766
rect 15108 18702 15160 18708
rect 15120 17882 15148 18702
rect 15108 17876 15160 17882
rect 15108 17818 15160 17824
rect 14924 17672 14976 17678
rect 14924 17614 14976 17620
rect 15016 17536 15068 17542
rect 14844 17462 14964 17490
rect 15016 17478 15068 17484
rect 14740 17332 14792 17338
rect 14740 17274 14792 17280
rect 14568 17202 14688 17218
rect 14556 17196 14688 17202
rect 14608 17190 14688 17196
rect 14830 17232 14886 17241
rect 14830 17167 14832 17176
rect 14556 17138 14608 17144
rect 14884 17167 14886 17176
rect 14832 17138 14884 17144
rect 14740 17128 14792 17134
rect 14646 17096 14702 17105
rect 14740 17070 14792 17076
rect 14646 17031 14702 17040
rect 14462 16552 14518 16561
rect 14462 16487 14518 16496
rect 14556 16516 14608 16522
rect 14096 16118 14148 16124
rect 13912 16108 13964 16114
rect 13912 16050 13964 16056
rect 14108 15978 14136 16118
rect 14292 16102 14412 16130
rect 14096 15972 14148 15978
rect 14096 15914 14148 15920
rect 14004 15700 14056 15706
rect 14004 15642 14056 15648
rect 13820 15360 13872 15366
rect 13820 15302 13872 15308
rect 13820 14952 13872 14958
rect 13820 14894 13872 14900
rect 13728 14816 13780 14822
rect 13728 14758 13780 14764
rect 13832 14278 13860 14894
rect 14016 14550 14044 15642
rect 14188 15496 14240 15502
rect 14188 15438 14240 15444
rect 14094 15056 14150 15065
rect 14094 14991 14096 15000
rect 14148 14991 14150 15000
rect 14096 14962 14148 14968
rect 14004 14544 14056 14550
rect 14004 14486 14056 14492
rect 13912 14476 13964 14482
rect 13912 14418 13964 14424
rect 13820 14272 13872 14278
rect 13820 14214 13872 14220
rect 13726 13968 13782 13977
rect 13924 13938 13952 14418
rect 13726 13903 13782 13912
rect 13912 13932 13964 13938
rect 13636 12776 13688 12782
rect 13636 12718 13688 12724
rect 13544 12708 13596 12714
rect 13544 12650 13596 12656
rect 13544 12300 13596 12306
rect 13544 12242 13596 12248
rect 13450 12200 13506 12209
rect 13450 12135 13506 12144
rect 13464 11354 13492 12135
rect 13556 11898 13584 12242
rect 13544 11892 13596 11898
rect 13544 11834 13596 11840
rect 13648 11744 13676 12718
rect 13740 11898 13768 13903
rect 13912 13874 13964 13880
rect 13820 13864 13872 13870
rect 13820 13806 13872 13812
rect 13832 13462 13860 13806
rect 14016 13802 14044 14486
rect 14200 14074 14228 15438
rect 14188 14068 14240 14074
rect 14188 14010 14240 14016
rect 14004 13796 14056 13802
rect 14004 13738 14056 13744
rect 13912 13524 13964 13530
rect 13912 13466 13964 13472
rect 13820 13456 13872 13462
rect 13820 13398 13872 13404
rect 13924 13308 13952 13466
rect 13832 13280 13952 13308
rect 13728 11892 13780 11898
rect 13728 11834 13780 11840
rect 13648 11716 13768 11744
rect 13634 11656 13690 11665
rect 13634 11591 13690 11600
rect 13320 11308 13400 11336
rect 13452 11348 13504 11354
rect 13268 11290 13320 11296
rect 13452 11290 13504 11296
rect 13174 10160 13230 10169
rect 12900 10124 12952 10130
rect 13174 10095 13230 10104
rect 12900 10066 12952 10072
rect 12912 9761 12940 10066
rect 13188 10062 13216 10095
rect 13176 10056 13228 10062
rect 13176 9998 13228 10004
rect 13084 9988 13136 9994
rect 13084 9930 13136 9936
rect 12898 9752 12954 9761
rect 12898 9687 12900 9696
rect 12952 9687 12954 9696
rect 12900 9658 12952 9664
rect 12912 8634 12940 9658
rect 13096 9586 13124 9930
rect 13464 9674 13492 11290
rect 13648 10810 13676 11591
rect 13636 10804 13688 10810
rect 13636 10746 13688 10752
rect 13464 9646 13676 9674
rect 13084 9580 13136 9586
rect 13084 9522 13136 9528
rect 13360 9580 13412 9586
rect 13360 9522 13412 9528
rect 13268 9376 13320 9382
rect 13268 9318 13320 9324
rect 12900 8628 12952 8634
rect 12900 8570 12952 8576
rect 12636 8486 12756 8514
rect 12808 8560 12860 8566
rect 12808 8502 12860 8508
rect 12532 7948 12584 7954
rect 12532 7890 12584 7896
rect 12544 7478 12572 7890
rect 12532 7472 12584 7478
rect 12532 7414 12584 7420
rect 12636 6798 12664 8486
rect 12716 8084 12768 8090
rect 12716 8026 12768 8032
rect 12624 6792 12676 6798
rect 12624 6734 12676 6740
rect 12728 6118 12756 8026
rect 12820 8022 12848 8502
rect 13084 8424 13136 8430
rect 13084 8366 13136 8372
rect 12992 8288 13044 8294
rect 12992 8230 13044 8236
rect 12808 8016 12860 8022
rect 12808 7958 12860 7964
rect 12900 7880 12952 7886
rect 12900 7822 12952 7828
rect 12806 7576 12862 7585
rect 12806 7511 12862 7520
rect 12820 6118 12848 7511
rect 12912 6390 12940 7822
rect 13004 7274 13032 8230
rect 12992 7268 13044 7274
rect 12992 7210 13044 7216
rect 13004 6730 13032 7210
rect 12992 6724 13044 6730
rect 12992 6666 13044 6672
rect 13096 6458 13124 8366
rect 13280 7857 13308 9318
rect 13372 8634 13400 9522
rect 13452 9172 13504 9178
rect 13452 9114 13504 9120
rect 13360 8628 13412 8634
rect 13360 8570 13412 8576
rect 13360 8424 13412 8430
rect 13360 8366 13412 8372
rect 13266 7848 13322 7857
rect 13266 7783 13322 7792
rect 13176 7404 13228 7410
rect 13176 7346 13228 7352
rect 13188 7002 13216 7346
rect 13176 6996 13228 7002
rect 13176 6938 13228 6944
rect 13280 6798 13308 7783
rect 13372 6798 13400 8366
rect 13464 8090 13492 9114
rect 13544 8968 13596 8974
rect 13544 8910 13596 8916
rect 13452 8084 13504 8090
rect 13452 8026 13504 8032
rect 13556 7886 13584 8910
rect 13648 8480 13676 9646
rect 13740 8634 13768 11716
rect 13832 11150 13860 13280
rect 14016 12374 14044 13738
rect 14200 13546 14228 14010
rect 14108 13518 14228 13546
rect 14108 13326 14136 13518
rect 14188 13456 14240 13462
rect 14188 13398 14240 13404
rect 14096 13320 14148 13326
rect 14096 13262 14148 13268
rect 14096 13184 14148 13190
rect 14096 13126 14148 13132
rect 14108 12986 14136 13126
rect 14096 12980 14148 12986
rect 14096 12922 14148 12928
rect 14200 12918 14228 13398
rect 14188 12912 14240 12918
rect 14188 12854 14240 12860
rect 14188 12640 14240 12646
rect 14188 12582 14240 12588
rect 14004 12368 14056 12374
rect 14004 12310 14056 12316
rect 14200 12238 14228 12582
rect 13912 12232 13964 12238
rect 13912 12174 13964 12180
rect 14188 12232 14240 12238
rect 14188 12174 14240 12180
rect 13924 12102 13952 12174
rect 13912 12096 13964 12102
rect 14096 12096 14148 12102
rect 13912 12038 13964 12044
rect 14002 12064 14058 12073
rect 14096 12038 14148 12044
rect 14002 11999 14058 12008
rect 13912 11756 13964 11762
rect 13912 11698 13964 11704
rect 13924 11218 13952 11698
rect 14016 11626 14044 11999
rect 14108 11762 14136 12038
rect 14096 11756 14148 11762
rect 14096 11698 14148 11704
rect 14004 11620 14056 11626
rect 14004 11562 14056 11568
rect 14200 11354 14228 12174
rect 14292 11694 14320 16102
rect 14372 15360 14424 15366
rect 14372 15302 14424 15308
rect 14384 13870 14412 15302
rect 14476 15026 14504 16487
rect 14556 16458 14608 16464
rect 14568 15978 14596 16458
rect 14660 16114 14688 17031
rect 14752 16674 14780 17070
rect 14936 16810 14964 17462
rect 15028 17202 15056 17478
rect 15106 17232 15162 17241
rect 15016 17196 15068 17202
rect 15212 17218 15240 18838
rect 15488 18834 15516 20334
rect 15580 19446 15608 20402
rect 15672 19961 15700 23598
rect 15764 22710 15792 24806
rect 15844 24608 15896 24614
rect 15844 24550 15896 24556
rect 15856 24138 15884 24550
rect 15844 24132 15896 24138
rect 15844 24074 15896 24080
rect 15936 24132 15988 24138
rect 15936 24074 15988 24080
rect 15948 23662 15976 24074
rect 15936 23656 15988 23662
rect 15936 23598 15988 23604
rect 16040 22778 16068 27406
rect 16132 26382 16160 27406
rect 16120 26376 16172 26382
rect 16120 26318 16172 26324
rect 16224 25945 16252 27814
rect 16316 26790 16344 28018
rect 16304 26784 16356 26790
rect 16304 26726 16356 26732
rect 16210 25936 16266 25945
rect 16210 25871 16266 25880
rect 16212 25832 16264 25838
rect 16212 25774 16264 25780
rect 16224 25158 16252 25774
rect 16212 25152 16264 25158
rect 16212 25094 16264 25100
rect 16224 24886 16252 25094
rect 16212 24880 16264 24886
rect 16212 24822 16264 24828
rect 16224 24206 16252 24822
rect 16212 24200 16264 24206
rect 16212 24142 16264 24148
rect 16120 23656 16172 23662
rect 16120 23598 16172 23604
rect 16028 22772 16080 22778
rect 16028 22714 16080 22720
rect 15752 22704 15804 22710
rect 15752 22646 15804 22652
rect 15658 19952 15714 19961
rect 15658 19887 15714 19896
rect 15660 19848 15712 19854
rect 15660 19790 15712 19796
rect 15568 19440 15620 19446
rect 15672 19417 15700 19790
rect 15568 19382 15620 19388
rect 15658 19408 15714 19417
rect 15382 18799 15438 18808
rect 15476 18828 15528 18834
rect 15476 18770 15528 18776
rect 15384 18760 15436 18766
rect 15384 18702 15436 18708
rect 15396 18426 15424 18702
rect 15384 18420 15436 18426
rect 15384 18362 15436 18368
rect 15384 18080 15436 18086
rect 15304 18028 15384 18034
rect 15304 18022 15436 18028
rect 15304 18006 15424 18022
rect 15304 17610 15332 18006
rect 15292 17604 15344 17610
rect 15292 17546 15344 17552
rect 15304 17270 15332 17546
rect 15162 17190 15240 17218
rect 15292 17264 15344 17270
rect 15292 17206 15344 17212
rect 15384 17196 15436 17202
rect 15106 17167 15162 17176
rect 15016 17138 15068 17144
rect 15384 17138 15436 17144
rect 15198 17096 15254 17105
rect 15016 17060 15068 17066
rect 15198 17031 15200 17040
rect 15016 17002 15068 17008
rect 15252 17031 15254 17040
rect 15200 17002 15252 17008
rect 15028 16946 15056 17002
rect 15028 16918 15240 16946
rect 14936 16782 15148 16810
rect 14752 16646 14964 16674
rect 14740 16584 14792 16590
rect 14738 16552 14740 16561
rect 14792 16552 14794 16561
rect 14738 16487 14794 16496
rect 14832 16516 14884 16522
rect 14832 16458 14884 16464
rect 14648 16108 14700 16114
rect 14648 16050 14700 16056
rect 14556 15972 14608 15978
rect 14556 15914 14608 15920
rect 14464 15020 14516 15026
rect 14464 14962 14516 14968
rect 14568 14414 14596 15914
rect 14660 15706 14688 16050
rect 14844 15706 14872 16458
rect 14936 16182 14964 16646
rect 15120 16522 15148 16782
rect 15108 16516 15160 16522
rect 15108 16458 15160 16464
rect 15016 16448 15068 16454
rect 15212 16425 15240 16918
rect 15396 16794 15424 17138
rect 15488 16998 15516 18770
rect 15580 18766 15608 19382
rect 15658 19343 15714 19352
rect 15764 18850 15792 22646
rect 15936 22024 15988 22030
rect 15936 21966 15988 21972
rect 16028 22024 16080 22030
rect 16028 21966 16080 21972
rect 15844 21888 15896 21894
rect 15842 21856 15844 21865
rect 15896 21856 15898 21865
rect 15842 21791 15898 21800
rect 15844 21548 15896 21554
rect 15948 21536 15976 21966
rect 16040 21690 16068 21966
rect 16028 21684 16080 21690
rect 16028 21626 16080 21632
rect 15896 21508 15976 21536
rect 15844 21490 15896 21496
rect 15844 21412 15896 21418
rect 15844 21354 15896 21360
rect 15672 18822 15792 18850
rect 15568 18760 15620 18766
rect 15568 18702 15620 18708
rect 15672 18442 15700 18822
rect 15752 18692 15804 18698
rect 15752 18634 15804 18640
rect 15580 18414 15700 18442
rect 15580 17746 15608 18414
rect 15764 18358 15792 18634
rect 15752 18352 15804 18358
rect 15752 18294 15804 18300
rect 15856 18290 15884 21354
rect 15948 20806 15976 21508
rect 16028 21548 16080 21554
rect 16028 21490 16080 21496
rect 15936 20800 15988 20806
rect 15936 20742 15988 20748
rect 15948 19854 15976 20742
rect 16040 20641 16068 21490
rect 16026 20632 16082 20641
rect 16026 20567 16082 20576
rect 16132 20584 16160 23598
rect 16316 22642 16344 26726
rect 16408 24138 16436 31826
rect 16396 24132 16448 24138
rect 16396 24074 16448 24080
rect 16500 23798 16528 33050
rect 16488 23792 16540 23798
rect 16488 23734 16540 23740
rect 16500 22710 16528 23734
rect 16488 22704 16540 22710
rect 16488 22646 16540 22652
rect 16304 22636 16356 22642
rect 16304 22578 16356 22584
rect 16212 21888 16264 21894
rect 16212 21830 16264 21836
rect 16224 21185 16252 21830
rect 16500 21486 16528 22646
rect 16488 21480 16540 21486
rect 16488 21422 16540 21428
rect 16304 21344 16356 21350
rect 16304 21286 16356 21292
rect 16210 21176 16266 21185
rect 16210 21111 16266 21120
rect 16040 20466 16068 20567
rect 16132 20556 16252 20584
rect 16028 20460 16080 20466
rect 16028 20402 16080 20408
rect 16120 20460 16172 20466
rect 16120 20402 16172 20408
rect 16132 20058 16160 20402
rect 16120 20052 16172 20058
rect 16120 19994 16172 20000
rect 16224 19854 16252 20556
rect 16316 20505 16344 21286
rect 16302 20496 16358 20505
rect 16302 20431 16358 20440
rect 16304 20392 16356 20398
rect 16304 20334 16356 20340
rect 16316 19922 16344 20334
rect 16394 19952 16450 19961
rect 16304 19916 16356 19922
rect 16394 19887 16450 19896
rect 16304 19858 16356 19864
rect 15936 19848 15988 19854
rect 15936 19790 15988 19796
rect 16212 19848 16264 19854
rect 16212 19790 16264 19796
rect 16028 19712 16080 19718
rect 16028 19654 16080 19660
rect 15936 19168 15988 19174
rect 15936 19110 15988 19116
rect 15948 18698 15976 19110
rect 16040 18698 16068 19654
rect 16120 18760 16172 18766
rect 16224 18748 16252 19790
rect 16172 18720 16252 18748
rect 16304 18760 16356 18766
rect 16302 18728 16304 18737
rect 16356 18728 16358 18737
rect 16120 18702 16172 18708
rect 15936 18692 15988 18698
rect 15936 18634 15988 18640
rect 16028 18692 16080 18698
rect 16302 18663 16358 18672
rect 16028 18634 16080 18640
rect 15660 18284 15712 18290
rect 15660 18226 15712 18232
rect 15844 18284 15896 18290
rect 15844 18226 15896 18232
rect 15568 17740 15620 17746
rect 15568 17682 15620 17688
rect 15672 17610 15700 18226
rect 16040 17626 16068 18634
rect 16302 17776 16358 17785
rect 16212 17740 16264 17746
rect 16302 17711 16358 17720
rect 16212 17682 16264 17688
rect 15660 17604 15712 17610
rect 15660 17546 15712 17552
rect 15844 17604 15896 17610
rect 16040 17598 16160 17626
rect 15844 17546 15896 17552
rect 15568 17128 15620 17134
rect 15568 17070 15620 17076
rect 15476 16992 15528 16998
rect 15476 16934 15528 16940
rect 15384 16788 15436 16794
rect 15384 16730 15436 16736
rect 15488 16658 15516 16934
rect 15580 16833 15608 17070
rect 15566 16824 15622 16833
rect 15566 16759 15622 16768
rect 15476 16652 15528 16658
rect 15476 16594 15528 16600
rect 15568 16448 15620 16454
rect 15016 16390 15068 16396
rect 15198 16416 15254 16425
rect 14924 16176 14976 16182
rect 14924 16118 14976 16124
rect 14648 15700 14700 15706
rect 14832 15700 14884 15706
rect 14648 15642 14700 15648
rect 14752 15660 14832 15688
rect 14660 15366 14688 15642
rect 14648 15360 14700 15366
rect 14648 15302 14700 15308
rect 14646 15056 14702 15065
rect 14752 15026 14780 15660
rect 14832 15642 14884 15648
rect 14936 15502 14964 16118
rect 15028 15570 15056 16390
rect 15568 16390 15620 16396
rect 15198 16351 15254 16360
rect 15106 16280 15162 16289
rect 15106 16215 15162 16224
rect 15292 16244 15344 16250
rect 15016 15564 15068 15570
rect 15016 15506 15068 15512
rect 14924 15496 14976 15502
rect 14924 15438 14976 15444
rect 14646 14991 14702 15000
rect 14740 15020 14792 15026
rect 14556 14408 14608 14414
rect 14556 14350 14608 14356
rect 14568 13870 14596 14350
rect 14372 13864 14424 13870
rect 14372 13806 14424 13812
rect 14556 13864 14608 13870
rect 14556 13806 14608 13812
rect 14384 13410 14412 13806
rect 14384 13394 14504 13410
rect 14372 13388 14504 13394
rect 14424 13382 14504 13388
rect 14372 13330 14424 13336
rect 14372 12844 14424 12850
rect 14372 12786 14424 12792
rect 14384 11914 14412 12786
rect 14476 12073 14504 13382
rect 14568 12170 14596 13806
rect 14660 13190 14688 14991
rect 14740 14962 14792 14968
rect 14832 14884 14884 14890
rect 14832 14826 14884 14832
rect 14740 14816 14792 14822
rect 14740 14758 14792 14764
rect 14752 14414 14780 14758
rect 14740 14408 14792 14414
rect 14740 14350 14792 14356
rect 14740 13252 14792 13258
rect 14740 13194 14792 13200
rect 14648 13184 14700 13190
rect 14648 13126 14700 13132
rect 14752 12782 14780 13194
rect 14648 12776 14700 12782
rect 14648 12718 14700 12724
rect 14740 12776 14792 12782
rect 14740 12718 14792 12724
rect 14660 12374 14688 12718
rect 14648 12368 14700 12374
rect 14648 12310 14700 12316
rect 14556 12164 14608 12170
rect 14556 12106 14608 12112
rect 14752 12102 14780 12718
rect 14844 12646 14872 14826
rect 14936 14278 14964 15438
rect 15016 15020 15068 15026
rect 15120 15008 15148 16215
rect 15292 16186 15344 16192
rect 15304 15745 15332 16186
rect 15580 16182 15608 16390
rect 15568 16176 15620 16182
rect 15568 16118 15620 16124
rect 15672 16114 15700 17546
rect 15752 17196 15804 17202
rect 15752 17138 15804 17144
rect 15764 16697 15792 17138
rect 15750 16688 15806 16697
rect 15750 16623 15806 16632
rect 15752 16516 15804 16522
rect 15752 16458 15804 16464
rect 15764 16289 15792 16458
rect 15750 16280 15806 16289
rect 15750 16215 15806 16224
rect 15660 16108 15712 16114
rect 15660 16050 15712 16056
rect 15856 15910 15884 17546
rect 16028 17536 16080 17542
rect 16028 17478 16080 17484
rect 16040 16590 16068 17478
rect 16028 16584 16080 16590
rect 16028 16526 16080 16532
rect 15844 15904 15896 15910
rect 15844 15846 15896 15852
rect 16028 15904 16080 15910
rect 16028 15846 16080 15852
rect 15290 15736 15346 15745
rect 15290 15671 15346 15680
rect 15290 15600 15346 15609
rect 15290 15535 15346 15544
rect 15304 15502 15332 15535
rect 16040 15502 16068 15846
rect 16132 15502 16160 17598
rect 15292 15496 15344 15502
rect 15292 15438 15344 15444
rect 15568 15496 15620 15502
rect 15568 15438 15620 15444
rect 16028 15496 16080 15502
rect 16028 15438 16080 15444
rect 16120 15496 16172 15502
rect 16120 15438 16172 15444
rect 15068 14980 15148 15008
rect 15016 14962 15068 14968
rect 15028 14890 15056 14962
rect 15016 14884 15068 14890
rect 15016 14826 15068 14832
rect 15108 14816 15160 14822
rect 15108 14758 15160 14764
rect 14924 14272 14976 14278
rect 14924 14214 14976 14220
rect 14936 12850 14964 14214
rect 15120 14006 15148 14758
rect 15200 14612 15252 14618
rect 15200 14554 15252 14560
rect 15212 14226 15240 14554
rect 15304 14346 15332 15438
rect 15382 15192 15438 15201
rect 15382 15127 15438 15136
rect 15396 15026 15424 15127
rect 15384 15020 15436 15026
rect 15384 14962 15436 14968
rect 15292 14340 15344 14346
rect 15292 14282 15344 14288
rect 15212 14198 15332 14226
rect 15200 14068 15252 14074
rect 15200 14010 15252 14016
rect 15108 14000 15160 14006
rect 15108 13942 15160 13948
rect 15108 13524 15160 13530
rect 15108 13466 15160 13472
rect 15120 12986 15148 13466
rect 15212 13326 15240 14010
rect 15304 13394 15332 14198
rect 15396 13818 15424 14962
rect 15396 13790 15516 13818
rect 15382 13696 15438 13705
rect 15382 13631 15438 13640
rect 15396 13530 15424 13631
rect 15384 13524 15436 13530
rect 15384 13466 15436 13472
rect 15292 13388 15344 13394
rect 15292 13330 15344 13336
rect 15200 13320 15252 13326
rect 15200 13262 15252 13268
rect 15292 13252 15344 13258
rect 15292 13194 15344 13200
rect 15108 12980 15160 12986
rect 15108 12922 15160 12928
rect 14924 12844 14976 12850
rect 14924 12786 14976 12792
rect 14832 12640 14884 12646
rect 14832 12582 14884 12588
rect 14936 12322 14964 12786
rect 15200 12776 15252 12782
rect 15200 12718 15252 12724
rect 15016 12436 15068 12442
rect 15212 12434 15240 12718
rect 15016 12378 15068 12384
rect 15120 12406 15240 12434
rect 15028 12345 15056 12378
rect 14844 12294 14964 12322
rect 15014 12336 15070 12345
rect 14740 12096 14792 12102
rect 14462 12064 14518 12073
rect 14740 12038 14792 12044
rect 14462 11999 14518 12008
rect 14384 11886 14596 11914
rect 14370 11792 14426 11801
rect 14370 11727 14372 11736
rect 14424 11727 14426 11736
rect 14372 11698 14424 11704
rect 14280 11688 14332 11694
rect 14280 11630 14332 11636
rect 14188 11348 14240 11354
rect 14188 11290 14240 11296
rect 13912 11212 13964 11218
rect 13912 11154 13964 11160
rect 13820 11144 13872 11150
rect 13820 11086 13872 11092
rect 13832 9654 13860 11086
rect 14292 11082 14320 11630
rect 14372 11552 14424 11558
rect 14568 11506 14596 11886
rect 14372 11494 14424 11500
rect 13912 11076 13964 11082
rect 13912 11018 13964 11024
rect 14280 11076 14332 11082
rect 14280 11018 14332 11024
rect 13820 9648 13872 9654
rect 13820 9590 13872 9596
rect 13820 8968 13872 8974
rect 13924 8956 13952 11018
rect 14096 11008 14148 11014
rect 14096 10950 14148 10956
rect 14108 10674 14136 10950
rect 14384 10674 14412 11494
rect 14476 11478 14596 11506
rect 14476 11150 14504 11478
rect 14556 11348 14608 11354
rect 14556 11290 14608 11296
rect 14568 11150 14596 11290
rect 14464 11144 14516 11150
rect 14464 11086 14516 11092
rect 14556 11144 14608 11150
rect 14556 11086 14608 11092
rect 14476 10674 14504 11086
rect 14096 10668 14148 10674
rect 14096 10610 14148 10616
rect 14372 10668 14424 10674
rect 14372 10610 14424 10616
rect 14464 10668 14516 10674
rect 14464 10610 14516 10616
rect 14004 10464 14056 10470
rect 14004 10406 14056 10412
rect 14016 10062 14044 10406
rect 14096 10192 14148 10198
rect 14476 10146 14504 10610
rect 14148 10140 14504 10146
rect 14096 10134 14504 10140
rect 14108 10118 14504 10134
rect 14004 10056 14056 10062
rect 14004 9998 14056 10004
rect 13872 8928 13952 8956
rect 13820 8910 13872 8916
rect 13728 8628 13780 8634
rect 13728 8570 13780 8576
rect 13728 8492 13780 8498
rect 13648 8452 13728 8480
rect 13728 8434 13780 8440
rect 13544 7880 13596 7886
rect 13544 7822 13596 7828
rect 13636 7880 13688 7886
rect 13636 7822 13688 7828
rect 13728 7880 13780 7886
rect 13728 7822 13780 7828
rect 13648 7546 13676 7822
rect 13636 7540 13688 7546
rect 13636 7482 13688 7488
rect 13740 6798 13768 7822
rect 13268 6792 13320 6798
rect 13268 6734 13320 6740
rect 13360 6792 13412 6798
rect 13360 6734 13412 6740
rect 13544 6792 13596 6798
rect 13544 6734 13596 6740
rect 13728 6792 13780 6798
rect 13728 6734 13780 6740
rect 13176 6656 13228 6662
rect 13372 6633 13400 6734
rect 13176 6598 13228 6604
rect 13358 6624 13414 6633
rect 13084 6452 13136 6458
rect 13084 6394 13136 6400
rect 12900 6384 12952 6390
rect 13188 6361 13216 6598
rect 13358 6559 13414 6568
rect 12900 6326 12952 6332
rect 13174 6352 13230 6361
rect 13174 6287 13230 6296
rect 12716 6112 12768 6118
rect 12716 6054 12768 6060
rect 12808 6112 12860 6118
rect 12808 6054 12860 6060
rect 12806 5944 12862 5953
rect 12806 5879 12862 5888
rect 12820 5710 12848 5879
rect 12256 5704 12308 5710
rect 12256 5646 12308 5652
rect 12808 5704 12860 5710
rect 12808 5646 12860 5652
rect 13084 5636 13136 5642
rect 13084 5578 13136 5584
rect 12348 5568 12400 5574
rect 12346 5536 12348 5545
rect 12400 5536 12402 5545
rect 12346 5471 12402 5480
rect 12990 5400 13046 5409
rect 12716 5364 12768 5370
rect 12990 5335 13046 5344
rect 12716 5306 12768 5312
rect 12072 5160 12124 5166
rect 12072 5102 12124 5108
rect 12164 5160 12216 5166
rect 12164 5102 12216 5108
rect 11704 5024 11756 5030
rect 11704 4966 11756 4972
rect 11716 4622 11744 4966
rect 11704 4616 11756 4622
rect 11704 4558 11756 4564
rect 11612 4548 11664 4554
rect 11612 4490 11664 4496
rect 11624 4321 11652 4490
rect 12084 4486 12112 5102
rect 12072 4480 12124 4486
rect 12072 4422 12124 4428
rect 11610 4312 11666 4321
rect 11610 4247 11612 4256
rect 11664 4247 11666 4256
rect 11612 4218 11664 4224
rect 12176 3738 12204 5102
rect 12440 5024 12492 5030
rect 12440 4966 12492 4972
rect 12164 3732 12216 3738
rect 12164 3674 12216 3680
rect 11980 3596 12032 3602
rect 11980 3538 12032 3544
rect 11520 3460 11572 3466
rect 11520 3402 11572 3408
rect 11244 3188 11296 3194
rect 11244 3130 11296 3136
rect 11992 3126 12020 3538
rect 12452 3466 12480 4966
rect 12728 4826 12756 5306
rect 12898 5264 12954 5273
rect 12898 5199 12900 5208
rect 12952 5199 12954 5208
rect 12900 5170 12952 5176
rect 13004 5166 13032 5335
rect 12992 5160 13044 5166
rect 12992 5102 13044 5108
rect 12900 5092 12952 5098
rect 12900 5034 12952 5040
rect 12716 4820 12768 4826
rect 12716 4762 12768 4768
rect 12912 4690 12940 5034
rect 12900 4684 12952 4690
rect 12900 4626 12952 4632
rect 12900 4480 12952 4486
rect 12900 4422 12952 4428
rect 12912 4214 12940 4422
rect 12900 4208 12952 4214
rect 12900 4150 12952 4156
rect 13096 3534 13124 5578
rect 13372 5302 13400 6559
rect 13556 6458 13584 6734
rect 13636 6656 13688 6662
rect 13636 6598 13688 6604
rect 13544 6452 13596 6458
rect 13544 6394 13596 6400
rect 13648 6338 13676 6598
rect 13556 6322 13676 6338
rect 13544 6316 13676 6322
rect 13596 6310 13676 6316
rect 13832 6304 13860 8910
rect 13912 8832 13964 8838
rect 13912 8774 13964 8780
rect 13924 8498 13952 8774
rect 14016 8498 14044 9998
rect 14188 9648 14240 9654
rect 14188 9590 14240 9596
rect 13912 8492 13964 8498
rect 13912 8434 13964 8440
rect 14004 8492 14056 8498
rect 14004 8434 14056 8440
rect 14016 7886 14044 8434
rect 14004 7880 14056 7886
rect 14004 7822 14056 7828
rect 14004 7200 14056 7206
rect 14004 7142 14056 7148
rect 14016 6798 14044 7142
rect 14200 6798 14228 9590
rect 14476 9466 14504 10118
rect 14568 9722 14596 11086
rect 14556 9716 14608 9722
rect 14556 9658 14608 9664
rect 14752 9586 14780 12038
rect 14844 11830 14872 12294
rect 15014 12271 15070 12280
rect 14924 12164 14976 12170
rect 14924 12106 14976 12112
rect 14832 11824 14884 11830
rect 14832 11766 14884 11772
rect 14936 11762 14964 12106
rect 15120 11898 15148 12406
rect 15304 12306 15332 13194
rect 15488 12434 15516 13790
rect 15580 13530 15608 15438
rect 15660 15020 15712 15026
rect 15660 14962 15712 14968
rect 15936 15020 15988 15026
rect 15936 14962 15988 14968
rect 16028 15020 16080 15026
rect 16028 14962 16080 14968
rect 15672 14618 15700 14962
rect 15948 14890 15976 14962
rect 15936 14884 15988 14890
rect 15936 14826 15988 14832
rect 15660 14612 15712 14618
rect 15660 14554 15712 14560
rect 15660 14408 15712 14414
rect 15660 14350 15712 14356
rect 15672 13734 15700 14350
rect 15660 13728 15712 13734
rect 15660 13670 15712 13676
rect 15568 13524 15620 13530
rect 15568 13466 15620 13472
rect 15672 12850 15700 13670
rect 15752 13184 15804 13190
rect 15752 13126 15804 13132
rect 15764 12850 15792 13126
rect 15660 12844 15712 12850
rect 15660 12786 15712 12792
rect 15752 12844 15804 12850
rect 15752 12786 15804 12792
rect 15844 12844 15896 12850
rect 15844 12786 15896 12792
rect 15856 12617 15884 12786
rect 15842 12608 15898 12617
rect 15842 12543 15898 12552
rect 15948 12458 15976 14826
rect 16040 14278 16068 14962
rect 16132 14550 16160 15438
rect 16224 15094 16252 17682
rect 16316 17678 16344 17711
rect 16304 17672 16356 17678
rect 16304 17614 16356 17620
rect 16304 17536 16356 17542
rect 16304 17478 16356 17484
rect 16316 16590 16344 17478
rect 16408 17134 16436 19887
rect 16396 17128 16448 17134
rect 16396 17070 16448 17076
rect 16304 16584 16356 16590
rect 16304 16526 16356 16532
rect 16396 15496 16448 15502
rect 16396 15438 16448 15444
rect 16212 15088 16264 15094
rect 16212 15030 16264 15036
rect 16302 15056 16358 15065
rect 16120 14544 16172 14550
rect 16120 14486 16172 14492
rect 16224 14346 16252 15030
rect 16302 14991 16358 15000
rect 16212 14340 16264 14346
rect 16212 14282 16264 14288
rect 16028 14272 16080 14278
rect 16080 14220 16160 14226
rect 16028 14214 16160 14220
rect 16040 14198 16160 14214
rect 16028 13932 16080 13938
rect 16028 13874 16080 13880
rect 16040 12986 16068 13874
rect 16132 13326 16160 14198
rect 16212 14068 16264 14074
rect 16212 14010 16264 14016
rect 16120 13320 16172 13326
rect 16120 13262 16172 13268
rect 16028 12980 16080 12986
rect 16028 12922 16080 12928
rect 15396 12406 15516 12434
rect 15856 12430 15976 12458
rect 15292 12300 15344 12306
rect 15292 12242 15344 12248
rect 15200 12096 15252 12102
rect 15200 12038 15252 12044
rect 15108 11892 15160 11898
rect 15108 11834 15160 11840
rect 14924 11756 14976 11762
rect 14924 11698 14976 11704
rect 14832 11688 14884 11694
rect 14832 11630 14884 11636
rect 14844 11354 14872 11630
rect 14832 11348 14884 11354
rect 14832 11290 14884 11296
rect 14936 11218 14964 11698
rect 15108 11552 15160 11558
rect 15028 11500 15108 11506
rect 15028 11494 15160 11500
rect 15028 11478 15148 11494
rect 14924 11212 14976 11218
rect 14924 11154 14976 11160
rect 14936 10606 14964 11154
rect 15028 10810 15056 11478
rect 15212 11150 15240 12038
rect 15200 11144 15252 11150
rect 15200 11086 15252 11092
rect 15292 11076 15344 11082
rect 15292 11018 15344 11024
rect 15304 10810 15332 11018
rect 15016 10804 15068 10810
rect 15016 10746 15068 10752
rect 15292 10804 15344 10810
rect 15292 10746 15344 10752
rect 15396 10656 15424 12406
rect 15476 12232 15528 12238
rect 15474 12200 15476 12209
rect 15660 12232 15712 12238
rect 15528 12200 15530 12209
rect 15660 12174 15712 12180
rect 15752 12232 15804 12238
rect 15856 12220 15884 12430
rect 15936 12300 15988 12306
rect 15936 12242 15988 12248
rect 15804 12192 15884 12220
rect 15752 12174 15804 12180
rect 15474 12135 15530 12144
rect 15568 12096 15620 12102
rect 15568 12038 15620 12044
rect 15580 11801 15608 12038
rect 15566 11792 15622 11801
rect 15566 11727 15622 11736
rect 15476 10668 15528 10674
rect 15396 10628 15476 10656
rect 15476 10610 15528 10616
rect 14832 10600 14884 10606
rect 14832 10542 14884 10548
rect 14924 10600 14976 10606
rect 14924 10542 14976 10548
rect 14844 9926 14872 10542
rect 15200 10464 15252 10470
rect 15200 10406 15252 10412
rect 15212 10305 15240 10406
rect 15198 10296 15254 10305
rect 15198 10231 15254 10240
rect 15292 10260 15344 10266
rect 15292 10202 15344 10208
rect 14832 9920 14884 9926
rect 14832 9862 14884 9868
rect 14844 9654 14872 9862
rect 14832 9648 14884 9654
rect 14832 9590 14884 9596
rect 14740 9580 14792 9586
rect 14740 9522 14792 9528
rect 15016 9580 15068 9586
rect 15016 9522 15068 9528
rect 14384 9438 14504 9466
rect 14554 9480 14610 9489
rect 14384 8362 14412 9438
rect 14554 9415 14556 9424
rect 14608 9415 14610 9424
rect 14556 9386 14608 9392
rect 14464 9376 14516 9382
rect 14464 9318 14516 9324
rect 14648 9376 14700 9382
rect 14648 9318 14700 9324
rect 14476 9110 14504 9318
rect 14464 9104 14516 9110
rect 14464 9046 14516 9052
rect 14660 8566 14688 9318
rect 14648 8560 14700 8566
rect 14648 8502 14700 8508
rect 14372 8356 14424 8362
rect 14372 8298 14424 8304
rect 14384 7886 14412 8298
rect 14280 7880 14332 7886
rect 14280 7822 14332 7828
rect 14372 7880 14424 7886
rect 14464 7880 14516 7886
rect 14372 7822 14424 7828
rect 14462 7848 14464 7857
rect 14516 7848 14518 7857
rect 14752 7834 14780 9522
rect 14924 8968 14976 8974
rect 14924 8910 14976 8916
rect 14832 8832 14884 8838
rect 14832 8774 14884 8780
rect 14936 8786 14964 8910
rect 15028 8906 15056 9522
rect 15200 8968 15252 8974
rect 15120 8916 15200 8922
rect 15304 8945 15332 10202
rect 15384 8968 15436 8974
rect 15120 8910 15252 8916
rect 15290 8936 15346 8945
rect 15016 8900 15068 8906
rect 15016 8842 15068 8848
rect 15120 8894 15240 8910
rect 14844 8566 14872 8774
rect 14936 8758 15056 8786
rect 14832 8560 14884 8566
rect 14832 8502 14884 8508
rect 14924 8424 14976 8430
rect 14924 8366 14976 8372
rect 14832 8016 14884 8022
rect 14832 7958 14884 7964
rect 14004 6792 14056 6798
rect 14004 6734 14056 6740
rect 14188 6792 14240 6798
rect 14188 6734 14240 6740
rect 13912 6316 13964 6322
rect 13832 6276 13912 6304
rect 13544 6258 13596 6264
rect 13912 6258 13964 6264
rect 13556 5642 13584 6258
rect 13636 6248 13688 6254
rect 13688 6196 13860 6202
rect 13636 6190 13860 6196
rect 13648 6174 13860 6190
rect 13832 6118 13860 6174
rect 13728 6112 13780 6118
rect 13728 6054 13780 6060
rect 13820 6112 13872 6118
rect 13820 6054 13872 6060
rect 13544 5636 13596 5642
rect 13544 5578 13596 5584
rect 13636 5568 13688 5574
rect 13636 5510 13688 5516
rect 13360 5296 13412 5302
rect 13360 5238 13412 5244
rect 13648 5098 13676 5510
rect 13740 5250 13768 6054
rect 13924 5778 13952 6258
rect 14016 6254 14044 6734
rect 14004 6248 14056 6254
rect 14004 6190 14056 6196
rect 14096 6248 14148 6254
rect 14096 6190 14148 6196
rect 13912 5772 13964 5778
rect 13912 5714 13964 5720
rect 13820 5636 13872 5642
rect 13820 5578 13872 5584
rect 13832 5409 13860 5578
rect 13818 5400 13874 5409
rect 13818 5335 13874 5344
rect 13820 5296 13872 5302
rect 13740 5244 13820 5250
rect 13740 5238 13872 5244
rect 13740 5222 13860 5238
rect 13912 5228 13964 5234
rect 13912 5170 13964 5176
rect 13924 5098 13952 5170
rect 13636 5092 13688 5098
rect 13636 5034 13688 5040
rect 13912 5092 13964 5098
rect 13912 5034 13964 5040
rect 13360 5024 13412 5030
rect 13360 4966 13412 4972
rect 13372 4146 13400 4966
rect 13820 4208 13872 4214
rect 13820 4150 13872 4156
rect 13360 4140 13412 4146
rect 13360 4082 13412 4088
rect 13084 3528 13136 3534
rect 13084 3470 13136 3476
rect 12440 3460 12492 3466
rect 12440 3402 12492 3408
rect 13832 3126 13860 4150
rect 13924 3670 13952 5034
rect 13912 3664 13964 3670
rect 13912 3606 13964 3612
rect 13912 3460 13964 3466
rect 13912 3402 13964 3408
rect 13924 3194 13952 3402
rect 13912 3188 13964 3194
rect 13912 3130 13964 3136
rect 11980 3120 12032 3126
rect 11980 3062 12032 3068
rect 13820 3120 13872 3126
rect 13820 3062 13872 3068
rect 10876 2984 10928 2990
rect 10876 2926 10928 2932
rect 10968 2984 11020 2990
rect 10968 2926 11020 2932
rect 10888 2582 10916 2926
rect 13820 2916 13872 2922
rect 13820 2858 13872 2864
rect 10876 2576 10928 2582
rect 10876 2518 10928 2524
rect 9312 2508 9364 2514
rect 9312 2450 9364 2456
rect 13832 2446 13860 2858
rect 13924 2446 13952 3130
rect 14016 2446 14044 6190
rect 14108 5914 14136 6190
rect 14096 5908 14148 5914
rect 14096 5850 14148 5856
rect 14200 5846 14228 6734
rect 14292 6458 14320 7822
rect 14462 7783 14518 7792
rect 14660 7806 14780 7834
rect 14556 7200 14608 7206
rect 14556 7142 14608 7148
rect 14464 6996 14516 7002
rect 14464 6938 14516 6944
rect 14476 6905 14504 6938
rect 14462 6896 14518 6905
rect 14462 6831 14518 6840
rect 14568 6730 14596 7142
rect 14660 6798 14688 7806
rect 14844 7750 14872 7958
rect 14936 7954 14964 8366
rect 14924 7948 14976 7954
rect 14924 7890 14976 7896
rect 14740 7744 14792 7750
rect 14740 7686 14792 7692
rect 14832 7744 14884 7750
rect 14832 7686 14884 7692
rect 14752 7410 14780 7686
rect 14936 7478 14964 7890
rect 15028 7750 15056 8758
rect 15120 7818 15148 8894
rect 15384 8910 15436 8916
rect 15290 8871 15346 8880
rect 15200 8288 15252 8294
rect 15200 8230 15252 8236
rect 15212 7886 15240 8230
rect 15200 7880 15252 7886
rect 15200 7822 15252 7828
rect 15108 7812 15160 7818
rect 15108 7754 15160 7760
rect 15016 7744 15068 7750
rect 15016 7686 15068 7692
rect 14924 7472 14976 7478
rect 14924 7414 14976 7420
rect 14740 7404 14792 7410
rect 14740 7346 14792 7352
rect 14936 6866 14964 7414
rect 14924 6860 14976 6866
rect 14924 6802 14976 6808
rect 14648 6792 14700 6798
rect 14648 6734 14700 6740
rect 14372 6724 14424 6730
rect 14372 6666 14424 6672
rect 14556 6724 14608 6730
rect 14556 6666 14608 6672
rect 14280 6452 14332 6458
rect 14280 6394 14332 6400
rect 14384 6322 14412 6666
rect 14464 6656 14516 6662
rect 14464 6598 14516 6604
rect 14476 6390 14504 6598
rect 14660 6390 14688 6734
rect 14464 6384 14516 6390
rect 14464 6326 14516 6332
rect 14648 6384 14700 6390
rect 14648 6326 14700 6332
rect 14372 6316 14424 6322
rect 14372 6258 14424 6264
rect 14556 6316 14608 6322
rect 14556 6258 14608 6264
rect 14188 5840 14240 5846
rect 14188 5782 14240 5788
rect 14188 5704 14240 5710
rect 14240 5664 14504 5692
rect 14188 5646 14240 5652
rect 14188 5568 14240 5574
rect 14372 5568 14424 5574
rect 14240 5528 14372 5556
rect 14188 5510 14240 5516
rect 14188 5160 14240 5166
rect 14188 5102 14240 5108
rect 14200 3738 14228 5102
rect 14292 4826 14320 5528
rect 14372 5510 14424 5516
rect 14372 5228 14424 5234
rect 14372 5170 14424 5176
rect 14384 5030 14412 5170
rect 14372 5024 14424 5030
rect 14372 4966 14424 4972
rect 14280 4820 14332 4826
rect 14280 4762 14332 4768
rect 14372 4616 14424 4622
rect 14372 4558 14424 4564
rect 14188 3732 14240 3738
rect 14188 3674 14240 3680
rect 14096 3392 14148 3398
rect 14096 3334 14148 3340
rect 14108 3058 14136 3334
rect 14200 3058 14228 3674
rect 14384 3534 14412 4558
rect 14476 3942 14504 5664
rect 14568 5642 14596 6258
rect 14660 5710 14688 6326
rect 14738 6080 14794 6089
rect 14738 6015 14794 6024
rect 14752 5846 14780 6015
rect 14740 5840 14792 5846
rect 14740 5782 14792 5788
rect 14648 5704 14700 5710
rect 14648 5646 14700 5652
rect 14738 5672 14794 5681
rect 14556 5636 14608 5642
rect 14738 5607 14740 5616
rect 14556 5578 14608 5584
rect 14792 5607 14794 5616
rect 14740 5578 14792 5584
rect 14832 5568 14884 5574
rect 14832 5510 14884 5516
rect 14844 5250 14872 5510
rect 14568 5222 14872 5250
rect 14464 3936 14516 3942
rect 14464 3878 14516 3884
rect 14280 3528 14332 3534
rect 14280 3470 14332 3476
rect 14372 3528 14424 3534
rect 14372 3470 14424 3476
rect 14292 3058 14320 3470
rect 14096 3052 14148 3058
rect 14096 2994 14148 3000
rect 14188 3052 14240 3058
rect 14188 2994 14240 3000
rect 14280 3052 14332 3058
rect 14280 2994 14332 3000
rect 14476 2922 14504 3878
rect 14568 3194 14596 5222
rect 14648 5160 14700 5166
rect 14648 5102 14700 5108
rect 14660 4622 14688 5102
rect 14740 5024 14792 5030
rect 14740 4966 14792 4972
rect 14648 4616 14700 4622
rect 14648 4558 14700 4564
rect 14752 4554 14780 4966
rect 14936 4622 14964 6802
rect 15014 6352 15070 6361
rect 15014 6287 15016 6296
rect 15068 6287 15070 6296
rect 15016 6256 15068 6262
rect 15016 6112 15068 6118
rect 15016 6054 15068 6060
rect 15028 5642 15056 6054
rect 15016 5636 15068 5642
rect 15016 5578 15068 5584
rect 14924 4616 14976 4622
rect 14924 4558 14976 4564
rect 14740 4548 14792 4554
rect 14740 4490 14792 4496
rect 14936 4214 14964 4558
rect 14924 4208 14976 4214
rect 14924 4150 14976 4156
rect 14738 4040 14794 4049
rect 14738 3975 14794 3984
rect 14556 3188 14608 3194
rect 14556 3130 14608 3136
rect 14752 3126 14780 3975
rect 14936 3602 14964 4150
rect 15028 4010 15056 5578
rect 15120 5234 15148 7754
rect 15198 6896 15254 6905
rect 15198 6831 15254 6840
rect 15212 6458 15240 6831
rect 15290 6624 15346 6633
rect 15290 6559 15346 6568
rect 15200 6452 15252 6458
rect 15200 6394 15252 6400
rect 15209 6316 15261 6322
rect 15304 6304 15332 6559
rect 15396 6361 15424 8910
rect 15261 6276 15332 6304
rect 15382 6352 15438 6361
rect 15382 6287 15438 6296
rect 15209 6258 15261 6264
rect 15198 6216 15254 6225
rect 15198 6151 15200 6160
rect 15252 6151 15254 6160
rect 15200 6122 15252 6128
rect 15304 5846 15332 6276
rect 15292 5840 15344 5846
rect 15292 5782 15344 5788
rect 15292 5568 15344 5574
rect 15292 5510 15344 5516
rect 15198 5400 15254 5409
rect 15198 5335 15254 5344
rect 15212 5234 15240 5335
rect 15108 5228 15160 5234
rect 15108 5170 15160 5176
rect 15200 5228 15252 5234
rect 15200 5170 15252 5176
rect 15120 5098 15148 5170
rect 15108 5092 15160 5098
rect 15108 5034 15160 5040
rect 15198 4176 15254 4185
rect 15198 4111 15254 4120
rect 15016 4004 15068 4010
rect 15016 3946 15068 3952
rect 14924 3596 14976 3602
rect 14924 3538 14976 3544
rect 14830 3496 14886 3505
rect 14830 3431 14886 3440
rect 14740 3120 14792 3126
rect 14740 3062 14792 3068
rect 14556 3052 14608 3058
rect 14556 2994 14608 3000
rect 14464 2916 14516 2922
rect 14464 2858 14516 2864
rect 14568 2582 14596 2994
rect 14752 2854 14780 3062
rect 14648 2848 14700 2854
rect 14648 2790 14700 2796
rect 14740 2848 14792 2854
rect 14740 2790 14792 2796
rect 14556 2576 14608 2582
rect 14556 2518 14608 2524
rect 14660 2446 14688 2790
rect 14752 2446 14780 2790
rect 14844 2650 14872 3431
rect 14936 3058 14964 3538
rect 14924 3052 14976 3058
rect 14924 2994 14976 3000
rect 15212 2650 15240 4111
rect 15304 3126 15332 5510
rect 15396 5370 15424 6287
rect 15488 5817 15516 10610
rect 15580 9926 15608 11727
rect 15568 9920 15620 9926
rect 15568 9862 15620 9868
rect 15672 9654 15700 12174
rect 15764 11014 15792 12174
rect 15948 11286 15976 12242
rect 16028 12164 16080 12170
rect 16028 12106 16080 12112
rect 16040 11558 16068 12106
rect 16028 11552 16080 11558
rect 16028 11494 16080 11500
rect 15936 11280 15988 11286
rect 15936 11222 15988 11228
rect 15752 11008 15804 11014
rect 15752 10950 15804 10956
rect 15844 10804 15896 10810
rect 15844 10746 15896 10752
rect 15750 10160 15806 10169
rect 15750 10095 15806 10104
rect 15660 9648 15712 9654
rect 15660 9590 15712 9596
rect 15764 8974 15792 10095
rect 15856 8974 15884 10746
rect 15948 9518 15976 11222
rect 16132 10062 16160 13262
rect 16224 13025 16252 14010
rect 16210 13016 16266 13025
rect 16210 12951 16266 12960
rect 16212 12096 16264 12102
rect 16212 12038 16264 12044
rect 16224 11354 16252 12038
rect 16212 11348 16264 11354
rect 16212 11290 16264 11296
rect 16210 10976 16266 10985
rect 16210 10911 16266 10920
rect 16120 10056 16172 10062
rect 16120 9998 16172 10004
rect 16120 9920 16172 9926
rect 16120 9862 16172 9868
rect 16132 9654 16160 9862
rect 16120 9648 16172 9654
rect 16120 9590 16172 9596
rect 16028 9580 16080 9586
rect 16028 9522 16080 9528
rect 15936 9512 15988 9518
rect 15936 9454 15988 9460
rect 15752 8968 15804 8974
rect 15752 8910 15804 8916
rect 15844 8968 15896 8974
rect 15844 8910 15896 8916
rect 15764 8634 15792 8910
rect 15936 8900 15988 8906
rect 15936 8842 15988 8848
rect 15752 8628 15804 8634
rect 15752 8570 15804 8576
rect 15752 8492 15804 8498
rect 15752 8434 15804 8440
rect 15568 6724 15620 6730
rect 15568 6666 15620 6672
rect 15580 6458 15608 6666
rect 15658 6488 15714 6497
rect 15568 6452 15620 6458
rect 15658 6423 15660 6432
rect 15568 6394 15620 6400
rect 15712 6423 15714 6432
rect 15660 6394 15712 6400
rect 15764 6322 15792 8434
rect 15948 6662 15976 8842
rect 16040 8090 16068 9522
rect 16132 8906 16160 9590
rect 16224 9178 16252 10911
rect 16316 10266 16344 14991
rect 16408 12170 16436 15438
rect 16396 12164 16448 12170
rect 16396 12106 16448 12112
rect 16304 10260 16356 10266
rect 16304 10202 16356 10208
rect 16212 9172 16264 9178
rect 16212 9114 16264 9120
rect 16120 8900 16172 8906
rect 16120 8842 16172 8848
rect 16210 8256 16266 8265
rect 16210 8191 16266 8200
rect 16028 8084 16080 8090
rect 16028 8026 16080 8032
rect 16040 7410 16068 8026
rect 16224 7546 16252 8191
rect 16304 7744 16356 7750
rect 16304 7686 16356 7692
rect 16212 7540 16264 7546
rect 16212 7482 16264 7488
rect 16028 7404 16080 7410
rect 16028 7346 16080 7352
rect 15936 6656 15988 6662
rect 15936 6598 15988 6604
rect 16040 6458 16068 7346
rect 16212 6656 16264 6662
rect 16212 6598 16264 6604
rect 16028 6452 16080 6458
rect 16028 6394 16080 6400
rect 16224 6322 16252 6598
rect 15752 6316 15804 6322
rect 15752 6258 15804 6264
rect 16028 6316 16080 6322
rect 16028 6258 16080 6264
rect 16212 6316 16264 6322
rect 16212 6258 16264 6264
rect 16040 5914 16068 6258
rect 16224 5953 16252 6258
rect 16210 5944 16266 5953
rect 16028 5908 16080 5914
rect 16210 5879 16266 5888
rect 16028 5850 16080 5856
rect 15474 5808 15530 5817
rect 15474 5743 15530 5752
rect 15658 5808 15714 5817
rect 15658 5743 15714 5752
rect 15672 5710 15700 5743
rect 15660 5704 15712 5710
rect 15660 5646 15712 5652
rect 15844 5704 15896 5710
rect 15844 5646 15896 5652
rect 15936 5704 15988 5710
rect 15936 5646 15988 5652
rect 16120 5704 16172 5710
rect 16120 5646 16172 5652
rect 15384 5364 15436 5370
rect 15384 5306 15436 5312
rect 15396 5234 15424 5306
rect 15384 5228 15436 5234
rect 15384 5170 15436 5176
rect 15396 5030 15424 5170
rect 15384 5024 15436 5030
rect 15384 4966 15436 4972
rect 15476 5024 15528 5030
rect 15476 4966 15528 4972
rect 15488 4146 15516 4966
rect 15856 4758 15884 5646
rect 15844 4752 15896 4758
rect 15844 4694 15896 4700
rect 15568 4480 15620 4486
rect 15568 4422 15620 4428
rect 15476 4140 15528 4146
rect 15476 4082 15528 4088
rect 15580 3534 15608 4422
rect 15658 4040 15714 4049
rect 15658 3975 15714 3984
rect 15672 3738 15700 3975
rect 15660 3732 15712 3738
rect 15660 3674 15712 3680
rect 15568 3528 15620 3534
rect 15568 3470 15620 3476
rect 15292 3120 15344 3126
rect 15292 3062 15344 3068
rect 14832 2644 14884 2650
rect 14832 2586 14884 2592
rect 15200 2644 15252 2650
rect 15200 2586 15252 2592
rect 15672 2446 15700 3674
rect 15856 3466 15884 4694
rect 15844 3460 15896 3466
rect 15844 3402 15896 3408
rect 15948 3194 15976 5646
rect 16132 5234 16160 5646
rect 16120 5228 16172 5234
rect 16120 5170 16172 5176
rect 16132 4622 16160 5170
rect 16210 4856 16266 4865
rect 16210 4791 16266 4800
rect 16028 4616 16080 4622
rect 16028 4558 16080 4564
rect 16120 4616 16172 4622
rect 16120 4558 16172 4564
rect 15936 3188 15988 3194
rect 15936 3130 15988 3136
rect 16040 2650 16068 4558
rect 16224 2650 16252 4791
rect 16316 4554 16344 7686
rect 16304 4548 16356 4554
rect 16304 4490 16356 4496
rect 16028 2644 16080 2650
rect 16028 2586 16080 2592
rect 16212 2644 16264 2650
rect 16212 2586 16264 2592
rect 7104 2440 7156 2446
rect 7104 2382 7156 2388
rect 8760 2440 8812 2446
rect 8760 2382 8812 2388
rect 9220 2440 9272 2446
rect 9220 2382 9272 2388
rect 13820 2440 13872 2446
rect 13820 2382 13872 2388
rect 13912 2440 13964 2446
rect 13912 2382 13964 2388
rect 14004 2440 14056 2446
rect 14004 2382 14056 2388
rect 14648 2440 14700 2446
rect 14648 2382 14700 2388
rect 14740 2440 14792 2446
rect 14740 2382 14792 2388
rect 15660 2440 15712 2446
rect 15660 2382 15712 2388
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 7116 800 7144 2382
rect 7748 2372 7800 2378
rect 7748 2314 7800 2320
rect 9680 2372 9732 2378
rect 9680 2314 9732 2320
rect 7760 800 7788 2314
rect 8392 2304 8444 2310
rect 8392 2246 8444 2252
rect 9036 2304 9088 2310
rect 9036 2246 9088 2252
rect 8404 800 8432 2246
rect 9048 800 9076 2246
rect 9692 800 9720 2314
rect 12900 2304 12952 2310
rect 12900 2246 12952 2252
rect 13544 2304 13596 2310
rect 13544 2246 13596 2252
rect 14188 2304 14240 2310
rect 14188 2246 14240 2252
rect 12912 800 12940 2246
rect 13556 800 13584 2246
rect 14200 800 14228 2246
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 9034 0 9090 800
rect 9678 0 9734 800
rect 12898 0 12954 800
rect 13542 0 13598 800
rect 14186 0 14242 800
<< via2 >>
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4880 32666 4936 32668
rect 4960 32666 5016 32668
rect 5040 32666 5096 32668
rect 5120 32666 5176 32668
rect 4880 32614 4926 32666
rect 4926 32614 4936 32666
rect 4960 32614 4990 32666
rect 4990 32614 5002 32666
rect 5002 32614 5016 32666
rect 5040 32614 5054 32666
rect 5054 32614 5066 32666
rect 5066 32614 5096 32666
rect 5120 32614 5130 32666
rect 5130 32614 5176 32666
rect 4880 32612 4936 32614
rect 4960 32612 5016 32614
rect 5040 32612 5096 32614
rect 5120 32612 5176 32614
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 7010 31864 7066 31920
rect 4880 31578 4936 31580
rect 4960 31578 5016 31580
rect 5040 31578 5096 31580
rect 5120 31578 5176 31580
rect 4880 31526 4926 31578
rect 4926 31526 4936 31578
rect 4960 31526 4990 31578
rect 4990 31526 5002 31578
rect 5002 31526 5016 31578
rect 5040 31526 5054 31578
rect 5054 31526 5066 31578
rect 5066 31526 5096 31578
rect 5120 31526 5130 31578
rect 5130 31526 5176 31578
rect 4880 31524 4936 31526
rect 4960 31524 5016 31526
rect 5040 31524 5096 31526
rect 5120 31524 5176 31526
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 7194 31728 7250 31784
rect 4880 30490 4936 30492
rect 4960 30490 5016 30492
rect 5040 30490 5096 30492
rect 5120 30490 5176 30492
rect 4880 30438 4926 30490
rect 4926 30438 4936 30490
rect 4960 30438 4990 30490
rect 4990 30438 5002 30490
rect 5002 30438 5016 30490
rect 5040 30438 5054 30490
rect 5054 30438 5066 30490
rect 5066 30438 5096 30490
rect 5120 30438 5130 30490
rect 5130 30438 5176 30490
rect 4880 30436 4936 30438
rect 4960 30436 5016 30438
rect 5040 30436 5096 30438
rect 5120 30436 5176 30438
rect 110 30096 166 30152
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4880 29402 4936 29404
rect 4960 29402 5016 29404
rect 5040 29402 5096 29404
rect 5120 29402 5176 29404
rect 4880 29350 4926 29402
rect 4926 29350 4936 29402
rect 4960 29350 4990 29402
rect 4990 29350 5002 29402
rect 5002 29350 5016 29402
rect 5040 29350 5054 29402
rect 5054 29350 5066 29402
rect 5066 29350 5096 29402
rect 5120 29350 5130 29402
rect 5130 29350 5176 29402
rect 4880 29348 4936 29350
rect 4960 29348 5016 29350
rect 5040 29348 5096 29350
rect 5120 29348 5176 29350
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 6918 29688 6974 29744
rect 7286 29688 7342 29744
rect 846 25336 902 25392
rect 846 21256 902 21312
rect 2778 27004 2780 27024
rect 2780 27004 2832 27024
rect 2832 27004 2834 27024
rect 2594 26424 2650 26480
rect 2778 26968 2834 27004
rect 4880 28314 4936 28316
rect 4960 28314 5016 28316
rect 5040 28314 5096 28316
rect 5120 28314 5176 28316
rect 4880 28262 4926 28314
rect 4926 28262 4936 28314
rect 4960 28262 4990 28314
rect 4990 28262 5002 28314
rect 5002 28262 5016 28314
rect 5040 28262 5054 28314
rect 5054 28262 5066 28314
rect 5066 28262 5096 28314
rect 5120 28262 5130 28314
rect 5130 28262 5176 28314
rect 4880 28260 4936 28262
rect 4960 28260 5016 28262
rect 5040 28260 5096 28262
rect 5120 28260 5176 28262
rect 2870 26832 2926 26888
rect 2778 26424 2834 26480
rect 3054 26696 3110 26752
rect 3514 26696 3570 26752
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 3422 24148 3424 24168
rect 3424 24148 3476 24168
rect 3476 24148 3478 24168
rect 3422 24112 3478 24148
rect 2226 20868 2282 20904
rect 2226 20848 2228 20868
rect 2228 20848 2280 20868
rect 2280 20848 2282 20868
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4880 27226 4936 27228
rect 4960 27226 5016 27228
rect 5040 27226 5096 27228
rect 5120 27226 5176 27228
rect 4880 27174 4926 27226
rect 4926 27174 4936 27226
rect 4960 27174 4990 27226
rect 4990 27174 5002 27226
rect 5002 27174 5016 27226
rect 5040 27174 5054 27226
rect 5054 27174 5066 27226
rect 5066 27174 5096 27226
rect 5120 27174 5130 27226
rect 5130 27174 5176 27226
rect 4880 27172 4936 27174
rect 4960 27172 5016 27174
rect 5040 27172 5096 27174
rect 5120 27172 5176 27174
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4802 26968 4858 27024
rect 5078 26832 5134 26888
rect 4880 26138 4936 26140
rect 4960 26138 5016 26140
rect 5040 26138 5096 26140
rect 5120 26138 5176 26140
rect 4880 26086 4926 26138
rect 4926 26086 4936 26138
rect 4960 26086 4990 26138
rect 4990 26086 5002 26138
rect 5002 26086 5016 26138
rect 5040 26086 5054 26138
rect 5054 26086 5066 26138
rect 5066 26086 5096 26138
rect 5120 26086 5130 26138
rect 5130 26086 5176 26138
rect 4880 26084 4936 26086
rect 4960 26084 5016 26086
rect 5040 26084 5096 26086
rect 5120 26084 5176 26086
rect 4880 25050 4936 25052
rect 4960 25050 5016 25052
rect 5040 25050 5096 25052
rect 5120 25050 5176 25052
rect 4880 24998 4926 25050
rect 4926 24998 4936 25050
rect 4960 24998 4990 25050
rect 4990 24998 5002 25050
rect 5002 24998 5016 25050
rect 5040 24998 5054 25050
rect 5054 24998 5066 25050
rect 5066 24998 5096 25050
rect 5120 24998 5130 25050
rect 5130 24998 5176 25050
rect 4880 24996 4936 24998
rect 4960 24996 5016 24998
rect 5040 24996 5096 24998
rect 5120 24996 5176 24998
rect 3974 24284 3976 24304
rect 3976 24284 4028 24304
rect 4028 24284 4030 24304
rect 3974 24248 4030 24284
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 2870 20884 2872 20904
rect 2872 20884 2924 20904
rect 2924 20884 2926 20904
rect 2870 20848 2926 20884
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 5906 26968 5962 27024
rect 4880 23962 4936 23964
rect 4960 23962 5016 23964
rect 5040 23962 5096 23964
rect 5120 23962 5176 23964
rect 4880 23910 4926 23962
rect 4926 23910 4936 23962
rect 4960 23910 4990 23962
rect 4990 23910 5002 23962
rect 5002 23910 5016 23962
rect 5040 23910 5054 23962
rect 5054 23910 5066 23962
rect 5066 23910 5096 23962
rect 5120 23910 5130 23962
rect 5130 23910 5176 23962
rect 4880 23908 4936 23910
rect 4960 23908 5016 23910
rect 5040 23908 5096 23910
rect 5120 23908 5176 23910
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 2410 17620 2412 17640
rect 2412 17620 2464 17640
rect 2464 17620 2466 17640
rect 2410 17584 2466 17620
rect 4880 22874 4936 22876
rect 4960 22874 5016 22876
rect 5040 22874 5096 22876
rect 5120 22874 5176 22876
rect 4880 22822 4926 22874
rect 4926 22822 4936 22874
rect 4960 22822 4990 22874
rect 4990 22822 5002 22874
rect 5002 22822 5016 22874
rect 5040 22822 5054 22874
rect 5054 22822 5066 22874
rect 5066 22822 5096 22874
rect 5120 22822 5130 22874
rect 5130 22822 5176 22874
rect 4880 22820 4936 22822
rect 4960 22820 5016 22822
rect 5040 22820 5096 22822
rect 5120 22820 5176 22822
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4158 20576 4214 20632
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4250 19216 4306 19272
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 3146 17196 3202 17232
rect 3146 17176 3148 17196
rect 3148 17176 3200 17196
rect 3200 17176 3202 17196
rect 2686 15544 2742 15600
rect 2870 15680 2926 15736
rect 2870 12008 2926 12064
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4880 21786 4936 21788
rect 4960 21786 5016 21788
rect 5040 21786 5096 21788
rect 5120 21786 5176 21788
rect 4880 21734 4926 21786
rect 4926 21734 4936 21786
rect 4960 21734 4990 21786
rect 4990 21734 5002 21786
rect 5002 21734 5016 21786
rect 5040 21734 5054 21786
rect 5054 21734 5066 21786
rect 5066 21734 5096 21786
rect 5120 21734 5130 21786
rect 5130 21734 5176 21786
rect 4880 21732 4936 21734
rect 4960 21732 5016 21734
rect 5040 21732 5096 21734
rect 5120 21732 5176 21734
rect 4880 20698 4936 20700
rect 4960 20698 5016 20700
rect 5040 20698 5096 20700
rect 5120 20698 5176 20700
rect 4880 20646 4926 20698
rect 4926 20646 4936 20698
rect 4960 20646 4990 20698
rect 4990 20646 5002 20698
rect 5002 20646 5016 20698
rect 5040 20646 5054 20698
rect 5054 20646 5066 20698
rect 5066 20646 5096 20698
rect 5120 20646 5130 20698
rect 5130 20646 5176 20698
rect 4880 20644 4936 20646
rect 4960 20644 5016 20646
rect 5040 20644 5096 20646
rect 5120 20644 5176 20646
rect 5170 19760 5226 19816
rect 4880 19610 4936 19612
rect 4960 19610 5016 19612
rect 5040 19610 5096 19612
rect 5120 19610 5176 19612
rect 4880 19558 4926 19610
rect 4926 19558 4936 19610
rect 4960 19558 4990 19610
rect 4990 19558 5002 19610
rect 5002 19558 5016 19610
rect 5040 19558 5054 19610
rect 5054 19558 5066 19610
rect 5066 19558 5096 19610
rect 5120 19558 5130 19610
rect 5130 19558 5176 19610
rect 4880 19556 4936 19558
rect 4960 19556 5016 19558
rect 5040 19556 5096 19558
rect 5120 19556 5176 19558
rect 5354 19760 5410 19816
rect 3238 15544 3294 15600
rect 3146 15408 3202 15464
rect 3882 17620 3884 17640
rect 3884 17620 3936 17640
rect 3936 17620 3938 17640
rect 3882 17584 3938 17620
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4066 15444 4068 15464
rect 4068 15444 4120 15464
rect 4120 15444 4122 15464
rect 4066 15408 4122 15444
rect 3606 13932 3662 13968
rect 3606 13912 3608 13932
rect 3608 13912 3660 13932
rect 3660 13912 3662 13932
rect 3422 13368 3478 13424
rect 3606 13640 3662 13696
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 5170 19372 5226 19408
rect 5170 19352 5172 19372
rect 5172 19352 5224 19372
rect 5224 19352 5226 19372
rect 4880 18522 4936 18524
rect 4960 18522 5016 18524
rect 5040 18522 5096 18524
rect 5120 18522 5176 18524
rect 4880 18470 4926 18522
rect 4926 18470 4936 18522
rect 4960 18470 4990 18522
rect 4990 18470 5002 18522
rect 5002 18470 5016 18522
rect 5040 18470 5054 18522
rect 5054 18470 5066 18522
rect 5066 18470 5096 18522
rect 5120 18470 5130 18522
rect 5130 18470 5176 18522
rect 4880 18468 4936 18470
rect 4960 18468 5016 18470
rect 5040 18468 5096 18470
rect 5120 18468 5176 18470
rect 5998 19352 6054 19408
rect 4880 17434 4936 17436
rect 4960 17434 5016 17436
rect 5040 17434 5096 17436
rect 5120 17434 5176 17436
rect 4880 17382 4926 17434
rect 4926 17382 4936 17434
rect 4960 17382 4990 17434
rect 4990 17382 5002 17434
rect 5002 17382 5016 17434
rect 5040 17382 5054 17434
rect 5054 17382 5066 17434
rect 5066 17382 5096 17434
rect 5120 17382 5130 17434
rect 5130 17382 5176 17434
rect 4880 17380 4936 17382
rect 4960 17380 5016 17382
rect 5040 17380 5096 17382
rect 5120 17380 5176 17382
rect 4880 16346 4936 16348
rect 4960 16346 5016 16348
rect 5040 16346 5096 16348
rect 5120 16346 5176 16348
rect 4880 16294 4926 16346
rect 4926 16294 4936 16346
rect 4960 16294 4990 16346
rect 4990 16294 5002 16346
rect 5002 16294 5016 16346
rect 5040 16294 5054 16346
rect 5054 16294 5066 16346
rect 5066 16294 5096 16346
rect 5120 16294 5130 16346
rect 5130 16294 5176 16346
rect 4880 16292 4936 16294
rect 4960 16292 5016 16294
rect 5040 16292 5096 16294
rect 5120 16292 5176 16294
rect 3882 13368 3938 13424
rect 3422 12300 3478 12336
rect 3422 12280 3424 12300
rect 3424 12280 3476 12300
rect 3476 12280 3478 12300
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4250 13404 4252 13424
rect 4252 13404 4304 13424
rect 4304 13404 4306 13424
rect 4250 13368 4306 13404
rect 4250 13268 4252 13288
rect 4252 13268 4304 13288
rect 4304 13268 4306 13288
rect 4250 13232 4306 13268
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4894 15444 4896 15464
rect 4896 15444 4948 15464
rect 4948 15444 4950 15464
rect 4894 15408 4950 15444
rect 5170 15544 5226 15600
rect 5078 15408 5134 15464
rect 4880 15258 4936 15260
rect 4960 15258 5016 15260
rect 5040 15258 5096 15260
rect 5120 15258 5176 15260
rect 4880 15206 4926 15258
rect 4926 15206 4936 15258
rect 4960 15206 4990 15258
rect 4990 15206 5002 15258
rect 5002 15206 5016 15258
rect 5040 15206 5054 15258
rect 5054 15206 5066 15258
rect 5066 15206 5096 15258
rect 5120 15206 5130 15258
rect 5130 15206 5176 15258
rect 4880 15204 4936 15206
rect 4960 15204 5016 15206
rect 5040 15204 5096 15206
rect 5120 15204 5176 15206
rect 5814 15272 5870 15328
rect 4880 14170 4936 14172
rect 4960 14170 5016 14172
rect 5040 14170 5096 14172
rect 5120 14170 5176 14172
rect 4880 14118 4926 14170
rect 4926 14118 4936 14170
rect 4960 14118 4990 14170
rect 4990 14118 5002 14170
rect 5002 14118 5016 14170
rect 5040 14118 5054 14170
rect 5054 14118 5066 14170
rect 5066 14118 5096 14170
rect 5120 14118 5130 14170
rect 5130 14118 5176 14170
rect 4880 14116 4936 14118
rect 4960 14116 5016 14118
rect 5040 14116 5096 14118
rect 5120 14116 5176 14118
rect 4802 13912 4858 13968
rect 4158 12008 4214 12064
rect 4880 13082 4936 13084
rect 4960 13082 5016 13084
rect 5040 13082 5096 13084
rect 5120 13082 5176 13084
rect 4880 13030 4926 13082
rect 4926 13030 4936 13082
rect 4960 13030 4990 13082
rect 4990 13030 5002 13082
rect 5002 13030 5016 13082
rect 5040 13030 5054 13082
rect 5054 13030 5066 13082
rect 5066 13030 5096 13082
rect 5120 13030 5130 13082
rect 5130 13030 5176 13082
rect 4880 13028 4936 13030
rect 4960 13028 5016 13030
rect 5040 13028 5096 13030
rect 5120 13028 5176 13030
rect 4894 12824 4950 12880
rect 4986 12416 5042 12472
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4526 11192 4582 11248
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4986 10668 5042 10704
rect 4986 10648 4988 10668
rect 4988 10648 5040 10668
rect 5040 10648 5042 10668
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 2962 6724 3018 6760
rect 2962 6704 2964 6724
rect 2964 6704 3016 6724
rect 3016 6704 3018 6724
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 5262 7792 5318 7848
rect 4066 7404 4122 7440
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 4066 7384 4068 7404
rect 4068 7384 4120 7404
rect 4120 7384 4122 7404
rect 5170 7384 5226 7440
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 5354 6724 5410 6760
rect 5354 6704 5356 6724
rect 5356 6704 5408 6724
rect 5408 6704 5410 6724
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 6366 14356 6368 14376
rect 6368 14356 6420 14376
rect 6420 14356 6422 14376
rect 6366 14320 6422 14356
rect 6734 14320 6790 14376
rect 6458 12416 6514 12472
rect 8114 29708 8170 29744
rect 8114 29688 8116 29708
rect 8116 29688 8168 29708
rect 8168 29688 8170 29708
rect 7654 25492 7710 25528
rect 7654 25472 7656 25492
rect 7656 25472 7708 25492
rect 7708 25472 7710 25492
rect 8114 25492 8170 25528
rect 8114 25472 8116 25492
rect 8116 25472 8168 25492
rect 8168 25472 8170 25492
rect 10506 30640 10562 30696
rect 10782 30368 10838 30424
rect 12806 32836 12862 32872
rect 15290 32852 15292 32872
rect 15292 32852 15344 32872
rect 15344 32852 15346 32872
rect 12806 32816 12808 32836
rect 12808 32816 12860 32836
rect 12860 32816 12862 32836
rect 11978 32136 12034 32192
rect 11702 31864 11758 31920
rect 11242 28600 11298 28656
rect 9494 23024 9550 23080
rect 10322 23296 10378 23352
rect 9678 22208 9734 22264
rect 9402 20712 9458 20768
rect 8850 15564 8906 15600
rect 8850 15544 8852 15564
rect 8852 15544 8904 15564
rect 8904 15544 8906 15564
rect 8758 15272 8814 15328
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 9310 16496 9366 16552
rect 9586 16108 9642 16144
rect 9586 16088 9588 16108
rect 9588 16088 9640 16108
rect 9640 16088 9642 16108
rect 9770 15444 9772 15464
rect 9772 15444 9824 15464
rect 9824 15444 9826 15464
rect 9770 15408 9826 15444
rect 10046 16088 10102 16144
rect 9954 15544 10010 15600
rect 9770 14320 9826 14376
rect 9126 12280 9182 12336
rect 9218 11500 9220 11520
rect 9220 11500 9272 11520
rect 9272 11500 9274 11520
rect 9218 11464 9274 11500
rect 9862 13368 9918 13424
rect 9862 12280 9918 12336
rect 11058 26560 11114 26616
rect 11610 29416 11666 29472
rect 12530 32680 12586 32736
rect 11794 26288 11850 26344
rect 10966 24928 11022 24984
rect 11242 23432 11298 23488
rect 11702 23432 11758 23488
rect 11978 24112 12034 24168
rect 11794 23296 11850 23352
rect 12162 24520 12218 24576
rect 12438 26288 12494 26344
rect 12806 26424 12862 26480
rect 12162 24112 12218 24168
rect 12254 23060 12256 23080
rect 12256 23060 12308 23080
rect 12308 23060 12310 23080
rect 12254 23024 12310 23060
rect 12162 22888 12218 22944
rect 12070 22752 12126 22808
rect 10598 15272 10654 15328
rect 11242 17856 11298 17912
rect 11058 15408 11114 15464
rect 7746 6024 7802 6080
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 8758 3984 8814 4040
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 11518 16632 11574 16688
rect 12530 22888 12586 22944
rect 13818 31864 13874 31920
rect 13634 31456 13690 31512
rect 14370 32272 14426 32328
rect 14278 31864 14334 31920
rect 14554 32272 14610 32328
rect 14554 31864 14610 31920
rect 15290 32816 15346 32852
rect 14094 30096 14150 30152
rect 12990 27648 13046 27704
rect 13450 26832 13506 26888
rect 12806 23568 12862 23624
rect 12438 22208 12494 22264
rect 12346 21140 12402 21176
rect 12346 21120 12348 21140
rect 12348 21120 12400 21140
rect 12400 21120 12402 21140
rect 12162 19372 12218 19408
rect 12162 19352 12164 19372
rect 12164 19352 12216 19372
rect 12216 19352 12218 19372
rect 12254 15544 12310 15600
rect 12990 21936 13046 21992
rect 13818 26324 13820 26344
rect 13820 26324 13872 26344
rect 13872 26324 13874 26344
rect 13818 26288 13874 26324
rect 13082 18400 13138 18456
rect 11794 15020 11850 15056
rect 11794 15000 11796 15020
rect 11796 15000 11848 15020
rect 11848 15000 11850 15020
rect 12530 15308 12532 15328
rect 12532 15308 12584 15328
rect 12584 15308 12586 15328
rect 12530 15272 12586 15308
rect 11610 14356 11612 14376
rect 11612 14356 11664 14376
rect 11664 14356 11666 14376
rect 11610 14320 11666 14356
rect 12254 12008 12310 12064
rect 10966 10920 11022 10976
rect 12070 9560 12126 9616
rect 11242 5752 11298 5808
rect 13266 16224 13322 16280
rect 12714 12144 12770 12200
rect 11978 5364 12034 5400
rect 11978 5344 11980 5364
rect 11980 5344 12032 5364
rect 12032 5344 12034 5364
rect 14922 32272 14978 32328
rect 15014 29008 15070 29064
rect 13910 25200 13966 25256
rect 13818 23296 13874 23352
rect 15382 30504 15438 30560
rect 15382 29960 15438 30016
rect 15842 32680 15898 32736
rect 15658 32136 15714 32192
rect 15566 32000 15622 32056
rect 16118 32136 16174 32192
rect 15382 27920 15438 27976
rect 14646 24384 14702 24440
rect 14462 23160 14518 23216
rect 13818 17584 13874 17640
rect 15106 24384 15162 24440
rect 15198 23840 15254 23896
rect 15934 30232 15990 30288
rect 15934 29164 15990 29200
rect 15934 29144 15936 29164
rect 15936 29144 15988 29164
rect 15988 29144 15990 29164
rect 16302 31340 16358 31376
rect 16302 31320 16304 31340
rect 16304 31320 16356 31340
rect 16356 31320 16358 31340
rect 16302 29280 16358 29336
rect 15566 25336 15622 25392
rect 15842 26324 15844 26344
rect 15844 26324 15896 26344
rect 15896 26324 15898 26344
rect 15842 26288 15898 26324
rect 15198 23160 15254 23216
rect 15290 22480 15346 22536
rect 14830 20596 14886 20632
rect 14830 20576 14832 20596
rect 14832 20576 14884 20596
rect 14884 20576 14886 20596
rect 14370 19352 14426 19408
rect 14186 19080 14242 19136
rect 14002 16532 14004 16552
rect 14004 16532 14056 16552
rect 14056 16532 14058 16552
rect 14002 16496 14058 16532
rect 15198 19760 15254 19816
rect 14830 17196 14886 17232
rect 14830 17176 14832 17196
rect 14832 17176 14884 17196
rect 14884 17176 14886 17196
rect 14646 17040 14702 17096
rect 14462 16496 14518 16552
rect 14094 15020 14150 15056
rect 14094 15000 14096 15020
rect 14096 15000 14148 15020
rect 14148 15000 14150 15020
rect 13726 13912 13782 13968
rect 13450 12144 13506 12200
rect 13634 11600 13690 11656
rect 13174 10104 13230 10160
rect 12898 9716 12954 9752
rect 12898 9696 12900 9716
rect 12900 9696 12952 9716
rect 12952 9696 12954 9716
rect 12806 7520 12862 7576
rect 13266 7792 13322 7848
rect 14002 12008 14058 12064
rect 15106 17176 15162 17232
rect 15382 18808 15438 18864
rect 16210 25880 16266 25936
rect 15658 19896 15714 19952
rect 15198 17060 15254 17096
rect 15198 17040 15200 17060
rect 15200 17040 15252 17060
rect 15252 17040 15254 17060
rect 14738 16532 14740 16552
rect 14740 16532 14792 16552
rect 14792 16532 14794 16552
rect 14738 16496 14794 16532
rect 15658 19352 15714 19408
rect 15842 21836 15844 21856
rect 15844 21836 15896 21856
rect 15896 21836 15898 21856
rect 15842 21800 15898 21836
rect 16026 20576 16082 20632
rect 16210 21120 16266 21176
rect 16302 20440 16358 20496
rect 16394 19896 16450 19952
rect 16302 18708 16304 18728
rect 16304 18708 16356 18728
rect 16356 18708 16358 18728
rect 16302 18672 16358 18708
rect 16302 17720 16358 17776
rect 15566 16768 15622 16824
rect 14646 15000 14702 15056
rect 15198 16360 15254 16416
rect 15106 16224 15162 16280
rect 15750 16632 15806 16688
rect 15750 16224 15806 16280
rect 15290 15680 15346 15736
rect 15290 15544 15346 15600
rect 15382 15136 15438 15192
rect 15382 13640 15438 13696
rect 14462 12008 14518 12064
rect 14370 11756 14426 11792
rect 14370 11736 14372 11756
rect 14372 11736 14424 11756
rect 14424 11736 14426 11756
rect 13358 6568 13414 6624
rect 13174 6296 13230 6352
rect 12806 5888 12862 5944
rect 12346 5516 12348 5536
rect 12348 5516 12400 5536
rect 12400 5516 12402 5536
rect 12346 5480 12402 5516
rect 12990 5344 13046 5400
rect 11610 4276 11666 4312
rect 11610 4256 11612 4276
rect 11612 4256 11664 4276
rect 11664 4256 11666 4276
rect 12898 5228 12954 5264
rect 12898 5208 12900 5228
rect 12900 5208 12952 5228
rect 12952 5208 12954 5228
rect 15014 12280 15070 12336
rect 15842 12552 15898 12608
rect 16302 15000 16358 15056
rect 15474 12180 15476 12200
rect 15476 12180 15528 12200
rect 15528 12180 15530 12200
rect 15474 12144 15530 12180
rect 15566 11736 15622 11792
rect 15198 10240 15254 10296
rect 14554 9444 14610 9480
rect 14554 9424 14556 9444
rect 14556 9424 14608 9444
rect 14608 9424 14610 9444
rect 14462 7828 14464 7848
rect 14464 7828 14516 7848
rect 14516 7828 14518 7848
rect 13818 5344 13874 5400
rect 14462 7792 14518 7828
rect 14462 6840 14518 6896
rect 15290 8880 15346 8936
rect 14738 6024 14794 6080
rect 14738 5636 14794 5672
rect 14738 5616 14740 5636
rect 14740 5616 14792 5636
rect 14792 5616 14794 5636
rect 15014 6314 15070 6352
rect 15014 6296 15016 6314
rect 15016 6296 15068 6314
rect 15068 6296 15070 6314
rect 14738 3984 14794 4040
rect 15198 6840 15254 6896
rect 15290 6568 15346 6624
rect 15382 6296 15438 6352
rect 15198 6180 15254 6216
rect 15198 6160 15200 6180
rect 15200 6160 15252 6180
rect 15252 6160 15254 6180
rect 15198 5344 15254 5400
rect 15198 4120 15254 4176
rect 14830 3440 14886 3496
rect 15750 10104 15806 10160
rect 16210 12960 16266 13016
rect 16210 10920 16266 10976
rect 15658 6452 15714 6488
rect 15658 6432 15660 6452
rect 15660 6432 15712 6452
rect 15712 6432 15714 6452
rect 16210 8200 16266 8256
rect 16210 5888 16266 5944
rect 15474 5752 15530 5808
rect 15658 5752 15714 5808
rect 15658 3984 15714 4040
rect 16210 4800 16266 4856
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
<< metal3 >>
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 12801 32874 12867 32877
rect 15285 32874 15351 32877
rect 12801 32872 15351 32874
rect 12801 32816 12806 32872
rect 12862 32816 15290 32872
rect 15346 32816 15351 32872
rect 12801 32814 15351 32816
rect 12801 32811 12867 32814
rect 15285 32811 15351 32814
rect 12525 32738 12591 32741
rect 15837 32738 15903 32741
rect 12525 32736 15903 32738
rect 12525 32680 12530 32736
rect 12586 32680 15842 32736
rect 15898 32680 15903 32736
rect 12525 32678 15903 32680
rect 12525 32675 12591 32678
rect 15837 32675 15903 32678
rect 4870 32672 5186 32673
rect 4870 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5186 32672
rect 4870 32607 5186 32608
rect 14365 32330 14431 32333
rect 14549 32330 14615 32333
rect 14917 32330 14983 32333
rect 14365 32328 14983 32330
rect 14365 32272 14370 32328
rect 14426 32272 14554 32328
rect 14610 32272 14922 32328
rect 14978 32272 14983 32328
rect 14365 32270 14983 32272
rect 14365 32267 14431 32270
rect 14549 32267 14615 32270
rect 14917 32267 14983 32270
rect 11973 32194 12039 32197
rect 15653 32194 15719 32197
rect 16113 32194 16179 32197
rect 11973 32192 16179 32194
rect 11973 32136 11978 32192
rect 12034 32136 15658 32192
rect 15714 32136 16118 32192
rect 16174 32136 16179 32192
rect 11973 32134 16179 32136
rect 11973 32131 12039 32134
rect 15653 32131 15719 32134
rect 16113 32131 16179 32134
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 15561 32058 15627 32061
rect 12390 32056 15627 32058
rect 12390 32000 15566 32056
rect 15622 32000 15627 32056
rect 12390 31998 15627 32000
rect 7005 31922 7071 31925
rect 8150 31922 8156 31924
rect 7005 31920 8156 31922
rect 7005 31864 7010 31920
rect 7066 31864 8156 31920
rect 7005 31862 8156 31864
rect 7005 31859 7071 31862
rect 8150 31860 8156 31862
rect 8220 31860 8226 31924
rect 11697 31922 11763 31925
rect 12390 31922 12450 31998
rect 15561 31995 15627 31998
rect 11697 31920 12450 31922
rect 11697 31864 11702 31920
rect 11758 31864 12450 31920
rect 11697 31862 12450 31864
rect 13813 31924 13879 31925
rect 13813 31920 13860 31924
rect 13924 31922 13930 31924
rect 14273 31922 14339 31925
rect 14549 31922 14615 31925
rect 13813 31864 13818 31920
rect 11697 31859 11763 31862
rect 13813 31860 13860 31864
rect 13924 31862 13970 31922
rect 14273 31920 14615 31922
rect 14273 31864 14278 31920
rect 14334 31864 14554 31920
rect 14610 31864 14615 31920
rect 14273 31862 14615 31864
rect 13924 31860 13930 31862
rect 13813 31859 13879 31860
rect 14273 31859 14339 31862
rect 14549 31859 14615 31862
rect 7189 31786 7255 31789
rect 7782 31786 7788 31788
rect 7189 31784 7788 31786
rect 7189 31728 7194 31784
rect 7250 31728 7788 31784
rect 7189 31726 7788 31728
rect 7189 31723 7255 31726
rect 7782 31724 7788 31726
rect 7852 31724 7858 31788
rect 4870 31584 5186 31585
rect 4870 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5186 31584
rect 4870 31519 5186 31520
rect 13486 31452 13492 31516
rect 13556 31514 13562 31516
rect 13629 31514 13695 31517
rect 13556 31512 13695 31514
rect 13556 31456 13634 31512
rect 13690 31456 13695 31512
rect 13556 31454 13695 31456
rect 13556 31452 13562 31454
rect 13629 31451 13695 31454
rect 0 31380 800 31408
rect 0 31316 796 31380
rect 860 31316 866 31380
rect 16297 31378 16363 31381
rect 16989 31378 17789 31408
rect 16297 31376 17789 31378
rect 16297 31320 16302 31376
rect 16358 31320 17789 31376
rect 16297 31318 17789 31320
rect 0 31288 800 31316
rect 16297 31315 16363 31318
rect 16989 31288 17789 31318
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 10501 30698 10567 30701
rect 16989 30698 17789 30728
rect 10501 30696 17789 30698
rect 10501 30640 10506 30696
rect 10562 30640 17789 30696
rect 10501 30638 17789 30640
rect 10501 30635 10567 30638
rect 16989 30608 17789 30638
rect 14222 30500 14228 30564
rect 14292 30562 14298 30564
rect 15377 30562 15443 30565
rect 14292 30560 15443 30562
rect 14292 30504 15382 30560
rect 15438 30504 15443 30560
rect 14292 30502 15443 30504
rect 14292 30500 14298 30502
rect 15377 30499 15443 30502
rect 4870 30496 5186 30497
rect 4870 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5186 30496
rect 4870 30431 5186 30432
rect 10777 30428 10843 30429
rect 10726 30426 10732 30428
rect 10686 30366 10732 30426
rect 10796 30426 10843 30428
rect 10796 30424 15210 30426
rect 10838 30368 15210 30424
rect 10726 30364 10732 30366
rect 10796 30366 15210 30368
rect 10796 30364 10843 30366
rect 10777 30363 10843 30364
rect 15150 30290 15210 30366
rect 15929 30290 15995 30293
rect 15150 30288 15995 30290
rect 15150 30232 15934 30288
rect 15990 30232 15995 30288
rect 15150 30230 15995 30232
rect 15929 30227 15995 30230
rect 105 30154 171 30157
rect 14089 30156 14155 30157
rect 790 30154 796 30156
rect 105 30152 796 30154
rect 105 30096 110 30152
rect 166 30096 796 30152
rect 105 30094 796 30096
rect 105 30091 171 30094
rect 790 30092 796 30094
rect 860 30092 866 30156
rect 14038 30092 14044 30156
rect 14108 30154 14155 30156
rect 14108 30152 14200 30154
rect 14150 30096 14200 30152
rect 14108 30094 14200 30096
rect 14108 30092 14155 30094
rect 14089 30091 14155 30092
rect 15377 30018 15443 30021
rect 16989 30018 17789 30048
rect 15377 30016 17789 30018
rect 15377 29960 15382 30016
rect 15438 29960 17789 30016
rect 15377 29958 17789 29960
rect 15377 29955 15443 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 16989 29928 17789 29958
rect 4210 29887 4526 29888
rect 6913 29746 6979 29749
rect 7281 29746 7347 29749
rect 8109 29746 8175 29749
rect 6913 29744 8175 29746
rect 6913 29688 6918 29744
rect 6974 29688 7286 29744
rect 7342 29688 8114 29744
rect 8170 29688 8175 29744
rect 6913 29686 8175 29688
rect 6913 29683 6979 29686
rect 7281 29683 7347 29686
rect 8109 29683 8175 29686
rect 11605 29474 11671 29477
rect 12014 29474 12020 29476
rect 11605 29472 12020 29474
rect 11605 29416 11610 29472
rect 11666 29416 12020 29472
rect 11605 29414 12020 29416
rect 11605 29411 11671 29414
rect 12014 29412 12020 29414
rect 12084 29412 12090 29476
rect 4870 29408 5186 29409
rect 4870 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5186 29408
rect 4870 29343 5186 29344
rect 16297 29338 16363 29341
rect 16989 29338 17789 29368
rect 16297 29336 17789 29338
rect 16297 29280 16302 29336
rect 16358 29280 17789 29336
rect 16297 29278 17789 29280
rect 16297 29275 16363 29278
rect 16989 29248 17789 29278
rect 9438 29140 9444 29204
rect 9508 29202 9514 29204
rect 15929 29202 15995 29205
rect 9508 29200 15995 29202
rect 9508 29144 15934 29200
rect 15990 29144 15995 29200
rect 9508 29142 15995 29144
rect 9508 29140 9514 29142
rect 15929 29139 15995 29142
rect 11830 29004 11836 29068
rect 11900 29066 11906 29068
rect 15009 29066 15075 29069
rect 11900 29064 15075 29066
rect 11900 29008 15014 29064
rect 15070 29008 15075 29064
rect 11900 29006 15075 29008
rect 11900 29004 11906 29006
rect 15009 29003 15075 29006
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 11237 28658 11303 28661
rect 16989 28658 17789 28688
rect 11237 28656 17789 28658
rect 11237 28600 11242 28656
rect 11298 28600 17789 28656
rect 11237 28598 17789 28600
rect 11237 28595 11303 28598
rect 16989 28568 17789 28598
rect 4870 28320 5186 28321
rect 4870 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5186 28320
rect 4870 28255 5186 28256
rect 15377 27978 15443 27981
rect 16989 27978 17789 28008
rect 15377 27976 17789 27978
rect 15377 27920 15382 27976
rect 15438 27920 17789 27976
rect 15377 27918 17789 27920
rect 15377 27915 15443 27918
rect 16989 27888 17789 27918
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 12566 27644 12572 27708
rect 12636 27706 12642 27708
rect 12985 27706 13051 27709
rect 12636 27704 13051 27706
rect 12636 27648 12990 27704
rect 13046 27648 13051 27704
rect 12636 27646 13051 27648
rect 12636 27644 12642 27646
rect 12985 27643 13051 27646
rect 13854 27236 13860 27300
rect 13924 27298 13930 27300
rect 16989 27298 17789 27328
rect 13924 27238 17789 27298
rect 13924 27236 13930 27238
rect 4870 27232 5186 27233
rect 4870 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5186 27232
rect 16989 27208 17789 27238
rect 4870 27167 5186 27168
rect 2773 27026 2839 27029
rect 4797 27026 4863 27029
rect 5901 27026 5967 27029
rect 2773 27024 5967 27026
rect 2773 26968 2778 27024
rect 2834 26968 4802 27024
rect 4858 26968 5906 27024
rect 5962 26968 5967 27024
rect 2773 26966 5967 26968
rect 2773 26963 2839 26966
rect 4797 26963 4863 26966
rect 5901 26963 5967 26966
rect 2865 26890 2931 26893
rect 5073 26890 5139 26893
rect 13445 26892 13511 26893
rect 13445 26890 13492 26892
rect 2865 26888 5139 26890
rect 2865 26832 2870 26888
rect 2926 26832 5078 26888
rect 5134 26832 5139 26888
rect 2865 26830 5139 26832
rect 13400 26888 13492 26890
rect 13400 26832 13450 26888
rect 13400 26830 13492 26832
rect 2865 26827 2931 26830
rect 5073 26827 5139 26830
rect 13445 26828 13492 26830
rect 13556 26828 13562 26892
rect 13445 26827 13511 26828
rect 3049 26754 3115 26757
rect 3509 26754 3575 26757
rect 3049 26752 3575 26754
rect 3049 26696 3054 26752
rect 3110 26696 3514 26752
rect 3570 26696 3575 26752
rect 3049 26694 3575 26696
rect 3049 26691 3115 26694
rect 3509 26691 3575 26694
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 11053 26618 11119 26621
rect 16989 26618 17789 26648
rect 11053 26616 17789 26618
rect 11053 26560 11058 26616
rect 11114 26560 17789 26616
rect 11053 26558 17789 26560
rect 11053 26555 11119 26558
rect 16989 26528 17789 26558
rect 2589 26482 2655 26485
rect 2773 26482 2839 26485
rect 2589 26480 2839 26482
rect 2589 26424 2594 26480
rect 2650 26424 2778 26480
rect 2834 26424 2839 26480
rect 2589 26422 2839 26424
rect 2589 26419 2655 26422
rect 2773 26419 2839 26422
rect 12801 26482 12867 26485
rect 14222 26482 14228 26484
rect 12801 26480 14228 26482
rect 12801 26424 12806 26480
rect 12862 26424 14228 26480
rect 12801 26422 14228 26424
rect 12801 26419 12867 26422
rect 14222 26420 14228 26422
rect 14292 26420 14298 26484
rect 11789 26346 11855 26349
rect 12433 26346 12499 26349
rect 13813 26346 13879 26349
rect 11789 26344 13879 26346
rect 11789 26288 11794 26344
rect 11850 26288 12438 26344
rect 12494 26288 13818 26344
rect 13874 26288 13879 26344
rect 11789 26286 13879 26288
rect 11789 26283 11855 26286
rect 12433 26283 12499 26286
rect 13813 26283 13879 26286
rect 14774 26284 14780 26348
rect 14844 26346 14850 26348
rect 15837 26346 15903 26349
rect 14844 26344 15903 26346
rect 14844 26288 15842 26344
rect 15898 26288 15903 26344
rect 14844 26286 15903 26288
rect 14844 26284 14850 26286
rect 15837 26283 15903 26286
rect 4870 26144 5186 26145
rect 4870 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5186 26144
rect 4870 26079 5186 26080
rect 16205 25938 16271 25941
rect 16989 25938 17789 25968
rect 16205 25936 17789 25938
rect 16205 25880 16210 25936
rect 16266 25880 17789 25936
rect 16205 25878 17789 25880
rect 16205 25875 16271 25878
rect 16989 25848 17789 25878
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 7649 25530 7715 25533
rect 8109 25532 8175 25533
rect 7782 25530 7788 25532
rect 7649 25528 7788 25530
rect 7649 25472 7654 25528
rect 7710 25472 7788 25528
rect 7649 25470 7788 25472
rect 7649 25467 7715 25470
rect 7782 25468 7788 25470
rect 7852 25468 7858 25532
rect 8109 25530 8156 25532
rect 8064 25528 8156 25530
rect 8064 25472 8114 25528
rect 8064 25470 8156 25472
rect 8109 25468 8156 25470
rect 8220 25468 8226 25532
rect 8109 25467 8175 25468
rect 841 25394 907 25397
rect 798 25392 907 25394
rect 798 25336 846 25392
rect 902 25336 907 25392
rect 798 25331 907 25336
rect 14590 25332 14596 25396
rect 14660 25394 14666 25396
rect 15561 25394 15627 25397
rect 14660 25392 15627 25394
rect 14660 25336 15566 25392
rect 15622 25336 15627 25392
rect 14660 25334 15627 25336
rect 14660 25332 14666 25334
rect 15561 25331 15627 25334
rect 798 25288 858 25331
rect 0 25198 858 25288
rect 13905 25258 13971 25261
rect 16989 25258 17789 25288
rect 13905 25256 17789 25258
rect 13905 25200 13910 25256
rect 13966 25200 17789 25256
rect 13905 25198 17789 25200
rect 0 25168 800 25198
rect 13905 25195 13971 25198
rect 16989 25168 17789 25198
rect 4870 25056 5186 25057
rect 4870 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5186 25056
rect 4870 24991 5186 24992
rect 10961 24988 11027 24989
rect 10910 24986 10916 24988
rect 10870 24926 10916 24986
rect 10980 24984 11027 24988
rect 11022 24928 11027 24984
rect 10910 24924 10916 24926
rect 10980 24924 11027 24928
rect 12198 24924 12204 24988
rect 12268 24986 12274 24988
rect 14038 24986 14044 24988
rect 12268 24926 14044 24986
rect 12268 24924 12274 24926
rect 14038 24924 14044 24926
rect 14108 24924 14114 24988
rect 10961 24923 11027 24924
rect 12157 24578 12223 24581
rect 16989 24578 17789 24608
rect 12157 24576 17789 24578
rect 12157 24520 12162 24576
rect 12218 24520 17789 24576
rect 12157 24518 17789 24520
rect 12157 24515 12223 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 16989 24488 17789 24518
rect 4210 24447 4526 24448
rect 14641 24442 14707 24445
rect 15101 24442 15167 24445
rect 14641 24440 15167 24442
rect 14641 24384 14646 24440
rect 14702 24384 15106 24440
rect 15162 24384 15167 24440
rect 14641 24382 15167 24384
rect 14641 24379 14707 24382
rect 15101 24379 15167 24382
rect 3969 24308 4035 24309
rect 3918 24306 3924 24308
rect 3878 24246 3924 24306
rect 3988 24304 4035 24308
rect 4030 24248 4035 24304
rect 3918 24244 3924 24246
rect 3988 24244 4035 24248
rect 3969 24243 4035 24244
rect 3182 24108 3188 24172
rect 3252 24170 3258 24172
rect 3417 24170 3483 24173
rect 3252 24168 3483 24170
rect 3252 24112 3422 24168
rect 3478 24112 3483 24168
rect 3252 24110 3483 24112
rect 3252 24108 3258 24110
rect 3417 24107 3483 24110
rect 11973 24170 12039 24173
rect 12157 24170 12223 24173
rect 11973 24168 12223 24170
rect 11973 24112 11978 24168
rect 12034 24112 12162 24168
rect 12218 24112 12223 24168
rect 11973 24110 12223 24112
rect 11973 24107 12039 24110
rect 12157 24107 12223 24110
rect 4870 23968 5186 23969
rect 4870 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5186 23968
rect 4870 23903 5186 23904
rect 15193 23898 15259 23901
rect 16989 23898 17789 23928
rect 15193 23896 17789 23898
rect 15193 23840 15198 23896
rect 15254 23840 17789 23896
rect 15193 23838 17789 23840
rect 15193 23835 15259 23838
rect 16989 23808 17789 23838
rect 12801 23626 12867 23629
rect 12934 23626 12940 23628
rect 12801 23624 12940 23626
rect 12801 23568 12806 23624
rect 12862 23568 12940 23624
rect 12801 23566 12940 23568
rect 12801 23563 12867 23566
rect 12934 23564 12940 23566
rect 13004 23564 13010 23628
rect 11237 23490 11303 23493
rect 11697 23490 11763 23493
rect 11237 23488 11763 23490
rect 11237 23432 11242 23488
rect 11298 23432 11702 23488
rect 11758 23432 11763 23488
rect 11237 23430 11763 23432
rect 11237 23427 11303 23430
rect 11697 23427 11763 23430
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 10317 23354 10383 23357
rect 11789 23354 11855 23357
rect 13813 23354 13879 23357
rect 10317 23352 13879 23354
rect 10317 23296 10322 23352
rect 10378 23296 11794 23352
rect 11850 23296 13818 23352
rect 13874 23296 13879 23352
rect 10317 23294 13879 23296
rect 10317 23291 10383 23294
rect 11789 23291 11855 23294
rect 13813 23291 13879 23294
rect 14457 23218 14523 23221
rect 14774 23218 14780 23220
rect 14457 23216 14780 23218
rect 14457 23160 14462 23216
rect 14518 23160 14780 23216
rect 14457 23158 14780 23160
rect 14457 23155 14523 23158
rect 14774 23156 14780 23158
rect 14844 23156 14850 23220
rect 15193 23218 15259 23221
rect 16989 23218 17789 23248
rect 15193 23216 17789 23218
rect 15193 23160 15198 23216
rect 15254 23160 17789 23216
rect 15193 23158 17789 23160
rect 15193 23155 15259 23158
rect 16989 23128 17789 23158
rect 9070 23020 9076 23084
rect 9140 23082 9146 23084
rect 9489 23082 9555 23085
rect 9140 23080 9555 23082
rect 9140 23024 9494 23080
rect 9550 23024 9555 23080
rect 9140 23022 9555 23024
rect 9140 23020 9146 23022
rect 9489 23019 9555 23022
rect 11646 23020 11652 23084
rect 11716 23082 11722 23084
rect 12249 23082 12315 23085
rect 11716 23080 12315 23082
rect 11716 23024 12254 23080
rect 12310 23024 12315 23080
rect 11716 23022 12315 23024
rect 11716 23020 11722 23022
rect 12249 23019 12315 23022
rect 12157 22946 12223 22949
rect 12525 22946 12591 22949
rect 12157 22944 12591 22946
rect 12157 22888 12162 22944
rect 12218 22888 12530 22944
rect 12586 22888 12591 22944
rect 12157 22886 12591 22888
rect 12157 22883 12223 22886
rect 12525 22883 12591 22886
rect 4870 22880 5186 22881
rect 4870 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5186 22880
rect 4870 22815 5186 22816
rect 11462 22748 11468 22812
rect 11532 22810 11538 22812
rect 12065 22810 12131 22813
rect 11532 22808 12131 22810
rect 11532 22752 12070 22808
rect 12126 22752 12131 22808
rect 11532 22750 12131 22752
rect 11532 22748 11538 22750
rect 12065 22747 12131 22750
rect 15285 22538 15351 22541
rect 16989 22538 17789 22568
rect 15285 22536 17789 22538
rect 15285 22480 15290 22536
rect 15346 22480 17789 22536
rect 15285 22478 17789 22480
rect 15285 22475 15351 22478
rect 16989 22448 17789 22478
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 9673 22266 9739 22269
rect 12433 22266 12499 22269
rect 9673 22264 12499 22266
rect 9673 22208 9678 22264
rect 9734 22208 12438 22264
rect 12494 22208 12499 22264
rect 9673 22206 12499 22208
rect 9673 22203 9739 22206
rect 12433 22203 12499 22206
rect 11830 22068 11836 22132
rect 11900 22130 11906 22132
rect 14774 22130 14780 22132
rect 11900 22070 14780 22130
rect 11900 22068 11906 22070
rect 14774 22068 14780 22070
rect 14844 22068 14850 22132
rect 12985 21994 13051 21997
rect 13118 21994 13124 21996
rect 12985 21992 13124 21994
rect 12985 21936 12990 21992
rect 13046 21936 13124 21992
rect 12985 21934 13124 21936
rect 12985 21931 13051 21934
rect 13118 21932 13124 21934
rect 13188 21932 13194 21996
rect 15837 21858 15903 21861
rect 16989 21858 17789 21888
rect 15837 21856 17789 21858
rect 15837 21800 15842 21856
rect 15898 21800 17789 21856
rect 15837 21798 17789 21800
rect 15837 21795 15903 21798
rect 4870 21792 5186 21793
rect 4870 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5186 21792
rect 16989 21768 17789 21798
rect 4870 21727 5186 21728
rect 12014 21388 12020 21452
rect 12084 21450 12090 21452
rect 13486 21450 13492 21452
rect 12084 21390 13492 21450
rect 12084 21388 12090 21390
rect 13486 21388 13492 21390
rect 13556 21388 13562 21452
rect 841 21314 907 21317
rect 798 21312 907 21314
rect 798 21256 846 21312
rect 902 21256 907 21312
rect 798 21251 907 21256
rect 798 21208 858 21251
rect 0 21118 858 21208
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 12341 21178 12407 21181
rect 12566 21178 12572 21180
rect 12341 21176 12572 21178
rect 12341 21120 12346 21176
rect 12402 21120 12572 21176
rect 12341 21118 12572 21120
rect 0 21088 800 21118
rect 12341 21115 12407 21118
rect 12566 21116 12572 21118
rect 12636 21116 12642 21180
rect 16205 21178 16271 21181
rect 16989 21178 17789 21208
rect 16205 21176 17789 21178
rect 16205 21120 16210 21176
rect 16266 21120 17789 21176
rect 16205 21118 17789 21120
rect 16205 21115 16271 21118
rect 16989 21088 17789 21118
rect 2221 20906 2287 20909
rect 2865 20906 2931 20909
rect 2221 20904 2931 20906
rect 2221 20848 2226 20904
rect 2282 20848 2870 20904
rect 2926 20848 2931 20904
rect 2221 20846 2931 20848
rect 2221 20843 2287 20846
rect 2865 20843 2931 20846
rect 9254 20708 9260 20772
rect 9324 20770 9330 20772
rect 9397 20770 9463 20773
rect 9324 20768 9463 20770
rect 9324 20712 9402 20768
rect 9458 20712 9463 20768
rect 9324 20710 9463 20712
rect 9324 20708 9330 20710
rect 9397 20707 9463 20710
rect 4870 20704 5186 20705
rect 4870 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5186 20704
rect 4870 20639 5186 20640
rect 3918 20572 3924 20636
rect 3988 20634 3994 20636
rect 4153 20634 4219 20637
rect 3988 20632 4219 20634
rect 3988 20576 4158 20632
rect 4214 20576 4219 20632
rect 3988 20574 4219 20576
rect 3988 20572 3994 20574
rect 4153 20571 4219 20574
rect 14825 20634 14891 20637
rect 16021 20634 16087 20637
rect 14825 20632 16087 20634
rect 14825 20576 14830 20632
rect 14886 20576 16026 20632
rect 16082 20576 16087 20632
rect 14825 20574 16087 20576
rect 14825 20571 14891 20574
rect 16021 20571 16087 20574
rect 16297 20498 16363 20501
rect 16989 20498 17789 20528
rect 16297 20496 17789 20498
rect 16297 20440 16302 20496
rect 16358 20440 17789 20496
rect 16297 20438 17789 20440
rect 16297 20435 16363 20438
rect 16989 20408 17789 20438
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 15653 19954 15719 19957
rect 16389 19954 16455 19957
rect 15653 19952 16455 19954
rect 15653 19896 15658 19952
rect 15714 19896 16394 19952
rect 16450 19896 16455 19952
rect 15653 19894 16455 19896
rect 15653 19891 15719 19894
rect 16389 19891 16455 19894
rect 5165 19818 5231 19821
rect 5349 19818 5415 19821
rect 5165 19816 5415 19818
rect 5165 19760 5170 19816
rect 5226 19760 5354 19816
rect 5410 19760 5415 19816
rect 5165 19758 5415 19760
rect 5165 19755 5231 19758
rect 5349 19755 5415 19758
rect 15193 19818 15259 19821
rect 16989 19818 17789 19848
rect 15193 19816 17789 19818
rect 15193 19760 15198 19816
rect 15254 19760 17789 19816
rect 15193 19758 17789 19760
rect 15193 19755 15259 19758
rect 16989 19728 17789 19758
rect 4870 19616 5186 19617
rect 4870 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5186 19616
rect 4870 19551 5186 19552
rect 5165 19410 5231 19413
rect 5993 19410 6059 19413
rect 12157 19412 12223 19413
rect 12157 19410 12204 19412
rect 5165 19408 6059 19410
rect 5165 19352 5170 19408
rect 5226 19352 5998 19408
rect 6054 19352 6059 19408
rect 5165 19350 6059 19352
rect 12112 19408 12204 19410
rect 12112 19352 12162 19408
rect 12112 19350 12204 19352
rect 5165 19347 5231 19350
rect 5993 19347 6059 19350
rect 12157 19348 12204 19350
rect 12268 19348 12274 19412
rect 14365 19410 14431 19413
rect 15653 19410 15719 19413
rect 14365 19408 15719 19410
rect 14365 19352 14370 19408
rect 14426 19352 15658 19408
rect 15714 19352 15719 19408
rect 14365 19350 15719 19352
rect 12157 19347 12223 19348
rect 14365 19347 14431 19350
rect 15653 19347 15719 19350
rect 3918 19212 3924 19276
rect 3988 19274 3994 19276
rect 4245 19274 4311 19277
rect 3988 19272 4311 19274
rect 3988 19216 4250 19272
rect 4306 19216 4311 19272
rect 3988 19214 4311 19216
rect 3988 19212 3994 19214
rect 4245 19211 4311 19214
rect 14181 19138 14247 19141
rect 16989 19138 17789 19168
rect 14181 19136 17789 19138
rect 14181 19080 14186 19136
rect 14242 19080 17789 19136
rect 14181 19078 17789 19080
rect 14181 19075 14247 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 16989 19048 17789 19078
rect 4210 19007 4526 19008
rect 15377 18868 15443 18869
rect 15326 18866 15332 18868
rect 15286 18806 15332 18866
rect 15396 18864 15443 18868
rect 15438 18808 15443 18864
rect 15326 18804 15332 18806
rect 15396 18804 15443 18808
rect 15377 18803 15443 18804
rect 13670 18668 13676 18732
rect 13740 18730 13746 18732
rect 16297 18730 16363 18733
rect 13740 18728 16363 18730
rect 13740 18672 16302 18728
rect 16358 18672 16363 18728
rect 13740 18670 16363 18672
rect 13740 18668 13746 18670
rect 16297 18667 16363 18670
rect 4870 18528 5186 18529
rect 4870 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5186 18528
rect 4870 18463 5186 18464
rect 13077 18458 13143 18461
rect 16989 18458 17789 18488
rect 13077 18456 17789 18458
rect 13077 18400 13082 18456
rect 13138 18400 17789 18456
rect 13077 18398 17789 18400
rect 13077 18395 13143 18398
rect 16989 18368 17789 18398
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 11237 17914 11303 17917
rect 13118 17914 13124 17916
rect 11237 17912 13124 17914
rect 11237 17856 11242 17912
rect 11298 17856 13124 17912
rect 11237 17854 13124 17856
rect 11237 17851 11303 17854
rect 13118 17852 13124 17854
rect 13188 17852 13194 17916
rect 10726 17716 10732 17780
rect 10796 17778 10802 17780
rect 16297 17778 16363 17781
rect 16989 17778 17789 17808
rect 10796 17776 16363 17778
rect 10796 17720 16302 17776
rect 16358 17720 16363 17776
rect 10796 17718 16363 17720
rect 10796 17716 10802 17718
rect 16297 17715 16363 17718
rect 16438 17718 17789 17778
rect 2405 17642 2471 17645
rect 3877 17642 3943 17645
rect 2405 17640 3943 17642
rect 2405 17584 2410 17640
rect 2466 17584 3882 17640
rect 3938 17584 3943 17640
rect 2405 17582 3943 17584
rect 2405 17579 2471 17582
rect 3877 17579 3943 17582
rect 13813 17642 13879 17645
rect 16438 17642 16498 17718
rect 16989 17688 17789 17718
rect 13813 17640 16498 17642
rect 13813 17584 13818 17640
rect 13874 17584 16498 17640
rect 13813 17582 16498 17584
rect 13813 17579 13879 17582
rect 4870 17440 5186 17441
rect 4870 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5186 17440
rect 4870 17375 5186 17376
rect 3141 17236 3207 17237
rect 3141 17234 3188 17236
rect 3096 17232 3188 17234
rect 3096 17176 3146 17232
rect 3096 17174 3188 17176
rect 3141 17172 3188 17174
rect 3252 17172 3258 17236
rect 14825 17234 14891 17237
rect 15101 17234 15167 17237
rect 14782 17232 15167 17234
rect 14782 17176 14830 17232
rect 14886 17176 15106 17232
rect 15162 17176 15167 17232
rect 14782 17174 15167 17176
rect 3141 17171 3207 17172
rect 14782 17171 14891 17174
rect 15101 17171 15167 17174
rect 14641 17098 14707 17101
rect 14782 17098 14842 17171
rect 14641 17096 14842 17098
rect 14641 17040 14646 17096
rect 14702 17040 14842 17096
rect 14641 17038 14842 17040
rect 15193 17098 15259 17101
rect 16989 17098 17789 17128
rect 15193 17096 17789 17098
rect 15193 17040 15198 17096
rect 15254 17040 17789 17096
rect 15193 17038 17789 17040
rect 14641 17035 14707 17038
rect 15193 17035 15259 17038
rect 16989 17008 17789 17038
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 14222 16764 14228 16828
rect 14292 16826 14298 16828
rect 15561 16826 15627 16829
rect 14292 16824 15627 16826
rect 14292 16768 15566 16824
rect 15622 16768 15627 16824
rect 14292 16766 15627 16768
rect 14292 16764 14298 16766
rect 15561 16763 15627 16766
rect 10910 16628 10916 16692
rect 10980 16690 10986 16692
rect 11513 16690 11579 16693
rect 10980 16688 11579 16690
rect 10980 16632 11518 16688
rect 11574 16632 11579 16688
rect 10980 16630 11579 16632
rect 10980 16628 10986 16630
rect 11513 16627 11579 16630
rect 14958 16628 14964 16692
rect 15028 16690 15034 16692
rect 15745 16690 15811 16693
rect 15028 16688 15811 16690
rect 15028 16632 15750 16688
rect 15806 16632 15811 16688
rect 15028 16630 15811 16632
rect 15028 16628 15034 16630
rect 15745 16627 15811 16630
rect 9305 16556 9371 16557
rect 9254 16554 9260 16556
rect 9214 16494 9260 16554
rect 9324 16552 9371 16556
rect 9366 16496 9371 16552
rect 9254 16492 9260 16494
rect 9324 16492 9371 16496
rect 9305 16491 9371 16492
rect 13997 16554 14063 16557
rect 14457 16554 14523 16557
rect 14733 16554 14799 16557
rect 13997 16552 14799 16554
rect 13997 16496 14002 16552
rect 14058 16496 14462 16552
rect 14518 16496 14738 16552
rect 14794 16496 14799 16552
rect 13997 16494 14799 16496
rect 13997 16491 14063 16494
rect 14457 16491 14523 16494
rect 14733 16491 14799 16494
rect 15193 16418 15259 16421
rect 16989 16418 17789 16448
rect 15193 16416 17789 16418
rect 15193 16360 15198 16416
rect 15254 16360 17789 16416
rect 15193 16358 17789 16360
rect 15193 16355 15259 16358
rect 4870 16352 5186 16353
rect 4870 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5186 16352
rect 16989 16328 17789 16358
rect 4870 16287 5186 16288
rect 13261 16282 13327 16285
rect 15101 16282 15167 16285
rect 15745 16282 15811 16285
rect 13261 16280 15811 16282
rect 13261 16224 13266 16280
rect 13322 16224 15106 16280
rect 15162 16224 15750 16280
rect 15806 16224 15811 16280
rect 13261 16222 15811 16224
rect 13261 16219 13327 16222
rect 15101 16219 15167 16222
rect 15745 16219 15811 16222
rect 9581 16146 9647 16149
rect 10041 16146 10107 16149
rect 9581 16144 10107 16146
rect 9581 16088 9586 16144
rect 9642 16088 10046 16144
rect 10102 16088 10107 16144
rect 9581 16086 10107 16088
rect 9581 16083 9647 16086
rect 9998 16083 10107 16086
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 2865 15738 2931 15741
rect 3182 15738 3188 15740
rect 2865 15736 3188 15738
rect 2865 15680 2870 15736
rect 2926 15680 3188 15736
rect 2865 15678 3188 15680
rect 2865 15675 2931 15678
rect 3182 15676 3188 15678
rect 3252 15676 3258 15740
rect 9998 15605 10058 16083
rect 15285 15738 15351 15741
rect 16989 15738 17789 15768
rect 15285 15736 17789 15738
rect 15285 15680 15290 15736
rect 15346 15680 17789 15736
rect 15285 15678 17789 15680
rect 15285 15675 15351 15678
rect 16989 15648 17789 15678
rect 2681 15602 2747 15605
rect 3233 15602 3299 15605
rect 5165 15602 5231 15605
rect 2681 15600 5231 15602
rect 2681 15544 2686 15600
rect 2742 15544 3238 15600
rect 3294 15544 5170 15600
rect 5226 15544 5231 15600
rect 2681 15542 5231 15544
rect 2681 15539 2747 15542
rect 3233 15539 3299 15542
rect 5165 15539 5231 15542
rect 8845 15602 8911 15605
rect 9949 15602 10058 15605
rect 8845 15600 10058 15602
rect 8845 15544 8850 15600
rect 8906 15544 9954 15600
rect 10010 15544 10058 15600
rect 8845 15542 10058 15544
rect 12249 15602 12315 15605
rect 15285 15604 15351 15605
rect 15285 15602 15332 15604
rect 12249 15600 15332 15602
rect 12249 15544 12254 15600
rect 12310 15544 15290 15600
rect 12249 15542 15332 15544
rect 8845 15539 8911 15542
rect 9949 15539 10015 15542
rect 12249 15539 12315 15542
rect 15285 15540 15332 15542
rect 15396 15540 15402 15604
rect 15285 15539 15351 15540
rect 3141 15466 3207 15469
rect 4061 15466 4127 15469
rect 3141 15464 4127 15466
rect 3141 15408 3146 15464
rect 3202 15408 4066 15464
rect 4122 15408 4127 15464
rect 3141 15406 4127 15408
rect 3141 15403 3207 15406
rect 4061 15403 4127 15406
rect 4654 15404 4660 15468
rect 4724 15466 4730 15468
rect 4889 15466 4955 15469
rect 4724 15464 4955 15466
rect 4724 15408 4894 15464
rect 4950 15408 4955 15464
rect 4724 15406 4955 15408
rect 4724 15404 4730 15406
rect 4889 15403 4955 15406
rect 5073 15466 5139 15469
rect 9765 15466 9831 15469
rect 11053 15466 11119 15469
rect 5073 15464 5826 15466
rect 5073 15408 5078 15464
rect 5134 15408 5826 15464
rect 5073 15406 5826 15408
rect 5073 15403 5139 15406
rect 5766 15333 5826 15406
rect 9765 15464 11119 15466
rect 9765 15408 9770 15464
rect 9826 15408 11058 15464
rect 11114 15408 11119 15464
rect 9765 15406 11119 15408
rect 9765 15403 9831 15406
rect 11053 15403 11119 15406
rect 5766 15332 5875 15333
rect 5758 15268 5764 15332
rect 5828 15330 5875 15332
rect 8753 15330 8819 15333
rect 10593 15330 10659 15333
rect 5828 15328 5920 15330
rect 5870 15272 5920 15328
rect 5828 15270 5920 15272
rect 8753 15328 10659 15330
rect 8753 15272 8758 15328
rect 8814 15272 10598 15328
rect 10654 15272 10659 15328
rect 8753 15270 10659 15272
rect 5828 15268 5875 15270
rect 5809 15267 5875 15268
rect 8753 15267 8819 15270
rect 10593 15267 10659 15270
rect 12525 15330 12591 15333
rect 12750 15330 12756 15332
rect 12525 15328 12756 15330
rect 12525 15272 12530 15328
rect 12586 15272 12756 15328
rect 12525 15270 12756 15272
rect 12525 15267 12591 15270
rect 12750 15268 12756 15270
rect 12820 15268 12826 15332
rect 4870 15264 5186 15265
rect 4870 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5186 15264
rect 4870 15199 5186 15200
rect 12198 15132 12204 15196
rect 12268 15194 12274 15196
rect 15377 15194 15443 15197
rect 12268 15192 15443 15194
rect 12268 15136 15382 15192
rect 15438 15136 15443 15192
rect 12268 15134 15443 15136
rect 12268 15132 12274 15134
rect 15377 15131 15443 15134
rect 11789 15058 11855 15061
rect 12014 15058 12020 15060
rect 11789 15056 12020 15058
rect 11789 15000 11794 15056
rect 11850 15000 12020 15056
rect 11789 14998 12020 15000
rect 11789 14995 11855 14998
rect 12014 14996 12020 14998
rect 12084 14996 12090 15060
rect 14089 15058 14155 15061
rect 14222 15058 14228 15060
rect 14089 15056 14228 15058
rect 14089 15000 14094 15056
rect 14150 15000 14228 15056
rect 14089 14998 14228 15000
rect 14089 14995 14155 14998
rect 14222 14996 14228 14998
rect 14292 15058 14298 15060
rect 14641 15058 14707 15061
rect 14292 15056 14707 15058
rect 14292 15000 14646 15056
rect 14702 15000 14707 15056
rect 14292 14998 14707 15000
rect 14292 14996 14298 14998
rect 14641 14995 14707 14998
rect 16297 15058 16363 15061
rect 16989 15058 17789 15088
rect 16297 15056 17789 15058
rect 16297 15000 16302 15056
rect 16358 15000 17789 15056
rect 16297 14998 17789 15000
rect 16297 14995 16363 14998
rect 16989 14968 17789 14998
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 3366 14316 3372 14380
rect 3436 14378 3442 14380
rect 6361 14378 6427 14381
rect 6729 14378 6795 14381
rect 3436 14376 6795 14378
rect 3436 14320 6366 14376
rect 6422 14320 6734 14376
rect 6790 14320 6795 14376
rect 3436 14318 6795 14320
rect 3436 14316 3442 14318
rect 6361 14315 6427 14318
rect 6729 14315 6795 14318
rect 9765 14378 9831 14381
rect 11605 14378 11671 14381
rect 16989 14378 17789 14408
rect 9765 14376 11671 14378
rect 9765 14320 9770 14376
rect 9826 14320 11610 14376
rect 11666 14320 11671 14376
rect 9765 14318 11671 14320
rect 9765 14315 9831 14318
rect 11605 14315 11671 14318
rect 13908 14318 17789 14378
rect 4870 14176 5186 14177
rect 4870 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5186 14176
rect 4870 14111 5186 14112
rect 3601 13970 3667 13973
rect 3734 13970 3740 13972
rect 3601 13968 3740 13970
rect 3601 13912 3606 13968
rect 3662 13912 3740 13968
rect 3601 13910 3740 13912
rect 3601 13907 3667 13910
rect 3734 13908 3740 13910
rect 3804 13970 3810 13972
rect 4797 13970 4863 13973
rect 3804 13968 4863 13970
rect 3804 13912 4802 13968
rect 4858 13912 4863 13968
rect 3804 13910 4863 13912
rect 3804 13908 3810 13910
rect 4797 13907 4863 13910
rect 13721 13970 13787 13973
rect 13908 13970 13968 14318
rect 16989 14288 17789 14318
rect 13721 13968 13968 13970
rect 13721 13912 13726 13968
rect 13782 13912 13968 13968
rect 13721 13910 13968 13912
rect 13721 13907 13787 13910
rect 3601 13698 3667 13701
rect 3918 13698 3924 13700
rect 3601 13696 3924 13698
rect 3601 13640 3606 13696
rect 3662 13640 3924 13696
rect 3601 13638 3924 13640
rect 3601 13635 3667 13638
rect 3918 13636 3924 13638
rect 3988 13636 3994 13700
rect 15377 13698 15443 13701
rect 16989 13698 17789 13728
rect 15377 13696 17789 13698
rect 15377 13640 15382 13696
rect 15438 13640 17789 13696
rect 15377 13638 17789 13640
rect 15377 13635 15443 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 16989 13608 17789 13638
rect 4210 13567 4526 13568
rect 3417 13424 3483 13429
rect 3417 13368 3422 13424
rect 3478 13368 3483 13424
rect 3417 13363 3483 13368
rect 3877 13426 3943 13429
rect 4245 13426 4311 13429
rect 3877 13424 4311 13426
rect 3877 13368 3882 13424
rect 3938 13368 4250 13424
rect 4306 13368 4311 13424
rect 3877 13366 4311 13368
rect 3877 13363 3943 13366
rect 4245 13363 4311 13366
rect 9857 13426 9923 13429
rect 11646 13426 11652 13428
rect 9857 13424 11652 13426
rect 9857 13368 9862 13424
rect 9918 13368 11652 13424
rect 9857 13366 11652 13368
rect 9857 13363 9923 13366
rect 11646 13364 11652 13366
rect 11716 13364 11722 13428
rect 3420 13290 3480 13363
rect 4245 13290 4311 13293
rect 3420 13288 4311 13290
rect 3420 13232 4250 13288
rect 4306 13232 4311 13288
rect 3420 13230 4311 13232
rect 4245 13227 4311 13230
rect 4870 13088 5186 13089
rect 4870 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5186 13088
rect 4870 13023 5186 13024
rect 16205 13018 16271 13021
rect 16989 13018 17789 13048
rect 16205 13016 17789 13018
rect 16205 12960 16210 13016
rect 16266 12960 17789 13016
rect 16205 12958 17789 12960
rect 16205 12955 16271 12958
rect 16989 12928 17789 12958
rect 4889 12882 4955 12885
rect 5758 12882 5764 12884
rect 4889 12880 5764 12882
rect 4889 12824 4894 12880
rect 4950 12824 5764 12880
rect 4889 12822 5764 12824
rect 4889 12819 4955 12822
rect 5758 12820 5764 12822
rect 5828 12820 5834 12884
rect 14406 12548 14412 12612
rect 14476 12610 14482 12612
rect 15837 12610 15903 12613
rect 14476 12608 15903 12610
rect 14476 12552 15842 12608
rect 15898 12552 15903 12608
rect 14476 12550 15903 12552
rect 14476 12548 14482 12550
rect 15837 12547 15903 12550
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 4981 12474 5047 12477
rect 6453 12474 6519 12477
rect 4981 12472 6519 12474
rect 4981 12416 4986 12472
rect 5042 12416 6458 12472
rect 6514 12416 6519 12472
rect 4981 12414 6519 12416
rect 4981 12411 5047 12414
rect 6453 12411 6519 12414
rect 3417 12340 3483 12341
rect 9121 12340 9187 12341
rect 3366 12276 3372 12340
rect 3436 12338 3483 12340
rect 9070 12338 9076 12340
rect 3436 12336 3528 12338
rect 3478 12280 3528 12336
rect 3436 12278 3528 12280
rect 9030 12278 9076 12338
rect 9140 12338 9187 12340
rect 9857 12338 9923 12341
rect 9140 12336 9923 12338
rect 9182 12280 9862 12336
rect 9918 12280 9923 12336
rect 3436 12276 3483 12278
rect 9070 12276 9076 12278
rect 9140 12278 9923 12280
rect 9140 12276 9187 12278
rect 3417 12275 3483 12276
rect 9121 12275 9187 12276
rect 9857 12275 9923 12278
rect 15009 12338 15075 12341
rect 16989 12338 17789 12368
rect 15009 12336 17789 12338
rect 15009 12280 15014 12336
rect 15070 12280 17789 12336
rect 15009 12278 17789 12280
rect 15009 12275 15075 12278
rect 16989 12248 17789 12278
rect 12709 12202 12775 12205
rect 12390 12200 12775 12202
rect 12390 12144 12714 12200
rect 12770 12144 12775 12200
rect 12390 12142 12775 12144
rect 2865 12066 2931 12069
rect 4153 12066 4219 12069
rect 2865 12064 4219 12066
rect 2865 12008 2870 12064
rect 2926 12008 4158 12064
rect 4214 12008 4219 12064
rect 2865 12006 4219 12008
rect 2865 12003 2931 12006
rect 4153 12003 4219 12006
rect 12249 12066 12315 12069
rect 12390 12066 12450 12142
rect 12709 12139 12775 12142
rect 13445 12202 13511 12205
rect 15469 12202 15535 12205
rect 13445 12200 15535 12202
rect 13445 12144 13450 12200
rect 13506 12144 15474 12200
rect 15530 12144 15535 12200
rect 13445 12142 15535 12144
rect 13445 12139 13511 12142
rect 15469 12139 15535 12142
rect 12249 12064 12450 12066
rect 12249 12008 12254 12064
rect 12310 12008 12450 12064
rect 12249 12006 12450 12008
rect 13997 12066 14063 12069
rect 14457 12066 14523 12069
rect 13997 12064 14523 12066
rect 13997 12008 14002 12064
rect 14058 12008 14462 12064
rect 14518 12008 14523 12064
rect 13997 12006 14523 12008
rect 12249 12003 12315 12006
rect 13997 12003 14063 12006
rect 14457 12003 14523 12006
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 14365 11794 14431 11797
rect 15561 11794 15627 11797
rect 14365 11792 15627 11794
rect 14365 11736 14370 11792
rect 14426 11736 15566 11792
rect 15622 11736 15627 11792
rect 14365 11734 15627 11736
rect 14365 11731 14431 11734
rect 15561 11731 15627 11734
rect 13629 11658 13695 11661
rect 16989 11658 17789 11688
rect 13629 11656 17789 11658
rect 13629 11600 13634 11656
rect 13690 11600 17789 11656
rect 13629 11598 17789 11600
rect 13629 11595 13695 11598
rect 16989 11568 17789 11598
rect 9070 11460 9076 11524
rect 9140 11522 9146 11524
rect 9213 11522 9279 11525
rect 9140 11520 9279 11522
rect 9140 11464 9218 11520
rect 9274 11464 9279 11520
rect 9140 11462 9279 11464
rect 9140 11460 9146 11462
rect 9213 11459 9279 11462
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 3734 11188 3740 11252
rect 3804 11250 3810 11252
rect 4521 11250 4587 11253
rect 3804 11248 4587 11250
rect 3804 11192 4526 11248
rect 4582 11192 4587 11248
rect 3804 11190 4587 11192
rect 3804 11188 3810 11190
rect 4521 11187 4587 11190
rect 10961 10978 11027 10981
rect 12566 10978 12572 10980
rect 10961 10976 12572 10978
rect 10961 10920 10966 10976
rect 11022 10920 12572 10976
rect 10961 10918 12572 10920
rect 10961 10915 11027 10918
rect 12566 10916 12572 10918
rect 12636 10916 12642 10980
rect 16205 10978 16271 10981
rect 16989 10978 17789 11008
rect 16205 10976 17789 10978
rect 16205 10920 16210 10976
rect 16266 10920 17789 10976
rect 16205 10918 17789 10920
rect 16205 10915 16271 10918
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 16989 10888 17789 10918
rect 4870 10847 5186 10848
rect 4654 10644 4660 10708
rect 4724 10706 4730 10708
rect 4981 10706 5047 10709
rect 4724 10704 5047 10706
rect 4724 10648 4986 10704
rect 5042 10648 5047 10704
rect 4724 10646 5047 10648
rect 4724 10644 4730 10646
rect 4981 10643 5047 10646
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 15193 10298 15259 10301
rect 16989 10298 17789 10328
rect 15193 10296 17789 10298
rect 15193 10240 15198 10296
rect 15254 10240 17789 10296
rect 15193 10238 17789 10240
rect 15193 10235 15259 10238
rect 16989 10208 17789 10238
rect 13169 10162 13235 10165
rect 13670 10162 13676 10164
rect 13169 10160 13676 10162
rect 13169 10104 13174 10160
rect 13230 10104 13676 10160
rect 13169 10102 13676 10104
rect 13169 10099 13235 10102
rect 13670 10100 13676 10102
rect 13740 10162 13746 10164
rect 15745 10162 15811 10165
rect 13740 10160 15811 10162
rect 13740 10104 15750 10160
rect 15806 10104 15811 10160
rect 13740 10102 15811 10104
rect 13740 10100 13746 10102
rect 15745 10099 15811 10102
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 12893 9756 12959 9757
rect 12893 9754 12940 9756
rect 12848 9752 12940 9754
rect 12848 9696 12898 9752
rect 12848 9694 12940 9696
rect 12893 9692 12940 9694
rect 13004 9692 13010 9756
rect 12893 9691 12959 9692
rect 12065 9618 12131 9621
rect 16989 9618 17789 9648
rect 12065 9616 17789 9618
rect 12065 9560 12070 9616
rect 12126 9560 17789 9616
rect 12065 9558 17789 9560
rect 12065 9555 12131 9558
rect 16989 9528 17789 9558
rect 13486 9420 13492 9484
rect 13556 9482 13562 9484
rect 14549 9482 14615 9485
rect 13556 9480 14615 9482
rect 13556 9424 14554 9480
rect 14610 9424 14615 9480
rect 13556 9422 14615 9424
rect 13556 9420 13562 9422
rect 14549 9419 14615 9422
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 15285 8938 15351 8941
rect 16989 8938 17789 8968
rect 15285 8936 17789 8938
rect 15285 8880 15290 8936
rect 15346 8880 17789 8936
rect 15285 8878 17789 8880
rect 15285 8875 15351 8878
rect 16989 8848 17789 8878
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 16205 8258 16271 8261
rect 16989 8258 17789 8288
rect 16205 8256 17789 8258
rect 16205 8200 16210 8256
rect 16266 8200 17789 8256
rect 16205 8198 17789 8200
rect 16205 8195 16271 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 16989 8168 17789 8198
rect 4210 8127 4526 8128
rect 5257 7850 5323 7853
rect 13261 7850 13327 7853
rect 14457 7850 14523 7853
rect 5257 7848 5458 7850
rect 5257 7792 5262 7848
rect 5318 7792 5458 7848
rect 5257 7790 5458 7792
rect 5257 7787 5323 7790
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 4061 7442 4127 7445
rect 5165 7442 5231 7445
rect 5398 7442 5458 7790
rect 13261 7848 14523 7850
rect 13261 7792 13266 7848
rect 13322 7792 14462 7848
rect 14518 7792 14523 7848
rect 13261 7790 14523 7792
rect 13261 7787 13327 7790
rect 14457 7787 14523 7790
rect 12801 7578 12867 7581
rect 16989 7578 17789 7608
rect 12801 7576 17789 7578
rect 12801 7520 12806 7576
rect 12862 7520 17789 7576
rect 12801 7518 17789 7520
rect 12801 7515 12867 7518
rect 16989 7488 17789 7518
rect 4061 7440 5458 7442
rect 4061 7384 4066 7440
rect 4122 7384 5170 7440
rect 5226 7384 5458 7440
rect 4061 7382 5458 7384
rect 4061 7379 4127 7382
rect 5165 7379 5231 7382
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 14457 6898 14523 6901
rect 14590 6898 14596 6900
rect 14457 6896 14596 6898
rect 14457 6840 14462 6896
rect 14518 6840 14596 6896
rect 14457 6838 14596 6840
rect 14457 6835 14523 6838
rect 14590 6836 14596 6838
rect 14660 6836 14666 6900
rect 15193 6898 15259 6901
rect 16989 6898 17789 6928
rect 15193 6896 17789 6898
rect 15193 6840 15198 6896
rect 15254 6840 17789 6896
rect 15193 6838 17789 6840
rect 15193 6835 15259 6838
rect 16989 6808 17789 6838
rect 2957 6762 3023 6765
rect 5349 6762 5415 6765
rect 2957 6760 5415 6762
rect 2957 6704 2962 6760
rect 3018 6704 5354 6760
rect 5410 6704 5415 6760
rect 2957 6702 5415 6704
rect 2957 6699 3023 6702
rect 5349 6699 5415 6702
rect 13353 6626 13419 6629
rect 15285 6626 15351 6629
rect 13353 6624 15351 6626
rect 13353 6568 13358 6624
rect 13414 6568 15290 6624
rect 15346 6568 15351 6624
rect 13353 6566 15351 6568
rect 13353 6563 13419 6566
rect 15285 6563 15351 6566
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 9438 6428 9444 6492
rect 9508 6490 9514 6492
rect 15653 6490 15719 6493
rect 9508 6488 15719 6490
rect 9508 6432 15658 6488
rect 15714 6432 15719 6488
rect 9508 6430 15719 6432
rect 9508 6428 9514 6430
rect 15653 6427 15719 6430
rect 13169 6354 13235 6357
rect 15009 6354 15075 6357
rect 15377 6354 15443 6357
rect 13169 6352 15443 6354
rect 13169 6296 13174 6352
rect 13230 6296 15014 6352
rect 15070 6296 15382 6352
rect 15438 6296 15443 6352
rect 13169 6294 15443 6296
rect 13169 6291 13235 6294
rect 15009 6291 15075 6294
rect 15377 6291 15443 6294
rect 15193 6218 15259 6221
rect 16989 6218 17789 6248
rect 15193 6216 17789 6218
rect 15193 6160 15198 6216
rect 15254 6160 17789 6216
rect 15193 6158 17789 6160
rect 15193 6155 15259 6158
rect 16989 6128 17789 6158
rect 7741 6082 7807 6085
rect 14733 6082 14799 6085
rect 7741 6080 14799 6082
rect 7741 6024 7746 6080
rect 7802 6024 14738 6080
rect 14794 6024 14799 6080
rect 7741 6022 14799 6024
rect 7741 6019 7807 6022
rect 14733 6019 14799 6022
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 12801 5946 12867 5949
rect 16205 5946 16271 5949
rect 12801 5944 16271 5946
rect 12801 5888 12806 5944
rect 12862 5888 16210 5944
rect 16266 5888 16271 5944
rect 12801 5886 16271 5888
rect 12801 5883 12867 5886
rect 16205 5883 16271 5886
rect 11237 5810 11303 5813
rect 15469 5810 15535 5813
rect 15653 5810 15719 5813
rect 11237 5808 15719 5810
rect 11237 5752 11242 5808
rect 11298 5752 15474 5808
rect 15530 5752 15658 5808
rect 15714 5752 15719 5808
rect 11237 5750 15719 5752
rect 11237 5747 11303 5750
rect 15469 5747 15535 5750
rect 15653 5747 15719 5750
rect 14733 5676 14799 5677
rect 14733 5674 14780 5676
rect 14688 5672 14780 5674
rect 14688 5616 14738 5672
rect 14688 5614 14780 5616
rect 14733 5612 14780 5614
rect 14844 5612 14850 5676
rect 14733 5611 14799 5612
rect 12341 5538 12407 5541
rect 16989 5538 17789 5568
rect 12341 5536 17789 5538
rect 12341 5480 12346 5536
rect 12402 5480 17789 5536
rect 12341 5478 17789 5480
rect 12341 5475 12407 5478
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 16989 5448 17789 5478
rect 4870 5407 5186 5408
rect 11973 5404 12039 5405
rect 11973 5402 12020 5404
rect 11928 5400 12020 5402
rect 11928 5344 11978 5400
rect 11928 5342 12020 5344
rect 11973 5340 12020 5342
rect 12084 5340 12090 5404
rect 12566 5340 12572 5404
rect 12636 5402 12642 5404
rect 12985 5402 13051 5405
rect 12636 5400 13051 5402
rect 12636 5344 12990 5400
rect 13046 5344 13051 5400
rect 12636 5342 13051 5344
rect 12636 5340 12642 5342
rect 11973 5339 12039 5340
rect 12985 5339 13051 5342
rect 13813 5402 13879 5405
rect 15193 5402 15259 5405
rect 13813 5400 15259 5402
rect 13813 5344 13818 5400
rect 13874 5344 15198 5400
rect 15254 5344 15259 5400
rect 13813 5342 15259 5344
rect 13813 5339 13879 5342
rect 15193 5339 15259 5342
rect 12750 5204 12756 5268
rect 12820 5266 12826 5268
rect 12893 5266 12959 5269
rect 12820 5264 12959 5266
rect 12820 5208 12898 5264
rect 12954 5208 12959 5264
rect 12820 5206 12959 5208
rect 12820 5204 12826 5206
rect 12893 5203 12959 5206
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 16205 4858 16271 4861
rect 16989 4858 17789 4888
rect 16205 4856 17789 4858
rect 16205 4800 16210 4856
rect 16266 4800 17789 4856
rect 16205 4798 17789 4800
rect 16205 4795 16271 4798
rect 16989 4768 17789 4798
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 11462 4252 11468 4316
rect 11532 4314 11538 4316
rect 11605 4314 11671 4317
rect 11532 4312 11671 4314
rect 11532 4256 11610 4312
rect 11666 4256 11671 4312
rect 11532 4254 11671 4256
rect 11532 4252 11538 4254
rect 11605 4251 11671 4254
rect 15193 4178 15259 4181
rect 16989 4178 17789 4208
rect 15193 4176 17789 4178
rect 15193 4120 15198 4176
rect 15254 4120 17789 4176
rect 15193 4118 17789 4120
rect 15193 4115 15259 4118
rect 16989 4088 17789 4118
rect 8753 4042 8819 4045
rect 9070 4042 9076 4044
rect 8753 4040 9076 4042
rect 8753 3984 8758 4040
rect 8814 3984 9076 4040
rect 8753 3982 9076 3984
rect 8753 3979 8819 3982
rect 9070 3980 9076 3982
rect 9140 3980 9146 4044
rect 14406 3980 14412 4044
rect 14476 4042 14482 4044
rect 14733 4042 14799 4045
rect 14476 4040 14799 4042
rect 14476 3984 14738 4040
rect 14794 3984 14799 4040
rect 14476 3982 14799 3984
rect 14476 3980 14482 3982
rect 14733 3979 14799 3982
rect 14958 3980 14964 4044
rect 15028 4042 15034 4044
rect 15653 4042 15719 4045
rect 15028 4040 15719 4042
rect 15028 3984 15658 4040
rect 15714 3984 15719 4040
rect 15028 3982 15719 3984
rect 15028 3980 15034 3982
rect 15653 3979 15719 3982
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 14825 3498 14891 3501
rect 16989 3498 17789 3528
rect 14825 3496 17789 3498
rect 14825 3440 14830 3496
rect 14886 3440 17789 3496
rect 14825 3438 17789 3440
rect 14825 3435 14891 3438
rect 16989 3408 17789 3438
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
<< via3 >>
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 4876 32668 4940 32672
rect 4876 32612 4880 32668
rect 4880 32612 4936 32668
rect 4936 32612 4940 32668
rect 4876 32608 4940 32612
rect 4956 32668 5020 32672
rect 4956 32612 4960 32668
rect 4960 32612 5016 32668
rect 5016 32612 5020 32668
rect 4956 32608 5020 32612
rect 5036 32668 5100 32672
rect 5036 32612 5040 32668
rect 5040 32612 5096 32668
rect 5096 32612 5100 32668
rect 5036 32608 5100 32612
rect 5116 32668 5180 32672
rect 5116 32612 5120 32668
rect 5120 32612 5176 32668
rect 5176 32612 5180 32668
rect 5116 32608 5180 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 8156 31860 8220 31924
rect 13860 31920 13924 31924
rect 13860 31864 13874 31920
rect 13874 31864 13924 31920
rect 13860 31860 13924 31864
rect 7788 31724 7852 31788
rect 4876 31580 4940 31584
rect 4876 31524 4880 31580
rect 4880 31524 4936 31580
rect 4936 31524 4940 31580
rect 4876 31520 4940 31524
rect 4956 31580 5020 31584
rect 4956 31524 4960 31580
rect 4960 31524 5016 31580
rect 5016 31524 5020 31580
rect 4956 31520 5020 31524
rect 5036 31580 5100 31584
rect 5036 31524 5040 31580
rect 5040 31524 5096 31580
rect 5096 31524 5100 31580
rect 5036 31520 5100 31524
rect 5116 31580 5180 31584
rect 5116 31524 5120 31580
rect 5120 31524 5176 31580
rect 5176 31524 5180 31580
rect 5116 31520 5180 31524
rect 13492 31452 13556 31516
rect 796 31316 860 31380
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 14228 30500 14292 30564
rect 4876 30492 4940 30496
rect 4876 30436 4880 30492
rect 4880 30436 4936 30492
rect 4936 30436 4940 30492
rect 4876 30432 4940 30436
rect 4956 30492 5020 30496
rect 4956 30436 4960 30492
rect 4960 30436 5016 30492
rect 5016 30436 5020 30492
rect 4956 30432 5020 30436
rect 5036 30492 5100 30496
rect 5036 30436 5040 30492
rect 5040 30436 5096 30492
rect 5096 30436 5100 30492
rect 5036 30432 5100 30436
rect 5116 30492 5180 30496
rect 5116 30436 5120 30492
rect 5120 30436 5176 30492
rect 5176 30436 5180 30492
rect 5116 30432 5180 30436
rect 10732 30424 10796 30428
rect 10732 30368 10782 30424
rect 10782 30368 10796 30424
rect 10732 30364 10796 30368
rect 796 30092 860 30156
rect 14044 30152 14108 30156
rect 14044 30096 14094 30152
rect 14094 30096 14108 30152
rect 14044 30092 14108 30096
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 12020 29412 12084 29476
rect 4876 29404 4940 29408
rect 4876 29348 4880 29404
rect 4880 29348 4936 29404
rect 4936 29348 4940 29404
rect 4876 29344 4940 29348
rect 4956 29404 5020 29408
rect 4956 29348 4960 29404
rect 4960 29348 5016 29404
rect 5016 29348 5020 29404
rect 4956 29344 5020 29348
rect 5036 29404 5100 29408
rect 5036 29348 5040 29404
rect 5040 29348 5096 29404
rect 5096 29348 5100 29404
rect 5036 29344 5100 29348
rect 5116 29404 5180 29408
rect 5116 29348 5120 29404
rect 5120 29348 5176 29404
rect 5176 29348 5180 29404
rect 5116 29344 5180 29348
rect 9444 29140 9508 29204
rect 11836 29004 11900 29068
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 4876 28316 4940 28320
rect 4876 28260 4880 28316
rect 4880 28260 4936 28316
rect 4936 28260 4940 28316
rect 4876 28256 4940 28260
rect 4956 28316 5020 28320
rect 4956 28260 4960 28316
rect 4960 28260 5016 28316
rect 5016 28260 5020 28316
rect 4956 28256 5020 28260
rect 5036 28316 5100 28320
rect 5036 28260 5040 28316
rect 5040 28260 5096 28316
rect 5096 28260 5100 28316
rect 5036 28256 5100 28260
rect 5116 28316 5180 28320
rect 5116 28260 5120 28316
rect 5120 28260 5176 28316
rect 5176 28260 5180 28316
rect 5116 28256 5180 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 12572 27644 12636 27708
rect 13860 27236 13924 27300
rect 4876 27228 4940 27232
rect 4876 27172 4880 27228
rect 4880 27172 4936 27228
rect 4936 27172 4940 27228
rect 4876 27168 4940 27172
rect 4956 27228 5020 27232
rect 4956 27172 4960 27228
rect 4960 27172 5016 27228
rect 5016 27172 5020 27228
rect 4956 27168 5020 27172
rect 5036 27228 5100 27232
rect 5036 27172 5040 27228
rect 5040 27172 5096 27228
rect 5096 27172 5100 27228
rect 5036 27168 5100 27172
rect 5116 27228 5180 27232
rect 5116 27172 5120 27228
rect 5120 27172 5176 27228
rect 5176 27172 5180 27228
rect 5116 27168 5180 27172
rect 13492 26888 13556 26892
rect 13492 26832 13506 26888
rect 13506 26832 13556 26888
rect 13492 26828 13556 26832
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 14228 26420 14292 26484
rect 14780 26284 14844 26348
rect 4876 26140 4940 26144
rect 4876 26084 4880 26140
rect 4880 26084 4936 26140
rect 4936 26084 4940 26140
rect 4876 26080 4940 26084
rect 4956 26140 5020 26144
rect 4956 26084 4960 26140
rect 4960 26084 5016 26140
rect 5016 26084 5020 26140
rect 4956 26080 5020 26084
rect 5036 26140 5100 26144
rect 5036 26084 5040 26140
rect 5040 26084 5096 26140
rect 5096 26084 5100 26140
rect 5036 26080 5100 26084
rect 5116 26140 5180 26144
rect 5116 26084 5120 26140
rect 5120 26084 5176 26140
rect 5176 26084 5180 26140
rect 5116 26080 5180 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 7788 25468 7852 25532
rect 8156 25528 8220 25532
rect 8156 25472 8170 25528
rect 8170 25472 8220 25528
rect 8156 25468 8220 25472
rect 14596 25332 14660 25396
rect 4876 25052 4940 25056
rect 4876 24996 4880 25052
rect 4880 24996 4936 25052
rect 4936 24996 4940 25052
rect 4876 24992 4940 24996
rect 4956 25052 5020 25056
rect 4956 24996 4960 25052
rect 4960 24996 5016 25052
rect 5016 24996 5020 25052
rect 4956 24992 5020 24996
rect 5036 25052 5100 25056
rect 5036 24996 5040 25052
rect 5040 24996 5096 25052
rect 5096 24996 5100 25052
rect 5036 24992 5100 24996
rect 5116 25052 5180 25056
rect 5116 24996 5120 25052
rect 5120 24996 5176 25052
rect 5176 24996 5180 25052
rect 5116 24992 5180 24996
rect 10916 24984 10980 24988
rect 10916 24928 10966 24984
rect 10966 24928 10980 24984
rect 10916 24924 10980 24928
rect 12204 24924 12268 24988
rect 14044 24924 14108 24988
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 3924 24304 3988 24308
rect 3924 24248 3974 24304
rect 3974 24248 3988 24304
rect 3924 24244 3988 24248
rect 3188 24108 3252 24172
rect 4876 23964 4940 23968
rect 4876 23908 4880 23964
rect 4880 23908 4936 23964
rect 4936 23908 4940 23964
rect 4876 23904 4940 23908
rect 4956 23964 5020 23968
rect 4956 23908 4960 23964
rect 4960 23908 5016 23964
rect 5016 23908 5020 23964
rect 4956 23904 5020 23908
rect 5036 23964 5100 23968
rect 5036 23908 5040 23964
rect 5040 23908 5096 23964
rect 5096 23908 5100 23964
rect 5036 23904 5100 23908
rect 5116 23964 5180 23968
rect 5116 23908 5120 23964
rect 5120 23908 5176 23964
rect 5176 23908 5180 23964
rect 5116 23904 5180 23908
rect 12940 23564 13004 23628
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 14780 23156 14844 23220
rect 9076 23020 9140 23084
rect 11652 23020 11716 23084
rect 4876 22876 4940 22880
rect 4876 22820 4880 22876
rect 4880 22820 4936 22876
rect 4936 22820 4940 22876
rect 4876 22816 4940 22820
rect 4956 22876 5020 22880
rect 4956 22820 4960 22876
rect 4960 22820 5016 22876
rect 5016 22820 5020 22876
rect 4956 22816 5020 22820
rect 5036 22876 5100 22880
rect 5036 22820 5040 22876
rect 5040 22820 5096 22876
rect 5096 22820 5100 22876
rect 5036 22816 5100 22820
rect 5116 22876 5180 22880
rect 5116 22820 5120 22876
rect 5120 22820 5176 22876
rect 5176 22820 5180 22876
rect 5116 22816 5180 22820
rect 11468 22748 11532 22812
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 11836 22068 11900 22132
rect 14780 22068 14844 22132
rect 13124 21932 13188 21996
rect 4876 21788 4940 21792
rect 4876 21732 4880 21788
rect 4880 21732 4936 21788
rect 4936 21732 4940 21788
rect 4876 21728 4940 21732
rect 4956 21788 5020 21792
rect 4956 21732 4960 21788
rect 4960 21732 5016 21788
rect 5016 21732 5020 21788
rect 4956 21728 5020 21732
rect 5036 21788 5100 21792
rect 5036 21732 5040 21788
rect 5040 21732 5096 21788
rect 5096 21732 5100 21788
rect 5036 21728 5100 21732
rect 5116 21788 5180 21792
rect 5116 21732 5120 21788
rect 5120 21732 5176 21788
rect 5176 21732 5180 21788
rect 5116 21728 5180 21732
rect 12020 21388 12084 21452
rect 13492 21388 13556 21452
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 12572 21116 12636 21180
rect 9260 20708 9324 20772
rect 4876 20700 4940 20704
rect 4876 20644 4880 20700
rect 4880 20644 4936 20700
rect 4936 20644 4940 20700
rect 4876 20640 4940 20644
rect 4956 20700 5020 20704
rect 4956 20644 4960 20700
rect 4960 20644 5016 20700
rect 5016 20644 5020 20700
rect 4956 20640 5020 20644
rect 5036 20700 5100 20704
rect 5036 20644 5040 20700
rect 5040 20644 5096 20700
rect 5096 20644 5100 20700
rect 5036 20640 5100 20644
rect 5116 20700 5180 20704
rect 5116 20644 5120 20700
rect 5120 20644 5176 20700
rect 5176 20644 5180 20700
rect 5116 20640 5180 20644
rect 3924 20572 3988 20636
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 4876 19612 4940 19616
rect 4876 19556 4880 19612
rect 4880 19556 4936 19612
rect 4936 19556 4940 19612
rect 4876 19552 4940 19556
rect 4956 19612 5020 19616
rect 4956 19556 4960 19612
rect 4960 19556 5016 19612
rect 5016 19556 5020 19612
rect 4956 19552 5020 19556
rect 5036 19612 5100 19616
rect 5036 19556 5040 19612
rect 5040 19556 5096 19612
rect 5096 19556 5100 19612
rect 5036 19552 5100 19556
rect 5116 19612 5180 19616
rect 5116 19556 5120 19612
rect 5120 19556 5176 19612
rect 5176 19556 5180 19612
rect 5116 19552 5180 19556
rect 12204 19408 12268 19412
rect 12204 19352 12218 19408
rect 12218 19352 12268 19408
rect 12204 19348 12268 19352
rect 3924 19212 3988 19276
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 15332 18864 15396 18868
rect 15332 18808 15382 18864
rect 15382 18808 15396 18864
rect 15332 18804 15396 18808
rect 13676 18668 13740 18732
rect 4876 18524 4940 18528
rect 4876 18468 4880 18524
rect 4880 18468 4936 18524
rect 4936 18468 4940 18524
rect 4876 18464 4940 18468
rect 4956 18524 5020 18528
rect 4956 18468 4960 18524
rect 4960 18468 5016 18524
rect 5016 18468 5020 18524
rect 4956 18464 5020 18468
rect 5036 18524 5100 18528
rect 5036 18468 5040 18524
rect 5040 18468 5096 18524
rect 5096 18468 5100 18524
rect 5036 18464 5100 18468
rect 5116 18524 5180 18528
rect 5116 18468 5120 18524
rect 5120 18468 5176 18524
rect 5176 18468 5180 18524
rect 5116 18464 5180 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 13124 17852 13188 17916
rect 10732 17716 10796 17780
rect 4876 17436 4940 17440
rect 4876 17380 4880 17436
rect 4880 17380 4936 17436
rect 4936 17380 4940 17436
rect 4876 17376 4940 17380
rect 4956 17436 5020 17440
rect 4956 17380 4960 17436
rect 4960 17380 5016 17436
rect 5016 17380 5020 17436
rect 4956 17376 5020 17380
rect 5036 17436 5100 17440
rect 5036 17380 5040 17436
rect 5040 17380 5096 17436
rect 5096 17380 5100 17436
rect 5036 17376 5100 17380
rect 5116 17436 5180 17440
rect 5116 17380 5120 17436
rect 5120 17380 5176 17436
rect 5176 17380 5180 17436
rect 5116 17376 5180 17380
rect 3188 17232 3252 17236
rect 3188 17176 3202 17232
rect 3202 17176 3252 17232
rect 3188 17172 3252 17176
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 14228 16764 14292 16828
rect 10916 16628 10980 16692
rect 14964 16628 15028 16692
rect 9260 16552 9324 16556
rect 9260 16496 9310 16552
rect 9310 16496 9324 16552
rect 9260 16492 9324 16496
rect 4876 16348 4940 16352
rect 4876 16292 4880 16348
rect 4880 16292 4936 16348
rect 4936 16292 4940 16348
rect 4876 16288 4940 16292
rect 4956 16348 5020 16352
rect 4956 16292 4960 16348
rect 4960 16292 5016 16348
rect 5016 16292 5020 16348
rect 4956 16288 5020 16292
rect 5036 16348 5100 16352
rect 5036 16292 5040 16348
rect 5040 16292 5096 16348
rect 5096 16292 5100 16348
rect 5036 16288 5100 16292
rect 5116 16348 5180 16352
rect 5116 16292 5120 16348
rect 5120 16292 5176 16348
rect 5176 16292 5180 16348
rect 5116 16288 5180 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 3188 15676 3252 15740
rect 15332 15600 15396 15604
rect 15332 15544 15346 15600
rect 15346 15544 15396 15600
rect 15332 15540 15396 15544
rect 4660 15404 4724 15468
rect 5764 15328 5828 15332
rect 5764 15272 5814 15328
rect 5814 15272 5828 15328
rect 5764 15268 5828 15272
rect 12756 15268 12820 15332
rect 4876 15260 4940 15264
rect 4876 15204 4880 15260
rect 4880 15204 4936 15260
rect 4936 15204 4940 15260
rect 4876 15200 4940 15204
rect 4956 15260 5020 15264
rect 4956 15204 4960 15260
rect 4960 15204 5016 15260
rect 5016 15204 5020 15260
rect 4956 15200 5020 15204
rect 5036 15260 5100 15264
rect 5036 15204 5040 15260
rect 5040 15204 5096 15260
rect 5096 15204 5100 15260
rect 5036 15200 5100 15204
rect 5116 15260 5180 15264
rect 5116 15204 5120 15260
rect 5120 15204 5176 15260
rect 5176 15204 5180 15260
rect 5116 15200 5180 15204
rect 12204 15132 12268 15196
rect 12020 14996 12084 15060
rect 14228 14996 14292 15060
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 3372 14316 3436 14380
rect 4876 14172 4940 14176
rect 4876 14116 4880 14172
rect 4880 14116 4936 14172
rect 4936 14116 4940 14172
rect 4876 14112 4940 14116
rect 4956 14172 5020 14176
rect 4956 14116 4960 14172
rect 4960 14116 5016 14172
rect 5016 14116 5020 14172
rect 4956 14112 5020 14116
rect 5036 14172 5100 14176
rect 5036 14116 5040 14172
rect 5040 14116 5096 14172
rect 5096 14116 5100 14172
rect 5036 14112 5100 14116
rect 5116 14172 5180 14176
rect 5116 14116 5120 14172
rect 5120 14116 5176 14172
rect 5176 14116 5180 14172
rect 5116 14112 5180 14116
rect 3740 13908 3804 13972
rect 3924 13636 3988 13700
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 11652 13364 11716 13428
rect 4876 13084 4940 13088
rect 4876 13028 4880 13084
rect 4880 13028 4936 13084
rect 4936 13028 4940 13084
rect 4876 13024 4940 13028
rect 4956 13084 5020 13088
rect 4956 13028 4960 13084
rect 4960 13028 5016 13084
rect 5016 13028 5020 13084
rect 4956 13024 5020 13028
rect 5036 13084 5100 13088
rect 5036 13028 5040 13084
rect 5040 13028 5096 13084
rect 5096 13028 5100 13084
rect 5036 13024 5100 13028
rect 5116 13084 5180 13088
rect 5116 13028 5120 13084
rect 5120 13028 5176 13084
rect 5176 13028 5180 13084
rect 5116 13024 5180 13028
rect 5764 12820 5828 12884
rect 14412 12548 14476 12612
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 3372 12336 3436 12340
rect 3372 12280 3422 12336
rect 3422 12280 3436 12336
rect 3372 12276 3436 12280
rect 9076 12336 9140 12340
rect 9076 12280 9126 12336
rect 9126 12280 9140 12336
rect 9076 12276 9140 12280
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 9076 11460 9140 11524
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 3740 11188 3804 11252
rect 12572 10916 12636 10980
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 4660 10644 4724 10708
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 13676 10100 13740 10164
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 12940 9752 13004 9756
rect 12940 9696 12954 9752
rect 12954 9696 13004 9752
rect 12940 9692 13004 9696
rect 13492 9420 13556 9484
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 14596 6836 14660 6900
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 9444 6428 9508 6492
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 14780 5672 14844 5676
rect 14780 5616 14794 5672
rect 14794 5616 14844 5672
rect 14780 5612 14844 5616
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 12020 5400 12084 5404
rect 12020 5344 12034 5400
rect 12034 5344 12084 5400
rect 12020 5340 12084 5344
rect 12572 5340 12636 5404
rect 12756 5204 12820 5268
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 11468 4252 11532 4316
rect 9076 3980 9140 4044
rect 14412 3980 14476 4044
rect 14964 3980 15028 4044
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
<< metal4 >>
rect 4208 33216 4528 33232
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 795 31380 861 31381
rect 795 31316 796 31380
rect 860 31316 861 31380
rect 795 31315 861 31316
rect 798 30157 858 31315
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 795 30156 861 30157
rect 795 30092 796 30156
rect 860 30092 861 30156
rect 795 30091 861 30092
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 3923 24308 3989 24309
rect 3923 24244 3924 24308
rect 3988 24244 3989 24308
rect 3923 24243 3989 24244
rect 3187 24172 3253 24173
rect 3187 24108 3188 24172
rect 3252 24108 3253 24172
rect 3187 24107 3253 24108
rect 3190 17237 3250 24107
rect 3926 20637 3986 24243
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 3923 20636 3989 20637
rect 3923 20572 3924 20636
rect 3988 20572 3989 20636
rect 3923 20571 3989 20572
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 3923 19276 3989 19277
rect 3923 19212 3924 19276
rect 3988 19212 3989 19276
rect 3923 19211 3989 19212
rect 3187 17236 3253 17237
rect 3187 17172 3188 17236
rect 3252 17172 3253 17236
rect 3187 17171 3253 17172
rect 3190 15741 3250 17171
rect 3187 15740 3253 15741
rect 3187 15676 3188 15740
rect 3252 15676 3253 15740
rect 3187 15675 3253 15676
rect 3190 15330 3250 15675
rect 3190 15270 3434 15330
rect 3374 14381 3434 15270
rect 3371 14380 3437 14381
rect 3371 14316 3372 14380
rect 3436 14316 3437 14380
rect 3371 14315 3437 14316
rect 3374 12341 3434 14315
rect 3739 13972 3805 13973
rect 3739 13908 3740 13972
rect 3804 13908 3805 13972
rect 3739 13907 3805 13908
rect 3371 12340 3437 12341
rect 3371 12276 3372 12340
rect 3436 12276 3437 12340
rect 3371 12275 3437 12276
rect 3742 11253 3802 13907
rect 3926 13701 3986 19211
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4868 32672 5188 33232
rect 4868 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5188 32672
rect 4868 31584 5188 32608
rect 8155 31924 8221 31925
rect 8155 31860 8156 31924
rect 8220 31860 8221 31924
rect 8155 31859 8221 31860
rect 13859 31924 13925 31925
rect 13859 31860 13860 31924
rect 13924 31860 13925 31924
rect 13859 31859 13925 31860
rect 7787 31788 7853 31789
rect 7787 31724 7788 31788
rect 7852 31724 7853 31788
rect 7787 31723 7853 31724
rect 4868 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5188 31584
rect 4868 30496 5188 31520
rect 4868 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5188 30496
rect 4868 29408 5188 30432
rect 4868 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5188 29408
rect 4868 28320 5188 29344
rect 4868 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5188 28320
rect 4868 27232 5188 28256
rect 4868 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5188 27232
rect 4868 26144 5188 27168
rect 4868 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5188 26144
rect 4868 25056 5188 26080
rect 7790 25533 7850 31723
rect 8158 25533 8218 31859
rect 13491 31516 13557 31517
rect 13491 31452 13492 31516
rect 13556 31452 13557 31516
rect 13491 31451 13557 31452
rect 10731 30428 10797 30429
rect 10731 30364 10732 30428
rect 10796 30364 10797 30428
rect 10731 30363 10797 30364
rect 9443 29204 9509 29205
rect 9443 29140 9444 29204
rect 9508 29140 9509 29204
rect 9443 29139 9509 29140
rect 7787 25532 7853 25533
rect 7787 25468 7788 25532
rect 7852 25468 7853 25532
rect 7787 25467 7853 25468
rect 8155 25532 8221 25533
rect 8155 25468 8156 25532
rect 8220 25468 8221 25532
rect 8155 25467 8221 25468
rect 4868 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5188 25056
rect 4868 23968 5188 24992
rect 4868 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5188 23968
rect 4868 22880 5188 23904
rect 9075 23084 9141 23085
rect 9075 23020 9076 23084
rect 9140 23020 9141 23084
rect 9075 23019 9141 23020
rect 4868 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5188 22880
rect 4868 21792 5188 22816
rect 4868 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5188 21792
rect 4868 20704 5188 21728
rect 4868 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5188 20704
rect 4868 19616 5188 20640
rect 4868 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5188 19616
rect 4868 18528 5188 19552
rect 4868 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5188 18528
rect 4868 17440 5188 18464
rect 4868 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5188 17440
rect 4868 16352 5188 17376
rect 4868 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5188 16352
rect 4659 15468 4725 15469
rect 4659 15404 4660 15468
rect 4724 15404 4725 15468
rect 4659 15403 4725 15404
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 3923 13700 3989 13701
rect 3923 13636 3924 13700
rect 3988 13636 3989 13700
rect 3923 13635 3989 13636
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 3739 11252 3805 11253
rect 3739 11188 3740 11252
rect 3804 11188 3805 11252
rect 3739 11187 3805 11188
rect 4208 10368 4528 11392
rect 4662 10709 4722 15403
rect 4868 15264 5188 16288
rect 5763 15332 5829 15333
rect 5763 15268 5764 15332
rect 5828 15268 5829 15332
rect 5763 15267 5829 15268
rect 4868 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5188 15264
rect 4868 14176 5188 15200
rect 4868 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5188 14176
rect 4868 13088 5188 14112
rect 4868 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5188 13088
rect 4868 12000 5188 13024
rect 5766 12885 5826 15267
rect 5763 12884 5829 12885
rect 5763 12820 5764 12884
rect 5828 12820 5829 12884
rect 5763 12819 5829 12820
rect 9078 12341 9138 23019
rect 9259 20772 9325 20773
rect 9259 20708 9260 20772
rect 9324 20708 9325 20772
rect 9259 20707 9325 20708
rect 9262 16557 9322 20707
rect 9259 16556 9325 16557
rect 9259 16492 9260 16556
rect 9324 16492 9325 16556
rect 9259 16491 9325 16492
rect 9075 12340 9141 12341
rect 9075 12276 9076 12340
rect 9140 12276 9141 12340
rect 9075 12275 9141 12276
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4868 10912 5188 11936
rect 9075 11524 9141 11525
rect 9075 11460 9076 11524
rect 9140 11460 9141 11524
rect 9075 11459 9141 11460
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4659 10708 4725 10709
rect 4659 10644 4660 10708
rect 4724 10644 4725 10708
rect 4659 10643 4725 10644
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 9824 5188 10848
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 5472 5188 6496
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 9078 4045 9138 11459
rect 9446 6493 9506 29139
rect 10734 17781 10794 30363
rect 12019 29476 12085 29477
rect 12019 29412 12020 29476
rect 12084 29412 12085 29476
rect 12019 29411 12085 29412
rect 11835 29068 11901 29069
rect 11835 29004 11836 29068
rect 11900 29004 11901 29068
rect 11835 29003 11901 29004
rect 10915 24988 10981 24989
rect 10915 24924 10916 24988
rect 10980 24924 10981 24988
rect 10915 24923 10981 24924
rect 10731 17780 10797 17781
rect 10731 17716 10732 17780
rect 10796 17716 10797 17780
rect 10731 17715 10797 17716
rect 10918 16693 10978 24923
rect 11651 23084 11717 23085
rect 11651 23020 11652 23084
rect 11716 23020 11717 23084
rect 11651 23019 11717 23020
rect 11467 22812 11533 22813
rect 11467 22748 11468 22812
rect 11532 22748 11533 22812
rect 11467 22747 11533 22748
rect 10915 16692 10981 16693
rect 10915 16628 10916 16692
rect 10980 16628 10981 16692
rect 10915 16627 10981 16628
rect 9443 6492 9509 6493
rect 9443 6428 9444 6492
rect 9508 6428 9509 6492
rect 9443 6427 9509 6428
rect 11470 4317 11530 22747
rect 11654 13429 11714 23019
rect 11838 22133 11898 29003
rect 11835 22132 11901 22133
rect 11835 22068 11836 22132
rect 11900 22068 11901 22132
rect 11835 22067 11901 22068
rect 12022 21453 12082 29411
rect 12571 27708 12637 27709
rect 12571 27644 12572 27708
rect 12636 27644 12637 27708
rect 12571 27643 12637 27644
rect 12203 24988 12269 24989
rect 12203 24924 12204 24988
rect 12268 24924 12269 24988
rect 12203 24923 12269 24924
rect 12019 21452 12085 21453
rect 12019 21388 12020 21452
rect 12084 21388 12085 21452
rect 12019 21387 12085 21388
rect 12206 20090 12266 24923
rect 12574 21181 12634 27643
rect 13494 26893 13554 31451
rect 13862 27301 13922 31859
rect 14227 30564 14293 30565
rect 14227 30500 14228 30564
rect 14292 30500 14293 30564
rect 14227 30499 14293 30500
rect 14043 30156 14109 30157
rect 14043 30092 14044 30156
rect 14108 30092 14109 30156
rect 14043 30091 14109 30092
rect 13859 27300 13925 27301
rect 13859 27236 13860 27300
rect 13924 27236 13925 27300
rect 13859 27235 13925 27236
rect 13491 26892 13557 26893
rect 13491 26828 13492 26892
rect 13556 26828 13557 26892
rect 13491 26827 13557 26828
rect 14046 24989 14106 30091
rect 14230 26485 14290 30499
rect 14227 26484 14293 26485
rect 14227 26420 14228 26484
rect 14292 26420 14293 26484
rect 14227 26419 14293 26420
rect 14779 26348 14845 26349
rect 14779 26284 14780 26348
rect 14844 26284 14845 26348
rect 14779 26283 14845 26284
rect 14595 25396 14661 25397
rect 14595 25332 14596 25396
rect 14660 25332 14661 25396
rect 14595 25331 14661 25332
rect 14043 24988 14109 24989
rect 14043 24924 14044 24988
rect 14108 24924 14109 24988
rect 14043 24923 14109 24924
rect 12939 23628 13005 23629
rect 12939 23564 12940 23628
rect 13004 23564 13005 23628
rect 12939 23563 13005 23564
rect 12571 21180 12637 21181
rect 12571 21116 12572 21180
rect 12636 21116 12637 21180
rect 12571 21115 12637 21116
rect 12022 20030 12266 20090
rect 12022 15061 12082 20030
rect 12203 19412 12269 19413
rect 12203 19348 12204 19412
rect 12268 19348 12269 19412
rect 12203 19347 12269 19348
rect 12206 15197 12266 19347
rect 12755 15332 12821 15333
rect 12755 15268 12756 15332
rect 12820 15268 12821 15332
rect 12755 15267 12821 15268
rect 12203 15196 12269 15197
rect 12203 15132 12204 15196
rect 12268 15132 12269 15196
rect 12203 15131 12269 15132
rect 12019 15060 12085 15061
rect 12019 14996 12020 15060
rect 12084 14996 12085 15060
rect 12019 14995 12085 14996
rect 11651 13428 11717 13429
rect 11651 13364 11652 13428
rect 11716 13364 11717 13428
rect 11651 13363 11717 13364
rect 12022 5405 12082 14995
rect 12571 10980 12637 10981
rect 12571 10916 12572 10980
rect 12636 10916 12637 10980
rect 12571 10915 12637 10916
rect 12574 5405 12634 10915
rect 12019 5404 12085 5405
rect 12019 5340 12020 5404
rect 12084 5340 12085 5404
rect 12019 5339 12085 5340
rect 12571 5404 12637 5405
rect 12571 5340 12572 5404
rect 12636 5340 12637 5404
rect 12571 5339 12637 5340
rect 12758 5269 12818 15267
rect 12942 9757 13002 23563
rect 13123 21996 13189 21997
rect 13123 21932 13124 21996
rect 13188 21932 13189 21996
rect 13123 21931 13189 21932
rect 13126 17917 13186 21931
rect 13491 21452 13557 21453
rect 13491 21388 13492 21452
rect 13556 21388 13557 21452
rect 13491 21387 13557 21388
rect 13123 17916 13189 17917
rect 13123 17852 13124 17916
rect 13188 17852 13189 17916
rect 13123 17851 13189 17852
rect 12939 9756 13005 9757
rect 12939 9692 12940 9756
rect 13004 9692 13005 9756
rect 12939 9691 13005 9692
rect 13494 9485 13554 21387
rect 13675 18732 13741 18733
rect 13675 18668 13676 18732
rect 13740 18668 13741 18732
rect 13675 18667 13741 18668
rect 13678 10165 13738 18667
rect 14227 16828 14293 16829
rect 14227 16764 14228 16828
rect 14292 16764 14293 16828
rect 14227 16763 14293 16764
rect 14230 15061 14290 16763
rect 14227 15060 14293 15061
rect 14227 14996 14228 15060
rect 14292 14996 14293 15060
rect 14227 14995 14293 14996
rect 14411 12612 14477 12613
rect 14411 12548 14412 12612
rect 14476 12548 14477 12612
rect 14411 12547 14477 12548
rect 13675 10164 13741 10165
rect 13675 10100 13676 10164
rect 13740 10100 13741 10164
rect 13675 10099 13741 10100
rect 13491 9484 13557 9485
rect 13491 9420 13492 9484
rect 13556 9420 13557 9484
rect 13491 9419 13557 9420
rect 12755 5268 12821 5269
rect 12755 5204 12756 5268
rect 12820 5204 12821 5268
rect 12755 5203 12821 5204
rect 11467 4316 11533 4317
rect 11467 4252 11468 4316
rect 11532 4252 11533 4316
rect 11467 4251 11533 4252
rect 14414 4045 14474 12547
rect 14598 6901 14658 25331
rect 14782 23221 14842 26283
rect 14779 23220 14845 23221
rect 14779 23156 14780 23220
rect 14844 23156 14845 23220
rect 14779 23155 14845 23156
rect 14779 22132 14845 22133
rect 14779 22068 14780 22132
rect 14844 22068 14845 22132
rect 14779 22067 14845 22068
rect 14595 6900 14661 6901
rect 14595 6836 14596 6900
rect 14660 6836 14661 6900
rect 14595 6835 14661 6836
rect 14782 5677 14842 22067
rect 15331 18868 15397 18869
rect 15331 18804 15332 18868
rect 15396 18804 15397 18868
rect 15331 18803 15397 18804
rect 14963 16692 15029 16693
rect 14963 16628 14964 16692
rect 15028 16628 15029 16692
rect 14963 16627 15029 16628
rect 14779 5676 14845 5677
rect 14779 5612 14780 5676
rect 14844 5612 14845 5676
rect 14779 5611 14845 5612
rect 14966 4045 15026 16627
rect 15334 15605 15394 18803
rect 15331 15604 15397 15605
rect 15331 15540 15332 15604
rect 15396 15540 15397 15604
rect 15331 15539 15397 15540
rect 9075 4044 9141 4045
rect 9075 3980 9076 4044
rect 9140 3980 9141 4044
rect 9075 3979 9141 3980
rect 14411 4044 14477 4045
rect 14411 3980 14412 4044
rect 14476 3980 14477 4044
rect 14411 3979 14477 3980
rect 14963 4044 15029 4045
rect 14963 3980 14964 4044
rect 15028 3980 15029 4044
rect 14963 3979 15029 3980
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
use sky130_fd_sc_hd__inv_2  _0527_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform -1 0 6256 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0528_
timestamp 1730882523
transform 1 0 11500 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0529_
timestamp 1730882523
transform 1 0 12236 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0530_
timestamp 1730882523
transform -1 0 13248 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0531_
timestamp 1730882523
transform -1 0 6900 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0532_
timestamp 1730882523
transform -1 0 9200 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0533_
timestamp 1730882523
transform 1 0 9936 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0534_
timestamp 1730882523
transform 1 0 4140 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0535_
timestamp 1730882523
transform -1 0 6624 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0536_
timestamp 1730882523
transform -1 0 9844 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0537_
timestamp 1730882523
transform 1 0 3772 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0538_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform -1 0 9752 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0539_
timestamp 1730882523
transform 1 0 7820 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _0540_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 10672 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0541_
timestamp 1730882523
transform -1 0 10212 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0542_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform -1 0 10764 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0543_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform -1 0 9752 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0544_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform -1 0 9384 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0545_
timestamp 1730882523
transform 1 0 7820 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0546_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 8188 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0547_
timestamp 1730882523
transform -1 0 4968 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0548_
timestamp 1730882523
transform -1 0 4600 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0549_
timestamp 1730882523
transform 1 0 3220 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0550_
timestamp 1730882523
transform -1 0 4784 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0551_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform -1 0 6072 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _0552_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 5152 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0553_
timestamp 1730882523
transform 1 0 3128 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _0554_
timestamp 1730882523
transform 1 0 3772 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _0555_
timestamp 1730882523
transform 1 0 3588 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _0556_
timestamp 1730882523
transform -1 0 3496 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_4  _0557_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform -1 0 5888 0 -1 18496
box -38 -48 2062 592
use sky130_fd_sc_hd__xor2_1  _0558_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 1748 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0559_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform -1 0 4416 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0560_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 3128 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0561_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform -1 0 3312 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0562_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 3036 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _0563_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 2392 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0564_
timestamp 1730882523
transform 1 0 3312 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _0565_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform -1 0 3404 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _0566_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform -1 0 4508 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nand2b_1  _0567_
timestamp 1730882523
transform -1 0 4416 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0568_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform -1 0 3404 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0569_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 3772 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0570_
timestamp 1730882523
transform 1 0 3404 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0571_
timestamp 1730882523
transform -1 0 3036 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _0572_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 3036 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0573_
timestamp 1730882523
transform -1 0 3680 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o311a_1  _0574_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform -1 0 4508 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a311o_1  _0575_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 3496 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0576_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 3772 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _0577_
timestamp 1730882523
transform 1 0 4508 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0578_
timestamp 1730882523
transform 1 0 2760 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0579_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 3128 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o22ai_1  _0580_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 4508 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0581_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform -1 0 4600 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0582_
timestamp 1730882523
transform 1 0 3680 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a22oi_4  _0583_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 3956 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__nand2_1  _0584_
timestamp 1730882523
transform 1 0 4968 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _0585_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 10948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0586_
timestamp 1730882523
transform 1 0 11316 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0587_
timestamp 1730882523
transform 1 0 11316 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0588_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 11592 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _0589_
timestamp 1730882523
transform -1 0 8740 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_2  _0590_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 8004 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0591_
timestamp 1730882523
transform -1 0 6164 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0592_
timestamp 1730882523
transform 1 0 8556 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _0593_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 9936 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0594_
timestamp 1730882523
transform -1 0 10212 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0595_
timestamp 1730882523
transform 1 0 10396 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _0596_
timestamp 1730882523
transform 1 0 10028 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0597_
timestamp 1730882523
transform 1 0 10396 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0598_
timestamp 1730882523
transform 1 0 8924 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0599_
timestamp 1730882523
transform 1 0 13248 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0600_
timestamp 1730882523
transform 1 0 10948 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0601_
timestamp 1730882523
transform -1 0 8832 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0602_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform -1 0 9384 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0603_
timestamp 1730882523
transform 1 0 8372 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0604_
timestamp 1730882523
transform 1 0 8372 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _0605_
timestamp 1730882523
transform 1 0 10212 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0606_
timestamp 1730882523
transform 1 0 10580 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0607_
timestamp 1730882523
transform 1 0 8464 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0608_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 10396 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0609_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform -1 0 8832 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0610_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 11132 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _0611_
timestamp 1730882523
transform 1 0 10856 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0612_
timestamp 1730882523
transform 1 0 11500 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0613_
timestamp 1730882523
transform 1 0 12144 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0614_
timestamp 1730882523
transform 1 0 7636 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0615_
timestamp 1730882523
transform 1 0 5704 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0616_
timestamp 1730882523
transform 1 0 4692 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0617_
timestamp 1730882523
transform -1 0 5980 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _0618_
timestamp 1730882523
transform 1 0 3128 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0619_
timestamp 1730882523
transform -1 0 3128 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0620_
timestamp 1730882523
transform 1 0 3220 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0621_
timestamp 1730882523
transform 1 0 3956 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0622_
timestamp 1730882523
transform -1 0 4416 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0623_
timestamp 1730882523
transform -1 0 4876 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _0624_
timestamp 1730882523
transform 1 0 3864 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0625_
timestamp 1730882523
transform 1 0 3036 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0626_
timestamp 1730882523
transform 1 0 2852 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0627_
timestamp 1730882523
transform 1 0 4508 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0628_
timestamp 1730882523
transform 1 0 4508 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0629_
timestamp 1730882523
transform 1 0 3220 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _0630_
timestamp 1730882523
transform -1 0 3680 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0631_
timestamp 1730882523
transform 1 0 3772 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0632_
timestamp 1730882523
transform -1 0 3864 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0633_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 3864 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0634_
timestamp 1730882523
transform -1 0 4508 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0635_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 3956 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0636_
timestamp 1730882523
transform -1 0 4692 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0637_
timestamp 1730882523
transform -1 0 4968 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _0638_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform -1 0 5428 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_4  _0639_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform -1 0 6256 0 -1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__o21a_1  _0640_
timestamp 1730882523
transform -1 0 3680 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _0641_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 3772 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _0642_
timestamp 1730882523
transform 1 0 3772 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_1  _0643_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform -1 0 2392 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__xor2_1  _0644_
timestamp 1730882523
transform -1 0 3588 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _0645_
timestamp 1730882523
transform -1 0 3128 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0646_
timestamp 1730882523
transform 1 0 2300 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0647_
timestamp 1730882523
transform -1 0 2300 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0648_
timestamp 1730882523
transform 1 0 2300 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _0649_
timestamp 1730882523
transform -1 0 2300 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _0650_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform -1 0 3220 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0651_
timestamp 1730882523
transform 1 0 2852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0652_
timestamp 1730882523
transform 1 0 2944 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _0653_
timestamp 1730882523
transform -1 0 2392 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _0654_
timestamp 1730882523
transform -1 0 2576 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _0655_
timestamp 1730882523
transform 1 0 1748 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0656_
timestamp 1730882523
transform -1 0 3588 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0657_
timestamp 1730882523
transform -1 0 3680 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0658_
timestamp 1730882523
transform -1 0 1748 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _0659_
timestamp 1730882523
transform -1 0 3312 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _0660_
timestamp 1730882523
transform -1 0 4232 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0661_
timestamp 1730882523
transform 1 0 4232 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0662_
timestamp 1730882523
transform 1 0 3772 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _0663_
timestamp 1730882523
transform 1 0 2484 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _0664_
timestamp 1730882523
transform -1 0 4876 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _0665_
timestamp 1730882523
transform 1 0 3956 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0666_
timestamp 1730882523
transform 1 0 5152 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0667_
timestamp 1730882523
transform -1 0 5796 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0668_
timestamp 1730882523
transform 1 0 5612 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _0669_
timestamp 1730882523
transform 1 0 4692 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _0670_
timestamp 1730882523
transform 1 0 6072 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0671_
timestamp 1730882523
transform 1 0 6348 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0672_
timestamp 1730882523
transform -1 0 5520 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _0673_
timestamp 1730882523
transform 1 0 4600 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0674_
timestamp 1730882523
transform 1 0 6624 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0675_
timestamp 1730882523
transform 1 0 4968 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _0676_
timestamp 1730882523
transform 1 0 5336 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0677_
timestamp 1730882523
transform -1 0 6900 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _0678_
timestamp 1730882523
transform 1 0 5520 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0679_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 5612 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _0680_
timestamp 1730882523
transform 1 0 4968 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _0681_
timestamp 1730882523
transform 1 0 8924 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _0682_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 8924 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _0683_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 9292 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0684_
timestamp 1730882523
transform -1 0 9200 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0685_
timestamp 1730882523
transform 1 0 9568 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_2  _0686_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform -1 0 9568 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0687_
timestamp 1730882523
transform 1 0 13708 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _0688_
timestamp 1730882523
transform 1 0 13340 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _0689_
timestamp 1730882523
transform 1 0 12880 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0690_
timestamp 1730882523
transform 1 0 14076 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0691_
timestamp 1730882523
transform 1 0 14076 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0692_
timestamp 1730882523
transform 1 0 13524 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0693_
timestamp 1730882523
transform -1 0 14812 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0694_
timestamp 1730882523
transform 1 0 14536 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0695_
timestamp 1730882523
transform 1 0 14076 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0696_
timestamp 1730882523
transform -1 0 14628 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0697_
timestamp 1730882523
transform -1 0 13432 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0698_
timestamp 1730882523
transform 1 0 13524 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0699_
timestamp 1730882523
transform 1 0 14076 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0700_
timestamp 1730882523
transform -1 0 14444 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0701_
timestamp 1730882523
transform -1 0 13984 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0702_
timestamp 1730882523
transform -1 0 13616 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0703_
timestamp 1730882523
transform 1 0 13892 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0704_
timestamp 1730882523
transform 1 0 13524 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0705_
timestamp 1730882523
transform 1 0 15548 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__and3_2  _0706_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 14076 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0707_
timestamp 1730882523
transform -1 0 14904 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0708_
timestamp 1730882523
transform -1 0 14996 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0709_
timestamp 1730882523
transform 1 0 15916 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0710_
timestamp 1730882523
transform 1 0 14904 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0711_
timestamp 1730882523
transform 1 0 15824 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0712_
timestamp 1730882523
transform 1 0 15548 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0713_
timestamp 1730882523
transform 1 0 14996 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0714_
timestamp 1730882523
transform 1 0 14812 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0715_
timestamp 1730882523
transform -1 0 16008 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0716_
timestamp 1730882523
transform 1 0 14904 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0717_
timestamp 1730882523
transform 1 0 14628 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0718_
timestamp 1730882523
transform -1 0 15548 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0719_
timestamp 1730882523
transform 1 0 15548 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0720_
timestamp 1730882523
transform 1 0 15548 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0721_
timestamp 1730882523
transform -1 0 12696 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0722_
timestamp 1730882523
transform 1 0 15548 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0723_
timestamp 1730882523
transform -1 0 16192 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0724_
timestamp 1730882523
transform -1 0 14812 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _0725_
timestamp 1730882523
transform 1 0 14076 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0726_
timestamp 1730882523
transform 1 0 13892 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0727_
timestamp 1730882523
transform -1 0 15272 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0728_
timestamp 1730882523
transform -1 0 16008 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0729_
timestamp 1730882523
transform 1 0 14812 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0730_
timestamp 1730882523
transform 1 0 15824 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0731_
timestamp 1730882523
transform -1 0 14904 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0732_
timestamp 1730882523
transform -1 0 16008 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0733_
timestamp 1730882523
transform 1 0 13248 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0734_
timestamp 1730882523
transform 1 0 14352 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0735_
timestamp 1730882523
transform -1 0 14904 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0736_
timestamp 1730882523
transform -1 0 13524 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0737_
timestamp 1730882523
transform 1 0 15456 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0738_
timestamp 1730882523
transform 1 0 15824 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0739_
timestamp 1730882523
transform -1 0 14904 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0740_
timestamp 1730882523
transform 1 0 13524 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0741_
timestamp 1730882523
transform 1 0 14720 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0742_
timestamp 1730882523
transform -1 0 14536 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0743_
timestamp 1730882523
transform -1 0 14812 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__and3_2  _0744_
timestamp 1730882523
transform 1 0 13248 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0745_
timestamp 1730882523
transform -1 0 13984 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0746_
timestamp 1730882523
transform -1 0 13524 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0747_
timestamp 1730882523
transform 1 0 15364 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0748_
timestamp 1730882523
transform 1 0 15548 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0749_
timestamp 1730882523
transform -1 0 13064 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0750_
timestamp 1730882523
transform -1 0 15640 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0751_
timestamp 1730882523
transform -1 0 14536 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0752_
timestamp 1730882523
transform 1 0 13340 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0753_
timestamp 1730882523
transform 1 0 14444 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0754_
timestamp 1730882523
transform 1 0 15456 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0755_
timestamp 1730882523
transform 1 0 13432 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0756_
timestamp 1730882523
transform 1 0 14076 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0757_
timestamp 1730882523
transform 1 0 15364 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0758_
timestamp 1730882523
transform 1 0 15088 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0759_
timestamp 1730882523
transform 1 0 13064 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0760_
timestamp 1730882523
transform 1 0 13248 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0761_
timestamp 1730882523
transform -1 0 13984 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0762_
timestamp 1730882523
transform 1 0 12972 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _0763_
timestamp 1730882523
transform -1 0 14260 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and2_2  _0764_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 13800 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _0765_
timestamp 1730882523
transform 1 0 14628 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0766_
timestamp 1730882523
transform -1 0 15548 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0767_
timestamp 1730882523
transform 1 0 14352 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0768_
timestamp 1730882523
transform 1 0 14996 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0769_
timestamp 1730882523
transform 1 0 15272 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0770_
timestamp 1730882523
transform 1 0 14076 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0771_
timestamp 1730882523
transform 1 0 14076 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0772_
timestamp 1730882523
transform 1 0 15916 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0773_
timestamp 1730882523
transform 1 0 15088 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0774_
timestamp 1730882523
transform -1 0 16192 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0775_
timestamp 1730882523
transform -1 0 14904 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0776_
timestamp 1730882523
transform -1 0 16284 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0777_
timestamp 1730882523
transform 1 0 14352 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0778_
timestamp 1730882523
transform -1 0 13156 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0779_
timestamp 1730882523
transform 1 0 14812 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0780_
timestamp 1730882523
transform -1 0 15824 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0781_
timestamp 1730882523
transform 1 0 14536 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0782_
timestamp 1730882523
transform -1 0 16100 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0783_
timestamp 1730882523
transform -1 0 16284 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0784_
timestamp 1730882523
transform 1 0 14260 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0785_
timestamp 1730882523
transform -1 0 13616 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0786_
timestamp 1730882523
transform -1 0 16284 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0787_
timestamp 1730882523
transform 1 0 15640 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0788_
timestamp 1730882523
transform 1 0 15456 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0789_
timestamp 1730882523
transform 1 0 12512 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0790_
timestamp 1730882523
transform -1 0 15180 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0791_
timestamp 1730882523
transform -1 0 16192 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0792_
timestamp 1730882523
transform 1 0 11132 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0793_
timestamp 1730882523
transform 1 0 12328 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0794_
timestamp 1730882523
transform 1 0 15640 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0795_
timestamp 1730882523
transform 1 0 15548 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0796_
timestamp 1730882523
transform 1 0 15640 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0797_
timestamp 1730882523
transform 1 0 12972 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0798_
timestamp 1730882523
transform -1 0 16192 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0799_
timestamp 1730882523
transform -1 0 15364 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0800_
timestamp 1730882523
transform 1 0 14076 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0801_
timestamp 1730882523
transform 1 0 14260 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0802_
timestamp 1730882523
transform -1 0 16192 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0803_
timestamp 1730882523
transform -1 0 16376 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0804_
timestamp 1730882523
transform 1 0 15088 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0805_
timestamp 1730882523
transform 1 0 11500 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0806_
timestamp 1730882523
transform 1 0 15548 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0807_
timestamp 1730882523
transform 1 0 14076 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0808_
timestamp 1730882523
transform 1 0 14444 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0809_
timestamp 1730882523
transform 1 0 11776 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0810_
timestamp 1730882523
transform 1 0 14076 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0811_
timestamp 1730882523
transform 1 0 15088 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0812_
timestamp 1730882523
transform 1 0 15088 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0813_
timestamp 1730882523
transform 1 0 13156 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0814_
timestamp 1730882523
transform 1 0 12420 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0815_
timestamp 1730882523
transform 1 0 13248 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0816_
timestamp 1730882523
transform 1 0 12604 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _0817_
timestamp 1730882523
transform 1 0 10764 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0818_
timestamp 1730882523
transform 1 0 12972 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _0819_
timestamp 1730882523
transform 1 0 11500 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0820_
timestamp 1730882523
transform 1 0 12512 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _0821_
timestamp 1730882523
transform 1 0 5796 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0822_
timestamp 1730882523
transform 1 0 6256 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0823_
timestamp 1730882523
transform 1 0 6716 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0824_
timestamp 1730882523
transform 1 0 8004 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0825_
timestamp 1730882523
transform -1 0 8096 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _0826_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 6992 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0827_
timestamp 1730882523
transform 1 0 8924 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0828_
timestamp 1730882523
transform -1 0 8188 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0829_
timestamp 1730882523
transform -1 0 8372 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0830_
timestamp 1730882523
transform 1 0 7544 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0831_
timestamp 1730882523
transform -1 0 11408 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0832_
timestamp 1730882523
transform -1 0 10580 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0833_
timestamp 1730882523
transform -1 0 11132 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0834_
timestamp 1730882523
transform -1 0 10120 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0835_
timestamp 1730882523
transform -1 0 8832 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0836_
timestamp 1730882523
transform 1 0 8924 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0837_
timestamp 1730882523
transform -1 0 10764 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0838_
timestamp 1730882523
transform -1 0 11316 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _0839_
timestamp 1730882523
transform 1 0 9384 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _0840_
timestamp 1730882523
transform 1 0 9200 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0841_
timestamp 1730882523
transform 1 0 6164 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0842_
timestamp 1730882523
transform 1 0 8740 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _0843_
timestamp 1730882523
transform 1 0 8924 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _0844_
timestamp 1730882523
transform 1 0 7452 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__o311a_1  _0845_
timestamp 1730882523
transform 1 0 6716 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0846_
timestamp 1730882523
transform 1 0 5428 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _0847_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform -1 0 7176 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0848_
timestamp 1730882523
transform 1 0 6716 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0849_
timestamp 1730882523
transform 1 0 9660 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0850_
timestamp 1730882523
transform 1 0 8004 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0851_
timestamp 1730882523
transform 1 0 12420 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0852_
timestamp 1730882523
transform 1 0 10120 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0853_
timestamp 1730882523
transform 1 0 10396 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0854_
timestamp 1730882523
transform 1 0 9568 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0855_
timestamp 1730882523
transform -1 0 12328 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0856_
timestamp 1730882523
transform 1 0 12328 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0857_
timestamp 1730882523
transform 1 0 10120 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0858_
timestamp 1730882523
transform 1 0 9016 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0859_
timestamp 1730882523
transform 1 0 11500 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0860_
timestamp 1730882523
transform 1 0 11132 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0861_
timestamp 1730882523
transform 1 0 10580 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0862_
timestamp 1730882523
transform 1 0 10120 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0863_
timestamp 1730882523
transform 1 0 9108 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0864_
timestamp 1730882523
transform 1 0 8280 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0865_
timestamp 1730882523
transform 1 0 5796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0866_
timestamp 1730882523
transform -1 0 8096 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0867_
timestamp 1730882523
transform 1 0 6348 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0868_
timestamp 1730882523
transform -1 0 6808 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _0869_
timestamp 1730882523
transform 1 0 5244 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0870_
timestamp 1730882523
transform 1 0 6256 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0871_
timestamp 1730882523
transform 1 0 5244 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _0872_
timestamp 1730882523
transform 1 0 5060 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0873_
timestamp 1730882523
transform 1 0 5796 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0874_
timestamp 1730882523
transform 1 0 5888 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0875_
timestamp 1730882523
transform 1 0 4140 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0876_
timestamp 1730882523
transform -1 0 6992 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o41ai_1  _0877_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform -1 0 6992 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _0878_
timestamp 1730882523
transform 1 0 6808 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _0879_
timestamp 1730882523
transform 1 0 6716 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0880_
timestamp 1730882523
transform -1 0 5980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0881_
timestamp 1730882523
transform -1 0 7544 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0882_
timestamp 1730882523
transform -1 0 7452 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _0883_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 4416 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0884_
timestamp 1730882523
transform 1 0 4784 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0885_
timestamp 1730882523
transform -1 0 6440 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0886_
timestamp 1730882523
transform 1 0 6440 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0887_
timestamp 1730882523
transform -1 0 5796 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0888_
timestamp 1730882523
transform 1 0 4600 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0889_
timestamp 1730882523
transform 1 0 5520 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0890_
timestamp 1730882523
transform -1 0 6808 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0891_
timestamp 1730882523
transform -1 0 5704 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0892_
timestamp 1730882523
transform 1 0 5612 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0893_
timestamp 1730882523
transform -1 0 5612 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0894_
timestamp 1730882523
transform 1 0 4140 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0895_
timestamp 1730882523
transform -1 0 5336 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0896_
timestamp 1730882523
transform 1 0 4416 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0897_
timestamp 1730882523
transform 1 0 4968 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0898_
timestamp 1730882523
transform -1 0 5888 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0899_
timestamp 1730882523
transform 1 0 5152 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0900_
timestamp 1730882523
transform 1 0 4968 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0901_
timestamp 1730882523
transform -1 0 6164 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0902_
timestamp 1730882523
transform 1 0 5428 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0903_
timestamp 1730882523
transform 1 0 5336 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0904_
timestamp 1730882523
transform 1 0 7268 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0905_
timestamp 1730882523
transform 1 0 6624 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0906_
timestamp 1730882523
transform 1 0 5980 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0907_
timestamp 1730882523
transform 1 0 8280 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0908_
timestamp 1730882523
transform 1 0 6900 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_1  _0909_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform -1 0 8648 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0910_
timestamp 1730882523
transform 1 0 8372 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0911_
timestamp 1730882523
transform -1 0 7728 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0912_
timestamp 1730882523
transform -1 0 8556 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0913_
timestamp 1730882523
transform 1 0 8096 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0914_
timestamp 1730882523
transform 1 0 9108 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0915_
timestamp 1730882523
transform 1 0 8924 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0916_
timestamp 1730882523
transform -1 0 8740 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _0917_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 8004 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0918_
timestamp 1730882523
transform -1 0 9200 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0919_
timestamp 1730882523
transform -1 0 7268 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0920_
timestamp 1730882523
transform -1 0 7268 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0921_
timestamp 1730882523
transform 1 0 8740 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0922_
timestamp 1730882523
transform -1 0 6164 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0923_
timestamp 1730882523
transform 1 0 6716 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0924_
timestamp 1730882523
transform 1 0 6532 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0925_
timestamp 1730882523
transform 1 0 5704 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0926_
timestamp 1730882523
transform -1 0 2208 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0927_
timestamp 1730882523
transform -1 0 3680 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0928_
timestamp 1730882523
transform -1 0 3956 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0929_
timestamp 1730882523
transform 1 0 3036 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0930_
timestamp 1730882523
transform -1 0 2668 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0931_
timestamp 1730882523
transform -1 0 4876 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0932_
timestamp 1730882523
transform -1 0 2760 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0933_
timestamp 1730882523
transform -1 0 2300 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0934_
timestamp 1730882523
transform -1 0 3496 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0935_
timestamp 1730882523
transform 1 0 2300 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0936_
timestamp 1730882523
transform -1 0 2208 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0937_
timestamp 1730882523
transform -1 0 1840 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0938_
timestamp 1730882523
transform -1 0 2116 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0939_
timestamp 1730882523
transform -1 0 2668 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0940_
timestamp 1730882523
transform -1 0 2208 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0941_
timestamp 1730882523
transform 1 0 1840 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0942_
timestamp 1730882523
transform 1 0 1472 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0943_
timestamp 1730882523
transform 1 0 2852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0944_
timestamp 1730882523
transform -1 0 3312 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0945_
timestamp 1730882523
transform -1 0 2944 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0946_
timestamp 1730882523
transform 1 0 4416 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0947_
timestamp 1730882523
transform -1 0 2760 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0948_
timestamp 1730882523
transform -1 0 2116 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0949_
timestamp 1730882523
transform 1 0 1472 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0950_
timestamp 1730882523
transform 1 0 2116 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0951_
timestamp 1730882523
transform 1 0 2852 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0952_
timestamp 1730882523
transform -1 0 2576 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0953_
timestamp 1730882523
transform -1 0 1656 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0954_
timestamp 1730882523
transform -1 0 2208 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0955_
timestamp 1730882523
transform -1 0 3680 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0956_
timestamp 1730882523
transform 1 0 3312 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0957_
timestamp 1730882523
transform 1 0 4140 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0958_
timestamp 1730882523
transform -1 0 3588 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0959_
timestamp 1730882523
transform 1 0 2576 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0960_
timestamp 1730882523
transform -1 0 5152 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0961_
timestamp 1730882523
transform -1 0 4140 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0962_
timestamp 1730882523
transform 1 0 3220 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0963_
timestamp 1730882523
transform 1 0 5244 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0964_
timestamp 1730882523
transform 1 0 2760 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0965_
timestamp 1730882523
transform -1 0 4416 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0966_
timestamp 1730882523
transform 1 0 10672 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0967_
timestamp 1730882523
transform -1 0 11408 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0968_
timestamp 1730882523
transform 1 0 11132 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0969_
timestamp 1730882523
transform 1 0 12328 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0970_
timestamp 1730882523
transform 1 0 10764 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0971_
timestamp 1730882523
transform 1 0 10396 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _0972_
timestamp 1730882523
transform 1 0 9292 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0973_
timestamp 1730882523
transform 1 0 10396 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0974_
timestamp 1730882523
transform -1 0 10396 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0975_
timestamp 1730882523
transform 1 0 10580 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0976_
timestamp 1730882523
transform 1 0 9660 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0977_
timestamp 1730882523
transform 1 0 10856 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0978_
timestamp 1730882523
transform 1 0 10948 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0979_
timestamp 1730882523
transform 1 0 10580 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0980_
timestamp 1730882523
transform -1 0 11592 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _0981_
timestamp 1730882523
transform 1 0 9752 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0982_
timestamp 1730882523
transform 1 0 9752 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0983_
timestamp 1730882523
transform 1 0 10488 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0984_
timestamp 1730882523
transform -1 0 13892 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0985_
timestamp 1730882523
transform -1 0 12052 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0986_
timestamp 1730882523
transform -1 0 12144 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0987_
timestamp 1730882523
transform 1 0 10212 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0988_
timestamp 1730882523
transform -1 0 11776 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0989_
timestamp 1730882523
transform -1 0 10856 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0990_
timestamp 1730882523
transform 1 0 10672 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0991_
timestamp 1730882523
transform -1 0 11868 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0992_
timestamp 1730882523
transform -1 0 10948 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0993_
timestamp 1730882523
transform 1 0 11960 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0994_
timestamp 1730882523
transform 1 0 11316 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _0995_
timestamp 1730882523
transform -1 0 10580 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0996_
timestamp 1730882523
transform 1 0 11316 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0997_
timestamp 1730882523
transform -1 0 11960 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0998_
timestamp 1730882523
transform 1 0 10580 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _0999_
timestamp 1730882523
transform -1 0 10580 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _1000_
timestamp 1730882523
transform -1 0 9660 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1001_
timestamp 1730882523
transform -1 0 9016 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1002_
timestamp 1730882523
transform -1 0 10948 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1003_
timestamp 1730882523
transform 1 0 12604 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1004_
timestamp 1730882523
transform 1 0 11960 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1005_
timestamp 1730882523
transform 1 0 12420 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1006_
timestamp 1730882523
transform 1 0 10948 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1007_
timestamp 1730882523
transform -1 0 11408 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1008_
timestamp 1730882523
transform -1 0 13984 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1009_
timestamp 1730882523
transform 1 0 12236 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _1010_
timestamp 1730882523
transform 1 0 10948 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1011_
timestamp 1730882523
transform -1 0 12420 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1012_
timestamp 1730882523
transform 1 0 9844 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1013_
timestamp 1730882523
transform 1 0 12512 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1014_
timestamp 1730882523
transform 1 0 12972 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__a2bb2o_1  _1015_
timestamp 1730882523
transform -1 0 11776 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a21boi_1  _1016_
timestamp 1730882523
transform -1 0 12328 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1017_
timestamp 1730882523
transform 1 0 11776 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1018_
timestamp 1730882523
transform 1 0 11868 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1019_
timestamp 1730882523
transform 1 0 12512 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1020_
timestamp 1730882523
transform 1 0 9568 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1021_
timestamp 1730882523
transform 1 0 10488 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _1022_
timestamp 1730882523
transform 1 0 9384 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1023_
timestamp 1730882523
transform 1 0 9292 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1024_
timestamp 1730882523
transform -1 0 10488 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1025_
timestamp 1730882523
transform 1 0 9200 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1026_
timestamp 1730882523
transform 1 0 8648 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1027_
timestamp 1730882523
transform 1 0 8924 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1028_
timestamp 1730882523
transform 1 0 8924 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_1  _1029_
timestamp 1730882523
transform 1 0 9660 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1030_
timestamp 1730882523
transform 1 0 9476 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1031_
timestamp 1730882523
transform 1 0 9752 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1032_
timestamp 1730882523
transform 1 0 10488 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1033_
timestamp 1730882523
transform -1 0 10672 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1034_
timestamp 1730882523
transform 1 0 9292 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1035_
timestamp 1730882523
transform -1 0 8924 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1036_
timestamp 1730882523
transform -1 0 8464 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1037_
timestamp 1730882523
transform 1 0 9292 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1038_
timestamp 1730882523
transform 1 0 8924 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _1039_
timestamp 1730882523
transform -1 0 8280 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1040_
timestamp 1730882523
transform 1 0 13432 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1041_
timestamp 1730882523
transform 1 0 11684 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _1042_
timestamp 1730882523
transform -1 0 13708 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1043_
timestamp 1730882523
transform 1 0 11500 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and4b_1  _1044_
timestamp 1730882523
transform -1 0 9660 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1045_
timestamp 1730882523
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1046_
timestamp 1730882523
transform 1 0 7268 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_1  _1047_
timestamp 1730882523
transform 1 0 8280 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1048_
timestamp 1730882523
transform 1 0 10396 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _1049_
timestamp 1730882523
transform 1 0 10764 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1050_
timestamp 1730882523
transform 1 0 11408 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1051_
timestamp 1730882523
transform 1 0 6348 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1052_
timestamp 1730882523
transform -1 0 8188 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1053_
timestamp 1730882523
transform 1 0 11500 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1054_
timestamp 1730882523
transform 1 0 12420 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1055_
timestamp 1730882523
transform -1 0 12696 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1056_
timestamp 1730882523
transform 1 0 12696 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1057_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 11408 0 1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1058_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 11776 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1059_
timestamp 1730882523
transform 1 0 1380 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1060_
timestamp 1730882523
transform 1 0 1472 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1061_
timestamp 1730882523
transform 1 0 1380 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1062_
timestamp 1730882523
transform 1 0 1472 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1063_
timestamp 1730882523
transform 1 0 2024 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1064_
timestamp 1730882523
transform 1 0 2760 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1065_
timestamp 1730882523
transform 1 0 3220 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1066_
timestamp 1730882523
transform 1 0 4048 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1067_
timestamp 1730882523
transform 1 0 4692 0 -1 27200
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1068_
timestamp 1730882523
transform 1 0 4784 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1069_
timestamp 1730882523
transform -1 0 6532 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1070_
timestamp 1730882523
transform -1 0 7820 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1071_
timestamp 1730882523
transform 1 0 5336 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1072_
timestamp 1730882523
transform 1 0 8004 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1073_
timestamp 1730882523
transform -1 0 8004 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1074_
timestamp 1730882523
transform 1 0 14076 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1075_
timestamp 1730882523
transform 1 0 14076 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1076_
timestamp 1730882523
transform -1 0 13616 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1077_
timestamp 1730882523
transform 1 0 13432 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1078_
timestamp 1730882523
transform 1 0 13156 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1079_
timestamp 1730882523
transform 1 0 14076 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1080_
timestamp 1730882523
transform -1 0 13892 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1081_
timestamp 1730882523
transform -1 0 14904 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1082_
timestamp 1730882523
transform 1 0 14904 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1083_
timestamp 1730882523
transform 1 0 14904 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1084_
timestamp 1730882523
transform 1 0 14904 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1085_
timestamp 1730882523
transform 1 0 14904 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1086_
timestamp 1730882523
transform 1 0 14904 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1087_
timestamp 1730882523
transform 1 0 14904 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1088_
timestamp 1730882523
transform 1 0 14904 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1089_
timestamp 1730882523
transform 1 0 14812 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1090_
timestamp 1730882523
transform 1 0 14904 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1091_
timestamp 1730882523
transform 1 0 14904 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1092_
timestamp 1730882523
transform 1 0 14076 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1093_
timestamp 1730882523
transform 1 0 14904 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1094_
timestamp 1730882523
transform -1 0 16100 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1095_
timestamp 1730882523
transform 1 0 14904 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1096_
timestamp 1730882523
transform -1 0 15548 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1097_
timestamp 1730882523
transform -1 0 16008 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1098_
timestamp 1730882523
transform 1 0 14904 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1099_
timestamp 1730882523
transform 1 0 14904 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1100_
timestamp 1730882523
transform 1 0 13064 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1101_
timestamp 1730882523
transform 1 0 14904 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1102_
timestamp 1730882523
transform 1 0 12696 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1103_
timestamp 1730882523
transform 1 0 14904 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1104_
timestamp 1730882523
transform 1 0 13064 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1105_
timestamp 1730882523
transform 1 0 13064 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1106_
timestamp 1730882523
transform 1 0 14444 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1107_
timestamp 1730882523
transform 1 0 14904 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1108_
timestamp 1730882523
transform 1 0 13524 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1109_
timestamp 1730882523
transform 1 0 14536 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1110_
timestamp 1730882523
transform 1 0 14904 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1111_
timestamp 1730882523
transform 1 0 14444 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1112_
timestamp 1730882523
transform 1 0 14076 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1113_
timestamp 1730882523
transform 1 0 13892 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1114_
timestamp 1730882523
transform 1 0 6900 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1115_
timestamp 1730882523
transform -1 0 13616 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1116_
timestamp 1730882523
transform -1 0 12972 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1117_
timestamp 1730882523
transform -1 0 12972 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1118_
timestamp 1730882523
transform -1 0 13432 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1119_
timestamp 1730882523
transform -1 0 13248 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1120_
timestamp 1730882523
transform -1 0 11408 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1121_
timestamp 1730882523
transform 1 0 10948 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1122_
timestamp 1730882523
transform -1 0 13340 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1123_
timestamp 1730882523
transform 1 0 11960 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1124_
timestamp 1730882523
transform 1 0 12052 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1125_
timestamp 1730882523
transform 1 0 12236 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1126_
timestamp 1730882523
transform -1 0 13064 0 -1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1127_
timestamp 1730882523
transform 1 0 11500 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1128_
timestamp 1730882523
transform 1 0 5520 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1129_
timestamp 1730882523
transform 1 0 6348 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1130_
timestamp 1730882523
transform 1 0 6440 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1131_
timestamp 1730882523
transform 1 0 6532 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1132_
timestamp 1730882523
transform 1 0 6808 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1133_
timestamp 1730882523
transform 1 0 8004 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1134_
timestamp 1730882523
transform 1 0 9660 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1135_
timestamp 1730882523
transform 1 0 8924 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1136_
timestamp 1730882523
transform 1 0 9568 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1137_
timestamp 1730882523
transform 1 0 8188 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1138_
timestamp 1730882523
transform 1 0 9660 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1139_
timestamp 1730882523
transform 1 0 9476 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1140_
timestamp 1730882523
transform -1 0 8832 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1141_
timestamp 1730882523
transform 1 0 5244 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1142_
timestamp 1730882523
transform 1 0 6348 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1143_
timestamp 1730882523
transform 1 0 5520 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1144_
timestamp 1730882523
transform 1 0 4784 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1145_
timestamp 1730882523
transform -1 0 6716 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1146_
timestamp 1730882523
transform 1 0 4784 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1147_
timestamp 1730882523
transform -1 0 6072 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1148_
timestamp 1730882523
transform 1 0 5244 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1149_
timestamp 1730882523
transform -1 0 8188 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1150_
timestamp 1730882523
transform -1 0 8096 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1151_
timestamp 1730882523
transform 1 0 6808 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1152_
timestamp 1730882523
transform -1 0 8096 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1153_
timestamp 1730882523
transform 1 0 8924 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1154_
timestamp 1730882523
transform 1 0 6900 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1155_
timestamp 1730882523
transform 1 0 6900 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1156_
timestamp 1730882523
transform -1 0 8372 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1157_
timestamp 1730882523
transform 1 0 8188 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1158_
timestamp 1730882523
transform 1 0 7912 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1159_
timestamp 1730882523
transform -1 0 8740 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1160_
timestamp 1730882523
transform 1 0 6348 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1161_
timestamp 1730882523
transform -1 0 7544 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1162_
timestamp 1730882523
transform 1 0 8372 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1163_
timestamp 1730882523
transform 1 0 9016 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1164_
timestamp 1730882523
transform 1 0 1380 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1165_
timestamp 1730882523
transform 1 0 3404 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1166_
timestamp 1730882523
transform 1 0 1564 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1167_
timestamp 1730882523
transform 1 0 1380 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1168_
timestamp 1730882523
transform 1 0 1380 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1169_
timestamp 1730882523
transform -1 0 2852 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1170_
timestamp 1730882523
transform 1 0 1380 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1171_
timestamp 1730882523
transform -1 0 2852 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1172_
timestamp 1730882523
transform 1 0 1564 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1173_
timestamp 1730882523
transform 1 0 1656 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1174_
timestamp 1730882523
transform -1 0 5244 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1175_
timestamp 1730882523
transform 1 0 3220 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1176_
timestamp 1730882523
transform 1 0 3772 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1177_
timestamp 1730882523
transform 1 0 11960 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1178_
timestamp 1730882523
transform 1 0 9844 0 -1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1179_
timestamp 1730882523
transform 1 0 8372 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1180_
timestamp 1730882523
transform 1 0 9476 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1181_
timestamp 1730882523
transform 1 0 9936 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1182_
timestamp 1730882523
transform 1 0 9200 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1183_
timestamp 1730882523
transform 1 0 11500 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1184_
timestamp 1730882523
transform -1 0 11500 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1185_
timestamp 1730882523
transform 1 0 10396 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1186_
timestamp 1730882523
transform 1 0 11960 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1187_
timestamp 1730882523
transform 1 0 11868 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1188_
timestamp 1730882523
transform 1 0 12328 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1189_
timestamp 1730882523
transform 1 0 12236 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1190_
timestamp 1730882523
transform 1 0 6440 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1191_
timestamp 1730882523
transform 1 0 7820 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1192_
timestamp 1730882523
transform 1 0 8004 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1193_
timestamp 1730882523
transform 1 0 8188 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1194_
timestamp 1730882523
transform 1 0 9016 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1195_
timestamp 1730882523
transform -1 0 10948 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1196_
timestamp 1730882523
transform 1 0 9752 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1197_
timestamp 1730882523
transform 1 0 9844 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1198_
timestamp 1730882523
transform 1 0 6900 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1199_
timestamp 1730882523
transform 1 0 6900 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1200_
timestamp 1730882523
transform 1 0 11500 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1201_
timestamp 1730882523
transform 1 0 11500 0 -1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1202_
timestamp 1730882523
transform 1 0 7084 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1203_
timestamp 1730882523
transform -1 0 8372 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1204_
timestamp 1730882523
transform 1 0 9752 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1205_
timestamp 1730882523
transform 1 0 11132 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1206_
timestamp 1730882523
transform 1 0 6900 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1207_
timestamp 1730882523
transform 1 0 12328 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _1208_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform -1 0 14444 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1209_
timestamp 1730882523
transform -1 0 14352 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1210_
timestamp 1730882523
transform 1 0 14628 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1211_
timestamp 1730882523
transform 1 0 13708 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1212_
timestamp 1730882523
transform -1 0 15548 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1213_
timestamp 1730882523
transform -1 0 15548 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1214_
timestamp 1730882523
transform -1 0 14536 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1215_
timestamp 1730882523
transform 1 0 8556 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 8924 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_clk ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform -1 0 5244 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_clk
timestamp 1730882523
transform -1 0 6900 0 1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_clk
timestamp 1730882523
transform 1 0 4600 0 1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_clk
timestamp 1730882523
transform 1 0 6992 0 -1 14144
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_clk
timestamp 1730882523
transform -1 0 11408 0 1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_clk
timestamp 1730882523
transform -1 0 13432 0 1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_clk
timestamp 1730882523
transform 1 0 11684 0 1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_clk
timestamp 1730882523
transform 1 0 14076 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_clk
timestamp 1730882523
transform 1 0 5612 0 1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_clk
timestamp 1730882523
transform 1 0 8188 0 -1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_clk
timestamp 1730882523
transform -1 0 6532 0 1 25024
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_clk
timestamp 1730882523
transform 1 0 7176 0 -1 26112
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_clk
timestamp 1730882523
transform 1 0 10948 0 1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_clk
timestamp 1730882523
transform 1 0 14076 0 1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_clk
timestamp 1730882523
transform -1 0 12512 0 -1 27200
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_clk
timestamp 1730882523
transform 1 0 13248 0 -1 26112
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_8  clkload0 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform -1 0 5520 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkinv_4  clkload1 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 5244 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__inv_6  clkload2 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 4600 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  clkload3
timestamp 1730882523
transform 1 0 7360 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__clkinvlp_4  clkload4 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 9844 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__inv_6  clkload5
timestamp 1730882523
transform 1 0 11684 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__clkinvlp_4  clkload6
timestamp 1730882523
transform 1 0 13432 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__inv_8  clkload7
timestamp 1730882523
transform 1 0 4784 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__inv_6  clkload8
timestamp 1730882523
transform 1 0 8924 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  clkload9
timestamp 1730882523
transform 1 0 5520 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_2  clkload10 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 7268 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__inv_6  clkload11
timestamp 1730882523
transform 1 0 11500 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__clkinvlp_4  clkload12
timestamp 1730882523
transform 1 0 13432 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkinvlp_4  clkload13
timestamp 1730882523
transform 1 0 10948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout58 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 3864 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout59
timestamp 1730882523
transform -1 0 6716 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout60
timestamp 1730882523
transform 1 0 3312 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout61
timestamp 1730882523
transform 1 0 2116 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout63
timestamp 1730882523
transform -1 0 6716 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout64 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 10856 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout65 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 9844 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout66
timestamp 1730882523
transform 1 0 9108 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout69
timestamp 1730882523
transform -1 0 9384 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout70
timestamp 1730882523
transform -1 0 3680 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout71 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform -1 0 8464 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  fanout72
timestamp 1730882523
transform -1 0 13524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout73
timestamp 1730882523
transform -1 0 4968 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout74 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 4508 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout75
timestamp 1730882523
transform -1 0 12972 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout76
timestamp 1730882523
transform -1 0 14168 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout77
timestamp 1730882523
transform -1 0 16376 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout78
timestamp 1730882523
transform -1 0 10672 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout79
timestamp 1730882523
transform -1 0 11040 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout80
timestamp 1730882523
transform -1 0 11316 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout81
timestamp 1730882523
transform 1 0 4048 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout82
timestamp 1730882523
transform 1 0 3496 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout83
timestamp 1730882523
transform 1 0 2392 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1730882523
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1730882523
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1730882523
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 6348 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65
timestamp 1730882523
transform 1 0 7084 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_91
timestamp 1730882523
transform 1 0 9476 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98
timestamp 1730882523
transform 1 0 10120 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1730882523
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1730882523
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_125 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 12604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_133
timestamp 1730882523
transform 1 0 13340 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1730882523
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_160
timestamp 1730882523
transform 1 0 15824 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1730882523
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1730882523
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1730882523
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1730882523
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1730882523
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1730882523
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1730882523
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_69 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 7452 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_91
timestamp 1730882523
transform 1 0 9476 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_99
timestamp 1730882523
transform 1 0 10212 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1730882523
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1730882523
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_125
timestamp 1730882523
transform 1 0 12604 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1730882523
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1730882523
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1730882523
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1730882523
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1730882523
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1730882523
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1730882523
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_77
timestamp 1730882523
transform 1 0 8188 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_85
timestamp 1730882523
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_116
timestamp 1730882523
transform 1 0 11776 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1730882523
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_149
timestamp 1730882523
transform 1 0 14812 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1730882523
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1730882523
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1730882523
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1730882523
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1730882523
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1730882523
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1730882523
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_69
timestamp 1730882523
transform 1 0 7452 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_93
timestamp 1730882523
transform 1 0 9660 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_146
timestamp 1730882523
transform 1 0 14536 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_163
timestamp 1730882523
transform 1 0 16100 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1730882523
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1730882523
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1730882523
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1730882523
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1730882523
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1730882523
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1730882523
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1730882523
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1730882523
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_110
timestamp 1730882523
transform 1 0 11224 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp 1730882523
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_165
timestamp 1730882523
transform 1 0 16284 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1730882523
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1730882523
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1730882523
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1730882523
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1730882523
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1730882523
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1730882523
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1730882523
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1730882523
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_93
timestamp 1730882523
transform 1 0 9660 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_104
timestamp 1730882523
transform 1 0 10672 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_113
timestamp 1730882523
transform 1 0 11500 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_164
timestamp 1730882523
transform 1 0 16192 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1730882523
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1730882523
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1730882523
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_61
timestamp 1730882523
transform 1 0 6716 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_73
timestamp 1730882523
transform 1 0 7820 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_81
timestamp 1730882523
transform 1 0 8556 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1730882523
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_97
timestamp 1730882523
transform 1 0 10028 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_101
timestamp 1730882523
transform 1 0 10396 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_108
timestamp 1730882523
transform 1 0 11040 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_114
timestamp 1730882523
transform 1 0 11592 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_155
timestamp 1730882523
transform 1 0 15364 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_164
timestamp 1730882523
transform 1 0 16192 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1730882523
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_15
timestamp 1730882523
transform 1 0 2484 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_44
timestamp 1730882523
transform 1 0 5152 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_53
timestamp 1730882523
transform 1 0 5980 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_63
timestamp 1730882523
transform 1 0 6900 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_75
timestamp 1730882523
transform 1 0 8004 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_87
timestamp 1730882523
transform 1 0 9108 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_98
timestamp 1730882523
transform 1 0 10120 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_120
timestamp 1730882523
transform 1 0 12144 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_140
timestamp 1730882523
transform 1 0 13984 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_165
timestamp 1730882523
transform 1 0 16284 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3
timestamp 1730882523
transform 1 0 1380 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_16
timestamp 1730882523
transform 1 0 2576 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_69
timestamp 1730882523
transform 1 0 7452 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_76
timestamp 1730882523
transform 1 0 8096 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_85
timestamp 1730882523
transform 1 0 8924 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_112
timestamp 1730882523
transform 1 0 11408 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_122
timestamp 1730882523
transform 1 0 12328 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_137
timestamp 1730882523
transform 1 0 13708 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_148
timestamp 1730882523
transform 1 0 14720 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_27
timestamp 1730882523
transform 1 0 3588 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_84
timestamp 1730882523
transform 1 0 8832 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 1730882523
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1730882523
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_36
timestamp 1730882523
transform 1 0 4416 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_70
timestamp 1730882523
transform 1 0 7544 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_90
timestamp 1730882523
transform 1 0 9384 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_137
timestamp 1730882523
transform 1 0 13708 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_149
timestamp 1730882523
transform 1 0 14812 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_27
timestamp 1730882523
transform 1 0 3588 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_52
timestamp 1730882523
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_62
timestamp 1730882523
transform 1 0 6808 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1730882523
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1730882523
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_141
timestamp 1730882523
transform 1 0 14076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_3
timestamp 1730882523
transform 1 0 1380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_16
timestamp 1730882523
transform 1 0 2576 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_22
timestamp 1730882523
transform 1 0 3128 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_35
timestamp 1730882523
transform 1 0 4324 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_44
timestamp 1730882523
transform 1 0 5152 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_121
timestamp 1730882523
transform 1 0 12236 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1730882523
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_146
timestamp 1730882523
transform 1 0 14536 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1730882523
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_15
timestamp 1730882523
transform 1 0 2484 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_37
timestamp 1730882523
transform 1 0 4508 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1730882523
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_62
timestamp 1730882523
transform 1 0 6808 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_93
timestamp 1730882523
transform 1 0 9660 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1730882523
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_153
timestamp 1730882523
transform 1 0 15180 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_165
timestamp 1730882523
transform 1 0 16284 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1730882523
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_15
timestamp 1730882523
transform 1 0 2484 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_21
timestamp 1730882523
transform 1 0 3036 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_29
timestamp 1730882523
transform 1 0 3772 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_80
timestamp 1730882523
transform 1 0 8464 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_93
timestamp 1730882523
transform 1 0 9660 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_103
timestamp 1730882523
transform 1 0 10580 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_14_125
timestamp 1730882523
transform 1 0 12604 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_3
timestamp 1730882523
transform 1 0 1380 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_18
timestamp 1730882523
transform 1 0 2760 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_30
timestamp 1730882523
transform 1 0 3864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_53
timestamp 1730882523
transform 1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_57
timestamp 1730882523
transform 1 0 6348 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_65
timestamp 1730882523
transform 1 0 7084 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_72
timestamp 1730882523
transform 1 0 7728 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_81
timestamp 1730882523
transform 1 0 8556 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_94
timestamp 1730882523
transform 1 0 9752 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_106
timestamp 1730882523
transform 1 0 10856 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_113
timestamp 1730882523
transform 1 0 11500 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_122
timestamp 1730882523
transform 1 0 12328 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_130
timestamp 1730882523
transform 1 0 13064 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_22
timestamp 1730882523
transform 1 0 3128 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_16_29
timestamp 1730882523
transform 1 0 3772 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_41
timestamp 1730882523
transform 1 0 4876 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_50
timestamp 1730882523
transform 1 0 5704 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_62
timestamp 1730882523
transform 1 0 6808 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_74
timestamp 1730882523
transform 1 0 7912 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_78
timestamp 1730882523
transform 1 0 8280 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1730882523
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_109
timestamp 1730882523
transform 1 0 11132 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_126
timestamp 1730882523
transform 1 0 12696 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_141
timestamp 1730882523
transform 1 0 14076 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_28
timestamp 1730882523
transform 1 0 3680 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_39
timestamp 1730882523
transform 1 0 4692 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1730882523
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_57
timestamp 1730882523
transform 1 0 6348 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_68
timestamp 1730882523
transform 1 0 7360 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_72
timestamp 1730882523
transform 1 0 7728 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_113
timestamp 1730882523
transform 1 0 11500 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_149
timestamp 1730882523
transform 1 0 14812 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_3
timestamp 1730882523
transform 1 0 1380 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_20
timestamp 1730882523
transform 1 0 2944 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_29
timestamp 1730882523
transform 1 0 3772 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1730882523
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_113
timestamp 1730882523
transform 1 0 11500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_165
timestamp 1730882523
transform 1 0 16284 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1730882523
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_34
timestamp 1730882523
transform 1 0 4232 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_52
timestamp 1730882523
transform 1 0 5888 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_99
timestamp 1730882523
transform 1 0 10212 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1730882523
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_122
timestamp 1730882523
transform 1 0 12328 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_164
timestamp 1730882523
transform 1 0 16192 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_19
timestamp 1730882523
transform 1 0 2852 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_37
timestamp 1730882523
transform 1 0 4508 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_49
timestamp 1730882523
transform 1 0 5612 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_53
timestamp 1730882523
transform 1 0 5980 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_70
timestamp 1730882523
transform 1 0 7544 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_81
timestamp 1730882523
transform 1 0 8556 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_85
timestamp 1730882523
transform 1 0 8924 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_93
timestamp 1730882523
transform 1 0 9660 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_134
timestamp 1730882523
transform 1 0 13432 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_164
timestamp 1730882523
transform 1 0 16192 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_3
timestamp 1730882523
transform 1 0 1380 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_7
timestamp 1730882523
transform 1 0 1748 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_11
timestamp 1730882523
transform 1 0 2116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_23
timestamp 1730882523
transform 1 0 3220 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1730882523
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_91
timestamp 1730882523
transform 1 0 9476 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_99
timestamp 1730882523
transform 1 0 10212 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_121
timestamp 1730882523
transform 1 0 12236 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1730882523
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_15
timestamp 1730882523
transform 1 0 2484 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_23
timestamp 1730882523
transform 1 0 3220 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1730882523
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_29
timestamp 1730882523
transform 1 0 3772 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_33
timestamp 1730882523
transform 1 0 4140 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_57
timestamp 1730882523
transform 1 0 6348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_64
timestamp 1730882523
transform 1 0 6992 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_94
timestamp 1730882523
transform 1 0 9752 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_23_3
timestamp 1730882523
transform 1 0 1380 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_23_12
timestamp 1730882523
transform 1 0 2208 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_18
timestamp 1730882523
transform 1 0 2760 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_30
timestamp 1730882523
transform 1 0 3864 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_38
timestamp 1730882523
transform 1 0 4600 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_57
timestamp 1730882523
transform 1 0 6348 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_74
timestamp 1730882523
transform 1 0 7912 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_137
timestamp 1730882523
transform 1 0 13708 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_165
timestamp 1730882523
transform 1 0 16284 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1730882523
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_12
timestamp 1730882523
transform 1 0 2208 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_45
timestamp 1730882523
transform 1 0 5244 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1730882523
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_107
timestamp 1730882523
transform 1 0 10948 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_130
timestamp 1730882523
transform 1 0 13064 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1730882523
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_41
timestamp 1730882523
transform 1 0 4876 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1730882523
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_57
timestamp 1730882523
transform 1 0 6348 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_72
timestamp 1730882523
transform 1 0 7728 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_80
timestamp 1730882523
transform 1 0 8464 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_118
timestamp 1730882523
transform 1 0 11960 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_138
timestamp 1730882523
transform 1 0 13800 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_19
timestamp 1730882523
transform 1 0 2852 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1730882523
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1730882523
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_85
timestamp 1730882523
transform 1 0 8924 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_97
timestamp 1730882523
transform 1 0 10028 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_112
timestamp 1730882523
transform 1 0 11408 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_124
timestamp 1730882523
transform 1 0 12512 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_128
timestamp 1730882523
transform 1 0 12880 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_165
timestamp 1730882523
transform 1 0 16284 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1730882523
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_21
timestamp 1730882523
transform 1 0 3036 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_41
timestamp 1730882523
transform 1 0 4876 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1730882523
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1730882523
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_69
timestamp 1730882523
transform 1 0 7452 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_77
timestamp 1730882523
transform 1 0 8188 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_93
timestamp 1730882523
transform 1 0 9660 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1730882523
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1730882523
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_125
timestamp 1730882523
transform 1 0 12604 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_155
timestamp 1730882523
transform 1 0 15364 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_163
timestamp 1730882523
transform 1 0 16100 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_13
timestamp 1730882523
transform 1 0 2300 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_32
timestamp 1730882523
transform 1 0 4048 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_36
timestamp 1730882523
transform 1 0 4416 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_42
timestamp 1730882523
transform 1 0 4968 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_49
timestamp 1730882523
transform 1 0 5612 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_61
timestamp 1730882523
transform 1 0 6716 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1730882523
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_105
timestamp 1730882523
transform 1 0 10764 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_117
timestamp 1730882523
transform 1 0 11868 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_130
timestamp 1730882523
transform 1 0 13064 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_3
timestamp 1730882523
transform 1 0 1380 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_11
timestamp 1730882523
transform 1 0 2116 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_16
timestamp 1730882523
transform 1 0 2576 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_28
timestamp 1730882523
transform 1 0 3680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_52
timestamp 1730882523
transform 1 0 5888 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_63
timestamp 1730882523
transform 1 0 6900 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_87
timestamp 1730882523
transform 1 0 9108 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_104
timestamp 1730882523
transform 1 0 10672 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_113
timestamp 1730882523
transform 1 0 11500 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1730882523
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1730882523
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1730882523
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1730882523
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_41
timestamp 1730882523
transform 1 0 4876 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_49
timestamp 1730882523
transform 1 0 5612 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_105
timestamp 1730882523
transform 1 0 10764 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_119
timestamp 1730882523
transform 1 0 12052 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1730882523
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_165
timestamp 1730882523
transform 1 0 16284 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1730882523
transform 1 0 1380 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_20
timestamp 1730882523
transform 1 0 2944 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_26
timestamp 1730882523
transform 1 0 3496 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_36
timestamp 1730882523
transform 1 0 4416 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_53
timestamp 1730882523
transform 1 0 5980 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_57
timestamp 1730882523
transform 1 0 6348 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_102
timestamp 1730882523
transform 1 0 10488 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_116
timestamp 1730882523
transform 1 0 11776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_149
timestamp 1730882523
transform 1 0 14812 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_19
timestamp 1730882523
transform 1 0 2852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_29
timestamp 1730882523
transform 1 0 3772 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_62
timestamp 1730882523
transform 1 0 6808 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1730882523
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_89
timestamp 1730882523
transform 1 0 9292 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_98
timestamp 1730882523
transform 1 0 10120 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_106
timestamp 1730882523
transform 1 0 10856 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_122
timestamp 1730882523
transform 1 0 12328 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_134
timestamp 1730882523
transform 1 0 13432 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_157
timestamp 1730882523
transform 1 0 15548 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_165
timestamp 1730882523
transform 1 0 16284 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_3
timestamp 1730882523
transform 1 0 1380 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_27
timestamp 1730882523
transform 1 0 3588 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_37
timestamp 1730882523
transform 1 0 4508 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_73
timestamp 1730882523
transform 1 0 7820 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_92
timestamp 1730882523
transform 1 0 9568 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_100
timestamp 1730882523
transform 1 0 10304 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1730882523
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_116
timestamp 1730882523
transform 1 0 11776 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_124
timestamp 1730882523
transform 1 0 12512 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_165
timestamp 1730882523
transform 1 0 16284 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_3
timestamp 1730882523
transform 1 0 1380 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1730882523
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_47
timestamp 1730882523
transform 1 0 5428 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_79
timestamp 1730882523
transform 1 0 8372 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1730882523
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_92
timestamp 1730882523
transform 1 0 9568 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_135
timestamp 1730882523
transform 1 0 13524 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1730882523
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_141
timestamp 1730882523
transform 1 0 14076 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_34_147
timestamp 1730882523
transform 1 0 14628 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_6
timestamp 1730882523
transform 1 0 1656 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_18
timestamp 1730882523
transform 1 0 2760 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_22
timestamp 1730882523
transform 1 0 3128 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_61
timestamp 1730882523
transform 1 0 6716 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_74
timestamp 1730882523
transform 1 0 7912 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_35_88
timestamp 1730882523
transform 1 0 9200 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1730882523
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_15
timestamp 1730882523
transform 1 0 2484 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_36_29
timestamp 1730882523
transform 1 0 3772 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_39
timestamp 1730882523
transform 1 0 4692 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_79
timestamp 1730882523
transform 1 0 8372 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1730882523
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_101
timestamp 1730882523
transform 1 0 10396 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_125
timestamp 1730882523
transform 1 0 12604 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_156
timestamp 1730882523
transform 1 0 15456 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_3
timestamp 1730882523
transform 1 0 1380 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_18
timestamp 1730882523
transform 1 0 2760 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_26
timestamp 1730882523
transform 1 0 3496 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_61
timestamp 1730882523
transform 1 0 6716 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1730882523
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_165
timestamp 1730882523
transform 1 0 16284 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1730882523
transform 1 0 1380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_42
timestamp 1730882523
transform 1 0 4968 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_78
timestamp 1730882523
transform 1 0 8280 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_38_85
timestamp 1730882523
transform 1 0 8924 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_165
timestamp 1730882523
transform 1 0 16284 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_30
timestamp 1730882523
transform 1 0 3864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_38
timestamp 1730882523
transform 1 0 4600 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1730882523
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1730882523
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_81
timestamp 1730882523
transform 1 0 8556 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_87
timestamp 1730882523
transform 1 0 9108 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_164
timestamp 1730882523
transform 1 0 16192 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_3
timestamp 1730882523
transform 1 0 1380 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_85
timestamp 1730882523
transform 1 0 8924 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_91
timestamp 1730882523
transform 1 0 9476 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_117
timestamp 1730882523
transform 1 0 11868 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_134
timestamp 1730882523
transform 1 0 13432 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_164
timestamp 1730882523
transform 1 0 16192 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_3
timestamp 1730882523
transform 1 0 1380 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_14
timestamp 1730882523
transform 1 0 2392 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_41
timestamp 1730882523
transform 1 0 4876 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1730882523
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_60
timestamp 1730882523
transform 1 0 6624 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_93
timestamp 1730882523
transform 1 0 9660 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_6
timestamp 1730882523
transform 1 0 1656 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_18
timestamp 1730882523
transform 1 0 2760 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_26
timestamp 1730882523
transform 1 0 3496 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1730882523
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_41
timestamp 1730882523
transform 1 0 4876 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_47
timestamp 1730882523
transform 1 0 5428 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_59
timestamp 1730882523
transform 1 0 6532 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_66
timestamp 1730882523
transform 1 0 7176 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_85
timestamp 1730882523
transform 1 0 8924 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_103
timestamp 1730882523
transform 1 0 10580 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1730882523
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_148
timestamp 1730882523
transform 1 0 14720 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1730882523
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_15
timestamp 1730882523
transform 1 0 2484 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_21
timestamp 1730882523
transform 1 0 3036 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_43_41
timestamp 1730882523
transform 1 0 4876 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_43_52
timestamp 1730882523
transform 1 0 5888 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_43_57
timestamp 1730882523
transform 1 0 6348 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_43_102
timestamp 1730882523
transform 1 0 10488 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_43_113
timestamp 1730882523
transform 1 0 11500 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_164
timestamp 1730882523
transform 1 0 16192 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_3
timestamp 1730882523
transform 1 0 1380 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_44_29
timestamp 1730882523
transform 1 0 3772 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_55
timestamp 1730882523
transform 1 0 6164 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_133
timestamp 1730882523
transform 1 0 13340 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_165
timestamp 1730882523
transform 1 0 16284 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_45_3
timestamp 1730882523
transform 1 0 1380 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_73
timestamp 1730882523
transform 1 0 7820 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_45_91
timestamp 1730882523
transform 1 0 9476 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_45_109
timestamp 1730882523
transform 1 0 11132 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_45_133
timestamp 1730882523
transform 1 0 13340 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_3
timestamp 1730882523
transform 1 0 1380 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_9
timestamp 1730882523
transform 1 0 1932 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_26
timestamp 1730882523
transform 1 0 3496 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_72
timestamp 1730882523
transform 1 0 7728 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_88
timestamp 1730882523
transform 1 0 9200 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_108
timestamp 1730882523
transform 1 0 11040 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_46_165
timestamp 1730882523
transform 1 0 16284 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1730882523
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_15
timestamp 1730882523
transform 1 0 2484 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_37
timestamp 1730882523
transform 1 0 4508 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_49
timestamp 1730882523
transform 1 0 5612 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1730882523
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_57
timestamp 1730882523
transform 1 0 6348 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_47_80
timestamp 1730882523
transform 1 0 8464 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_47_92
timestamp 1730882523
transform 1 0 9568 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_100
timestamp 1730882523
transform 1 0 10304 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1730882523
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_15
timestamp 1730882523
transform 1 0 2484 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_23
timestamp 1730882523
transform 1 0 3220 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1730882523
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1730882523
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_53
timestamp 1730882523
transform 1 0 5980 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_67
timestamp 1730882523
transform 1 0 7268 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_48_78
timestamp 1730882523
transform 1 0 8280 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_90
timestamp 1730882523
transform 1 0 9384 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_113
timestamp 1730882523
transform 1 0 11500 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_138
timestamp 1730882523
transform 1 0 13800 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_149
timestamp 1730882523
transform 1 0 14812 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1730882523
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1730882523
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1730882523
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1730882523
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1730882523
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1730882523
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_57
timestamp 1730882523
transform 1 0 6348 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_49_66
timestamp 1730882523
transform 1 0 7176 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_89
timestamp 1730882523
transform 1 0 9292 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1730882523
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1730882523
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1730882523
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1730882523
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_41
timestamp 1730882523
transform 1 0 4876 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_49
timestamp 1730882523
transform 1 0 5612 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1730882523
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_50_134
timestamp 1730882523
transform 1 0 13432 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_50_165
timestamp 1730882523
transform 1 0 16284 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1730882523
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1730882523
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1730882523
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_39
timestamp 1730882523
transform 1 0 4692 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_73
timestamp 1730882523
transform 1 0 7820 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1730882523
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1730882523
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1730882523
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1730882523
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1730882523
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1730882523
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_53
timestamp 1730882523
transform 1 0 5980 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1730882523
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_52_149
timestamp 1730882523
transform 1 0 14812 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1730882523
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1730882523
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1730882523
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1730882523
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1730882523
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1730882523
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_57
timestamp 1730882523
transform 1 0 6348 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_53_109
timestamp 1730882523
transform 1 0 11132 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1730882523
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1730882523
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1730882523
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1730882523
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1730882523
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_53
timestamp 1730882523
transform 1 0 5980 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_57
timestamp 1730882523
transform 1 0 6348 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1730882523
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_118
timestamp 1730882523
transform 1 0 11960 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_54_157
timestamp 1730882523
transform 1 0 15548 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_54_165
timestamp 1730882523
transform 1 0 16284 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1730882523
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1730882523
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1730882523
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1730882523
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1730882523
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1730882523
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_57
timestamp 1730882523
transform 1 0 6348 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1730882523
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_81
timestamp 1730882523
transform 1 0 8556 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_88
timestamp 1730882523
transform 1 0 9200 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_121
timestamp 1730882523
transform 1 0 12236 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_139
timestamp 1730882523
transform 1 0 13892 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_164
timestamp 1730882523
transform 1 0 16192 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1730882523
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1730882523
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1730882523
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1730882523
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1730882523
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_53
timestamp 1730882523
transform 1 0 5980 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_57
timestamp 1730882523
transform 1 0 6348 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_69
timestamp 1730882523
transform 1 0 7452 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1730882523
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1730882523
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1730882523
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_97
timestamp 1730882523
transform 1 0 10028 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_56_156
timestamp 1730882523
transform 1 0 15456 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_164
timestamp 1730882523
transform 1 0 16192 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 6900 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1730882523
transform 1 0 7360 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1730882523
transform 1 0 10672 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1730882523
transform 1 0 9108 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1730882523
transform 1 0 9936 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1730882523
transform -1 0 13892 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1730882523
transform -1 0 13984 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1730882523
transform -1 0 14076 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1730882523
transform -1 0 10580 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1730882523
transform 1 0 10580 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1730882523
transform -1 0 14076 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1730882523
transform 1 0 11500 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1730882523
transform -1 0 15272 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1730882523
transform -1 0 13892 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1730882523
transform 1 0 13156 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1730882523
transform -1 0 13708 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1730882523
transform -1 0 8004 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1730882523
transform -1 0 12236 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1730882523
transform -1 0 12236 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1730882523
transform -1 0 14536 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1730882523
transform -1 0 8832 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1730882523
transform 1 0 10672 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1730882523
transform -1 0 10672 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1730882523
transform 1 0 12696 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1730882523
transform -1 0 11132 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1730882523
transform -1 0 15548 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1730882523
transform -1 0 14536 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1730882523
transform -1 0 10580 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1730882523
transform -1 0 14444 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1730882523
transform -1 0 14720 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1730882523
transform 1 0 11592 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1730882523
transform -1 0 14812 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1730882523
transform 1 0 11316 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1730882523
transform -1 0 7728 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1730882523
transform 1 0 6440 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 1730882523
transform 1 0 6072 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 1730882523
transform -1 0 8556 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 1730882523
transform -1 0 10580 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 1730882523
transform -1 0 7452 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 1730882523
transform -1 0 10212 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 1730882523
transform 1 0 6164 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 1730882523
transform -1 0 8832 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 1730882523
transform -1 0 9568 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 1730882523
transform -1 0 14812 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 1730882523
transform 1 0 8372 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 1730882523
transform -1 0 9660 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 1730882523
transform -1 0 8832 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 1730882523
transform -1 0 11224 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 1730882523
transform -1 0 8832 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 1730882523
transform 1 0 8004 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 1730882523
transform -1 0 14812 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 1730882523
transform -1 0 8280 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 1730882523
transform 1 0 10948 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 1730882523
transform -1 0 9660 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 1730882523
transform -1 0 14812 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold56
timestamp 1730882523
transform -1 0 13156 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp 1730882523
transform -1 0 9936 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1730882523
transform 1 0 1380 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1730882523
transform -1 0 1656 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input3
timestamp 1730882523
transform -1 0 16376 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1730882523
transform 1 0 8096 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5
timestamp 1730882523
transform 1 0 7176 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1730882523
transform -1 0 16376 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1730882523
transform 1 0 9752 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  max_cap67
timestamp 1730882523
transform -1 0 15180 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  max_cap68
timestamp 1730882523
transform -1 0 13984 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp 1730882523
transform 1 0 14628 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 1730882523
transform 1 0 14996 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1730882523
transform -1 0 10672 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 1730882523
transform -1 0 13340 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1730882523
transform 1 0 16008 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 1730882523
transform 1 0 16008 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 1730882523
transform 1 0 15180 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 1730882523
transform -1 0 8832 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 1730882523
transform -1 0 9476 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output17
timestamp 1730882523
transform -1 0 14076 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp 1730882523
transform 1 0 15088 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp 1730882523
transform -1 0 13984 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp 1730882523
transform -1 0 13892 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp 1730882523
transform -1 0 14168 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 1730882523
transform 1 0 16008 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 1730882523
transform -1 0 12236 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 1730882523
transform -1 0 13984 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 1730882523
transform 1 0 16008 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 1730882523
transform -1 0 12604 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 1730882523
transform -1 0 12236 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 1730882523
transform 1 0 14996 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 1730882523
transform -1 0 13984 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 1730882523
transform -1 0 11960 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 1730882523
transform -1 0 13340 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp 1730882523
transform -1 0 14628 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 1730882523
transform -1 0 13248 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 1730882523
transform 1 0 16008 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp 1730882523
transform -1 0 13524 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp 1730882523
transform 1 0 16008 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output37
timestamp 1730882523
transform -1 0 12696 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output38
timestamp 1730882523
transform -1 0 13892 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output39
timestamp 1730882523
transform 1 0 14536 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output40
timestamp 1730882523
transform -1 0 13064 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp 1730882523
transform -1 0 14444 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp 1730882523
transform 1 0 16008 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp 1730882523
transform -1 0 11500 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output44
timestamp 1730882523
transform 1 0 15640 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp 1730882523
transform -1 0 12420 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp 1730882523
transform -1 0 12880 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp 1730882523
transform -1 0 10120 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp 1730882523
transform -1 0 15456 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp 1730882523
transform -1 0 13984 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp 1730882523
transform -1 0 11316 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp 1730882523
transform 1 0 11500 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp 1730882523
transform 1 0 16008 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp 1730882523
transform -1 0 12512 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp 1730882523
transform -1 0 13708 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp 1730882523
transform -1 0 11408 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp 1730882523
transform 1 0 13616 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp 1730882523
transform -1 0 8188 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_57
timestamp 1730882523
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1730882523
transform -1 0 16652 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_58
timestamp 1730882523
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1730882523
transform -1 0 16652 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_59
timestamp 1730882523
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1730882523
transform -1 0 16652 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_60
timestamp 1730882523
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1730882523
transform -1 0 16652 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_61
timestamp 1730882523
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1730882523
transform -1 0 16652 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_62
timestamp 1730882523
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1730882523
transform -1 0 16652 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_63
timestamp 1730882523
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1730882523
transform -1 0 16652 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_64
timestamp 1730882523
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1730882523
transform -1 0 16652 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_65
timestamp 1730882523
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1730882523
transform -1 0 16652 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_66
timestamp 1730882523
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1730882523
transform -1 0 16652 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_67
timestamp 1730882523
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1730882523
transform -1 0 16652 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_68
timestamp 1730882523
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1730882523
transform -1 0 16652 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_69
timestamp 1730882523
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1730882523
transform -1 0 16652 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_70
timestamp 1730882523
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1730882523
transform -1 0 16652 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_71
timestamp 1730882523
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1730882523
transform -1 0 16652 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_72
timestamp 1730882523
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1730882523
transform -1 0 16652 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_73
timestamp 1730882523
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1730882523
transform -1 0 16652 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_74
timestamp 1730882523
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1730882523
transform -1 0 16652 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_75
timestamp 1730882523
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1730882523
transform -1 0 16652 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_76
timestamp 1730882523
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1730882523
transform -1 0 16652 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_77
timestamp 1730882523
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1730882523
transform -1 0 16652 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_78
timestamp 1730882523
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1730882523
transform -1 0 16652 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_79
timestamp 1730882523
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1730882523
transform -1 0 16652 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_80
timestamp 1730882523
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1730882523
transform -1 0 16652 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_81
timestamp 1730882523
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1730882523
transform -1 0 16652 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_82
timestamp 1730882523
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1730882523
transform -1 0 16652 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_83
timestamp 1730882523
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1730882523
transform -1 0 16652 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_84
timestamp 1730882523
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1730882523
transform -1 0 16652 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_85
timestamp 1730882523
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1730882523
transform -1 0 16652 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_86
timestamp 1730882523
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1730882523
transform -1 0 16652 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_87
timestamp 1730882523
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1730882523
transform -1 0 16652 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_88
timestamp 1730882523
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1730882523
transform -1 0 16652 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_89
timestamp 1730882523
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1730882523
transform -1 0 16652 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_90
timestamp 1730882523
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1730882523
transform -1 0 16652 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_91
timestamp 1730882523
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 1730882523
transform -1 0 16652 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_92
timestamp 1730882523
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 1730882523
transform -1 0 16652 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_93
timestamp 1730882523
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 1730882523
transform -1 0 16652 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_94
timestamp 1730882523
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 1730882523
transform -1 0 16652 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_95
timestamp 1730882523
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 1730882523
transform -1 0 16652 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_96
timestamp 1730882523
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp 1730882523
transform -1 0 16652 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_97
timestamp 1730882523
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp 1730882523
transform -1 0 16652 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_98
timestamp 1730882523
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp 1730882523
transform -1 0 16652 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Left_99
timestamp 1730882523
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Right_42
timestamp 1730882523
transform -1 0 16652 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Left_100
timestamp 1730882523
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Right_43
timestamp 1730882523
transform -1 0 16652 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Left_101
timestamp 1730882523
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Right_44
timestamp 1730882523
transform -1 0 16652 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Left_102
timestamp 1730882523
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Right_45
timestamp 1730882523
transform -1 0 16652 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Left_103
timestamp 1730882523
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Right_46
timestamp 1730882523
transform -1 0 16652 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Left_104
timestamp 1730882523
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Right_47
timestamp 1730882523
transform -1 0 16652 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Left_105
timestamp 1730882523
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Right_48
timestamp 1730882523
transform -1 0 16652 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Left_106
timestamp 1730882523
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Right_49
timestamp 1730882523
transform -1 0 16652 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Left_107
timestamp 1730882523
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Right_50
timestamp 1730882523
transform -1 0 16652 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Left_108
timestamp 1730882523
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Right_51
timestamp 1730882523
transform -1 0 16652 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Left_109
timestamp 1730882523
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Right_52
timestamp 1730882523
transform -1 0 16652 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Left_110
timestamp 1730882523
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Right_53
timestamp 1730882523
transform -1 0 16652 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Left_111
timestamp 1730882523
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Right_54
timestamp 1730882523
transform -1 0 16652 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Left_112
timestamp 1730882523
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Right_55
timestamp 1730882523
transform -1 0 16652 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Left_113
timestamp 1730882523
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Right_56
timestamp 1730882523
transform -1 0 16652 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_114 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_115
timestamp 1730882523
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_116
timestamp 1730882523
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_117
timestamp 1730882523
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_118
timestamp 1730882523
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_119
timestamp 1730882523
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_120
timestamp 1730882523
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_121
timestamp 1730882523
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_122
timestamp 1730882523
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_123
timestamp 1730882523
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_124
timestamp 1730882523
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_125
timestamp 1730882523
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_126
timestamp 1730882523
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_127
timestamp 1730882523
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_128
timestamp 1730882523
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_129
timestamp 1730882523
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_130
timestamp 1730882523
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_131
timestamp 1730882523
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_132
timestamp 1730882523
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_133
timestamp 1730882523
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_134
timestamp 1730882523
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_135
timestamp 1730882523
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_136
timestamp 1730882523
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_137
timestamp 1730882523
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_138
timestamp 1730882523
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_139
timestamp 1730882523
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_140
timestamp 1730882523
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_141
timestamp 1730882523
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_142
timestamp 1730882523
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_143
timestamp 1730882523
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_144
timestamp 1730882523
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_145
timestamp 1730882523
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_146
timestamp 1730882523
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_147
timestamp 1730882523
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_148
timestamp 1730882523
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_149
timestamp 1730882523
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_150
timestamp 1730882523
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_151
timestamp 1730882523
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_152
timestamp 1730882523
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_153
timestamp 1730882523
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_154
timestamp 1730882523
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_155
timestamp 1730882523
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_156
timestamp 1730882523
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_157
timestamp 1730882523
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_158
timestamp 1730882523
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_159
timestamp 1730882523
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_160
timestamp 1730882523
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_161
timestamp 1730882523
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_162
timestamp 1730882523
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_163
timestamp 1730882523
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_164
timestamp 1730882523
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_165
timestamp 1730882523
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_166
timestamp 1730882523
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_167
timestamp 1730882523
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_168
timestamp 1730882523
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_169
timestamp 1730882523
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_170
timestamp 1730882523
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_171
timestamp 1730882523
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_172
timestamp 1730882523
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_173
timestamp 1730882523
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_174
timestamp 1730882523
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_175
timestamp 1730882523
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_176
timestamp 1730882523
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_177
timestamp 1730882523
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_178
timestamp 1730882523
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_179
timestamp 1730882523
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_180
timestamp 1730882523
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_181
timestamp 1730882523
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_182
timestamp 1730882523
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_183
timestamp 1730882523
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_184
timestamp 1730882523
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_185
timestamp 1730882523
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_186
timestamp 1730882523
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_187
timestamp 1730882523
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_188
timestamp 1730882523
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_189
timestamp 1730882523
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_190
timestamp 1730882523
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_191
timestamp 1730882523
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_192
timestamp 1730882523
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_193
timestamp 1730882523
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_194
timestamp 1730882523
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_195
timestamp 1730882523
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_196
timestamp 1730882523
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_197
timestamp 1730882523
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_198
timestamp 1730882523
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_199
timestamp 1730882523
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_200
timestamp 1730882523
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_201
timestamp 1730882523
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_202
timestamp 1730882523
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_203
timestamp 1730882523
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_204
timestamp 1730882523
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_205
timestamp 1730882523
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_206
timestamp 1730882523
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_207
timestamp 1730882523
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_208
timestamp 1730882523
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_209
timestamp 1730882523
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_210
timestamp 1730882523
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_211
timestamp 1730882523
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_212
timestamp 1730882523
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_213
timestamp 1730882523
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_214
timestamp 1730882523
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_215
timestamp 1730882523
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_216
timestamp 1730882523
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_217
timestamp 1730882523
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_218
timestamp 1730882523
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_219
timestamp 1730882523
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_220
timestamp 1730882523
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_221
timestamp 1730882523
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_222
timestamp 1730882523
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_223
timestamp 1730882523
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_224
timestamp 1730882523
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_225
timestamp 1730882523
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_226
timestamp 1730882523
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_227
timestamp 1730882523
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_228
timestamp 1730882523
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_229
timestamp 1730882523
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_230
timestamp 1730882523
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_231
timestamp 1730882523
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_232
timestamp 1730882523
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_233
timestamp 1730882523
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_234
timestamp 1730882523
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_235
timestamp 1730882523
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_236
timestamp 1730882523
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_237
timestamp 1730882523
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_238
timestamp 1730882523
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_239
timestamp 1730882523
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_240
timestamp 1730882523
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_241
timestamp 1730882523
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_242
timestamp 1730882523
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_243
timestamp 1730882523
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_244
timestamp 1730882523
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_245
timestamp 1730882523
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_246
timestamp 1730882523
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_247
timestamp 1730882523
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_248
timestamp 1730882523
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_249
timestamp 1730882523
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_250
timestamp 1730882523
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_251
timestamp 1730882523
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_252
timestamp 1730882523
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_253
timestamp 1730882523
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_254
timestamp 1730882523
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_255
timestamp 1730882523
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_256
timestamp 1730882523
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_257
timestamp 1730882523
transform 1 0 6256 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_258
timestamp 1730882523
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_259
timestamp 1730882523
transform 1 0 11408 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_260
timestamp 1730882523
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  wire62
timestamp 1730882523
transform -1 0 6900 0 -1 11968
box -38 -48 314 592
<< labels >>
flabel metal4 s 4868 2128 5188 33232 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4208 2128 4528 33232 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 21088 800 21208 0 FreeSans 480 0 0 0 b0
port 2 nsew signal input
flabel metal3 s 0 25168 800 25288 0 FreeSans 480 0 0 0 b1
port 3 nsew signal input
flabel metal3 s 0 31288 800 31408 0 FreeSans 480 0 0 0 clk
port 4 nsew signal input
flabel metal3 s 16989 31288 17789 31408 0 FreeSans 480 0 0 0 compr
port 5 nsew signal input
flabel metal3 s 16989 3408 17789 3528 0 FreeSans 480 0 0 0 dac[0]
port 6 nsew signal output
flabel metal3 s 16989 17008 17789 17128 0 FreeSans 480 0 0 0 dac[1]
port 7 nsew signal output
flabel metal3 s 16989 30608 17789 30728 0 FreeSans 480 0 0 0 dac[2]
port 8 nsew signal output
flabel metal3 s 16989 18368 17789 18488 0 FreeSans 480 0 0 0 dac[3]
port 9 nsew signal output
flabel metal3 s 16989 21088 17789 21208 0 FreeSans 480 0 0 0 dac[4]
port 10 nsew signal output
flabel metal3 s 16989 12928 17789 13048 0 FreeSans 480 0 0 0 dac[5]
port 11 nsew signal output
flabel metal3 s 16989 13608 17789 13728 0 FreeSans 480 0 0 0 dac[6]
port 12 nsew signal output
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 dac[7]
port 13 nsew signal output
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 dac_coupl
port 14 nsew signal output
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 m0
port 15 nsew signal input
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 m1
port 16 nsew signal input
flabel metal3 s 16989 17688 17789 17808 0 FreeSans 480 0 0 0 reg0[0]
port 17 nsew signal output
flabel metal3 s 16989 29928 17789 30048 0 FreeSans 480 0 0 0 reg0[1]
port 18 nsew signal output
flabel metal2 s 14830 34714 14886 35514 0 FreeSans 224 90 0 0 reg0[2]
port 19 nsew signal output
flabel metal3 s 16989 14288 17789 14408 0 FreeSans 480 0 0 0 reg0[3]
port 20 nsew signal output
flabel metal3 s 16989 25168 17789 25288 0 FreeSans 480 0 0 0 reg0[4]
port 21 nsew signal output
flabel metal3 s 16989 14968 17789 15088 0 FreeSans 480 0 0 0 reg0[5]
port 22 nsew signal output
flabel metal2 s 15474 34714 15530 35514 0 FreeSans 224 90 0 0 reg0[6]
port 23 nsew signal output
flabel metal3 s 16989 22448 17789 22568 0 FreeSans 480 0 0 0 reg0[7]
port 24 nsew signal output
flabel metal3 s 16989 4768 17789 4888 0 FreeSans 480 0 0 0 reg1[0]
port 25 nsew signal output
flabel metal3 s 16989 5448 17789 5568 0 FreeSans 480 0 0 0 reg1[1]
port 26 nsew signal output
flabel metal3 s 16989 9528 17789 9648 0 FreeSans 480 0 0 0 reg1[2]
port 27 nsew signal output
flabel metal3 s 16989 4088 17789 4208 0 FreeSans 480 0 0 0 reg1[3]
port 28 nsew signal output
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 reg1[4]
port 29 nsew signal output
flabel metal3 s 16989 12248 17789 12368 0 FreeSans 480 0 0 0 reg1[5]
port 30 nsew signal output
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 reg1[6]
port 31 nsew signal output
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 reg1[7]
port 32 nsew signal output
flabel metal3 s 16989 8848 17789 8968 0 FreeSans 480 0 0 0 reg2[0]
port 33 nsew signal output
flabel metal3 s 16989 8168 17789 8288 0 FreeSans 480 0 0 0 reg2[1]
port 34 nsew signal output
flabel metal3 s 16989 10208 17789 10328 0 FreeSans 480 0 0 0 reg2[2]
port 35 nsew signal output
flabel metal3 s 16989 10888 17789 11008 0 FreeSans 480 0 0 0 reg2[3]
port 36 nsew signal output
flabel metal3 s 16989 6128 17789 6248 0 FreeSans 480 0 0 0 reg2[4]
port 37 nsew signal output
flabel metal3 s 16989 11568 17789 11688 0 FreeSans 480 0 0 0 reg2[5]
port 38 nsew signal output
flabel metal3 s 16989 6808 17789 6928 0 FreeSans 480 0 0 0 reg2[6]
port 39 nsew signal output
flabel metal3 s 16989 7488 17789 7608 0 FreeSans 480 0 0 0 reg2[7]
port 40 nsew signal output
flabel metal3 s 16989 19048 17789 19168 0 FreeSans 480 0 0 0 reg3[0]
port 41 nsew signal output
flabel metal3 s 16989 25848 17789 25968 0 FreeSans 480 0 0 0 reg3[1]
port 42 nsew signal output
flabel metal3 s 16989 28568 17789 28688 0 FreeSans 480 0 0 0 reg3[2]
port 43 nsew signal output
flabel metal3 s 16989 21768 17789 21888 0 FreeSans 480 0 0 0 reg3[3]
port 44 nsew signal output
flabel metal3 s 16989 24488 17789 24608 0 FreeSans 480 0 0 0 reg3[4]
port 45 nsew signal output
flabel metal3 s 16989 15648 17789 15768 0 FreeSans 480 0 0 0 reg3[5]
port 46 nsew signal output
flabel metal3 s 16989 27888 17789 28008 0 FreeSans 480 0 0 0 reg3[6]
port 47 nsew signal output
flabel metal3 s 16989 23128 17789 23248 0 FreeSans 480 0 0 0 reg3[7]
port 48 nsew signal output
flabel metal3 s 16989 19728 17789 19848 0 FreeSans 480 0 0 0 reg4[0]
port 49 nsew signal output
flabel metal3 s 16989 26528 17789 26648 0 FreeSans 480 0 0 0 reg4[1]
port 50 nsew signal output
flabel metal2 s 12898 34714 12954 35514 0 FreeSans 224 90 0 0 reg4[2]
port 51 nsew signal output
flabel metal3 s 16989 20408 17789 20528 0 FreeSans 480 0 0 0 reg4[3]
port 52 nsew signal output
flabel metal3 s 16989 23808 17789 23928 0 FreeSans 480 0 0 0 reg4[4]
port 53 nsew signal output
flabel metal3 s 16989 16328 17789 16448 0 FreeSans 480 0 0 0 reg4[5]
port 54 nsew signal output
flabel metal2 s 13542 34714 13598 35514 0 FreeSans 224 90 0 0 reg4[6]
port 55 nsew signal output
flabel metal3 s 16989 27208 17789 27328 0 FreeSans 480 0 0 0 reg4[7]
port 56 nsew signal output
flabel metal3 s 16989 29248 17789 29368 0 FreeSans 480 0 0 0 rst
port 57 nsew signal input
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 rx
port 58 nsew signal input
flabel metal2 s 7746 34714 7802 35514 0 FreeSans 224 90 0 0 tx
port 59 nsew signal output
rlabel metal1 8878 32640 8878 32640 0 VGND
rlabel metal1 8878 33184 8878 33184 0 VPWR
rlabel via1 11725 4590 11725 4590 0 _0000_
rlabel metal1 12139 14314 12139 14314 0 _0001_
rlabel metal1 1600 19822 1600 19822 0 _0002_
rlabel metal1 2111 20502 2111 20502 0 _0003_
rlabel metal1 1656 23290 1656 23290 0 _0004_
rlabel via1 1789 24174 1789 24174 0 _0005_
rlabel metal2 2438 27098 2438 27098 0 _0006_
rlabel metal2 2622 27302 2622 27302 0 _0007_
rlabel via1 3537 26962 3537 26962 0 _0008_
rlabel metal2 4646 26928 4646 26928 0 _0009_
rlabel metal1 5198 26214 5198 26214 0 _0010_
rlabel metal1 5239 23698 5239 23698 0 _0011_
rlabel via1 6214 23086 6214 23086 0 _0012_
rlabel metal1 7410 20502 7410 20502 0 _0013_
rlabel via1 5653 19822 5653 19822 0 _0014_
rlabel metal1 8643 3094 8643 3094 0 _0015_
rlabel metal1 11132 13906 11132 13906 0 _0016_
rlabel metal1 14260 19482 14260 19482 0 _0017_
rlabel metal1 14577 27370 14577 27370 0 _0018_
rlabel metal1 13616 30634 13616 30634 0 _0019_
rlabel metal1 13554 20502 13554 20502 0 _0020_
rlabel metal1 13795 23766 13795 23766 0 _0021_
rlabel metal1 14152 16490 14152 16490 0 _0022_
rlabel via1 13574 32402 13574 32402 0 _0023_
rlabel metal1 15180 26554 15180 26554 0 _0024_
rlabel metal1 14996 18938 14996 18938 0 _0025_
rlabel metal1 15405 27030 15405 27030 0 _0026_
rlabel metal2 14858 30226 14858 30226 0 _0027_
rlabel metal1 14996 20570 14996 20570 0 _0028_
rlabel metal2 15502 24582 15502 24582 0 _0029_
rlabel metal1 15405 16150 15405 16150 0 _0030_
rlabel metal2 15594 30022 15594 30022 0 _0031_
rlabel metal1 14934 23018 14934 23018 0 _0032_
rlabel metal1 15026 8534 15026 8534 0 _0033_
rlabel via1 15221 7854 15221 7854 0 _0034_
rlabel metal1 14290 9962 14290 9962 0 _0035_
rlabel metal1 15026 10710 15026 10710 0 _0036_
rlabel metal1 15644 4114 15644 4114 0 _0037_
rlabel metal2 14858 11492 14858 11492 0 _0038_
rlabel metal1 15000 4522 15000 4522 0 _0039_
rlabel metal1 15230 7378 15230 7378 0 _0040_
rlabel metal1 15405 3502 15405 3502 0 _0041_
rlabel metal2 15594 6562 15594 6562 0 _0042_
rlabel metal2 13386 9078 13386 9078 0 _0043_
rlabel metal1 15267 3094 15267 3094 0 _0044_
rlabel metal1 13565 3026 13565 3026 0 _0045_
rlabel via1 15221 11118 15221 11118 0 _0046_
rlabel via1 13381 4114 13381 4114 0 _0047_
rlabel metal1 13110 6970 13110 6970 0 _0048_
rlabel metal1 14490 17850 14490 17850 0 _0049_
rlabel metal2 15318 28322 15318 28322 0 _0050_
rlabel metal1 13979 31314 13979 31314 0 _0051_
rlabel metal1 14991 13974 14991 13974 0 _0052_
rlabel metal1 15042 24582 15042 24582 0 _0053_
rlabel via1 14761 14382 14761 14382 0 _0054_
rlabel metal1 14628 32198 14628 32198 0 _0055_
rlabel metal1 14393 22610 14393 22610 0 _0056_
rlabel metal1 13524 22202 13524 22202 0 _0057_
rlabel metal1 12604 27098 12604 27098 0 _0058_
rlabel metal2 12374 30838 12374 30838 0 _0059_
rlabel metal1 13068 24106 13068 24106 0 _0060_
rlabel metal1 13033 25942 13033 25942 0 _0061_
rlabel metal1 11331 11798 11331 11798 0 _0062_
rlabel metal2 11822 30192 11822 30192 0 _0063_
rlabel metal1 13120 26350 13120 26350 0 _0064_
rlabel metal1 12374 12614 12374 12614 0 _0065_
rlabel metal1 12834 12682 12834 12682 0 _0066_
rlabel metal1 12599 29206 12599 29206 0 _0067_
rlabel metal1 12849 4182 12849 4182 0 _0068_
rlabel metal1 12604 8602 12604 8602 0 _0069_
rlabel metal1 5929 27370 5929 27370 0 _0070_
rlabel metal1 6803 26962 6803 26962 0 _0071_
rlabel via1 6757 31722 6757 31722 0 _0072_
rlabel metal2 6578 25636 6578 25636 0 _0073_
rlabel metal1 7176 24378 7176 24378 0 _0074_
rlabel metal1 8096 26554 8096 26554 0 _0075_
rlabel metal1 10074 30906 10074 30906 0 _0076_
rlabel metal1 9425 26350 9425 26350 0 _0077_
rlabel metal1 10483 27438 10483 27438 0 _0078_
rlabel metal2 9062 25670 9062 25670 0 _0079_
rlabel metal1 10575 31790 10575 31790 0 _0080_
rlabel metal2 10166 28934 10166 28934 0 _0081_
rlabel via1 8514 24174 8514 24174 0 _0082_
rlabel viali 5561 5678 5561 5678 0 _0083_
rlabel metal2 7038 7174 7038 7174 0 _0084_
rlabel metal1 5883 6698 5883 6698 0 _0085_
rlabel metal1 5239 7378 5239 7378 0 _0086_
rlabel metal2 6394 9826 6394 9826 0 _0087_
rlabel metal1 5152 11866 5152 11866 0 _0088_
rlabel metal1 5382 12954 5382 12954 0 _0089_
rlabel via1 5561 16558 5561 16558 0 _0090_
rlabel metal2 6026 16354 6026 16354 0 _0091_
rlabel metal1 7502 15470 7502 15470 0 _0092_
rlabel metal2 7314 11866 7314 11866 0 _0093_
rlabel metal2 8326 13124 8326 13124 0 _0094_
rlabel metal1 8786 9044 8786 9044 0 _0095_
rlabel metal1 7447 8942 7447 8942 0 _0096_
rlabel metal1 7677 8534 7677 8534 0 _0097_
rlabel metal1 8152 9554 8152 9554 0 _0098_
rlabel via1 8505 31314 8505 31314 0 _0099_
rlabel metal1 8126 30294 8126 30294 0 _0100_
rlabel metal1 8520 29138 8520 29138 0 _0101_
rlabel metal1 6624 29274 6624 29274 0 _0102_
rlabel metal1 6394 30022 6394 30022 0 _0103_
rlabel metal1 1656 15674 1656 15674 0 _0104_
rlabel metal1 3680 16762 3680 16762 0 _0105_
rlabel via1 1881 17170 1881 17170 0 _0106_
rlabel metal1 1600 16558 1600 16558 0 _0107_
rlabel metal1 1656 12954 1656 12954 0 _0108_
rlabel metal1 2632 11730 2632 11730 0 _0109_
rlabel metal2 1702 10914 1702 10914 0 _0110_
rlabel metal2 2530 7548 2530 7548 0 _0111_
rlabel via1 1881 7854 1881 7854 0 _0112_
rlabel metal1 3174 7480 3174 7480 0 _0113_
rlabel metal1 4834 5610 4834 5610 0 _0114_
rlabel metal1 3342 6358 3342 6358 0 _0115_
rlabel metal1 4365 6766 4365 6766 0 _0116_
rlabel via1 12277 13294 12277 13294 0 _0117_
rlabel metal2 10442 3638 10442 3638 0 _0118_
rlabel metal1 10902 22712 10902 22712 0 _0119_
rlabel metal2 9798 21318 9798 21318 0 _0120_
rlabel metal1 11546 23528 11546 23528 0 _0121_
rlabel metal1 10626 23290 10626 23290 0 _0122_
rlabel metal1 11592 23290 11592 23290 0 _0123_
rlabel metal1 11868 13158 11868 13158 0 _0124_
rlabel metal1 10672 26010 10672 26010 0 _0125_
rlabel metal2 12466 4216 12466 4216 0 _0126_
rlabel metal1 12236 17850 12236 17850 0 _0127_
rlabel metal2 13018 28322 13018 28322 0 _0128_
rlabel via1 12553 18734 12553 18734 0 _0129_
rlabel metal1 8510 12614 8510 12614 0 _0130_
rlabel via1 8321 13906 8321 13906 0 _0131_
rlabel metal1 9103 14994 9103 14994 0 _0132_
rlabel metal1 9425 19414 9425 19414 0 _0133_
rlabel via1 10630 7786 10630 7786 0 _0134_
rlabel metal1 9874 4522 9874 4522 0 _0135_
rlabel metal1 9742 3502 9742 3502 0 _0136_
rlabel metal1 8740 22202 8740 22202 0 _0137_
rlabel metal1 8326 19890 8326 19890 0 _0138_
rlabel via1 11817 7854 11817 7854 0 _0139_
rlabel metal1 11592 6970 11592 6970 0 _0140_
rlabel metal1 7360 17850 7360 17850 0 _0141_
rlabel metal1 8372 20026 8372 20026 0 _0142_
rlabel metal2 10442 9078 10442 9078 0 _0143_
rlabel metal2 11454 9554 11454 9554 0 _0144_
rlabel metal2 7590 18598 7590 18598 0 _0145_
rlabel metal1 12696 21114 12696 21114 0 _0146_
rlabel metal1 7176 25262 7176 25262 0 _0147_
rlabel metal1 11684 24174 11684 24174 0 _0148_
rlabel metal1 13386 16116 13386 16116 0 _0149_
rlabel metal1 13432 15402 13432 15402 0 _0150_
rlabel metal2 8786 18632 8786 18632 0 _0151_
rlabel metal1 9016 17306 9016 17306 0 _0152_
rlabel metal1 12880 15402 12880 15402 0 _0153_
rlabel metal2 3634 13005 3634 13005 0 _0154_
rlabel metal2 7314 13124 7314 13124 0 _0155_
rlabel metal2 12466 22151 12466 22151 0 _0156_
rlabel via2 3910 17629 3910 17629 0 _0157_
rlabel metal1 8602 7310 8602 7310 0 _0158_
rlabel metal1 10994 7786 10994 7786 0 _0159_
rlabel metal2 13662 7684 13662 7684 0 _0160_
rlabel metal1 10442 5338 10442 5338 0 _0161_
rlabel metal2 10994 9418 10994 9418 0 _0162_
rlabel metal1 8188 7310 8188 7310 0 _0163_
rlabel metal1 8472 8806 8472 8806 0 _0164_
rlabel metal1 4600 17850 4600 17850 0 _0165_
rlabel metal1 4474 9622 4474 9622 0 _0166_
rlabel metal2 3634 9316 3634 9316 0 _0167_
rlabel metal1 3496 9622 3496 9622 0 _0168_
rlabel metal1 4738 9486 4738 9486 0 _0169_
rlabel metal2 5382 18819 5382 18819 0 _0170_
rlabel metal1 3956 9690 3956 9690 0 _0171_
rlabel metal1 4600 9690 4600 9690 0 _0172_
rlabel metal1 4462 19482 4462 19482 0 _0173_
rlabel metal1 3220 19142 3220 19142 0 _0174_
rlabel metal2 3772 20740 3772 20740 0 _0175_
rlabel metal2 2392 22080 2392 22080 0 _0176_
rlabel metal1 2990 12750 2990 12750 0 _0177_
rlabel metal1 3220 12410 3220 12410 0 _0178_
rlabel metal1 3220 13430 3220 13430 0 _0179_
rlabel metal1 3910 12920 3910 12920 0 _0180_
rlabel metal1 4002 15504 4002 15504 0 _0181_
rlabel via2 4278 13277 4278 13277 0 _0182_
rlabel metal1 3634 15470 3634 15470 0 _0183_
rlabel metal1 3956 13702 3956 13702 0 _0184_
rlabel metal2 4002 16354 4002 16354 0 _0185_
rlabel metal2 3818 16762 3818 16762 0 _0186_
rlabel metal1 4186 14450 4186 14450 0 _0187_
rlabel metal2 3726 13260 3726 13260 0 _0188_
rlabel metal1 4094 12750 4094 12750 0 _0189_
rlabel metal1 4232 13430 4232 13430 0 _0190_
rlabel metal1 4508 13362 4508 13362 0 _0191_
rlabel metal2 4186 12988 4186 12988 0 _0192_
rlabel metal1 3588 12614 3588 12614 0 _0193_
rlabel metal1 4508 8942 4508 8942 0 _0194_
rlabel metal1 4324 9146 4324 9146 0 _0195_
rlabel metal1 3220 9690 3220 9690 0 _0196_
rlabel metal1 2254 15674 2254 15674 0 _0197_
rlabel metal1 4692 15674 4692 15674 0 _0198_
rlabel viali 3946 13940 3946 13940 0 _0199_
rlabel metal2 4094 12172 4094 12172 0 _0200_
rlabel metal1 3082 16490 3082 16490 0 _0201_
rlabel metal1 13478 8976 13478 8976 0 _0202_
rlabel via1 11554 3434 11554 3434 0 _0203_
rlabel metal1 11960 3706 11960 3706 0 _0204_
rlabel metal1 8786 18598 8786 18598 0 _0205_
rlabel via2 8786 15300 8786 15300 0 _0206_
rlabel metal1 6394 18224 6394 18224 0 _0207_
rlabel metal1 9936 17238 9936 17238 0 _0208_
rlabel metal1 12190 20910 12190 20910 0 _0209_
rlabel metal1 10994 15878 10994 15878 0 _0210_
rlabel metal1 10672 15130 10672 15130 0 _0211_
rlabel metal2 10626 14297 10626 14297 0 _0212_
rlabel metal1 10718 14552 10718 14552 0 _0213_
rlabel metal2 10626 15810 10626 15810 0 _0214_
rlabel metal1 11178 14484 11178 14484 0 _0215_
rlabel metal2 11914 16286 11914 16286 0 _0216_
rlabel metal1 8891 10982 8891 10982 0 _0217_
rlabel metal2 8970 9690 8970 9690 0 _0218_
rlabel metal2 9890 13345 9890 13345 0 _0219_
rlabel metal1 9798 18054 9798 18054 0 _0220_
rlabel metal2 11638 20910 11638 20910 0 _0221_
rlabel metal2 11730 16286 11730 16286 0 _0222_
rlabel metal1 9614 17136 9614 17136 0 _0223_
rlabel metal1 10764 17306 10764 17306 0 _0224_
rlabel metal1 11454 15402 11454 15402 0 _0225_
rlabel metal1 12558 14892 12558 14892 0 _0226_
rlabel metal1 12604 23018 12604 23018 0 _0227_
rlabel metal1 12374 15130 12374 15130 0 _0228_
rlabel metal1 6256 19142 6256 19142 0 _0229_
rlabel metal1 5796 19346 5796 19346 0 _0230_
rlabel metal2 5934 19550 5934 19550 0 _0231_
rlabel metal1 4278 20468 4278 20468 0 _0232_
rlabel metal2 3358 21318 3358 21318 0 _0233_
rlabel metal1 3266 21488 3266 21488 0 _0234_
rlabel metal1 3864 21318 3864 21318 0 _0235_
rlabel metal2 4140 23086 4140 23086 0 _0236_
rlabel metal1 4370 22610 4370 22610 0 _0237_
rlabel metal1 4646 23018 4646 23018 0 _0238_
rlabel metal1 4554 21930 4554 21930 0 _0239_
rlabel metal2 4370 21828 4370 21828 0 _0240_
rlabel metal1 4554 22576 4554 22576 0 _0241_
rlabel metal2 4876 21862 4876 21862 0 _0242_
rlabel metal1 4669 21998 4669 21998 0 _0243_
rlabel metal1 4002 23052 4002 23052 0 _0244_
rlabel metal1 3542 24106 3542 24106 0 _0245_
rlabel metal3 4071 20604 4071 20604 0 _0246_
rlabel metal2 3818 23290 3818 23290 0 _0247_
rlabel metal2 3910 21794 3910 21794 0 _0248_
rlabel metal1 4508 22066 4508 22066 0 _0249_
rlabel metal2 4646 21148 4646 21148 0 _0250_
rlabel metal2 4140 20026 4140 20026 0 _0251_
rlabel metal1 4830 19346 4830 19346 0 _0252_
rlabel metal1 5336 19482 5336 19482 0 _0253_
rlabel metal1 6624 21522 6624 21522 0 _0254_
rlabel metal2 3634 20230 3634 20230 0 _0255_
rlabel metal1 4416 20570 4416 20570 0 _0256_
rlabel metal1 5198 22746 5198 22746 0 _0257_
rlabel metal2 2990 20604 2990 20604 0 _0258_
rlabel metal2 2898 23392 2898 23392 0 _0259_
rlabel metal1 2300 22474 2300 22474 0 _0260_
rlabel metal1 2103 23018 2103 23018 0 _0261_
rlabel metal1 3174 24140 3174 24140 0 _0262_
rlabel metal2 2990 24004 2990 24004 0 _0263_
rlabel metal2 1886 24548 1886 24548 0 _0264_
rlabel metal1 2116 26554 2116 26554 0 _0265_
rlabel metal1 2070 26792 2070 26792 0 _0266_
rlabel metal2 1702 26724 1702 26724 0 _0267_
rlabel metal1 2655 26418 2655 26418 0 _0268_
rlabel via1 5392 26010 5392 26010 0 _0269_
rlabel metal2 3818 27676 3818 27676 0 _0270_
rlabel metal1 3094 27030 3094 27030 0 _0271_
rlabel metal1 4370 25806 4370 25806 0 _0272_
rlabel metal2 5842 25330 5842 25330 0 _0273_
rlabel metal1 5704 25874 5704 25874 0 _0274_
rlabel metal1 5658 26010 5658 26010 0 _0275_
rlabel metal1 6256 22066 6256 22066 0 _0276_
rlabel metal1 5474 24752 5474 24752 0 _0277_
rlabel metal1 5302 24242 5302 24242 0 _0278_
rlabel metal2 6762 21420 6762 21420 0 _0279_
rlabel metal2 5566 23324 5566 23324 0 _0280_
rlabel metal1 6176 20842 6176 20842 0 _0281_
rlabel metal1 5578 21590 5578 21590 0 _0282_
rlabel metal2 9614 4284 9614 4284 0 _0283_
rlabel metal2 12742 30464 12742 30464 0 _0284_
rlabel metal1 9668 10982 9668 10982 0 _0285_
rlabel metal1 13662 14382 13662 14382 0 _0286_
rlabel metal1 14398 14246 14398 14246 0 _0287_
rlabel via1 14122 17187 14122 17187 0 _0288_
rlabel metal1 13570 16524 13570 16524 0 _0289_
rlabel metal2 14490 18326 14490 18326 0 _0290_
rlabel metal2 14306 29002 14306 29002 0 _0291_
rlabel metal2 14812 32742 14812 32742 0 _0292_
rlabel metal2 12926 20604 12926 20604 0 _0293_
rlabel metal1 14582 24138 14582 24138 0 _0294_
rlabel metal1 13754 16150 13754 16150 0 _0295_
rlabel metal1 13800 30158 13800 30158 0 _0296_
rlabel metal1 16054 26316 16054 26316 0 _0297_
rlabel metal1 16146 19822 16146 19822 0 _0298_
rlabel metal1 15640 17578 15640 17578 0 _0299_
rlabel metal1 15318 18768 15318 18768 0 _0300_
rlabel metal1 15870 18394 15870 18394 0 _0301_
rlabel metal1 16146 22746 16146 22746 0 _0302_
rlabel metal1 15364 32742 15364 32742 0 _0303_
rlabel metal2 15410 20910 15410 20910 0 _0304_
rlabel metal2 15042 24004 15042 24004 0 _0305_
rlabel metal2 16054 17034 16054 17034 0 _0306_
rlabel metal1 16054 29682 16054 29682 0 _0307_
rlabel metal2 14306 23324 14306 23324 0 _0308_
rlabel metal2 16054 19176 16054 19176 0 _0309_
rlabel metal1 13524 6290 13524 6290 0 _0310_
rlabel metal1 14628 12818 14628 12818 0 _0311_
rlabel metal1 15318 8908 15318 8908 0 _0312_
rlabel metal1 14398 8500 14398 8500 0 _0313_
rlabel metal1 13754 10064 13754 10064 0 _0314_
rlabel metal2 14398 11084 14398 11084 0 _0315_
rlabel metal1 15962 5236 15962 5236 0 _0316_
rlabel metal1 14398 11186 14398 11186 0 _0317_
rlabel metal2 15226 5287 15226 5287 0 _0318_
rlabel metal1 14214 6426 14214 6426 0 _0319_
rlabel metal1 13340 15334 13340 15334 0 _0320_
rlabel metal1 13754 11050 13754 11050 0 _0321_
rlabel metal1 13432 11322 13432 11322 0 _0322_
rlabel metal1 15916 2618 15916 2618 0 _0323_
rlabel metal1 13386 5882 13386 5882 0 _0324_
rlabel metal1 13892 8466 13892 8466 0 _0325_
rlabel metal1 15410 3162 15410 3162 0 _0326_
rlabel metal1 14582 3570 14582 3570 0 _0327_
rlabel metal1 15732 9622 15732 9622 0 _0328_
rlabel metal1 13800 5202 13800 5202 0 _0329_
rlabel metal2 13570 6596 13570 6596 0 _0330_
rlabel metal2 14214 14756 14214 14756 0 _0331_
rlabel metal1 15502 17680 15502 17680 0 _0332_
rlabel metal2 14950 21420 14950 21420 0 _0333_
rlabel metal1 14858 17680 14858 17680 0 _0334_
rlabel metal2 15778 29580 15778 29580 0 _0335_
rlabel metal1 14582 32436 14582 32436 0 _0336_
rlabel metal1 16008 14586 16008 14586 0 _0337_
rlabel metal2 14398 25262 14398 25262 0 _0338_
rlabel metal1 14858 14960 14858 14960 0 _0339_
rlabel metal1 15318 32436 15318 32436 0 _0340_
rlabel metal1 15226 22474 15226 22474 0 _0341_
rlabel metal1 15134 17306 15134 17306 0 _0342_
rlabel metal1 14858 18700 14858 18700 0 _0343_
rlabel metal1 14214 18938 14214 18938 0 _0344_
rlabel via2 15686 6443 15686 6443 0 _0345_
rlabel metal1 16146 31926 16146 31926 0 _0346_
rlabel metal1 13202 26962 13202 26962 0 _0347_
rlabel via2 14582 9435 14582 9435 0 _0348_
rlabel metal3 12075 31892 12075 31892 0 _0349_
rlabel metal1 12834 30124 12834 30124 0 _0350_
rlabel metal1 16192 20026 16192 20026 0 _0351_
rlabel metal1 14858 12682 14858 12682 0 _0352_
rlabel metal1 15410 20570 15410 20570 0 _0353_
rlabel metal2 15594 24752 15594 24752 0 _0354_
rlabel metal2 14766 5933 14766 5933 0 _0355_
rlabel metal1 14306 25126 14306 25126 0 _0356_
rlabel metal2 15594 14484 15594 14484 0 _0357_
rlabel metal1 15732 15470 15732 15470 0 _0358_
rlabel metal1 12190 12818 12190 12818 0 _0359_
rlabel metal1 15824 32742 15824 32742 0 _0360_
rlabel metal1 14674 5576 14674 5576 0 _0361_
rlabel metal1 14168 28934 14168 28934 0 _0362_
rlabel metal1 14582 6970 14582 6970 0 _0363_
rlabel metal1 15502 23494 15502 23494 0 _0364_
rlabel metal2 15134 26656 15134 26656 0 _0365_
rlabel metal2 12926 4862 12926 4862 0 _0366_
rlabel metal2 13110 7412 13110 7412 0 _0367_
rlabel metal2 7314 27302 7314 27302 0 _0368_
rlabel metal1 6946 28118 6946 28118 0 _0369_
rlabel metal2 8050 24276 8050 24276 0 _0370_
rlabel metal3 7521 31756 7521 31756 0 _0371_
rlabel metal1 8924 29614 8924 29614 0 _0372_
rlabel metal1 8234 32402 8234 32402 0 _0373_
rlabel metal1 8050 31382 8050 31382 0 _0374_
rlabel metal1 8096 30702 8096 30702 0 _0375_
rlabel metal1 10948 29274 10948 29274 0 _0376_
rlabel metal2 9982 30294 9982 30294 0 _0377_
rlabel metal1 10534 29818 10534 29818 0 _0378_
rlabel metal1 9752 29614 9752 29614 0 _0379_
rlabel metal1 9016 28662 9016 28662 0 _0380_
rlabel metal1 9706 28730 9706 28730 0 _0381_
rlabel metal1 9798 30056 9798 30056 0 _0382_
rlabel metal1 10304 30158 10304 30158 0 _0383_
rlabel metal2 9890 29818 9890 29818 0 _0384_
rlabel metal1 9384 29818 9384 29818 0 _0385_
rlabel metal1 8556 31790 8556 31790 0 _0386_
rlabel metal1 8970 28186 8970 28186 0 _0387_
rlabel metal1 8510 30906 8510 30906 0 _0388_
rlabel metal1 7452 31450 7452 31450 0 _0389_
rlabel metal1 6946 28526 6946 28526 0 _0390_
rlabel metal1 9752 26010 9752 26010 0 _0391_
rlabel metal1 12466 30770 12466 30770 0 _0392_
rlabel metal1 10442 12920 10442 12920 0 _0393_
rlabel metal1 12282 27336 12282 27336 0 _0394_
rlabel metal2 10166 24786 10166 24786 0 _0395_
rlabel metal2 11546 31008 11546 31008 0 _0396_
rlabel metal1 10580 28186 10580 28186 0 _0397_
rlabel metal1 8924 23290 8924 23290 0 _0398_
rlabel metal2 5658 13532 5658 13532 0 _0399_
rlabel metal1 7682 6698 7682 6698 0 _0400_
rlabel metal2 5566 7378 5566 7378 0 _0401_
rlabel metal1 5658 8500 5658 8500 0 _0402_
rlabel metal1 5428 12614 5428 12614 0 _0403_
rlabel metal1 5750 12852 5750 12852 0 _0404_
rlabel metal1 5428 12818 5428 12818 0 _0405_
rlabel metal2 5842 13328 5842 13328 0 _0406_
rlabel metal2 6210 15266 6210 15266 0 _0407_
rlabel via1 6670 13787 6670 13787 0 _0408_
rlabel metal1 6762 13804 6762 13804 0 _0409_
rlabel metal2 6946 14076 6946 14076 0 _0410_
rlabel metal1 7038 14042 7038 14042 0 _0411_
rlabel metal1 7452 13158 7452 13158 0 _0412_
rlabel metal1 8234 12716 8234 12716 0 _0413_
rlabel metal1 7160 6698 7160 6698 0 _0414_
rlabel metal2 4738 8058 4738 8058 0 _0415_
rlabel metal1 5796 7990 5796 7990 0 _0416_
rlabel metal1 5934 8058 5934 8058 0 _0417_
rlabel metal2 6578 10268 6578 10268 0 _0418_
rlabel metal1 6240 9622 6240 9622 0 _0419_
rlabel metal1 4922 14246 4922 14246 0 _0420_
rlabel metal1 5428 11526 5428 11526 0 _0421_
rlabel metal1 4692 12682 4692 12682 0 _0422_
rlabel metal1 4784 12614 4784 12614 0 _0423_
rlabel metal1 5198 16762 5198 16762 0 _0424_
rlabel metal1 5428 15674 5428 15674 0 _0425_
rlabel metal1 6394 16082 6394 16082 0 _0426_
rlabel metal2 5842 16422 5842 16422 0 _0427_
rlabel metal2 5750 15538 5750 15538 0 _0428_
rlabel metal1 7038 15912 7038 15912 0 _0429_
rlabel metal1 6578 12750 6578 12750 0 _0430_
rlabel metal1 7925 11866 7925 11866 0 _0431_
rlabel metal1 9016 10098 9016 10098 0 _0432_
rlabel metal2 8418 32028 8418 32028 0 _0433_
rlabel metal1 9246 29172 9246 29172 0 _0434_
rlabel metal1 6762 29036 6762 29036 0 _0435_
rlabel metal2 8970 28934 8970 28934 0 _0436_
rlabel metal1 6256 28526 6256 28526 0 _0437_
rlabel metal1 7038 29172 7038 29172 0 _0438_
rlabel metal2 3358 16286 3358 16286 0 _0439_
rlabel metal2 3542 16320 3542 16320 0 _0440_
rlabel metal2 2530 16252 2530 16252 0 _0441_
rlabel metal2 4738 15419 4738 15419 0 _0442_
rlabel metal1 2530 15130 2530 15130 0 _0443_
rlabel metal1 2024 14994 2024 14994 0 _0444_
rlabel metal2 2162 16524 2162 16524 0 _0445_
rlabel metal1 1840 15130 1840 15130 0 _0446_
rlabel metal1 1932 12954 1932 12954 0 _0447_
rlabel metal1 2024 12886 2024 12886 0 _0448_
rlabel metal2 2254 11968 2254 11968 0 _0449_
rlabel metal1 2438 11254 2438 11254 0 _0450_
rlabel metal1 3036 11322 3036 11322 0 _0451_
rlabel metal1 2438 10642 2438 10642 0 _0452_
rlabel metal1 3128 10642 3128 10642 0 _0453_
rlabel metal1 2300 10574 2300 10574 0 _0454_
rlabel via1 2354 6698 2354 6698 0 _0455_
rlabel metal1 1426 7446 1426 7446 0 _0456_
rlabel metal2 1610 8228 1610 8228 0 _0457_
rlabel metal2 1518 8160 1518 8160 0 _0458_
rlabel metal1 3182 6630 3182 6630 0 _0459_
rlabel metal2 4186 7956 4186 7956 0 _0460_
rlabel metal1 3810 7514 3810 7514 0 _0461_
rlabel metal1 3266 6222 3266 6222 0 _0462_
rlabel metal2 5474 7378 5474 7378 0 _0463_
rlabel metal1 4278 6630 4278 6630 0 _0464_
rlabel via1 2998 6698 2998 6698 0 _0465_
rlabel metal1 10948 14586 10948 14586 0 _0466_
rlabel metal2 12466 14348 12466 14348 0 _0467_
rlabel metal2 12834 14144 12834 14144 0 _0468_
rlabel via1 10994 4250 10994 4250 0 _0469_
rlabel metal2 9430 17612 9430 17612 0 _0470_
rlabel metal1 11500 20842 11500 20842 0 _0471_
rlabel metal1 10580 22202 10580 22202 0 _0472_
rlabel metal1 10258 18938 10258 18938 0 _0473_
rlabel metal2 10902 19924 10902 19924 0 _0474_
rlabel metal1 11132 18734 11132 18734 0 _0475_
rlabel metal1 10488 20570 10488 20570 0 _0476_
rlabel metal1 11178 23086 11178 23086 0 _0477_
rlabel metal2 10166 18857 10166 18857 0 _0478_
rlabel metal1 11224 21522 11224 21522 0 _0479_
rlabel metal1 11132 23290 11132 23290 0 _0480_
rlabel metal1 11868 23290 11868 23290 0 _0481_
rlabel metal2 11730 19142 11730 19142 0 _0482_
rlabel metal2 11638 19584 11638 19584 0 _0483_
rlabel metal1 9982 19788 9982 19788 0 _0484_
rlabel metal1 11362 23290 11362 23290 0 _0485_
rlabel metal2 11730 21318 11730 21318 0 _0486_
rlabel metal1 11822 22202 11822 22202 0 _0487_
rlabel metal1 11546 13192 11546 13192 0 _0488_
rlabel metal2 11546 16439 11546 16439 0 _0489_
rlabel metal2 10442 15946 10442 15946 0 _0490_
rlabel via1 9141 18666 9141 18666 0 _0491_
rlabel metal1 9890 15028 9890 15028 0 _0492_
rlabel metal4 12604 8160 12604 8160 0 _0493_
rlabel metal1 12052 15470 12052 15470 0 _0494_
rlabel metal3 12673 15300 12673 15300 0 _0495_
rlabel metal2 11730 18156 11730 18156 0 _0496_
rlabel metal2 13938 18020 13938 18020 0 _0497_
rlabel metal1 13064 17510 13064 17510 0 _0498_
rlabel metal2 11914 21114 11914 21114 0 _0499_
rlabel metal3 12811 27676 12811 27676 0 _0500_
rlabel metal2 12558 23902 12558 23902 0 _0501_
rlabel metal2 13110 25908 13110 25908 0 _0502_
rlabel metal1 11776 19822 11776 19822 0 _0503_
rlabel metal2 13110 19482 13110 19482 0 _0504_
rlabel metal2 11914 19142 11914 19142 0 _0505_
rlabel metal1 12742 19482 12742 19482 0 _0506_
rlabel metal1 9890 16014 9890 16014 0 _0507_
rlabel metal1 9522 16592 9522 16592 0 _0508_
rlabel metal2 9430 16388 9430 16388 0 _0509_
rlabel metal2 9338 14042 9338 14042 0 _0510_
rlabel metal1 9844 12206 9844 12206 0 _0511_
rlabel metal1 9200 12410 9200 12410 0 _0512_
rlabel metal1 9476 19822 9476 19822 0 _0513_
rlabel metal1 10258 5678 10258 5678 0 _0514_
rlabel metal2 9522 4828 9522 4828 0 _0515_
rlabel metal1 8464 4114 8464 4114 0 _0516_
rlabel via3 9315 16524 9315 16524 0 _0517_
rlabel metal2 12374 8602 12374 8602 0 _0518_
rlabel metal1 13110 7752 13110 7752 0 _0519_
rlabel metal1 8924 18938 8924 18938 0 _0520_
rlabel metal1 7314 17578 7314 17578 0 _0521_
rlabel metal1 11684 6426 11684 6426 0 _0522_
rlabel metal2 7958 18020 7958 18020 0 _0523_
rlabel metal2 13294 21148 13294 21148 0 _0524_
rlabel metal1 12696 21046 12696 21046 0 _0525_
rlabel metal2 13202 21964 13202 21964 0 _0526_
rlabel metal3 751 21148 751 21148 0 b0
rlabel metal3 751 25228 751 25228 0 b1
rlabel metal1 8970 17680 8970 17680 0 clk
rlabel metal1 13708 21930 13708 21930 0 clknet_0_clk
rlabel metal1 1610 7990 1610 7990 0 clknet_4_0_0_clk
rlabel metal1 1472 24174 1472 24174 0 clknet_4_10_0_clk
rlabel metal1 6693 31790 6693 31790 0 clknet_4_11_0_clk
rlabel metal1 9384 21522 9384 21522 0 clknet_4_12_0_clk
rlabel metal1 14398 18190 14398 18190 0 clknet_4_13_0_clk
rlabel metal1 12742 28084 12742 28084 0 clknet_4_14_0_clk
rlabel metal2 14950 27778 14950 27778 0 clknet_4_15_0_clk
rlabel metal1 5336 5678 5336 5678 0 clknet_4_1_0_clk
rlabel metal1 1426 13430 1426 13430 0 clknet_4_2_0_clk
rlabel metal1 8096 15538 8096 15538 0 clknet_4_3_0_clk
rlabel metal2 9890 3808 9890 3808 0 clknet_4_4_0_clk
rlabel metal2 12558 8160 12558 8160 0 clknet_4_5_0_clk
rlabel metal1 14122 9996 14122 9996 0 clknet_4_6_0_clk
rlabel metal1 14536 14382 14536 14382 0 clknet_4_7_0_clk
rlabel metal1 1472 20366 1472 20366 0 clknet_4_8_0_clk
rlabel metal2 6946 18768 6946 18768 0 clknet_4_9_0_clk
rlabel via2 16330 31331 16330 31331 0 compr
rlabel metal1 8096 15130 8096 15130 0 control.baud_clk
rlabel metal1 3542 16082 3542 16082 0 control.baud_rate_gen.count\[0\]
rlabel metal2 4140 10540 4140 10540 0 control.baud_rate_gen.count\[10\]
rlabel metal2 3450 6528 3450 6528 0 control.baud_rate_gen.count\[11\]
rlabel metal1 5198 8942 5198 8942 0 control.baud_rate_gen.count\[12\]
rlabel metal2 4094 16762 4094 16762 0 control.baud_rate_gen.count\[1\]
rlabel metal1 3312 17782 3312 17782 0 control.baud_rate_gen.count\[2\]
rlabel metal1 3129 17646 3129 17646 0 control.baud_rate_gen.count\[3\]
rlabel metal2 2438 13362 2438 13362 0 control.baud_rate_gen.count\[4\]
rlabel metal2 1518 12002 1518 12002 0 control.baud_rate_gen.count\[5\]
rlabel metal1 2852 12138 2852 12138 0 control.baud_rate_gen.count\[6\]
rlabel metal2 2346 8704 2346 8704 0 control.baud_rate_gen.count\[7\]
rlabel metal1 2645 8874 2645 8874 0 control.baud_rate_gen.count\[8\]
rlabel metal1 3266 7854 3266 7854 0 control.baud_rate_gen.count\[9\]
rlabel metal1 6660 14994 6660 14994 0 control.baud_rate_gen.n805_o
rlabel metal1 8510 18836 8510 18836 0 control.n576_q\[0\]
rlabel metal1 7038 18598 7038 18598 0 control.n576_q\[1\]
rlabel metal1 8372 19482 8372 19482 0 control.n576_q\[2\]
rlabel metal1 8418 21114 8418 21114 0 control.n579_q
rlabel metal1 9246 16082 9246 16082 0 control.n588_o
rlabel metal2 14214 4080 14214 4080 0 control.n598_o
rlabel metal1 13938 18156 13938 18156 0 control.n600_o
rlabel metal1 14444 29138 14444 29138 0 control.n602_o
rlabel metal2 13938 19006 13938 19006 0 control.n604_o
rlabel metal1 14398 21420 14398 21420 0 control.n606_o
rlabel metal1 13800 13430 13800 13430 0 control.n608_o
rlabel metal1 13248 14246 13248 14246 0 control.n610_o
rlabel metal1 10028 12750 10028 12750 0 control.n612_o
rlabel via1 9798 23086 9798 23086 0 control.n633_o
rlabel metal1 10994 21012 10994 21012 0 control.n635_o
rlabel metal2 11362 27744 11362 27744 0 control.n637_o
rlabel metal2 10626 24038 10626 24038 0 control.n639_o
rlabel metal2 13018 26350 13018 26350 0 control.n641_o
rlabel metal1 10810 12954 10810 12954 0 control.n643_o
rlabel metal1 12696 30566 12696 30566 0 control.n645_o
rlabel metal2 10442 24242 10442 24242 0 control.n647_o
rlabel metal1 9844 19822 9844 19822 0 control.n651_o
rlabel metal1 10120 18802 10120 18802 0 control.n653_o
rlabel metal3 15924 3468 15924 3468 0 dac[0]
rlabel via2 15226 17051 15226 17051 0 dac[1]
rlabel metal2 10442 32241 10442 32241 0 dac[2]
rlabel metal2 13110 17867 13110 17867 0 dac[3]
rlabel metal2 16238 21505 16238 21505 0 dac[4]
rlabel metal2 16238 13515 16238 13515 0 dac[5]
rlabel metal2 15410 13583 15410 13583 0 dac[6]
rlabel metal2 8418 1520 8418 1520 0 dac[7]
rlabel metal2 9062 1520 9062 1520 0 dac_coupl
rlabel metal2 7774 1554 7774 1554 0 m0
rlabel metal2 7130 1588 7130 1588 0 m1
rlabel metal1 14076 13770 14076 13770 0 n119_q\[0\]
rlabel metal1 14076 15334 14076 15334 0 n119_q\[1\]
rlabel metal1 14812 29614 14812 29614 0 n119_q\[2\]
rlabel metal1 8372 22202 8372 22202 0 n120_q
rlabel metal2 9522 22712 9522 22712 0 n126_q\[0\]
rlabel metal1 13478 27880 13478 27880 0 n126_q\[1\]
rlabel metal1 13846 30838 13846 30838 0 n126_q\[2\]
rlabel metal2 12006 24820 12006 24820 0 n126_q\[3\]
rlabel metal1 12880 25670 12880 25670 0 n126_q\[4\]
rlabel metal2 10810 13362 10810 13362 0 n126_q\[5\]
rlabel metal2 12834 30464 12834 30464 0 n126_q\[6\]
rlabel metal1 12926 28152 12926 28152 0 n126_q\[7\]
rlabel metal1 6762 22950 6762 22950 0 n127_q
rlabel metal1 2530 19448 2530 19448 0 net1
rlabel metal1 12926 30158 12926 30158 0 net10
rlabel metal2 6946 29308 6946 29308 0 net100
rlabel metal1 11316 32266 11316 32266 0 net101
rlabel metal1 11086 28526 11086 28526 0 net102
rlabel metal1 13478 20910 13478 20910 0 net103
rlabel metal2 8510 26860 8510 26860 0 net104
rlabel metal1 11500 31858 11500 31858 0 net105
rlabel metal2 10074 6426 10074 6426 0 net106
rlabel metal1 13294 21998 13294 21998 0 net107
rlabel metal1 10258 26962 10258 26962 0 net108
rlabel metal1 14766 26010 14766 26010 0 net109
rlabel metal2 13294 17884 13294 17884 0 net11
rlabel metal2 13570 27642 13570 27642 0 net110
rlabel metal1 9706 25126 9706 25126 0 net111
rlabel metal1 13570 28186 13570 28186 0 net112
rlabel metal1 13432 5338 13432 5338 0 net113
rlabel metal2 12834 27948 12834 27948 0 net114
rlabel metal1 10902 26010 10902 26010 0 net115
rlabel metal2 12098 24412 12098 24412 0 net116
rlabel metal2 7038 26384 7038 26384 0 net117
rlabel metal1 7038 26010 7038 26010 0 net118
rlabel metal2 6578 12988 6578 12988 0 net119
rlabel metal1 15778 21658 15778 21658 0 net12
rlabel via1 7778 12818 7778 12818 0 net120
rlabel metal1 9660 21862 9660 21862 0 net121
rlabel metal1 6440 30362 6440 30362 0 net122
rlabel metal1 9292 12818 9292 12818 0 net123
rlabel metal1 7360 18666 7360 18666 0 net124
rlabel metal2 7958 20026 7958 20026 0 net125
rlabel metal2 8878 20706 8878 20706 0 net126
rlabel metal1 13570 29614 13570 29614 0 net127
rlabel metal2 9062 10166 9062 10166 0 net128
rlabel metal1 8418 10098 8418 10098 0 net129
rlabel metal1 15778 12954 15778 12954 0 net13
rlabel metal1 8280 8058 8280 8058 0 net130
rlabel metal2 9706 6834 9706 6834 0 net131
rlabel metal3 7613 31892 7613 31892 0 net132
rlabel metal1 8924 29274 8924 29274 0 net133
rlabel metal1 13156 12954 13156 12954 0 net134
rlabel metal1 7268 24174 7268 24174 0 net135
rlabel metal2 11086 20604 11086 20604 0 net136
rlabel metal1 9062 31994 9062 31994 0 net137
rlabel metal1 13892 12954 13892 12954 0 net138
rlabel metal2 12282 24752 12282 24752 0 net139
rlabel metal2 15226 13668 15226 13668 0 net14
rlabel metal1 9200 6834 9200 6834 0 net140
rlabel metal1 8694 3366 8694 3366 0 net15
rlabel metal1 9338 2414 9338 2414 0 net16
rlabel metal2 15318 17408 15318 17408 0 net17
rlabel metal1 15456 31790 15456 31790 0 net18
rlabel metal2 14306 32623 14306 32623 0 net19
rlabel metal2 3542 24956 3542 24956 0 net2
rlabel metal1 15594 12784 15594 12784 0 net20
rlabel metal1 16284 25126 16284 25126 0 net21
rlabel metal1 15962 14246 15962 14246 0 net22
rlabel metal1 12190 32844 12190 32844 0 net23
rlabel metal1 14536 21998 14536 21998 0 net24
rlabel metal1 15640 2414 15640 2414 0 net25
rlabel metal2 16238 6460 16238 6460 0 net26
rlabel metal1 14306 9010 14306 9010 0 net27
rlabel metal1 14904 2414 14904 2414 0 net28
rlabel metal1 14352 3162 14352 3162 0 net29
rlabel metal1 12788 20910 12788 20910 0 net3
rlabel metal1 15594 13226 15594 13226 0 net30
rlabel metal1 13570 2414 13570 2414 0 net31
rlabel metal1 14306 2414 14306 2414 0 net32
rlabel metal1 16284 18734 16284 18734 0 net33
rlabel metal1 16192 8058 16192 8058 0 net34
rlabel metal2 14858 10098 14858 10098 0 net35
rlabel metal2 14352 16116 14352 16116 0 net36
rlabel metal2 15042 4794 15042 4794 0 net37
rlabel metal1 16376 15470 16376 15470 0 net38
rlabel metal1 14398 5644 14398 5644 0 net39
rlabel metal1 8648 2550 8648 2550 0 net4
rlabel metal1 14490 6698 14490 6698 0 net40
rlabel metal1 15272 18326 15272 18326 0 net41
rlabel metal2 16330 24684 16330 24684 0 net42
rlabel metal1 15870 32402 15870 32402 0 net43
rlabel metal1 16146 20774 16146 20774 0 net44
rlabel metal1 14536 23766 14536 23766 0 net45
rlabel metal1 14950 15878 14950 15878 0 net46
rlabel metal1 10304 28526 10304 28526 0 net47
rlabel metal1 15686 23766 15686 23766 0 net48
rlabel metal1 13984 19822 13984 19822 0 net49
rlabel metal1 8418 2482 8418 2482 0 net5
rlabel metal1 15410 27302 15410 27302 0 net50
rlabel metal2 11546 32436 11546 32436 0 net51
rlabel metal1 16008 20434 16008 20434 0 net52
rlabel metal1 13754 24208 13754 24208 0 net53
rlabel metal1 14076 16082 14076 16082 0 net54
rlabel metal2 11362 32708 11362 32708 0 net55
rlabel metal2 13478 26809 13478 26809 0 net56
rlabel metal2 8142 32334 8142 32334 0 net57
rlabel metal1 4922 12886 4922 12886 0 net58
rlabel metal1 4922 26418 4922 26418 0 net59
rlabel metal1 10948 32878 10948 32878 0 net6
rlabel metal1 1886 15402 1886 15402 0 net60
rlabel metal2 2346 17170 2346 17170 0 net61
rlabel metal1 7360 10778 7360 10778 0 net62
rlabel metal1 2806 27098 2806 27098 0 net63
rlabel metal1 13110 12784 13110 12784 0 net64
rlabel metal1 13018 23698 13018 23698 0 net65
rlabel metal1 11500 31790 11500 31790 0 net66
rlabel metal1 15134 12784 15134 12784 0 net67
rlabel metal1 15870 17136 15870 17136 0 net68
rlabel metal2 9982 21454 9982 21454 0 net69
rlabel metal1 10488 2550 10488 2550 0 net7
rlabel metal1 5060 21454 5060 21454 0 net70
rlabel metal2 2622 25585 2622 25585 0 net71
rlabel metal2 14674 29206 14674 29206 0 net72
rlabel metal1 4922 9146 4922 9146 0 net73
rlabel metal1 4784 19210 4784 19210 0 net74
rlabel metal2 9154 3774 9154 3774 0 net75
rlabel metal1 13938 7854 13938 7854 0 net76
rlabel metal2 12696 8500 12696 8500 0 net77
rlabel metal1 12006 32300 12006 32300 0 net78
rlabel metal2 10810 32606 10810 32606 0 net79
rlabel metal1 14536 2822 14536 2822 0 net8
rlabel metal1 11132 21454 11132 21454 0 net80
rlabel metal1 2369 19346 2369 19346 0 net81
rlabel via2 3174 17187 3174 17187 0 net82
rlabel metal1 2438 15436 2438 15436 0 net83
rlabel metal2 7590 21794 7590 21794 0 net84
rlabel metal1 8372 10234 8372 10234 0 net85
rlabel metal2 10994 23358 10994 23358 0 net86
rlabel metal2 9798 3944 9798 3944 0 net87
rlabel metal2 10626 22780 10626 22780 0 net88
rlabel metal2 12190 29818 12190 29818 0 net89
rlabel metal2 15042 17340 15042 17340 0 net9
rlabel metal1 13018 30362 13018 30362 0 net90
rlabel metal1 13156 19346 13156 19346 0 net91
rlabel metal1 8602 7378 8602 7378 0 net92
rlabel metal1 11316 13294 11316 13294 0 net93
rlabel metal1 13018 17646 13018 17646 0 net94
rlabel metal1 12052 12954 12052 12954 0 net95
rlabel metal1 13754 27098 13754 27098 0 net96
rlabel metal1 12972 13906 12972 13906 0 net97
rlabel metal2 13386 25024 13386 25024 0 net98
rlabel metal1 12788 14994 12788 14994 0 net99
rlabel metal2 13846 17459 13846 17459 0 reg0[0]
rlabel metal1 15364 29002 15364 29002 0 reg0[1]
rlabel metal1 14306 33082 14306 33082 0 reg0[2]
rlabel metal3 13846 13940 13846 13940 0 reg0[3]
rlabel metal2 13938 24939 13938 24939 0 reg0[4]
rlabel metal3 16660 15028 16660 15028 0 reg0[5]
rlabel metal1 12052 32742 12052 32742 0 reg0[6]
rlabel metal1 14352 21862 14352 21862 0 reg0[7]
rlabel metal3 16614 4828 16614 4828 0 reg1[0]
rlabel via2 12374 5525 12374 5525 0 reg1[1]
rlabel metal1 12052 5882 12052 5882 0 reg1[2]
rlabel metal3 16108 4148 16108 4148 0 reg1[3]
rlabel metal2 13570 1520 13570 1520 0 reg1[4]
rlabel metal2 15042 12359 15042 12359 0 reg1[5]
rlabel metal2 12926 1520 12926 1520 0 reg1[6]
rlabel metal2 14214 1520 14214 1520 0 reg1[7]
rlabel metal1 14168 10234 14168 10234 0 reg2[0]
rlabel metal2 16238 7871 16238 7871 0 reg2[1]
rlabel metal1 14122 10506 14122 10506 0 reg2[2]
rlabel metal2 16238 10047 16238 10047 0 reg2[3]
rlabel metal1 13846 6154 13846 6154 0 reg2[4]
rlabel metal2 13662 11203 13662 11203 0 reg2[5]
rlabel metal1 14996 6426 14996 6426 0 reg2[6]
rlabel metal2 12834 6817 12834 6817 0 reg2[7]
rlabel metal2 14214 18751 14214 18751 0 reg3[0]
rlabel metal2 16238 26877 16238 26877 0 reg3[1]
rlabel metal2 11270 27965 11270 27965 0 reg3[2]
rlabel via2 15870 21845 15870 21845 0 reg3[3]
rlabel metal2 12190 24837 12190 24837 0 reg3[4]
rlabel metal1 13984 16218 13984 16218 0 reg3[5]
rlabel metal1 12466 28560 12466 28560 0 reg3[6]
rlabel metal3 16108 23188 16108 23188 0 reg3[7]
rlabel metal1 14490 19686 14490 19686 0 reg4[0]
rlabel metal2 11086 26027 11086 26027 0 reg4[1]
rlabel metal2 12926 33908 12926 33908 0 reg4[2]
rlabel metal1 16284 21318 16284 21318 0 reg4[3]
rlabel metal1 14214 23562 14214 23562 0 reg4[4]
rlabel metal1 14260 17034 14260 17034 0 reg4[5]
rlabel metal2 13570 33874 13570 33874 0 reg4[6]
rlabel via3 13869 31892 13869 31892 0 reg4[7]
rlabel metal2 16330 29223 16330 29223 0 rst
rlabel metal2 9706 1554 9706 1554 0 rx
rlabel metal1 7866 33082 7866 33082 0 tx
rlabel metal1 8372 9146 8372 9146 0 uart_receive.baud_clk
rlabel metal2 8602 10302 8602 10302 0 uart_receive.baud_clk2
rlabel metal2 11178 8092 11178 8092 0 uart_receive.baud_clk3
rlabel metal1 5612 7786 5612 7786 0 uart_receive.baud_rate_gen.count\[0\]
rlabel metal1 6210 12852 6210 12852 0 uart_receive.baud_rate_gen.count\[10\]
rlabel metal1 6302 14246 6302 14246 0 uart_receive.baud_rate_gen.count\[11\]
rlabel metal2 6026 7446 6026 7446 0 uart_receive.baud_rate_gen.count\[1\]
rlabel metal2 6118 7616 6118 7616 0 uart_receive.baud_rate_gen.count\[2\]
rlabel metal1 5980 7854 5980 7854 0 uart_receive.baud_rate_gen.count\[3\]
rlabel metal1 6118 11866 6118 11866 0 uart_receive.baud_rate_gen.count\[4\]
rlabel metal1 6072 14382 6072 14382 0 uart_receive.baud_rate_gen.count\[5\]
rlabel metal1 4922 14042 4922 14042 0 uart_receive.baud_rate_gen.count\[6\]
rlabel metal2 6302 15946 6302 15946 0 uart_receive.baud_rate_gen.count\[7\]
rlabel metal2 5934 16966 5934 16966 0 uart_receive.baud_rate_gen.count\[8\]
rlabel metal1 7038 15674 7038 15674 0 uart_receive.baud_rate_gen.count\[9\]
rlabel metal1 8326 7514 8326 7514 0 uart_receive.n328_o\[0\]
rlabel metal1 8786 7276 8786 7276 0 uart_receive.n328_o\[1\]
rlabel metal1 7084 10030 7084 10030 0 uart_receive.n345_q
rlabel metal1 9706 10676 9706 10676 0 uart_receive.n346_q\[0\]
rlabel metal1 10626 7174 10626 7174 0 uart_receive.n346_q\[1\]
rlabel metal1 13018 8058 13018 8058 0 uart_receive.n352_o
rlabel metal1 13110 7854 13110 7854 0 uart_receive.n354_o
rlabel metal1 10304 8058 10304 8058 0 uart_receive.n360_o
rlabel metal1 12788 12750 12788 12750 0 uart_receive.n370_o
rlabel metal1 13708 12750 13708 12750 0 uart_receive.n372_o
rlabel metal1 14398 32436 14398 32436 0 uart_receive.n374_o
rlabel metal2 15410 15079 15410 15079 0 uart_receive.n376_o
rlabel metal1 14076 4590 14076 4590 0 uart_receive.n378_o
rlabel metal1 13846 16558 13846 16558 0 uart_receive.n380_o
rlabel metal1 15088 32402 15088 32402 0 uart_receive.n382_o
rlabel metal1 13708 21046 13708 21046 0 uart_receive.n384_o
rlabel metal1 6624 27302 6624 27302 0 uart_transmit.baud_clk
rlabel via1 2262 22746 2262 22746 0 uart_transmit.baud_rate_gen.count\[0\]
rlabel metal1 5980 21590 5980 21590 0 uart_transmit.baud_rate_gen.count\[10\]
rlabel metal1 6578 20910 6578 20910 0 uart_transmit.baud_rate_gen.count\[11\]
rlabel metal1 6532 20026 6532 20026 0 uart_transmit.baud_rate_gen.count\[12\]
rlabel metal1 2300 22406 2300 22406 0 uart_transmit.baud_rate_gen.count\[1\]
rlabel metal1 2346 22644 2346 22644 0 uart_transmit.baud_rate_gen.count\[2\]
rlabel metal2 3082 23868 3082 23868 0 uart_transmit.baud_rate_gen.count\[3\]
rlabel metal1 4002 24106 4002 24106 0 uart_transmit.baud_rate_gen.count\[4\]
rlabel metal2 4002 26928 4002 26928 0 uart_transmit.baud_rate_gen.count\[5\]
rlabel metal1 4692 27098 4692 27098 0 uart_transmit.baud_rate_gen.count\[6\]
rlabel metal1 4876 24718 4876 24718 0 uart_transmit.baud_rate_gen.count\[7\]
rlabel metal1 5482 20366 5482 20366 0 uart_transmit.baud_rate_gen.count\[8\]
rlabel metal1 6072 23494 6072 23494 0 uart_transmit.baud_rate_gen.count\[9\]
rlabel metal1 8832 25330 8832 25330 0 uart_transmit.n167_o
rlabel metal1 8326 28050 8326 28050 0 uart_transmit.n224_q
rlabel metal2 7866 25670 7866 25670 0 uart_transmit.n226_q\[0\]
rlabel metal1 6946 32368 6946 32368 0 uart_transmit.n226_q\[1\]
rlabel metal1 9476 31790 9476 31790 0 uart_transmit.n227_q\[0\]
rlabel metal2 8510 30770 8510 30770 0 uart_transmit.n227_q\[1\]
rlabel metal2 10166 30498 10166 30498 0 uart_transmit.n227_q\[2\]
rlabel metal1 6946 29682 6946 29682 0 uart_transmit.n227_q\[3\]
rlabel metal2 6118 31076 6118 31076 0 uart_transmit.n227_q\[4\]
rlabel metal2 8786 27268 8786 27268 0 uart_transmit.n231_o
rlabel metal1 11592 31450 11592 31450 0 uart_transmit.n232_o
rlabel metal2 10350 28016 10350 28016 0 uart_transmit.n233_o
rlabel metal2 11638 28084 11638 28084 0 uart_transmit.n234_o
rlabel metal1 9430 26010 9430 26010 0 uart_transmit.n235_o
rlabel metal1 11040 31926 11040 31926 0 uart_transmit.n236_o
rlabel metal1 10856 29002 10856 29002 0 uart_transmit.n237_o
<< properties >>
string FIXED_BBOX 0 0 17789 35514
<< end >>
