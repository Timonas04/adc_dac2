VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_tim2305_adc_dac
  CLASS BLOCK ;
  FOREIGN tt_um_tim2305_adc_dac ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 240.000000 ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.200000 ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.200000 ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.200000 ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.200000 ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.200000 ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.200000 ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.200000 ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.200000 ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 112.465 219.150 113.275 219.290 ;
        RECT 112.275 218.980 113.275 219.150 ;
        RECT 112.465 217.920 113.275 218.980 ;
        RECT 112.465 217.770 113.275 217.910 ;
        RECT 112.275 217.600 113.275 217.770 ;
        RECT 112.465 212.400 113.275 217.600 ;
        RECT 112.465 212.250 113.275 212.390 ;
        RECT 112.275 212.080 113.275 212.250 ;
        RECT 112.465 208.720 113.275 212.080 ;
        RECT 112.305 208.455 112.415 208.575 ;
        RECT 112.465 208.110 113.145 208.250 ;
        RECT 112.275 207.940 113.145 208.110 ;
        RECT 112.465 207.765 113.145 207.940 ;
        RECT 112.465 206.420 113.375 207.765 ;
        RECT 112.550 205.970 113.335 206.400 ;
        RECT 112.305 205.695 112.415 205.815 ;
        RECT 112.465 204.145 113.375 205.490 ;
        RECT 112.465 203.970 113.145 204.145 ;
        RECT 112.275 203.800 113.145 203.970 ;
        RECT 112.465 203.660 113.145 203.800 ;
        RECT 112.465 203.510 113.145 203.650 ;
        RECT 112.275 203.340 113.145 203.510 ;
        RECT 112.465 200.135 113.145 203.340 ;
        RECT 112.465 199.225 113.365 200.135 ;
        RECT 112.465 197.690 113.145 199.225 ;
        RECT 112.465 196.340 113.375 197.690 ;
        RECT 112.465 194.945 113.375 196.290 ;
        RECT 112.465 194.770 113.145 194.945 ;
        RECT 112.275 194.600 113.145 194.770 ;
        RECT 112.465 194.460 113.145 194.600 ;
        RECT 112.310 194.140 112.420 194.300 ;
        RECT 112.550 193.090 113.335 193.520 ;
        RECT 112.310 192.760 112.420 192.920 ;
        RECT 112.465 192.010 113.145 192.150 ;
        RECT 112.275 191.840 113.145 192.010 ;
        RECT 112.465 191.665 113.145 191.840 ;
        RECT 112.465 190.320 113.375 191.665 ;
        RECT 112.465 189.260 113.245 190.310 ;
        RECT 112.275 189.090 113.245 189.260 ;
        RECT 112.465 188.940 113.245 189.090 ;
        RECT 112.310 188.620 112.420 188.780 ;
        RECT 112.465 187.870 113.145 188.010 ;
        RECT 112.275 187.700 113.145 187.870 ;
        RECT 112.465 186.190 113.145 187.700 ;
        RECT 112.465 185.260 113.375 186.190 ;
        RECT 112.305 184.995 112.415 185.115 ;
        RECT 112.465 183.730 113.275 184.790 ;
        RECT 112.275 183.560 113.275 183.730 ;
        RECT 112.465 183.420 113.275 183.560 ;
      LAYER nwell ;
        RECT 113.665 183.225 116.495 219.485 ;
      LAYER pwell ;
        RECT 116.885 219.150 117.695 219.290 ;
        RECT 117.905 219.150 118.715 219.290 ;
        RECT 116.885 218.980 118.715 219.150 ;
        RECT 116.885 217.920 117.695 218.980 ;
        RECT 117.905 217.920 118.715 218.980 ;
        RECT 116.785 216.565 117.695 217.910 ;
        RECT 117.015 216.390 117.695 216.565 ;
        RECT 117.905 216.520 118.815 217.870 ;
        RECT 117.015 216.220 117.885 216.390 ;
        RECT 117.015 216.080 117.695 216.220 ;
        RECT 117.740 215.760 117.850 215.920 ;
        RECT 116.785 214.735 117.695 215.150 ;
        RECT 117.905 214.985 118.585 216.520 ;
        RECT 116.785 214.565 117.885 214.735 ;
        RECT 116.785 214.220 117.695 214.565 ;
        RECT 117.015 211.250 117.695 214.220 ;
        RECT 117.905 214.075 118.805 214.985 ;
        RECT 116.885 210.870 117.695 211.010 ;
        RECT 117.905 210.870 118.585 214.075 ;
        RECT 116.885 210.700 118.585 210.870 ;
        RECT 116.885 207.340 117.695 210.700 ;
        RECT 117.905 210.560 118.585 210.700 ;
        RECT 117.905 210.410 118.715 210.550 ;
        RECT 117.715 210.240 118.715 210.410 ;
        RECT 116.885 207.190 117.695 207.330 ;
        RECT 116.885 207.020 117.885 207.190 ;
        RECT 116.885 205.960 117.695 207.020 ;
        RECT 117.905 206.880 118.715 210.240 ;
        RECT 117.745 206.615 117.855 206.735 ;
        RECT 117.990 205.970 118.775 206.400 ;
        RECT 116.785 204.560 117.695 205.910 ;
        RECT 117.905 205.810 118.585 205.950 ;
        RECT 117.715 205.640 118.585 205.810 ;
        RECT 117.015 203.025 117.695 204.560 ;
        RECT 116.795 202.115 117.695 203.025 ;
        RECT 117.015 198.910 117.695 202.115 ;
        RECT 117.015 198.740 117.885 198.910 ;
        RECT 117.015 198.600 117.695 198.740 ;
        RECT 116.785 198.175 117.695 198.590 ;
        RECT 116.785 198.005 117.885 198.175 ;
        RECT 116.785 197.660 117.695 198.005 ;
        RECT 117.015 194.690 117.695 197.660 ;
        RECT 117.905 196.845 118.585 205.640 ;
        RECT 117.905 196.610 118.715 196.750 ;
        RECT 117.715 196.440 118.715 196.610 ;
        RECT 117.905 195.380 118.715 196.440 ;
        RECT 117.905 195.230 118.685 195.370 ;
        RECT 117.715 195.060 118.685 195.230 ;
        RECT 117.740 194.140 117.850 194.300 ;
        RECT 117.905 194.000 118.685 195.060 ;
        RECT 117.905 193.850 118.685 193.990 ;
        RECT 117.715 193.680 118.685 193.850 ;
        RECT 116.825 193.090 117.610 193.520 ;
        RECT 116.785 192.055 117.695 192.975 ;
        RECT 117.905 192.620 118.685 193.680 ;
        RECT 117.905 192.470 118.685 192.610 ;
        RECT 117.715 192.300 118.685 192.470 ;
        RECT 117.015 189.710 117.695 192.055 ;
        RECT 117.905 191.240 118.685 192.300 ;
        RECT 117.905 191.090 118.685 191.230 ;
        RECT 117.715 190.920 118.685 191.090 ;
        RECT 117.905 189.860 118.685 190.920 ;
        RECT 117.015 189.540 117.885 189.710 ;
        RECT 117.015 189.510 117.695 189.540 ;
        RECT 117.740 189.080 117.850 189.240 ;
        RECT 117.905 188.795 118.815 189.830 ;
        RECT 117.715 188.625 118.815 188.795 ;
        RECT 117.905 188.480 118.815 188.625 ;
        RECT 116.785 186.030 117.695 188.470 ;
        RECT 117.905 188.330 118.815 188.390 ;
        RECT 117.715 188.160 118.815 188.330 ;
        RECT 116.785 185.860 117.885 186.030 ;
        RECT 116.785 185.720 117.695 185.860 ;
        RECT 117.740 185.400 117.850 185.560 ;
        RECT 117.905 184.940 118.815 188.160 ;
        RECT 116.885 183.730 117.695 184.790 ;
        RECT 117.905 183.730 118.715 184.790 ;
        RECT 116.885 183.560 118.715 183.730 ;
        RECT 116.885 183.420 117.695 183.560 ;
        RECT 117.905 183.420 118.715 183.560 ;
      LAYER nwell ;
        RECT 119.105 183.225 121.935 219.485 ;
      LAYER pwell ;
        RECT 122.325 219.150 123.135 219.290 ;
        RECT 123.345 219.150 124.155 219.290 ;
        RECT 122.325 218.980 124.155 219.150 ;
        RECT 122.325 217.920 123.135 218.980 ;
        RECT 123.345 217.920 124.155 218.980 ;
        RECT 122.225 216.565 123.135 217.910 ;
        RECT 123.345 217.770 124.025 217.910 ;
        RECT 123.155 217.600 124.025 217.770 ;
        RECT 122.455 216.390 123.135 216.565 ;
        RECT 122.455 216.220 123.325 216.390 ;
        RECT 122.455 216.080 123.135 216.220 ;
        RECT 123.180 215.760 123.290 215.920 ;
        RECT 122.455 215.010 123.135 215.040 ;
        RECT 122.455 214.840 123.325 215.010 ;
        RECT 122.455 212.495 123.135 214.840 ;
        RECT 122.225 211.575 123.135 212.495 ;
        RECT 123.345 214.395 124.025 217.600 ;
        RECT 123.345 213.485 124.245 214.395 ;
        RECT 123.345 211.950 124.025 213.485 ;
        RECT 123.180 211.160 123.290 211.320 ;
        RECT 123.345 210.600 124.255 211.950 ;
        RECT 122.455 210.410 123.135 210.440 ;
        RECT 123.345 210.410 124.155 210.550 ;
        RECT 122.455 210.240 124.155 210.410 ;
        RECT 122.455 207.895 123.135 210.240 ;
        RECT 122.225 206.975 123.135 207.895 ;
        RECT 123.345 206.880 124.155 210.240 ;
        RECT 122.455 203.670 123.135 206.640 ;
        RECT 123.185 206.615 123.295 206.735 ;
        RECT 123.430 205.970 124.215 206.400 ;
        RECT 123.345 205.810 124.025 205.950 ;
        RECT 123.155 205.640 124.025 205.810 ;
        RECT 122.225 203.325 123.135 203.670 ;
        RECT 122.225 203.155 123.325 203.325 ;
        RECT 122.225 202.740 123.135 203.155 ;
        RECT 122.325 202.590 123.135 202.730 ;
        RECT 122.325 202.420 123.325 202.590 ;
        RECT 123.345 202.435 124.025 205.640 ;
        RECT 122.325 200.900 123.135 202.420 ;
        RECT 123.345 201.525 124.245 202.435 ;
        RECT 122.455 200.750 123.135 200.890 ;
        RECT 122.455 200.580 123.325 200.750 ;
        RECT 122.455 197.375 123.135 200.580 ;
        RECT 123.345 199.990 124.025 201.525 ;
        RECT 123.345 198.640 124.255 199.990 ;
        RECT 123.345 198.445 124.025 198.590 ;
        RECT 123.155 198.275 124.025 198.445 ;
        RECT 122.235 196.465 123.135 197.375 ;
        RECT 122.455 194.930 123.135 196.465 ;
        RECT 123.345 196.745 124.025 198.275 ;
        RECT 123.345 195.380 124.255 196.745 ;
        RECT 123.345 195.230 124.155 195.370 ;
        RECT 123.155 195.060 124.155 195.230 ;
        RECT 122.225 193.580 123.135 194.930 ;
        RECT 122.265 193.090 123.050 193.520 ;
        RECT 122.225 192.655 123.135 193.070 ;
        RECT 122.225 192.485 123.325 192.655 ;
        RECT 123.345 192.620 124.155 195.060 ;
        RECT 122.225 192.140 123.135 192.485 ;
        RECT 123.185 192.355 123.295 192.475 ;
        RECT 122.455 189.170 123.135 192.140 ;
        RECT 123.345 192.010 124.025 192.040 ;
        RECT 123.155 191.840 124.025 192.010 ;
        RECT 123.345 189.495 124.025 191.840 ;
        RECT 122.355 188.790 123.135 188.930 ;
        RECT 122.355 188.620 123.325 188.790 ;
        RECT 122.355 187.560 123.135 188.620 ;
        RECT 123.345 188.575 124.255 189.495 ;
        RECT 123.345 188.330 124.255 188.390 ;
        RECT 123.155 188.160 124.255 188.330 ;
        RECT 122.225 186.605 123.135 187.550 ;
        RECT 122.425 185.115 123.105 186.605 ;
        RECT 123.345 185.390 124.255 188.160 ;
        RECT 122.425 184.945 123.325 185.115 ;
        RECT 122.425 184.800 123.105 184.945 ;
        RECT 122.325 183.730 123.135 184.790 ;
        RECT 123.345 183.730 124.155 184.790 ;
        RECT 122.325 183.560 124.155 183.730 ;
        RECT 122.325 183.420 123.135 183.560 ;
        RECT 123.345 183.420 124.155 183.560 ;
      LAYER nwell ;
        RECT 124.545 183.225 127.375 219.485 ;
      LAYER pwell ;
        RECT 127.765 219.150 128.575 219.290 ;
        RECT 128.785 219.150 129.595 219.290 ;
        RECT 127.765 218.980 129.595 219.150 ;
        RECT 127.765 217.920 128.575 218.980 ;
        RECT 128.785 217.920 129.595 218.980 ;
        RECT 127.665 216.565 128.575 217.910 ;
        RECT 128.785 217.770 129.595 217.910 ;
        RECT 128.595 217.600 129.595 217.770 ;
        RECT 127.895 216.390 128.575 216.565 ;
        RECT 128.785 216.540 129.595 217.600 ;
        RECT 128.785 216.390 129.465 216.420 ;
        RECT 127.895 216.220 129.465 216.390 ;
        RECT 127.895 216.080 128.575 216.220 ;
        RECT 128.625 215.815 128.735 215.935 ;
        RECT 127.665 215.195 128.575 215.610 ;
        RECT 127.665 215.025 128.765 215.195 ;
        RECT 127.665 214.680 128.575 215.025 ;
        RECT 127.895 211.710 128.575 214.680 ;
        RECT 128.785 213.875 129.465 216.220 ;
        RECT 128.785 212.955 129.695 213.875 ;
        RECT 128.785 211.835 129.695 212.755 ;
        RECT 127.895 211.330 128.575 211.470 ;
        RECT 127.895 211.160 128.765 211.330 ;
        RECT 127.895 207.955 128.575 211.160 ;
        RECT 128.785 209.490 129.465 211.835 ;
        RECT 128.595 209.320 129.465 209.490 ;
        RECT 128.785 209.290 129.465 209.320 ;
        RECT 128.785 209.030 129.595 209.170 ;
        RECT 128.595 208.860 129.595 209.030 ;
        RECT 127.675 207.045 128.575 207.955 ;
        RECT 127.895 205.510 128.575 207.045 ;
        RECT 128.785 206.420 129.595 208.860 ;
        RECT 128.870 205.970 129.655 206.400 ;
        RECT 127.665 204.160 128.575 205.510 ;
        RECT 128.785 204.895 129.695 205.930 ;
        RECT 128.595 204.725 129.695 204.895 ;
        RECT 128.785 204.580 129.695 204.725 ;
        RECT 127.665 203.695 128.575 204.110 ;
        RECT 127.665 203.525 128.765 203.695 ;
        RECT 127.665 203.180 128.575 203.525 ;
        RECT 127.895 200.210 128.575 203.180 ;
        RECT 128.785 200.750 129.695 204.500 ;
        RECT 128.595 200.580 129.695 200.750 ;
        RECT 128.785 200.440 129.695 200.580 ;
        RECT 127.665 198.955 128.575 199.875 ;
        RECT 127.895 196.610 128.575 198.955 ;
        RECT 128.785 199.415 129.695 200.335 ;
        RECT 128.785 197.070 129.465 199.415 ;
        RECT 128.595 196.900 129.465 197.070 ;
        RECT 128.785 196.870 129.465 196.900 ;
        RECT 128.785 196.610 129.595 196.750 ;
        RECT 127.895 196.440 129.595 196.610 ;
        RECT 127.895 196.410 128.575 196.440 ;
        RECT 127.765 196.150 128.575 196.290 ;
        RECT 127.765 195.980 128.765 196.150 ;
        RECT 127.765 193.540 128.575 195.980 ;
        RECT 128.785 195.380 129.595 196.440 ;
        RECT 128.785 194.420 129.695 195.370 ;
        RECT 127.705 193.090 128.490 193.520 ;
        RECT 127.665 190.175 128.575 192.780 ;
        RECT 128.815 192.015 129.495 194.420 ;
        RECT 128.595 191.845 129.495 192.015 ;
        RECT 128.815 191.700 129.495 191.845 ;
        RECT 128.785 191.545 129.695 191.690 ;
        RECT 128.595 191.375 129.695 191.545 ;
        RECT 128.785 190.340 129.695 191.375 ;
        RECT 127.665 190.160 128.765 190.175 ;
        RECT 128.785 190.160 129.565 190.310 ;
        RECT 127.665 190.005 129.565 190.160 ;
        RECT 127.665 189.860 128.575 190.005 ;
        RECT 128.595 189.990 129.565 190.005 ;
        RECT 128.620 189.540 128.730 189.700 ;
        RECT 128.785 188.940 129.565 189.990 ;
        RECT 127.665 185.570 128.575 188.790 ;
        RECT 128.785 185.570 129.695 188.790 ;
        RECT 127.665 185.400 129.695 185.570 ;
        RECT 127.665 185.340 128.575 185.400 ;
        RECT 128.785 185.340 129.695 185.400 ;
        RECT 128.625 184.995 128.735 185.115 ;
        RECT 127.765 183.730 128.575 184.790 ;
        RECT 128.785 183.730 129.595 184.790 ;
        RECT 127.765 183.560 129.595 183.730 ;
        RECT 127.765 183.420 128.575 183.560 ;
        RECT 128.785 183.420 129.595 183.560 ;
      LAYER nwell ;
        RECT 129.985 183.225 132.815 219.485 ;
      LAYER pwell ;
        RECT 133.205 219.150 134.015 219.290 ;
        RECT 134.225 219.150 135.035 219.290 ;
        RECT 133.205 218.980 135.035 219.150 ;
        RECT 133.205 217.920 134.015 218.980 ;
        RECT 134.225 217.920 135.035 218.980 ;
        RECT 133.105 216.520 134.015 217.870 ;
        RECT 134.225 217.495 135.135 217.910 ;
        RECT 134.035 217.325 135.135 217.495 ;
        RECT 133.335 214.985 134.015 216.520 ;
        RECT 133.115 214.075 134.015 214.985 ;
        RECT 133.335 210.870 134.015 214.075 ;
        RECT 134.225 216.980 135.135 217.325 ;
        RECT 134.225 214.010 134.905 216.980 ;
        RECT 134.225 213.630 134.905 213.770 ;
        RECT 134.035 213.460 134.905 213.630 ;
        RECT 133.335 210.700 134.205 210.870 ;
        RECT 133.335 210.560 134.015 210.700 ;
        RECT 133.205 210.410 134.015 210.550 ;
        RECT 133.205 210.240 134.205 210.410 ;
        RECT 134.225 210.255 134.905 213.460 ;
        RECT 133.205 207.800 134.015 210.240 ;
        RECT 134.225 209.345 135.125 210.255 ;
        RECT 134.225 207.810 134.905 209.345 ;
        RECT 134.065 207.535 134.175 207.655 ;
        RECT 133.335 207.190 134.015 207.330 ;
        RECT 133.335 207.020 134.205 207.190 ;
        RECT 133.335 198.225 134.015 207.020 ;
        RECT 134.225 206.460 135.135 207.810 ;
        RECT 134.310 205.970 135.095 206.400 ;
        RECT 134.225 205.810 134.905 205.950 ;
        RECT 134.035 205.640 134.905 205.810 ;
        RECT 134.225 202.435 134.905 205.640 ;
        RECT 134.225 201.525 135.125 202.435 ;
        RECT 134.225 199.990 134.905 201.525 ;
        RECT 134.225 198.640 135.135 199.990 ;
        RECT 134.065 198.335 134.175 198.455 ;
        RECT 133.105 197.115 134.015 198.035 ;
        RECT 133.335 194.770 134.015 197.115 ;
        RECT 134.225 196.765 135.135 198.130 ;
        RECT 134.225 195.235 134.905 196.765 ;
        RECT 134.035 195.065 134.905 195.235 ;
        RECT 134.225 194.920 134.905 195.065 ;
        RECT 133.335 194.600 134.205 194.770 ;
        RECT 133.335 194.570 134.015 194.600 ;
        RECT 134.060 194.140 134.170 194.300 ;
        RECT 134.225 193.850 135.135 193.910 ;
        RECT 134.035 193.680 135.135 193.850 ;
        RECT 133.145 193.090 133.930 193.520 ;
        RECT 133.305 192.935 133.985 193.060 ;
        RECT 133.305 192.765 134.205 192.935 ;
        RECT 133.305 191.735 133.985 192.765 ;
        RECT 133.105 190.780 134.015 191.735 ;
        RECT 134.225 190.910 135.135 193.680 ;
        RECT 133.205 190.630 134.015 190.770 ;
        RECT 133.205 190.625 134.205 190.630 ;
        RECT 134.225 190.625 135.135 190.770 ;
        RECT 133.205 190.460 135.135 190.625 ;
        RECT 133.205 188.020 134.015 190.460 ;
        RECT 134.035 190.455 135.135 190.460 ;
        RECT 134.225 189.420 135.135 190.455 ;
        RECT 134.065 189.135 134.175 189.255 ;
        RECT 134.225 188.790 135.135 188.850 ;
        RECT 134.035 188.620 135.135 188.790 ;
        RECT 134.065 187.755 134.175 187.875 ;
        RECT 133.105 186.495 134.015 187.530 ;
        RECT 133.105 186.325 134.205 186.495 ;
        RECT 133.105 186.180 134.015 186.325 ;
        RECT 133.235 185.110 134.015 186.170 ;
        RECT 134.225 185.400 135.135 188.620 ;
        RECT 134.065 185.110 134.175 185.115 ;
        RECT 133.235 184.940 134.205 185.110 ;
        RECT 133.235 184.800 134.015 184.940 ;
        RECT 133.205 183.730 134.015 184.790 ;
        RECT 134.225 183.730 135.035 184.790 ;
        RECT 133.205 183.560 135.035 183.730 ;
        RECT 133.205 183.420 134.015 183.560 ;
        RECT 134.225 183.420 135.035 183.560 ;
      LAYER nwell ;
        RECT 135.425 183.225 138.255 219.485 ;
      LAYER pwell ;
        RECT 138.645 219.150 139.455 219.290 ;
        RECT 139.665 219.150 140.475 219.290 ;
        RECT 138.645 218.980 140.475 219.150 ;
        RECT 138.645 217.920 139.455 218.980 ;
        RECT 139.665 217.920 140.475 218.980 ;
        RECT 138.545 216.565 139.455 217.910 ;
        RECT 139.665 217.770 140.345 217.910 ;
        RECT 139.475 217.600 140.345 217.770 ;
        RECT 138.775 216.390 139.455 216.565 ;
        RECT 138.775 216.220 139.645 216.390 ;
        RECT 138.775 216.080 139.455 216.220 ;
        RECT 138.545 215.655 139.455 216.070 ;
        RECT 138.545 215.485 139.645 215.655 ;
        RECT 138.545 215.140 139.455 215.485 ;
        RECT 138.775 212.170 139.455 215.140 ;
        RECT 139.665 214.395 140.345 217.600 ;
        RECT 139.665 213.485 140.565 214.395 ;
        RECT 139.665 211.950 140.345 213.485 ;
        RECT 138.645 211.790 139.455 211.930 ;
        RECT 138.645 211.620 139.645 211.790 ;
        RECT 138.645 210.560 139.455 211.620 ;
        RECT 139.665 210.600 140.575 211.950 ;
        RECT 138.775 201.670 139.455 210.465 ;
        RECT 139.665 209.535 140.575 210.455 ;
        RECT 139.665 207.190 140.345 209.535 ;
        RECT 139.475 207.020 140.345 207.190 ;
        RECT 139.665 206.990 140.345 207.020 ;
        RECT 139.505 206.615 139.615 206.735 ;
        RECT 139.750 205.970 140.535 206.400 ;
        RECT 139.665 205.535 140.575 205.950 ;
        RECT 139.475 205.365 140.575 205.535 ;
        RECT 139.665 205.020 140.575 205.365 ;
        RECT 139.665 202.050 140.345 205.020 ;
        RECT 139.505 201.670 139.615 201.675 ;
        RECT 138.775 201.500 139.645 201.670 ;
        RECT 138.775 201.360 139.455 201.500 ;
        RECT 138.545 200.335 139.455 201.255 ;
        RECT 139.475 201.205 139.645 201.210 ;
        RECT 139.475 201.040 140.345 201.205 ;
        RECT 138.775 197.990 139.455 200.335 ;
        RECT 139.665 200.300 140.345 201.040 ;
        RECT 139.665 199.370 140.575 200.300 ;
        RECT 139.665 197.990 140.575 199.040 ;
        RECT 138.775 197.820 140.575 197.990 ;
        RECT 138.775 197.790 139.455 197.820 ;
        RECT 139.665 197.690 140.575 197.820 ;
        RECT 138.645 197.530 139.455 197.670 ;
        RECT 139.665 197.530 140.345 197.670 ;
        RECT 138.645 197.360 140.345 197.530 ;
        RECT 138.645 196.300 139.455 197.360 ;
        RECT 138.745 196.145 139.425 196.290 ;
        RECT 138.745 195.975 139.645 196.145 ;
        RECT 138.745 194.485 139.425 195.975 ;
        RECT 138.545 193.540 139.455 194.485 ;
        RECT 139.665 194.155 140.345 197.360 ;
        RECT 138.585 193.090 139.370 193.520 ;
        RECT 139.665 193.245 140.565 194.155 ;
        RECT 138.545 192.930 139.455 192.990 ;
        RECT 138.545 192.760 139.645 192.930 ;
        RECT 138.545 189.540 139.455 192.760 ;
        RECT 139.665 191.710 140.345 193.245 ;
        RECT 139.665 190.360 140.575 191.710 ;
        RECT 139.505 190.055 139.615 190.175 ;
        RECT 139.475 189.705 139.645 189.710 ;
        RECT 139.475 189.540 140.345 189.705 ;
        RECT 138.545 189.250 139.455 189.310 ;
        RECT 138.545 189.080 139.645 189.250 ;
        RECT 138.545 185.860 139.455 189.080 ;
        RECT 139.665 188.800 140.345 189.540 ;
        RECT 139.665 187.870 140.575 188.800 ;
        RECT 139.665 187.410 140.445 187.550 ;
        RECT 139.475 187.240 140.445 187.410 ;
        RECT 139.665 186.180 140.445 187.240 ;
        RECT 139.500 185.400 139.610 185.560 ;
        RECT 139.665 185.120 140.445 186.170 ;
        RECT 139.475 184.950 140.445 185.120 ;
        RECT 139.665 184.800 140.445 184.950 ;
        RECT 138.645 183.730 139.455 184.790 ;
        RECT 139.665 183.730 140.475 184.790 ;
        RECT 138.645 183.560 140.475 183.730 ;
        RECT 138.645 183.420 139.455 183.560 ;
        RECT 139.665 183.420 140.475 183.560 ;
      LAYER nwell ;
        RECT 140.865 183.225 143.695 219.485 ;
      LAYER pwell ;
        RECT 144.085 219.150 144.895 219.290 ;
        RECT 145.105 219.150 145.915 219.290 ;
        RECT 144.085 218.980 145.915 219.150 ;
        RECT 144.085 217.920 144.895 218.980 ;
        RECT 145.105 217.920 145.915 218.980 ;
        RECT 144.085 217.770 144.895 217.910 ;
        RECT 145.105 217.770 145.915 217.910 ;
        RECT 144.085 217.600 145.915 217.770 ;
        RECT 144.085 214.240 144.895 217.600 ;
        RECT 144.945 213.975 145.055 214.095 ;
        RECT 143.985 212.380 144.895 213.730 ;
        RECT 145.105 212.400 145.915 217.600 ;
        RECT 144.215 210.845 144.895 212.380 ;
        RECT 144.950 212.080 145.060 212.240 ;
        RECT 145.105 211.330 145.785 211.470 ;
        RECT 144.915 211.160 145.785 211.330 ;
        RECT 143.995 209.935 144.895 210.845 ;
        RECT 144.215 206.730 144.895 209.935 ;
        RECT 145.105 210.985 145.785 211.160 ;
        RECT 145.105 209.640 146.015 210.985 ;
        RECT 145.105 206.730 146.015 209.500 ;
        RECT 144.215 206.560 146.015 206.730 ;
        RECT 144.215 206.420 144.895 206.560 ;
        RECT 145.105 206.500 146.015 206.560 ;
        RECT 144.215 206.270 144.895 206.410 ;
        RECT 144.215 206.100 145.085 206.270 ;
        RECT 144.215 202.895 144.895 206.100 ;
        RECT 145.190 205.970 145.975 206.400 ;
        RECT 144.950 205.640 145.060 205.800 ;
        RECT 145.105 204.890 145.785 204.920 ;
        RECT 144.915 204.720 145.785 204.890 ;
        RECT 143.995 201.985 144.895 202.895 ;
        RECT 144.215 200.450 144.895 201.985 ;
        RECT 145.105 202.375 145.785 204.720 ;
        RECT 145.105 201.455 146.015 202.375 ;
        RECT 144.950 201.040 145.060 201.200 ;
        RECT 143.985 199.100 144.895 200.450 ;
        RECT 145.105 199.085 146.015 200.430 ;
        RECT 145.105 198.910 145.785 199.085 ;
        RECT 144.915 198.740 145.785 198.910 ;
        RECT 143.985 197.810 144.895 198.740 ;
        RECT 145.105 198.600 145.785 198.740 ;
        RECT 145.105 198.450 145.785 198.480 ;
        RECT 144.915 198.280 145.785 198.450 ;
        RECT 144.215 197.070 144.895 197.810 ;
        RECT 144.215 196.905 145.085 197.070 ;
        RECT 144.915 196.900 145.085 196.905 ;
        RECT 144.215 196.610 144.895 196.750 ;
        RECT 144.215 196.440 145.085 196.610 ;
        RECT 144.215 196.265 144.895 196.440 ;
        RECT 143.985 194.920 144.895 196.265 ;
        RECT 145.105 195.935 145.785 198.280 ;
        RECT 145.105 195.015 146.015 195.935 ;
        RECT 143.985 194.770 144.895 194.900 ;
        RECT 143.985 194.760 145.085 194.770 ;
        RECT 145.105 194.760 145.885 194.910 ;
        RECT 143.985 194.600 145.885 194.760 ;
        RECT 143.985 193.550 144.895 194.600 ;
        RECT 144.915 194.590 145.885 194.600 ;
        RECT 145.105 193.540 145.885 194.590 ;
        RECT 144.025 193.090 144.810 193.520 ;
        RECT 145.190 193.090 145.975 193.520 ;
        RECT 143.985 192.930 144.895 192.990 ;
        RECT 143.985 192.760 145.085 192.930 ;
        RECT 143.985 189.990 144.895 192.760 ;
        RECT 145.105 190.805 146.015 192.150 ;
        RECT 145.105 190.630 145.785 190.805 ;
        RECT 144.915 190.460 145.785 190.630 ;
        RECT 145.105 190.320 145.785 190.460 ;
        RECT 145.105 190.170 145.915 190.310 ;
        RECT 144.915 190.000 145.915 190.170 ;
        RECT 144.215 189.710 144.895 189.740 ;
        RECT 144.215 189.540 145.085 189.710 ;
        RECT 144.215 187.195 144.895 189.540 ;
        RECT 145.105 188.940 145.915 190.000 ;
        RECT 145.105 187.870 145.885 188.930 ;
        RECT 144.915 187.700 145.885 187.870 ;
        RECT 145.105 187.560 145.885 187.700 ;
        RECT 143.985 186.275 144.895 187.195 ;
        RECT 145.105 186.490 145.885 187.550 ;
        RECT 144.915 186.320 145.885 186.490 ;
        RECT 145.105 186.180 145.885 186.320 ;
        RECT 144.115 185.120 144.895 186.170 ;
        RECT 145.105 185.120 145.885 186.170 ;
        RECT 144.115 184.950 145.885 185.120 ;
        RECT 144.115 184.800 144.895 184.950 ;
        RECT 145.105 184.800 145.885 184.950 ;
        RECT 144.085 183.730 144.895 184.790 ;
        RECT 145.105 183.730 145.915 184.790 ;
        RECT 144.085 183.560 145.915 183.730 ;
        RECT 144.085 183.420 144.895 183.560 ;
        RECT 145.105 183.420 145.915 183.560 ;
      LAYER nwell ;
        RECT 146.305 183.225 147.910 219.485 ;
        RECT 11.910 172.445 90.030 174.050 ;
      LAYER pwell ;
        RECT 12.105 171.245 13.475 172.055 ;
        RECT 13.485 171.245 18.995 172.055 ;
        RECT 19.005 171.245 24.515 172.055 ;
        RECT 24.995 171.330 25.425 172.115 ;
        RECT 25.445 171.245 30.955 172.055 ;
        RECT 30.965 171.245 36.475 172.055 ;
        RECT 36.485 171.245 37.855 172.055 ;
        RECT 37.875 171.330 38.305 172.115 ;
        RECT 38.325 171.245 43.835 172.055 ;
        RECT 43.845 171.245 45.675 172.055 ;
        RECT 45.685 171.925 47.030 172.155 ;
        RECT 45.685 171.245 47.515 171.925 ;
        RECT 47.525 171.245 50.275 172.055 ;
        RECT 50.755 171.330 51.185 172.115 ;
        RECT 51.205 171.245 56.715 172.055 ;
        RECT 56.725 171.245 58.095 172.055 ;
        RECT 58.105 171.925 59.450 172.155 ;
        RECT 59.945 171.925 61.290 172.155 ;
        RECT 61.785 171.925 63.130 172.155 ;
        RECT 58.105 171.245 59.935 171.925 ;
        RECT 59.945 171.245 61.775 171.925 ;
        RECT 61.785 171.245 63.615 171.925 ;
        RECT 63.635 171.330 64.065 172.115 ;
        RECT 64.570 171.925 65.915 172.155 ;
        RECT 64.085 171.245 65.915 171.925 ;
        RECT 65.925 171.925 67.270 172.155 ;
        RECT 68.075 171.925 69.005 172.155 ;
        RECT 70.375 171.925 71.305 172.155 ;
        RECT 72.675 171.925 73.605 172.155 ;
        RECT 74.665 171.925 76.010 172.155 ;
        RECT 65.925 171.245 67.755 171.925 ;
        RECT 68.075 171.245 69.910 171.925 ;
        RECT 70.375 171.245 72.210 171.925 ;
        RECT 72.675 171.245 74.510 171.925 ;
        RECT 74.665 171.245 76.495 171.925 ;
        RECT 76.515 171.330 76.945 172.115 ;
        RECT 78.015 171.925 78.945 172.155 ;
        RECT 80.315 171.925 81.245 172.155 ;
        RECT 82.615 171.925 83.545 172.155 ;
        RECT 77.110 171.245 78.945 171.925 ;
        RECT 79.410 171.245 81.245 171.925 ;
        RECT 81.710 171.245 83.545 171.925 ;
        RECT 84.325 171.245 87.535 172.155 ;
        RECT 88.465 171.245 89.835 172.055 ;
        RECT 12.245 171.035 12.415 171.245 ;
        RECT 13.625 171.035 13.795 171.245 ;
        RECT 19.145 171.035 19.315 171.245 ;
        RECT 24.665 171.195 24.835 171.225 ;
        RECT 24.660 171.085 24.835 171.195 ;
        RECT 24.665 171.035 24.835 171.085 ;
        RECT 25.585 171.055 25.755 171.245 ;
        RECT 30.185 171.035 30.355 171.225 ;
        RECT 31.105 171.055 31.275 171.245 ;
        RECT 35.705 171.035 35.875 171.225 ;
        RECT 36.625 171.055 36.795 171.245 ;
        RECT 37.540 171.085 37.660 171.195 ;
        RECT 38.465 171.035 38.635 171.245 ;
        RECT 40.300 171.035 40.470 171.225 ;
        RECT 43.985 171.035 44.155 171.245 ;
        RECT 47.205 171.055 47.375 171.245 ;
        RECT 47.665 171.055 47.835 171.245 ;
        RECT 51.345 171.225 51.515 171.245 ;
        RECT 49.505 171.035 49.675 171.225 ;
        RECT 50.420 171.085 50.540 171.195 ;
        RECT 51.340 171.055 51.515 171.225 ;
        RECT 51.340 171.035 51.510 171.055 ;
        RECT 52.725 171.035 52.895 171.225 ;
        RECT 56.865 171.055 57.035 171.245 ;
        RECT 59.625 171.035 59.795 171.245 ;
        RECT 60.085 171.035 60.255 171.225 ;
        RECT 61.465 171.055 61.635 171.245 ;
        RECT 63.305 171.055 63.475 171.245 ;
        RECT 64.225 171.055 64.395 171.245 ;
        RECT 67.445 171.035 67.615 171.245 ;
        RECT 69.745 171.225 69.910 171.245 ;
        RECT 72.045 171.225 72.210 171.245 ;
        RECT 74.345 171.225 74.510 171.245 ;
        RECT 67.915 171.080 68.075 171.190 ;
        RECT 69.745 171.055 69.915 171.225 ;
        RECT 72.045 171.055 72.215 171.225 ;
        RECT 74.345 171.055 74.515 171.225 ;
        RECT 75.725 171.035 75.895 171.225 ;
        RECT 76.185 171.055 76.355 171.245 ;
        RECT 77.110 171.225 77.275 171.245 ;
        RECT 79.410 171.225 79.575 171.245 ;
        RECT 81.710 171.225 81.875 171.245 ;
        RECT 77.105 171.055 77.280 171.225 ;
        RECT 79.405 171.055 79.575 171.225 ;
        RECT 77.110 171.035 77.280 171.055 ;
        RECT 80.790 171.035 80.960 171.225 ;
        RECT 81.705 171.055 81.875 171.225 ;
        RECT 84.000 171.085 84.120 171.195 ;
        RECT 84.465 171.055 84.635 171.245 ;
        RECT 87.225 171.035 87.395 171.225 ;
        RECT 87.695 171.080 87.855 171.200 ;
        RECT 89.525 171.035 89.695 171.245 ;
        RECT 12.105 170.225 13.475 171.035 ;
        RECT 13.485 170.225 18.995 171.035 ;
        RECT 19.005 170.225 24.515 171.035 ;
        RECT 24.525 170.225 30.035 171.035 ;
        RECT 30.045 170.225 35.555 171.035 ;
        RECT 35.565 170.225 37.395 171.035 ;
        RECT 37.875 170.165 38.305 170.950 ;
        RECT 38.325 170.225 40.155 171.035 ;
        RECT 40.175 170.125 43.835 171.035 ;
        RECT 43.845 170.225 49.355 171.035 ;
        RECT 49.365 170.225 51.195 171.035 ;
        RECT 51.225 170.125 52.575 171.035 ;
        RECT 52.585 170.225 58.095 171.035 ;
        RECT 58.105 170.355 59.935 171.035 ;
        RECT 60.055 170.355 63.520 171.035 ;
        RECT 58.105 170.125 59.450 170.355 ;
        RECT 62.600 170.125 63.520 170.355 ;
        RECT 63.635 170.165 64.065 170.950 ;
        RECT 64.180 170.355 67.645 171.035 ;
        RECT 68.725 170.355 76.035 171.035 ;
        RECT 64.180 170.125 65.100 170.355 ;
        RECT 68.725 170.125 70.075 170.355 ;
        RECT 71.610 170.135 72.520 170.355 ;
        RECT 76.965 170.125 80.440 171.035 ;
        RECT 80.645 170.125 84.120 171.035 ;
        RECT 84.325 170.125 87.535 171.035 ;
        RECT 88.465 170.225 89.835 171.035 ;
      LAYER nwell ;
        RECT 11.910 167.005 90.030 169.835 ;
      LAYER pwell ;
        RECT 100.450 167.190 106.550 176.980 ;
        RECT 100.450 167.160 106.560 167.190 ;
        RECT 100.650 166.760 101.810 167.160 ;
        RECT 12.105 165.805 13.475 166.615 ;
        RECT 13.485 165.805 18.995 166.615 ;
        RECT 19.005 165.805 24.515 166.615 ;
        RECT 24.995 165.890 25.425 166.675 ;
        RECT 25.445 165.805 30.955 166.615 ;
        RECT 30.965 165.805 36.475 166.615 ;
        RECT 36.485 165.805 38.315 166.615 ;
        RECT 42.300 166.485 43.210 166.705 ;
        RECT 44.745 166.485 46.095 166.715 ;
        RECT 38.785 165.805 46.095 166.485 ;
        RECT 46.455 166.485 47.385 166.715 ;
        RECT 46.455 165.805 48.290 166.485 ;
        RECT 48.445 165.805 50.275 166.715 ;
        RECT 50.755 165.890 51.185 166.675 ;
        RECT 51.300 166.485 52.220 166.715 ;
        RECT 58.400 166.485 59.310 166.705 ;
        RECT 60.845 166.485 62.195 166.715 ;
        RECT 51.300 165.805 54.765 166.485 ;
        RECT 54.885 165.805 62.195 166.485 ;
        RECT 62.245 166.485 63.175 166.715 ;
        RECT 67.345 166.485 68.695 166.715 ;
        RECT 70.230 166.485 71.140 166.705 ;
        RECT 75.150 166.485 76.495 166.715 ;
        RECT 62.245 165.805 66.145 166.485 ;
        RECT 67.345 165.805 74.655 166.485 ;
        RECT 74.665 165.805 76.495 166.485 ;
        RECT 76.515 165.890 76.945 166.675 ;
        RECT 80.480 166.485 81.390 166.705 ;
        RECT 82.925 166.485 84.275 166.715 ;
        RECT 76.965 165.805 84.275 166.485 ;
        RECT 84.785 165.805 87.995 166.715 ;
        RECT 88.465 165.805 89.835 166.615 ;
        RECT 12.245 165.595 12.415 165.805 ;
        RECT 13.625 165.595 13.795 165.805 ;
        RECT 19.145 165.595 19.315 165.805 ;
        RECT 24.665 165.755 24.835 165.785 ;
        RECT 24.660 165.645 24.835 165.755 ;
        RECT 24.665 165.595 24.835 165.645 ;
        RECT 25.585 165.615 25.755 165.805 ;
        RECT 30.185 165.595 30.355 165.785 ;
        RECT 31.105 165.615 31.275 165.805 ;
        RECT 35.705 165.595 35.875 165.785 ;
        RECT 36.625 165.615 36.795 165.805 ;
        RECT 38.465 165.755 38.635 165.785 ;
        RECT 37.540 165.645 37.660 165.755 ;
        RECT 38.460 165.645 38.635 165.755 ;
        RECT 38.465 165.595 38.635 165.645 ;
        RECT 38.925 165.615 39.095 165.805 ;
        RECT 48.125 165.785 48.290 165.805 ;
        RECT 43.525 165.595 43.695 165.785 ;
        RECT 43.990 165.595 44.160 165.785 ;
        RECT 47.665 165.595 47.835 165.785 ;
        RECT 48.125 165.615 48.295 165.785 ;
        RECT 49.960 165.615 50.130 165.805 ;
        RECT 50.420 165.645 50.540 165.755 ;
        RECT 54.565 165.615 54.735 165.805 ;
        RECT 55.025 165.595 55.195 165.805 ;
        RECT 62.385 165.595 62.555 165.785 ;
        RECT 62.660 165.615 62.830 165.805 ;
        RECT 66.535 165.650 66.695 165.760 ;
        RECT 71.125 165.595 71.295 165.785 ;
        RECT 73.885 165.595 74.055 165.785 ;
        RECT 74.345 165.595 74.515 165.805 ;
        RECT 74.805 165.615 74.975 165.805 ;
        RECT 77.105 165.615 77.275 165.805 ;
        RECT 81.705 165.615 81.875 165.785 ;
        RECT 84.460 165.645 84.580 165.755 ;
        RECT 84.925 165.615 85.095 165.805 ;
        RECT 88.170 165.755 88.340 165.785 ;
        RECT 88.140 165.645 88.340 165.755 ;
        RECT 88.170 165.615 88.340 165.645 ;
        RECT 81.710 165.595 81.875 165.615 ;
        RECT 88.170 165.595 88.280 165.615 ;
        RECT 89.525 165.595 89.695 165.805 ;
        RECT 12.105 164.785 13.475 165.595 ;
        RECT 13.485 164.785 18.995 165.595 ;
        RECT 19.005 164.785 24.515 165.595 ;
        RECT 24.525 164.785 30.035 165.595 ;
        RECT 30.045 164.785 35.555 165.595 ;
        RECT 35.565 164.785 37.395 165.595 ;
        RECT 37.875 164.725 38.305 165.510 ;
        RECT 38.325 164.785 40.155 165.595 ;
        RECT 40.260 164.915 43.725 165.595 ;
        RECT 43.845 164.915 47.430 165.595 ;
        RECT 47.525 164.915 54.835 165.595 ;
        RECT 54.885 164.915 62.195 165.595 ;
        RECT 40.260 164.685 41.180 164.915 ;
        RECT 43.845 164.685 44.765 164.915 ;
        RECT 51.040 164.695 51.950 164.915 ;
        RECT 53.485 164.685 54.835 164.915 ;
        RECT 58.400 164.695 59.310 164.915 ;
        RECT 60.845 164.685 62.195 164.915 ;
        RECT 62.245 164.785 63.615 165.595 ;
        RECT 63.635 164.725 64.065 165.510 ;
        RECT 64.125 164.915 71.435 165.595 ;
        RECT 71.455 164.915 74.195 165.595 ;
        RECT 74.205 164.915 81.515 165.595 ;
        RECT 81.710 164.915 83.545 165.595 ;
        RECT 64.125 164.685 65.475 164.915 ;
        RECT 67.010 164.695 67.920 164.915 ;
        RECT 77.720 164.695 78.630 164.915 ;
        RECT 80.165 164.685 81.515 164.915 ;
        RECT 82.615 164.685 83.545 164.915 ;
        RECT 83.865 164.915 88.280 165.595 ;
        RECT 83.865 164.685 87.795 164.915 ;
        RECT 88.465 164.785 89.835 165.595 ;
        RECT 103.770 165.080 106.560 167.160 ;
      LAYER nwell ;
        RECT 11.910 161.565 90.030 164.395 ;
        RECT 101.660 162.970 106.500 165.080 ;
        RECT 107.780 164.740 117.970 176.990 ;
      LAYER pwell ;
        RECT 120.330 167.140 126.430 176.930 ;
        RECT 120.330 167.110 126.440 167.140 ;
        RECT 120.530 166.710 121.690 167.110 ;
        RECT 123.650 165.030 126.440 167.110 ;
      LAYER nwell ;
        RECT 121.540 162.920 126.380 165.030 ;
        RECT 127.660 164.690 137.850 176.940 ;
      LAYER pwell ;
        RECT 140.360 167.190 146.460 176.980 ;
        RECT 140.360 167.160 146.470 167.190 ;
        RECT 140.560 166.760 141.720 167.160 ;
        RECT 143.680 165.080 146.470 167.160 ;
      LAYER nwell ;
        RECT 141.570 162.970 146.410 165.080 ;
        RECT 147.690 164.740 157.880 176.990 ;
      LAYER pwell ;
        RECT 12.105 160.365 13.475 161.175 ;
        RECT 13.485 160.365 18.995 161.175 ;
        RECT 19.005 160.365 24.515 161.175 ;
        RECT 24.995 160.450 25.425 161.235 ;
        RECT 25.445 160.365 30.955 161.175 ;
        RECT 30.965 160.365 36.475 161.175 ;
        RECT 36.985 161.045 38.335 161.275 ;
        RECT 39.870 161.045 40.780 161.265 ;
        RECT 45.445 161.185 46.395 161.275 ;
        RECT 36.985 160.365 44.295 161.045 ;
        RECT 44.465 160.365 46.395 161.185 ;
        RECT 46.775 160.365 50.275 161.275 ;
        RECT 50.755 160.450 51.185 161.235 ;
        RECT 51.205 160.365 54.415 161.275 ;
        RECT 54.425 161.075 55.370 161.275 ;
        RECT 54.425 160.395 57.175 161.075 ;
        RECT 57.185 161.045 58.115 161.275 ;
        RECT 64.840 161.045 65.750 161.265 ;
        RECT 67.285 161.045 68.635 161.275 ;
        RECT 54.425 160.365 55.370 160.395 ;
        RECT 12.245 160.155 12.415 160.365 ;
        RECT 13.625 160.155 13.795 160.365 ;
        RECT 19.145 160.155 19.315 160.365 ;
        RECT 24.665 160.315 24.835 160.345 ;
        RECT 24.660 160.205 24.835 160.315 ;
        RECT 24.665 160.155 24.835 160.205 ;
        RECT 25.585 160.175 25.755 160.365 ;
        RECT 30.185 160.155 30.355 160.345 ;
        RECT 31.105 160.175 31.275 160.365 ;
        RECT 33.860 160.155 34.030 160.345 ;
        RECT 35.245 160.155 35.415 160.345 ;
        RECT 36.620 160.205 36.740 160.315 ;
        RECT 38.465 160.155 38.635 160.345 ;
        RECT 43.985 160.175 44.155 160.365 ;
        RECT 44.465 160.345 44.615 160.365 ;
        RECT 46.775 160.345 46.910 160.365 ;
        RECT 44.445 160.175 44.615 160.345 ;
        RECT 45.820 160.205 45.940 160.315 ;
        RECT 46.285 160.155 46.455 160.345 ;
        RECT 46.740 160.175 46.910 160.345 ;
        RECT 50.420 160.205 50.540 160.315 ;
        RECT 51.335 160.175 51.505 160.365 ;
        RECT 12.105 159.345 13.475 160.155 ;
        RECT 13.485 159.345 18.995 160.155 ;
        RECT 19.005 159.345 24.515 160.155 ;
        RECT 24.525 159.345 30.035 160.155 ;
        RECT 30.045 159.345 33.715 160.155 ;
        RECT 33.745 159.245 35.095 160.155 ;
        RECT 35.115 159.245 37.845 160.155 ;
        RECT 37.875 159.285 38.305 160.070 ;
        RECT 38.325 159.475 45.635 160.155 ;
        RECT 46.145 159.475 53.455 160.155 ;
        RECT 53.650 160.125 53.820 160.345 ;
        RECT 56.860 160.175 57.030 160.395 ;
        RECT 57.185 160.365 61.085 161.045 ;
        RECT 61.325 160.365 68.635 161.045 ;
        RECT 68.685 161.045 69.615 161.275 ;
        RECT 72.920 161.045 73.840 161.275 ;
        RECT 68.685 160.365 72.585 161.045 ;
        RECT 72.920 160.365 76.385 161.045 ;
        RECT 76.515 160.450 76.945 161.235 ;
        RECT 76.965 160.365 80.440 161.275 ;
        RECT 84.620 161.045 85.530 161.265 ;
        RECT 87.065 161.045 88.415 161.275 ;
        RECT 81.105 160.365 88.415 161.045 ;
        RECT 88.465 160.365 89.835 161.175 ;
        RECT 57.600 160.175 57.770 160.365 ;
        RECT 56.225 160.125 57.175 160.155 ;
        RECT 41.840 159.255 42.750 159.475 ;
        RECT 44.285 159.245 45.635 159.475 ;
        RECT 49.660 159.255 50.570 159.475 ;
        RECT 52.105 159.245 53.455 159.475 ;
        RECT 53.505 159.445 57.175 160.125 ;
        RECT 56.225 159.245 57.175 159.445 ;
        RECT 57.185 160.125 58.120 160.155 ;
        RECT 60.080 160.125 60.250 160.345 ;
        RECT 61.465 160.175 61.635 160.365 ;
        RECT 62.845 160.155 63.015 160.345 ;
        RECT 63.300 160.205 63.420 160.315 ;
        RECT 64.500 160.155 64.670 160.345 ;
        RECT 68.640 160.155 68.810 160.345 ;
        RECT 69.100 160.175 69.270 160.365 ;
        RECT 76.185 160.345 76.355 160.365 ;
        RECT 75.725 160.155 75.895 160.345 ;
        RECT 76.185 160.175 76.360 160.345 ;
        RECT 77.110 160.175 77.280 160.365 ;
        RECT 80.785 160.315 80.955 160.345 ;
        RECT 80.780 160.205 80.955 160.315 ;
        RECT 76.190 160.155 76.360 160.175 ;
        RECT 80.785 160.155 80.955 160.205 ;
        RECT 81.245 160.155 81.415 160.365 ;
        RECT 89.525 160.155 89.695 160.365 ;
        RECT 57.185 159.925 60.250 160.125 ;
        RECT 57.185 159.445 60.395 159.925 ;
        RECT 57.185 159.245 58.135 159.445 ;
        RECT 59.465 159.245 60.395 159.445 ;
        RECT 60.405 159.475 63.155 160.155 ;
        RECT 60.405 159.245 61.335 159.475 ;
        RECT 63.635 159.285 64.065 160.070 ;
        RECT 64.085 159.475 67.985 160.155 ;
        RECT 68.225 159.475 72.125 160.155 ;
        RECT 72.460 159.475 75.925 160.155 ;
        RECT 64.085 159.245 65.015 159.475 ;
        RECT 68.225 159.245 69.155 159.475 ;
        RECT 72.460 159.245 73.380 159.475 ;
        RECT 76.045 159.245 79.520 160.155 ;
        RECT 79.725 159.375 81.095 160.155 ;
        RECT 81.105 159.475 88.415 160.155 ;
        RECT 84.620 159.255 85.530 159.475 ;
        RECT 87.065 159.245 88.415 159.475 ;
        RECT 88.465 159.345 89.835 160.155 ;
      LAYER nwell ;
        RECT 11.910 156.125 90.030 158.955 ;
      LAYER pwell ;
        RECT 12.105 154.925 13.475 155.735 ;
        RECT 13.485 154.925 18.995 155.735 ;
        RECT 19.005 154.925 24.515 155.735 ;
        RECT 24.995 155.010 25.425 155.795 ;
        RECT 25.445 154.925 30.955 155.735 ;
        RECT 30.965 154.925 34.635 155.735 ;
        RECT 35.105 155.635 36.060 155.835 ;
        RECT 35.105 154.955 37.385 155.635 ;
        RECT 38.455 155.605 39.385 155.835 ;
        RECT 35.105 154.925 36.060 154.955 ;
        RECT 12.245 154.715 12.415 154.925 ;
        RECT 13.625 154.715 13.795 154.925 ;
        RECT 19.145 154.715 19.315 154.925 ;
        RECT 24.665 154.875 24.835 154.905 ;
        RECT 24.660 154.765 24.835 154.875 ;
        RECT 24.665 154.715 24.835 154.765 ;
        RECT 25.585 154.735 25.755 154.925 ;
        RECT 30.185 154.715 30.355 154.905 ;
        RECT 31.105 154.735 31.275 154.925 ;
        RECT 34.780 154.765 34.900 154.875 ;
        RECT 35.705 154.715 35.875 154.905 ;
        RECT 37.090 154.735 37.260 154.955 ;
        RECT 37.550 154.925 39.385 155.605 ;
        RECT 39.705 155.635 40.650 155.835 ;
        RECT 41.985 155.635 42.915 155.835 ;
        RECT 39.705 155.155 42.915 155.635 ;
        RECT 43.020 155.605 43.940 155.835 ;
        RECT 49.260 155.605 50.180 155.835 ;
        RECT 39.705 154.955 42.775 155.155 ;
        RECT 39.705 154.925 40.650 154.955 ;
        RECT 37.550 154.905 37.715 154.925 ;
        RECT 37.545 154.875 37.715 154.905 ;
        RECT 37.540 154.765 37.715 154.875 ;
        RECT 37.545 154.735 37.715 154.765 ;
        RECT 38.475 154.760 38.635 154.870 ;
        RECT 39.390 154.715 39.560 154.905 ;
        RECT 42.605 154.875 42.775 154.955 ;
        RECT 43.020 154.925 46.485 155.605 ;
        RECT 46.715 154.925 50.180 155.605 ;
        RECT 50.755 155.010 51.185 155.795 ;
        RECT 51.205 154.925 52.555 155.835 ;
        RECT 52.585 154.925 56.060 155.835 ;
        RECT 56.265 155.635 57.215 155.835 ;
        RECT 58.545 155.635 59.475 155.835 ;
        RECT 56.265 155.155 59.475 155.635 ;
        RECT 59.485 155.605 60.415 155.835 ;
        RECT 56.265 154.955 59.330 155.155 ;
        RECT 56.265 154.925 57.200 154.955 ;
        RECT 42.600 154.765 42.775 154.875 ;
        RECT 42.605 154.735 42.775 154.765 ;
        RECT 46.285 154.735 46.455 154.925 ;
        RECT 46.745 154.735 46.915 154.925 ;
        RECT 49.965 154.715 50.135 154.905 ;
        RECT 50.425 154.875 50.595 154.905 ;
        RECT 50.420 154.765 50.595 154.875 ;
        RECT 50.425 154.715 50.595 154.765 ;
        RECT 52.270 154.735 52.440 154.925 ;
        RECT 52.730 154.735 52.900 154.925 ;
        RECT 53.195 154.760 53.355 154.870 ;
        RECT 54.105 154.715 54.275 154.905 ;
        RECT 59.160 154.735 59.330 154.955 ;
        RECT 59.485 154.925 62.235 155.605 ;
        RECT 62.245 154.925 65.455 155.835 ;
        RECT 65.465 155.605 66.395 155.835 ;
        RECT 69.605 155.605 70.535 155.835 ;
        RECT 75.255 155.605 76.185 155.835 ;
        RECT 65.465 154.925 69.365 155.605 ;
        RECT 69.605 154.925 73.505 155.605 ;
        RECT 74.350 154.925 76.185 155.605 ;
        RECT 76.515 155.010 76.945 155.795 ;
        RECT 77.060 155.605 77.980 155.835 ;
        RECT 77.060 154.925 80.525 155.605 ;
        RECT 80.645 154.925 84.120 155.835 ;
        RECT 84.325 154.925 87.800 155.835 ;
        RECT 88.465 154.925 89.835 155.735 ;
        RECT 61.925 154.735 62.095 154.925 ;
        RECT 62.375 154.735 62.545 154.925 ;
        RECT 63.305 154.715 63.475 154.905 ;
        RECT 65.880 154.735 66.050 154.925 ;
        RECT 67.445 154.715 67.615 154.905 ;
        RECT 67.905 154.715 68.075 154.905 ;
        RECT 70.020 154.735 70.190 154.925 ;
        RECT 74.350 154.905 74.515 154.925 ;
        RECT 73.880 154.765 74.000 154.875 ;
        RECT 74.345 154.735 74.515 154.905 ;
        RECT 78.485 154.715 78.655 154.905 ;
        RECT 78.935 154.715 79.105 154.905 ;
        RECT 80.325 154.735 80.495 154.925 ;
        RECT 80.790 154.735 80.960 154.925 ;
        RECT 82.165 154.715 82.335 154.905 ;
        RECT 83.995 154.715 84.165 154.905 ;
        RECT 84.470 154.735 84.640 154.925 ;
        RECT 88.135 154.715 88.305 154.905 ;
        RECT 89.525 154.715 89.695 154.925 ;
        RECT 12.105 153.905 13.475 154.715 ;
        RECT 13.485 153.905 18.995 154.715 ;
        RECT 19.005 153.905 24.515 154.715 ;
        RECT 24.525 153.905 30.035 154.715 ;
        RECT 30.045 153.905 35.555 154.715 ;
        RECT 35.565 153.905 37.395 154.715 ;
        RECT 37.875 153.845 38.305 154.630 ;
        RECT 39.245 153.805 42.165 154.715 ;
        RECT 42.965 154.035 50.275 154.715 ;
        RECT 42.965 153.805 44.315 154.035 ;
        RECT 45.850 153.815 46.760 154.035 ;
        RECT 50.295 153.805 53.025 154.715 ;
        RECT 53.965 154.035 61.275 154.715 ;
        RECT 57.480 153.815 58.390 154.035 ;
        RECT 59.925 153.805 61.275 154.035 ;
        RECT 61.325 154.035 63.615 154.715 ;
        RECT 61.325 153.805 62.245 154.035 ;
        RECT 63.635 153.845 64.065 154.630 ;
        RECT 64.180 154.035 67.645 154.715 ;
        RECT 67.765 154.035 75.075 154.715 ;
        RECT 64.180 153.805 65.100 154.035 ;
        RECT 71.280 153.815 72.190 154.035 ;
        RECT 73.725 153.805 75.075 154.035 ;
        RECT 75.220 154.035 78.685 154.715 ;
        RECT 75.220 153.805 76.140 154.035 ;
        RECT 78.805 153.805 82.015 154.715 ;
        RECT 82.025 154.035 83.855 154.715 ;
        RECT 82.510 153.805 83.855 154.035 ;
        RECT 83.865 153.805 87.075 154.715 ;
        RECT 87.085 153.935 88.455 154.715 ;
        RECT 88.465 153.905 89.835 154.715 ;
      LAYER nwell ;
        RECT 11.910 150.685 90.030 153.515 ;
      LAYER pwell ;
        RECT 100.450 152.190 106.550 161.980 ;
        RECT 100.450 152.160 106.560 152.190 ;
        RECT 100.650 151.760 101.810 152.160 ;
        RECT 12.105 149.485 13.475 150.295 ;
        RECT 13.485 149.485 18.995 150.295 ;
        RECT 19.005 149.485 22.675 150.295 ;
        RECT 23.145 149.485 24.975 150.165 ;
        RECT 24.995 149.570 25.425 150.355 ;
        RECT 25.445 149.485 30.955 150.295 ;
        RECT 30.965 149.485 36.475 150.295 ;
        RECT 36.485 149.485 40.155 150.295 ;
        RECT 40.175 149.485 41.525 150.395 ;
        RECT 41.545 149.485 42.895 150.395 ;
        RECT 42.925 149.485 44.295 150.295 ;
        RECT 44.400 150.165 45.320 150.395 ;
        RECT 44.400 149.485 47.865 150.165 ;
        RECT 47.985 149.485 49.355 150.295 ;
        RECT 49.385 149.485 50.735 150.395 ;
        RECT 50.755 149.570 51.185 150.355 ;
        RECT 52.575 150.165 53.495 150.395 ;
        RECT 51.205 149.485 53.495 150.165 ;
        RECT 53.505 149.485 55.335 150.295 ;
        RECT 55.345 150.165 56.690 150.395 ;
        RECT 57.185 150.165 58.115 150.395 ;
        RECT 55.345 149.485 57.175 150.165 ;
        RECT 57.185 149.485 61.085 150.165 ;
        RECT 61.325 149.485 63.415 150.295 ;
        RECT 67.200 150.165 68.120 150.395 ;
        RECT 71.740 150.165 72.650 150.385 ;
        RECT 74.185 150.165 75.535 150.395 ;
        RECT 64.655 149.485 68.120 150.165 ;
        RECT 68.225 149.485 75.535 150.165 ;
        RECT 76.515 149.570 76.945 150.355 ;
        RECT 77.160 149.485 80.635 150.395 ;
        RECT 84.620 150.165 85.530 150.385 ;
        RECT 87.065 150.165 88.415 150.395 ;
        RECT 81.105 149.485 88.415 150.165 ;
        RECT 88.465 149.485 89.835 150.295 ;
        RECT 103.770 150.080 106.560 152.160 ;
        RECT 12.245 149.275 12.415 149.485 ;
        RECT 13.625 149.275 13.795 149.485 ;
        RECT 19.145 149.275 19.315 149.485 ;
        RECT 20.525 149.275 20.695 149.465 ;
        RECT 22.820 149.325 22.940 149.435 ;
        RECT 24.665 149.295 24.835 149.485 ;
        RECT 25.585 149.295 25.755 149.485 ;
        RECT 27.890 149.275 28.060 149.465 ;
        RECT 29.265 149.275 29.435 149.465 ;
        RECT 31.105 149.295 31.275 149.485 ;
        RECT 34.785 149.275 34.955 149.465 ;
        RECT 36.625 149.295 36.795 149.485 ;
        RECT 40.305 149.465 40.475 149.485 ;
        RECT 37.540 149.325 37.660 149.435 ;
        RECT 38.465 149.275 38.635 149.465 ;
        RECT 40.300 149.295 40.475 149.465 ;
        RECT 40.300 149.275 40.470 149.295 ;
        RECT 41.690 149.275 41.860 149.465 ;
        RECT 42.610 149.295 42.780 149.485 ;
        RECT 43.065 149.295 43.235 149.485 ;
        RECT 47.205 149.295 47.375 149.465 ;
        RECT 47.665 149.295 47.835 149.485 ;
        RECT 48.125 149.295 48.295 149.485 ;
        RECT 47.205 149.275 47.370 149.295 ;
        RECT 48.575 149.275 48.745 149.465 ;
        RECT 49.045 149.275 49.215 149.465 ;
        RECT 50.420 149.295 50.590 149.485 ;
        RECT 50.700 149.275 50.870 149.465 ;
        RECT 51.345 149.295 51.515 149.485 ;
        RECT 53.645 149.295 53.815 149.485 ;
        RECT 54.565 149.275 54.735 149.465 ;
        RECT 56.865 149.295 57.035 149.485 ;
        RECT 57.600 149.295 57.770 149.485 ;
        RECT 58.245 149.275 58.415 149.465 ;
        RECT 59.900 149.275 60.070 149.465 ;
        RECT 61.465 149.295 61.635 149.485 ;
        RECT 64.220 149.325 64.340 149.435 ;
        RECT 64.685 149.295 64.855 149.485 ;
        RECT 68.365 149.295 68.535 149.485 ;
        RECT 71.125 149.275 71.295 149.465 ;
        RECT 71.860 149.275 72.030 149.465 ;
        RECT 75.735 149.330 75.895 149.440 ;
        RECT 78.945 149.275 79.115 149.465 ;
        RECT 80.320 149.295 80.490 149.485 ;
        RECT 80.780 149.325 80.900 149.435 ;
        RECT 81.245 149.295 81.415 149.485 ;
        RECT 82.625 149.275 82.795 149.465 ;
        RECT 83.090 149.275 83.260 149.465 ;
        RECT 86.765 149.275 86.935 149.465 ;
        RECT 89.525 149.275 89.695 149.485 ;
        RECT 12.105 148.465 13.475 149.275 ;
        RECT 13.485 148.465 18.995 149.275 ;
        RECT 19.005 148.465 20.375 149.275 ;
        RECT 20.385 148.595 27.695 149.275 ;
        RECT 23.900 148.375 24.810 148.595 ;
        RECT 26.345 148.365 27.695 148.595 ;
        RECT 27.745 148.365 29.095 149.275 ;
        RECT 29.125 148.465 34.635 149.275 ;
        RECT 34.645 148.465 37.395 149.275 ;
        RECT 37.875 148.405 38.305 149.190 ;
        RECT 38.325 148.465 40.155 149.275 ;
        RECT 40.185 148.365 41.535 149.275 ;
        RECT 41.545 148.595 45.130 149.275 ;
        RECT 45.535 148.595 47.370 149.275 ;
        RECT 41.545 148.365 42.465 148.595 ;
        RECT 45.535 148.365 46.465 148.595 ;
        RECT 47.525 148.495 48.895 149.275 ;
        RECT 48.905 148.465 50.275 149.275 ;
        RECT 50.285 148.595 54.185 149.275 ;
        RECT 50.285 148.365 51.215 148.595 ;
        RECT 54.425 148.465 58.095 149.275 ;
        RECT 58.105 148.465 59.475 149.275 ;
        RECT 59.485 148.595 63.385 149.275 ;
        RECT 59.485 148.365 60.415 148.595 ;
        RECT 63.635 148.405 64.065 149.190 ;
        RECT 64.125 148.595 71.435 149.275 ;
        RECT 71.445 148.595 75.345 149.275 ;
        RECT 75.680 148.595 79.145 149.275 ;
        RECT 79.360 148.595 82.825 149.275 ;
        RECT 64.125 148.365 65.475 148.595 ;
        RECT 67.010 148.375 67.920 148.595 ;
        RECT 71.445 148.365 72.375 148.595 ;
        RECT 75.680 148.365 76.600 148.595 ;
        RECT 79.360 148.365 80.280 148.595 ;
        RECT 82.945 148.365 86.420 149.275 ;
        RECT 86.625 148.595 88.455 149.275 ;
        RECT 87.110 148.365 88.455 148.595 ;
        RECT 88.465 148.465 89.835 149.275 ;
      LAYER nwell ;
        RECT 11.910 145.245 90.030 148.075 ;
        RECT 101.660 147.970 106.500 150.080 ;
        RECT 107.780 149.740 117.970 161.990 ;
      LAYER pwell ;
        RECT 120.330 152.190 126.430 161.980 ;
        RECT 120.330 152.160 126.440 152.190 ;
        RECT 120.530 151.760 121.690 152.160 ;
        RECT 123.650 150.080 126.440 152.160 ;
      LAYER nwell ;
        RECT 121.540 147.970 126.380 150.080 ;
        RECT 127.660 149.740 137.850 161.990 ;
      LAYER pwell ;
        RECT 140.410 152.140 146.510 161.930 ;
        RECT 140.410 152.110 146.520 152.140 ;
        RECT 140.610 151.710 141.770 152.110 ;
        RECT 143.730 150.030 146.520 152.110 ;
      LAYER nwell ;
        RECT 141.620 147.920 146.460 150.030 ;
        RECT 147.740 149.690 157.930 161.940 ;
      LAYER pwell ;
        RECT 12.105 144.045 13.475 144.855 ;
        RECT 13.485 144.045 16.235 144.855 ;
        RECT 20.220 144.725 21.130 144.945 ;
        RECT 22.665 144.725 24.015 144.955 ;
        RECT 16.705 144.045 24.015 144.725 ;
        RECT 24.995 144.130 25.425 144.915 ;
        RECT 25.445 144.045 26.795 144.955 ;
        RECT 30.340 144.725 31.250 144.945 ;
        RECT 32.785 144.725 34.135 144.955 ;
        RECT 37.700 144.725 38.610 144.945 ;
        RECT 40.145 144.725 41.495 144.955 ;
        RECT 26.825 144.045 34.135 144.725 ;
        RECT 34.185 144.045 41.495 144.725 ;
        RECT 41.640 144.725 42.560 144.955 ;
        RECT 41.640 144.045 45.105 144.725 ;
        RECT 45.225 144.045 47.055 144.855 ;
        RECT 47.160 144.725 48.080 144.955 ;
        RECT 47.160 144.045 50.625 144.725 ;
        RECT 50.755 144.130 51.185 144.915 ;
        RECT 51.205 144.045 52.555 144.955 ;
        RECT 52.585 144.045 54.415 144.855 ;
        RECT 57.940 144.725 58.850 144.945 ;
        RECT 60.385 144.725 61.735 144.955 ;
        RECT 54.425 144.045 61.735 144.725 ;
        RECT 62.245 144.725 63.590 144.955 ;
        RECT 67.285 144.725 68.215 144.955 ;
        RECT 62.245 144.045 64.075 144.725 ;
        RECT 64.315 144.045 68.215 144.725 ;
        RECT 68.225 144.725 69.155 144.955 ;
        RECT 72.365 144.725 73.295 144.955 ;
        RECT 68.225 144.045 72.125 144.725 ;
        RECT 72.365 144.045 76.265 144.725 ;
        RECT 76.515 144.130 76.945 144.915 ;
        RECT 80.480 144.725 81.390 144.945 ;
        RECT 82.925 144.725 84.275 144.955 ;
        RECT 76.965 144.045 84.275 144.725 ;
        RECT 84.325 144.045 87.800 144.955 ;
        RECT 88.465 144.045 89.835 144.855 ;
        RECT 12.245 143.835 12.415 144.045 ;
        RECT 13.625 143.995 13.795 144.045 ;
        RECT 13.620 143.885 13.795 143.995 ;
        RECT 13.625 143.855 13.795 143.885 ;
        RECT 15.000 143.835 15.170 144.025 ;
        RECT 15.465 143.835 15.635 144.025 ;
        RECT 16.380 143.885 16.500 143.995 ;
        RECT 16.845 143.855 17.015 144.045 ;
        RECT 19.145 143.835 19.315 144.025 ;
        RECT 22.825 143.835 22.995 144.025 ;
        RECT 24.215 143.890 24.375 144.000 ;
        RECT 25.590 143.855 25.760 144.045 ;
        RECT 26.965 143.855 27.135 144.045 ;
        RECT 30.185 143.835 30.355 144.025 ;
        RECT 34.325 143.855 34.495 144.045 ;
        RECT 38.465 143.835 38.635 144.025 ;
        RECT 44.905 143.855 45.075 144.045 ;
        RECT 45.365 143.855 45.535 144.045 ;
        RECT 45.835 143.880 45.995 143.990 ;
        RECT 46.745 143.835 46.915 144.025 ;
        RECT 50.425 143.855 50.595 144.045 ;
        RECT 51.350 143.855 51.520 144.045 ;
        RECT 52.725 143.855 52.895 144.045 ;
        RECT 54.100 143.885 54.220 143.995 ;
        RECT 54.565 143.855 54.735 144.045 ;
        RECT 54.840 143.835 55.010 144.025 ;
        RECT 61.925 143.995 62.095 144.025 ;
        RECT 61.920 143.885 62.095 143.995 ;
        RECT 61.925 143.835 62.095 143.885 ;
        RECT 62.385 143.835 62.555 144.025 ;
        RECT 63.765 143.855 63.935 144.045 ;
        RECT 67.630 143.855 67.800 144.045 ;
        RECT 68.640 143.855 68.810 144.045 ;
        RECT 68.825 143.835 68.995 144.025 ;
        RECT 69.560 143.835 69.730 144.025 ;
        RECT 72.780 143.855 72.950 144.045 ;
        RECT 73.420 143.885 73.540 143.995 ;
        RECT 77.105 143.855 77.275 144.045 ;
        RECT 80.785 143.835 80.955 144.025 ;
        RECT 81.245 143.835 81.415 144.025 ;
        RECT 84.470 143.855 84.640 144.045 ;
        RECT 88.140 143.885 88.260 143.995 ;
        RECT 89.525 143.835 89.695 144.045 ;
        RECT 12.105 143.025 13.475 143.835 ;
        RECT 13.965 142.925 15.315 143.835 ;
        RECT 15.325 143.155 18.995 143.835 ;
        RECT 19.005 143.155 22.675 143.835 ;
        RECT 22.685 143.155 29.995 143.835 ;
        RECT 30.045 143.155 37.775 143.835 ;
        RECT 18.065 142.925 18.995 143.155 ;
        RECT 21.745 142.925 22.675 143.155 ;
        RECT 26.200 142.935 27.110 143.155 ;
        RECT 28.645 142.925 29.995 143.155 ;
        RECT 33.560 142.935 34.470 143.155 ;
        RECT 36.005 142.925 37.775 143.155 ;
        RECT 37.875 142.965 38.305 143.750 ;
        RECT 38.325 143.155 45.635 143.835 ;
        RECT 46.605 143.155 53.915 143.835 ;
        RECT 41.840 142.935 42.750 143.155 ;
        RECT 44.285 142.925 45.635 143.155 ;
        RECT 50.120 142.935 51.030 143.155 ;
        RECT 52.565 142.925 53.915 143.155 ;
        RECT 54.425 143.155 58.325 143.835 ;
        RECT 58.660 143.155 62.125 143.835 ;
        RECT 54.425 142.925 55.355 143.155 ;
        RECT 58.660 142.925 59.580 143.155 ;
        RECT 62.245 143.025 63.615 143.835 ;
        RECT 63.635 142.965 64.065 143.750 ;
        RECT 64.320 143.155 69.135 143.835 ;
        RECT 69.145 143.155 73.045 143.835 ;
        RECT 73.785 143.155 81.095 143.835 ;
        RECT 81.105 143.155 88.415 143.835 ;
        RECT 69.145 142.925 70.075 143.155 ;
        RECT 73.785 142.925 75.135 143.155 ;
        RECT 76.670 142.935 77.580 143.155 ;
        RECT 84.620 142.935 85.530 143.155 ;
        RECT 87.065 142.925 88.415 143.155 ;
        RECT 88.465 143.025 89.835 143.835 ;
      LAYER nwell ;
        RECT 11.910 139.805 90.030 142.635 ;
      LAYER pwell ;
        RECT 12.105 138.605 13.475 139.415 ;
        RECT 13.485 138.605 16.235 139.415 ;
        RECT 16.245 138.605 19.415 139.515 ;
        RECT 19.465 139.285 20.395 139.515 ;
        RECT 19.465 138.605 23.135 139.285 ;
        RECT 23.145 138.605 24.960 139.515 ;
        RECT 24.995 138.690 25.425 139.475 ;
        RECT 29.105 139.285 30.035 139.515 ;
        RECT 32.785 139.285 33.715 139.515 ;
        RECT 26.365 138.605 30.035 139.285 ;
        RECT 30.045 138.605 33.715 139.285 ;
        RECT 33.725 138.605 35.540 139.515 ;
        RECT 35.580 138.605 37.395 139.515 ;
        RECT 37.885 138.605 39.235 139.515 ;
        RECT 42.760 139.285 43.670 139.505 ;
        RECT 45.205 139.285 46.555 139.515 ;
        RECT 39.245 138.605 46.555 139.285 ;
        RECT 46.605 139.285 47.535 139.515 ;
        RECT 46.605 138.605 50.505 139.285 ;
        RECT 50.755 138.690 51.185 139.475 ;
        RECT 54.720 139.285 55.630 139.505 ;
        RECT 57.165 139.285 58.515 139.515 ;
        RECT 62.080 139.285 62.990 139.505 ;
        RECT 64.525 139.285 65.875 139.515 ;
        RECT 51.205 138.605 58.515 139.285 ;
        RECT 58.565 138.605 65.875 139.285 ;
        RECT 65.965 139.285 67.315 139.515 ;
        RECT 68.850 139.285 69.760 139.505 ;
        RECT 75.255 139.285 76.185 139.515 ;
        RECT 65.965 138.605 73.275 139.285 ;
        RECT 74.350 138.605 76.185 139.285 ;
        RECT 76.515 138.690 76.945 139.475 ;
        RECT 77.060 139.285 77.980 139.515 ;
        RECT 80.740 139.285 81.660 139.515 ;
        RECT 77.060 138.605 80.525 139.285 ;
        RECT 80.740 138.605 84.205 139.285 ;
        RECT 84.325 138.605 87.800 139.515 ;
        RECT 88.465 138.605 89.835 139.415 ;
        RECT 12.245 138.395 12.415 138.605 ;
        RECT 13.625 138.395 13.795 138.605 ;
        RECT 19.145 138.395 19.315 138.605 ;
        RECT 21.900 138.445 22.020 138.555 ;
        RECT 22.825 138.415 22.995 138.605 ;
        RECT 24.205 138.395 24.375 138.585 ;
        RECT 24.665 138.415 24.835 138.605 ;
        RECT 25.595 138.450 25.755 138.560 ;
        RECT 26.505 138.415 26.675 138.605 ;
        RECT 27.425 138.395 27.595 138.585 ;
        RECT 30.185 138.415 30.355 138.605 ;
        RECT 30.645 138.395 30.815 138.585 ;
        RECT 31.105 138.395 31.275 138.585 ;
        RECT 32.485 138.395 32.655 138.585 ;
        RECT 34.790 138.395 34.960 138.585 ;
        RECT 35.245 138.415 35.415 138.605 ;
        RECT 35.705 138.415 35.875 138.605 ;
        RECT 37.545 138.555 37.715 138.585 ;
        RECT 36.160 138.445 36.280 138.555 ;
        RECT 37.540 138.445 37.715 138.555 ;
        RECT 37.545 138.395 37.715 138.445 ;
        RECT 38.000 138.415 38.170 138.605 ;
        RECT 38.460 138.445 38.580 138.555 ;
        RECT 38.925 138.395 39.095 138.585 ;
        RECT 39.385 138.415 39.555 138.605 ;
        RECT 42.605 138.395 42.775 138.585 ;
        RECT 47.020 138.415 47.190 138.605 ;
        RECT 47.665 138.395 47.835 138.585 ;
        RECT 51.345 138.415 51.515 138.605 ;
        RECT 55.300 138.395 55.470 138.585 ;
        RECT 58.705 138.415 58.875 138.605 ;
        RECT 59.160 138.445 59.280 138.555 ;
        RECT 59.900 138.395 60.070 138.585 ;
        RECT 64.225 138.395 64.395 138.585 ;
        RECT 72.505 138.395 72.675 138.585 ;
        RECT 72.965 138.395 73.135 138.605 ;
        RECT 74.350 138.585 74.515 138.605 ;
        RECT 73.435 138.450 73.595 138.560 ;
        RECT 74.345 138.415 74.515 138.585 ;
        RECT 78.300 138.395 78.470 138.585 ;
        RECT 80.325 138.415 80.495 138.605 ;
        RECT 82.155 138.395 82.325 138.585 ;
        RECT 84.005 138.415 84.175 138.605 ;
        RECT 84.470 138.415 84.640 138.605 ;
        RECT 87.225 138.415 87.395 138.585 ;
        RECT 87.695 138.440 87.855 138.550 ;
        RECT 88.140 138.445 88.260 138.555 ;
        RECT 87.225 138.395 87.390 138.415 ;
        RECT 89.525 138.395 89.695 138.605 ;
        RECT 12.105 137.585 13.475 138.395 ;
        RECT 13.485 137.585 18.995 138.395 ;
        RECT 19.005 137.585 21.755 138.395 ;
        RECT 22.225 137.715 24.515 138.395 ;
        RECT 24.525 137.715 27.735 138.395 ;
        RECT 22.225 137.485 23.145 137.715 ;
        RECT 24.525 137.485 25.660 137.715 ;
        RECT 27.745 137.485 30.915 138.395 ;
        RECT 30.965 137.585 32.335 138.395 ;
        RECT 32.345 137.715 34.635 138.395 ;
        RECT 33.715 137.485 34.635 137.715 ;
        RECT 34.645 137.485 35.995 138.395 ;
        RECT 36.495 137.485 37.845 138.395 ;
        RECT 37.875 137.525 38.305 138.310 ;
        RECT 38.895 137.715 42.360 138.395 ;
        RECT 42.465 137.715 47.280 138.395 ;
        RECT 47.525 137.715 54.835 138.395 ;
        RECT 41.440 137.485 42.360 137.715 ;
        RECT 51.040 137.495 51.950 137.715 ;
        RECT 53.485 137.485 54.835 137.715 ;
        RECT 54.885 137.715 58.785 138.395 ;
        RECT 59.485 137.715 63.385 138.395 ;
        RECT 54.885 137.485 55.815 137.715 ;
        RECT 59.485 137.485 60.415 137.715 ;
        RECT 63.635 137.525 64.065 138.310 ;
        RECT 64.085 137.585 65.455 138.395 ;
        RECT 65.505 137.715 72.815 138.395 ;
        RECT 72.825 137.715 77.640 138.395 ;
        RECT 77.885 137.715 81.785 138.395 ;
        RECT 65.505 137.485 66.855 137.715 ;
        RECT 68.390 137.495 69.300 137.715 ;
        RECT 77.885 137.485 78.815 137.715 ;
        RECT 82.025 137.485 85.235 138.395 ;
        RECT 85.555 137.715 87.390 138.395 ;
        RECT 85.555 137.485 86.485 137.715 ;
        RECT 88.465 137.585 89.835 138.395 ;
      LAYER nwell ;
        RECT 11.910 134.365 90.030 137.195 ;
      LAYER pwell ;
        RECT 100.450 137.140 106.550 146.930 ;
        RECT 100.450 137.110 106.560 137.140 ;
        RECT 100.650 136.710 101.810 137.110 ;
        RECT 103.770 135.030 106.560 137.110 ;
        RECT 12.105 133.165 13.475 133.975 ;
        RECT 13.485 133.165 14.855 133.945 ;
        RECT 14.865 133.165 20.375 133.975 ;
        RECT 20.385 133.165 24.055 133.975 ;
        RECT 24.995 133.250 25.425 134.035 ;
        RECT 25.445 133.165 30.955 133.975 ;
        RECT 30.965 133.165 33.715 133.975 ;
        RECT 34.420 133.165 39.235 133.845 ;
        RECT 39.735 133.165 42.455 134.075 ;
        RECT 44.765 133.875 45.720 134.075 ;
        RECT 43.390 133.165 44.755 133.845 ;
        RECT 44.765 133.195 47.045 133.875 ;
        RECT 47.160 133.845 48.080 134.075 ;
        RECT 44.765 133.165 45.720 133.195 ;
        RECT 12.245 132.955 12.415 133.165 ;
        RECT 13.625 132.955 13.795 133.165 ;
        RECT 15.005 132.975 15.175 133.165 ;
        RECT 18.225 132.955 18.395 133.145 ;
        RECT 18.685 132.955 18.855 133.145 ;
        RECT 20.525 132.975 20.695 133.165 ;
        RECT 24.205 132.955 24.375 133.145 ;
        RECT 25.585 132.975 25.755 133.165 ;
        RECT 28.345 132.955 28.515 133.145 ;
        RECT 30.645 132.975 30.815 133.145 ;
        RECT 30.645 132.955 30.795 132.975 ;
        RECT 31.105 132.955 31.275 133.165 ;
        RECT 33.860 132.955 34.030 133.145 ;
        RECT 34.325 132.975 34.495 133.145 ;
        RECT 37.540 133.005 37.660 133.115 ;
        RECT 38.470 132.955 38.640 133.145 ;
        RECT 38.925 132.975 39.095 133.165 ;
        RECT 39.380 133.005 39.500 133.115 ;
        RECT 39.855 133.000 40.015 133.110 ;
        RECT 40.765 132.955 40.935 133.145 ;
        RECT 42.145 132.975 42.315 133.165 ;
        RECT 42.600 133.005 42.720 133.115 ;
        RECT 43.065 132.975 43.235 133.145 ;
        RECT 46.750 132.975 46.920 133.195 ;
        RECT 47.160 133.165 50.625 133.845 ;
        RECT 50.755 133.250 51.185 134.035 ;
        RECT 51.665 133.845 52.595 134.075 ;
        RECT 55.900 133.845 56.820 134.075 ;
        RECT 51.665 133.165 55.565 133.845 ;
        RECT 55.900 133.165 59.365 133.845 ;
        RECT 59.485 133.165 61.315 133.975 ;
        RECT 61.325 133.845 62.670 134.075 ;
        RECT 65.820 133.845 66.740 134.075 ;
        RECT 61.325 133.165 63.155 133.845 ;
        RECT 63.275 133.165 66.740 133.845 ;
        RECT 66.845 133.845 68.190 134.075 ;
        RECT 68.780 133.845 69.700 134.075 ;
        RECT 75.020 133.845 75.940 134.075 ;
        RECT 66.845 133.165 68.675 133.845 ;
        RECT 68.780 133.165 72.245 133.845 ;
        RECT 72.475 133.165 75.940 133.845 ;
        RECT 76.515 133.250 76.945 134.035 ;
        RECT 76.965 133.165 80.175 134.075 ;
        RECT 84.620 133.845 85.530 134.065 ;
        RECT 87.065 133.845 88.415 134.075 ;
        RECT 81.105 133.165 88.415 133.845 ;
        RECT 88.465 133.165 89.835 133.975 ;
        RECT 48.400 132.955 48.570 133.145 ;
        RECT 50.425 132.975 50.595 133.165 ;
        RECT 51.340 133.005 51.460 133.115 ;
        RECT 52.080 132.975 52.250 133.165 ;
        RECT 52.265 132.955 52.435 133.145 ;
        RECT 55.025 132.955 55.195 133.145 ;
        RECT 56.405 132.955 56.575 133.145 ;
        RECT 59.165 132.975 59.335 133.165 ;
        RECT 59.625 132.975 59.795 133.165 ;
        RECT 62.845 132.975 63.015 133.165 ;
        RECT 63.305 132.975 63.475 133.165 ;
        RECT 64.225 132.955 64.395 133.145 ;
        RECT 68.365 132.975 68.535 133.165 ;
        RECT 71.860 132.955 72.030 133.145 ;
        RECT 72.045 132.975 72.215 133.165 ;
        RECT 72.505 132.975 72.675 133.165 ;
        RECT 77.095 133.145 77.265 133.165 ;
        RECT 76.180 133.005 76.300 133.115 ;
        RECT 77.095 132.975 77.275 133.145 ;
        RECT 80.335 133.010 80.495 133.120 ;
        RECT 77.105 132.955 77.275 132.975 ;
        RECT 80.780 132.955 80.950 133.145 ;
        RECT 81.245 132.955 81.415 133.165 ;
        RECT 89.525 132.955 89.695 133.165 ;
        RECT 12.105 132.145 13.475 132.955 ;
        RECT 13.485 132.145 14.855 132.955 ;
        RECT 14.865 132.275 18.535 132.955 ;
        RECT 14.865 132.045 15.795 132.275 ;
        RECT 18.545 132.145 24.055 132.955 ;
        RECT 24.065 132.275 25.895 132.955 ;
        RECT 24.550 132.045 25.895 132.275 ;
        RECT 25.905 132.045 28.655 132.955 ;
        RECT 28.865 132.135 30.795 132.955 ;
        RECT 30.965 132.145 32.795 132.955 ;
        RECT 28.865 132.045 29.815 132.135 ;
        RECT 32.825 132.045 34.175 132.955 ;
        RECT 34.590 132.275 37.015 132.955 ;
        RECT 37.875 132.085 38.305 132.870 ;
        RECT 38.325 132.045 39.675 132.955 ;
        RECT 40.625 132.275 47.935 132.955 ;
        RECT 44.140 132.055 45.050 132.275 ;
        RECT 46.585 132.045 47.935 132.275 ;
        RECT 47.985 132.275 51.885 132.955 ;
        RECT 52.125 132.275 54.865 132.955 ;
        RECT 47.985 132.045 48.915 132.275 ;
        RECT 54.885 132.145 56.255 132.955 ;
        RECT 56.265 132.275 63.575 132.955 ;
        RECT 59.780 132.055 60.690 132.275 ;
        RECT 62.225 132.045 63.575 132.275 ;
        RECT 63.635 132.085 64.065 132.870 ;
        RECT 64.085 132.275 71.395 132.955 ;
        RECT 67.600 132.055 68.510 132.275 ;
        RECT 70.045 132.045 71.395 132.275 ;
        RECT 71.445 132.275 75.345 132.955 ;
        RECT 75.585 132.275 77.415 132.955 ;
        RECT 71.445 132.045 72.375 132.275 ;
        RECT 75.585 132.045 76.930 132.275 ;
        RECT 77.620 132.045 81.095 132.955 ;
        RECT 81.105 132.275 88.415 132.955 ;
        RECT 84.620 132.055 85.530 132.275 ;
        RECT 87.065 132.045 88.415 132.275 ;
        RECT 88.465 132.145 89.835 132.955 ;
      LAYER nwell ;
        RECT 101.660 132.920 106.500 135.030 ;
        RECT 107.780 134.690 117.970 146.940 ;
      LAYER pwell ;
        RECT 120.330 137.140 126.430 146.930 ;
        RECT 120.330 137.110 126.440 137.140 ;
        RECT 120.530 136.710 121.690 137.110 ;
        RECT 123.650 135.030 126.440 137.110 ;
      LAYER nwell ;
        RECT 121.540 132.920 126.380 135.030 ;
        RECT 127.660 134.690 137.850 146.940 ;
      LAYER pwell ;
        RECT 140.360 137.140 146.460 146.930 ;
        RECT 140.360 137.110 146.470 137.140 ;
        RECT 140.560 136.710 141.720 137.110 ;
        RECT 143.680 135.030 146.470 137.110 ;
      LAYER nwell ;
        RECT 141.570 132.920 146.410 135.030 ;
        RECT 147.690 134.690 157.880 146.940 ;
        RECT 11.910 128.925 90.030 131.755 ;
      LAYER pwell ;
        RECT 12.105 127.725 13.475 128.535 ;
        RECT 17.460 128.405 18.370 128.625 ;
        RECT 19.905 128.405 21.255 128.635 ;
        RECT 13.945 127.725 21.255 128.405 ;
        RECT 21.305 127.725 22.655 128.635 ;
        RECT 23.140 127.955 24.975 128.635 ;
        RECT 23.140 127.725 24.830 127.955 ;
        RECT 24.995 127.810 25.425 128.595 ;
        RECT 25.465 127.725 26.815 128.635 ;
        RECT 32.325 128.405 33.255 128.635 ;
        RECT 36.005 128.405 36.935 128.635 ;
        RECT 39.020 128.405 40.155 128.635 ;
        RECT 26.825 127.725 29.565 128.405 ;
        RECT 29.585 127.725 33.255 128.405 ;
        RECT 33.265 127.725 36.935 128.405 ;
        RECT 36.945 127.725 40.155 128.405 ;
        RECT 40.265 127.725 43.375 128.635 ;
        RECT 43.425 128.405 44.775 128.635 ;
        RECT 46.310 128.405 47.220 128.625 ;
        RECT 43.425 127.725 50.735 128.405 ;
        RECT 50.755 127.810 51.185 128.595 ;
        RECT 51.205 127.725 53.955 128.535 ;
        RECT 54.435 127.725 55.785 128.635 ;
        RECT 55.825 127.725 57.175 128.635 ;
        RECT 57.185 128.405 58.115 128.635 ;
        RECT 61.325 128.405 62.670 128.635 ;
        RECT 57.185 127.725 61.085 128.405 ;
        RECT 61.325 127.725 63.155 128.405 ;
        RECT 63.165 127.725 64.515 128.635 ;
        RECT 64.545 127.725 65.895 128.635 ;
        RECT 66.425 128.405 67.775 128.635 ;
        RECT 69.310 128.405 70.220 128.625 ;
        RECT 75.255 128.405 76.185 128.635 ;
        RECT 66.425 127.725 73.735 128.405 ;
        RECT 74.350 127.725 76.185 128.405 ;
        RECT 76.515 127.810 76.945 128.595 ;
        RECT 76.965 127.725 80.440 128.635 ;
        RECT 80.840 127.725 84.315 128.635 ;
        RECT 84.325 127.725 87.535 128.635 ;
        RECT 88.465 127.725 89.835 128.535 ;
        RECT 12.245 127.515 12.415 127.725 ;
        RECT 13.625 127.675 13.795 127.705 ;
        RECT 13.620 127.565 13.795 127.675 ;
        RECT 13.625 127.515 13.795 127.565 ;
        RECT 14.085 127.535 14.255 127.725 ;
        RECT 20.990 127.515 21.160 127.705 ;
        RECT 21.450 127.535 21.620 127.725 ;
        RECT 24.660 127.535 24.830 127.725 ;
        RECT 25.580 127.515 25.750 127.725 ;
        RECT 26.040 127.565 26.160 127.675 ;
        RECT 26.505 127.515 26.675 127.705 ;
        RECT 26.965 127.535 27.135 127.725 ;
        RECT 29.725 127.535 29.895 127.725 ;
        RECT 30.645 127.515 30.815 127.705 ;
        RECT 33.405 127.535 33.575 127.725 ;
        RECT 37.085 127.535 37.255 127.725 ;
        RECT 38.465 127.515 38.635 127.705 ;
        RECT 40.305 127.535 40.475 127.725 ;
        RECT 43.985 127.515 44.155 127.705 ;
        RECT 49.505 127.515 49.675 127.705 ;
        RECT 50.425 127.535 50.595 127.725 ;
        RECT 51.345 127.535 51.515 127.725 ;
        RECT 52.260 127.565 52.380 127.675 ;
        RECT 52.725 127.515 52.895 127.705 ;
        RECT 54.100 127.565 54.220 127.675 ;
        RECT 55.485 127.535 55.655 127.725 ;
        RECT 55.940 127.535 56.110 127.725 ;
        RECT 57.600 127.535 57.770 127.725 ;
        RECT 60.085 127.515 60.255 127.705 ;
        RECT 62.845 127.535 63.015 127.725 ;
        RECT 64.230 127.535 64.400 127.725 ;
        RECT 65.610 127.535 65.780 127.725 ;
        RECT 66.060 127.565 66.180 127.675 ;
        RECT 66.985 127.515 67.155 127.705 ;
        RECT 68.825 127.515 68.995 127.705 ;
        RECT 69.285 127.515 69.455 127.705 ;
        RECT 72.505 127.515 72.675 127.705 ;
        RECT 73.425 127.535 73.595 127.725 ;
        RECT 74.350 127.705 74.515 127.725 ;
        RECT 73.880 127.565 74.000 127.675 ;
        RECT 74.345 127.535 74.515 127.705 ;
        RECT 77.110 127.535 77.280 127.725 ;
        RECT 79.865 127.535 80.035 127.705 ;
        RECT 79.870 127.515 80.035 127.535 ;
        RECT 82.165 127.515 82.335 127.705 ;
        RECT 84.000 127.535 84.170 127.725 ;
        RECT 87.225 127.535 87.395 127.725 ;
        RECT 87.695 127.560 87.855 127.680 ;
        RECT 87.225 127.515 87.390 127.535 ;
        RECT 89.525 127.515 89.695 127.725 ;
        RECT 12.105 126.705 13.475 127.515 ;
        RECT 13.485 126.835 20.795 127.515 ;
        RECT 17.000 126.615 17.910 126.835 ;
        RECT 19.445 126.605 20.795 126.835 ;
        RECT 20.845 126.605 22.195 127.515 ;
        RECT 22.420 126.605 25.895 127.515 ;
        RECT 26.365 126.605 29.575 127.515 ;
        RECT 30.505 126.835 37.815 127.515 ;
        RECT 34.020 126.615 34.930 126.835 ;
        RECT 36.465 126.605 37.815 126.835 ;
        RECT 37.875 126.645 38.305 127.430 ;
        RECT 38.325 126.705 43.835 127.515 ;
        RECT 43.845 126.705 49.355 127.515 ;
        RECT 49.365 126.705 52.115 127.515 ;
        RECT 52.585 126.835 59.895 127.515 ;
        RECT 60.055 126.835 63.520 127.515 ;
        RECT 56.100 126.615 57.010 126.835 ;
        RECT 58.545 126.605 59.895 126.835 ;
        RECT 62.600 126.605 63.520 126.835 ;
        RECT 63.635 126.645 64.065 127.430 ;
        RECT 64.085 126.605 67.295 127.515 ;
        RECT 67.305 126.835 69.135 127.515 ;
        RECT 67.305 126.605 68.650 126.835 ;
        RECT 69.145 126.605 72.355 127.515 ;
        RECT 72.365 126.835 79.675 127.515 ;
        RECT 79.870 126.835 81.705 127.515 ;
        RECT 75.880 126.615 76.790 126.835 ;
        RECT 78.325 126.605 79.675 126.835 ;
        RECT 80.775 126.605 81.705 126.835 ;
        RECT 82.025 126.605 85.235 127.515 ;
        RECT 85.555 126.835 87.390 127.515 ;
        RECT 85.555 126.605 86.485 126.835 ;
        RECT 88.465 126.705 89.835 127.515 ;
      LAYER nwell ;
        RECT 11.910 123.485 90.030 126.315 ;
      LAYER pwell ;
        RECT 12.105 122.285 13.475 123.095 ;
        RECT 14.405 122.965 15.335 123.195 ;
        RECT 14.405 122.285 18.075 122.965 ;
        RECT 18.085 122.285 19.435 123.195 ;
        RECT 19.465 122.965 20.600 123.195 ;
        RECT 24.020 122.995 24.975 123.195 ;
        RECT 19.465 122.285 22.675 122.965 ;
        RECT 22.695 122.315 24.975 122.995 ;
        RECT 24.995 122.370 25.425 123.155 ;
        RECT 12.245 122.075 12.415 122.285 ;
        RECT 13.625 122.075 13.795 122.265 ;
        RECT 17.765 122.075 17.935 122.285 ;
        RECT 18.230 122.265 18.400 122.285 ;
        RECT 18.225 122.095 18.400 122.265 ;
        RECT 20.520 122.125 20.640 122.235 ;
        RECT 18.225 122.075 18.395 122.095 ;
        RECT 20.985 122.075 21.155 122.265 ;
        RECT 22.365 122.095 22.535 122.285 ;
        RECT 22.820 122.095 22.990 122.315 ;
        RECT 24.020 122.285 24.975 122.315 ;
        RECT 25.640 122.285 29.115 123.195 ;
        RECT 30.175 122.965 31.105 123.195 ;
        RECT 29.270 122.285 31.105 122.965 ;
        RECT 31.925 122.965 33.275 123.195 ;
        RECT 34.810 122.965 35.720 123.185 ;
        RECT 39.285 122.965 40.635 123.195 ;
        RECT 42.170 122.965 43.080 123.185 ;
        RECT 31.925 122.285 39.235 122.965 ;
        RECT 39.285 122.285 46.595 122.965 ;
        RECT 46.605 122.285 47.955 123.195 ;
        RECT 47.985 122.285 50.735 123.095 ;
        RECT 50.755 122.370 51.185 123.155 ;
        RECT 52.125 122.965 53.055 123.195 ;
        RECT 58.920 122.965 59.840 123.195 ;
        RECT 52.125 122.285 56.025 122.965 ;
        RECT 56.375 122.285 59.840 122.965 ;
        RECT 59.945 122.285 63.155 123.195 ;
        RECT 63.165 122.285 64.995 123.195 ;
        RECT 65.005 122.285 66.835 123.195 ;
        RECT 66.845 122.285 70.055 123.195 ;
        RECT 72.720 122.965 73.640 123.195 ;
        RECT 70.175 122.285 73.640 122.965 ;
        RECT 73.745 122.285 75.835 123.095 ;
        RECT 76.515 122.370 76.945 123.155 ;
        RECT 77.160 122.285 80.635 123.195 ;
        RECT 84.160 122.965 85.070 123.185 ;
        RECT 86.605 122.965 87.955 123.195 ;
        RECT 80.645 122.285 87.955 122.965 ;
        RECT 88.465 122.285 89.835 123.095 ;
        RECT 24.205 122.075 24.375 122.265 ;
        RECT 12.105 121.265 13.475 122.075 ;
        RECT 13.485 121.265 16.235 122.075 ;
        RECT 16.245 121.165 18.060 122.075 ;
        RECT 18.085 121.395 20.375 122.075 ;
        RECT 19.455 121.165 20.375 121.395 ;
        RECT 20.945 121.165 24.055 122.075 ;
        RECT 24.065 121.265 25.895 122.075 ;
        RECT 26.045 122.045 26.215 122.265 ;
        RECT 28.800 122.095 28.970 122.285 ;
        RECT 29.270 122.265 29.435 122.285 ;
        RECT 29.260 122.095 29.435 122.265 ;
        RECT 31.565 122.235 31.735 122.265 ;
        RECT 31.560 122.125 31.735 122.235 ;
        RECT 28.170 122.045 29.115 122.075 ;
        RECT 29.260 122.045 29.430 122.095 ;
        RECT 31.565 122.075 31.735 122.125 ;
        RECT 34.790 122.075 34.960 122.265 ;
        RECT 38.925 122.095 39.095 122.285 ;
        RECT 39.845 122.075 40.015 122.265 ;
        RECT 40.315 122.120 40.475 122.230 ;
        RECT 41.225 122.075 41.395 122.265 ;
        RECT 46.285 122.095 46.455 122.285 ;
        RECT 46.750 122.095 46.920 122.285 ;
        RECT 48.125 122.095 48.295 122.285 ;
        RECT 48.585 122.075 48.755 122.265 ;
        RECT 51.355 122.130 51.515 122.240 ;
        RECT 52.540 122.095 52.710 122.285 ;
        RECT 56.405 122.095 56.575 122.285 ;
        RECT 59.165 122.075 59.335 122.265 ;
        RECT 59.625 122.075 59.795 122.265 ;
        RECT 60.085 122.095 60.255 122.285 ;
        RECT 62.855 122.120 63.015 122.230 ;
        RECT 63.310 122.095 63.480 122.285 ;
        RECT 64.225 122.075 64.395 122.265 ;
        RECT 66.520 122.095 66.690 122.285 ;
        RECT 69.745 122.095 69.915 122.285 ;
        RECT 70.205 122.095 70.375 122.285 ;
        RECT 73.885 122.095 74.055 122.285 ;
        RECT 74.345 122.075 74.515 122.265 ;
        RECT 75.730 122.075 75.900 122.265 ;
        RECT 76.185 122.075 76.355 122.265 ;
        RECT 80.320 122.095 80.490 122.285 ;
        RECT 80.785 122.095 80.955 122.285 ;
        RECT 85.385 122.095 85.555 122.265 ;
        RECT 85.845 122.095 86.015 122.265 ;
        RECT 88.140 122.125 88.260 122.235 ;
        RECT 85.385 122.075 85.550 122.095 ;
        RECT 30.460 122.045 31.415 122.075 ;
        RECT 26.045 121.845 29.115 122.045 ;
        RECT 25.905 121.365 29.115 121.845 ;
        RECT 29.135 121.365 31.415 122.045 ;
        RECT 25.905 121.165 26.835 121.365 ;
        RECT 28.170 121.165 29.115 121.365 ;
        RECT 30.460 121.165 31.415 121.365 ;
        RECT 31.465 121.165 34.635 122.075 ;
        RECT 34.645 121.165 37.565 122.075 ;
        RECT 37.875 121.205 38.305 121.990 ;
        RECT 38.325 121.395 40.155 122.075 ;
        RECT 41.085 121.395 48.395 122.075 ;
        RECT 48.445 121.395 55.755 122.075 ;
        RECT 44.600 121.175 45.510 121.395 ;
        RECT 47.045 121.165 48.395 121.395 ;
        RECT 51.960 121.175 52.870 121.395 ;
        RECT 54.405 121.165 55.755 121.395 ;
        RECT 55.900 121.395 59.365 122.075 ;
        RECT 55.900 121.165 56.820 121.395 ;
        RECT 59.485 121.165 62.695 122.075 ;
        RECT 63.635 121.205 64.065 121.990 ;
        RECT 64.135 121.165 67.295 122.075 ;
        RECT 67.345 121.395 74.655 122.075 ;
        RECT 67.345 121.165 68.695 121.395 ;
        RECT 70.230 121.175 71.140 121.395 ;
        RECT 74.665 121.165 76.015 122.075 ;
        RECT 76.045 121.395 83.355 122.075 ;
        RECT 79.560 121.175 80.470 121.395 ;
        RECT 82.005 121.165 83.355 121.395 ;
        RECT 83.715 121.395 85.550 122.075 ;
        RECT 85.850 122.075 86.015 122.095 ;
        RECT 89.525 122.075 89.695 122.285 ;
        RECT 100.450 122.140 106.550 131.930 ;
        RECT 100.450 122.110 106.560 122.140 ;
        RECT 85.850 121.395 87.685 122.075 ;
        RECT 83.715 121.165 84.645 121.395 ;
        RECT 86.755 121.165 87.685 121.395 ;
        RECT 88.465 121.265 89.835 122.075 ;
        RECT 100.650 121.710 101.810 122.110 ;
      LAYER nwell ;
        RECT 11.910 118.045 90.030 120.875 ;
      LAYER pwell ;
        RECT 103.770 120.030 106.560 122.110 ;
      LAYER nwell ;
        RECT 101.660 117.920 106.500 120.030 ;
        RECT 107.780 119.690 117.970 131.940 ;
      LAYER pwell ;
        RECT 120.330 122.200 126.430 131.990 ;
        RECT 120.330 122.170 126.440 122.200 ;
        RECT 120.530 121.770 121.690 122.170 ;
        RECT 123.650 120.090 126.440 122.170 ;
      LAYER nwell ;
        RECT 121.540 117.980 126.380 120.090 ;
        RECT 127.660 119.750 137.850 132.000 ;
      LAYER pwell ;
        RECT 140.360 122.200 146.460 131.990 ;
        RECT 140.360 122.170 146.470 122.200 ;
        RECT 140.560 121.770 141.720 122.170 ;
        RECT 143.680 120.090 146.470 122.170 ;
      LAYER nwell ;
        RECT 141.570 117.980 146.410 120.090 ;
        RECT 147.690 119.750 157.880 132.000 ;
      LAYER pwell ;
        RECT 12.105 116.845 13.475 117.655 ;
        RECT 13.485 116.845 18.995 117.655 ;
        RECT 19.005 116.845 21.755 117.655 ;
        RECT 21.865 116.845 24.975 117.755 ;
        RECT 24.995 116.930 25.425 117.715 ;
        RECT 26.365 116.845 30.020 117.755 ;
        RECT 30.670 116.845 34.540 117.755 ;
        RECT 34.645 116.845 39.460 117.525 ;
        RECT 39.725 116.845 41.075 117.755 ;
        RECT 44.600 117.525 45.510 117.745 ;
        RECT 47.045 117.525 48.395 117.755 ;
        RECT 41.085 116.845 48.395 117.525 ;
        RECT 48.445 116.845 50.275 117.655 ;
        RECT 50.755 116.930 51.185 117.715 ;
        RECT 51.205 117.525 52.135 117.755 ;
        RECT 51.205 116.845 55.105 117.525 ;
        RECT 55.345 116.845 58.555 117.755 ;
        RECT 60.165 117.665 61.115 117.755 ;
        RECT 59.185 116.845 61.115 117.665 ;
        RECT 61.325 116.845 66.140 117.525 ;
        RECT 66.385 116.845 69.305 117.755 ;
        RECT 73.725 117.525 74.655 117.755 ;
        RECT 70.755 116.845 74.655 117.525 ;
        RECT 74.665 117.525 76.010 117.755 ;
        RECT 74.665 116.845 76.495 117.525 ;
        RECT 76.515 116.930 76.945 117.715 ;
        RECT 82.025 117.525 83.370 117.755 ;
        RECT 85.270 117.525 86.615 117.755 ;
        RECT 87.110 117.525 88.455 117.755 ;
        RECT 76.965 116.845 81.780 117.525 ;
        RECT 82.025 116.845 83.855 117.525 ;
        RECT 84.785 116.845 86.615 117.525 ;
        RECT 86.625 116.845 88.455 117.525 ;
        RECT 88.465 116.845 89.835 117.655 ;
        RECT 12.245 116.635 12.415 116.845 ;
        RECT 13.625 116.825 13.795 116.845 ;
        RECT 13.625 116.655 13.805 116.825 ;
        RECT 13.635 116.635 13.805 116.655 ;
        RECT 15.005 116.635 15.175 116.825 ;
        RECT 19.145 116.655 19.315 116.845 ;
        RECT 21.905 116.825 22.075 116.845 ;
        RECT 20.520 116.685 20.640 116.795 ;
        RECT 21.900 116.655 22.075 116.825 ;
        RECT 22.360 116.685 22.480 116.795 ;
        RECT 21.900 116.635 22.070 116.655 ;
        RECT 22.825 116.635 22.995 116.825 ;
        RECT 25.595 116.690 25.755 116.800 ;
        RECT 26.035 116.635 26.205 116.825 ;
        RECT 26.510 116.655 26.680 116.845 ;
        RECT 30.670 116.825 30.815 116.845 ;
        RECT 30.180 116.685 30.300 116.795 ;
        RECT 30.645 116.655 30.815 116.825 ;
        RECT 31.105 116.655 31.275 116.825 ;
        RECT 31.105 116.635 31.270 116.655 ;
        RECT 31.565 116.635 31.735 116.825 ;
        RECT 34.785 116.655 34.955 116.845 ;
        RECT 39.840 116.825 40.010 116.845 ;
        RECT 35.245 116.635 35.415 116.825 ;
        RECT 39.840 116.655 40.015 116.825 ;
        RECT 40.315 116.680 40.475 116.790 ;
        RECT 39.845 116.635 40.015 116.655 ;
        RECT 41.225 116.635 41.395 116.845 ;
        RECT 44.910 116.635 45.080 116.825 ;
        RECT 46.285 116.635 46.455 116.825 ;
        RECT 47.665 116.635 47.835 116.825 ;
        RECT 48.585 116.655 48.755 116.845 ;
        RECT 50.420 116.685 50.540 116.795 ;
        RECT 51.620 116.655 51.790 116.845 ;
        RECT 52.725 116.635 52.895 116.825 ;
        RECT 54.105 116.635 54.275 116.825 ;
        RECT 58.255 116.655 58.425 116.845 ;
        RECT 59.185 116.825 59.335 116.845 ;
        RECT 61.465 116.825 61.635 116.845 ;
        RECT 58.700 116.685 58.820 116.795 ;
        RECT 59.165 116.655 59.335 116.825 ;
        RECT 61.460 116.655 61.635 116.825 ;
        RECT 64.225 116.655 64.395 116.825 ;
        RECT 66.530 116.655 66.700 116.845 ;
        RECT 12.105 115.825 13.475 116.635 ;
        RECT 13.485 115.855 14.855 116.635 ;
        RECT 14.865 115.825 20.375 116.635 ;
        RECT 20.865 115.725 22.215 116.635 ;
        RECT 22.685 115.725 25.895 116.635 ;
        RECT 25.905 115.725 29.115 116.635 ;
        RECT 29.435 115.955 31.270 116.635 ;
        RECT 31.425 115.955 35.095 116.635 ;
        RECT 29.435 115.725 30.365 115.955 ;
        RECT 34.165 115.725 35.095 115.955 ;
        RECT 35.115 115.725 37.845 116.635 ;
        RECT 37.875 115.765 38.305 116.550 ;
        RECT 38.325 115.955 40.155 116.635 ;
        RECT 41.195 115.955 44.660 116.635 ;
        RECT 43.740 115.725 44.660 115.955 ;
        RECT 44.765 115.725 46.115 116.635 ;
        RECT 46.145 115.825 47.515 116.635 ;
        RECT 47.525 115.955 52.340 116.635 ;
        RECT 52.585 115.825 53.955 116.635 ;
        RECT 53.965 115.955 61.275 116.635 ;
        RECT 61.460 116.605 61.630 116.655 ;
        RECT 64.235 116.635 64.395 116.655 ;
        RECT 68.365 116.635 68.535 116.825 ;
        RECT 69.755 116.690 69.915 116.800 ;
        RECT 74.070 116.655 74.240 116.845 ;
        RECT 76.185 116.655 76.355 116.845 ;
        RECT 77.105 116.655 77.275 116.845 ;
        RECT 78.945 116.635 79.115 116.825 ;
        RECT 79.410 116.635 79.580 116.825 ;
        RECT 83.085 116.635 83.255 116.825 ;
        RECT 83.545 116.655 83.715 116.845 ;
        RECT 84.015 116.690 84.175 116.800 ;
        RECT 84.925 116.655 85.095 116.845 ;
        RECT 86.305 116.655 86.475 116.825 ;
        RECT 86.305 116.635 86.470 116.655 ;
        RECT 86.765 116.635 86.935 116.845 ;
        RECT 89.525 116.635 89.695 116.845 ;
        RECT 62.660 116.605 63.615 116.635 ;
        RECT 57.480 115.735 58.390 115.955 ;
        RECT 59.925 115.725 61.275 115.955 ;
        RECT 61.335 115.925 63.615 116.605 ;
        RECT 62.660 115.725 63.615 115.925 ;
        RECT 63.635 115.765 64.065 116.550 ;
        RECT 64.235 115.725 67.890 116.635 ;
        RECT 68.225 115.955 75.535 116.635 ;
        RECT 71.740 115.735 72.650 115.955 ;
        RECT 74.185 115.725 75.535 115.955 ;
        RECT 75.680 115.955 79.145 116.635 ;
        RECT 75.680 115.725 76.600 115.955 ;
        RECT 79.265 115.725 82.740 116.635 ;
        RECT 82.945 115.855 84.315 116.635 ;
        RECT 84.635 115.955 86.470 116.635 ;
        RECT 86.625 115.955 88.455 116.635 ;
        RECT 84.635 115.725 85.565 115.955 ;
        RECT 87.110 115.725 88.455 115.955 ;
        RECT 88.465 115.825 89.835 116.635 ;
      LAYER nwell ;
        RECT 11.910 112.605 90.030 115.435 ;
      LAYER pwell ;
        RECT 12.105 111.405 13.475 112.215 ;
        RECT 13.955 112.085 16.955 112.315 ;
        RECT 18.545 112.085 19.475 112.315 ;
        RECT 13.955 111.995 18.535 112.085 ;
        RECT 13.945 111.635 18.535 111.995 ;
        RECT 13.945 111.445 14.875 111.635 ;
        RECT 13.955 111.405 14.875 111.445 ;
        RECT 16.965 111.405 18.535 111.635 ;
        RECT 18.545 111.405 22.215 112.085 ;
        RECT 22.225 111.635 24.060 112.315 ;
        RECT 22.370 111.405 24.060 111.635 ;
        RECT 24.995 111.490 25.425 112.275 ;
        RECT 25.445 112.085 26.370 112.315 ;
        RECT 29.785 112.085 33.715 112.315 ;
        RECT 36.925 112.085 37.855 112.315 ;
        RECT 25.445 111.405 29.115 112.085 ;
        RECT 29.300 111.405 33.715 112.085 ;
        RECT 34.185 111.405 37.855 112.085 ;
        RECT 37.865 111.405 40.975 112.315 ;
        RECT 44.600 112.085 45.510 112.305 ;
        RECT 47.045 112.085 48.395 112.315 ;
        RECT 41.085 111.405 48.395 112.085 ;
        RECT 48.445 111.405 50.275 112.215 ;
        RECT 50.755 111.490 51.185 112.275 ;
        RECT 51.255 111.405 54.415 112.315 ;
        RECT 55.425 111.405 58.425 112.315 ;
        RECT 58.565 111.405 59.915 112.315 ;
        RECT 59.945 111.405 61.295 112.315 ;
        RECT 63.980 112.085 64.900 112.315 ;
        RECT 61.435 111.405 64.900 112.085 ;
        RECT 65.200 111.405 68.675 112.315 ;
        RECT 68.705 111.405 70.055 112.315 ;
        RECT 70.065 112.085 70.995 112.315 ;
        RECT 70.065 111.405 73.965 112.085 ;
        RECT 74.205 111.405 76.035 112.215 ;
        RECT 76.515 111.490 76.945 112.275 ;
        RECT 77.735 112.085 78.665 112.315 ;
        RECT 77.735 111.405 79.570 112.085 ;
        RECT 79.725 111.405 81.095 112.215 ;
        RECT 84.620 112.085 85.530 112.305 ;
        RECT 87.065 112.085 88.415 112.315 ;
        RECT 81.105 111.405 88.415 112.085 ;
        RECT 88.465 111.405 89.835 112.215 ;
        RECT 12.245 111.195 12.415 111.405 ;
        RECT 13.620 111.245 13.740 111.355 ;
        RECT 14.085 111.195 14.255 111.385 ;
        RECT 18.225 111.215 18.395 111.405 ;
        RECT 21.905 111.215 22.075 111.405 ;
        RECT 22.370 111.215 22.540 111.405 ;
        RECT 24.205 111.195 24.375 111.385 ;
        RECT 24.660 111.350 24.780 111.355 ;
        RECT 24.660 111.245 24.835 111.350 ;
        RECT 24.675 111.240 24.835 111.245 ;
        RECT 12.105 110.385 13.475 111.195 ;
        RECT 13.945 110.515 21.255 111.195 ;
        RECT 17.460 110.295 18.370 110.515 ;
        RECT 19.905 110.285 21.255 110.515 ;
        RECT 21.305 110.285 24.475 111.195 ;
        RECT 25.590 111.165 25.760 111.405 ;
        RECT 29.300 111.385 29.410 111.405 ;
        RECT 29.240 111.350 29.410 111.385 ;
        RECT 29.240 111.240 29.435 111.350 ;
        RECT 33.860 111.245 33.980 111.355 ;
        RECT 29.240 111.215 29.410 111.240 ;
        RECT 34.325 111.215 34.495 111.405 ;
        RECT 37.540 111.195 37.710 111.385 ;
        RECT 40.765 111.215 40.935 111.405 ;
        RECT 41.225 111.215 41.395 111.405 ;
        RECT 45.365 111.195 45.535 111.385 ;
        RECT 45.825 111.195 45.995 111.385 ;
        RECT 48.585 111.215 48.755 111.405 ;
        RECT 50.425 111.355 50.595 111.385 ;
        RECT 50.420 111.245 50.595 111.355 ;
        RECT 50.425 111.195 50.595 111.245 ;
        RECT 51.345 111.215 51.515 111.405 ;
        RECT 54.105 111.195 54.275 111.385 ;
        RECT 54.565 111.195 54.735 111.385 ;
        RECT 55.485 111.215 55.655 111.405 ;
        RECT 58.245 111.195 58.415 111.385 ;
        RECT 58.710 111.215 58.880 111.405 ;
        RECT 59.630 111.195 59.800 111.385 ;
        RECT 61.010 111.215 61.180 111.405 ;
        RECT 61.465 111.215 61.635 111.405 ;
        RECT 62.855 111.240 63.015 111.350 ;
        RECT 64.225 111.195 64.395 111.385 ;
        RECT 65.605 111.195 65.775 111.385 ;
        RECT 68.360 111.215 68.530 111.405 ;
        RECT 68.820 111.215 68.990 111.405 ;
        RECT 69.295 111.240 69.455 111.350 ;
        RECT 70.480 111.215 70.650 111.405 ;
        RECT 73.420 111.195 73.590 111.385 ;
        RECT 73.885 111.195 74.055 111.385 ;
        RECT 74.345 111.215 74.515 111.405 ;
        RECT 79.405 111.385 79.570 111.405 ;
        RECT 76.180 111.245 76.300 111.355 ;
        RECT 77.100 111.245 77.220 111.355 ;
        RECT 79.405 111.215 79.575 111.385 ;
        RECT 79.865 111.215 80.035 111.405 ;
        RECT 81.245 111.385 81.415 111.405 ;
        RECT 81.245 111.215 81.420 111.385 ;
        RECT 81.250 111.195 81.420 111.215 ;
        RECT 84.915 111.195 85.085 111.385 ;
        RECT 88.140 111.245 88.260 111.355 ;
        RECT 89.525 111.195 89.695 111.405 ;
        RECT 28.165 111.165 29.115 111.195 ;
        RECT 25.445 110.485 29.115 111.165 ;
        RECT 28.165 110.285 29.115 110.485 ;
        RECT 30.295 110.285 37.855 111.195 ;
        RECT 37.875 110.325 38.305 111.110 ;
        RECT 38.365 110.515 45.675 111.195 ;
        RECT 38.365 110.285 39.715 110.515 ;
        RECT 41.250 110.295 42.160 110.515 ;
        RECT 45.685 110.385 47.055 111.195 ;
        RECT 47.160 110.515 50.625 111.195 ;
        RECT 50.840 110.515 54.305 111.195 ;
        RECT 47.160 110.285 48.080 110.515 ;
        RECT 50.840 110.285 51.760 110.515 ;
        RECT 54.425 110.385 58.095 111.195 ;
        RECT 58.105 110.385 59.475 111.195 ;
        RECT 59.485 110.285 62.405 111.195 ;
        RECT 63.635 110.325 64.065 111.110 ;
        RECT 64.095 110.285 65.445 111.195 ;
        RECT 65.465 110.385 69.135 111.195 ;
        RECT 70.260 110.285 73.735 111.195 ;
        RECT 73.745 110.515 81.055 111.195 ;
        RECT 77.260 110.295 78.170 110.515 ;
        RECT 79.705 110.285 81.055 110.515 ;
        RECT 81.105 110.285 84.580 111.195 ;
        RECT 84.785 110.285 87.995 111.195 ;
        RECT 88.465 110.385 89.835 111.195 ;
      LAYER nwell ;
        RECT 11.910 107.165 90.030 109.995 ;
      LAYER pwell ;
        RECT 100.400 107.200 106.500 116.990 ;
        RECT 100.400 107.170 106.510 107.200 ;
        RECT 12.105 105.965 13.475 106.775 ;
        RECT 17.000 106.645 17.910 106.865 ;
        RECT 19.445 106.645 20.795 106.875 ;
        RECT 13.485 105.965 20.795 106.645 ;
        RECT 20.845 105.965 22.215 106.775 ;
        RECT 22.225 105.965 24.975 106.875 ;
        RECT 24.995 106.050 25.425 106.835 ;
        RECT 25.445 105.965 27.275 106.775 ;
        RECT 27.285 106.675 28.230 106.875 ;
        RECT 27.285 105.995 30.035 106.675 ;
        RECT 27.285 105.965 28.230 105.995 ;
        RECT 12.245 105.755 12.415 105.965 ;
        RECT 13.625 105.755 13.795 105.965 ;
        RECT 15.465 105.755 15.635 105.945 ;
        RECT 18.685 105.755 18.855 105.945 ;
        RECT 20.985 105.775 21.155 105.965 ;
        RECT 21.440 105.805 21.560 105.915 ;
        RECT 23.740 105.755 23.910 105.945 ;
        RECT 24.200 105.805 24.320 105.915 ;
        RECT 24.665 105.755 24.835 105.965 ;
        RECT 25.585 105.775 25.755 105.965 ;
        RECT 27.425 105.755 27.595 105.945 ;
        RECT 28.805 105.755 28.975 105.945 ;
        RECT 29.720 105.775 29.890 105.995 ;
        RECT 30.145 105.965 33.255 106.875 ;
        RECT 36.780 106.645 37.690 106.865 ;
        RECT 39.225 106.645 40.575 106.875 ;
        RECT 33.265 105.965 40.575 106.645 ;
        RECT 40.625 105.965 44.295 106.775 ;
        RECT 44.500 105.965 47.975 106.875 ;
        RECT 47.985 105.965 50.275 106.875 ;
        RECT 50.755 106.050 51.185 106.835 ;
        RECT 51.205 105.965 53.035 106.875 ;
        RECT 53.965 105.965 57.175 106.875 ;
        RECT 57.185 105.965 60.855 106.775 ;
        RECT 64.535 106.645 65.455 106.875 ;
        RECT 61.870 105.965 65.455 106.645 ;
        RECT 65.475 106.645 67.435 106.875 ;
        RECT 65.475 105.965 67.925 106.645 ;
        RECT 68.225 105.965 73.735 106.775 ;
        RECT 74.665 106.645 76.010 106.875 ;
        RECT 74.665 105.965 76.495 106.645 ;
        RECT 76.515 106.050 76.945 106.835 ;
        RECT 80.480 106.645 81.390 106.865 ;
        RECT 82.925 106.645 84.275 106.875 ;
        RECT 76.965 105.965 84.275 106.645 ;
        RECT 84.785 105.965 87.995 106.875 ;
        RECT 88.465 105.965 89.835 106.775 ;
        RECT 100.600 106.770 101.760 107.170 ;
        RECT 30.185 105.775 30.355 105.965 ;
        RECT 33.405 105.755 33.575 105.965 ;
        RECT 12.105 104.945 13.475 105.755 ;
        RECT 13.485 104.945 15.315 105.755 ;
        RECT 15.365 104.845 18.535 105.755 ;
        RECT 18.545 105.075 21.285 105.755 ;
        RECT 22.220 105.525 23.910 105.755 ;
        RECT 22.220 104.845 24.055 105.525 ;
        RECT 24.525 105.075 27.275 105.755 ;
        RECT 26.345 104.845 27.275 105.075 ;
        RECT 27.295 104.845 28.645 105.755 ;
        RECT 28.665 104.945 30.495 105.755 ;
        RECT 30.635 104.845 33.635 105.755 ;
        RECT 33.725 105.725 34.670 105.755 ;
        RECT 36.160 105.725 36.330 105.945 ;
        RECT 36.625 105.755 36.795 105.945 ;
        RECT 38.465 105.755 38.635 105.945 ;
        RECT 40.765 105.775 40.935 105.965 ;
        RECT 41.225 105.755 41.395 105.945 ;
        RECT 47.660 105.775 47.830 105.965 ;
        RECT 48.125 105.775 48.295 105.965 ;
        RECT 33.725 105.045 36.475 105.725 ;
        RECT 33.725 104.845 34.670 105.045 ;
        RECT 36.485 104.945 37.855 105.755 ;
        RECT 37.875 104.885 38.305 105.670 ;
        RECT 38.325 104.945 41.075 105.755 ;
        RECT 41.085 105.075 48.395 105.755 ;
        RECT 48.590 105.725 48.760 105.945 ;
        RECT 50.420 105.805 50.540 105.915 ;
        RECT 51.350 105.775 51.520 105.965 ;
        RECT 51.805 105.755 51.975 105.945 ;
        RECT 53.195 105.810 53.355 105.920 ;
        RECT 54.095 105.775 54.265 105.965 ;
        RECT 57.325 105.775 57.495 105.965 ;
        RECT 65.140 105.945 65.310 105.965 ;
        RECT 67.905 105.945 67.925 105.965 ;
        RECT 59.160 105.805 59.280 105.915 ;
        RECT 60.540 105.755 60.710 105.945 ;
        RECT 61.005 105.755 61.175 105.945 ;
        RECT 65.140 105.775 65.320 105.945 ;
        RECT 65.600 105.805 65.720 105.915 ;
        RECT 65.150 105.755 65.320 105.775 ;
        RECT 66.065 105.755 66.235 105.945 ;
        RECT 67.905 105.775 68.075 105.945 ;
        RECT 68.365 105.775 68.535 105.965 ;
        RECT 69.560 105.755 69.730 105.945 ;
        RECT 73.895 105.810 74.055 105.920 ;
        RECT 76.185 105.775 76.355 105.965 ;
        RECT 77.105 105.945 77.275 105.965 ;
        RECT 76.645 105.755 76.815 105.945 ;
        RECT 77.105 105.775 77.280 105.945 ;
        RECT 80.780 105.805 80.900 105.915 ;
        RECT 77.110 105.755 77.280 105.775 ;
        RECT 81.245 105.755 81.415 105.945 ;
        RECT 84.460 105.805 84.580 105.915 ;
        RECT 84.925 105.775 85.095 105.965 ;
        RECT 88.140 105.805 88.260 105.915 ;
        RECT 89.525 105.755 89.695 105.965 ;
        RECT 50.720 105.725 51.655 105.755 ;
        RECT 48.590 105.525 51.655 105.725 ;
        RECT 44.600 104.855 45.510 105.075 ;
        RECT 47.045 104.845 48.395 105.075 ;
        RECT 48.445 105.045 51.655 105.525 ;
        RECT 51.665 105.075 58.975 105.755 ;
        RECT 48.445 104.845 49.375 105.045 ;
        RECT 50.705 104.845 51.655 105.045 ;
        RECT 55.180 104.855 56.090 105.075 ;
        RECT 57.625 104.845 58.975 105.075 ;
        RECT 59.505 104.845 60.855 105.755 ;
        RECT 60.875 104.845 63.605 105.755 ;
        RECT 63.635 104.885 64.065 105.670 ;
        RECT 64.085 104.845 65.435 105.755 ;
        RECT 65.925 104.845 69.135 105.755 ;
        RECT 69.145 105.075 73.045 105.755 ;
        RECT 73.380 105.075 76.845 105.755 ;
        RECT 69.145 104.845 70.075 105.075 ;
        RECT 73.380 104.845 74.300 105.075 ;
        RECT 76.965 104.845 80.440 105.755 ;
        RECT 81.105 105.075 88.415 105.755 ;
        RECT 84.620 104.855 85.530 105.075 ;
        RECT 87.065 104.845 88.415 105.075 ;
        RECT 88.465 104.945 89.835 105.755 ;
        RECT 103.720 105.090 106.510 107.170 ;
      LAYER nwell ;
        RECT 11.910 101.725 90.030 104.555 ;
        RECT 101.610 102.980 106.450 105.090 ;
        RECT 107.730 104.750 117.920 117.000 ;
      LAYER pwell ;
        RECT 120.330 107.200 126.430 116.990 ;
        RECT 120.330 107.170 126.440 107.200 ;
        RECT 120.530 106.770 121.690 107.170 ;
        RECT 123.650 105.090 126.440 107.170 ;
      LAYER nwell ;
        RECT 121.540 102.980 126.380 105.090 ;
        RECT 127.660 104.750 137.850 117.000 ;
      LAYER pwell ;
        RECT 140.360 107.200 146.460 116.990 ;
        RECT 140.360 107.170 146.470 107.200 ;
        RECT 140.560 106.770 141.720 107.170 ;
        RECT 143.680 105.090 146.470 107.170 ;
      LAYER nwell ;
        RECT 141.570 102.980 146.410 105.090 ;
        RECT 147.690 104.750 157.880 117.000 ;
      LAYER pwell ;
        RECT 12.105 100.525 13.475 101.335 ;
        RECT 13.485 100.525 18.995 101.335 ;
        RECT 19.005 100.525 24.515 101.335 ;
        RECT 24.995 100.610 25.425 101.395 ;
        RECT 25.445 100.525 30.955 101.335 ;
        RECT 30.965 100.525 34.635 101.335 ;
        RECT 34.645 100.525 36.015 101.335 ;
        RECT 36.045 100.525 37.395 101.435 ;
        RECT 40.060 101.205 40.980 101.435 ;
        RECT 37.515 100.525 40.980 101.205 ;
        RECT 41.125 101.205 42.475 101.435 ;
        RECT 44.010 101.205 44.920 101.425 ;
        RECT 41.125 100.525 48.435 101.205 ;
        RECT 48.545 100.525 50.735 101.435 ;
        RECT 50.755 100.610 51.185 101.395 ;
        RECT 51.205 101.205 52.135 101.435 ;
        RECT 56.705 101.205 57.635 101.435 ;
        RECT 59.465 101.205 60.395 101.435 ;
        RECT 51.205 100.525 54.875 101.205 ;
        RECT 54.885 100.525 57.635 101.205 ;
        RECT 57.645 100.525 60.395 101.205 ;
        RECT 61.475 100.525 65.130 101.435 ;
        RECT 65.485 100.525 66.835 101.435 ;
        RECT 71.280 101.205 72.190 101.425 ;
        RECT 73.725 101.205 75.075 101.435 ;
        RECT 67.765 100.525 75.075 101.205 ;
        RECT 75.125 100.525 76.495 101.305 ;
        RECT 76.515 100.610 76.945 101.395 ;
        RECT 77.885 100.525 81.095 101.435 ;
        RECT 81.105 100.525 84.580 101.435 ;
        RECT 84.785 100.525 87.995 101.435 ;
        RECT 88.465 100.525 89.835 101.335 ;
        RECT 12.245 100.315 12.415 100.525 ;
        RECT 13.625 100.315 13.795 100.525 ;
        RECT 17.315 100.360 17.475 100.470 ;
        RECT 18.230 100.315 18.400 100.505 ;
        RECT 19.145 100.335 19.315 100.525 ;
        RECT 19.605 100.315 19.775 100.505 ;
        RECT 24.660 100.365 24.780 100.475 ;
        RECT 25.135 100.360 25.295 100.470 ;
        RECT 25.585 100.335 25.755 100.525 ;
        RECT 31.105 100.335 31.275 100.525 ;
        RECT 34.785 100.335 34.955 100.525 ;
        RECT 35.705 100.315 35.875 100.505 ;
        RECT 36.165 100.315 36.335 100.505 ;
        RECT 37.080 100.335 37.250 100.525 ;
        RECT 37.545 100.335 37.715 100.525 ;
        RECT 38.460 100.315 38.630 100.505 ;
        RECT 40.765 100.315 40.935 100.505 ;
        RECT 41.235 100.360 41.395 100.470 ;
        RECT 42.145 100.315 42.315 100.505 ;
        RECT 48.125 100.335 48.295 100.525 ;
        RECT 49.505 100.315 49.675 100.505 ;
        RECT 50.420 100.335 50.590 100.525 ;
        RECT 52.275 100.360 52.435 100.470 ;
        RECT 53.190 100.315 53.360 100.505 ;
        RECT 54.565 100.335 54.735 100.525 ;
        RECT 55.025 100.335 55.195 100.525 ;
        RECT 57.785 100.505 57.955 100.525 ;
        RECT 61.475 100.505 61.635 100.525 ;
        RECT 55.485 100.315 55.655 100.505 ;
        RECT 57.785 100.335 57.960 100.505 ;
        RECT 60.095 100.360 60.255 100.470 ;
        RECT 60.555 100.370 60.715 100.480 ;
        RECT 61.465 100.335 61.635 100.505 ;
        RECT 57.790 100.315 57.960 100.335 ;
        RECT 63.305 100.315 63.475 100.505 ;
        RECT 64.225 100.315 64.395 100.505 ;
        RECT 65.600 100.335 65.770 100.525 ;
        RECT 66.065 100.315 66.235 100.505 ;
        RECT 66.995 100.370 67.155 100.480 ;
        RECT 67.905 100.335 68.075 100.525 ;
        RECT 76.185 100.335 76.355 100.525 ;
        RECT 76.645 100.315 76.815 100.505 ;
        RECT 77.115 100.370 77.275 100.480 ;
        RECT 78.015 100.335 78.185 100.525 ;
        RECT 78.485 100.315 78.655 100.505 ;
        RECT 78.945 100.315 79.115 100.505 ;
        RECT 81.250 100.335 81.420 100.525 ;
        RECT 86.305 100.335 86.475 100.505 ;
        RECT 87.685 100.335 87.855 100.525 ;
        RECT 88.140 100.365 88.260 100.475 ;
        RECT 86.310 100.315 86.475 100.335 ;
        RECT 89.525 100.315 89.695 100.525 ;
        RECT 12.105 99.505 13.475 100.315 ;
        RECT 13.485 99.505 17.155 100.315 ;
        RECT 18.085 99.405 19.435 100.315 ;
        RECT 19.465 99.505 24.975 100.315 ;
        RECT 25.940 99.405 35.960 100.315 ;
        RECT 36.025 99.505 37.855 100.315 ;
        RECT 37.875 99.445 38.305 100.230 ;
        RECT 38.345 99.405 39.695 100.315 ;
        RECT 39.715 99.405 41.065 100.315 ;
        RECT 42.005 99.635 49.315 100.315 ;
        RECT 49.365 99.635 52.115 100.315 ;
        RECT 45.520 99.415 46.430 99.635 ;
        RECT 47.965 99.405 49.315 99.635 ;
        RECT 51.185 99.405 52.115 99.635 ;
        RECT 53.045 99.405 55.235 100.315 ;
        RECT 55.345 99.635 57.635 100.315 ;
        RECT 57.645 99.635 59.920 100.315 ;
        RECT 56.715 99.405 57.635 99.635 ;
        RECT 58.550 99.405 59.920 99.635 ;
        RECT 60.875 99.405 63.605 100.315 ;
        RECT 63.635 99.445 64.065 100.230 ;
        RECT 64.085 99.505 65.915 100.315 ;
        RECT 65.925 99.635 73.235 100.315 ;
        RECT 69.440 99.415 70.350 99.635 ;
        RECT 71.885 99.405 73.235 99.635 ;
        RECT 73.380 99.635 76.845 100.315 ;
        RECT 76.965 99.635 78.795 100.315 ;
        RECT 78.805 99.635 86.115 100.315 ;
        RECT 86.310 99.635 88.145 100.315 ;
        RECT 73.380 99.405 74.300 99.635 ;
        RECT 76.965 99.405 78.310 99.635 ;
        RECT 82.320 99.415 83.230 99.635 ;
        RECT 84.765 99.405 86.115 99.635 ;
        RECT 87.215 99.405 88.145 99.635 ;
        RECT 88.465 99.505 89.835 100.315 ;
      LAYER nwell ;
        RECT 11.910 96.285 90.030 99.115 ;
      LAYER pwell ;
        RECT 12.105 95.085 13.475 95.895 ;
        RECT 13.485 95.765 14.405 95.995 ;
        RECT 15.785 95.765 16.705 95.995 ;
        RECT 13.485 95.085 15.775 95.765 ;
        RECT 15.785 95.085 18.075 95.765 ;
        RECT 18.565 95.085 19.915 95.995 ;
        RECT 22.670 95.765 23.595 95.995 ;
        RECT 19.925 95.085 23.595 95.765 ;
        RECT 23.605 95.085 24.955 95.995 ;
        RECT 24.995 95.170 25.425 95.955 ;
        RECT 25.455 95.085 26.805 95.995 ;
        RECT 26.825 95.085 28.655 95.895 ;
        RECT 29.435 95.765 30.365 95.995 ;
        RECT 29.435 95.085 31.270 95.765 ;
        RECT 32.345 95.315 34.180 95.995 ;
        RECT 12.245 94.875 12.415 95.085 ;
        RECT 13.635 94.920 13.795 95.030 ;
        RECT 14.545 94.875 14.715 95.065 ;
        RECT 15.465 94.895 15.635 95.085 ;
        RECT 17.765 94.895 17.935 95.085 ;
        RECT 18.220 94.925 18.340 95.035 ;
        RECT 19.600 94.895 19.770 95.085 ;
        RECT 21.900 94.925 22.020 95.035 ;
        RECT 23.280 94.875 23.450 95.085 ;
        RECT 23.745 94.875 23.915 95.065 ;
        RECT 24.670 94.895 24.840 95.085 ;
        RECT 25.585 94.895 25.755 95.085 ;
        RECT 26.965 94.895 27.135 95.085 ;
        RECT 31.105 95.065 31.270 95.085 ;
        RECT 32.490 95.085 34.180 95.315 ;
        RECT 34.645 95.085 40.155 95.895 ;
        RECT 40.165 95.085 42.915 95.895 ;
        RECT 42.925 95.085 44.275 95.995 ;
        RECT 44.305 95.085 47.515 95.995 ;
        RECT 47.525 95.085 50.275 95.995 ;
        RECT 50.755 95.170 51.185 95.955 ;
        RECT 51.205 95.085 60.310 95.765 ;
        RECT 60.405 95.085 65.915 95.895 ;
        RECT 65.925 95.085 67.755 95.895 ;
        RECT 67.765 95.765 68.695 95.995 ;
        RECT 67.765 95.085 71.665 95.765 ;
        RECT 71.905 95.085 73.275 95.895 ;
        RECT 73.285 95.085 76.495 95.995 ;
        RECT 76.515 95.170 76.945 95.955 ;
        RECT 76.965 95.085 78.335 95.865 ;
        RECT 78.345 95.085 81.820 95.995 ;
        RECT 82.335 95.765 83.265 95.995 ;
        RECT 85.375 95.765 86.305 95.995 ;
        RECT 82.335 95.085 84.170 95.765 ;
        RECT 32.490 95.065 32.660 95.085 ;
        RECT 28.800 94.925 28.920 95.035 ;
        RECT 31.105 94.875 31.275 95.065 ;
        RECT 31.575 94.930 31.735 95.040 ;
        RECT 32.485 94.895 32.660 95.065 ;
        RECT 34.785 94.895 34.955 95.085 ;
        RECT 32.485 94.875 32.655 94.895 ;
        RECT 37.085 94.875 37.255 95.065 ;
        RECT 37.540 94.925 37.660 95.035 ;
        RECT 38.465 94.875 38.635 95.065 ;
        RECT 40.305 94.895 40.475 95.085 ;
        RECT 43.070 94.895 43.240 95.085 ;
        RECT 43.985 94.875 44.155 95.065 ;
        RECT 47.205 94.895 47.375 95.085 ;
        RECT 47.665 94.875 47.835 95.085 ;
        RECT 12.105 94.065 13.475 94.875 ;
        RECT 14.405 94.195 21.715 94.875 ;
        RECT 17.920 93.975 18.830 94.195 ;
        RECT 20.365 93.965 21.715 94.195 ;
        RECT 22.245 93.965 23.595 94.875 ;
        RECT 23.605 94.195 30.915 94.875 ;
        RECT 27.120 93.975 28.030 94.195 ;
        RECT 29.565 93.965 30.915 94.195 ;
        RECT 30.965 94.065 32.335 94.875 ;
        RECT 32.345 94.195 34.635 94.875 ;
        RECT 33.715 93.965 34.635 94.195 ;
        RECT 34.655 93.965 37.385 94.875 ;
        RECT 37.875 94.005 38.305 94.790 ;
        RECT 38.325 94.065 43.835 94.875 ;
        RECT 43.845 94.065 47.515 94.875 ;
        RECT 47.525 94.065 48.895 94.875 ;
        RECT 49.040 94.845 49.210 95.065 ;
        RECT 50.420 94.925 50.540 95.035 ;
        RECT 51.345 94.895 51.515 95.085 ;
        RECT 52.265 94.875 52.435 95.065 ;
        RECT 54.560 94.875 54.730 95.065 ;
        RECT 55.025 94.875 55.195 95.065 ;
        RECT 56.410 94.875 56.580 95.065 ;
        RECT 58.710 94.875 58.880 95.065 ;
        RECT 60.545 94.895 60.715 95.085 ;
        RECT 61.010 94.875 61.180 95.065 ;
        RECT 63.300 94.925 63.420 95.035 ;
        RECT 64.225 94.875 64.395 95.065 ;
        RECT 66.065 94.895 66.235 95.085 ;
        RECT 68.180 94.895 68.350 95.085 ;
        RECT 69.745 94.875 69.915 95.065 ;
        RECT 72.045 94.895 72.215 95.085 ;
        RECT 72.965 94.875 73.135 95.065 ;
        RECT 74.805 94.875 74.975 95.065 ;
        RECT 76.185 94.895 76.355 95.085 ;
        RECT 76.645 94.875 76.815 95.065 ;
        RECT 77.105 94.895 77.275 95.085 ;
        RECT 78.490 94.895 78.660 95.085 ;
        RECT 84.005 95.065 84.170 95.085 ;
        RECT 84.470 95.085 86.305 95.765 ;
        RECT 86.625 95.765 87.970 95.995 ;
        RECT 86.625 95.085 88.455 95.765 ;
        RECT 88.465 95.085 89.835 95.895 ;
        RECT 84.470 95.065 84.635 95.085 ;
        RECT 77.110 94.875 77.275 94.895 ;
        RECT 81.240 94.875 81.410 95.065 ;
        RECT 81.705 94.875 81.875 95.065 ;
        RECT 83.540 94.925 83.660 95.035 ;
        RECT 84.005 94.895 84.175 95.065 ;
        RECT 84.465 94.895 84.635 95.065 ;
        RECT 86.765 94.875 86.935 95.065 ;
        RECT 87.225 94.875 87.395 95.065 ;
        RECT 88.145 94.895 88.315 95.085 ;
        RECT 89.525 94.875 89.695 95.085 ;
        RECT 50.240 94.845 51.195 94.875 ;
        RECT 48.915 94.165 51.195 94.845 ;
        RECT 50.240 93.965 51.195 94.165 ;
        RECT 51.215 93.965 52.565 94.875 ;
        RECT 53.040 94.645 54.730 94.875 ;
        RECT 53.040 93.965 54.875 94.645 ;
        RECT 54.885 94.065 56.255 94.875 ;
        RECT 56.265 94.195 58.540 94.875 ;
        RECT 57.170 93.965 58.540 94.195 ;
        RECT 58.565 93.965 60.775 94.875 ;
        RECT 60.865 93.965 63.075 94.875 ;
        RECT 63.635 94.005 64.065 94.790 ;
        RECT 64.085 94.065 69.595 94.875 ;
        RECT 69.605 94.065 71.435 94.875 ;
        RECT 71.445 94.195 73.275 94.875 ;
        RECT 73.285 94.195 75.115 94.875 ;
        RECT 75.125 94.195 76.955 94.875 ;
        RECT 77.110 94.195 78.945 94.875 ;
        RECT 71.445 93.965 72.790 94.195 ;
        RECT 73.285 93.965 74.630 94.195 ;
        RECT 75.125 93.965 76.470 94.195 ;
        RECT 78.015 93.965 78.945 94.195 ;
        RECT 79.365 93.965 81.555 94.875 ;
        RECT 81.565 94.195 83.395 94.875 ;
        RECT 82.050 93.965 83.395 94.195 ;
        RECT 83.865 93.965 87.075 94.875 ;
        RECT 87.085 94.065 88.455 94.875 ;
        RECT 88.465 94.065 89.835 94.875 ;
      LAYER nwell ;
        RECT 11.910 90.845 90.030 93.675 ;
        RECT 99.800 92.735 112.970 100.575 ;
      LAYER pwell ;
        RECT 134.270 96.400 158.480 102.920 ;
        RECT 12.105 89.645 13.475 90.455 ;
        RECT 17.000 90.325 17.910 90.545 ;
        RECT 19.445 90.325 20.795 90.555 ;
        RECT 23.840 90.325 24.975 90.555 ;
        RECT 13.485 89.645 20.795 90.325 ;
        RECT 21.765 89.645 24.975 90.325 ;
        RECT 24.995 89.730 25.425 90.515 ;
        RECT 25.445 89.645 28.655 90.555 ;
        RECT 28.675 89.645 31.415 90.325 ;
        RECT 31.445 89.645 32.795 90.555 ;
        RECT 36.320 90.325 37.230 90.545 ;
        RECT 38.765 90.325 40.115 90.555 ;
        RECT 32.805 89.645 40.115 90.325 ;
        RECT 40.205 90.325 41.555 90.555 ;
        RECT 43.090 90.325 44.000 90.545 ;
        RECT 40.205 89.645 47.515 90.325 ;
        RECT 47.525 89.645 50.275 90.455 ;
        RECT 50.755 89.730 51.185 90.515 ;
        RECT 51.205 89.645 53.035 90.455 ;
        RECT 53.065 89.645 54.415 90.555 ;
        RECT 55.795 90.325 56.715 90.555 ;
        RECT 54.425 89.645 56.715 90.325 ;
        RECT 57.185 90.355 58.140 90.555 ;
        RECT 57.185 89.675 59.465 90.355 ;
        RECT 57.185 89.645 58.140 89.675 ;
        RECT 12.245 89.435 12.415 89.645 ;
        RECT 13.625 89.435 13.795 89.645 ;
        RECT 20.995 89.490 21.155 89.600 ;
        RECT 21.905 89.455 22.075 89.645 ;
        RECT 23.745 89.435 23.915 89.625 ;
        RECT 25.585 89.455 25.755 89.645 ;
        RECT 26.045 89.455 26.215 89.625 ;
        RECT 26.045 89.435 26.210 89.455 ;
        RECT 28.340 89.435 28.510 89.625 ;
        RECT 30.645 89.455 30.815 89.625 ;
        RECT 31.105 89.595 31.275 89.645 ;
        RECT 31.100 89.485 31.275 89.595 ;
        RECT 31.105 89.455 31.275 89.485 ;
        RECT 31.560 89.625 31.730 89.645 ;
        RECT 31.560 89.455 31.735 89.625 ;
        RECT 32.945 89.455 33.115 89.645 ;
        RECT 30.645 89.435 30.795 89.455 ;
        RECT 31.565 89.435 31.735 89.455 ;
        RECT 12.105 88.625 13.475 89.435 ;
        RECT 13.485 88.755 20.795 89.435 ;
        RECT 17.000 88.535 17.910 88.755 ;
        RECT 19.445 88.525 20.795 88.755 ;
        RECT 20.845 88.755 24.055 89.435 ;
        RECT 24.375 88.755 26.210 89.435 ;
        RECT 26.820 89.205 28.510 89.435 ;
        RECT 20.845 88.525 21.980 88.755 ;
        RECT 24.375 88.525 25.305 88.755 ;
        RECT 26.820 88.525 28.655 89.205 ;
        RECT 28.865 88.615 30.795 89.435 ;
        RECT 31.425 88.755 33.715 89.435 ;
        RECT 33.870 89.405 34.040 89.625 ;
        RECT 37.095 89.480 37.255 89.590 ;
        RECT 38.465 89.435 38.635 89.625 ;
        RECT 36.000 89.405 36.935 89.435 ;
        RECT 33.870 89.205 36.935 89.405 ;
        RECT 28.865 88.525 29.815 88.615 ;
        RECT 32.795 88.525 33.715 88.755 ;
        RECT 33.725 88.725 36.935 89.205 ;
        RECT 33.725 88.525 34.655 88.725 ;
        RECT 35.985 88.525 36.935 88.725 ;
        RECT 37.875 88.565 38.305 89.350 ;
        RECT 38.325 88.625 39.695 89.435 ;
        RECT 39.850 89.405 40.020 89.625 ;
        RECT 43.065 89.455 43.235 89.625 ;
        RECT 43.070 89.435 43.235 89.455 ;
        RECT 45.365 89.435 45.535 89.625 ;
        RECT 47.205 89.455 47.375 89.645 ;
        RECT 47.665 89.455 47.835 89.645 ;
        RECT 51.345 89.625 51.515 89.645 ;
        RECT 49.045 89.435 49.215 89.625 ;
        RECT 50.420 89.485 50.540 89.595 ;
        RECT 51.340 89.455 51.515 89.625 ;
        RECT 53.180 89.625 53.350 89.645 ;
        RECT 53.180 89.455 53.355 89.625 ;
        RECT 51.340 89.435 51.510 89.455 ;
        RECT 53.185 89.435 53.355 89.455 ;
        RECT 53.645 89.435 53.815 89.625 ;
        RECT 54.565 89.455 54.735 89.645 ;
        RECT 59.170 89.625 59.340 89.675 ;
        RECT 59.485 89.645 61.315 90.555 ;
        RECT 62.375 90.325 63.305 90.555 ;
        RECT 61.470 89.645 63.305 90.325 ;
        RECT 63.625 89.645 69.135 90.455 ;
        RECT 69.145 89.645 70.975 90.455 ;
        RECT 71.455 89.645 72.805 90.555 ;
        RECT 73.020 89.645 76.495 90.555 ;
        RECT 76.515 89.730 76.945 90.515 ;
        RECT 80.480 90.325 81.390 90.545 ;
        RECT 82.925 90.325 84.275 90.555 ;
        RECT 76.965 89.645 84.275 90.325 ;
        RECT 84.325 89.645 87.800 90.555 ;
        RECT 88.465 89.645 89.835 90.455 ;
        RECT 56.860 89.485 56.980 89.595 ;
        RECT 41.980 89.405 42.915 89.435 ;
        RECT 39.850 89.205 42.915 89.405 ;
        RECT 39.705 88.725 42.915 89.205 ;
        RECT 43.070 88.755 44.905 89.435 ;
        RECT 39.705 88.525 40.635 88.725 ;
        RECT 41.965 88.525 42.915 88.725 ;
        RECT 43.975 88.525 44.905 88.755 ;
        RECT 45.225 88.625 48.895 89.435 ;
        RECT 48.905 88.625 50.275 89.435 ;
        RECT 50.305 88.525 51.655 89.435 ;
        RECT 51.665 88.755 53.495 89.435 ;
        RECT 51.665 88.525 53.010 88.755 ;
        RECT 53.585 88.525 56.585 89.435 ;
        RECT 56.725 89.405 57.680 89.435 ;
        RECT 58.710 89.405 58.880 89.625 ;
        RECT 59.160 89.455 59.340 89.625 ;
        RECT 59.630 89.455 59.800 89.645 ;
        RECT 61.470 89.625 61.635 89.645 ;
        RECT 59.160 89.405 59.330 89.455 ;
        RECT 61.465 89.435 61.635 89.625 ;
        RECT 63.765 89.455 63.935 89.645 ;
        RECT 66.065 89.435 66.235 89.625 ;
        RECT 66.525 89.435 66.695 89.625 ;
        RECT 67.905 89.435 68.075 89.625 ;
        RECT 69.285 89.455 69.455 89.645 ;
        RECT 70.665 89.435 70.835 89.625 ;
        RECT 71.130 89.595 71.300 89.625 ;
        RECT 71.120 89.485 71.300 89.595 ;
        RECT 71.130 89.435 71.300 89.485 ;
        RECT 72.505 89.455 72.675 89.645 ;
        RECT 73.430 89.435 73.600 89.625 ;
        RECT 75.735 89.480 75.895 89.590 ;
        RECT 76.180 89.455 76.350 89.645 ;
        RECT 77.105 89.455 77.275 89.645 ;
        RECT 78.485 89.455 78.655 89.625 ;
        RECT 80.785 89.455 80.955 89.625 ;
        RECT 78.485 89.435 78.650 89.455 ;
        RECT 80.785 89.435 80.935 89.455 ;
        RECT 81.245 89.435 81.415 89.625 ;
        RECT 84.470 89.455 84.640 89.645 ;
        RECT 88.140 89.485 88.260 89.595 ;
        RECT 89.525 89.435 89.695 89.645 ;
        RECT 60.360 89.405 61.315 89.435 ;
        RECT 56.725 88.725 59.005 89.405 ;
        RECT 59.035 88.725 61.315 89.405 ;
        RECT 61.325 88.755 63.615 89.435 ;
        RECT 56.725 88.525 57.680 88.725 ;
        RECT 60.360 88.525 61.315 88.725 ;
        RECT 62.695 88.525 63.615 88.755 ;
        RECT 63.635 88.565 64.065 89.350 ;
        RECT 64.085 88.755 66.375 89.435 ;
        RECT 64.085 88.525 65.005 88.755 ;
        RECT 66.385 88.625 67.755 89.435 ;
        RECT 67.775 88.525 69.125 89.435 ;
        RECT 69.145 88.755 70.975 89.435 ;
        RECT 70.985 88.755 73.260 89.435 ;
        RECT 69.145 88.525 70.490 88.755 ;
        RECT 71.890 88.525 73.260 88.755 ;
        RECT 73.285 88.525 75.495 89.435 ;
        RECT 76.815 88.755 78.650 89.435 ;
        RECT 76.815 88.525 77.745 88.755 ;
        RECT 79.005 88.615 80.935 89.435 ;
        RECT 81.105 88.755 88.415 89.435 ;
        RECT 79.005 88.525 79.955 88.615 ;
        RECT 84.620 88.535 85.530 88.755 ;
        RECT 87.065 88.525 88.415 88.755 ;
        RECT 88.465 88.625 89.835 89.435 ;
        RECT 99.810 88.235 112.980 92.025 ;
      LAYER nwell ;
        RECT 11.910 85.405 90.030 88.235 ;
      LAYER pwell ;
        RECT 12.105 84.205 13.475 85.015 ;
        RECT 14.405 84.915 15.355 85.115 ;
        RECT 16.685 84.915 17.615 85.115 ;
        RECT 14.405 84.435 17.615 84.915 ;
        RECT 18.545 84.915 19.475 85.115 ;
        RECT 20.810 84.915 21.755 85.115 ;
        RECT 18.545 84.435 21.755 84.915 ;
        RECT 21.765 84.915 22.695 85.115 ;
        RECT 24.025 84.915 24.975 85.115 ;
        RECT 21.765 84.435 24.975 84.915 ;
        RECT 14.405 84.235 17.470 84.435 ;
        RECT 14.405 84.205 15.340 84.235 ;
        RECT 12.245 83.995 12.415 84.205 ;
        RECT 13.625 83.995 13.795 84.185 ;
        RECT 17.300 83.995 17.470 84.235 ;
        RECT 18.685 84.235 21.755 84.435 ;
        RECT 17.765 83.995 17.935 84.185 ;
        RECT 18.685 84.015 18.855 84.235 ;
        RECT 20.810 84.205 21.755 84.235 ;
        RECT 21.910 84.235 24.975 84.435 ;
        RECT 24.995 84.290 25.425 85.075 ;
        RECT 20.060 83.995 20.230 84.185 ;
        RECT 20.525 83.995 20.695 84.185 ;
        RECT 21.910 84.015 22.080 84.235 ;
        RECT 24.040 84.205 24.975 84.235 ;
        RECT 25.640 84.205 29.115 85.115 ;
        RECT 29.125 84.205 31.415 85.115 ;
        RECT 31.445 84.205 32.795 85.115 ;
        RECT 34.035 84.885 34.965 85.115 ;
        RECT 34.035 84.205 35.870 84.885 ;
        RECT 36.025 84.205 39.680 85.115 ;
        RECT 39.745 84.885 41.095 85.115 ;
        RECT 42.630 84.885 43.540 85.105 ;
        RECT 47.065 84.915 48.015 85.115 ;
        RECT 49.345 84.915 50.275 85.115 ;
        RECT 39.745 84.205 47.055 84.885 ;
        RECT 47.065 84.435 50.275 84.915 ;
        RECT 47.065 84.235 50.130 84.435 ;
        RECT 50.755 84.290 51.185 85.075 ;
        RECT 47.065 84.205 48.000 84.235 ;
        RECT 26.045 83.995 26.215 84.185 ;
        RECT 28.800 84.015 28.970 84.205 ;
        RECT 29.265 84.015 29.435 84.205 ;
        RECT 29.725 83.995 29.895 84.185 ;
        RECT 31.560 84.015 31.730 84.205 ;
        RECT 35.705 84.185 35.870 84.205 ;
        RECT 32.945 84.015 33.115 84.185 ;
        RECT 33.405 84.015 33.575 84.185 ;
        RECT 35.705 84.015 35.875 84.185 ;
        RECT 36.170 84.015 36.340 84.205 ;
        RECT 38.460 84.045 38.580 84.155 ;
        RECT 32.945 83.995 33.110 84.015 ;
        RECT 12.105 83.185 13.475 83.995 ;
        RECT 13.485 83.185 16.235 83.995 ;
        RECT 16.265 83.085 17.615 83.995 ;
        RECT 17.625 83.185 18.995 83.995 ;
        RECT 19.025 83.085 20.375 83.995 ;
        RECT 20.385 83.185 25.895 83.995 ;
        RECT 25.905 83.185 29.575 83.995 ;
        RECT 29.585 83.185 30.955 83.995 ;
        RECT 31.275 83.315 33.110 83.995 ;
        RECT 33.425 83.995 33.575 84.015 ;
        RECT 35.710 83.995 35.875 84.015 ;
        RECT 38.925 83.995 39.095 84.185 ;
        RECT 46.285 83.995 46.455 84.185 ;
        RECT 46.745 84.015 46.915 84.205 ;
        RECT 47.665 83.995 47.835 84.185 ;
        RECT 49.960 84.015 50.130 84.235 ;
        RECT 51.205 84.205 53.035 85.115 ;
        RECT 53.045 84.205 56.255 85.115 ;
        RECT 56.275 84.205 57.625 85.115 ;
        RECT 57.840 84.205 61.315 85.115 ;
        RECT 62.395 84.205 66.050 85.115 ;
        RECT 66.385 84.205 69.595 85.115 ;
        RECT 70.655 84.885 71.585 85.115 ;
        RECT 74.165 84.915 75.575 85.115 ;
        RECT 69.750 84.205 71.585 84.885 ;
        RECT 72.840 84.235 75.575 84.915 ;
        RECT 76.515 84.290 76.945 85.075 ;
        RECT 78.305 84.915 79.715 85.115 ;
        RECT 76.980 84.235 79.715 84.915 ;
        RECT 50.420 84.045 50.540 84.155 ;
        RECT 51.350 84.015 51.520 84.205 ;
        RECT 53.185 84.015 53.355 84.205 ;
        RECT 55.030 83.995 55.200 84.185 ;
        RECT 56.405 84.015 56.575 84.205 ;
        RECT 58.700 83.995 58.870 84.185 ;
        RECT 61.000 84.015 61.170 84.205 ;
        RECT 62.395 84.185 62.555 84.205 ;
        RECT 61.475 84.050 61.635 84.160 ;
        RECT 62.385 84.015 62.555 84.185 ;
        RECT 63.300 83.995 63.470 84.185 ;
        RECT 64.225 83.995 64.395 84.185 ;
        RECT 66.525 84.015 66.695 84.205 ;
        RECT 69.750 84.185 69.915 84.205 ;
        RECT 67.720 83.995 67.890 84.185 ;
        RECT 69.745 84.015 69.915 84.185 ;
        RECT 72.055 84.050 72.215 84.160 ;
        RECT 72.965 84.015 73.135 84.235 ;
        RECT 74.180 84.205 75.575 84.235 ;
        RECT 74.805 83.995 74.975 84.185 ;
        RECT 75.260 84.045 75.380 84.155 ;
        RECT 75.725 84.015 75.895 84.185 ;
        RECT 77.105 84.015 77.275 84.235 ;
        RECT 78.320 84.205 79.715 84.235 ;
        RECT 79.725 84.205 81.915 85.115 ;
        RECT 82.025 84.205 85.235 85.115 ;
        RECT 85.245 84.205 88.455 85.115 ;
        RECT 88.465 84.205 89.835 85.015 ;
        RECT 75.755 83.995 75.895 84.015 ;
        RECT 78.490 83.995 78.660 84.185 ;
        RECT 79.870 84.015 80.040 84.205 ;
        RECT 82.155 84.185 82.325 84.205 ;
        RECT 82.155 84.015 82.340 84.185 ;
        RECT 82.170 83.995 82.340 84.015 ;
        RECT 87.685 84.015 87.855 84.185 ;
        RECT 88.145 84.155 88.315 84.205 ;
        RECT 88.140 84.045 88.315 84.155 ;
        RECT 88.145 84.015 88.315 84.045 ;
        RECT 87.685 83.995 87.850 84.015 ;
        RECT 89.525 83.995 89.695 84.205 ;
        RECT 31.275 83.085 32.205 83.315 ;
        RECT 33.425 83.175 35.355 83.995 ;
        RECT 35.710 83.315 37.545 83.995 ;
        RECT 34.405 83.085 35.355 83.175 ;
        RECT 36.615 83.085 37.545 83.315 ;
        RECT 37.875 83.125 38.305 83.910 ;
        RECT 38.785 83.315 46.095 83.995 ;
        RECT 42.300 83.095 43.210 83.315 ;
        RECT 44.745 83.085 46.095 83.315 ;
        RECT 46.145 83.185 47.515 83.995 ;
        RECT 47.525 83.315 54.835 83.995 ;
        RECT 51.040 83.095 51.950 83.315 ;
        RECT 53.485 83.085 54.835 83.315 ;
        RECT 54.885 83.085 58.555 83.995 ;
        RECT 58.585 83.085 59.935 83.995 ;
        RECT 60.140 83.085 63.615 83.995 ;
        RECT 63.635 83.125 64.065 83.910 ;
        RECT 64.085 83.085 67.295 83.995 ;
        RECT 67.305 83.315 71.205 83.995 ;
        RECT 71.540 83.315 75.005 83.995 ;
        RECT 67.305 83.085 68.235 83.315 ;
        RECT 71.540 83.085 72.460 83.315 ;
        RECT 75.755 83.175 78.325 83.995 ;
        RECT 76.735 83.085 78.325 83.175 ;
        RECT 78.345 83.085 81.820 83.995 ;
        RECT 82.025 83.085 85.500 83.995 ;
        RECT 86.015 83.315 87.850 83.995 ;
        RECT 86.015 83.085 86.945 83.315 ;
        RECT 88.465 83.185 89.835 83.995 ;
      LAYER nwell ;
        RECT 11.910 79.965 90.030 82.795 ;
      LAYER pwell ;
        RECT 99.810 80.745 113.660 87.965 ;
        RECT 12.105 78.765 13.475 79.575 ;
        RECT 13.485 78.765 18.995 79.575 ;
        RECT 19.005 78.765 22.675 79.575 ;
        RECT 23.155 78.765 24.505 79.675 ;
        RECT 24.995 78.850 25.425 79.635 ;
        RECT 25.445 78.765 27.275 79.575 ;
        RECT 27.805 78.765 29.575 79.675 ;
        RECT 29.635 78.765 32.795 79.675 ;
        RECT 32.805 78.765 35.555 79.675 ;
        RECT 35.565 78.765 38.315 79.675 ;
        RECT 38.795 78.765 41.525 79.675 ;
        RECT 41.545 78.765 43.375 79.575 ;
        RECT 47.090 79.445 50.700 79.675 ;
        RECT 43.790 78.765 46.215 79.445 ;
        RECT 46.605 78.765 50.700 79.445 ;
        RECT 50.755 78.850 51.185 79.635 ;
        RECT 51.205 79.445 52.135 79.675 ;
        RECT 51.205 78.765 55.105 79.445 ;
        RECT 55.345 78.765 56.715 79.575 ;
        RECT 56.725 79.475 57.655 79.675 ;
        RECT 58.985 79.475 59.935 79.675 ;
        RECT 61.280 79.475 62.235 79.675 ;
        RECT 56.725 78.995 59.935 79.475 ;
        RECT 56.870 78.795 59.935 78.995 ;
        RECT 59.955 78.795 62.235 79.475 ;
        RECT 12.245 78.555 12.415 78.765 ;
        RECT 13.625 78.555 13.795 78.765 ;
        RECT 15.460 78.605 15.580 78.715 ;
        RECT 16.850 78.555 17.020 78.745 ;
        RECT 17.305 78.555 17.475 78.745 ;
        RECT 19.145 78.575 19.315 78.765 ;
        RECT 22.820 78.710 22.940 78.715 ;
        RECT 22.820 78.605 22.995 78.710 ;
        RECT 22.835 78.600 22.995 78.605 ;
        RECT 23.285 78.575 23.455 78.765 ;
        RECT 23.740 78.555 23.910 78.745 ;
        RECT 24.660 78.605 24.780 78.715 ;
        RECT 25.125 78.555 25.295 78.745 ;
        RECT 25.585 78.575 25.755 78.765 ;
        RECT 27.425 78.715 27.595 78.745 ;
        RECT 27.420 78.605 27.595 78.715 ;
        RECT 27.425 78.575 27.595 78.605 ;
        RECT 29.260 78.575 29.430 78.765 ;
        RECT 29.725 78.575 29.895 78.765 ;
        RECT 32.945 78.575 33.115 78.765 ;
        RECT 35.705 78.575 35.875 78.765 ;
        RECT 41.225 78.745 41.395 78.765 ;
        RECT 27.445 78.555 27.595 78.575 ;
        RECT 36.625 78.555 36.795 78.745 ;
        RECT 37.095 78.600 37.255 78.710 ;
        RECT 38.460 78.605 38.580 78.715 ;
        RECT 41.220 78.575 41.395 78.745 ;
        RECT 41.220 78.555 41.390 78.575 ;
        RECT 41.685 78.555 41.855 78.765 ;
        RECT 46.750 78.745 46.920 78.765 ;
        RECT 43.525 78.575 43.695 78.745 ;
        RECT 46.745 78.575 46.920 78.745 ;
        RECT 51.620 78.575 51.790 78.765 ;
        RECT 46.745 78.555 46.915 78.575 ;
        RECT 54.105 78.555 54.275 78.745 ;
        RECT 55.485 78.575 55.655 78.765 ;
        RECT 56.870 78.575 57.040 78.795 ;
        RECT 59.000 78.765 59.935 78.795 ;
        RECT 57.325 78.575 57.495 78.745 ;
        RECT 57.795 78.600 57.955 78.710 ;
        RECT 58.705 78.575 58.875 78.745 ;
        RECT 60.080 78.575 60.250 78.795 ;
        RECT 61.280 78.765 62.235 78.795 ;
        RECT 62.245 78.765 65.455 79.675 ;
        RECT 68.980 79.445 69.890 79.665 ;
        RECT 71.425 79.445 72.775 79.675 ;
        RECT 73.875 79.445 74.805 79.675 ;
        RECT 65.465 78.765 72.775 79.445 ;
        RECT 72.970 78.765 74.805 79.445 ;
        RECT 75.135 78.765 76.485 79.675 ;
        RECT 76.515 78.850 76.945 79.635 ;
        RECT 76.965 78.765 78.735 79.675 ;
        RECT 82.320 79.445 83.230 79.665 ;
        RECT 84.765 79.445 86.115 79.675 ;
        RECT 87.215 79.445 88.145 79.675 ;
        RECT 78.805 78.765 86.115 79.445 ;
        RECT 86.310 78.765 88.145 79.445 ;
        RECT 88.465 78.765 89.835 79.575 ;
        RECT 57.325 78.555 57.490 78.575 ;
        RECT 12.105 77.745 13.475 78.555 ;
        RECT 13.485 77.745 15.315 78.555 ;
        RECT 15.785 77.645 17.135 78.555 ;
        RECT 17.165 77.745 22.675 78.555 ;
        RECT 23.625 77.645 24.975 78.555 ;
        RECT 24.985 77.875 27.275 78.555 ;
        RECT 26.355 77.645 27.275 77.875 ;
        RECT 27.445 77.735 29.375 78.555 ;
        RECT 28.425 77.645 29.375 77.735 ;
        RECT 29.625 77.875 36.935 78.555 ;
        RECT 29.625 77.645 30.975 77.875 ;
        RECT 32.510 77.655 33.420 77.875 ;
        RECT 37.875 77.685 38.305 78.470 ;
        RECT 38.470 77.645 41.535 78.555 ;
        RECT 41.545 77.875 46.360 78.555 ;
        RECT 46.605 77.875 53.915 78.555 ;
        RECT 50.120 77.655 51.030 77.875 ;
        RECT 52.565 77.645 53.915 77.875 ;
        RECT 53.965 77.745 55.335 78.555 ;
        RECT 55.655 77.875 57.490 78.555 ;
        RECT 58.725 78.555 58.875 78.575 ;
        RECT 61.005 78.555 61.175 78.745 ;
        RECT 62.385 78.575 62.555 78.765 ;
        RECT 64.225 78.555 64.395 78.745 ;
        RECT 65.605 78.575 65.775 78.765 ;
        RECT 72.970 78.745 73.135 78.765 ;
        RECT 67.900 78.605 68.020 78.715 ;
        RECT 68.640 78.555 68.810 78.745 ;
        RECT 72.965 78.575 73.135 78.745 ;
        RECT 75.265 78.575 75.435 78.765 ;
        RECT 75.725 78.555 75.895 78.745 ;
        RECT 77.110 78.575 77.280 78.765 ;
        RECT 77.560 78.555 77.730 78.745 ;
        RECT 78.025 78.555 78.195 78.745 ;
        RECT 78.945 78.575 79.115 78.765 ;
        RECT 86.310 78.745 86.475 78.765 ;
        RECT 79.405 78.555 79.575 78.745 ;
        RECT 86.305 78.575 86.475 78.745 ;
        RECT 86.765 78.555 86.935 78.745 ;
        RECT 89.525 78.555 89.695 78.765 ;
        RECT 55.655 77.645 56.585 77.875 ;
        RECT 58.725 77.735 60.655 78.555 ;
        RECT 60.865 77.875 63.605 78.555 ;
        RECT 59.705 77.645 60.655 77.735 ;
        RECT 63.635 77.685 64.065 78.470 ;
        RECT 64.195 77.875 67.660 78.555 ;
        RECT 66.740 77.645 67.660 77.875 ;
        RECT 68.225 77.875 72.125 78.555 ;
        RECT 72.460 77.875 75.925 78.555 ;
        RECT 68.225 77.645 69.155 77.875 ;
        RECT 72.460 77.645 73.380 77.875 ;
        RECT 76.105 77.645 77.875 78.555 ;
        RECT 77.885 77.775 79.255 78.555 ;
        RECT 79.265 77.875 86.575 78.555 ;
        RECT 86.625 77.875 88.455 78.555 ;
        RECT 82.780 77.655 83.690 77.875 ;
        RECT 85.225 77.645 86.575 77.875 ;
        RECT 87.110 77.645 88.455 77.875 ;
        RECT 88.465 77.745 89.835 78.555 ;
      LAYER nwell ;
        RECT 11.910 74.525 90.030 77.355 ;
      LAYER pwell ;
        RECT 99.810 74.755 110.700 80.745 ;
        RECT 12.105 73.325 13.475 74.135 ;
        RECT 17.000 74.005 17.910 74.225 ;
        RECT 19.445 74.005 20.795 74.235 ;
        RECT 13.485 73.325 20.795 74.005 ;
        RECT 21.305 73.325 23.120 74.235 ;
        RECT 23.145 73.325 24.975 74.235 ;
        RECT 24.995 73.410 25.425 74.195 ;
        RECT 25.445 73.325 29.105 74.235 ;
        RECT 29.585 73.325 34.400 74.005 ;
        RECT 34.645 73.325 36.475 74.135 ;
        RECT 39.600 74.005 40.520 74.235 ;
        RECT 43.345 74.035 44.295 74.235 ;
        RECT 37.055 73.325 40.520 74.005 ;
        RECT 40.625 73.355 44.295 74.035 ;
        RECT 12.245 73.115 12.415 73.325 ;
        RECT 13.625 73.135 13.795 73.325 ;
        RECT 17.305 73.115 17.475 73.305 ;
        RECT 19.605 73.135 19.775 73.305 ;
        RECT 20.980 73.165 21.100 73.275 ;
        RECT 19.605 73.115 19.770 73.135 ;
        RECT 21.445 73.115 21.615 73.305 ;
        RECT 21.905 73.135 22.075 73.305 ;
        RECT 22.825 73.135 22.995 73.325 ;
        RECT 21.925 73.115 22.075 73.135 ;
        RECT 24.205 73.115 24.375 73.305 ;
        RECT 24.660 73.135 24.830 73.325 ;
        RECT 27.895 73.160 28.055 73.270 ;
        RECT 12.105 72.305 13.475 73.115 ;
        RECT 14.405 72.435 17.615 73.115 ;
        RECT 17.935 72.435 19.770 73.115 ;
        RECT 14.405 72.205 15.540 72.435 ;
        RECT 17.935 72.205 18.865 72.435 ;
        RECT 19.925 72.205 21.740 73.115 ;
        RECT 21.925 72.295 23.855 73.115 ;
        RECT 22.905 72.205 23.855 72.295 ;
        RECT 24.065 72.205 27.735 73.115 ;
        RECT 28.810 73.085 28.980 73.325 ;
        RECT 29.260 73.165 29.380 73.275 ;
        RECT 29.725 73.135 29.895 73.325 ;
        RECT 32.025 73.135 32.195 73.305 ;
        RECT 34.785 73.135 34.955 73.325 ;
        RECT 36.160 73.165 36.280 73.275 ;
        RECT 32.035 73.115 32.195 73.135 ;
        RECT 36.620 73.115 36.790 73.305 ;
        RECT 37.085 73.135 37.255 73.325 ;
        RECT 39.385 73.115 39.555 73.305 ;
        RECT 40.770 73.135 40.940 73.355 ;
        RECT 43.345 73.325 44.295 73.355 ;
        RECT 44.305 73.325 45.675 74.135 ;
        RECT 45.780 74.005 46.700 74.235 ;
        RECT 45.780 73.325 49.245 74.005 ;
        RECT 49.365 73.325 50.735 74.135 ;
        RECT 50.755 73.410 51.185 74.195 ;
        RECT 51.205 73.325 54.875 74.135 ;
        RECT 56.290 74.005 57.635 74.235 ;
        RECT 55.805 73.325 57.635 74.005 ;
        RECT 57.645 73.325 59.475 74.235 ;
        RECT 62.140 74.005 63.060 74.235 ;
        RECT 59.595 73.325 63.060 74.005 ;
        RECT 63.165 73.325 66.375 74.235 ;
        RECT 69.900 74.005 70.810 74.225 ;
        RECT 72.345 74.005 73.695 74.235 ;
        RECT 66.385 73.325 73.695 74.005 ;
        RECT 74.665 74.005 76.010 74.235 ;
        RECT 74.665 73.325 76.495 74.005 ;
        RECT 76.515 73.410 76.945 74.195 ;
        RECT 77.060 74.005 77.980 74.235 ;
        RECT 82.970 74.005 84.315 74.235 ;
        RECT 77.060 73.325 80.525 74.005 ;
        RECT 80.645 73.325 82.475 74.005 ;
        RECT 82.485 73.325 84.315 74.005 ;
        RECT 84.325 73.325 87.535 74.235 ;
        RECT 88.465 73.325 89.835 74.135 ;
        RECT 44.445 73.135 44.615 73.325 ;
        RECT 46.745 73.115 46.915 73.305 ;
        RECT 49.045 73.135 49.215 73.325 ;
        RECT 49.505 73.135 49.675 73.325 ;
        RECT 49.505 73.115 49.525 73.135 ;
        RECT 50.240 73.115 50.410 73.305 ;
        RECT 51.345 73.135 51.515 73.325 ;
        RECT 55.035 73.170 55.195 73.280 ;
        RECT 55.945 73.135 56.115 73.325 ;
        RECT 57.325 73.115 57.495 73.305 ;
        RECT 57.795 73.160 57.955 73.270 ;
        RECT 58.980 73.115 59.150 73.305 ;
        RECT 59.160 73.135 59.330 73.325 ;
        RECT 59.625 73.135 59.795 73.325 ;
        RECT 62.855 73.160 63.015 73.270 ;
        RECT 63.305 73.135 63.475 73.325 ;
        RECT 64.500 73.115 64.670 73.305 ;
        RECT 66.525 73.135 66.695 73.325 ;
        RECT 68.360 73.165 68.480 73.275 ;
        RECT 69.100 73.115 69.270 73.305 ;
        RECT 73.240 73.115 73.410 73.305 ;
        RECT 73.895 73.170 74.055 73.280 ;
        RECT 76.185 73.135 76.355 73.325 ;
        RECT 80.325 73.115 80.495 73.325 ;
        RECT 82.165 73.135 82.335 73.325 ;
        RECT 82.625 73.305 82.795 73.325 ;
        RECT 82.620 73.135 82.795 73.305 ;
        RECT 82.620 73.115 82.790 73.135 ;
        RECT 83.085 73.115 83.255 73.305 ;
        RECT 84.465 73.115 84.635 73.305 ;
        RECT 87.225 73.135 87.395 73.325 ;
        RECT 87.695 73.160 87.855 73.280 ;
        RECT 89.525 73.115 89.695 73.325 ;
        RECT 30.940 73.085 31.875 73.115 ;
        RECT 28.810 72.885 31.875 73.085 ;
        RECT 28.665 72.405 31.875 72.885 ;
        RECT 28.665 72.205 29.595 72.405 ;
        RECT 30.925 72.205 31.875 72.405 ;
        RECT 32.035 72.205 35.690 73.115 ;
        RECT 36.505 72.205 37.855 73.115 ;
        RECT 37.875 72.245 38.305 73.030 ;
        RECT 38.335 72.205 39.685 73.115 ;
        RECT 39.745 72.435 47.055 73.115 ;
        RECT 47.075 72.435 49.525 73.115 ;
        RECT 49.825 72.435 53.725 73.115 ;
        RECT 54.060 72.435 57.525 73.115 ;
        RECT 58.565 72.435 62.465 73.115 ;
        RECT 39.745 72.205 41.095 72.435 ;
        RECT 42.630 72.215 43.540 72.435 ;
        RECT 47.075 72.205 49.035 72.435 ;
        RECT 49.825 72.205 50.755 72.435 ;
        RECT 54.060 72.205 54.980 72.435 ;
        RECT 58.565 72.205 59.495 72.435 ;
        RECT 63.635 72.245 64.065 73.030 ;
        RECT 64.085 72.435 67.985 73.115 ;
        RECT 68.685 72.435 72.585 73.115 ;
        RECT 72.825 72.435 76.725 73.115 ;
        RECT 77.060 72.435 80.525 73.115 ;
        RECT 64.085 72.205 65.015 72.435 ;
        RECT 68.685 72.205 69.615 72.435 ;
        RECT 72.825 72.205 73.755 72.435 ;
        RECT 77.060 72.205 77.980 72.435 ;
        RECT 80.745 72.205 82.935 73.115 ;
        RECT 82.945 72.335 84.315 73.115 ;
        RECT 84.325 72.205 87.535 73.115 ;
        RECT 88.465 72.305 89.835 73.115 ;
      LAYER nwell ;
        RECT 11.910 69.085 90.030 71.915 ;
      LAYER pwell ;
        RECT 12.105 67.885 13.475 68.695 ;
        RECT 13.960 67.885 15.775 68.795 ;
        RECT 17.155 68.565 18.075 68.795 ;
        RECT 15.785 67.885 18.075 68.565 ;
        RECT 18.085 68.565 19.220 68.795 ;
        RECT 18.085 67.885 21.295 68.565 ;
        RECT 22.225 67.885 24.975 68.795 ;
        RECT 24.995 67.970 25.425 68.755 ;
        RECT 25.445 67.885 27.275 68.695 ;
        RECT 29.360 68.565 30.495 68.795 ;
        RECT 34.020 68.565 34.930 68.785 ;
        RECT 36.465 68.565 37.815 68.795 ;
        RECT 27.285 67.885 30.495 68.565 ;
        RECT 30.505 67.885 37.815 68.565 ;
        RECT 37.875 67.885 40.605 68.795 ;
        RECT 44.140 68.565 45.050 68.785 ;
        RECT 46.585 68.565 47.935 68.795 ;
        RECT 49.035 68.565 49.965 68.795 ;
        RECT 40.625 67.885 47.935 68.565 ;
        RECT 48.130 67.885 49.965 68.565 ;
        RECT 50.755 67.970 51.185 68.755 ;
        RECT 51.215 67.885 52.565 68.795 ;
        RECT 52.585 68.565 53.515 68.795 ;
        RECT 56.765 68.565 58.115 68.795 ;
        RECT 59.650 68.565 60.560 68.785 ;
        RECT 64.545 68.565 65.890 68.795 ;
        RECT 69.900 68.565 70.810 68.785 ;
        RECT 72.345 68.565 73.695 68.795 ;
        RECT 52.585 67.885 56.485 68.565 ;
        RECT 56.765 67.885 64.075 68.565 ;
        RECT 64.545 67.885 66.375 68.565 ;
        RECT 66.385 67.885 73.695 68.565 ;
        RECT 73.745 67.885 75.835 68.695 ;
        RECT 76.515 67.970 76.945 68.755 ;
        RECT 76.965 67.885 81.780 68.565 ;
        RECT 82.025 67.885 85.500 68.795 ;
        RECT 86.755 68.565 87.685 68.795 ;
        RECT 85.850 67.885 87.685 68.565 ;
        RECT 88.465 67.885 89.835 68.695 ;
        RECT 12.245 67.675 12.415 67.885 ;
        RECT 13.620 67.725 13.740 67.835 ;
        RECT 14.085 67.695 14.255 67.885 ;
        RECT 15.925 67.695 16.095 67.885 ;
        RECT 20.525 67.675 20.695 67.865 ;
        RECT 20.985 67.695 21.155 67.885 ;
        RECT 21.455 67.730 21.615 67.840 ;
        RECT 22.365 67.695 22.535 67.885 ;
        RECT 22.825 67.675 22.995 67.865 ;
        RECT 23.285 67.675 23.455 67.865 ;
        RECT 25.120 67.725 25.240 67.835 ;
        RECT 25.585 67.695 25.755 67.885 ;
        RECT 27.425 67.695 27.595 67.885 ;
        RECT 28.345 67.675 28.515 67.865 ;
        RECT 28.810 67.675 28.980 67.865 ;
        RECT 30.185 67.675 30.355 67.865 ;
        RECT 30.645 67.695 30.815 67.885 ;
        RECT 12.105 66.865 13.475 67.675 ;
        RECT 13.525 66.995 20.835 67.675 ;
        RECT 20.845 66.995 23.135 67.675 ;
        RECT 23.145 66.995 24.975 67.675 ;
        RECT 13.525 66.765 14.875 66.995 ;
        RECT 16.410 66.775 17.320 66.995 ;
        RECT 20.845 66.765 21.765 66.995 ;
        RECT 25.445 66.765 28.655 67.675 ;
        RECT 28.665 66.765 30.015 67.675 ;
        RECT 30.045 66.865 31.415 67.675 ;
        RECT 31.425 67.645 32.360 67.675 ;
        RECT 34.320 67.645 34.490 67.865 ;
        RECT 34.785 67.675 34.955 67.865 ;
        RECT 37.540 67.725 37.660 67.835 ;
        RECT 38.005 67.695 38.175 67.885 ;
        RECT 38.465 67.675 38.635 67.865 ;
        RECT 39.845 67.675 40.015 67.865 ;
        RECT 40.765 67.695 40.935 67.885 ;
        RECT 48.130 67.865 48.295 67.885 ;
        RECT 41.225 67.675 41.395 67.865 ;
        RECT 43.525 67.675 43.695 67.865 ;
        RECT 45.360 67.725 45.480 67.835 ;
        RECT 45.825 67.675 45.995 67.865 ;
        RECT 48.125 67.695 48.295 67.865 ;
        RECT 50.420 67.725 50.540 67.835 ;
        RECT 52.265 67.695 52.435 67.885 ;
        RECT 53.000 67.695 53.170 67.885 ;
        RECT 53.190 67.675 53.360 67.865 ;
        RECT 63.305 67.675 63.475 67.865 ;
        RECT 63.765 67.695 63.935 67.885 ;
        RECT 64.225 67.835 64.395 67.865 ;
        RECT 64.220 67.725 64.395 67.835 ;
        RECT 64.225 67.675 64.395 67.725 ;
        RECT 66.065 67.695 66.235 67.885 ;
        RECT 66.525 67.695 66.695 67.885 ;
        RECT 66.985 67.675 67.155 67.865 ;
        RECT 73.885 67.695 74.055 67.885 ;
        RECT 75.725 67.675 75.895 67.865 ;
        RECT 76.185 67.695 76.355 67.865 ;
        RECT 77.105 67.695 77.275 67.885 ;
        RECT 78.485 67.695 78.655 67.865 ;
        RECT 80.780 67.725 80.900 67.835 ;
        RECT 76.205 67.675 76.355 67.695 ;
        RECT 78.490 67.675 78.655 67.695 ;
        RECT 81.245 67.675 81.415 67.865 ;
        RECT 82.170 67.695 82.340 67.885 ;
        RECT 85.850 67.865 86.015 67.885 ;
        RECT 85.845 67.695 86.015 67.865 ;
        RECT 88.140 67.725 88.260 67.835 ;
        RECT 89.525 67.675 89.695 67.885 ;
        RECT 31.425 67.445 34.490 67.645 ;
        RECT 31.425 66.965 34.635 67.445 ;
        RECT 31.425 66.765 32.375 66.965 ;
        RECT 33.705 66.765 34.635 66.965 ;
        RECT 34.655 66.765 37.385 67.675 ;
        RECT 37.875 66.805 38.305 67.590 ;
        RECT 38.325 66.865 39.695 67.675 ;
        RECT 39.705 66.895 41.075 67.675 ;
        RECT 41.085 66.995 43.375 67.675 ;
        RECT 42.455 66.765 43.375 66.995 ;
        RECT 43.385 66.865 45.215 67.675 ;
        RECT 45.685 66.995 52.995 67.675 ;
        RECT 49.200 66.775 50.110 66.995 ;
        RECT 51.645 66.765 52.995 66.995 ;
        RECT 53.045 66.765 56.160 67.675 ;
        RECT 56.305 66.995 63.615 67.675 ;
        RECT 56.305 66.765 57.655 66.995 ;
        RECT 59.190 66.775 60.100 66.995 ;
        RECT 63.635 66.805 64.065 67.590 ;
        RECT 64.085 66.865 66.835 67.675 ;
        RECT 66.845 66.995 74.155 67.675 ;
        RECT 70.360 66.775 71.270 66.995 ;
        RECT 72.805 66.765 74.155 66.995 ;
        RECT 74.205 66.995 76.035 67.675 ;
        RECT 74.205 66.765 75.550 66.995 ;
        RECT 76.205 66.855 78.135 67.675 ;
        RECT 78.490 66.995 80.325 67.675 ;
        RECT 81.105 66.995 88.415 67.675 ;
        RECT 77.185 66.765 78.135 66.855 ;
        RECT 79.395 66.765 80.325 66.995 ;
        RECT 84.620 66.775 85.530 66.995 ;
        RECT 87.065 66.765 88.415 66.995 ;
        RECT 88.465 66.865 89.835 67.675 ;
      LAYER nwell ;
        RECT 11.910 63.645 90.030 66.475 ;
      LAYER pwell ;
        RECT 12.105 62.445 13.475 63.255 ;
        RECT 17.000 63.125 17.910 63.345 ;
        RECT 19.445 63.125 20.795 63.355 ;
        RECT 13.485 62.445 20.795 63.125 ;
        RECT 20.845 62.445 22.195 63.355 ;
        RECT 22.225 62.445 24.975 63.255 ;
        RECT 24.995 62.530 25.425 63.315 ;
        RECT 25.445 62.445 28.195 63.255 ;
        RECT 28.205 62.445 29.555 63.355 ;
        RECT 29.605 62.445 30.955 63.355 ;
        RECT 30.965 62.445 32.795 63.255 ;
        RECT 32.805 63.125 33.725 63.355 ;
        RECT 32.805 62.445 35.095 63.125 ;
        RECT 35.105 62.445 40.615 63.255 ;
        RECT 40.625 62.445 46.135 63.255 ;
        RECT 46.145 62.445 47.975 63.255 ;
        RECT 49.815 63.125 50.735 63.355 ;
        RECT 48.445 62.445 50.735 63.125 ;
        RECT 50.755 62.530 51.185 63.315 ;
        RECT 52.575 63.155 53.930 63.355 ;
        RECT 51.250 63.125 53.930 63.155 ;
        RECT 55.795 63.125 56.715 63.355 ;
        RECT 51.250 62.475 54.415 63.125 ;
        RECT 52.575 62.445 54.415 62.475 ;
        RECT 54.425 62.445 56.715 63.125 ;
        RECT 56.725 62.445 62.235 63.255 ;
        RECT 62.245 62.445 64.995 63.255 ;
        RECT 65.005 62.445 69.820 63.125 ;
        RECT 70.065 62.445 71.895 63.255 ;
        RECT 72.005 62.445 74.195 63.355 ;
        RECT 74.405 63.265 75.355 63.355 ;
        RECT 74.405 62.445 76.335 63.265 ;
        RECT 76.515 62.530 76.945 63.315 ;
        RECT 77.620 62.445 81.095 63.355 ;
        RECT 84.620 63.125 85.530 63.345 ;
        RECT 87.065 63.125 88.415 63.355 ;
        RECT 81.105 62.445 88.415 63.125 ;
        RECT 88.465 62.445 89.835 63.255 ;
        RECT 12.245 62.235 12.415 62.445 ;
        RECT 13.625 62.235 13.795 62.445 ;
        RECT 16.845 62.235 17.015 62.425 ;
        RECT 17.305 62.235 17.475 62.425 ;
        RECT 20.060 62.235 20.230 62.425 ;
        RECT 20.525 62.235 20.695 62.425 ;
        RECT 20.990 62.255 21.160 62.445 ;
        RECT 22.365 62.255 22.535 62.445 ;
        RECT 25.585 62.255 25.755 62.445 ;
        RECT 26.040 62.285 26.160 62.395 ;
        RECT 26.510 62.235 26.680 62.425 ;
        RECT 29.270 62.255 29.440 62.445 ;
        RECT 29.720 62.255 29.890 62.445 ;
        RECT 31.105 62.255 31.275 62.445 ;
        RECT 34.325 62.255 34.495 62.425 ;
        RECT 34.785 62.255 34.955 62.445 ;
        RECT 35.245 62.255 35.415 62.445 ;
        RECT 34.330 62.235 34.495 62.255 ;
        RECT 36.625 62.235 36.795 62.425 ;
        RECT 38.465 62.235 38.635 62.425 ;
        RECT 40.765 62.255 40.935 62.445 ;
        RECT 42.145 62.235 42.315 62.425 ;
        RECT 44.905 62.235 45.075 62.425 ;
        RECT 45.365 62.235 45.535 62.425 ;
        RECT 46.285 62.255 46.455 62.445 ;
        RECT 48.120 62.285 48.240 62.395 ;
        RECT 48.585 62.255 48.755 62.445 ;
        RECT 49.040 62.235 49.210 62.425 ;
        RECT 49.505 62.235 49.675 62.425 ;
        RECT 53.185 62.255 53.355 62.425 ;
        RECT 54.105 62.255 54.275 62.445 ;
        RECT 54.565 62.255 54.735 62.445 ;
        RECT 53.185 62.235 53.350 62.255 ;
        RECT 55.020 62.235 55.190 62.425 ;
        RECT 55.485 62.235 55.655 62.425 ;
        RECT 56.865 62.255 57.035 62.445 ;
        RECT 61.005 62.235 61.175 62.425 ;
        RECT 62.385 62.255 62.555 62.445 ;
        RECT 64.235 62.280 64.395 62.390 ;
        RECT 65.145 62.235 65.315 62.445 ;
        RECT 68.365 62.235 68.535 62.425 ;
        RECT 70.205 62.255 70.375 62.445 ;
        RECT 73.880 62.425 74.050 62.445 ;
        RECT 76.185 62.425 76.335 62.445 ;
        RECT 72.040 62.285 72.160 62.395 ;
        RECT 73.880 62.255 74.055 62.425 ;
        RECT 73.885 62.235 74.055 62.255 ;
        RECT 75.725 62.235 75.895 62.425 ;
        RECT 76.185 62.255 76.355 62.425 ;
        RECT 77.095 62.235 77.265 62.425 ;
        RECT 80.780 62.235 80.950 62.445 ;
        RECT 81.245 62.235 81.415 62.445 ;
        RECT 89.525 62.235 89.695 62.445 ;
        RECT 12.105 61.425 13.475 62.235 ;
        RECT 13.485 61.425 14.855 62.235 ;
        RECT 14.865 61.555 17.155 62.235 ;
        RECT 17.165 61.555 18.995 62.235 ;
        RECT 14.865 61.325 15.785 61.555 ;
        RECT 19.025 61.325 20.375 62.235 ;
        RECT 20.385 61.425 25.895 62.235 ;
        RECT 26.365 61.325 34.115 62.235 ;
        RECT 34.330 61.555 36.165 62.235 ;
        RECT 35.235 61.325 36.165 61.555 ;
        RECT 36.485 61.425 37.855 62.235 ;
        RECT 37.875 61.365 38.305 62.150 ;
        RECT 38.325 61.425 41.995 62.235 ;
        RECT 42.005 61.425 43.375 62.235 ;
        RECT 43.385 61.325 45.200 62.235 ;
        RECT 45.225 61.425 47.975 62.235 ;
        RECT 48.005 61.325 49.355 62.235 ;
        RECT 49.365 61.425 51.195 62.235 ;
        RECT 51.515 61.555 53.350 62.235 ;
        RECT 51.515 61.325 52.445 61.555 ;
        RECT 53.505 61.325 55.335 62.235 ;
        RECT 55.345 61.425 60.855 62.235 ;
        RECT 60.865 61.425 63.615 62.235 ;
        RECT 63.635 61.365 64.065 62.150 ;
        RECT 65.055 61.325 68.215 62.235 ;
        RECT 68.225 61.425 71.895 62.235 ;
        RECT 72.365 61.555 74.195 62.235 ;
        RECT 74.205 61.555 76.035 62.235 ;
        RECT 72.365 61.325 73.710 61.555 ;
        RECT 74.205 61.325 75.550 61.555 ;
        RECT 76.045 61.455 77.415 62.235 ;
        RECT 77.620 61.325 81.095 62.235 ;
        RECT 81.105 61.555 88.415 62.235 ;
        RECT 84.620 61.335 85.530 61.555 ;
        RECT 87.065 61.325 88.415 61.555 ;
        RECT 88.465 61.425 89.835 62.235 ;
      LAYER nwell ;
        RECT 11.910 58.205 90.030 61.035 ;
      LAYER pwell ;
        RECT 12.105 57.005 13.475 57.815 ;
        RECT 13.485 57.005 18.995 57.815 ;
        RECT 19.005 57.005 21.755 57.815 ;
        RECT 22.235 57.005 24.965 57.915 ;
        RECT 24.995 57.090 25.425 57.875 ;
        RECT 32.845 57.685 34.195 57.915 ;
        RECT 35.730 57.685 36.640 57.905 ;
        RECT 40.165 57.715 41.095 57.915 ;
        RECT 42.425 57.715 43.375 57.915 ;
        RECT 25.905 57.005 27.735 57.685 ;
        RECT 27.980 57.005 32.795 57.685 ;
        RECT 32.845 57.005 40.155 57.685 ;
        RECT 40.165 57.235 43.375 57.715 ;
        RECT 46.040 57.685 46.960 57.915 ;
        RECT 40.310 57.035 43.375 57.235 ;
        RECT 12.245 56.795 12.415 57.005 ;
        RECT 13.625 56.795 13.795 57.005 ;
        RECT 19.145 56.795 19.315 57.005 ;
        RECT 20.530 56.795 20.700 56.985 ;
        RECT 21.900 56.845 22.020 56.955 ;
        RECT 22.365 56.795 22.535 57.005 ;
        RECT 25.585 56.955 25.755 56.985 ;
        RECT 25.580 56.845 25.755 56.955 ;
        RECT 25.585 56.795 25.755 56.845 ;
        RECT 26.045 56.815 26.215 57.005 ;
        RECT 29.275 56.840 29.435 56.950 ;
        RECT 32.485 56.815 32.655 57.005 ;
        RECT 33.865 56.815 34.035 56.985 ;
        RECT 33.865 56.795 34.010 56.815 ;
        RECT 36.625 56.795 36.795 56.985 ;
        RECT 37.095 56.840 37.255 56.950 ;
        RECT 39.845 56.815 40.015 57.005 ;
        RECT 40.310 56.985 40.480 57.035 ;
        RECT 42.440 57.005 43.375 57.035 ;
        RECT 43.495 57.005 46.960 57.685 ;
        RECT 47.080 57.005 48.895 57.915 ;
        RECT 49.385 57.005 50.735 57.915 ;
        RECT 50.755 57.090 51.185 57.875 ;
        RECT 51.300 57.685 52.220 57.915 ;
        RECT 55.900 57.685 56.820 57.915 ;
        RECT 51.300 57.005 54.765 57.685 ;
        RECT 55.900 57.005 59.365 57.685 ;
        RECT 59.485 57.005 62.235 57.815 ;
        RECT 65.760 57.685 66.670 57.905 ;
        RECT 68.205 57.685 69.555 57.915 ;
        RECT 62.245 57.005 69.555 57.685 ;
        RECT 69.605 57.005 70.975 57.815 ;
        RECT 70.985 57.685 72.330 57.915 ;
        RECT 70.985 57.005 72.815 57.685 ;
        RECT 72.825 57.005 76.300 57.915 ;
        RECT 76.515 57.090 76.945 57.875 ;
        RECT 80.480 57.685 81.390 57.905 ;
        RECT 82.925 57.685 84.275 57.915 ;
        RECT 76.965 57.005 84.275 57.685 ;
        RECT 84.635 57.685 85.565 57.915 ;
        RECT 87.110 57.685 88.455 57.915 ;
        RECT 84.635 57.005 86.470 57.685 ;
        RECT 86.625 57.005 88.455 57.685 ;
        RECT 88.465 57.005 89.835 57.815 ;
        RECT 40.305 56.815 40.480 56.985 ;
        RECT 40.760 56.845 40.880 56.955 ;
        RECT 43.525 56.815 43.695 57.005 ;
        RECT 47.205 56.815 47.375 57.005 ;
        RECT 40.305 56.795 40.475 56.815 ;
        RECT 48.125 56.795 48.295 56.985 ;
        RECT 48.585 56.795 48.755 56.985 ;
        RECT 49.040 56.845 49.160 56.955 ;
        RECT 50.420 56.815 50.590 57.005 ;
        RECT 52.265 56.795 52.435 56.985 ;
        RECT 54.565 56.815 54.735 57.005 ;
        RECT 55.035 56.955 55.195 56.960 ;
        RECT 55.020 56.850 55.195 56.955 ;
        RECT 55.020 56.845 55.140 56.850 ;
        RECT 55.485 56.795 55.655 56.985 ;
        RECT 59.165 56.815 59.335 57.005 ;
        RECT 59.625 56.815 59.795 57.005 ;
        RECT 62.385 56.815 62.555 57.005 ;
        RECT 63.300 56.845 63.420 56.955 ;
        RECT 64.225 56.795 64.395 56.985 ;
        RECT 69.745 56.815 69.915 57.005 ;
        RECT 72.045 56.795 72.215 56.985 ;
        RECT 72.505 56.815 72.675 57.005 ;
        RECT 72.970 56.815 73.140 57.005 ;
        RECT 77.105 56.815 77.275 57.005 ;
        RECT 86.305 56.985 86.470 57.005 ;
        RECT 82.165 56.795 82.335 56.985 ;
        RECT 82.635 56.840 82.795 56.950 ;
        RECT 83.545 56.815 83.715 56.985 ;
        RECT 85.845 56.815 86.015 56.985 ;
        RECT 86.305 56.815 86.475 56.985 ;
        RECT 86.765 56.815 86.935 57.005 ;
        RECT 88.140 56.845 88.260 56.955 ;
        RECT 83.550 56.795 83.715 56.815 ;
        RECT 85.850 56.795 86.015 56.815 ;
        RECT 89.525 56.795 89.695 57.005 ;
        RECT 12.105 55.985 13.475 56.795 ;
        RECT 13.485 55.985 18.995 56.795 ;
        RECT 19.005 55.985 20.375 56.795 ;
        RECT 20.385 55.885 22.215 56.795 ;
        RECT 22.325 55.885 25.435 56.795 ;
        RECT 25.445 56.115 29.115 56.795 ;
        RECT 28.185 55.885 29.115 56.115 ;
        RECT 30.140 55.885 34.010 56.795 ;
        RECT 34.185 56.115 36.935 56.795 ;
        RECT 34.185 55.885 35.115 56.115 ;
        RECT 37.875 55.925 38.305 56.710 ;
        RECT 38.325 56.115 40.615 56.795 ;
        RECT 41.125 56.115 48.435 56.795 ;
        RECT 48.555 56.115 52.020 56.795 ;
        RECT 38.325 55.885 39.245 56.115 ;
        RECT 41.125 55.885 42.475 56.115 ;
        RECT 44.010 55.895 44.920 56.115 ;
        RECT 51.100 55.885 52.020 56.115 ;
        RECT 52.125 55.885 54.875 56.795 ;
        RECT 55.345 56.115 63.075 56.795 ;
        RECT 58.860 55.895 59.770 56.115 ;
        RECT 61.305 55.885 63.075 56.115 ;
        RECT 63.635 55.925 64.065 56.710 ;
        RECT 64.085 56.115 71.815 56.795 ;
        RECT 71.905 56.115 79.215 56.795 ;
        RECT 67.600 55.895 68.510 56.115 ;
        RECT 70.045 55.885 71.815 56.115 ;
        RECT 75.420 55.895 76.330 56.115 ;
        RECT 77.865 55.885 79.215 56.115 ;
        RECT 79.265 55.885 82.475 56.795 ;
        RECT 83.550 56.115 85.385 56.795 ;
        RECT 85.850 56.115 87.685 56.795 ;
        RECT 84.455 55.885 85.385 56.115 ;
        RECT 86.755 55.885 87.685 56.115 ;
        RECT 88.465 55.985 89.835 56.795 ;
      LAYER nwell ;
        RECT 11.910 52.765 90.030 55.595 ;
      LAYER pwell ;
        RECT 12.105 51.565 13.475 52.375 ;
        RECT 13.485 51.565 15.315 52.375 ;
        RECT 15.325 52.245 16.245 52.475 ;
        RECT 15.325 51.565 17.615 52.245 ;
        RECT 17.625 51.565 19.440 52.475 ;
        RECT 19.465 51.565 22.215 52.375 ;
        RECT 23.735 52.245 24.665 52.475 ;
        RECT 22.830 51.565 24.665 52.245 ;
        RECT 24.995 51.650 25.425 52.435 ;
        RECT 27.250 52.275 28.195 52.475 ;
        RECT 25.445 51.595 28.195 52.275 ;
        RECT 12.245 51.355 12.415 51.565 ;
        RECT 13.625 51.375 13.795 51.565 ;
        RECT 17.305 51.375 17.475 51.565 ;
        RECT 19.145 51.375 19.315 51.565 ;
        RECT 19.605 51.375 19.775 51.565 ;
        RECT 22.830 51.545 22.995 51.565 ;
        RECT 20.525 51.355 20.695 51.545 ;
        RECT 20.985 51.355 21.155 51.545 ;
        RECT 22.360 51.405 22.480 51.515 ;
        RECT 22.825 51.375 22.995 51.545 ;
        RECT 23.290 51.355 23.460 51.545 ;
        RECT 24.665 51.355 24.835 51.545 ;
        RECT 25.590 51.375 25.760 51.595 ;
        RECT 27.250 51.565 28.195 51.595 ;
        RECT 29.125 51.565 32.335 52.475 ;
        RECT 44.600 52.245 45.510 52.465 ;
        RECT 47.045 52.245 48.395 52.475 ;
        RECT 49.815 52.245 50.735 52.475 ;
        RECT 33.210 51.565 35.635 52.245 ;
        RECT 36.260 51.565 41.075 52.245 ;
        RECT 41.085 51.565 48.395 52.245 ;
        RECT 48.445 51.565 50.735 52.245 ;
        RECT 50.755 51.650 51.185 52.435 ;
        RECT 54.720 52.245 55.630 52.465 ;
        RECT 57.165 52.245 58.515 52.475 ;
        RECT 63.625 52.245 64.555 52.475 ;
        RECT 75.080 52.275 76.035 52.475 ;
        RECT 51.205 51.565 58.515 52.245 ;
        RECT 58.800 51.565 63.615 52.245 ;
        RECT 63.625 51.565 67.525 52.245 ;
        RECT 68.920 51.565 73.735 52.245 ;
        RECT 73.755 51.595 76.035 52.275 ;
        RECT 76.515 51.650 76.945 52.435 ;
        RECT 77.275 52.245 78.205 52.475 ;
        RECT 28.355 51.410 28.515 51.520 ;
        RECT 29.265 51.375 29.435 51.565 ;
        RECT 30.185 51.375 30.355 51.545 ;
        RECT 30.185 51.355 30.350 51.375 ;
        RECT 30.645 51.355 30.815 51.545 ;
        RECT 32.480 51.405 32.600 51.515 ;
        RECT 32.945 51.355 33.115 51.545 ;
        RECT 36.165 51.355 36.335 51.545 ;
        RECT 40.305 51.375 40.475 51.545 ;
        RECT 40.765 51.515 40.935 51.565 ;
        RECT 40.760 51.405 40.935 51.515 ;
        RECT 40.765 51.375 40.935 51.405 ;
        RECT 40.305 51.355 40.455 51.375 ;
        RECT 41.225 51.355 41.395 51.565 ;
        RECT 48.585 51.355 48.755 51.565 ;
        RECT 51.345 51.375 51.515 51.565 ;
        RECT 55.945 51.355 56.115 51.545 ;
        RECT 58.980 51.355 59.150 51.545 ;
        RECT 62.855 51.400 63.015 51.510 ;
        RECT 63.305 51.375 63.475 51.565 ;
        RECT 64.040 51.375 64.210 51.565 ;
        RECT 73.425 51.545 73.595 51.565 ;
        RECT 64.235 51.400 64.395 51.510 ;
        RECT 65.420 51.355 65.590 51.545 ;
        RECT 67.915 51.410 68.075 51.520 ;
        RECT 69.560 51.355 69.730 51.545 ;
        RECT 73.425 51.375 73.600 51.545 ;
        RECT 73.880 51.375 74.050 51.595 ;
        RECT 75.080 51.565 76.035 51.595 ;
        RECT 77.275 51.565 79.110 52.245 ;
        RECT 79.265 51.565 80.635 52.375 ;
        RECT 80.645 51.565 84.120 52.475 ;
        RECT 84.635 52.245 85.565 52.475 ;
        RECT 87.110 52.245 88.455 52.475 ;
        RECT 84.635 51.565 86.470 52.245 ;
        RECT 86.625 51.565 88.455 52.245 ;
        RECT 88.465 51.565 89.835 52.375 ;
        RECT 78.945 51.545 79.110 51.565 ;
        RECT 76.180 51.405 76.300 51.515 ;
        RECT 77.100 51.405 77.220 51.515 ;
        RECT 78.945 51.375 79.115 51.545 ;
        RECT 79.405 51.375 79.575 51.565 ;
        RECT 80.790 51.545 80.960 51.565 ;
        RECT 86.305 51.545 86.470 51.565 ;
        RECT 80.780 51.375 80.960 51.545 ;
        RECT 73.430 51.355 73.600 51.375 ;
        RECT 80.780 51.355 80.950 51.375 ;
        RECT 81.245 51.355 81.415 51.545 ;
        RECT 86.305 51.375 86.475 51.545 ;
        RECT 86.765 51.375 86.935 51.565 ;
        RECT 89.525 51.355 89.695 51.565 ;
        RECT 12.105 50.545 13.475 51.355 ;
        RECT 13.525 50.675 20.835 51.355 ;
        RECT 20.845 50.675 23.135 51.355 ;
        RECT 13.525 50.445 14.875 50.675 ;
        RECT 16.410 50.455 17.320 50.675 ;
        RECT 22.215 50.445 23.135 50.675 ;
        RECT 23.145 50.445 24.495 51.355 ;
        RECT 24.525 50.545 28.195 51.355 ;
        RECT 28.515 50.675 30.350 51.355 ;
        RECT 30.505 50.675 32.795 51.355 ;
        RECT 28.515 50.445 29.445 50.675 ;
        RECT 31.875 50.445 32.795 50.675 ;
        RECT 32.885 50.445 35.885 51.355 ;
        RECT 36.025 50.545 37.855 51.355 ;
        RECT 37.875 50.485 38.305 51.270 ;
        RECT 38.525 50.535 40.455 51.355 ;
        RECT 41.085 50.675 48.395 51.355 ;
        RECT 48.445 50.675 55.755 51.355 ;
        RECT 38.525 50.445 39.475 50.535 ;
        RECT 44.600 50.455 45.510 50.675 ;
        RECT 47.045 50.445 48.395 50.675 ;
        RECT 51.960 50.455 52.870 50.675 ;
        RECT 54.405 50.445 55.755 50.675 ;
        RECT 55.805 50.545 57.895 51.355 ;
        RECT 58.565 50.675 62.465 51.355 ;
        RECT 58.565 50.445 59.495 50.675 ;
        RECT 63.635 50.485 64.065 51.270 ;
        RECT 65.005 50.675 68.905 51.355 ;
        RECT 69.145 50.675 73.045 51.355 ;
        RECT 65.005 50.445 65.935 50.675 ;
        RECT 69.145 50.445 70.075 50.675 ;
        RECT 73.285 50.445 76.760 51.355 ;
        RECT 77.620 50.445 81.095 51.355 ;
        RECT 81.105 50.675 88.415 51.355 ;
        RECT 84.620 50.455 85.530 50.675 ;
        RECT 87.065 50.445 88.415 50.675 ;
        RECT 88.465 50.545 89.835 51.355 ;
      LAYER nwell ;
        RECT 11.910 47.325 90.030 50.155 ;
      LAYER pwell ;
        RECT 12.105 46.125 13.475 46.935 ;
        RECT 17.920 46.805 18.830 47.025 ;
        RECT 20.365 46.805 21.715 47.035 ;
        RECT 14.405 46.125 21.715 46.805 ;
        RECT 21.765 46.805 22.900 47.035 ;
        RECT 21.765 46.125 24.975 46.805 ;
        RECT 24.995 46.210 25.425 46.995 ;
        RECT 25.445 46.125 27.260 47.035 ;
        RECT 27.285 46.125 28.635 47.035 ;
        RECT 28.665 46.125 32.335 46.935 ;
        RECT 32.345 46.835 33.295 47.035 ;
        RECT 34.625 46.835 35.555 47.035 ;
        RECT 32.345 46.355 35.555 46.835 ;
        RECT 35.565 46.805 36.700 47.035 ;
        RECT 32.345 46.155 35.410 46.355 ;
        RECT 32.345 46.125 33.280 46.155 ;
        RECT 12.245 45.915 12.415 46.125 ;
        RECT 14.545 46.105 14.715 46.125 ;
        RECT 13.635 45.970 13.795 46.080 ;
        RECT 14.540 45.935 14.715 46.105 ;
        RECT 14.540 45.915 14.710 45.935 ;
        RECT 15.005 45.915 15.175 46.105 ;
        RECT 24.205 45.915 24.375 46.105 ;
        RECT 24.665 46.075 24.835 46.125 ;
        RECT 24.660 45.965 24.835 46.075 ;
        RECT 24.665 45.935 24.835 45.965 ;
        RECT 26.965 45.935 27.135 46.125 ;
        RECT 27.430 45.935 27.600 46.125 ;
        RECT 28.805 46.105 28.975 46.125 ;
        RECT 28.340 45.915 28.510 46.105 ;
        RECT 28.805 45.935 28.980 46.105 ;
        RECT 28.810 45.915 28.980 45.935 ;
        RECT 30.645 45.915 30.815 46.105 ;
        RECT 35.240 45.935 35.410 46.155 ;
        RECT 35.565 46.125 38.775 46.805 ;
        RECT 38.785 46.125 41.705 47.035 ;
        RECT 42.315 46.805 43.245 47.035 ;
        RECT 42.315 46.125 44.150 46.805 ;
        RECT 44.305 46.125 45.675 46.935 ;
        RECT 45.705 46.125 47.055 47.035 ;
        RECT 47.160 46.805 48.080 47.035 ;
        RECT 47.160 46.125 50.625 46.805 ;
        RECT 50.755 46.210 51.185 46.995 ;
        RECT 51.205 46.835 52.160 47.035 ;
        RECT 51.205 46.155 53.485 46.835 ;
        RECT 54.005 46.805 55.355 47.035 ;
        RECT 56.890 46.805 57.800 47.025 ;
        RECT 62.665 46.835 64.045 47.035 ;
        RECT 51.205 46.125 52.160 46.155 ;
        RECT 38.465 45.915 38.635 46.125 ;
        RECT 38.930 45.935 39.100 46.125 ;
        RECT 43.985 46.105 44.150 46.125 ;
        RECT 43.985 45.935 44.155 46.105 ;
        RECT 44.445 45.935 44.615 46.125 ;
        RECT 45.820 46.105 45.990 46.125 ;
        RECT 45.820 45.935 46.000 46.105 ;
        RECT 45.830 45.915 46.000 45.935 ;
        RECT 47.665 45.915 47.835 46.105 ;
        RECT 50.425 45.935 50.595 46.125 ;
        RECT 50.895 45.960 51.055 46.070 ;
        RECT 51.805 45.915 51.975 46.105 ;
        RECT 53.190 45.935 53.360 46.155 ;
        RECT 54.005 46.125 61.315 46.805 ;
        RECT 61.340 46.155 64.045 46.835 ;
        RECT 67.600 46.805 68.510 47.025 ;
        RECT 70.045 46.805 71.815 47.035 ;
        RECT 53.640 45.965 53.760 46.075 ;
        RECT 61.005 45.935 61.175 46.125 ;
        RECT 61.465 45.935 61.635 46.155 ;
        RECT 62.665 46.125 64.045 46.155 ;
        RECT 64.085 46.125 71.815 46.805 ;
        RECT 71.905 46.835 72.850 47.035 ;
        RECT 74.185 46.835 75.115 47.035 ;
        RECT 71.905 46.355 75.115 46.835 ;
        RECT 71.905 46.155 74.975 46.355 ;
        RECT 71.905 46.125 72.850 46.155 ;
        RECT 62.385 45.915 62.555 46.105 ;
        RECT 62.855 45.960 63.015 46.070 ;
        RECT 64.225 45.915 64.395 46.125 ;
        RECT 72.045 45.915 72.215 46.105 ;
        RECT 74.805 45.935 74.975 46.155 ;
        RECT 75.125 46.125 76.495 46.935 ;
        RECT 76.515 46.210 76.945 46.995 ;
        RECT 77.160 46.125 80.635 47.035 ;
        RECT 84.620 46.805 85.530 47.025 ;
        RECT 87.065 46.805 88.415 47.035 ;
        RECT 81.105 46.125 88.415 46.805 ;
        RECT 88.465 46.125 89.835 46.935 ;
        RECT 75.265 45.935 75.435 46.125 ;
        RECT 80.320 45.935 80.490 46.125 ;
        RECT 80.780 45.965 80.900 46.075 ;
        RECT 81.245 45.935 81.415 46.125 ;
        RECT 86.305 45.915 86.475 46.105 ;
        RECT 86.765 45.915 86.935 46.105 ;
        RECT 89.525 45.915 89.695 46.125 ;
        RECT 12.105 45.105 13.475 45.915 ;
        RECT 13.505 45.005 14.855 45.915 ;
        RECT 14.865 45.235 22.175 45.915 ;
        RECT 18.380 45.015 19.290 45.235 ;
        RECT 20.825 45.005 22.175 45.235 ;
        RECT 22.225 45.235 24.515 45.915 ;
        RECT 22.225 45.005 23.145 45.235 ;
        RECT 25.180 45.005 28.655 45.915 ;
        RECT 28.665 45.005 30.495 45.915 ;
        RECT 30.505 45.235 37.815 45.915 ;
        RECT 34.020 45.015 34.930 45.235 ;
        RECT 36.465 45.005 37.815 45.235 ;
        RECT 37.875 45.045 38.305 45.830 ;
        RECT 38.325 45.235 45.635 45.915 ;
        RECT 41.840 45.015 42.750 45.235 ;
        RECT 44.285 45.005 45.635 45.235 ;
        RECT 45.685 45.005 47.515 45.915 ;
        RECT 47.625 45.005 50.735 45.915 ;
        RECT 51.665 45.235 58.975 45.915 ;
        RECT 55.180 45.015 56.090 45.235 ;
        RECT 57.625 45.005 58.975 45.235 ;
        RECT 59.120 45.235 62.585 45.915 ;
        RECT 59.120 45.005 60.040 45.235 ;
        RECT 63.635 45.045 64.065 45.830 ;
        RECT 64.085 45.235 71.815 45.915 ;
        RECT 71.905 45.235 79.215 45.915 ;
        RECT 67.600 45.015 68.510 45.235 ;
        RECT 70.045 45.005 71.815 45.235 ;
        RECT 75.420 45.015 76.330 45.235 ;
        RECT 77.865 45.005 79.215 45.235 ;
        RECT 79.305 45.235 86.615 45.915 ;
        RECT 86.625 45.235 88.455 45.915 ;
        RECT 79.305 45.005 80.655 45.235 ;
        RECT 82.190 45.015 83.100 45.235 ;
        RECT 87.110 45.005 88.455 45.235 ;
        RECT 88.465 45.105 89.835 45.915 ;
      LAYER nwell ;
        RECT 11.910 41.885 90.030 44.715 ;
      LAYER pwell ;
        RECT 12.105 40.685 13.475 41.495 ;
        RECT 13.985 40.685 17.155 41.595 ;
        RECT 18.535 41.365 19.455 41.595 ;
        RECT 21.755 41.365 22.675 41.595 ;
        RECT 24.055 41.365 24.975 41.595 ;
        RECT 17.165 40.685 19.455 41.365 ;
        RECT 20.385 40.685 22.675 41.365 ;
        RECT 22.685 40.685 24.975 41.365 ;
        RECT 24.995 40.770 25.425 41.555 ;
        RECT 28.960 41.365 29.870 41.585 ;
        RECT 31.405 41.365 32.755 41.595 ;
        RECT 25.445 40.685 32.755 41.365 ;
        RECT 32.805 40.685 34.155 41.595 ;
        RECT 37.700 41.365 38.610 41.585 ;
        RECT 40.145 41.365 41.495 41.595 ;
        RECT 34.185 40.685 41.495 41.365 ;
        RECT 41.545 41.365 42.465 41.595 ;
        RECT 41.545 40.685 43.835 41.365 ;
        RECT 43.845 40.685 45.675 41.495 ;
        RECT 45.685 40.685 47.035 41.595 ;
        RECT 47.065 40.685 50.735 41.495 ;
        RECT 50.755 40.770 51.185 41.555 ;
        RECT 51.205 40.685 52.575 41.495 ;
        RECT 52.680 41.365 53.600 41.595 ;
        RECT 56.360 41.365 57.280 41.595 ;
        RECT 62.685 41.365 63.615 41.595 ;
        RECT 52.680 40.685 56.145 41.365 ;
        RECT 56.360 40.685 59.825 41.365 ;
        RECT 59.945 40.685 63.615 41.365 ;
        RECT 64.085 41.365 65.015 41.595 ;
        RECT 64.085 40.685 67.985 41.365 ;
        RECT 68.225 40.685 69.595 41.495 ;
        RECT 69.605 41.365 70.950 41.595 ;
        RECT 69.605 40.685 71.435 41.365 ;
        RECT 71.445 40.685 74.920 41.595 ;
        RECT 75.125 40.685 76.495 41.495 ;
        RECT 76.515 40.770 76.945 41.555 ;
        RECT 76.965 40.685 80.175 41.595 ;
        RECT 84.620 41.365 85.530 41.585 ;
        RECT 87.065 41.365 88.415 41.595 ;
        RECT 81.105 40.685 88.415 41.365 ;
        RECT 88.465 40.685 89.835 41.495 ;
        RECT 12.245 40.475 12.415 40.685 ;
        RECT 13.625 40.635 13.795 40.665 ;
        RECT 13.620 40.525 13.795 40.635 ;
        RECT 13.625 40.475 13.795 40.525 ;
        RECT 14.085 40.495 14.255 40.685 ;
        RECT 17.305 40.495 17.475 40.685 ;
        RECT 19.140 40.525 19.260 40.635 ;
        RECT 19.605 40.475 19.775 40.665 ;
        RECT 20.525 40.495 20.695 40.685 ;
        RECT 22.825 40.475 22.995 40.685 ;
        RECT 25.585 40.495 25.755 40.685 ;
        RECT 32.025 40.475 32.195 40.665 ;
        RECT 32.485 40.475 32.655 40.665 ;
        RECT 32.950 40.495 33.120 40.685 ;
        RECT 34.325 40.495 34.495 40.685 ;
        RECT 36.165 40.475 36.335 40.665 ;
        RECT 36.625 40.475 36.795 40.665 ;
        RECT 38.465 40.475 38.635 40.665 ;
        RECT 41.225 40.475 41.395 40.665 ;
        RECT 43.525 40.495 43.695 40.685 ;
        RECT 43.985 40.495 44.155 40.685 ;
        RECT 46.750 40.665 46.920 40.685 ;
        RECT 46.745 40.495 46.920 40.665 ;
        RECT 47.205 40.495 47.375 40.685 ;
        RECT 51.345 40.495 51.515 40.685 ;
        RECT 46.745 40.475 46.915 40.495 ;
        RECT 52.265 40.475 52.435 40.665 ;
        RECT 55.030 40.475 55.200 40.665 ;
        RECT 55.490 40.475 55.660 40.665 ;
        RECT 55.945 40.495 56.115 40.685 ;
        RECT 57.335 40.520 57.495 40.630 ;
        RECT 59.625 40.495 59.795 40.685 ;
        RECT 60.085 40.475 60.255 40.685 ;
        RECT 12.105 39.665 13.475 40.475 ;
        RECT 13.485 39.665 18.995 40.475 ;
        RECT 19.505 39.565 22.675 40.475 ;
        RECT 22.685 39.795 29.995 40.475 ;
        RECT 26.200 39.575 27.110 39.795 ;
        RECT 28.645 39.565 29.995 39.795 ;
        RECT 30.045 39.795 32.335 40.475 ;
        RECT 30.045 39.565 30.965 39.795 ;
        RECT 32.345 39.665 33.715 40.475 ;
        RECT 33.725 39.795 36.475 40.475 ;
        RECT 33.725 39.565 34.655 39.795 ;
        RECT 36.485 39.665 37.855 40.475 ;
        RECT 37.875 39.605 38.305 40.390 ;
        RECT 38.335 39.565 41.065 40.475 ;
        RECT 41.085 39.665 46.595 40.475 ;
        RECT 46.605 39.665 52.115 40.475 ;
        RECT 52.125 39.665 53.955 40.475 ;
        RECT 53.965 39.565 55.315 40.475 ;
        RECT 55.345 39.565 57.175 40.475 ;
        RECT 58.105 39.795 60.395 40.475 ;
        RECT 60.550 40.445 60.720 40.665 ;
        RECT 63.760 40.525 63.880 40.635 ;
        RECT 62.680 40.445 63.615 40.475 ;
        RECT 60.550 40.245 63.615 40.445 ;
        RECT 64.225 40.445 64.395 40.665 ;
        RECT 64.500 40.495 64.670 40.685 ;
        RECT 67.455 40.520 67.615 40.630 ;
        RECT 68.365 40.495 68.535 40.685 ;
        RECT 69.745 40.475 69.915 40.665 ;
        RECT 71.125 40.495 71.295 40.685 ;
        RECT 71.590 40.665 71.760 40.685 ;
        RECT 71.585 40.495 71.760 40.665 ;
        RECT 73.885 40.495 74.055 40.665 ;
        RECT 75.265 40.495 75.435 40.685 ;
        RECT 76.185 40.495 76.355 40.665 ;
        RECT 76.640 40.525 76.760 40.635 ;
        RECT 77.105 40.495 77.275 40.685 ;
        RECT 78.945 40.495 79.115 40.665 ;
        RECT 71.585 40.475 71.755 40.495 ;
        RECT 73.885 40.475 74.050 40.495 ;
        RECT 76.185 40.475 76.350 40.495 ;
        RECT 78.945 40.475 79.110 40.495 ;
        RECT 79.405 40.475 79.575 40.665 ;
        RECT 80.335 40.530 80.495 40.640 ;
        RECT 81.245 40.495 81.415 40.685 ;
        RECT 84.460 40.475 84.630 40.665 ;
        RECT 87.685 40.475 87.855 40.665 ;
        RECT 88.140 40.525 88.260 40.635 ;
        RECT 89.525 40.475 89.695 40.685 ;
        RECT 66.350 40.445 67.295 40.475 ;
        RECT 58.105 39.565 59.025 39.795 ;
        RECT 60.405 39.765 63.615 40.245 ;
        RECT 60.405 39.565 61.335 39.765 ;
        RECT 62.665 39.565 63.615 39.765 ;
        RECT 63.635 39.605 64.065 40.390 ;
        RECT 64.225 40.245 67.295 40.445 ;
        RECT 64.085 39.765 67.295 40.245 ;
        RECT 64.085 39.565 65.015 39.765 ;
        RECT 66.350 39.565 67.295 39.765 ;
        RECT 68.225 39.795 70.055 40.475 ;
        RECT 70.065 39.795 71.895 40.475 ;
        RECT 72.215 39.795 74.050 40.475 ;
        RECT 74.515 39.795 76.350 40.475 ;
        RECT 77.275 39.795 79.110 40.475 ;
        RECT 79.265 39.795 81.095 40.475 ;
        RECT 68.225 39.565 69.570 39.795 ;
        RECT 70.065 39.565 71.410 39.795 ;
        RECT 72.215 39.565 73.145 39.795 ;
        RECT 74.515 39.565 75.445 39.795 ;
        RECT 77.275 39.565 78.205 39.795 ;
        RECT 79.750 39.565 81.095 39.795 ;
        RECT 81.300 39.565 84.775 40.475 ;
        RECT 84.785 39.565 87.995 40.475 ;
        RECT 88.465 39.665 89.835 40.475 ;
      LAYER nwell ;
        RECT 11.910 36.445 90.030 39.275 ;
      LAYER pwell ;
        RECT 12.105 35.245 13.475 36.055 ;
        RECT 13.485 35.245 18.995 36.055 ;
        RECT 19.005 35.245 24.515 36.055 ;
        RECT 24.995 35.330 25.425 36.115 ;
        RECT 25.485 35.925 26.835 36.155 ;
        RECT 28.370 35.925 29.280 36.145 ;
        RECT 36.320 35.925 37.230 36.145 ;
        RECT 38.765 35.925 40.115 36.155 ;
        RECT 25.485 35.245 32.795 35.925 ;
        RECT 32.805 35.245 40.115 35.925 ;
        RECT 40.165 35.245 45.675 36.055 ;
        RECT 45.685 35.245 49.355 36.055 ;
        RECT 49.365 35.245 50.735 36.055 ;
        RECT 50.755 35.330 51.185 36.115 ;
        RECT 51.205 35.245 56.715 36.055 ;
        RECT 56.725 35.245 58.555 36.055 ;
        RECT 59.045 35.245 60.395 36.155 ;
        RECT 60.405 35.245 61.755 36.155 ;
        RECT 61.785 35.245 63.155 36.055 ;
        RECT 63.175 35.245 64.525 36.155 ;
        RECT 64.545 35.245 65.915 36.055 ;
        RECT 65.925 35.925 67.270 36.155 ;
        RECT 67.765 35.925 69.110 36.155 ;
        RECT 69.915 35.925 70.845 36.155 ;
        RECT 72.955 35.925 73.885 36.155 ;
        RECT 75.255 35.925 76.185 36.155 ;
        RECT 65.925 35.245 67.755 35.925 ;
        RECT 67.765 35.245 69.595 35.925 ;
        RECT 69.915 35.245 71.750 35.925 ;
        RECT 12.245 35.035 12.415 35.245 ;
        RECT 13.625 35.035 13.795 35.245 ;
        RECT 19.145 35.035 19.315 35.245 ;
        RECT 24.665 35.195 24.835 35.225 ;
        RECT 24.660 35.085 24.835 35.195 ;
        RECT 24.665 35.035 24.835 35.085 ;
        RECT 30.185 35.035 30.355 35.225 ;
        RECT 32.485 35.055 32.655 35.245 ;
        RECT 32.945 35.055 33.115 35.245 ;
        RECT 35.705 35.035 35.875 35.225 ;
        RECT 37.540 35.085 37.660 35.195 ;
        RECT 38.465 35.035 38.635 35.225 ;
        RECT 40.305 35.055 40.475 35.245 ;
        RECT 43.985 35.035 44.155 35.225 ;
        RECT 45.825 35.055 45.995 35.245 ;
        RECT 49.505 35.035 49.675 35.245 ;
        RECT 51.345 35.055 51.515 35.245 ;
        RECT 55.025 35.035 55.195 35.225 ;
        RECT 56.865 35.055 57.035 35.245 ;
        RECT 57.330 35.035 57.500 35.225 ;
        RECT 58.700 35.085 58.820 35.195 ;
        RECT 59.160 35.055 59.330 35.245 ;
        RECT 60.550 35.225 60.720 35.245 ;
        RECT 59.625 35.055 59.795 35.225 ;
        RECT 60.080 35.085 60.200 35.195 ;
        RECT 60.545 35.055 60.720 35.225 ;
        RECT 61.925 35.055 62.095 35.245 ;
        RECT 63.305 35.055 63.475 35.245 ;
        RECT 64.220 35.085 64.340 35.195 ;
        RECT 64.685 35.055 64.855 35.245 ;
        RECT 59.625 35.035 59.790 35.055 ;
        RECT 12.105 34.225 13.475 35.035 ;
        RECT 13.485 34.225 18.995 35.035 ;
        RECT 19.005 34.225 24.515 35.035 ;
        RECT 24.525 34.225 30.035 35.035 ;
        RECT 30.045 34.225 35.555 35.035 ;
        RECT 35.565 34.225 37.395 35.035 ;
        RECT 37.875 34.165 38.305 34.950 ;
        RECT 38.325 34.225 43.835 35.035 ;
        RECT 43.845 34.225 49.355 35.035 ;
        RECT 49.365 34.225 54.875 35.035 ;
        RECT 54.885 34.225 56.255 35.035 ;
        RECT 56.265 34.125 57.615 35.035 ;
        RECT 57.955 34.355 59.790 35.035 ;
        RECT 60.545 35.005 60.715 35.055 ;
        RECT 64.960 35.035 65.130 35.225 ;
        RECT 67.445 35.055 67.615 35.245 ;
        RECT 69.100 35.035 69.270 35.225 ;
        RECT 69.285 35.055 69.455 35.245 ;
        RECT 71.585 35.225 71.750 35.245 ;
        RECT 72.050 35.245 73.885 35.925 ;
        RECT 74.350 35.245 76.185 35.925 ;
        RECT 76.515 35.330 76.945 36.115 ;
        RECT 76.965 35.245 80.175 36.155 ;
        RECT 80.185 35.245 83.395 36.155 ;
        RECT 83.865 35.245 87.340 36.155 ;
        RECT 88.465 35.245 89.835 36.055 ;
        RECT 72.050 35.225 72.215 35.245 ;
        RECT 74.350 35.225 74.515 35.245 ;
        RECT 71.585 35.055 71.755 35.225 ;
        RECT 72.045 35.055 72.215 35.225 ;
        RECT 72.970 35.035 73.140 35.225 ;
        RECT 74.345 35.055 74.515 35.225 ;
        RECT 77.105 35.055 77.275 35.245 ;
        RECT 79.865 35.035 80.035 35.225 ;
        RECT 80.330 35.035 80.500 35.225 ;
        RECT 83.085 35.055 83.255 35.245 ;
        RECT 83.540 35.085 83.660 35.195 ;
        RECT 84.010 35.035 84.180 35.245 ;
        RECT 87.695 35.080 87.855 35.200 ;
        RECT 89.525 35.035 89.695 35.245 ;
        RECT 62.670 35.005 63.615 35.035 ;
        RECT 60.545 34.805 63.615 35.005 ;
        RECT 57.955 34.125 58.885 34.355 ;
        RECT 60.405 34.325 63.615 34.805 ;
        RECT 60.405 34.125 61.335 34.325 ;
        RECT 62.670 34.125 63.615 34.325 ;
        RECT 63.635 34.165 64.065 34.950 ;
        RECT 64.545 34.355 68.445 35.035 ;
        RECT 68.685 34.355 72.585 35.035 ;
        RECT 64.545 34.125 65.475 34.355 ;
        RECT 68.685 34.125 69.615 34.355 ;
        RECT 72.825 34.125 76.300 35.035 ;
        RECT 76.600 34.355 80.065 35.035 ;
        RECT 76.600 34.125 77.520 34.355 ;
        RECT 80.185 34.125 83.660 35.035 ;
        RECT 83.865 34.125 87.340 35.035 ;
        RECT 88.465 34.225 89.835 35.035 ;
      LAYER nwell ;
        RECT 11.910 31.005 90.030 33.835 ;
      LAYER pwell ;
        RECT 12.105 29.805 13.475 30.615 ;
        RECT 13.485 29.805 18.995 30.615 ;
        RECT 19.005 29.805 24.515 30.615 ;
        RECT 24.995 29.890 25.425 30.675 ;
        RECT 25.445 29.805 30.955 30.615 ;
        RECT 30.965 29.805 36.475 30.615 ;
        RECT 36.485 29.805 41.995 30.615 ;
        RECT 42.005 29.805 47.515 30.615 ;
        RECT 47.525 29.805 50.275 30.615 ;
        RECT 50.755 29.890 51.185 30.675 ;
        RECT 51.205 29.805 53.035 30.715 ;
        RECT 54.185 30.625 55.135 30.715 ;
        RECT 53.205 29.805 55.135 30.625 ;
        RECT 58.860 30.485 59.770 30.705 ;
        RECT 61.305 30.485 62.655 30.715 ;
        RECT 67.140 30.485 68.050 30.705 ;
        RECT 69.585 30.485 71.355 30.715 ;
        RECT 55.345 29.805 62.655 30.485 ;
        RECT 63.625 29.805 71.355 30.485 ;
        RECT 71.445 30.485 72.375 30.715 ;
        RECT 71.445 29.805 75.345 30.485 ;
        RECT 76.515 29.890 76.945 30.675 ;
        RECT 77.005 30.485 78.355 30.715 ;
        RECT 79.890 30.485 80.800 30.705 ;
        RECT 77.005 29.805 84.315 30.485 ;
        RECT 84.325 29.805 87.800 30.715 ;
        RECT 88.465 29.805 89.835 30.615 ;
        RECT 12.245 29.595 12.415 29.805 ;
        RECT 13.625 29.595 13.795 29.805 ;
        RECT 19.145 29.595 19.315 29.805 ;
        RECT 24.665 29.755 24.835 29.785 ;
        RECT 24.660 29.645 24.835 29.755 ;
        RECT 24.665 29.595 24.835 29.645 ;
        RECT 25.585 29.615 25.755 29.805 ;
        RECT 30.185 29.595 30.355 29.785 ;
        RECT 31.105 29.615 31.275 29.805 ;
        RECT 35.705 29.595 35.875 29.785 ;
        RECT 36.625 29.615 36.795 29.805 ;
        RECT 37.540 29.645 37.660 29.755 ;
        RECT 38.465 29.595 38.635 29.785 ;
        RECT 42.145 29.615 42.315 29.805 ;
        RECT 43.985 29.595 44.155 29.785 ;
        RECT 47.665 29.615 47.835 29.805 ;
        RECT 48.585 29.615 48.755 29.785 ;
        RECT 50.420 29.645 50.540 29.755 ;
        RECT 50.885 29.615 51.055 29.785 ;
        RECT 48.585 29.595 48.750 29.615 ;
        RECT 50.885 29.595 51.035 29.615 ;
        RECT 51.350 29.595 51.520 29.805 ;
        RECT 53.205 29.785 53.355 29.805 ;
        RECT 53.185 29.615 53.355 29.785 ;
        RECT 55.035 29.640 55.195 29.750 ;
        RECT 55.485 29.615 55.655 29.805 ;
        RECT 55.945 29.595 56.115 29.785 ;
        RECT 62.855 29.650 63.015 29.760 ;
        RECT 63.765 29.615 63.935 29.805 ;
        RECT 71.585 29.595 71.755 29.785 ;
        RECT 71.860 29.615 72.030 29.805 ;
        RECT 72.045 29.595 72.215 29.785 ;
        RECT 75.735 29.650 75.895 29.760 ;
        RECT 79.400 29.645 79.520 29.755 ;
        RECT 84.005 29.615 84.175 29.805 ;
        RECT 84.470 29.615 84.640 29.805 ;
        RECT 86.765 29.595 86.935 29.785 ;
        RECT 87.225 29.595 87.395 29.785 ;
        RECT 88.140 29.645 88.260 29.755 ;
        RECT 89.525 29.595 89.695 29.805 ;
        RECT 12.105 28.785 13.475 29.595 ;
        RECT 13.485 28.785 18.995 29.595 ;
        RECT 19.005 28.785 24.515 29.595 ;
        RECT 24.525 28.785 30.035 29.595 ;
        RECT 30.045 28.785 35.555 29.595 ;
        RECT 35.565 28.785 37.395 29.595 ;
        RECT 37.875 28.725 38.305 29.510 ;
        RECT 38.325 28.785 43.835 29.595 ;
        RECT 43.845 28.785 46.595 29.595 ;
        RECT 46.915 28.915 48.750 29.595 ;
        RECT 46.915 28.685 47.845 28.915 ;
        RECT 49.105 28.775 51.035 29.595 ;
        RECT 49.105 28.685 50.055 28.775 ;
        RECT 51.205 28.685 54.875 29.595 ;
        RECT 55.805 28.915 63.535 29.595 ;
        RECT 59.320 28.695 60.230 28.915 ;
        RECT 61.765 28.685 63.535 28.915 ;
        RECT 63.635 28.725 64.065 29.510 ;
        RECT 64.165 28.915 71.895 29.595 ;
        RECT 71.905 28.915 79.215 29.595 ;
        RECT 64.165 28.685 65.935 28.915 ;
        RECT 67.470 28.695 68.380 28.915 ;
        RECT 75.420 28.695 76.330 28.915 ;
        RECT 77.865 28.685 79.215 28.915 ;
        RECT 79.765 28.915 87.075 29.595 ;
        RECT 79.765 28.685 81.115 28.915 ;
        RECT 82.650 28.695 83.560 28.915 ;
        RECT 87.085 28.785 88.455 29.595 ;
        RECT 88.465 28.785 89.835 29.595 ;
      LAYER nwell ;
        RECT 11.910 25.565 90.030 28.395 ;
      LAYER pwell ;
        RECT 12.105 24.365 13.475 25.175 ;
        RECT 13.485 24.365 18.995 25.175 ;
        RECT 19.005 24.365 24.515 25.175 ;
        RECT 24.995 24.450 25.425 25.235 ;
        RECT 25.445 24.365 30.955 25.175 ;
        RECT 30.965 24.365 36.475 25.175 ;
        RECT 36.485 24.365 41.995 25.175 ;
        RECT 42.005 24.365 47.515 25.175 ;
        RECT 47.525 24.365 49.355 25.175 ;
        RECT 49.365 24.365 50.735 25.145 ;
        RECT 50.755 24.450 51.185 25.235 ;
        RECT 54.780 25.045 55.700 25.275 ;
        RECT 59.320 25.045 60.230 25.265 ;
        RECT 61.765 25.045 63.115 25.275 ;
        RECT 64.535 25.045 65.455 25.275 ;
        RECT 69.900 25.045 70.810 25.265 ;
        RECT 72.345 25.045 73.695 25.275 ;
        RECT 74.795 25.045 75.725 25.275 ;
        RECT 52.235 24.365 55.700 25.045 ;
        RECT 55.805 24.365 63.115 25.045 ;
        RECT 63.165 24.365 65.455 25.045 ;
        RECT 66.385 24.365 73.695 25.045 ;
        RECT 73.890 24.365 75.725 25.045 ;
        RECT 76.515 24.450 76.945 25.235 ;
        RECT 76.965 24.365 80.440 25.275 ;
        RECT 84.620 25.045 85.530 25.265 ;
        RECT 87.065 25.045 88.415 25.275 ;
        RECT 81.105 24.365 88.415 25.045 ;
        RECT 88.465 24.365 89.835 25.175 ;
        RECT 12.245 24.155 12.415 24.365 ;
        RECT 13.625 24.155 13.795 24.365 ;
        RECT 19.145 24.155 19.315 24.365 ;
        RECT 24.665 24.315 24.835 24.345 ;
        RECT 24.660 24.205 24.835 24.315 ;
        RECT 24.665 24.155 24.835 24.205 ;
        RECT 25.585 24.175 25.755 24.365 ;
        RECT 30.185 24.155 30.355 24.345 ;
        RECT 31.105 24.175 31.275 24.365 ;
        RECT 35.705 24.155 35.875 24.345 ;
        RECT 36.625 24.175 36.795 24.365 ;
        RECT 37.540 24.205 37.660 24.315 ;
        RECT 38.465 24.155 38.635 24.345 ;
        RECT 42.145 24.175 42.315 24.365 ;
        RECT 43.985 24.155 44.155 24.345 ;
        RECT 46.745 24.155 46.915 24.345 ;
        RECT 47.665 24.175 47.835 24.365 ;
        RECT 50.425 24.175 50.595 24.365 ;
        RECT 51.355 24.210 51.515 24.320 ;
        RECT 52.265 24.175 52.435 24.365 ;
        RECT 54.105 24.155 54.275 24.345 ;
        RECT 55.945 24.175 56.115 24.365 ;
        RECT 57.795 24.200 57.955 24.310 ;
        RECT 58.980 24.155 59.150 24.345 ;
        RECT 62.855 24.200 63.015 24.310 ;
        RECT 63.305 24.175 63.475 24.365 ;
        RECT 64.225 24.155 64.395 24.345 ;
        RECT 65.615 24.210 65.775 24.320 ;
        RECT 66.525 24.175 66.695 24.365 ;
        RECT 73.890 24.345 74.055 24.365 ;
        RECT 69.740 24.205 69.860 24.315 ;
        RECT 70.205 24.155 70.375 24.345 ;
        RECT 73.885 24.175 74.055 24.345 ;
        RECT 76.180 24.205 76.300 24.315 ;
        RECT 77.110 24.175 77.280 24.365 ;
        RECT 77.565 24.155 77.735 24.345 ;
        RECT 78.945 24.175 79.115 24.345 ;
        RECT 80.780 24.205 80.900 24.315 ;
        RECT 78.950 24.155 79.115 24.175 ;
        RECT 81.245 24.155 81.415 24.365 ;
        RECT 89.525 24.155 89.695 24.365 ;
        RECT 12.105 23.345 13.475 24.155 ;
        RECT 13.485 23.345 18.995 24.155 ;
        RECT 19.005 23.345 24.515 24.155 ;
        RECT 24.525 23.345 30.035 24.155 ;
        RECT 30.045 23.345 35.555 24.155 ;
        RECT 35.565 23.345 37.395 24.155 ;
        RECT 37.875 23.285 38.305 24.070 ;
        RECT 38.325 23.345 43.835 24.155 ;
        RECT 43.845 23.345 46.595 24.155 ;
        RECT 46.605 23.475 53.915 24.155 ;
        RECT 50.120 23.255 51.030 23.475 ;
        RECT 52.565 23.245 53.915 23.475 ;
        RECT 53.965 23.345 57.635 24.155 ;
        RECT 58.565 23.475 62.465 24.155 ;
        RECT 58.565 23.245 59.495 23.475 ;
        RECT 63.635 23.285 64.065 24.070 ;
        RECT 64.085 23.345 69.595 24.155 ;
        RECT 70.065 23.475 77.375 24.155 ;
        RECT 73.580 23.255 74.490 23.475 ;
        RECT 76.025 23.245 77.375 23.475 ;
        RECT 77.425 23.375 78.795 24.155 ;
        RECT 78.950 23.475 80.785 24.155 ;
        RECT 81.105 23.475 88.415 24.155 ;
        RECT 79.855 23.245 80.785 23.475 ;
        RECT 84.620 23.255 85.530 23.475 ;
        RECT 87.065 23.245 88.415 23.475 ;
        RECT 88.465 23.345 89.835 24.155 ;
      LAYER nwell ;
        RECT 11.910 20.125 90.030 22.955 ;
      LAYER pwell ;
        RECT 12.105 18.925 13.475 19.735 ;
        RECT 13.485 18.925 18.995 19.735 ;
        RECT 19.005 18.925 24.515 19.735 ;
        RECT 24.995 19.010 25.425 19.795 ;
        RECT 25.445 18.925 30.955 19.735 ;
        RECT 30.965 18.925 36.475 19.735 ;
        RECT 36.485 18.925 37.855 19.735 ;
        RECT 37.875 19.010 38.305 19.795 ;
        RECT 38.325 18.925 41.995 19.735 ;
        RECT 43.125 19.605 47.055 19.835 ;
        RECT 48.905 19.605 50.250 19.835 ;
        RECT 42.640 18.925 47.055 19.605 ;
        RECT 47.065 18.925 48.895 19.605 ;
        RECT 48.905 18.925 50.735 19.605 ;
        RECT 50.755 19.010 51.185 19.795 ;
        RECT 52.125 19.605 53.470 19.835 ;
        RECT 52.125 18.925 53.955 19.605 ;
        RECT 53.965 18.925 55.335 19.735 ;
        RECT 55.345 18.925 57.175 19.605 ;
        RECT 57.185 18.925 62.695 19.735 ;
        RECT 63.635 19.010 64.065 19.795 ;
        RECT 64.085 18.925 69.595 19.735 ;
        RECT 69.605 18.925 71.435 19.735 ;
        RECT 71.445 19.605 72.790 19.835 ;
        RECT 71.445 18.925 73.275 19.605 ;
        RECT 73.285 18.925 74.655 19.735 ;
        RECT 74.665 19.605 76.010 19.835 ;
        RECT 74.665 18.925 76.495 19.605 ;
        RECT 76.515 19.010 76.945 19.795 ;
        RECT 77.885 19.605 79.230 19.835 ;
        RECT 80.210 19.605 81.555 19.835 ;
        RECT 82.050 19.605 83.395 19.835 ;
        RECT 84.455 19.605 85.385 19.835 ;
        RECT 87.110 19.605 88.455 19.835 ;
        RECT 77.885 18.925 79.715 19.605 ;
        RECT 79.725 18.925 81.555 19.605 ;
        RECT 81.565 18.925 83.395 19.605 ;
        RECT 83.550 18.925 85.385 19.605 ;
        RECT 86.625 18.925 88.455 19.605 ;
        RECT 88.465 18.925 89.835 19.735 ;
        RECT 12.245 18.735 12.415 18.925 ;
        RECT 13.625 18.735 13.795 18.925 ;
        RECT 19.145 18.735 19.315 18.925 ;
        RECT 24.660 18.765 24.780 18.875 ;
        RECT 25.585 18.735 25.755 18.925 ;
        RECT 31.105 18.735 31.275 18.925 ;
        RECT 36.625 18.735 36.795 18.925 ;
        RECT 38.465 18.735 38.635 18.925 ;
        RECT 42.640 18.905 42.750 18.925 ;
        RECT 42.140 18.765 42.260 18.875 ;
        RECT 42.580 18.735 42.750 18.905 ;
        RECT 47.205 18.735 47.375 18.925 ;
        RECT 50.425 18.735 50.595 18.925 ;
        RECT 51.355 18.770 51.515 18.880 ;
        RECT 53.645 18.735 53.815 18.925 ;
        RECT 54.105 18.735 54.275 18.925 ;
        RECT 55.485 18.735 55.655 18.925 ;
        RECT 57.325 18.735 57.495 18.925 ;
        RECT 62.855 18.770 63.015 18.880 ;
        RECT 64.225 18.735 64.395 18.925 ;
        RECT 69.745 18.735 69.915 18.925 ;
        RECT 72.965 18.735 73.135 18.925 ;
        RECT 73.425 18.735 73.595 18.925 ;
        RECT 76.185 18.735 76.355 18.925 ;
        RECT 77.115 18.770 77.275 18.880 ;
        RECT 79.405 18.735 79.575 18.925 ;
        RECT 79.865 18.735 80.035 18.925 ;
        RECT 81.705 18.735 81.875 18.925 ;
        RECT 83.550 18.905 83.715 18.925 ;
        RECT 83.545 18.735 83.715 18.905 ;
        RECT 85.855 18.770 86.015 18.880 ;
        RECT 86.765 18.735 86.935 18.925 ;
        RECT 89.525 18.735 89.695 18.925 ;
      LAYER li1 ;
        RECT 112.275 219.210 112.445 219.295 ;
        RECT 114.995 219.210 115.165 219.295 ;
        RECT 117.715 219.210 117.885 219.295 ;
        RECT 120.435 219.210 120.605 219.295 ;
        RECT 123.155 219.210 123.325 219.295 ;
        RECT 125.875 219.210 126.045 219.295 ;
        RECT 128.595 219.210 128.765 219.295 ;
        RECT 131.315 219.210 131.485 219.295 ;
        RECT 134.035 219.210 134.205 219.295 ;
        RECT 136.755 219.210 136.925 219.295 ;
        RECT 139.475 219.210 139.645 219.295 ;
        RECT 142.195 219.210 142.365 219.295 ;
        RECT 144.915 219.210 145.085 219.295 ;
        RECT 147.635 219.210 147.805 219.295 ;
        RECT 112.275 218.690 113.735 219.210 ;
        RECT 112.275 218.000 113.195 218.690 ;
        RECT 113.905 218.520 116.255 219.210 ;
        RECT 116.425 218.690 119.175 219.210 ;
        RECT 113.365 218.000 116.795 218.520 ;
        RECT 116.965 218.000 118.635 218.690 ;
        RECT 119.345 218.520 121.695 219.210 ;
        RECT 121.865 218.690 124.615 219.210 ;
        RECT 118.805 218.000 122.235 218.520 ;
        RECT 122.405 218.000 124.075 218.690 ;
        RECT 124.785 218.520 127.135 219.210 ;
        RECT 127.305 218.690 130.055 219.210 ;
        RECT 124.245 218.000 127.675 218.520 ;
        RECT 127.845 218.000 129.515 218.690 ;
        RECT 130.225 218.520 132.575 219.210 ;
        RECT 132.745 218.690 135.495 219.210 ;
        RECT 129.685 218.000 133.115 218.520 ;
        RECT 133.285 218.000 134.955 218.690 ;
        RECT 135.665 218.520 138.015 219.210 ;
        RECT 138.185 218.690 140.935 219.210 ;
        RECT 135.125 218.000 138.555 218.520 ;
        RECT 138.725 218.000 140.395 218.690 ;
        RECT 141.105 218.520 143.455 219.210 ;
        RECT 143.625 218.690 146.375 219.210 ;
        RECT 140.565 218.000 143.995 218.520 ;
        RECT 144.165 218.000 145.835 218.690 ;
        RECT 146.545 218.520 147.805 219.210 ;
        RECT 146.005 218.000 147.805 218.520 ;
        RECT 112.275 217.830 112.445 218.000 ;
        RECT 114.995 217.830 115.165 218.000 ;
        RECT 112.275 216.245 112.990 217.830 ;
        RECT 114.560 217.825 115.165 217.830 ;
        RECT 117.715 217.825 117.885 218.000 ;
        RECT 114.560 217.565 116.315 217.825 ;
        RECT 116.875 217.565 117.885 217.825 ;
        RECT 118.540 217.780 119.375 217.830 ;
        RECT 114.560 216.965 115.165 217.565 ;
        RECT 115.335 217.220 117.545 217.390 ;
        RECT 115.335 217.135 116.240 217.220 ;
        RECT 116.970 217.135 117.545 217.220 ;
        RECT 117.715 217.280 117.885 217.565 ;
        RECT 118.105 217.770 119.375 217.780 ;
        RECT 120.435 217.825 120.605 218.000 ;
        RECT 123.155 217.825 123.325 218.000 ;
        RECT 125.875 217.825 126.045 218.000 ;
        RECT 128.595 217.830 128.765 218.000 ;
        RECT 131.315 217.830 131.485 218.000 ;
        RECT 128.595 217.825 130.055 217.830 ;
        RECT 118.105 217.660 120.220 217.770 ;
        RECT 118.105 217.605 118.665 217.660 ;
        RECT 119.245 217.615 120.220 217.660 ;
        RECT 118.105 217.450 118.625 217.605 ;
        RECT 117.715 217.110 118.495 217.280 ;
        RECT 116.475 216.965 116.805 217.050 ;
        RECT 117.715 216.965 117.885 217.110 ;
        RECT 114.560 216.635 115.925 216.965 ;
        RECT 116.095 216.795 117.165 216.965 ;
        RECT 112.275 215.905 113.820 216.245 ;
        RECT 112.275 212.485 112.990 215.905 ;
        RECT 114.560 214.560 115.165 216.635 ;
        RECT 116.095 216.420 116.265 216.795 ;
        RECT 115.335 216.250 116.265 216.420 ;
        RECT 116.445 216.160 116.815 216.515 ;
        RECT 116.995 216.420 117.165 216.795 ;
        RECT 117.335 216.635 117.885 216.965 ;
        RECT 118.795 216.940 119.125 217.490 ;
        RECT 119.295 217.440 120.220 217.615 ;
        RECT 120.435 217.565 121.755 217.825 ;
        RECT 122.315 217.565 123.325 217.825 ;
        RECT 123.585 217.570 124.045 217.740 ;
        RECT 120.435 217.270 120.605 217.565 ;
        RECT 123.155 217.400 123.325 217.565 ;
        RECT 119.425 217.100 120.605 217.270 ;
        RECT 120.775 217.220 122.985 217.390 ;
        RECT 120.775 217.135 121.680 217.220 ;
        RECT 122.410 217.135 122.985 217.220 ;
        RECT 116.995 216.250 117.545 216.420 ;
        RECT 117.715 216.350 117.885 216.635 ;
        RECT 118.100 216.930 119.125 216.940 ;
        RECT 120.435 216.965 120.605 217.100 ;
        RECT 123.155 217.070 123.705 217.400 ;
        RECT 123.875 217.305 124.045 217.570 ;
        RECT 124.215 217.475 124.865 217.825 ;
        RECT 125.035 217.570 125.705 217.740 ;
        RECT 125.035 217.305 125.205 217.570 ;
        RECT 125.875 217.565 127.195 217.825 ;
        RECT 127.755 217.565 130.055 217.825 ;
        RECT 125.875 217.400 126.045 217.565 ;
        RECT 123.875 217.075 125.205 217.305 ;
        RECT 125.375 217.070 126.045 217.400 ;
        RECT 126.215 217.220 128.425 217.390 ;
        RECT 126.215 217.135 127.120 217.220 ;
        RECT 127.850 217.135 128.425 217.220 ;
        RECT 128.595 217.310 130.055 217.565 ;
        RECT 121.915 216.965 122.245 217.050 ;
        RECT 123.155 216.965 123.325 217.070 ;
        RECT 118.100 216.740 120.265 216.930 ;
        RECT 118.100 216.610 118.625 216.740 ;
        RECT 119.330 216.590 120.265 216.740 ;
        RECT 120.435 216.635 121.365 216.965 ;
        RECT 121.535 216.795 122.605 216.965 ;
        RECT 117.715 216.140 118.415 216.350 ;
        RECT 115.335 214.895 117.545 215.065 ;
        RECT 115.335 214.730 116.305 214.895 ;
        RECT 116.975 214.810 117.545 214.895 ;
        RECT 116.475 214.640 116.805 214.725 ;
        RECT 117.715 214.640 117.885 216.140 ;
        RECT 118.795 215.865 119.125 216.570 ;
        RECT 119.330 216.035 119.705 216.590 ;
        RECT 120.435 216.360 120.605 216.635 ;
        RECT 121.535 216.420 121.705 216.795 ;
        RECT 119.935 216.045 120.605 216.360 ;
        RECT 120.775 216.250 121.705 216.420 ;
        RECT 121.885 216.160 122.255 216.515 ;
        RECT 122.435 216.420 122.605 216.795 ;
        RECT 122.775 216.635 123.325 216.965 ;
        RECT 125.875 216.965 126.045 217.070 ;
        RECT 127.355 216.965 127.685 217.050 ;
        RECT 128.595 216.965 129.515 217.310 ;
        RECT 130.225 217.270 131.485 217.830 ;
        RECT 132.545 217.780 133.380 217.830 ;
        RECT 132.545 217.770 133.815 217.780 ;
        RECT 131.700 217.660 133.815 217.770 ;
        RECT 131.700 217.615 132.675 217.660 ;
        RECT 131.700 217.440 132.625 217.615 ;
        RECT 133.255 217.605 133.815 217.660 ;
        RECT 130.225 217.140 132.495 217.270 ;
        RECT 123.585 216.715 125.705 216.900 ;
        RECT 123.155 216.460 123.325 216.635 ;
        RECT 125.875 216.635 126.805 216.965 ;
        RECT 126.975 216.795 128.045 216.965 ;
        RECT 122.435 216.250 122.985 216.420 ;
        RECT 123.155 216.210 123.785 216.460 ;
        RECT 123.955 216.265 124.905 216.545 ;
        RECT 125.875 216.475 126.045 216.635 ;
        RECT 125.415 216.210 126.045 216.475 ;
        RECT 126.975 216.420 127.145 216.795 ;
        RECT 126.215 216.250 127.145 216.420 ;
        RECT 118.165 215.695 120.135 215.865 ;
        RECT 118.165 215.080 118.335 215.695 ;
        RECT 118.505 215.205 119.795 215.525 ;
        RECT 118.505 215.060 118.835 215.205 ;
        RECT 114.560 214.425 116.305 214.560 ;
        RECT 116.475 214.470 117.145 214.640 ;
        RECT 113.310 214.390 116.305 214.425 ;
        RECT 113.310 214.075 115.165 214.390 ;
        RECT 116.475 214.220 116.805 214.245 ;
        RECT 114.560 212.485 115.165 214.075 ;
        RECT 112.275 212.310 112.445 212.485 ;
        RECT 114.995 212.310 115.165 212.485 ;
        RECT 112.275 210.660 113.735 212.310 ;
        RECT 113.905 212.020 115.165 212.310 ;
        RECT 115.335 214.050 116.805 214.220 ;
        RECT 115.335 212.360 115.505 214.050 ;
        RECT 116.975 213.885 117.145 214.470 ;
        RECT 117.315 214.325 117.885 214.640 ;
        RECT 118.165 214.675 118.335 214.910 ;
        RECT 119.045 214.845 119.765 215.035 ;
        RECT 119.965 214.980 120.135 215.695 ;
        RECT 119.935 214.675 120.265 214.755 ;
        RECT 118.165 214.505 120.265 214.675 ;
        RECT 117.315 214.310 118.385 214.325 ;
        RECT 117.715 213.955 118.385 214.310 ;
        RECT 118.565 214.045 118.865 214.505 ;
        RECT 120.435 214.500 120.605 216.045 ;
        RECT 120.775 214.670 121.455 214.955 ;
        RECT 120.435 214.335 121.065 214.500 ;
        RECT 119.045 214.165 119.375 214.335 ;
        RECT 119.635 214.230 121.065 214.335 ;
        RECT 119.635 214.165 120.605 214.230 ;
        RECT 116.975 213.880 117.545 213.885 ;
        RECT 115.675 213.710 117.545 213.880 ;
        RECT 115.675 212.755 115.845 213.710 ;
        RECT 116.015 213.370 116.985 213.540 ;
        RECT 116.015 212.720 116.185 213.370 ;
        RECT 117.180 213.355 117.545 213.710 ;
        RECT 117.205 213.165 117.375 213.170 ;
        RECT 116.385 212.890 117.545 213.165 ;
        RECT 116.015 212.530 117.545 212.720 ;
        RECT 115.335 212.190 116.360 212.360 ;
        RECT 117.715 212.350 117.885 213.955 ;
        RECT 118.565 213.845 118.895 214.045 ;
        RECT 119.115 213.995 119.375 214.165 ;
        RECT 119.115 213.825 120.160 213.995 ;
        RECT 119.115 213.635 119.285 213.825 ;
        RECT 118.165 213.465 119.285 213.635 ;
        RECT 118.165 212.960 118.335 213.465 ;
        RECT 119.455 213.295 119.820 213.655 ;
        RECT 118.535 213.125 119.820 213.295 ;
        RECT 118.535 212.770 118.755 213.125 ;
        RECT 118.165 212.600 118.335 212.765 ;
        RECT 118.925 212.715 119.520 212.955 ;
        RECT 119.990 212.890 120.160 213.825 ;
        RECT 118.165 212.545 118.605 212.600 ;
        RECT 119.710 212.545 120.265 212.680 ;
        RECT 118.165 212.430 120.265 212.545 ;
        RECT 120.435 212.440 120.605 214.165 ;
        RECT 121.235 214.210 121.455 214.670 ;
        RECT 121.625 214.380 122.185 215.070 ;
        RECT 122.355 214.670 122.985 214.955 ;
        RECT 122.355 214.210 122.525 214.670 ;
        RECT 123.155 214.515 123.325 216.210 ;
        RECT 123.915 216.040 125.280 216.095 ;
        RECT 123.605 215.925 125.705 216.040 ;
        RECT 123.605 215.870 124.045 215.925 ;
        RECT 123.605 215.705 123.775 215.870 ;
        RECT 125.150 215.790 125.705 215.925 ;
        RECT 123.605 215.005 123.775 215.510 ;
        RECT 123.975 215.345 124.195 215.700 ;
        RECT 124.365 215.515 124.960 215.755 ;
        RECT 123.975 215.175 125.260 215.345 ;
        RECT 123.605 214.835 124.725 215.005 ;
        RECT 124.555 214.645 124.725 214.835 ;
        RECT 124.895 214.815 125.260 215.175 ;
        RECT 125.430 214.645 125.600 215.580 ;
        RECT 123.155 214.500 123.825 214.515 ;
        RECT 122.695 214.230 123.825 214.500 ;
        RECT 121.235 214.000 122.525 214.210 ;
        RECT 123.155 214.145 123.825 214.230 ;
        RECT 124.005 214.425 124.335 214.625 ;
        RECT 124.555 214.475 125.600 214.645 ;
        RECT 125.875 215.020 126.045 216.210 ;
        RECT 127.325 216.160 127.695 216.515 ;
        RECT 127.875 216.420 128.045 216.795 ;
        RECT 128.215 216.635 129.515 216.965 ;
        RECT 128.595 216.620 129.515 216.635 ;
        RECT 129.685 217.100 132.495 217.140 ;
        RECT 129.685 216.620 131.485 217.100 ;
        RECT 132.795 216.940 133.125 217.490 ;
        RECT 133.295 217.450 133.815 217.605 ;
        RECT 134.035 217.400 134.205 218.000 ;
        RECT 136.755 217.825 136.925 218.000 ;
        RECT 139.475 217.825 139.645 218.000 ;
        RECT 142.195 217.830 142.365 218.000 ;
        RECT 144.915 217.830 145.085 218.000 ;
        RECT 147.635 217.830 147.805 218.000 ;
        RECT 134.375 217.655 136.585 217.825 ;
        RECT 134.375 217.570 134.945 217.655 ;
        RECT 135.615 217.490 136.585 217.655 ;
        RECT 136.755 217.565 138.075 217.825 ;
        RECT 138.635 217.565 139.645 217.825 ;
        RECT 139.905 217.570 140.365 217.740 ;
        RECT 135.115 217.400 135.445 217.485 ;
        RECT 134.035 217.280 134.605 217.400 ;
        RECT 133.425 217.110 134.605 217.280 ;
        RECT 134.035 217.070 134.605 217.110 ;
        RECT 134.775 217.230 135.445 217.400 ;
        RECT 136.755 217.320 136.925 217.565 ;
        RECT 139.475 217.400 139.645 217.565 ;
        RECT 132.795 216.930 133.820 216.940 ;
        RECT 127.875 216.250 128.425 216.420 ;
        RECT 128.595 215.880 128.765 216.620 ;
        RECT 128.935 216.050 129.565 216.335 ;
        RECT 128.595 215.610 129.225 215.880 ;
        RECT 126.215 215.355 128.425 215.525 ;
        RECT 126.215 215.190 127.185 215.355 ;
        RECT 127.855 215.270 128.425 215.355 ;
        RECT 127.355 215.100 127.685 215.185 ;
        RECT 128.595 215.100 128.765 215.610 ;
        RECT 129.395 215.590 129.565 216.050 ;
        RECT 129.735 215.760 130.295 216.450 ;
        RECT 131.315 216.360 131.485 216.620 ;
        RECT 131.655 216.740 133.820 216.930 ;
        RECT 131.655 216.590 132.590 216.740 ;
        RECT 133.295 216.610 133.820 216.740 ;
        RECT 130.465 216.050 131.145 216.335 ;
        RECT 130.465 215.590 130.685 216.050 ;
        RECT 131.315 216.045 131.985 216.360 ;
        RECT 131.315 215.880 131.485 216.045 ;
        RECT 132.215 216.035 132.590 216.590 ;
        RECT 130.855 215.610 131.485 215.880 ;
        RECT 132.795 215.865 133.125 216.570 ;
        RECT 134.035 216.350 134.205 217.070 ;
        RECT 134.775 216.645 134.945 217.230 ;
        RECT 135.615 217.150 136.925 217.320 ;
        RECT 135.115 216.980 135.445 217.005 ;
        RECT 135.115 216.810 136.585 216.980 ;
        RECT 133.505 216.140 134.205 216.350 ;
        RECT 129.395 215.380 130.685 215.590 ;
        RECT 125.875 214.850 127.185 215.020 ;
        RECT 127.355 214.930 128.025 215.100 ;
        RECT 120.775 213.430 122.985 213.830 ;
        RECT 120.775 212.960 121.455 213.240 ;
        RECT 121.235 212.565 121.455 212.960 ;
        RECT 121.625 212.735 122.185 213.430 ;
        RECT 122.355 212.960 122.985 213.240 ;
        RECT 122.355 212.565 122.525 212.960 ;
        RECT 118.475 212.375 119.840 212.430 ;
        RECT 113.905 211.850 115.925 212.020 ;
        RECT 113.905 210.930 115.165 211.850 ;
        RECT 115.515 211.440 115.925 211.615 ;
        RECT 116.170 211.610 116.360 212.190 ;
        RECT 116.735 211.620 116.905 212.330 ;
        RECT 117.180 212.260 117.885 212.350 ;
        RECT 120.435 212.260 121.065 212.440 ;
        RECT 117.180 212.010 118.345 212.260 ;
        RECT 117.180 211.840 117.885 212.010 ;
        RECT 118.515 211.925 119.465 212.205 ;
        RECT 119.975 212.115 121.065 212.260 ;
        RECT 121.235 212.115 122.525 212.565 ;
        RECT 123.155 212.440 123.325 214.145 ;
        RECT 124.005 213.965 124.305 214.425 ;
        RECT 124.555 214.305 124.815 214.475 ;
        RECT 125.875 214.305 126.045 214.850 ;
        RECT 127.355 214.680 127.685 214.705 ;
        RECT 124.485 214.135 124.815 214.305 ;
        RECT 125.075 214.135 126.045 214.305 ;
        RECT 123.605 213.795 125.705 213.965 ;
        RECT 123.605 213.560 123.775 213.795 ;
        RECT 125.375 213.715 125.705 213.795 ;
        RECT 124.485 213.435 125.205 213.625 ;
        RECT 123.605 212.775 123.775 213.390 ;
        RECT 123.945 213.265 124.275 213.410 ;
        RECT 123.945 212.945 125.235 213.265 ;
        RECT 125.405 212.775 125.575 213.490 ;
        RECT 123.605 212.605 125.575 212.775 ;
        RECT 122.695 212.330 123.325 212.440 ;
        RECT 122.695 212.120 123.855 212.330 ;
        RECT 122.695 212.115 123.325 212.120 ;
        RECT 119.975 211.995 120.605 212.115 ;
        RECT 121.915 212.010 122.245 212.115 ;
        RECT 116.735 211.440 117.510 211.620 ;
        RECT 115.515 211.375 117.510 211.440 ;
        RECT 117.715 211.400 117.885 211.840 ;
        RECT 118.145 211.570 120.265 211.755 ;
        RECT 120.435 211.400 120.605 211.995 ;
        RECT 120.775 211.840 121.745 211.945 ;
        RECT 122.415 211.840 122.985 211.945 ;
        RECT 120.775 211.560 122.985 211.840 ;
        RECT 115.515 211.100 116.905 211.375 ;
        RECT 117.715 211.070 118.265 211.400 ;
        RECT 118.435 211.165 119.765 211.395 ;
        RECT 117.715 210.930 117.885 211.070 ;
        RECT 112.275 208.800 113.215 210.660 ;
        RECT 113.905 210.490 116.255 210.930 ;
        RECT 113.385 209.110 116.255 210.490 ;
        RECT 116.425 210.470 117.885 210.930 ;
        RECT 118.435 210.900 118.605 211.165 ;
        RECT 118.145 210.730 118.605 210.900 ;
        RECT 118.775 210.645 119.425 210.995 ;
        RECT 119.595 210.900 119.765 211.165 ;
        RECT 119.935 211.070 120.605 211.400 ;
        RECT 119.595 210.730 120.265 210.900 ;
        RECT 120.435 210.470 120.605 211.070 ;
        RECT 123.155 211.360 123.325 212.115 ;
        RECT 124.235 211.900 124.565 212.605 ;
        RECT 125.875 212.480 126.045 214.135 ;
        RECT 126.215 214.510 127.685 214.680 ;
        RECT 126.215 212.820 126.385 214.510 ;
        RECT 127.855 214.345 128.025 214.930 ;
        RECT 128.195 214.770 128.765 215.100 ;
        RECT 128.935 214.810 131.145 215.210 ;
        RECT 127.855 214.340 128.425 214.345 ;
        RECT 126.555 214.170 128.425 214.340 ;
        RECT 126.555 213.215 126.725 214.170 ;
        RECT 126.895 213.830 127.865 214.000 ;
        RECT 126.895 213.180 127.065 213.830 ;
        RECT 128.060 213.815 128.425 214.170 ;
        RECT 128.595 213.820 128.765 214.770 ;
        RECT 128.935 214.340 129.565 214.620 ;
        RECT 129.395 213.945 129.565 214.340 ;
        RECT 129.735 214.115 130.295 214.810 ;
        RECT 130.465 214.340 131.145 214.620 ;
        RECT 130.465 213.945 130.685 214.340 ;
        RECT 128.085 213.625 128.255 213.630 ;
        RECT 127.265 213.350 128.425 213.625 ;
        RECT 128.595 213.495 129.225 213.820 ;
        RECT 129.395 213.495 130.685 213.945 ;
        RECT 131.315 214.335 131.485 215.610 ;
        RECT 131.785 215.695 133.755 215.865 ;
        RECT 131.785 214.980 131.955 215.695 ;
        RECT 132.125 215.205 133.415 215.525 ;
        RECT 133.085 215.060 133.415 215.205 ;
        RECT 133.585 215.080 133.755 215.695 ;
        RECT 134.035 215.110 134.205 216.140 ;
        RECT 134.375 216.640 134.945 216.645 ;
        RECT 134.375 216.470 136.245 216.640 ;
        RECT 134.375 216.115 134.740 216.470 ;
        RECT 134.935 216.130 135.905 216.300 ;
        RECT 134.545 215.925 134.715 215.930 ;
        RECT 134.375 215.650 135.535 215.925 ;
        RECT 135.735 215.480 135.905 216.130 ;
        RECT 136.075 215.515 136.245 216.470 ;
        RECT 134.375 215.290 135.905 215.480 ;
        RECT 136.415 215.120 136.585 216.810 ;
        RECT 132.155 214.845 132.875 215.035 ;
        RECT 131.655 214.675 131.985 214.755 ;
        RECT 133.585 214.675 133.755 214.910 ;
        RECT 131.655 214.505 133.755 214.675 ;
        RECT 134.035 214.600 134.740 215.110 ;
        RECT 131.315 214.165 132.285 214.335 ;
        RECT 132.545 214.165 132.875 214.335 ;
        RECT 131.315 213.820 131.485 214.165 ;
        RECT 132.545 213.995 132.805 214.165 ;
        RECT 133.055 214.045 133.355 214.505 ;
        RECT 134.035 214.325 134.205 214.600 ;
        RECT 135.015 214.380 135.185 215.090 ;
        RECT 130.855 213.495 131.485 213.820 ;
        RECT 126.895 212.990 128.425 213.180 ;
        RECT 126.215 212.650 127.240 212.820 ;
        RECT 128.595 212.810 128.765 213.495 ;
        RECT 129.675 213.390 130.005 213.495 ;
        RECT 128.935 213.220 129.505 213.325 ;
        RECT 130.175 213.220 131.145 213.325 ;
        RECT 128.935 212.940 131.145 213.220 ;
        RECT 124.770 211.880 125.145 212.435 ;
        RECT 125.875 212.425 126.805 212.480 ;
        RECT 125.375 212.310 126.805 212.425 ;
        RECT 125.375 212.110 126.045 212.310 ;
        RECT 123.540 211.730 124.065 211.860 ;
        RECT 124.770 211.730 125.705 211.880 ;
        RECT 123.540 211.540 125.705 211.730 ;
        RECT 123.540 211.530 124.565 211.540 ;
        RECT 123.155 211.190 123.935 211.360 ;
        RECT 123.155 210.470 123.325 211.190 ;
        RECT 123.545 210.865 124.065 211.020 ;
        RECT 124.235 210.980 124.565 211.530 ;
        RECT 125.875 211.370 126.045 212.110 ;
        RECT 126.395 211.900 126.805 212.075 ;
        RECT 127.050 212.070 127.240 212.650 ;
        RECT 127.615 212.080 127.785 212.790 ;
        RECT 128.060 212.300 128.765 212.810 ;
        RECT 128.935 212.490 131.145 212.770 ;
        RECT 128.935 212.385 129.505 212.490 ;
        RECT 130.175 212.385 131.145 212.490 ;
        RECT 128.595 212.215 128.765 212.300 ;
        RECT 129.675 212.215 130.005 212.320 ;
        RECT 131.315 212.260 131.485 213.495 ;
        RECT 131.760 213.825 132.805 213.995 ;
        RECT 133.025 213.845 133.355 214.045 ;
        RECT 133.535 213.955 134.205 214.325 ;
        RECT 134.410 214.200 135.185 214.380 ;
        RECT 135.560 214.950 136.585 215.120 ;
        RECT 136.755 216.965 136.925 217.150 ;
        RECT 137.095 217.220 139.305 217.390 ;
        RECT 137.095 217.135 138.000 217.220 ;
        RECT 138.730 217.135 139.305 217.220 ;
        RECT 139.475 217.070 140.025 217.400 ;
        RECT 140.195 217.305 140.365 217.570 ;
        RECT 140.535 217.475 141.185 217.825 ;
        RECT 141.355 217.570 142.025 217.740 ;
        RECT 141.355 217.305 141.525 217.570 ;
        RECT 142.195 217.400 143.455 217.830 ;
        RECT 140.195 217.075 141.525 217.305 ;
        RECT 141.695 217.070 143.455 217.400 ;
        RECT 138.235 216.965 138.565 217.050 ;
        RECT 139.475 216.965 139.645 217.070 ;
        RECT 136.755 216.635 137.685 216.965 ;
        RECT 137.855 216.795 138.925 216.965 ;
        RECT 136.755 215.480 136.925 216.635 ;
        RECT 137.855 216.420 138.025 216.795 ;
        RECT 137.095 216.250 138.025 216.420 ;
        RECT 138.205 216.160 138.575 216.515 ;
        RECT 138.755 216.420 138.925 216.795 ;
        RECT 139.095 216.635 139.645 216.965 ;
        RECT 139.905 216.715 142.025 216.900 ;
        RECT 139.475 216.460 139.645 216.635 ;
        RECT 138.755 216.250 139.305 216.420 ;
        RECT 139.475 216.210 140.105 216.460 ;
        RECT 140.275 216.265 141.225 216.545 ;
        RECT 142.195 216.475 143.455 217.070 ;
        RECT 141.735 216.210 143.455 216.475 ;
        RECT 137.095 215.815 139.305 215.985 ;
        RECT 137.095 215.650 138.065 215.815 ;
        RECT 138.735 215.730 139.305 215.815 ;
        RECT 138.235 215.560 138.565 215.645 ;
        RECT 139.475 215.560 139.645 216.210 ;
        RECT 140.235 216.040 141.600 216.095 ;
        RECT 139.925 215.925 142.025 216.040 ;
        RECT 139.925 215.870 140.365 215.925 ;
        RECT 139.925 215.705 140.095 215.870 ;
        RECT 141.470 215.790 142.025 215.925 ;
        RECT 142.195 216.010 143.455 216.210 ;
        RECT 143.625 216.245 145.630 217.830 ;
        RECT 143.625 216.180 146.460 216.245 ;
        RECT 136.755 215.310 138.065 215.480 ;
        RECT 138.235 215.390 138.905 215.560 ;
        RECT 135.560 214.370 135.750 214.950 ;
        RECT 136.755 214.780 136.925 215.310 ;
        RECT 138.235 215.140 138.565 215.165 ;
        RECT 135.995 214.610 136.925 214.780 ;
        RECT 135.995 214.200 136.405 214.375 ;
        RECT 134.410 214.135 136.405 214.200 ;
        RECT 131.760 212.890 131.930 213.825 ;
        RECT 132.100 213.295 132.465 213.655 ;
        RECT 132.635 213.635 132.805 213.825 ;
        RECT 132.635 213.465 133.755 213.635 ;
        RECT 132.100 213.125 133.385 213.295 ;
        RECT 132.400 212.715 132.995 212.955 ;
        RECT 133.165 212.770 133.385 213.125 ;
        RECT 133.585 212.960 133.755 213.465 ;
        RECT 134.035 213.260 134.205 213.955 ;
        RECT 135.015 213.860 136.405 214.135 ;
        RECT 134.465 213.430 134.925 213.600 ;
        RECT 134.035 212.930 134.585 213.260 ;
        RECT 134.755 213.165 134.925 213.430 ;
        RECT 135.095 213.335 135.745 213.685 ;
        RECT 135.915 213.430 136.585 213.600 ;
        RECT 135.915 213.165 136.085 213.430 ;
        RECT 136.755 213.260 136.925 214.610 ;
        RECT 134.755 212.935 136.085 213.165 ;
        RECT 136.255 212.940 136.925 213.260 ;
        RECT 137.095 214.970 138.565 215.140 ;
        RECT 137.095 213.280 137.265 214.970 ;
        RECT 138.735 214.805 138.905 215.390 ;
        RECT 139.075 215.230 139.645 215.560 ;
        RECT 138.735 214.800 139.305 214.805 ;
        RECT 137.435 214.630 139.305 214.800 ;
        RECT 137.435 213.675 137.605 214.630 ;
        RECT 137.775 214.290 138.745 214.460 ;
        RECT 137.775 213.640 137.945 214.290 ;
        RECT 138.940 214.275 139.305 214.630 ;
        RECT 139.475 214.515 139.645 215.230 ;
        RECT 139.925 215.005 140.095 215.510 ;
        RECT 140.295 215.345 140.515 215.700 ;
        RECT 140.685 215.515 141.280 215.755 ;
        RECT 140.295 215.175 141.580 215.345 ;
        RECT 139.925 214.835 141.045 215.005 ;
        RECT 140.875 214.645 141.045 214.835 ;
        RECT 141.215 214.815 141.580 215.175 ;
        RECT 141.750 214.645 141.920 215.580 ;
        RECT 139.475 214.145 140.145 214.515 ;
        RECT 140.325 214.425 140.655 214.625 ;
        RECT 140.875 214.475 141.920 214.645 ;
        RECT 138.965 214.085 139.135 214.090 ;
        RECT 138.145 213.810 139.305 214.085 ;
        RECT 137.775 213.450 139.305 213.640 ;
        RECT 137.095 213.110 138.120 213.280 ;
        RECT 139.475 213.270 139.645 214.145 ;
        RECT 140.325 213.965 140.625 214.425 ;
        RECT 140.875 214.305 141.135 214.475 ;
        RECT 142.195 214.320 143.975 216.010 ;
        RECT 144.145 215.905 146.460 216.180 ;
        RECT 144.145 214.320 145.630 215.905 ;
        RECT 147.200 214.425 147.805 217.830 ;
        RECT 142.195 214.305 142.365 214.320 ;
        RECT 140.805 214.135 141.135 214.305 ;
        RECT 141.395 214.135 142.365 214.305 ;
        RECT 139.925 213.795 142.025 213.965 ;
        RECT 139.925 213.560 140.095 213.795 ;
        RECT 141.695 213.715 142.025 213.795 ;
        RECT 140.805 213.435 141.525 213.625 ;
        RECT 136.255 212.930 137.685 212.940 ;
        RECT 131.655 212.545 132.210 212.680 ;
        RECT 133.585 212.600 133.755 212.765 ;
        RECT 133.315 212.545 133.755 212.600 ;
        RECT 131.655 212.430 133.755 212.545 ;
        RECT 132.080 212.375 133.445 212.430 ;
        RECT 134.035 212.320 134.205 212.930 ;
        RECT 136.755 212.770 137.685 212.930 ;
        RECT 134.465 212.575 136.585 212.760 ;
        RECT 134.035 212.260 134.665 212.320 ;
        RECT 131.315 212.215 131.945 212.260 ;
        RECT 127.615 211.900 128.390 212.080 ;
        RECT 126.395 211.835 128.390 211.900 ;
        RECT 128.595 211.890 129.225 212.215 ;
        RECT 126.395 211.560 127.785 211.835 ;
        RECT 124.865 211.200 126.045 211.370 ;
        RECT 123.545 210.810 124.105 210.865 ;
        RECT 124.735 210.855 125.660 211.030 ;
        RECT 124.685 210.810 125.660 210.855 ;
        RECT 123.545 210.700 125.660 210.810 ;
        RECT 125.875 210.960 126.045 211.200 ;
        RECT 126.215 211.130 126.885 211.300 ;
        RECT 123.545 210.690 124.815 210.700 ;
        RECT 123.980 210.640 124.815 210.690 ;
        RECT 125.875 210.630 126.545 210.960 ;
        RECT 126.715 210.865 126.885 211.130 ;
        RECT 127.055 211.035 127.705 211.385 ;
        RECT 127.875 211.130 128.335 211.300 ;
        RECT 127.875 210.865 128.045 211.130 ;
        RECT 128.595 210.960 128.765 211.890 ;
        RECT 129.395 211.765 130.685 212.215 ;
        RECT 130.855 211.995 131.945 212.215 ;
        RECT 130.855 211.890 131.485 211.995 ;
        RECT 132.455 211.925 133.405 212.205 ;
        RECT 133.575 212.070 134.665 212.260 ;
        RECT 134.835 212.125 135.785 212.405 ;
        RECT 136.755 212.335 136.925 212.770 ;
        RECT 136.295 212.070 136.925 212.335 ;
        RECT 133.575 212.010 134.205 212.070 ;
        RECT 129.395 211.370 129.565 211.765 ;
        RECT 128.935 211.090 129.565 211.370 ;
        RECT 126.715 210.635 128.045 210.865 ;
        RECT 128.215 210.630 128.765 210.960 ;
        RECT 129.735 210.900 130.295 211.595 ;
        RECT 130.465 211.370 130.685 211.765 ;
        RECT 131.315 211.400 131.485 211.890 ;
        RECT 131.655 211.570 133.775 211.755 ;
        RECT 134.035 211.400 134.205 212.010 ;
        RECT 134.795 211.900 136.160 211.955 ;
        RECT 134.485 211.785 136.585 211.900 ;
        RECT 134.485 211.730 134.925 211.785 ;
        RECT 134.485 211.565 134.655 211.730 ;
        RECT 136.030 211.650 136.585 211.785 ;
        RECT 136.755 211.850 136.925 212.070 ;
        RECT 137.275 212.360 137.685 212.535 ;
        RECT 137.930 212.530 138.120 213.110 ;
        RECT 138.495 212.540 138.665 213.250 ;
        RECT 138.940 212.760 139.645 213.270 ;
        RECT 138.495 212.360 139.270 212.540 ;
        RECT 137.275 212.295 139.270 212.360 ;
        RECT 139.475 212.330 139.645 212.760 ;
        RECT 139.925 212.775 140.095 213.390 ;
        RECT 140.265 213.265 140.595 213.410 ;
        RECT 140.265 212.945 141.555 213.265 ;
        RECT 141.725 212.775 141.895 213.490 ;
        RECT 139.925 212.605 141.895 212.775 ;
        RECT 142.195 213.130 142.365 214.135 ;
        RECT 143.425 213.640 144.260 213.690 ;
        RECT 143.425 213.630 144.695 213.640 ;
        RECT 142.580 213.520 144.695 213.630 ;
        RECT 142.580 213.475 143.555 213.520 ;
        RECT 142.580 213.300 143.505 213.475 ;
        RECT 144.135 213.465 144.695 213.520 ;
        RECT 142.195 212.960 143.375 213.130 ;
        RECT 137.275 212.020 138.665 212.295 ;
        RECT 139.475 212.120 140.175 212.330 ;
        RECT 139.475 211.850 139.645 212.120 ;
        RECT 140.555 211.900 140.885 212.605 ;
        RECT 141.090 211.880 141.465 212.435 ;
        RECT 142.195 212.425 142.365 212.960 ;
        RECT 143.675 212.800 144.005 213.350 ;
        RECT 144.175 213.310 144.695 213.465 ;
        RECT 144.915 213.140 145.630 214.320 ;
        RECT 145.950 214.075 147.805 214.425 ;
        RECT 144.305 212.970 145.630 213.140 ;
        RECT 143.675 212.790 144.700 212.800 ;
        RECT 142.535 212.600 144.700 212.790 ;
        RECT 142.535 212.450 143.470 212.600 ;
        RECT 144.175 212.470 144.700 212.600 ;
        RECT 144.915 212.485 145.630 212.970 ;
        RECT 147.200 212.485 147.805 214.075 ;
        RECT 141.695 212.220 142.365 212.425 ;
        RECT 141.695 212.110 142.865 212.220 ;
        RECT 142.195 211.905 142.865 212.110 ;
        RECT 130.465 211.090 131.145 211.370 ;
        RECT 131.315 211.070 131.985 211.400 ;
        RECT 132.155 211.165 133.485 211.395 ;
        RECT 125.875 210.470 126.045 210.630 ;
        RECT 116.425 209.280 119.175 210.470 ;
        RECT 113.385 208.800 116.775 209.110 ;
        RECT 112.275 207.695 112.445 208.800 ;
        RECT 112.615 207.910 113.165 208.080 ;
        RECT 112.275 207.365 112.825 207.695 ;
        RECT 112.995 207.535 113.165 207.910 ;
        RECT 113.345 207.815 113.715 208.170 ;
        RECT 113.895 207.910 114.825 208.080 ;
        RECT 113.895 207.535 114.065 207.910 ;
        RECT 114.995 207.695 116.775 208.800 ;
        RECT 112.995 207.365 114.065 207.535 ;
        RECT 114.235 207.420 116.775 207.695 ;
        RECT 116.945 208.820 119.175 209.280 ;
        RECT 119.345 209.900 120.605 210.470 ;
        RECT 120.775 210.070 121.455 210.355 ;
        RECT 119.345 209.630 121.065 209.900 ;
        RECT 116.945 207.420 118.655 208.820 ;
        RECT 119.345 208.650 120.605 209.630 ;
        RECT 121.235 209.610 121.455 210.070 ;
        RECT 121.625 209.780 122.185 210.470 ;
        RECT 122.355 210.070 122.985 210.355 ;
        RECT 122.355 209.610 122.525 210.070 ;
        RECT 123.155 209.900 124.615 210.470 ;
        RECT 122.695 209.630 124.615 209.900 ;
        RECT 121.235 209.400 122.525 209.610 ;
        RECT 120.775 208.830 122.985 209.230 ;
        RECT 114.235 207.365 115.165 207.420 ;
        RECT 112.275 206.765 112.445 207.365 ;
        RECT 113.355 207.280 113.685 207.365 ;
        RECT 114.995 207.250 115.165 207.365 ;
        RECT 117.715 207.250 118.655 207.420 ;
        RECT 112.615 207.110 113.190 207.195 ;
        RECT 113.920 207.110 114.825 207.195 ;
        RECT 112.615 206.940 114.825 207.110 ;
        RECT 114.995 206.765 116.255 207.250 ;
        RECT 112.275 206.505 113.285 206.765 ;
        RECT 113.845 206.560 116.255 206.765 ;
        RECT 116.425 206.960 118.655 207.250 ;
        RECT 118.825 207.840 120.605 208.650 ;
        RECT 120.775 208.360 121.455 208.640 ;
        RECT 121.235 207.965 121.455 208.360 ;
        RECT 121.625 208.135 122.185 208.830 ;
        RECT 123.155 208.820 124.615 209.630 ;
        RECT 124.785 210.035 126.045 210.470 ;
        RECT 126.215 210.275 128.335 210.460 ;
        RECT 124.785 209.770 126.505 210.035 ;
        RECT 127.015 209.825 127.965 210.105 ;
        RECT 128.595 210.100 128.765 210.630 ;
        RECT 128.935 210.500 131.145 210.900 ;
        RECT 131.315 210.470 131.485 211.070 ;
        RECT 132.155 210.900 132.325 211.165 ;
        RECT 131.655 210.730 132.325 210.900 ;
        RECT 132.495 210.645 133.145 210.995 ;
        RECT 133.315 210.900 133.485 211.165 ;
        RECT 133.655 211.070 134.205 211.400 ;
        RECT 133.315 210.730 133.775 210.900 ;
        RECT 134.035 210.470 134.205 211.070 ;
        RECT 134.485 210.865 134.655 211.370 ;
        RECT 134.855 211.205 135.075 211.560 ;
        RECT 135.245 211.375 135.840 211.615 ;
        RECT 134.855 211.035 136.140 211.205 ;
        RECT 134.485 210.695 135.605 210.865 ;
        RECT 135.435 210.505 135.605 210.695 ;
        RECT 135.775 210.675 136.140 211.035 ;
        RECT 136.310 210.505 136.480 211.440 ;
        RECT 129.395 210.120 130.685 210.330 ;
        RECT 128.595 210.020 129.225 210.100 ;
        RECT 128.135 209.830 129.225 210.020 ;
        RECT 128.135 209.770 128.765 209.830 ;
        RECT 122.355 208.360 122.985 208.640 ;
        RECT 122.355 207.965 122.525 208.360 ;
        RECT 118.825 207.515 121.065 207.840 ;
        RECT 121.235 207.515 122.525 207.965 ;
        RECT 123.155 207.840 124.095 208.820 ;
        RECT 124.785 208.650 126.045 209.770 ;
        RECT 126.640 209.600 128.005 209.655 ;
        RECT 126.215 209.485 128.315 209.600 ;
        RECT 126.215 209.350 126.770 209.485 ;
        RECT 127.875 209.430 128.315 209.485 ;
        RECT 122.695 207.515 124.095 207.840 ;
        RECT 118.825 206.960 120.605 207.515 ;
        RECT 121.915 207.410 122.245 207.515 ;
        RECT 120.775 207.240 121.745 207.345 ;
        RECT 122.415 207.240 122.985 207.345 ;
        RECT 120.775 206.960 122.985 207.240 ;
        RECT 123.155 206.960 124.095 207.515 ;
        RECT 124.265 207.865 126.045 208.650 ;
        RECT 126.320 208.205 126.490 209.140 ;
        RECT 126.960 209.075 127.555 209.315 ;
        RECT 128.145 209.265 128.315 209.430 ;
        RECT 127.725 208.905 127.945 209.260 ;
        RECT 128.595 209.090 128.765 209.770 ;
        RECT 129.395 209.660 129.565 210.120 ;
        RECT 128.935 209.375 129.565 209.660 ;
        RECT 129.735 209.260 130.295 209.950 ;
        RECT 130.465 209.660 130.685 210.120 ;
        RECT 131.315 210.100 132.575 210.470 ;
        RECT 130.855 209.830 132.575 210.100 ;
        RECT 130.465 209.375 131.145 209.660 ;
        RECT 131.315 209.090 132.575 209.830 ;
        RECT 132.745 210.375 134.205 210.470 ;
        RECT 132.745 210.005 134.705 210.375 ;
        RECT 134.885 210.285 135.215 210.485 ;
        RECT 135.435 210.335 136.480 210.505 ;
        RECT 136.755 211.160 138.015 211.850 ;
        RECT 138.185 211.360 139.645 211.850 ;
        RECT 139.860 211.730 140.385 211.860 ;
        RECT 141.090 211.730 142.025 211.880 ;
        RECT 139.860 211.540 142.025 211.730 ;
        RECT 139.860 211.530 140.885 211.540 ;
        RECT 138.185 211.330 140.255 211.360 ;
        RECT 138.725 211.190 140.255 211.330 ;
        RECT 136.755 210.640 138.555 211.160 ;
        RECT 138.725 210.640 139.645 211.190 ;
        RECT 139.865 210.865 140.385 211.020 ;
        RECT 140.555 210.980 140.885 211.530 ;
        RECT 142.195 211.370 142.365 211.905 ;
        RECT 143.095 211.895 143.470 212.450 ;
        RECT 143.675 211.725 144.005 212.430 ;
        RECT 144.915 212.210 145.085 212.485 ;
        RECT 144.385 212.000 145.085 212.210 ;
        RECT 141.185 211.200 142.365 211.370 ;
        RECT 139.865 210.810 140.425 210.865 ;
        RECT 141.055 210.855 141.980 211.030 ;
        RECT 141.005 210.810 141.980 210.855 ;
        RECT 139.865 210.700 141.980 210.810 ;
        RECT 139.865 210.690 141.135 210.700 ;
        RECT 140.300 210.640 141.135 210.690 ;
        RECT 136.755 210.380 136.925 210.640 ;
        RECT 139.475 210.380 139.645 210.640 ;
        RECT 132.745 209.260 134.205 210.005 ;
        RECT 134.885 209.825 135.185 210.285 ;
        RECT 135.435 210.165 135.695 210.335 ;
        RECT 136.755 210.165 137.670 210.380 ;
        RECT 135.365 209.995 135.695 210.165 ;
        RECT 135.955 210.110 137.670 210.165 ;
        RECT 135.955 209.995 136.925 210.110 ;
        RECT 134.485 209.655 136.585 209.825 ;
        RECT 134.485 209.420 134.655 209.655 ;
        RECT 136.255 209.575 136.585 209.655 ;
        RECT 135.365 209.295 136.085 209.485 ;
        RECT 136.755 209.480 136.925 209.995 ;
        RECT 137.840 209.940 138.825 210.380 ;
        RECT 138.995 210.080 139.645 210.380 ;
        RECT 139.815 210.190 142.025 210.470 ;
        RECT 139.815 210.085 140.385 210.190 ;
        RECT 141.055 210.085 142.025 210.190 ;
        RECT 142.195 210.195 142.365 211.200 ;
        RECT 142.665 211.555 144.635 211.725 ;
        RECT 142.665 210.840 142.835 211.555 ;
        RECT 143.005 211.065 144.295 211.385 ;
        RECT 143.965 210.920 144.295 211.065 ;
        RECT 144.465 210.940 144.635 211.555 ;
        RECT 144.915 210.915 145.085 212.000 ;
        RECT 145.255 211.130 145.805 211.300 ;
        RECT 143.035 210.705 143.755 210.895 ;
        RECT 142.535 210.535 142.865 210.615 ;
        RECT 144.465 210.535 144.635 210.770 ;
        RECT 142.535 210.365 144.635 210.535 ;
        RECT 144.915 210.585 145.465 210.915 ;
        RECT 145.635 210.755 145.805 211.130 ;
        RECT 145.985 211.035 146.355 211.390 ;
        RECT 146.535 211.130 147.465 211.300 ;
        RECT 146.535 210.755 146.705 211.130 ;
        RECT 147.635 210.915 147.805 212.485 ;
        RECT 145.635 210.585 146.705 210.755 ;
        RECT 146.875 210.585 147.805 210.915 ;
        RECT 137.100 209.910 138.825 209.940 ;
        RECT 139.475 209.915 139.645 210.080 ;
        RECT 142.195 210.025 143.165 210.195 ;
        RECT 143.425 210.025 143.755 210.195 ;
        RECT 140.555 209.915 140.885 210.020 ;
        RECT 142.195 209.915 142.365 210.025 ;
        RECT 137.100 209.650 139.280 209.910 ;
        RECT 126.660 208.735 127.945 208.905 ;
        RECT 126.660 208.375 127.025 208.735 ;
        RECT 128.145 208.565 128.315 209.070 ;
        RECT 127.195 208.395 128.315 208.565 ;
        RECT 127.195 208.205 127.365 208.395 ;
        RECT 126.320 208.035 127.365 208.205 ;
        RECT 127.105 207.865 127.365 208.035 ;
        RECT 127.585 207.985 127.915 208.185 ;
        RECT 128.595 208.075 130.055 209.090 ;
        RECT 124.265 207.695 126.845 207.865 ;
        RECT 127.105 207.695 127.435 207.865 ;
        RECT 124.265 206.960 126.045 207.695 ;
        RECT 127.615 207.525 127.915 207.985 ;
        RECT 128.095 207.880 130.055 208.075 ;
        RECT 130.225 207.880 133.095 209.090 ;
        RECT 133.265 208.190 134.205 209.260 ;
        RECT 134.485 208.635 134.655 209.250 ;
        RECT 134.825 209.125 135.155 209.270 ;
        RECT 134.825 208.805 136.115 209.125 ;
        RECT 136.285 208.635 136.455 209.350 ;
        RECT 134.485 208.465 136.455 208.635 ;
        RECT 136.755 209.225 137.655 209.480 ;
        RECT 136.755 208.610 136.930 209.225 ;
        RECT 137.840 209.215 138.825 209.650 ;
        RECT 139.475 209.590 140.105 209.915 ;
        RECT 139.475 209.480 139.645 209.590 ;
        RECT 138.995 209.220 139.645 209.480 ;
        RECT 137.840 209.040 138.065 209.215 ;
        RECT 137.100 208.780 138.065 209.040 ;
        RECT 133.265 207.980 134.735 208.190 ;
        RECT 133.265 207.880 134.205 207.980 ;
        RECT 128.095 207.705 129.535 207.880 ;
        RECT 130.225 207.710 131.485 207.880 ;
        RECT 126.215 207.355 128.315 207.525 ;
        RECT 126.215 207.275 126.545 207.355 ;
        RECT 116.425 206.730 117.885 206.960 ;
        RECT 113.845 206.505 116.795 206.560 ;
        RECT 112.275 206.330 112.445 206.505 ;
        RECT 114.995 206.330 116.795 206.505 ;
        RECT 112.275 206.040 113.170 206.330 ;
        RECT 113.830 206.040 116.795 206.330 ;
        RECT 116.965 206.330 117.885 206.730 ;
        RECT 120.435 206.330 120.605 206.960 ;
        RECT 116.965 206.040 118.610 206.330 ;
        RECT 119.270 206.040 120.605 206.330 ;
        RECT 120.955 206.515 122.345 206.790 ;
        RECT 120.955 206.450 122.950 206.515 ;
        RECT 120.955 206.275 121.365 206.450 ;
        RECT 112.275 205.405 112.445 206.040 ;
        RECT 114.995 205.405 115.165 206.040 ;
        RECT 117.715 205.870 117.885 206.040 ;
        RECT 120.435 205.870 121.365 206.040 ;
        RECT 116.225 205.820 117.060 205.870 ;
        RECT 116.225 205.810 117.495 205.820 ;
        RECT 115.380 205.700 117.495 205.810 ;
        RECT 115.380 205.655 116.355 205.700 ;
        RECT 115.380 205.480 116.305 205.655 ;
        RECT 116.935 205.645 117.495 205.700 ;
        RECT 112.275 205.145 113.285 205.405 ;
        RECT 113.845 205.310 115.165 205.405 ;
        RECT 113.845 205.145 116.175 205.310 ;
        RECT 112.275 204.545 112.445 205.145 ;
        RECT 114.995 205.140 116.175 205.145 ;
        RECT 112.615 204.800 114.825 204.970 ;
        RECT 112.615 204.715 113.190 204.800 ;
        RECT 113.920 204.715 114.825 204.800 ;
        RECT 113.355 204.545 113.685 204.630 ;
        RECT 114.995 204.545 115.165 205.140 ;
        RECT 116.475 204.980 116.805 205.530 ;
        RECT 116.975 205.490 117.495 205.645 ;
        RECT 117.715 205.565 118.395 205.870 ;
        RECT 117.715 205.320 117.885 205.565 ;
        RECT 118.565 205.555 119.125 205.870 ;
        RECT 120.435 205.860 120.605 205.870 ;
        RECT 119.625 205.565 120.605 205.860 ;
        RECT 121.610 205.700 121.800 206.280 ;
        RECT 117.105 205.150 117.885 205.320 ;
        RECT 116.475 204.970 117.500 204.980 ;
        RECT 115.335 204.780 117.500 204.970 ;
        RECT 115.335 204.630 116.270 204.780 ;
        RECT 116.975 204.650 117.500 204.780 ;
        RECT 117.715 204.965 117.885 205.150 ;
        RECT 118.065 205.140 120.265 205.385 ;
        RECT 118.065 205.135 119.125 205.140 ;
        RECT 117.715 204.705 118.410 204.965 ;
        RECT 112.275 204.215 112.825 204.545 ;
        RECT 112.995 204.375 114.065 204.545 ;
        RECT 112.275 203.140 112.445 204.215 ;
        RECT 112.995 204.000 113.165 204.375 ;
        RECT 112.615 203.830 113.165 204.000 ;
        RECT 113.345 203.740 113.715 204.095 ;
        RECT 113.895 204.000 114.065 204.375 ;
        RECT 114.235 204.400 115.165 204.545 ;
        RECT 114.235 204.215 115.665 204.400 ;
        RECT 114.995 204.085 115.665 204.215 ;
        RECT 113.895 203.830 114.825 204.000 ;
        RECT 112.705 203.310 113.165 203.480 ;
        RECT 112.275 202.810 112.825 203.140 ;
        RECT 112.995 203.045 113.165 203.310 ;
        RECT 113.335 203.215 113.985 203.565 ;
        RECT 114.155 203.310 114.825 203.480 ;
        RECT 114.155 203.045 114.325 203.310 ;
        RECT 114.995 203.140 115.165 204.085 ;
        RECT 115.895 204.075 116.270 204.630 ;
        RECT 116.475 203.905 116.805 204.610 ;
        RECT 117.715 204.390 117.885 204.705 ;
        RECT 118.875 204.525 119.125 205.135 ;
        RECT 120.435 204.965 120.605 205.565 ;
        RECT 119.625 204.705 120.605 204.965 ;
        RECT 117.185 204.180 117.885 204.390 ;
        RECT 118.065 204.275 120.260 204.525 ;
        RECT 117.715 204.105 117.885 204.180 ;
        RECT 112.995 202.815 114.325 203.045 ;
        RECT 114.495 202.810 115.165 203.140 ;
        RECT 115.465 203.735 117.435 203.905 ;
        RECT 115.465 203.020 115.635 203.735 ;
        RECT 115.805 203.245 117.095 203.565 ;
        RECT 116.765 203.100 117.095 203.245 ;
        RECT 117.265 203.120 117.435 203.735 ;
        RECT 117.715 203.845 118.445 204.105 ;
        RECT 117.715 203.245 117.885 203.845 ;
        RECT 118.080 203.415 118.705 203.675 ;
        RECT 115.835 202.885 116.555 203.075 ;
        RECT 117.715 202.985 118.365 203.245 ;
        RECT 112.275 202.200 112.445 202.810 ;
        RECT 112.705 202.455 114.825 202.640 ;
        RECT 114.995 202.375 115.165 202.810 ;
        RECT 115.335 202.715 115.665 202.795 ;
        RECT 117.265 202.715 117.435 202.950 ;
        RECT 115.335 202.545 117.435 202.715 ;
        RECT 112.275 201.950 112.905 202.200 ;
        RECT 113.075 202.005 114.025 202.285 ;
        RECT 114.995 202.215 115.965 202.375 ;
        RECT 114.535 202.205 115.965 202.215 ;
        RECT 116.225 202.205 116.555 202.375 ;
        RECT 114.535 201.950 115.165 202.205 ;
        RECT 116.225 202.035 116.485 202.205 ;
        RECT 116.735 202.085 117.035 202.545 ;
        RECT 117.715 202.385 117.885 202.985 ;
        RECT 118.535 202.815 118.705 203.415 ;
        RECT 118.080 202.555 118.705 202.815 ;
        RECT 117.715 202.365 118.365 202.385 ;
        RECT 112.275 200.255 112.445 201.950 ;
        RECT 113.035 201.780 114.400 201.835 ;
        RECT 112.725 201.665 114.825 201.780 ;
        RECT 112.725 201.610 113.165 201.665 ;
        RECT 112.725 201.445 112.895 201.610 ;
        RECT 114.270 201.530 114.825 201.665 ;
        RECT 112.725 200.745 112.895 201.250 ;
        RECT 113.095 201.085 113.315 201.440 ;
        RECT 113.485 201.255 114.080 201.495 ;
        RECT 113.095 200.915 114.380 201.085 ;
        RECT 112.725 200.575 113.845 200.745 ;
        RECT 113.675 200.385 113.845 200.575 ;
        RECT 114.015 200.555 114.380 200.915 ;
        RECT 114.550 200.385 114.720 201.320 ;
        RECT 112.275 199.885 112.945 200.255 ;
        RECT 113.125 200.165 113.455 200.365 ;
        RECT 113.675 200.215 114.720 200.385 ;
        RECT 114.995 200.300 115.165 201.950 ;
        RECT 115.440 201.865 116.485 202.035 ;
        RECT 116.705 201.885 117.035 202.085 ;
        RECT 117.215 202.125 118.365 202.365 ;
        RECT 117.215 201.995 117.885 202.125 ;
        RECT 115.440 200.930 115.610 201.865 ;
        RECT 115.780 201.335 116.145 201.695 ;
        RECT 116.315 201.675 116.485 201.865 ;
        RECT 116.315 201.505 117.435 201.675 ;
        RECT 115.780 201.165 117.065 201.335 ;
        RECT 116.080 200.755 116.675 200.995 ;
        RECT 116.845 200.810 117.065 201.165 ;
        RECT 117.265 201.000 117.435 201.505 ;
        RECT 117.715 201.525 117.885 201.995 ;
        RECT 118.535 201.955 118.705 202.555 ;
        RECT 118.080 201.695 118.705 201.955 ;
        RECT 117.715 201.280 118.365 201.525 ;
        RECT 115.335 200.585 115.890 200.720 ;
        RECT 117.265 200.640 117.435 200.805 ;
        RECT 116.995 200.585 117.435 200.640 ;
        RECT 115.335 200.470 117.435 200.585 ;
        RECT 117.715 200.665 117.885 201.280 ;
        RECT 118.535 201.110 118.705 201.695 ;
        RECT 118.080 200.835 118.705 201.110 ;
        RECT 115.760 200.415 117.125 200.470 ;
        RECT 117.715 200.420 118.365 200.665 ;
        RECT 117.715 200.300 117.885 200.420 ;
        RECT 112.275 198.070 112.445 199.885 ;
        RECT 113.125 199.705 113.425 200.165 ;
        RECT 113.675 200.045 113.935 200.215 ;
        RECT 114.995 200.045 115.625 200.300 ;
        RECT 113.605 199.875 113.935 200.045 ;
        RECT 114.195 200.035 115.625 200.045 ;
        RECT 114.195 199.875 115.165 200.035 ;
        RECT 116.135 199.965 117.085 200.245 ;
        RECT 117.255 200.050 117.885 200.300 ;
        RECT 118.535 200.250 118.705 200.835 ;
        RECT 112.725 199.535 114.825 199.705 ;
        RECT 112.725 199.300 112.895 199.535 ;
        RECT 114.495 199.455 114.825 199.535 ;
        RECT 114.995 199.440 115.165 199.875 ;
        RECT 117.715 199.810 117.885 200.050 ;
        RECT 118.080 199.990 118.705 200.250 ;
        RECT 115.335 199.610 117.455 199.795 ;
        RECT 117.715 199.560 118.365 199.810 ;
        RECT 117.715 199.440 117.885 199.560 ;
        RECT 113.605 199.175 114.325 199.365 ;
        RECT 112.725 198.515 112.895 199.130 ;
        RECT 113.065 199.005 113.395 199.150 ;
        RECT 113.065 198.685 114.355 199.005 ;
        RECT 114.525 198.515 114.695 199.230 ;
        RECT 112.725 198.345 114.695 198.515 ;
        RECT 114.995 199.110 115.665 199.440 ;
        RECT 115.835 199.205 117.165 199.435 ;
        RECT 112.275 197.860 112.975 198.070 ;
        RECT 112.275 197.100 112.445 197.860 ;
        RECT 113.355 197.640 113.685 198.345 ;
        RECT 113.890 197.620 114.265 198.175 ;
        RECT 114.995 198.165 115.165 199.110 ;
        RECT 115.835 198.940 116.005 199.205 ;
        RECT 115.335 198.770 116.005 198.940 ;
        RECT 116.175 198.685 116.825 199.035 ;
        RECT 116.995 198.940 117.165 199.205 ;
        RECT 117.335 199.110 117.885 199.440 ;
        RECT 118.535 199.390 118.705 199.990 ;
        RECT 118.080 199.130 118.705 199.390 ;
        RECT 117.715 198.950 117.885 199.110 ;
        RECT 116.995 198.770 117.455 198.940 ;
        RECT 117.715 198.700 118.365 198.950 ;
        RECT 115.335 198.335 117.545 198.505 ;
        RECT 115.335 198.170 116.305 198.335 ;
        RECT 116.975 198.250 117.545 198.335 ;
        RECT 114.495 198.000 115.165 198.165 ;
        RECT 116.475 198.080 116.805 198.165 ;
        RECT 117.715 198.090 117.885 198.700 ;
        RECT 118.535 198.530 118.705 199.130 ;
        RECT 118.080 198.270 118.705 198.530 ;
        RECT 118.535 198.095 118.705 198.270 ;
        RECT 118.875 198.265 119.125 204.275 ;
        RECT 120.435 204.105 120.605 204.705 ;
        RECT 119.635 203.845 120.605 204.105 ;
        RECT 119.295 203.415 120.260 203.675 ;
        RECT 120.430 203.500 120.605 203.845 ;
        RECT 120.775 205.530 121.800 205.700 ;
        RECT 122.175 206.270 122.950 206.450 ;
        RECT 123.155 206.330 123.325 206.960 ;
        RECT 125.875 206.330 126.045 206.960 ;
        RECT 122.175 205.560 122.345 206.270 ;
        RECT 123.155 206.050 124.050 206.330 ;
        RECT 122.620 206.040 124.050 206.050 ;
        RECT 124.710 206.040 126.045 206.330 ;
        RECT 126.345 206.335 126.515 207.050 ;
        RECT 126.715 206.995 127.435 207.185 ;
        RECT 128.145 207.120 128.315 207.355 ;
        RECT 127.645 206.825 127.975 206.970 ;
        RECT 126.685 206.505 127.975 206.825 ;
        RECT 128.145 206.335 128.315 206.950 ;
        RECT 126.345 206.165 128.315 206.335 ;
        RECT 128.595 206.500 129.535 207.705 ;
        RECT 129.705 207.240 131.485 207.710 ;
        RECT 134.035 207.250 134.205 207.880 ;
        RECT 135.115 207.760 135.445 208.465 ;
        RECT 136.755 208.365 137.655 208.610 ;
        RECT 135.650 207.740 136.025 208.295 ;
        RECT 136.755 208.285 136.930 208.365 ;
        RECT 136.255 207.970 136.930 208.285 ;
        RECT 137.825 208.180 138.065 208.780 ;
        RECT 136.755 207.750 136.930 207.970 ;
        RECT 137.100 207.920 138.065 208.180 ;
        RECT 134.420 207.590 134.945 207.720 ;
        RECT 135.650 207.590 136.585 207.740 ;
        RECT 134.420 207.400 136.585 207.590 ;
        RECT 136.755 207.505 137.655 207.750 ;
        RECT 134.420 207.390 135.445 207.400 ;
        RECT 129.705 206.945 132.295 207.240 ;
        RECT 129.705 206.500 131.485 206.945 ;
        RECT 132.795 206.935 133.355 207.250 ;
        RECT 133.525 207.220 134.205 207.250 ;
        RECT 133.525 207.050 134.815 207.220 ;
        RECT 133.525 206.945 134.205 207.050 ;
        RECT 131.655 206.520 133.855 206.765 ;
        RECT 128.595 206.330 128.765 206.500 ;
        RECT 131.315 206.345 131.485 206.500 ;
        RECT 132.795 206.515 133.855 206.520 ;
        RECT 131.315 206.330 132.295 206.345 ;
        RECT 122.620 205.540 123.325 206.040 ;
        RECT 125.875 205.985 126.045 206.040 ;
        RECT 123.585 205.610 124.045 205.780 ;
        RECT 120.775 203.840 120.945 205.530 ;
        RECT 123.155 205.440 123.325 205.540 ;
        RECT 121.455 205.170 122.985 205.360 ;
        RECT 121.115 204.180 121.285 205.135 ;
        RECT 121.455 204.520 121.625 205.170 ;
        RECT 123.155 205.110 123.705 205.440 ;
        RECT 123.875 205.345 124.045 205.610 ;
        RECT 124.215 205.515 124.865 205.865 ;
        RECT 125.035 205.610 125.705 205.780 ;
        RECT 125.875 205.670 126.545 205.985 ;
        RECT 125.035 205.345 125.205 205.610 ;
        RECT 125.875 205.440 126.045 205.670 ;
        RECT 126.775 205.440 127.150 205.995 ;
        RECT 127.355 205.460 127.685 206.165 ;
        RECT 128.595 206.040 129.490 206.330 ;
        RECT 130.150 206.085 132.295 206.330 ;
        RECT 130.150 206.040 131.485 206.085 ;
        RECT 128.595 205.890 128.765 206.040 ;
        RECT 128.065 205.860 128.765 205.890 ;
        RECT 128.065 205.680 129.575 205.860 ;
        RECT 128.595 205.590 129.575 205.680 ;
        RECT 123.875 205.115 125.205 205.345 ;
        RECT 125.375 205.110 126.045 205.440 ;
        RECT 121.825 204.725 122.985 205.000 ;
        RECT 121.965 204.720 122.135 204.725 ;
        RECT 121.455 204.350 122.425 204.520 ;
        RECT 122.620 204.180 122.985 204.535 ;
        RECT 121.115 204.010 122.985 204.180 ;
        RECT 122.415 204.005 122.985 204.010 ;
        RECT 123.155 204.500 123.325 205.110 ;
        RECT 123.585 204.755 125.705 204.940 ;
        RECT 125.875 204.930 126.045 205.110 ;
        RECT 126.215 205.290 127.150 205.440 ;
        RECT 127.855 205.290 128.380 205.420 ;
        RECT 126.215 205.100 128.380 205.290 ;
        RECT 127.355 205.090 128.380 205.100 ;
        RECT 125.875 204.760 127.055 204.930 ;
        RECT 123.155 204.250 123.785 204.500 ;
        RECT 123.955 204.305 124.905 204.585 ;
        RECT 125.875 204.515 126.045 204.760 ;
        RECT 125.415 204.250 126.045 204.515 ;
        RECT 126.260 204.415 127.185 204.590 ;
        RECT 127.355 204.540 127.685 205.090 ;
        RECT 128.595 204.920 128.765 205.590 ;
        RECT 129.755 205.520 130.005 205.870 ;
        RECT 131.315 205.860 131.485 206.040 ;
        RECT 132.795 205.905 133.045 206.515 ;
        RECT 134.035 206.345 134.205 206.945 ;
        RECT 134.425 206.725 134.945 206.880 ;
        RECT 135.115 206.840 135.445 207.390 ;
        RECT 136.755 207.230 136.930 207.505 ;
        RECT 137.825 207.320 138.065 207.920 ;
        RECT 135.745 207.060 136.930 207.230 ;
        RECT 137.100 207.060 138.065 207.320 ;
        RECT 136.755 206.890 136.930 207.060 ;
        RECT 134.425 206.670 134.985 206.725 ;
        RECT 135.615 206.715 136.540 206.890 ;
        RECT 135.565 206.670 136.540 206.715 ;
        RECT 134.425 206.560 136.540 206.670 ;
        RECT 136.755 206.645 137.655 206.890 ;
        RECT 134.425 206.550 135.695 206.560 ;
        RECT 134.860 206.500 135.695 206.550 ;
        RECT 133.510 206.330 134.205 206.345 ;
        RECT 136.755 206.330 136.930 206.645 ;
        RECT 137.825 206.475 138.065 207.060 ;
        RECT 133.510 206.085 134.930 206.330 ;
        RECT 134.035 206.040 134.930 206.085 ;
        RECT 135.590 206.045 136.930 206.330 ;
        RECT 137.100 206.215 138.065 206.475 ;
        RECT 135.590 206.040 137.655 206.045 ;
        RECT 130.175 205.530 131.485 205.860 ;
        RECT 131.660 205.655 133.855 205.905 ;
        RECT 131.315 205.485 131.485 205.530 ;
        RECT 128.935 205.350 129.575 205.420 ;
        RECT 128.935 205.180 130.345 205.350 ;
        RECT 128.935 205.090 129.575 205.180 ;
        RECT 127.985 204.750 129.575 204.920 ;
        RECT 128.595 204.680 129.575 204.750 ;
        RECT 127.855 204.425 128.375 204.580 ;
        RECT 126.260 204.370 127.235 204.415 ;
        RECT 127.815 204.370 128.375 204.425 ;
        RECT 126.260 204.260 128.375 204.370 ;
        RECT 120.775 203.670 122.245 203.840 ;
        RECT 121.915 203.645 122.245 203.670 ;
        RECT 119.295 202.815 119.535 203.415 ;
        RECT 120.430 203.330 121.745 203.500 ;
        RECT 122.415 203.420 122.585 204.005 ;
        RECT 123.155 203.580 123.325 204.250 ;
        RECT 123.915 204.080 125.280 204.135 ;
        RECT 123.605 203.965 125.705 204.080 ;
        RECT 123.605 203.910 124.045 203.965 ;
        RECT 123.605 203.745 123.775 203.910 ;
        RECT 125.150 203.830 125.705 203.965 ;
        RECT 120.430 203.245 120.605 203.330 ;
        RECT 119.705 202.985 120.605 203.245 ;
        RECT 121.915 203.250 122.585 203.420 ;
        RECT 122.755 203.250 123.325 203.580 ;
        RECT 121.915 203.165 122.245 203.250 ;
        RECT 119.295 202.555 120.260 202.815 ;
        RECT 120.430 202.650 120.605 202.985 ;
        RECT 120.775 202.995 121.745 203.160 ;
        RECT 122.415 202.995 122.985 203.080 ;
        RECT 120.775 202.825 122.985 202.995 ;
        RECT 123.155 202.650 123.325 203.250 ;
        RECT 123.605 203.045 123.775 203.550 ;
        RECT 123.975 203.385 124.195 203.740 ;
        RECT 124.365 203.555 124.960 203.795 ;
        RECT 123.975 203.215 125.260 203.385 ;
        RECT 123.605 202.875 124.725 203.045 ;
        RECT 124.555 202.685 124.725 202.875 ;
        RECT 124.895 202.855 125.260 203.215 ;
        RECT 125.430 202.685 125.600 203.620 ;
        RECT 119.295 201.955 119.535 202.555 ;
        RECT 120.430 202.385 121.695 202.650 ;
        RECT 119.705 202.125 121.695 202.385 ;
        RECT 119.295 201.695 120.260 201.955 ;
        RECT 120.430 201.730 121.695 202.125 ;
        RECT 121.865 202.555 123.325 202.650 ;
        RECT 121.865 202.185 123.825 202.555 ;
        RECT 124.005 202.465 124.335 202.665 ;
        RECT 124.555 202.515 125.600 202.685 ;
        RECT 125.875 203.520 126.045 204.250 ;
        RECT 127.105 204.250 128.375 204.260 ;
        RECT 127.105 204.200 127.940 204.250 ;
        RECT 126.215 203.855 128.425 204.025 ;
        RECT 126.215 203.690 127.185 203.855 ;
        RECT 127.855 203.770 128.425 203.855 ;
        RECT 128.595 203.890 128.765 204.680 ;
        RECT 129.755 204.660 130.005 205.010 ;
        RECT 130.175 205.000 130.345 205.180 ;
        RECT 131.315 205.225 132.285 205.485 ;
        RECT 130.175 204.670 131.130 205.000 ;
        RECT 131.315 204.625 131.490 205.225 ;
        RECT 131.660 204.795 132.625 205.055 ;
        RECT 128.935 204.060 129.585 204.390 ;
        RECT 127.355 203.600 127.685 203.685 ;
        RECT 128.595 203.600 129.225 203.890 ;
        RECT 125.875 203.350 127.185 203.520 ;
        RECT 127.355 203.430 128.025 203.600 ;
        RECT 121.865 201.900 123.325 202.185 ;
        RECT 124.005 202.005 124.305 202.465 ;
        RECT 124.555 202.345 124.815 202.515 ;
        RECT 125.875 202.345 126.045 203.350 ;
        RECT 127.355 203.180 127.685 203.205 ;
        RECT 124.485 202.175 124.815 202.345 ;
        RECT 125.075 202.175 126.045 202.345 ;
        RECT 119.295 201.095 119.535 201.695 ;
        RECT 120.430 201.525 122.215 201.730 ;
        RECT 119.705 201.265 122.215 201.525 ;
        RECT 119.295 200.835 120.260 201.095 ;
        RECT 120.430 200.980 122.215 201.265 ;
        RECT 122.385 200.980 123.325 201.900 ;
        RECT 123.605 201.835 125.705 202.005 ;
        RECT 123.605 201.600 123.775 201.835 ;
        RECT 125.375 201.755 125.705 201.835 ;
        RECT 124.485 201.475 125.205 201.665 ;
        RECT 119.295 200.250 119.535 200.835 ;
        RECT 120.430 200.665 120.605 200.980 ;
        RECT 119.705 200.420 120.605 200.665 ;
        RECT 120.775 200.550 121.445 200.720 ;
        RECT 120.430 200.380 120.605 200.420 ;
        RECT 119.295 199.990 120.260 200.250 ;
        RECT 120.430 200.050 121.105 200.380 ;
        RECT 121.275 200.285 121.445 200.550 ;
        RECT 121.615 200.455 122.265 200.805 ;
        RECT 122.435 200.550 122.895 200.720 ;
        RECT 122.435 200.285 122.605 200.550 ;
        RECT 123.155 200.380 123.325 200.980 ;
        RECT 123.605 200.815 123.775 201.430 ;
        RECT 123.945 201.305 124.275 201.450 ;
        RECT 123.945 200.985 125.235 201.305 ;
        RECT 125.405 200.815 125.575 201.530 ;
        RECT 123.605 200.645 125.575 200.815 ;
        RECT 125.875 200.980 126.045 202.175 ;
        RECT 126.215 203.010 127.685 203.180 ;
        RECT 126.215 201.320 126.385 203.010 ;
        RECT 127.855 202.845 128.025 203.430 ;
        RECT 128.195 203.560 129.225 203.600 ;
        RECT 128.195 203.270 128.765 203.560 ;
        RECT 129.415 203.345 129.585 204.060 ;
        RECT 129.755 203.920 130.005 204.430 ;
        RECT 131.315 204.370 132.215 204.625 ;
        RECT 130.195 204.365 132.215 204.370 ;
        RECT 130.195 204.040 131.490 204.365 ;
        RECT 132.385 204.195 132.625 204.795 ;
        RECT 131.315 203.765 131.490 204.040 ;
        RECT 131.660 203.935 132.625 204.195 ;
        RECT 127.855 202.840 128.425 202.845 ;
        RECT 126.555 202.670 128.425 202.840 ;
        RECT 126.555 201.715 126.725 202.670 ;
        RECT 126.895 202.330 127.865 202.500 ;
        RECT 126.895 201.680 127.065 202.330 ;
        RECT 128.060 202.315 128.425 202.670 ;
        RECT 128.595 202.815 128.765 203.270 ;
        RECT 128.935 203.015 129.585 203.345 ;
        RECT 129.755 203.340 131.070 203.710 ;
        RECT 131.315 203.505 132.215 203.765 ;
        RECT 128.595 202.485 129.225 202.815 ;
        RECT 127.405 202.125 127.575 202.130 ;
        RECT 127.265 201.850 128.425 202.125 ;
        RECT 126.895 201.490 128.425 201.680 ;
        RECT 128.595 201.320 128.765 202.485 ;
        RECT 129.415 202.260 129.585 203.015 ;
        RECT 129.755 202.840 131.070 203.170 ;
        RECT 131.315 202.905 131.490 203.505 ;
        RECT 132.385 203.335 132.625 203.935 ;
        RECT 131.660 203.075 132.625 203.335 ;
        RECT 131.315 202.645 132.215 202.905 ;
        RECT 129.755 202.300 131.070 202.630 ;
        RECT 129.095 202.090 129.585 202.260 ;
        RECT 128.950 201.590 129.585 201.920 ;
        RECT 129.755 201.710 129.965 202.130 ;
        RECT 131.315 202.045 131.490 202.645 ;
        RECT 132.385 202.475 132.625 203.075 ;
        RECT 131.660 202.215 132.625 202.475 ;
        RECT 130.135 201.780 131.145 202.030 ;
        RECT 131.315 201.800 132.215 202.045 ;
        RECT 129.395 201.540 129.585 201.590 ;
        RECT 130.135 201.540 130.425 201.780 ;
        RECT 131.315 201.610 131.490 201.800 ;
        RECT 132.385 201.630 132.625 202.215 ;
        RECT 126.215 201.150 127.240 201.320 ;
        RECT 128.595 201.310 129.225 201.320 ;
        RECT 125.875 200.810 126.805 200.980 ;
        RECT 121.275 200.055 122.605 200.285 ;
        RECT 122.775 200.370 123.325 200.380 ;
        RECT 122.775 200.160 123.855 200.370 ;
        RECT 122.775 200.050 123.325 200.160 ;
        RECT 119.295 199.390 119.535 199.990 ;
        RECT 120.430 199.805 120.605 200.050 ;
        RECT 119.705 199.560 120.605 199.805 ;
        RECT 120.775 199.695 122.895 199.880 ;
        RECT 120.430 199.455 120.605 199.560 ;
        RECT 119.295 199.130 120.260 199.390 ;
        RECT 120.430 199.190 121.065 199.455 ;
        RECT 121.575 199.245 122.525 199.525 ;
        RECT 123.155 199.440 123.325 200.050 ;
        RECT 124.235 199.940 124.565 200.645 ;
        RECT 124.770 199.920 125.145 200.475 ;
        RECT 125.875 200.465 126.045 200.810 ;
        RECT 125.375 200.150 126.045 200.465 ;
        RECT 123.540 199.770 124.065 199.900 ;
        RECT 124.770 199.770 125.705 199.920 ;
        RECT 123.540 199.580 125.705 199.770 ;
        RECT 123.540 199.570 124.565 199.580 ;
        RECT 122.695 199.400 123.325 199.440 ;
        RECT 122.695 199.230 123.935 199.400 ;
        RECT 122.695 199.190 123.325 199.230 ;
        RECT 119.295 198.530 119.535 199.130 ;
        RECT 120.430 198.945 120.605 199.190 ;
        RECT 121.200 199.020 122.565 199.075 ;
        RECT 119.705 198.700 120.605 198.945 ;
        RECT 120.775 198.905 122.875 199.020 ;
        RECT 120.775 198.770 121.330 198.905 ;
        RECT 122.435 198.850 122.875 198.905 ;
        RECT 119.295 198.270 120.260 198.530 ;
        RECT 119.295 198.095 119.520 198.270 ;
        RECT 117.715 198.080 118.365 198.090 ;
        RECT 114.495 197.850 116.305 198.000 ;
        RECT 116.475 197.910 117.145 198.080 ;
        RECT 114.995 197.830 116.305 197.850 ;
        RECT 112.660 197.470 113.185 197.600 ;
        RECT 113.890 197.470 114.825 197.620 ;
        RECT 112.660 197.280 114.825 197.470 ;
        RECT 112.660 197.270 113.685 197.280 ;
        RECT 112.275 196.930 113.055 197.100 ;
        RECT 112.275 196.205 112.445 196.930 ;
        RECT 112.665 196.605 113.185 196.760 ;
        RECT 113.355 196.720 113.685 197.270 ;
        RECT 114.995 197.110 115.165 197.830 ;
        RECT 116.475 197.660 116.805 197.685 ;
        RECT 113.985 196.940 115.165 197.110 ;
        RECT 112.665 196.550 113.225 196.605 ;
        RECT 113.855 196.595 114.780 196.770 ;
        RECT 113.805 196.550 114.780 196.595 ;
        RECT 112.665 196.440 114.780 196.550 ;
        RECT 112.665 196.430 113.935 196.440 ;
        RECT 113.100 196.380 113.935 196.430 ;
        RECT 114.995 196.205 115.165 196.940 ;
        RECT 112.275 195.945 113.285 196.205 ;
        RECT 113.845 195.945 115.165 196.205 ;
        RECT 112.275 195.345 112.445 195.945 ;
        RECT 112.615 195.600 114.825 195.770 ;
        RECT 112.615 195.515 113.190 195.600 ;
        RECT 113.920 195.515 114.825 195.600 ;
        RECT 114.995 195.460 115.165 195.945 ;
        RECT 115.335 197.490 116.805 197.660 ;
        RECT 115.335 195.800 115.505 197.490 ;
        RECT 116.975 197.325 117.145 197.910 ;
        RECT 117.315 197.830 118.365 198.080 ;
        RECT 117.315 197.750 117.885 197.830 ;
        RECT 116.975 197.320 117.545 197.325 ;
        RECT 115.675 197.150 117.545 197.320 ;
        RECT 115.675 196.195 115.845 197.150 ;
        RECT 116.015 196.810 116.985 196.980 ;
        RECT 116.015 196.160 116.185 196.810 ;
        RECT 117.180 196.795 117.545 197.150 ;
        RECT 117.715 197.230 117.885 197.750 ;
        RECT 118.535 197.660 119.520 198.095 ;
        RECT 120.430 198.085 120.605 198.700 ;
        RECT 119.705 197.830 120.605 198.085 ;
        RECT 118.080 197.400 120.260 197.660 ;
        RECT 118.535 197.370 120.260 197.400 ;
        RECT 117.715 196.930 118.365 197.230 ;
        RECT 118.535 196.930 119.520 197.370 ;
        RECT 120.435 197.285 120.605 197.830 ;
        RECT 120.880 197.625 121.050 198.560 ;
        RECT 121.520 198.495 122.115 198.735 ;
        RECT 122.705 198.685 122.875 198.850 ;
        RECT 122.285 198.325 122.505 198.680 ;
        RECT 123.155 198.500 123.325 199.190 ;
        RECT 123.545 198.905 124.065 199.060 ;
        RECT 124.235 199.020 124.565 199.570 ;
        RECT 125.875 199.410 126.045 200.150 ;
        RECT 126.395 200.400 126.805 200.575 ;
        RECT 127.050 200.570 127.240 201.150 ;
        RECT 127.615 200.580 127.785 201.290 ;
        RECT 128.060 201.150 129.225 201.310 ;
        RECT 129.395 201.280 130.425 201.540 ;
        RECT 130.595 201.280 131.490 201.610 ;
        RECT 131.660 201.370 132.625 201.630 ;
        RECT 129.395 201.170 129.965 201.280 ;
        RECT 128.060 200.800 128.765 201.150 ;
        RECT 129.755 200.960 129.965 201.170 ;
        RECT 131.315 201.185 131.490 201.280 ;
        RECT 127.615 200.400 128.390 200.580 ;
        RECT 126.395 200.335 128.390 200.400 ;
        RECT 126.395 200.060 127.785 200.335 ;
        RECT 126.215 199.610 128.425 199.890 ;
        RECT 126.215 199.505 127.185 199.610 ;
        RECT 127.855 199.505 128.425 199.610 ;
        RECT 128.595 199.795 128.765 200.800 ;
        RECT 128.935 200.790 129.565 200.860 ;
        RECT 130.135 200.790 131.145 201.045 ;
        RECT 128.935 200.520 131.145 200.790 ;
        RECT 131.315 200.940 132.215 201.185 ;
        RECT 128.935 200.070 131.145 200.350 ;
        RECT 128.935 199.965 129.505 200.070 ;
        RECT 130.175 199.965 131.145 200.070 ;
        RECT 131.315 200.325 131.490 200.940 ;
        RECT 132.385 200.770 132.625 201.370 ;
        RECT 131.660 200.510 132.625 200.770 ;
        RECT 131.315 200.080 132.215 200.325 ;
        RECT 129.675 199.795 130.005 199.900 ;
        RECT 131.315 199.795 131.490 200.080 ;
        RECT 132.385 199.910 132.625 200.510 ;
        RECT 128.595 199.470 129.225 199.795 ;
        RECT 124.865 199.335 126.045 199.410 ;
        RECT 127.355 199.335 127.685 199.440 ;
        RECT 128.595 199.335 128.765 199.470 ;
        RECT 124.865 199.240 126.505 199.335 ;
        RECT 123.545 198.850 124.105 198.905 ;
        RECT 124.735 198.895 125.660 199.070 ;
        RECT 124.685 198.850 125.660 198.895 ;
        RECT 123.545 198.740 125.660 198.850 ;
        RECT 125.875 199.010 126.505 199.240 ;
        RECT 123.545 198.730 124.815 198.740 ;
        RECT 123.980 198.680 124.815 198.730 ;
        RECT 121.220 198.155 122.505 198.325 ;
        RECT 121.220 197.795 121.585 198.155 ;
        RECT 122.705 197.985 122.875 198.490 ;
        RECT 121.755 197.815 122.875 197.985 ;
        RECT 123.155 198.170 123.830 198.500 ;
        RECT 124.685 198.445 124.855 198.450 ;
        RECT 121.755 197.625 121.925 197.815 ;
        RECT 120.880 197.455 121.925 197.625 ;
        RECT 121.665 197.285 121.925 197.455 ;
        RECT 122.145 197.405 122.475 197.605 ;
        RECT 123.155 197.495 123.325 198.170 ;
        RECT 124.005 198.145 124.855 198.445 ;
        RECT 125.025 198.250 125.685 198.420 ;
        RECT 123.520 197.975 123.895 198.000 ;
        RECT 125.025 197.975 125.255 198.250 ;
        RECT 125.875 198.080 126.045 199.010 ;
        RECT 126.675 198.885 127.965 199.335 ;
        RECT 128.135 199.010 128.765 199.335 ;
        RECT 126.675 198.490 126.895 198.885 ;
        RECT 126.215 198.210 126.895 198.490 ;
        RECT 123.520 197.760 125.255 197.975 ;
        RECT 120.435 197.200 121.405 197.285 ;
        RECT 119.690 197.115 121.405 197.200 ;
        RECT 121.665 197.115 121.995 197.285 ;
        RECT 119.690 196.930 120.605 197.115 ;
        RECT 122.175 196.945 122.475 197.405 ;
        RECT 122.655 197.125 123.325 197.495 ;
        RECT 124.045 197.740 125.255 197.760 ;
        RECT 125.425 197.750 126.045 198.080 ;
        RECT 127.065 198.020 127.625 198.715 ;
        RECT 127.795 198.490 127.965 198.885 ;
        RECT 127.795 198.210 128.425 198.490 ;
        RECT 123.510 197.310 123.850 197.480 ;
        RECT 124.045 197.420 124.375 197.740 ;
        RECT 117.715 196.670 117.885 196.930 ;
        RECT 120.435 196.670 120.605 196.930 ;
        RECT 120.775 196.775 122.875 196.945 ;
        RECT 120.775 196.695 121.105 196.775 ;
        RECT 116.525 196.605 116.695 196.610 ;
        RECT 116.385 196.330 117.545 196.605 ;
        RECT 116.015 195.970 117.545 196.160 ;
        RECT 117.715 196.150 119.175 196.670 ;
        RECT 115.335 195.630 116.360 195.800 ;
        RECT 117.715 195.790 118.635 196.150 ;
        RECT 119.345 195.980 120.605 196.670 ;
        RECT 113.355 195.345 113.685 195.430 ;
        RECT 114.995 195.345 115.925 195.460 ;
        RECT 112.275 195.015 112.825 195.345 ;
        RECT 112.995 195.175 114.065 195.345 ;
        RECT 112.275 193.450 112.445 195.015 ;
        RECT 112.995 194.800 113.165 195.175 ;
        RECT 112.615 194.630 113.165 194.800 ;
        RECT 113.345 194.540 113.715 194.895 ;
        RECT 113.895 194.800 114.065 195.175 ;
        RECT 114.235 195.290 115.925 195.345 ;
        RECT 114.235 195.015 115.165 195.290 ;
        RECT 113.895 194.630 114.825 194.800 ;
        RECT 114.995 193.450 115.165 195.015 ;
        RECT 115.515 194.880 115.925 195.055 ;
        RECT 116.170 195.050 116.360 195.630 ;
        RECT 116.735 195.060 116.905 195.770 ;
        RECT 117.180 195.460 118.635 195.790 ;
        RECT 118.805 195.460 120.605 195.980 ;
        RECT 120.905 195.755 121.075 196.470 ;
        RECT 121.275 196.415 121.995 196.605 ;
        RECT 122.705 196.540 122.875 196.775 ;
        RECT 123.155 196.720 123.325 197.125 ;
        RECT 123.655 197.250 123.850 197.310 ;
        RECT 124.545 197.265 125.660 197.550 ;
        RECT 124.545 197.250 124.715 197.265 ;
        RECT 123.655 197.080 124.715 197.250 ;
        RECT 125.875 197.220 126.045 197.750 ;
        RECT 126.215 197.620 128.425 198.020 ;
        RECT 128.595 197.680 128.765 199.010 ;
        RECT 129.395 199.345 130.685 199.795 ;
        RECT 130.855 199.470 131.490 199.795 ;
        RECT 131.660 199.650 132.625 199.910 ;
        RECT 129.395 198.950 129.565 199.345 ;
        RECT 128.935 198.670 129.565 198.950 ;
        RECT 129.735 198.480 130.295 199.175 ;
        RECT 130.465 198.950 130.685 199.345 ;
        RECT 131.315 199.465 131.490 199.470 ;
        RECT 132.400 199.475 132.625 199.650 ;
        RECT 132.795 199.645 133.045 205.655 ;
        RECT 134.035 205.485 134.205 206.040 ;
        RECT 134.465 205.610 134.925 205.780 ;
        RECT 133.475 205.440 134.205 205.485 ;
        RECT 133.475 205.225 134.585 205.440 ;
        RECT 134.035 205.110 134.585 205.225 ;
        RECT 134.755 205.345 134.925 205.610 ;
        RECT 135.095 205.515 135.745 205.865 ;
        RECT 136.755 205.785 137.655 206.040 ;
        RECT 135.915 205.610 136.585 205.780 ;
        RECT 135.915 205.345 136.085 205.610 ;
        RECT 136.755 205.440 136.930 205.785 ;
        RECT 137.825 205.615 138.065 206.215 ;
        RECT 134.755 205.115 136.085 205.345 ;
        RECT 136.255 205.185 136.930 205.440 ;
        RECT 137.100 205.355 138.065 205.615 ;
        RECT 136.255 205.110 137.655 205.185 ;
        RECT 133.215 204.795 133.840 205.055 ;
        RECT 133.215 204.195 133.385 204.795 ;
        RECT 134.035 204.625 134.205 205.110 ;
        RECT 134.465 204.755 136.585 204.940 ;
        RECT 136.755 204.925 137.655 205.110 ;
        RECT 133.555 204.500 134.205 204.625 ;
        RECT 133.555 204.365 134.665 204.500 ;
        RECT 134.035 204.250 134.665 204.365 ;
        RECT 134.835 204.305 135.785 204.585 ;
        RECT 136.755 204.515 136.930 204.925 ;
        RECT 137.825 204.755 138.065 205.355 ;
        RECT 136.295 204.325 136.930 204.515 ;
        RECT 137.100 204.495 138.065 204.755 ;
        RECT 136.295 204.250 137.655 204.325 ;
        RECT 133.215 203.935 133.840 204.195 ;
        RECT 133.215 203.335 133.385 203.935 ;
        RECT 134.035 203.765 134.205 204.250 ;
        RECT 134.795 204.080 136.160 204.135 ;
        RECT 133.555 203.505 134.205 203.765 ;
        RECT 134.485 203.965 136.585 204.080 ;
        RECT 134.485 203.910 134.925 203.965 ;
        RECT 134.485 203.745 134.655 203.910 ;
        RECT 136.030 203.830 136.585 203.965 ;
        RECT 136.755 204.065 137.655 204.250 ;
        RECT 133.215 203.075 133.840 203.335 ;
        RECT 133.215 202.490 133.385 203.075 ;
        RECT 134.035 202.905 134.205 203.505 ;
        RECT 133.555 202.660 134.205 202.905 ;
        RECT 134.485 203.045 134.655 203.550 ;
        RECT 134.855 203.385 135.075 203.740 ;
        RECT 135.245 203.555 135.840 203.795 ;
        RECT 134.855 203.215 136.140 203.385 ;
        RECT 134.485 202.875 135.605 203.045 ;
        RECT 135.435 202.685 135.605 202.875 ;
        RECT 135.775 202.855 136.140 203.215 ;
        RECT 136.310 202.685 136.480 203.620 ;
        RECT 134.035 202.555 134.205 202.660 ;
        RECT 133.215 202.215 133.840 202.490 ;
        RECT 133.215 201.630 133.385 202.215 ;
        RECT 134.035 202.185 134.705 202.555 ;
        RECT 134.885 202.465 135.215 202.665 ;
        RECT 135.435 202.515 136.480 202.685 ;
        RECT 136.755 203.465 136.930 204.065 ;
        RECT 137.825 203.895 138.065 204.495 ;
        RECT 137.100 203.635 138.065 203.895 ;
        RECT 136.755 203.205 137.725 203.465 ;
        RECT 136.755 202.605 136.925 203.205 ;
        RECT 138.235 203.035 138.485 209.045 ;
        RECT 138.655 209.040 138.825 209.215 ;
        RECT 138.655 208.780 139.280 209.040 ;
        RECT 138.655 208.180 138.825 208.780 ;
        RECT 139.475 208.610 139.645 209.220 ;
        RECT 140.275 209.465 141.565 209.915 ;
        RECT 141.735 209.590 142.365 209.915 ;
        RECT 143.425 209.855 143.685 210.025 ;
        RECT 143.935 209.905 144.235 210.365 ;
        RECT 144.915 210.185 145.085 210.585 ;
        RECT 145.995 210.500 146.325 210.585 ;
        RECT 140.275 209.070 140.445 209.465 ;
        RECT 139.815 208.790 140.445 209.070 ;
        RECT 138.995 208.360 139.645 208.610 ;
        RECT 140.615 208.600 141.175 209.295 ;
        RECT 141.345 209.070 141.565 209.465 ;
        RECT 141.345 208.790 142.025 209.070 ;
        RECT 138.655 207.920 139.280 208.180 ;
        RECT 138.655 207.320 138.825 207.920 ;
        RECT 139.475 207.800 139.645 208.360 ;
        RECT 139.815 208.200 142.025 208.600 ;
        RECT 142.195 208.120 142.365 209.590 ;
        RECT 142.640 209.685 143.685 209.855 ;
        RECT 143.905 209.705 144.235 209.905 ;
        RECT 144.415 209.985 145.085 210.185 ;
        RECT 145.255 210.330 145.830 210.415 ;
        RECT 146.560 210.330 147.465 210.415 ;
        RECT 145.255 210.160 147.465 210.330 ;
        RECT 147.635 209.985 147.805 210.585 ;
        RECT 144.415 209.815 145.925 209.985 ;
        RECT 144.915 209.725 145.925 209.815 ;
        RECT 146.485 209.725 147.805 209.985 ;
        RECT 142.640 208.750 142.810 209.685 ;
        RECT 142.980 209.155 143.345 209.515 ;
        RECT 143.515 209.495 143.685 209.685 ;
        RECT 143.515 209.325 144.635 209.495 ;
        RECT 142.980 208.985 144.265 209.155 ;
        RECT 143.280 208.575 143.875 208.815 ;
        RECT 144.045 208.630 144.265 208.985 ;
        RECT 144.465 208.820 144.635 209.325 ;
        RECT 142.535 208.405 143.090 208.540 ;
        RECT 144.465 208.460 144.635 208.625 ;
        RECT 144.195 208.405 144.635 208.460 ;
        RECT 142.535 208.290 144.635 208.405 ;
        RECT 144.915 208.490 145.085 209.725 ;
        RECT 145.255 209.380 146.665 209.550 ;
        RECT 147.635 209.540 147.805 209.725 ;
        RECT 145.255 209.060 145.825 209.380 ;
        RECT 145.255 208.660 145.825 208.890 ;
        RECT 145.995 208.805 146.325 209.210 ;
        RECT 146.495 209.030 146.665 209.380 ;
        RECT 146.835 209.210 147.805 209.540 ;
        RECT 146.495 208.780 147.465 209.030 ;
        RECT 142.960 208.235 144.325 208.290 ;
        RECT 144.915 208.120 145.485 208.490 ;
        RECT 140.275 207.820 141.565 208.030 ;
        RECT 139.475 207.750 140.105 207.800 ;
        RECT 138.995 207.530 140.105 207.750 ;
        RECT 138.995 207.500 139.645 207.530 ;
        RECT 138.655 207.060 139.280 207.320 ;
        RECT 138.655 206.475 138.825 207.060 ;
        RECT 139.475 206.890 139.645 207.500 ;
        RECT 140.275 207.360 140.445 207.820 ;
        RECT 139.815 207.075 140.445 207.360 ;
        RECT 140.615 206.960 141.175 207.650 ;
        RECT 141.345 207.360 141.565 207.820 ;
        RECT 142.195 207.855 142.825 208.120 ;
        RECT 144.455 208.070 145.485 208.120 ;
        RECT 142.195 207.800 142.365 207.855 ;
        RECT 141.735 207.530 142.365 207.800 ;
        RECT 143.335 207.785 144.285 208.065 ;
        RECT 144.455 207.870 145.085 208.070 ;
        RECT 145.655 207.900 145.825 208.660 ;
        RECT 145.995 208.340 147.125 208.590 ;
        RECT 141.345 207.075 142.025 207.360 ;
        RECT 142.195 207.260 142.365 207.530 ;
        RECT 142.535 207.430 144.655 207.615 ;
        RECT 144.915 207.560 145.085 207.870 ;
        RECT 145.255 207.730 145.825 207.900 ;
        RECT 145.995 207.940 147.125 208.140 ;
        RECT 145.995 207.895 146.325 207.940 ;
        RECT 147.295 207.770 147.465 208.780 ;
        RECT 144.915 207.260 145.825 207.560 ;
        RECT 145.995 207.320 146.275 207.710 ;
        RECT 146.445 207.600 147.465 207.770 ;
        RECT 138.995 206.645 139.645 206.890 ;
        RECT 138.655 206.200 139.280 206.475 ;
        RECT 139.475 206.330 139.645 206.645 ;
        RECT 142.195 206.930 142.865 207.260 ;
        RECT 143.035 207.025 144.365 207.255 ;
        RECT 142.195 206.330 142.365 206.930 ;
        RECT 143.035 206.760 143.205 207.025 ;
        RECT 142.535 206.590 143.205 206.760 ;
        RECT 143.375 206.505 144.025 206.855 ;
        RECT 144.195 206.760 144.365 207.025 ;
        RECT 144.535 207.110 145.825 207.260 ;
        RECT 146.445 207.150 146.615 207.600 ;
        RECT 147.635 207.430 147.805 209.210 ;
        RECT 144.535 206.930 145.085 207.110 ;
        RECT 145.995 206.980 146.615 207.150 ;
        RECT 146.785 207.115 147.805 207.430 ;
        RECT 144.195 206.590 144.655 206.760 ;
        RECT 138.655 205.615 138.825 206.200 ;
        RECT 139.475 206.040 140.370 206.330 ;
        RECT 141.030 206.040 142.365 206.330 ;
        RECT 144.915 206.330 145.085 206.930 ;
        RECT 145.265 206.810 145.825 206.940 ;
        RECT 146.835 206.810 147.465 206.940 ;
        RECT 145.265 206.500 147.465 206.810 ;
        RECT 147.635 206.330 147.805 207.115 ;
        RECT 142.535 206.070 143.205 206.240 ;
        RECT 139.475 206.030 139.645 206.040 ;
        RECT 138.995 205.785 139.645 206.030 ;
        RECT 142.195 205.900 142.365 206.040 ;
        RECT 138.655 205.355 139.280 205.615 ;
        RECT 139.475 205.440 139.645 205.785 ;
        RECT 139.815 205.695 142.025 205.865 ;
        RECT 139.815 205.610 140.385 205.695 ;
        RECT 141.055 205.530 142.025 205.695 ;
        RECT 142.195 205.570 142.865 205.900 ;
        RECT 143.035 205.805 143.205 206.070 ;
        RECT 143.375 205.975 144.025 206.325 ;
        RECT 144.195 206.070 144.655 206.240 ;
        RECT 144.195 205.805 144.365 206.070 ;
        RECT 144.915 206.040 145.810 206.330 ;
        RECT 146.470 206.040 147.805 206.330 ;
        RECT 144.915 205.900 145.085 206.040 ;
        RECT 143.035 205.575 144.365 205.805 ;
        RECT 144.535 205.570 145.085 205.900 ;
        RECT 140.555 205.440 140.885 205.525 ;
        RECT 138.655 204.755 138.825 205.355 ;
        RECT 139.475 205.185 140.045 205.440 ;
        RECT 138.995 205.110 140.045 205.185 ;
        RECT 140.215 205.270 140.885 205.440 ;
        RECT 142.195 205.360 142.365 205.570 ;
        RECT 138.995 204.925 139.645 205.110 ;
        RECT 138.655 204.495 139.280 204.755 ;
        RECT 138.655 203.895 138.825 204.495 ;
        RECT 139.475 204.325 139.645 204.925 ;
        RECT 140.215 204.685 140.385 205.270 ;
        RECT 141.055 205.190 142.365 205.360 ;
        RECT 142.535 205.215 144.655 205.400 ;
        RECT 140.555 205.020 140.885 205.045 ;
        RECT 140.555 204.850 142.025 205.020 ;
        RECT 138.995 204.065 139.645 204.325 ;
        RECT 139.815 204.680 140.385 204.685 ;
        RECT 139.815 204.510 141.685 204.680 ;
        RECT 139.815 204.155 140.180 204.510 ;
        RECT 140.375 204.170 141.345 204.340 ;
        RECT 138.655 203.635 139.280 203.895 ;
        RECT 139.475 203.465 139.645 204.065 ;
        RECT 140.665 203.965 140.835 203.970 ;
        RECT 139.815 203.690 140.975 203.965 ;
        RECT 141.175 203.520 141.345 204.170 ;
        RECT 141.515 203.555 141.685 204.510 ;
        RECT 138.915 203.205 139.645 203.465 ;
        RECT 139.815 203.330 141.345 203.520 ;
        RECT 139.475 203.150 139.645 203.205 ;
        RECT 141.855 203.160 142.025 204.850 ;
        RECT 137.100 202.785 139.295 203.035 ;
        RECT 134.035 202.045 134.205 202.185 ;
        RECT 133.555 201.800 134.205 202.045 ;
        RECT 134.885 202.005 135.185 202.465 ;
        RECT 135.435 202.345 135.695 202.515 ;
        RECT 136.755 202.345 137.735 202.605 ;
        RECT 135.365 202.175 135.695 202.345 ;
        RECT 135.955 202.175 136.925 202.345 ;
        RECT 133.215 201.370 133.840 201.630 ;
        RECT 133.215 200.770 133.385 201.370 ;
        RECT 134.035 201.190 134.205 201.800 ;
        RECT 134.485 201.835 136.585 202.005 ;
        RECT 134.485 201.600 134.655 201.835 ;
        RECT 136.255 201.755 136.585 201.835 ;
        RECT 136.755 201.745 136.925 202.175 ;
        RECT 138.235 202.175 138.485 202.785 ;
        RECT 139.475 202.640 140.180 203.150 ;
        RECT 139.475 202.605 139.645 202.640 ;
        RECT 138.950 202.345 139.645 202.605 ;
        RECT 140.455 202.420 140.625 203.130 ;
        RECT 138.235 202.170 139.295 202.175 ;
        RECT 137.095 201.925 139.295 202.170 ;
        RECT 135.365 201.475 136.085 201.665 ;
        RECT 133.555 200.940 134.205 201.190 ;
        RECT 133.215 200.510 133.840 200.770 ;
        RECT 133.215 199.910 133.385 200.510 ;
        RECT 134.035 200.370 134.205 200.940 ;
        RECT 134.485 200.815 134.655 201.430 ;
        RECT 134.825 201.305 135.155 201.450 ;
        RECT 134.825 200.985 136.115 201.305 ;
        RECT 136.285 200.815 136.455 201.530 ;
        RECT 134.485 200.645 136.455 200.815 ;
        RECT 136.755 201.450 137.735 201.745 ;
        RECT 136.755 200.715 136.925 201.450 ;
        RECT 138.235 201.440 138.795 201.755 ;
        RECT 139.475 201.745 139.645 202.345 ;
        RECT 139.850 202.240 140.625 202.420 ;
        RECT 141.000 202.990 142.025 203.160 ;
        RECT 142.195 204.975 142.365 205.190 ;
        RECT 142.195 204.710 142.825 204.975 ;
        RECT 143.335 204.765 144.285 205.045 ;
        RECT 144.915 204.960 145.085 205.570 ;
        RECT 144.455 204.710 145.085 204.960 ;
        RECT 141.000 202.410 141.190 202.990 ;
        RECT 142.195 202.820 142.365 204.710 ;
        RECT 142.960 204.540 144.325 204.595 ;
        RECT 142.535 204.425 144.635 204.540 ;
        RECT 142.535 204.290 143.090 204.425 ;
        RECT 144.195 204.370 144.635 204.425 ;
        RECT 142.640 203.145 142.810 204.080 ;
        RECT 143.280 204.015 143.875 204.255 ;
        RECT 144.465 204.205 144.635 204.370 ;
        RECT 144.915 204.380 145.085 204.710 ;
        RECT 145.255 204.550 145.885 204.835 ;
        RECT 144.045 203.845 144.265 204.200 ;
        RECT 144.915 204.110 145.545 204.380 ;
        RECT 142.980 203.675 144.265 203.845 ;
        RECT 142.980 203.315 143.345 203.675 ;
        RECT 144.465 203.505 144.635 204.010 ;
        RECT 143.515 203.335 144.635 203.505 ;
        RECT 143.515 203.145 143.685 203.335 ;
        RECT 142.640 202.975 143.685 203.145 ;
        RECT 141.435 202.805 142.365 202.820 ;
        RECT 143.425 202.805 143.685 202.975 ;
        RECT 143.905 202.925 144.235 203.125 ;
        RECT 144.915 203.015 145.085 204.110 ;
        RECT 145.715 204.090 145.885 204.550 ;
        RECT 146.055 204.260 146.615 204.950 ;
        RECT 146.785 204.550 147.465 204.835 ;
        RECT 146.785 204.090 147.005 204.550 ;
        RECT 147.635 204.380 147.805 206.040 ;
        RECT 147.175 204.110 147.805 204.380 ;
        RECT 145.715 203.880 147.005 204.090 ;
        RECT 145.255 203.310 147.465 203.710 ;
        RECT 141.435 202.650 143.165 202.805 ;
        RECT 142.195 202.635 143.165 202.650 ;
        RECT 143.425 202.635 143.755 202.805 ;
        RECT 141.435 202.240 141.845 202.415 ;
        RECT 139.850 202.175 141.845 202.240 ;
        RECT 140.455 201.900 141.845 202.175 ;
        RECT 138.965 201.440 139.645 201.745 ;
        RECT 137.095 200.990 139.305 201.270 ;
        RECT 137.095 200.885 138.065 200.990 ;
        RECT 138.735 200.885 139.305 200.990 ;
        RECT 139.475 201.105 139.645 201.440 ;
        RECT 139.475 200.865 140.155 201.105 ;
        RECT 138.235 200.715 138.565 200.820 ;
        RECT 139.475 200.715 139.645 200.865 ;
        RECT 140.325 200.855 140.885 201.210 ;
        RECT 134.035 200.330 134.735 200.370 ;
        RECT 133.555 200.160 134.735 200.330 ;
        RECT 133.555 200.080 134.205 200.160 ;
        RECT 133.215 199.650 133.840 199.910 ;
        RECT 133.215 199.475 133.385 199.650 ;
        RECT 131.315 199.210 132.215 199.465 ;
        RECT 130.465 198.670 131.145 198.950 ;
        RECT 131.315 198.580 131.485 199.210 ;
        RECT 132.400 199.040 133.385 199.475 ;
        RECT 134.035 199.470 134.205 200.080 ;
        RECT 135.115 199.940 135.445 200.645 ;
        RECT 135.650 199.920 136.025 200.475 ;
        RECT 136.755 200.465 137.385 200.715 ;
        RECT 136.255 200.390 137.385 200.465 ;
        RECT 136.255 200.150 136.925 200.390 ;
        RECT 134.420 199.770 134.945 199.900 ;
        RECT 135.650 199.770 136.585 199.920 ;
        RECT 134.420 199.580 136.585 199.770 ;
        RECT 134.420 199.570 135.445 199.580 ;
        RECT 133.555 199.400 134.205 199.470 ;
        RECT 133.555 199.230 134.815 199.400 ;
        RECT 133.555 199.210 134.205 199.230 ;
        RECT 131.660 198.780 133.840 199.040 ;
        RECT 131.660 198.750 133.385 198.780 ;
        RECT 128.935 198.080 131.145 198.480 ;
        RECT 131.315 198.310 132.230 198.580 ;
        RECT 132.400 198.310 133.385 198.750 ;
        RECT 134.035 198.610 134.205 199.210 ;
        RECT 134.425 198.905 134.945 199.060 ;
        RECT 135.115 199.020 135.445 199.570 ;
        RECT 136.755 199.410 136.925 200.150 ;
        RECT 137.555 200.265 138.845 200.715 ;
        RECT 139.015 200.390 139.645 200.715 ;
        RECT 141.055 200.695 141.400 201.085 ;
        RECT 142.195 200.925 142.365 202.635 ;
        RECT 143.935 202.465 144.235 202.925 ;
        RECT 144.415 202.645 145.085 203.015 ;
        RECT 145.255 202.840 145.885 203.120 ;
        RECT 142.535 202.295 144.635 202.465 ;
        RECT 142.535 202.215 142.865 202.295 ;
        RECT 142.665 201.275 142.835 201.990 ;
        RECT 143.035 201.935 143.755 202.125 ;
        RECT 144.465 202.060 144.635 202.295 ;
        RECT 144.915 202.320 145.085 202.645 ;
        RECT 145.715 202.445 145.885 202.840 ;
        RECT 146.055 202.615 146.615 203.310 ;
        RECT 146.785 202.840 147.465 203.120 ;
        RECT 146.785 202.445 147.005 202.840 ;
        RECT 144.915 201.995 145.545 202.320 ;
        RECT 145.715 201.995 147.005 202.445 ;
        RECT 147.635 202.320 147.805 204.110 ;
        RECT 147.175 201.995 147.805 202.320 ;
        RECT 143.965 201.765 144.295 201.910 ;
        RECT 143.005 201.445 144.295 201.765 ;
        RECT 144.465 201.275 144.635 201.890 ;
        RECT 142.665 201.105 144.635 201.275 ;
        RECT 141.055 200.685 141.225 200.695 ;
        RECT 139.825 200.515 141.225 200.685 ;
        RECT 139.825 200.405 140.155 200.515 ;
        RECT 137.555 199.870 137.775 200.265 ;
        RECT 137.095 199.590 137.775 199.870 ;
        RECT 135.745 199.240 136.925 199.410 ;
        RECT 137.945 199.400 138.505 200.095 ;
        RECT 138.675 199.870 138.845 200.265 ;
        RECT 139.475 200.175 139.645 200.390 ;
        RECT 139.475 199.960 140.155 200.175 ;
        RECT 140.325 200.080 140.885 200.345 ;
        RECT 138.675 199.590 139.305 199.870 ;
        RECT 134.425 198.850 134.985 198.905 ;
        RECT 135.615 198.895 136.540 199.070 ;
        RECT 135.565 198.850 136.540 198.895 ;
        RECT 134.425 198.740 136.540 198.850 ;
        RECT 134.425 198.730 135.695 198.740 ;
        RECT 134.860 198.680 135.695 198.730 ;
        RECT 133.555 198.310 134.205 198.610 ;
        RECT 129.395 197.700 130.685 197.910 ;
        RECT 126.675 197.240 127.965 197.450 ;
        RECT 122.205 196.245 122.535 196.390 ;
        RECT 121.245 195.925 122.535 196.245 ;
        RECT 122.705 195.755 122.875 196.370 ;
        RECT 120.905 195.585 122.875 195.755 ;
        RECT 123.155 196.320 123.820 196.720 ;
        RECT 124.185 196.690 124.715 197.080 ;
        RECT 123.155 195.730 123.325 196.320 ;
        RECT 124.185 196.260 124.565 196.690 ;
        RECT 124.885 196.395 125.195 197.090 ;
        RECT 125.875 197.085 126.505 197.220 ;
        RECT 125.405 196.950 126.505 197.085 ;
        RECT 125.405 196.400 126.045 196.950 ;
        RECT 126.675 196.780 126.895 197.240 ;
        RECT 126.215 196.495 126.895 196.780 ;
        RECT 123.495 196.090 124.015 196.150 ;
        RECT 124.820 196.090 125.605 196.220 ;
        RECT 123.495 195.915 125.605 196.090 ;
        RECT 125.875 196.210 126.045 196.400 ;
        RECT 127.065 196.380 127.625 197.070 ;
        RECT 127.795 196.780 127.965 197.240 ;
        RECT 128.595 197.410 129.225 197.680 ;
        RECT 128.595 197.220 128.765 197.410 ;
        RECT 129.395 197.240 129.565 197.700 ;
        RECT 128.135 196.950 128.765 197.220 ;
        RECT 128.935 196.955 129.565 197.240 ;
        RECT 127.795 196.495 128.425 196.780 ;
        RECT 128.595 196.670 128.765 196.950 ;
        RECT 129.735 196.840 130.295 197.530 ;
        RECT 130.465 197.240 130.685 197.700 ;
        RECT 131.315 197.680 131.485 198.310 ;
        RECT 134.035 198.050 134.205 198.310 ;
        RECT 136.755 198.600 136.925 199.240 ;
        RECT 137.095 199.000 139.305 199.400 ;
        RECT 139.475 198.910 139.645 199.960 ;
        RECT 141.055 199.830 141.225 200.515 ;
        RECT 142.195 200.610 142.865 200.925 ;
        RECT 142.195 200.210 142.365 200.610 ;
        RECT 143.095 200.380 143.470 200.935 ;
        RECT 143.675 200.400 144.005 201.105 ;
        RECT 144.915 200.830 145.085 201.995 ;
        RECT 145.995 201.890 146.325 201.995 ;
        RECT 145.255 201.720 145.825 201.825 ;
        RECT 146.495 201.720 147.465 201.825 ;
        RECT 145.255 201.440 147.465 201.720 ;
        RECT 144.385 200.620 145.085 200.830 ;
        RECT 141.395 199.880 142.365 200.210 ;
        RECT 142.535 200.230 143.470 200.380 ;
        RECT 144.175 200.230 144.700 200.360 ;
        RECT 142.535 200.040 144.700 200.230 ;
        RECT 139.815 199.490 140.385 199.790 ;
        RECT 140.555 199.660 141.225 199.830 ;
        RECT 142.195 199.870 142.365 199.880 ;
        RECT 143.675 200.030 144.700 200.040 ;
        RECT 144.915 200.345 145.085 200.620 ;
        RECT 147.635 200.345 147.805 201.995 ;
        RECT 144.915 200.085 145.925 200.345 ;
        RECT 146.485 200.085 147.805 200.345 ;
        RECT 141.405 199.490 142.025 199.710 ;
        RECT 139.815 199.175 142.025 199.490 ;
        RECT 142.195 199.700 143.375 199.870 ;
        RECT 142.195 198.910 142.365 199.700 ;
        RECT 142.580 199.355 143.505 199.530 ;
        RECT 143.675 199.480 144.005 200.030 ;
        RECT 144.915 199.860 145.085 200.085 ;
        RECT 144.305 199.690 145.085 199.860 ;
        RECT 144.175 199.365 144.695 199.520 ;
        RECT 142.580 199.310 143.555 199.355 ;
        RECT 144.135 199.310 144.695 199.365 ;
        RECT 142.580 199.200 144.695 199.310 ;
        RECT 143.425 199.190 144.695 199.200 ;
        RECT 144.915 199.485 145.085 199.690 ;
        RECT 145.255 199.740 147.465 199.910 ;
        RECT 145.255 199.655 145.830 199.740 ;
        RECT 146.560 199.655 147.465 199.740 ;
        RECT 145.995 199.485 146.325 199.570 ;
        RECT 147.635 199.485 147.805 200.085 ;
        RECT 143.425 199.140 144.260 199.190 ;
        RECT 144.915 199.155 145.465 199.485 ;
        RECT 145.635 199.315 146.705 199.485 ;
        RECT 137.555 198.620 138.845 198.830 ;
        RECT 136.755 198.330 137.385 198.600 ;
        RECT 136.755 198.050 136.925 198.330 ;
        RECT 137.555 198.160 137.775 198.620 ;
        RECT 130.855 197.495 131.485 197.680 ;
        RECT 131.655 197.770 133.865 198.050 ;
        RECT 131.655 197.665 132.625 197.770 ;
        RECT 133.295 197.665 133.865 197.770 ;
        RECT 134.035 197.780 134.840 198.050 ;
        RECT 135.800 197.780 136.925 198.050 ;
        RECT 137.095 197.875 137.775 198.160 ;
        RECT 132.795 197.495 133.125 197.600 ;
        RECT 134.035 197.495 134.205 197.780 ;
        RECT 130.855 197.410 131.945 197.495 ;
        RECT 130.465 196.955 131.145 197.240 ;
        RECT 131.315 197.170 131.945 197.410 ;
        RECT 131.315 196.670 131.485 197.170 ;
        RECT 128.595 196.210 130.055 196.670 ;
        RECT 125.875 195.730 127.135 196.210 ;
        RECT 117.180 195.280 117.885 195.460 ;
        RECT 116.735 194.880 117.510 195.060 ;
        RECT 115.515 194.815 117.510 194.880 ;
        RECT 117.715 194.850 117.885 195.280 ;
        RECT 120.435 195.405 120.605 195.460 ;
        RECT 118.055 195.030 118.605 195.200 ;
        RECT 115.515 194.540 116.905 194.815 ;
        RECT 117.715 194.520 118.265 194.850 ;
        RECT 118.435 194.705 118.605 195.030 ;
        RECT 118.785 194.940 119.155 195.270 ;
        RECT 119.335 195.030 120.265 195.200 ;
        RECT 120.435 195.090 121.105 195.405 ;
        RECT 119.335 194.705 119.505 195.030 ;
        RECT 120.435 194.850 120.605 195.090 ;
        RECT 121.335 194.860 121.710 195.415 ;
        RECT 121.915 194.880 122.245 195.585 ;
        RECT 123.155 195.460 123.960 195.730 ;
        RECT 124.920 195.460 127.135 195.730 ;
        RECT 123.155 195.310 123.325 195.460 ;
        RECT 122.625 195.290 123.325 195.310 ;
        RECT 125.875 195.290 127.135 195.460 ;
        RECT 122.625 195.100 124.615 195.290 ;
        RECT 118.435 194.535 119.505 194.705 ;
        RECT 117.715 193.470 117.885 194.520 ;
        RECT 118.860 194.420 119.190 194.535 ;
        RECT 119.675 194.520 120.605 194.850 ;
        RECT 120.775 194.710 121.710 194.860 ;
        RECT 122.415 194.710 122.940 194.840 ;
        RECT 120.775 194.520 122.940 194.710 ;
        RECT 120.435 194.350 120.605 194.520 ;
        RECT 121.915 194.510 122.940 194.520 ;
        RECT 118.055 194.250 118.560 194.340 ;
        RECT 119.360 194.250 120.265 194.350 ;
        RECT 118.055 194.080 120.265 194.250 ;
        RECT 120.435 194.180 121.615 194.350 ;
        RECT 118.055 193.650 118.605 193.820 ;
        RECT 117.715 193.450 118.265 193.470 ;
        RECT 112.275 193.160 113.170 193.450 ;
        RECT 113.830 193.160 116.330 193.450 ;
        RECT 116.990 193.160 118.265 193.450 ;
        RECT 112.275 191.595 112.445 193.160 ;
        RECT 114.995 192.435 115.165 193.160 ;
        RECT 117.715 193.140 118.265 193.160 ;
        RECT 118.435 193.325 118.605 193.650 ;
        RECT 118.785 193.560 119.155 193.890 ;
        RECT 119.335 193.650 120.265 193.820 ;
        RECT 119.335 193.325 119.505 193.650 ;
        RECT 120.435 193.470 120.605 194.180 ;
        RECT 120.820 193.835 121.745 194.010 ;
        RECT 121.915 193.960 122.245 194.510 ;
        RECT 123.155 194.340 124.615 195.100 ;
        RECT 122.545 194.170 124.615 194.340 ;
        RECT 123.155 194.080 124.615 194.170 ;
        RECT 124.785 194.830 127.135 195.290 ;
        RECT 127.305 196.150 130.055 196.210 ;
        RECT 127.305 195.460 129.515 196.150 ;
        RECT 130.225 195.980 131.485 196.670 ;
        RECT 132.115 197.045 133.405 197.495 ;
        RECT 133.575 197.190 134.205 197.495 ;
        RECT 134.375 197.420 136.485 197.595 ;
        RECT 134.375 197.360 134.895 197.420 ;
        RECT 135.700 197.290 136.485 197.420 ;
        RECT 136.755 197.590 136.925 197.780 ;
        RECT 137.945 197.760 138.505 198.450 ;
        RECT 138.675 198.160 138.845 198.620 ;
        RECT 139.475 198.700 140.465 198.910 ;
        RECT 141.055 198.700 142.365 198.910 ;
        RECT 139.475 198.600 139.645 198.700 ;
        RECT 139.015 198.330 139.645 198.600 ;
        RECT 138.675 197.875 139.305 198.160 ;
        RECT 139.475 198.030 139.645 198.330 ;
        RECT 139.815 198.280 142.025 198.530 ;
        RECT 139.815 198.200 140.445 198.280 ;
        RECT 141.045 198.200 142.025 198.280 ;
        RECT 142.195 198.230 142.365 198.700 ;
        RECT 142.535 198.620 144.745 198.935 ;
        RECT 142.535 198.400 143.155 198.620 ;
        RECT 143.335 198.280 144.005 198.450 ;
        RECT 144.175 198.320 144.745 198.620 ;
        RECT 139.475 197.800 140.465 198.030 ;
        RECT 139.475 197.590 139.645 197.800 ;
        RECT 140.635 197.780 140.885 198.110 ;
        RECT 142.195 198.030 143.165 198.230 ;
        RECT 141.055 197.900 143.165 198.030 ;
        RECT 141.055 197.800 142.365 197.900 ;
        RECT 133.575 197.170 134.700 197.190 ;
        RECT 132.115 196.650 132.335 197.045 ;
        RECT 131.655 196.370 132.335 196.650 ;
        RECT 132.505 196.180 133.065 196.875 ;
        RECT 133.235 196.650 133.405 197.045 ;
        RECT 134.035 196.790 134.700 197.170 ;
        RECT 135.065 196.820 135.445 197.250 ;
        RECT 133.235 196.370 133.865 196.650 ;
        RECT 129.685 195.460 131.485 195.980 ;
        RECT 131.655 195.780 133.865 196.180 ;
        RECT 127.305 195.000 128.765 195.460 ;
        RECT 131.315 195.380 131.485 195.460 ;
        RECT 132.115 195.400 133.405 195.610 ;
        RECT 129.095 195.120 131.145 195.290 ;
        RECT 129.095 195.015 129.440 195.120 ;
        RECT 130.175 195.015 131.145 195.120 ;
        RECT 131.315 195.110 131.945 195.380 ;
        RECT 122.415 193.845 122.935 194.000 ;
        RECT 120.820 193.790 121.795 193.835 ;
        RECT 122.375 193.790 122.935 193.845 ;
        RECT 120.820 193.680 122.935 193.790 ;
        RECT 121.665 193.670 122.935 193.680 ;
        RECT 121.665 193.620 122.500 193.670 ;
        RECT 118.435 193.155 119.505 193.325 ;
        RECT 119.675 193.450 120.605 193.470 ;
        RECT 123.155 193.450 124.095 194.080 ;
        RECT 124.785 193.910 127.655 194.830 ;
        RECT 119.675 193.160 121.770 193.450 ;
        RECT 122.430 193.160 124.095 193.450 ;
        RECT 115.335 192.710 117.545 192.990 ;
        RECT 115.335 192.605 116.305 192.710 ;
        RECT 116.975 192.605 117.545 192.710 ;
        RECT 116.475 192.435 116.805 192.540 ;
        RECT 117.715 192.435 117.885 193.140 ;
        RECT 118.860 193.040 119.190 193.155 ;
        RECT 119.675 193.140 120.605 193.160 ;
        RECT 118.055 192.870 118.560 192.960 ;
        RECT 119.360 192.870 120.265 192.970 ;
        RECT 118.055 192.700 120.265 192.870 ;
        RECT 114.995 192.110 115.625 192.435 ;
        RECT 112.615 191.810 113.165 191.980 ;
        RECT 112.275 191.265 112.825 191.595 ;
        RECT 112.995 191.435 113.165 191.810 ;
        RECT 113.345 191.715 113.715 192.070 ;
        RECT 113.895 191.810 114.825 191.980 ;
        RECT 113.895 191.435 114.065 191.810 ;
        RECT 114.995 191.595 115.165 192.110 ;
        RECT 112.995 191.265 114.065 191.435 ;
        RECT 114.235 191.265 115.165 191.595 ;
        RECT 115.795 191.985 117.085 192.435 ;
        RECT 117.255 192.110 117.885 192.435 ;
        RECT 118.055 192.270 118.605 192.440 ;
        RECT 115.795 191.590 116.015 191.985 ;
        RECT 115.335 191.310 116.015 191.590 ;
        RECT 112.275 190.665 112.445 191.265 ;
        RECT 113.355 191.180 113.685 191.265 ;
        RECT 112.615 191.010 113.190 191.095 ;
        RECT 113.920 191.010 114.825 191.095 ;
        RECT 112.615 190.840 114.825 191.010 ;
        RECT 114.995 190.665 115.165 191.265 ;
        RECT 116.185 191.120 116.745 191.815 ;
        RECT 116.915 191.590 117.085 191.985 ;
        RECT 117.715 192.090 117.885 192.110 ;
        RECT 117.715 191.760 118.265 192.090 ;
        RECT 118.435 191.945 118.605 192.270 ;
        RECT 118.785 192.180 119.155 192.510 ;
        RECT 120.435 192.480 120.605 193.140 ;
        RECT 120.775 192.815 122.985 192.985 ;
        RECT 120.775 192.650 121.745 192.815 ;
        RECT 122.415 192.730 122.985 192.815 ;
        RECT 123.155 192.700 124.095 193.160 ;
        RECT 124.265 193.620 127.655 193.910 ;
        RECT 127.825 194.825 128.765 195.000 ;
        RECT 129.675 194.845 130.005 194.950 ;
        RECT 127.825 194.445 129.165 194.825 ;
        RECT 129.335 194.675 130.345 194.845 ;
        RECT 131.315 194.805 131.485 195.110 ;
        RECT 132.115 194.940 132.335 195.400 ;
        RECT 127.825 193.935 128.765 194.445 ;
        RECT 129.335 194.275 129.505 194.675 ;
        RECT 128.985 194.105 129.505 194.275 ;
        RECT 129.675 194.125 130.005 194.505 ;
        RECT 130.175 194.355 130.345 194.675 ;
        RECT 130.515 194.525 131.485 194.805 ;
        RECT 131.655 194.655 132.335 194.940 ;
        RECT 132.505 194.540 133.065 195.230 ;
        RECT 133.235 194.940 133.405 195.400 ;
        RECT 134.035 195.380 134.205 196.790 ;
        RECT 135.065 196.430 135.595 196.820 ;
        RECT 134.535 196.260 135.595 196.430 ;
        RECT 135.765 196.420 136.075 197.115 ;
        RECT 136.755 197.110 138.015 197.590 ;
        RECT 136.285 196.900 138.015 197.110 ;
        RECT 138.185 197.160 139.645 197.590 ;
        RECT 139.905 197.330 140.365 197.500 ;
        RECT 138.185 197.070 140.025 197.160 ;
        RECT 136.285 196.425 138.555 196.900 ;
        RECT 134.535 196.200 134.730 196.260 ;
        RECT 134.390 196.030 134.730 196.200 ;
        RECT 135.425 196.245 135.595 196.260 ;
        RECT 136.755 196.380 138.555 196.425 ;
        RECT 138.725 196.830 140.025 197.070 ;
        RECT 140.195 197.065 140.365 197.330 ;
        RECT 140.535 197.235 141.185 197.585 ;
        RECT 141.355 197.330 142.025 197.500 ;
        RECT 141.355 197.065 141.525 197.330 ;
        RECT 142.195 197.160 142.365 197.800 ;
        RECT 143.335 197.595 143.505 198.280 ;
        RECT 144.915 198.150 145.085 199.155 ;
        RECT 145.635 198.940 145.805 199.315 ;
        RECT 145.255 198.770 145.805 198.940 ;
        RECT 145.985 198.680 146.355 199.035 ;
        RECT 146.535 198.940 146.705 199.315 ;
        RECT 146.875 199.155 147.805 199.485 ;
        RECT 146.535 198.770 147.465 198.940 ;
        RECT 143.675 197.765 144.235 198.030 ;
        RECT 144.405 197.940 145.085 198.150 ;
        RECT 145.255 198.110 145.885 198.395 ;
        RECT 144.405 197.935 145.545 197.940 ;
        RECT 144.405 197.595 144.735 197.705 ;
        RECT 143.335 197.425 144.735 197.595 ;
        RECT 144.915 197.670 145.545 197.935 ;
        RECT 143.335 197.415 143.505 197.425 ;
        RECT 140.195 196.835 141.525 197.065 ;
        RECT 141.695 196.830 142.365 197.160 ;
        RECT 143.160 197.025 143.505 197.415 ;
        RECT 143.675 196.900 144.235 197.255 ;
        RECT 144.915 197.245 145.085 197.670 ;
        RECT 145.715 197.650 145.885 198.110 ;
        RECT 146.055 197.820 146.615 198.510 ;
        RECT 146.785 198.110 147.465 198.395 ;
        RECT 146.785 197.650 147.005 198.110 ;
        RECT 147.635 197.940 147.805 199.155 ;
        RECT 147.175 197.670 147.805 197.940 ;
        RECT 145.715 197.440 147.005 197.650 ;
        RECT 144.405 197.005 145.085 197.245 ;
        RECT 138.725 196.380 139.645 196.830 ;
        RECT 139.905 196.475 142.025 196.660 ;
        RECT 134.925 195.770 135.255 196.090 ;
        RECT 135.425 195.960 136.540 196.245 ;
        RECT 134.925 195.750 136.135 195.770 ;
        RECT 136.755 195.760 136.925 196.380 ;
        RECT 139.475 196.220 139.645 196.380 ;
        RECT 134.400 195.535 136.135 195.750 ;
        RECT 134.400 195.510 134.775 195.535 ;
        RECT 133.575 195.340 134.205 195.380 ;
        RECT 133.575 195.110 134.710 195.340 ;
        RECT 134.035 195.010 134.710 195.110 ;
        RECT 134.885 195.065 135.735 195.365 ;
        RECT 135.905 195.260 136.135 195.535 ;
        RECT 136.305 195.430 136.925 195.760 ;
        RECT 135.905 195.090 136.565 195.260 ;
        RECT 134.885 195.060 135.055 195.065 ;
        RECT 133.235 194.655 133.865 194.940 ;
        RECT 130.175 194.185 130.635 194.355 ;
        RECT 127.825 193.620 129.165 193.935 ;
        RECT 124.265 193.450 126.045 193.620 ;
        RECT 128.595 193.605 129.165 193.620 ;
        RECT 128.595 193.450 128.765 193.605 ;
        RECT 124.265 193.160 127.210 193.450 ;
        RECT 127.870 193.160 128.765 193.450 ;
        RECT 129.335 193.430 129.505 194.105 ;
        RECT 128.985 193.260 129.505 193.430 ;
        RECT 129.675 193.215 130.295 193.955 ;
        RECT 124.265 192.700 126.045 193.160 ;
        RECT 128.595 193.060 128.765 193.160 ;
        RECT 121.915 192.560 122.245 192.645 ;
        RECT 123.155 192.560 123.325 192.700 ;
        RECT 119.335 192.270 120.265 192.440 ;
        RECT 120.435 192.310 121.745 192.480 ;
        RECT 121.915 192.390 122.585 192.560 ;
        RECT 119.335 191.945 119.505 192.270 ;
        RECT 120.435 192.090 120.605 192.310 ;
        RECT 121.915 192.140 122.245 192.165 ;
        RECT 118.435 191.775 119.505 191.945 ;
        RECT 116.915 191.310 117.545 191.590 ;
        RECT 115.335 190.720 117.545 191.120 ;
        RECT 112.275 190.405 113.285 190.665 ;
        RECT 113.845 190.405 115.165 190.665 ;
        RECT 117.715 190.710 117.885 191.760 ;
        RECT 118.860 191.660 119.190 191.775 ;
        RECT 119.675 191.760 120.605 192.090 ;
        RECT 118.055 191.490 118.560 191.580 ;
        RECT 119.360 191.490 120.265 191.590 ;
        RECT 118.055 191.320 120.265 191.490 ;
        RECT 118.055 190.890 118.605 191.060 ;
        RECT 112.275 189.790 112.445 190.405 ;
        RECT 114.995 190.320 115.165 190.405 ;
        RECT 115.795 190.340 117.085 190.550 ;
        RECT 112.615 190.050 114.825 190.230 ;
        RECT 112.615 189.970 113.120 190.050 ;
        RECT 113.920 189.960 114.825 190.050 ;
        RECT 114.995 190.050 115.625 190.320 ;
        RECT 112.275 189.460 112.825 189.790 ;
        RECT 113.420 189.775 113.750 189.880 ;
        RECT 114.995 189.790 115.165 190.050 ;
        RECT 115.795 189.880 116.015 190.340 ;
        RECT 112.995 189.605 114.065 189.775 ;
        RECT 112.275 187.925 112.445 189.460 ;
        RECT 112.995 189.280 113.165 189.605 ;
        RECT 112.615 189.110 113.165 189.280 ;
        RECT 113.345 189.040 113.715 189.380 ;
        RECT 113.895 189.280 114.065 189.605 ;
        RECT 114.235 189.460 115.165 189.790 ;
        RECT 115.335 189.595 116.015 189.880 ;
        RECT 116.185 189.480 116.745 190.170 ;
        RECT 116.915 189.880 117.085 190.340 ;
        RECT 117.715 190.380 118.265 190.710 ;
        RECT 118.435 190.565 118.605 190.890 ;
        RECT 118.785 190.800 119.155 191.130 ;
        RECT 119.335 190.890 120.265 191.060 ;
        RECT 119.335 190.565 119.505 190.890 ;
        RECT 120.435 190.710 120.605 191.760 ;
        RECT 118.435 190.395 119.505 190.565 ;
        RECT 117.715 190.320 117.885 190.380 ;
        RECT 117.255 190.050 117.885 190.320 ;
        RECT 118.860 190.280 119.190 190.395 ;
        RECT 119.675 190.380 120.605 190.710 ;
        RECT 116.915 189.595 117.545 189.880 ;
        RECT 117.715 189.760 117.885 190.050 ;
        RECT 118.055 190.110 118.560 190.200 ;
        RECT 119.360 190.110 120.265 190.210 ;
        RECT 118.055 189.940 120.265 190.110 ;
        RECT 120.435 189.940 120.605 190.380 ;
        RECT 120.775 191.970 122.245 192.140 ;
        RECT 120.775 190.280 120.945 191.970 ;
        RECT 122.415 191.805 122.585 192.390 ;
        RECT 122.755 192.230 123.325 192.560 ;
        RECT 122.415 191.800 122.985 191.805 ;
        RECT 121.115 191.630 122.985 191.800 ;
        RECT 121.115 190.675 121.285 191.630 ;
        RECT 121.455 191.290 122.425 191.460 ;
        RECT 121.455 190.640 121.625 191.290 ;
        RECT 122.620 191.275 122.985 191.630 ;
        RECT 123.155 191.500 123.325 192.230 ;
        RECT 123.495 191.670 124.125 191.955 ;
        RECT 123.155 191.230 123.785 191.500 ;
        RECT 122.645 191.085 122.815 191.090 ;
        RECT 121.825 190.810 122.985 191.085 ;
        RECT 121.455 190.450 122.985 190.640 ;
        RECT 120.775 190.110 121.800 190.280 ;
        RECT 123.155 190.270 123.325 191.230 ;
        RECT 123.955 191.210 124.125 191.670 ;
        RECT 124.295 191.380 124.855 192.070 ;
        RECT 125.025 191.670 125.705 191.955 ;
        RECT 125.875 191.700 126.045 192.700 ;
        RECT 126.685 192.690 128.025 192.815 ;
        RECT 126.255 192.645 128.025 192.690 ;
        RECT 128.595 192.730 129.265 193.060 ;
        RECT 130.465 193.045 130.635 194.185 ;
        RECT 128.595 192.660 128.765 192.730 ;
        RECT 126.255 192.360 126.855 192.645 ;
        RECT 127.025 192.230 127.685 192.475 ;
        RECT 126.265 191.930 126.855 192.180 ;
        RECT 127.855 192.160 128.025 192.645 ;
        RECT 128.195 192.330 128.765 192.660 ;
        RECT 129.675 192.535 130.005 192.945 ;
        RECT 130.175 192.725 130.635 193.045 ;
        RECT 125.025 191.210 125.245 191.670 ;
        RECT 125.875 191.500 126.515 191.700 ;
        RECT 125.415 191.370 126.515 191.500 ;
        RECT 125.415 191.230 126.045 191.370 ;
        RECT 123.955 191.000 125.245 191.210 ;
        RECT 123.495 190.430 125.705 190.830 ;
        RECT 125.875 190.700 126.045 191.230 ;
        RECT 126.685 191.140 126.855 191.930 ;
        RECT 127.025 191.750 127.685 192.015 ;
        RECT 127.855 191.830 128.365 192.160 ;
        RECT 128.595 192.120 128.765 192.330 ;
        RECT 128.985 192.530 130.005 192.535 ;
        RECT 128.985 192.290 130.600 192.530 ;
        RECT 130.805 192.305 131.095 194.355 ;
        RECT 131.315 193.450 131.485 194.525 ;
        RECT 134.035 193.450 134.205 195.010 ;
        RECT 136.755 194.380 136.925 195.430 ;
        RECT 137.145 194.550 137.435 196.205 ;
        RECT 137.605 195.885 138.065 196.205 ;
        RECT 137.605 194.785 137.775 195.885 ;
        RECT 138.235 195.855 138.805 196.205 ;
        RECT 139.475 196.200 140.105 196.220 ;
        RECT 138.975 195.970 140.105 196.200 ;
        RECT 140.275 196.025 141.225 196.305 ;
        RECT 142.195 196.235 142.365 196.830 ;
        RECT 142.535 196.410 143.465 196.580 ;
        RECT 141.735 196.195 142.365 196.235 ;
        RECT 141.735 195.970 143.125 196.195 ;
        RECT 138.975 195.870 139.645 195.970 ;
        RECT 137.945 194.975 138.565 195.685 ;
        RECT 138.735 195.500 139.255 195.670 ;
        RECT 137.605 194.615 138.065 194.785 ;
        RECT 136.755 194.100 137.725 194.380 ;
        RECT 137.895 194.230 138.065 194.615 ;
        RECT 138.235 194.400 138.565 194.805 ;
        RECT 138.735 194.800 138.905 195.500 ;
        RECT 139.475 195.300 139.645 195.870 ;
        RECT 142.195 195.865 143.125 195.970 ;
        RECT 143.295 196.035 143.465 196.410 ;
        RECT 143.645 196.315 144.015 196.670 ;
        RECT 144.195 196.410 144.745 196.580 ;
        RECT 144.195 196.035 144.365 196.410 ;
        RECT 144.915 196.195 145.085 197.005 ;
        RECT 145.255 196.870 147.465 197.270 ;
        RECT 145.255 196.400 145.885 196.680 ;
        RECT 143.295 195.865 144.365 196.035 ;
        RECT 144.535 195.880 145.085 196.195 ;
        RECT 145.715 196.005 145.885 196.400 ;
        RECT 146.055 196.175 146.615 196.870 ;
        RECT 146.785 196.400 147.465 196.680 ;
        RECT 146.785 196.005 147.005 196.400 ;
        RECT 144.535 195.865 145.545 195.880 ;
        RECT 140.235 195.800 141.600 195.855 ;
        RECT 139.925 195.685 142.025 195.800 ;
        RECT 139.925 195.630 140.365 195.685 ;
        RECT 139.925 195.465 140.095 195.630 ;
        RECT 141.470 195.550 142.025 195.685 ;
        RECT 139.075 194.970 139.645 195.300 ;
        RECT 138.735 194.630 139.255 194.800 ;
        RECT 138.735 194.230 138.905 194.630 ;
        RECT 139.475 194.460 139.645 194.970 ;
        RECT 139.925 194.765 140.095 195.270 ;
        RECT 140.295 195.105 140.515 195.460 ;
        RECT 140.685 195.275 141.280 195.515 ;
        RECT 140.295 194.935 141.580 195.105 ;
        RECT 139.925 194.595 141.045 194.765 ;
        RECT 134.385 193.600 136.585 193.910 ;
        RECT 134.385 193.470 134.945 193.600 ;
        RECT 135.955 193.470 136.585 193.600 ;
        RECT 131.315 193.160 132.650 193.450 ;
        RECT 133.310 193.300 134.205 193.450 ;
        RECT 136.755 193.450 136.925 194.100 ;
        RECT 137.895 194.060 138.905 194.230 ;
        RECT 139.075 194.275 139.645 194.460 ;
        RECT 140.875 194.405 141.045 194.595 ;
        RECT 141.215 194.575 141.580 194.935 ;
        RECT 141.750 194.405 141.920 195.340 ;
        RECT 139.075 194.080 140.145 194.275 ;
        RECT 138.235 193.960 138.565 194.060 ;
        RECT 139.475 193.905 140.145 194.080 ;
        RECT 140.325 194.185 140.655 194.385 ;
        RECT 140.875 194.235 141.920 194.405 ;
        RECT 142.195 195.265 142.365 195.865 ;
        RECT 143.675 195.780 144.005 195.865 ;
        RECT 142.535 195.610 143.440 195.695 ;
        RECT 144.170 195.610 144.745 195.695 ;
        RECT 142.535 195.440 144.745 195.610 ;
        RECT 144.915 195.555 145.545 195.865 ;
        RECT 145.715 195.555 147.005 196.005 ;
        RECT 147.635 195.880 147.805 197.670 ;
        RECT 147.175 195.555 147.805 195.880 ;
        RECT 144.915 195.265 145.085 195.555 ;
        RECT 145.995 195.450 146.325 195.555 ;
        RECT 142.195 195.005 143.515 195.265 ;
        RECT 144.075 195.005 145.085 195.265 ;
        RECT 142.195 194.790 142.365 195.005 ;
        RECT 142.195 194.560 143.505 194.790 ;
        RECT 137.095 193.790 138.065 193.890 ;
        RECT 138.800 193.790 139.145 193.890 ;
        RECT 137.095 193.620 139.145 193.790 ;
        RECT 139.475 193.450 139.645 193.905 ;
        RECT 140.325 193.725 140.625 194.185 ;
        RECT 140.875 194.065 141.135 194.235 ;
        RECT 142.195 194.065 142.365 194.560 ;
        RECT 143.675 194.480 143.925 194.810 ;
        RECT 144.915 194.790 145.085 195.005 ;
        RECT 145.255 195.280 145.825 195.385 ;
        RECT 146.495 195.280 147.465 195.385 ;
        RECT 145.255 195.000 147.465 195.280 ;
        RECT 144.095 194.560 145.085 194.790 ;
        RECT 145.255 194.570 145.805 194.740 ;
        RECT 144.915 194.390 145.085 194.560 ;
        RECT 140.805 193.895 141.135 194.065 ;
        RECT 141.395 193.895 142.365 194.065 ;
        RECT 142.535 194.310 143.515 194.390 ;
        RECT 144.115 194.310 144.745 194.390 ;
        RECT 142.535 194.060 144.745 194.310 ;
        RECT 144.915 194.060 145.465 194.390 ;
        RECT 145.635 194.245 145.805 194.570 ;
        RECT 145.985 194.470 146.355 194.810 ;
        RECT 146.535 194.570 147.465 194.750 ;
        RECT 146.535 194.245 146.705 194.570 ;
        RECT 147.635 194.390 147.805 195.555 ;
        RECT 145.635 194.075 146.705 194.245 ;
        RECT 142.195 193.890 142.365 193.895 ;
        RECT 144.915 193.890 145.085 194.060 ;
        RECT 146.060 193.970 146.390 194.075 ;
        RECT 146.875 194.060 147.805 194.390 ;
        RECT 133.310 193.160 134.945 193.300 ;
        RECT 135.115 193.260 135.735 193.430 ;
        RECT 136.755 193.295 138.090 193.450 ;
        RECT 131.315 192.120 131.485 193.160 ;
        RECT 127.025 191.270 127.685 191.555 ;
        RECT 126.265 190.890 126.855 191.140 ;
        RECT 127.025 190.880 127.685 191.095 ;
        RECT 127.355 190.790 127.685 190.880 ;
        RECT 125.875 190.450 127.185 190.700 ;
        RECT 127.855 190.620 128.025 191.830 ;
        RECT 128.595 191.780 129.265 192.120 ;
        RECT 129.435 191.780 130.005 192.120 ;
        RECT 130.240 191.780 131.485 192.120 ;
        RECT 131.705 191.800 131.995 192.990 ;
        RECT 132.165 192.645 132.625 192.970 ;
        RECT 132.795 192.645 133.125 192.990 ;
        RECT 133.295 192.720 133.815 192.975 ;
        RECT 134.035 192.850 134.945 193.160 ;
        RECT 132.165 191.970 132.335 192.645 ;
        RECT 132.505 192.280 133.125 192.475 ;
        RECT 132.165 191.800 132.625 191.970 ;
        RECT 128.595 191.590 128.765 191.780 ;
        RECT 131.315 191.630 131.485 191.780 ;
        RECT 128.595 191.350 129.575 191.590 ;
        RECT 128.595 190.780 128.765 191.350 ;
        RECT 129.755 191.260 130.005 191.610 ;
        RECT 130.175 191.270 131.130 191.600 ;
        RECT 131.315 191.350 132.285 191.630 ;
        RECT 132.455 191.480 132.625 191.800 ;
        RECT 132.795 191.650 133.125 192.280 ;
        RECT 133.295 192.050 133.465 192.720 ;
        RECT 134.035 192.550 134.205 192.850 ;
        RECT 135.115 192.700 135.395 193.090 ;
        RECT 135.565 192.810 135.735 193.260 ;
        RECT 135.905 193.160 138.090 193.295 ;
        RECT 138.750 193.160 139.645 193.450 ;
        RECT 139.925 193.555 142.025 193.725 ;
        RECT 139.925 193.320 140.095 193.555 ;
        RECT 141.695 193.475 142.025 193.555 ;
        RECT 142.195 193.680 143.505 193.890 ;
        RECT 144.095 193.680 145.085 193.890 ;
        RECT 142.195 193.450 142.365 193.680 ;
        RECT 144.915 193.450 145.085 193.680 ;
        RECT 145.255 193.800 145.760 193.880 ;
        RECT 146.560 193.800 147.465 193.890 ;
        RECT 145.255 193.620 147.465 193.800 ;
        RECT 147.635 193.450 147.805 194.060 ;
        RECT 140.805 193.195 141.525 193.385 ;
        RECT 135.905 192.980 136.925 193.160 ;
        RECT 133.635 192.340 134.205 192.550 ;
        RECT 134.375 192.510 134.945 192.680 ;
        RECT 135.565 192.640 136.585 192.810 ;
        RECT 133.635 192.220 134.605 192.340 ;
        RECT 133.295 191.880 133.815 192.050 ;
        RECT 134.035 191.920 134.605 192.220 ;
        RECT 133.295 191.480 133.465 191.880 ;
        RECT 134.035 191.710 134.205 191.920 ;
        RECT 134.775 191.750 134.945 192.510 ;
        RECT 135.115 192.470 135.445 192.515 ;
        RECT 135.115 192.270 136.245 192.470 ;
        RECT 135.115 191.820 136.245 192.070 ;
        RECT 128.935 191.090 129.575 191.180 ;
        RECT 130.175 191.090 130.345 191.270 ;
        RECT 128.935 190.920 130.345 191.090 ;
        RECT 128.935 190.850 129.575 190.920 ;
        RECT 127.355 190.450 128.025 190.620 ;
        RECT 128.195 190.680 128.765 190.780 ;
        RECT 128.195 190.450 129.575 190.680 ;
        RECT 120.435 189.770 121.365 189.940 ;
        RECT 117.715 189.490 118.695 189.760 ;
        RECT 113.895 189.100 114.825 189.280 ;
        RECT 114.995 188.380 115.165 189.460 ;
        RECT 117.715 188.820 117.885 189.490 ;
        RECT 118.875 189.420 119.125 189.770 ;
        RECT 120.435 189.760 120.605 189.770 ;
        RECT 119.295 189.430 120.605 189.760 ;
        RECT 118.055 189.250 118.695 189.320 ;
        RECT 118.055 189.080 119.465 189.250 ;
        RECT 118.055 188.990 118.695 189.080 ;
        RECT 117.715 188.580 118.695 188.820 ;
        RECT 114.995 188.050 115.885 188.380 ;
        RECT 116.185 188.160 116.725 188.390 ;
        RECT 116.525 188.060 116.725 188.160 ;
        RECT 116.895 188.050 117.545 188.390 ;
        RECT 112.275 187.590 112.950 187.925 ;
        RECT 112.275 186.165 112.445 187.590 ;
        RECT 113.125 187.570 113.975 187.870 ;
        RECT 114.145 187.670 114.805 187.840 ;
        RECT 112.640 187.400 113.015 187.420 ;
        RECT 114.145 187.400 114.375 187.670 ;
        RECT 114.995 187.500 115.165 188.050 ;
        RECT 115.410 187.750 116.705 187.870 ;
        RECT 115.410 187.655 116.725 187.750 ;
        RECT 112.640 187.180 114.375 187.400 ;
        RECT 113.165 187.165 114.375 187.180 ;
        RECT 114.545 187.170 115.165 187.500 ;
        RECT 112.630 186.730 112.970 186.900 ;
        RECT 113.165 186.865 113.495 187.165 ;
        RECT 112.775 186.695 112.970 186.730 ;
        RECT 113.665 186.710 114.780 186.995 ;
        RECT 114.995 186.960 115.165 187.170 ;
        RECT 115.335 187.130 116.325 187.460 ;
        RECT 116.525 187.420 116.725 187.655 ;
        RECT 116.895 187.540 117.085 188.050 ;
        RECT 117.715 187.880 117.885 188.580 ;
        RECT 118.875 188.560 119.125 188.910 ;
        RECT 119.295 188.900 119.465 189.080 ;
        RECT 119.295 188.570 120.250 188.900 ;
        RECT 120.435 188.410 120.605 189.430 ;
        RECT 120.955 189.360 121.365 189.535 ;
        RECT 121.610 189.530 121.800 190.110 ;
        RECT 122.175 189.540 122.345 190.250 ;
        RECT 122.620 189.760 123.325 190.270 ;
        RECT 123.495 189.960 124.125 190.240 ;
        RECT 122.175 189.360 122.950 189.540 ;
        RECT 120.955 189.295 122.950 189.360 ;
        RECT 123.155 189.440 123.325 189.760 ;
        RECT 123.955 189.565 124.125 189.960 ;
        RECT 124.295 189.735 124.855 190.430 ;
        RECT 125.025 189.960 125.705 190.240 ;
        RECT 125.025 189.565 125.245 189.960 ;
        RECT 120.955 189.020 122.345 189.295 ;
        RECT 123.155 189.115 123.785 189.440 ;
        RECT 123.955 189.115 125.245 189.565 ;
        RECT 125.875 189.440 126.045 190.450 ;
        RECT 127.355 190.310 127.685 190.450 ;
        RECT 128.595 190.410 129.575 190.450 ;
        RECT 126.255 190.140 127.105 190.280 ;
        RECT 127.870 190.140 128.380 190.280 ;
        RECT 126.255 189.950 128.380 190.140 ;
        RECT 125.415 189.115 126.045 189.440 ;
        RECT 120.775 188.590 121.705 188.760 ;
        RECT 118.250 188.135 120.265 188.390 ;
        RECT 118.250 188.030 118.625 188.135 ;
        RECT 119.280 188.050 120.265 188.135 ;
        RECT 120.435 188.080 121.365 188.410 ;
        RECT 121.535 188.265 121.705 188.590 ;
        RECT 121.885 188.500 122.255 188.830 ;
        RECT 122.435 188.590 122.985 188.760 ;
        RECT 122.435 188.265 122.605 188.590 ;
        RECT 123.155 188.410 123.325 189.115 ;
        RECT 124.235 189.010 124.565 189.115 ;
        RECT 123.495 188.840 124.065 188.945 ;
        RECT 124.735 188.840 125.705 188.945 ;
        RECT 123.495 188.560 125.705 188.840 ;
        RECT 125.875 188.635 126.045 189.115 ;
        RECT 128.595 189.790 128.765 190.410 ;
        RECT 129.755 190.400 130.005 190.750 ;
        RECT 131.315 190.740 131.485 191.350 ;
        RECT 132.455 191.310 133.465 191.480 ;
        RECT 133.635 191.330 134.205 191.710 ;
        RECT 134.375 191.520 134.945 191.750 ;
        RECT 136.415 191.630 136.585 192.640 ;
        RECT 132.795 191.205 133.125 191.310 ;
        RECT 131.655 191.035 132.625 191.140 ;
        RECT 133.360 191.035 133.705 191.140 ;
        RECT 131.655 190.865 133.705 191.035 ;
        RECT 130.175 190.690 131.485 190.740 ;
        RECT 134.035 190.690 134.205 191.330 ;
        RECT 134.375 191.030 134.945 191.350 ;
        RECT 135.115 191.200 135.445 191.605 ;
        RECT 135.615 191.380 136.585 191.630 ;
        RECT 136.755 192.480 136.925 192.980 ;
        RECT 137.095 192.735 139.110 192.990 ;
        RECT 137.095 192.650 138.080 192.735 ;
        RECT 138.735 192.630 139.110 192.735 ;
        RECT 138.235 192.480 138.565 192.565 ;
        RECT 136.755 192.070 137.355 192.480 ;
        RECT 137.525 192.215 138.565 192.480 ;
        RECT 139.475 192.365 139.645 193.160 ;
        RECT 139.925 192.535 140.095 193.150 ;
        RECT 140.265 193.025 140.595 193.170 ;
        RECT 140.265 192.705 141.555 193.025 ;
        RECT 141.725 192.535 141.895 193.250 ;
        RECT 139.925 192.365 141.895 192.535 ;
        RECT 142.195 193.160 143.530 193.450 ;
        RECT 144.190 193.160 145.810 193.450 ;
        RECT 146.470 193.160 147.805 193.450 ;
        RECT 142.195 192.375 142.365 193.160 ;
        RECT 142.535 192.680 144.735 192.990 ;
        RECT 142.535 192.550 143.165 192.680 ;
        RECT 144.175 192.550 144.735 192.680 ;
        RECT 135.615 191.030 135.785 191.380 ;
        RECT 136.755 191.325 136.925 192.070 ;
        RECT 136.755 191.200 137.345 191.325 ;
        RECT 134.375 190.860 135.785 191.030 ;
        RECT 135.955 190.995 137.345 191.200 ;
        RECT 137.525 191.205 137.695 192.215 ;
        RECT 138.735 192.195 139.645 192.365 ;
        RECT 139.475 192.090 139.645 192.195 ;
        RECT 137.865 191.545 138.035 192.000 ;
        RECT 138.235 191.715 138.565 192.045 ;
        RECT 138.735 191.745 139.110 191.915 ;
        RECT 139.475 191.880 140.175 192.090 ;
        RECT 138.735 191.545 138.905 191.745 ;
        RECT 137.865 191.375 138.905 191.545 ;
        RECT 137.525 191.035 139.305 191.205 ;
        RECT 139.475 191.120 139.645 191.880 ;
        RECT 140.555 191.660 140.885 192.365 ;
        RECT 141.090 191.640 141.465 192.195 ;
        RECT 142.195 192.185 143.215 192.375 ;
        RECT 141.695 192.060 143.215 192.185 ;
        RECT 143.385 192.340 144.005 192.510 ;
        RECT 144.915 192.380 145.085 193.160 ;
        RECT 141.695 191.870 142.365 192.060 ;
        RECT 143.385 191.890 143.555 192.340 ;
        RECT 139.860 191.490 140.385 191.620 ;
        RECT 141.090 191.490 142.025 191.640 ;
        RECT 139.860 191.300 142.025 191.490 ;
        RECT 139.860 191.290 140.885 191.300 ;
        RECT 135.955 190.870 136.925 190.995 ;
        RECT 130.175 190.410 132.575 190.690 ;
        RECT 128.935 189.970 129.485 190.140 ;
        RECT 128.595 189.460 129.145 189.790 ;
        RECT 129.315 189.645 129.485 189.970 ;
        RECT 129.665 189.870 130.035 190.210 ;
        RECT 130.215 189.970 131.145 190.150 ;
        RECT 130.215 189.645 130.385 189.970 ;
        RECT 131.315 189.790 132.575 190.410 ;
        RECT 129.315 189.475 130.385 189.645 ;
        RECT 121.535 188.095 122.605 188.265 ;
        RECT 117.255 187.765 117.885 187.880 ;
        RECT 118.795 187.880 119.125 187.965 ;
        RECT 120.435 187.880 120.605 188.080 ;
        RECT 121.850 187.980 122.180 188.095 ;
        RECT 122.775 188.080 123.325 188.410 ;
        RECT 117.255 187.710 118.625 187.765 ;
        RECT 117.715 187.595 118.625 187.710 ;
        RECT 118.795 187.615 119.835 187.880 ;
        RECT 113.665 186.695 113.835 186.710 ;
        RECT 112.775 186.525 113.835 186.695 ;
        RECT 112.275 185.770 112.940 186.165 ;
        RECT 113.305 186.135 113.835 186.525 ;
        RECT 112.275 184.710 112.445 185.770 ;
        RECT 113.305 185.710 113.685 186.135 ;
        RECT 114.005 185.840 114.315 186.535 ;
        RECT 114.995 186.530 115.940 186.960 ;
        RECT 114.525 186.250 115.940 186.530 ;
        RECT 116.110 186.595 116.325 187.130 ;
        RECT 116.495 186.780 116.725 187.250 ;
        RECT 116.895 187.210 117.165 187.540 ;
        RECT 117.280 187.075 117.545 187.080 ;
        RECT 117.275 187.070 117.545 187.075 ;
        RECT 117.265 187.065 117.545 187.070 ;
        RECT 117.260 187.060 117.545 187.065 ;
        RECT 117.250 187.055 117.545 187.060 ;
        RECT 117.245 187.045 117.545 187.055 ;
        RECT 117.235 187.035 117.545 187.045 ;
        RECT 117.225 187.020 117.545 187.035 ;
        RECT 116.895 186.720 117.545 187.020 ;
        RECT 116.895 186.595 117.085 186.720 ;
        RECT 116.110 186.310 117.085 186.595 ;
        RECT 117.715 186.480 117.885 187.595 ;
        RECT 118.250 187.145 118.625 187.315 ;
        RECT 118.455 186.945 118.625 187.145 ;
        RECT 118.795 187.115 119.125 187.445 ;
        RECT 119.325 186.945 119.495 187.400 ;
        RECT 118.455 186.775 119.495 186.945 ;
        RECT 119.665 186.605 119.835 187.615 ;
        RECT 120.005 187.470 120.605 187.880 ;
        RECT 120.775 187.810 121.680 187.910 ;
        RECT 122.480 187.810 122.985 187.900 ;
        RECT 120.775 187.640 122.985 187.810 ;
        RECT 123.155 187.780 123.325 188.080 ;
        RECT 123.505 188.080 125.705 188.390 ;
        RECT 123.505 187.950 124.065 188.080 ;
        RECT 125.075 187.950 125.705 188.080 ;
        RECT 125.875 188.305 127.145 188.635 ;
        RECT 120.435 186.990 120.605 187.470 ;
        RECT 120.775 187.300 122.825 187.470 ;
        RECT 120.775 187.200 121.745 187.300 ;
        RECT 122.480 187.200 122.825 187.300 ;
        RECT 123.155 187.330 124.065 187.780 ;
        RECT 124.235 187.740 124.855 187.910 ;
        RECT 125.875 187.775 126.045 188.305 ;
        RECT 127.395 188.205 127.605 188.850 ;
        RECT 127.775 188.365 128.410 188.695 ;
        RECT 121.915 187.030 122.245 187.130 ;
        RECT 120.435 186.725 121.405 186.990 ;
        RECT 117.255 186.310 117.885 186.480 ;
        RECT 118.055 186.435 119.835 186.605 ;
        RECT 114.525 185.845 115.165 186.250 ;
        RECT 116.770 186.080 117.545 186.140 ;
        RECT 112.615 185.535 113.135 185.600 ;
        RECT 113.940 185.535 114.725 185.665 ;
        RECT 112.615 185.360 114.725 185.535 ;
        RECT 114.995 184.710 115.165 185.845 ;
        RECT 115.335 185.800 117.545 186.080 ;
        RECT 117.715 185.705 117.885 186.310 ;
        RECT 118.055 185.875 118.705 186.205 ;
        RECT 117.715 185.535 118.355 185.705 ;
        RECT 117.715 184.710 117.885 185.535 ;
        RECT 118.535 185.365 118.705 185.875 ;
        RECT 118.875 185.695 119.085 186.265 ;
        RECT 119.255 186.225 119.835 186.435 ;
        RECT 120.015 186.710 121.405 186.725 ;
        RECT 121.575 186.860 122.585 187.030 ;
        RECT 123.155 187.010 123.325 187.330 ;
        RECT 124.235 187.180 124.515 187.570 ;
        RECT 124.685 187.290 124.855 187.740 ;
        RECT 125.025 187.460 126.045 187.775 ;
        RECT 126.215 187.505 127.225 187.830 ;
        RECT 125.875 187.335 126.045 187.460 ;
        RECT 120.015 186.395 120.605 186.710 ;
        RECT 119.255 185.900 120.265 186.225 ;
        RECT 118.070 185.035 118.705 185.365 ;
        RECT 118.875 184.880 119.085 185.525 ;
        RECT 120.435 185.425 120.605 186.395 ;
        RECT 119.335 185.095 120.605 185.425 ;
        RECT 120.435 184.710 120.605 185.095 ;
        RECT 120.825 184.885 121.115 186.540 ;
        RECT 121.575 186.475 121.745 186.860 ;
        RECT 121.285 186.305 121.745 186.475 ;
        RECT 121.285 185.205 121.455 186.305 ;
        RECT 121.915 186.285 122.245 186.690 ;
        RECT 122.415 186.460 122.585 186.860 ;
        RECT 122.755 186.820 123.325 187.010 ;
        RECT 123.495 186.990 124.065 187.160 ;
        RECT 124.685 187.120 125.705 187.290 ;
        RECT 122.755 186.630 123.725 186.820 ;
        RECT 122.415 186.290 122.935 186.460 ;
        RECT 123.155 186.400 123.725 186.630 ;
        RECT 121.625 185.405 122.245 186.115 ;
        RECT 122.415 185.590 122.585 186.290 ;
        RECT 123.155 186.120 123.325 186.400 ;
        RECT 123.895 186.230 124.065 186.990 ;
        RECT 124.235 186.950 124.565 186.995 ;
        RECT 124.235 186.750 125.365 186.950 ;
        RECT 124.235 186.300 125.365 186.550 ;
        RECT 122.755 185.790 123.325 186.120 ;
        RECT 123.495 186.000 124.065 186.230 ;
        RECT 125.535 186.110 125.705 187.120 ;
        RECT 122.415 185.420 122.935 185.590 ;
        RECT 121.285 184.885 121.745 185.205 ;
        RECT 121.915 184.885 122.485 185.235 ;
        RECT 123.155 185.220 123.325 185.790 ;
        RECT 123.495 185.510 124.065 185.830 ;
        RECT 124.235 185.680 124.565 186.085 ;
        RECT 124.735 185.860 125.705 186.110 ;
        RECT 125.875 187.005 126.465 187.335 ;
        RECT 126.645 187.295 127.225 187.505 ;
        RECT 127.395 187.465 127.605 188.035 ;
        RECT 127.775 187.855 127.945 188.365 ;
        RECT 128.595 188.195 128.765 189.460 ;
        RECT 129.740 189.370 130.070 189.475 ;
        RECT 130.555 189.460 132.575 189.790 ;
        RECT 132.745 190.670 134.205 190.690 ;
        RECT 132.745 190.430 135.015 190.670 ;
        RECT 132.745 189.760 134.205 190.430 ;
        RECT 135.195 190.340 135.445 190.690 ;
        RECT 135.615 190.350 136.570 190.680 ;
        RECT 134.375 190.170 135.015 190.260 ;
        RECT 135.615 190.170 135.785 190.350 ;
        RECT 134.375 190.000 135.785 190.170 ;
        RECT 136.755 190.025 136.925 190.870 ;
        RECT 137.525 190.825 138.105 191.035 ;
        RECT 139.475 190.950 140.255 191.120 ;
        RECT 137.095 190.500 138.105 190.825 ;
        RECT 138.275 190.295 138.485 190.865 ;
        RECT 138.655 190.475 139.305 190.805 ;
        RECT 134.375 189.930 135.015 190.000 ;
        RECT 132.745 189.490 135.015 189.760 ;
        RECT 132.745 189.480 134.205 189.490 ;
        RECT 135.195 189.480 135.445 189.830 ;
        RECT 136.755 189.820 138.025 190.025 ;
        RECT 135.615 189.695 138.025 189.820 ;
        RECT 135.615 189.490 136.925 189.695 ;
        RECT 131.315 189.310 132.575 189.460 ;
        RECT 128.935 189.200 129.440 189.280 ;
        RECT 130.240 189.200 131.145 189.290 ;
        RECT 128.935 189.020 131.145 189.200 ;
        RECT 128.950 188.365 129.585 188.695 ;
        RECT 128.125 188.025 129.235 188.195 ;
        RECT 127.775 187.525 128.425 187.855 ;
        RECT 126.645 187.125 128.425 187.295 ;
        RECT 125.875 186.260 126.045 187.005 ;
        RECT 124.735 185.510 124.905 185.860 ;
        RECT 125.875 185.850 126.475 186.260 ;
        RECT 126.645 186.115 126.815 187.125 ;
        RECT 126.985 186.785 128.025 186.955 ;
        RECT 126.985 186.330 127.155 186.785 ;
        RECT 127.355 186.285 127.685 186.615 ;
        RECT 127.855 186.585 128.025 186.785 ;
        RECT 127.855 186.415 128.230 186.585 ;
        RECT 128.595 186.135 128.765 188.025 ;
        RECT 129.415 187.855 129.585 188.365 ;
        RECT 129.755 188.205 129.965 188.850 ;
        RECT 131.315 188.635 133.095 189.310 ;
        RECT 130.215 188.305 133.095 188.635 ;
        RECT 131.315 188.100 133.095 188.305 ;
        RECT 133.265 188.225 134.205 189.480 ;
        RECT 134.570 188.595 136.585 188.850 ;
        RECT 134.570 188.490 134.945 188.595 ;
        RECT 135.600 188.510 136.585 188.595 ;
        RECT 136.755 188.800 136.925 189.490 ;
        RECT 138.275 189.480 138.485 190.125 ;
        RECT 138.655 189.965 138.825 190.475 ;
        RECT 139.475 190.305 139.645 190.950 ;
        RECT 139.865 190.625 140.385 190.780 ;
        RECT 140.555 190.740 140.885 191.290 ;
        RECT 142.195 191.130 142.365 191.870 ;
        RECT 141.185 190.960 142.365 191.130 ;
        RECT 139.865 190.570 140.425 190.625 ;
        RECT 141.055 190.615 141.980 190.790 ;
        RECT 141.005 190.570 141.980 190.615 ;
        RECT 139.865 190.460 141.980 190.570 ;
        RECT 139.865 190.450 141.135 190.460 ;
        RECT 140.300 190.400 141.135 190.450 ;
        RECT 139.005 190.135 139.645 190.305 ;
        RECT 138.655 189.635 139.290 189.965 ;
        RECT 139.475 189.605 139.645 190.135 ;
        RECT 142.195 190.280 142.365 190.960 ;
        RECT 142.535 191.720 143.555 191.890 ;
        RECT 143.725 191.780 144.005 192.170 ;
        RECT 144.175 192.065 145.085 192.380 ;
        RECT 147.635 192.065 147.805 193.160 ;
        RECT 144.175 191.930 145.925 192.065 ;
        RECT 144.915 191.805 145.925 191.930 ;
        RECT 146.485 191.805 147.805 192.065 ;
        RECT 142.535 190.710 142.705 191.720 ;
        RECT 143.675 191.550 144.005 191.595 ;
        RECT 142.875 191.350 144.005 191.550 ;
        RECT 144.175 191.590 144.745 191.760 ;
        RECT 142.875 190.900 144.005 191.150 ;
        RECT 144.175 190.830 144.345 191.590 ;
        RECT 144.915 191.420 145.085 191.805 ;
        RECT 144.515 191.205 145.085 191.420 ;
        RECT 145.255 191.460 147.465 191.630 ;
        RECT 145.255 191.375 145.830 191.460 ;
        RECT 146.560 191.375 147.465 191.460 ;
        RECT 145.995 191.205 146.325 191.290 ;
        RECT 147.635 191.205 147.805 191.805 ;
        RECT 144.515 191.000 145.465 191.205 ;
        RECT 144.915 190.875 145.465 191.000 ;
        RECT 145.635 191.035 146.705 191.205 ;
        RECT 142.535 190.460 143.505 190.710 ;
        RECT 142.195 189.950 143.165 190.280 ;
        RECT 143.335 190.110 143.505 190.460 ;
        RECT 143.675 190.280 144.005 190.685 ;
        RECT 144.175 190.600 144.745 190.830 ;
        RECT 144.175 190.110 144.745 190.430 ;
        RECT 139.475 189.365 140.155 189.605 ;
        RECT 137.095 189.055 139.110 189.310 ;
        RECT 137.095 188.970 138.080 189.055 ;
        RECT 138.735 188.950 139.110 189.055 ;
        RECT 138.235 188.800 138.565 188.885 ;
        RECT 135.115 188.340 135.445 188.425 ;
        RECT 136.755 188.390 137.355 188.800 ;
        RECT 137.525 188.535 138.565 188.800 ;
        RECT 139.475 188.685 139.645 189.365 ;
        RECT 140.325 189.355 140.885 189.710 ;
        RECT 141.055 189.195 141.400 189.585 ;
        RECT 142.195 189.200 142.365 189.950 ;
        RECT 143.335 189.940 144.745 190.110 ;
        RECT 144.915 190.230 145.085 190.875 ;
        RECT 145.635 190.660 145.805 191.035 ;
        RECT 145.255 190.490 145.805 190.660 ;
        RECT 145.985 190.400 146.355 190.755 ;
        RECT 146.535 190.660 146.705 191.035 ;
        RECT 146.875 190.875 147.805 191.205 ;
        RECT 146.535 190.490 147.465 190.660 ;
        RECT 147.635 190.230 147.805 190.875 ;
        RECT 142.535 189.370 143.215 189.655 ;
        RECT 141.055 189.185 141.225 189.195 ;
        RECT 139.825 189.015 141.225 189.185 ;
        RECT 139.825 188.905 140.155 189.015 ;
        RECT 138.735 188.675 139.645 188.685 ;
        RECT 136.755 188.340 136.925 188.390 ;
        RECT 133.265 188.100 134.945 188.225 ;
        RECT 128.935 187.525 129.585 187.855 ;
        RECT 129.755 187.465 129.965 188.035 ;
        RECT 130.135 187.505 131.145 187.830 ;
        RECT 130.135 187.295 130.715 187.505 ;
        RECT 131.315 187.460 131.485 188.100 ;
        RECT 134.035 188.055 134.945 188.100 ;
        RECT 135.115 188.075 136.155 188.340 ;
        RECT 131.315 187.335 132.625 187.460 ;
        RECT 128.935 187.125 130.715 187.295 ;
        RECT 129.335 186.785 130.375 186.955 ;
        RECT 129.335 186.585 129.505 186.785 ;
        RECT 129.130 186.415 129.505 186.585 ;
        RECT 129.675 186.285 130.005 186.615 ;
        RECT 130.205 186.330 130.375 186.785 ;
        RECT 126.645 185.850 127.685 186.115 ;
        RECT 127.855 185.965 129.505 186.135 ;
        RECT 130.545 186.115 130.715 187.125 ;
        RECT 130.895 187.130 132.625 187.335 ;
        RECT 130.895 187.005 131.485 187.130 ;
        RECT 132.795 187.120 133.045 187.470 ;
        RECT 134.035 187.460 134.205 188.055 ;
        RECT 134.570 187.605 134.945 187.775 ;
        RECT 133.225 187.190 134.205 187.460 ;
        RECT 134.775 187.405 134.945 187.605 ;
        RECT 135.115 187.575 135.445 187.905 ;
        RECT 135.645 187.405 135.815 187.860 ;
        RECT 134.775 187.235 135.815 187.405 ;
        RECT 131.315 186.260 131.485 187.005 ;
        RECT 133.225 186.950 133.865 187.020 ;
        RECT 132.455 186.780 133.865 186.950 ;
        RECT 132.455 186.600 132.625 186.780 ;
        RECT 133.225 186.690 133.865 186.780 ;
        RECT 131.670 186.270 132.625 186.600 ;
        RECT 132.795 186.260 133.045 186.610 ;
        RECT 134.035 186.520 134.205 187.190 ;
        RECT 135.985 187.065 136.155 188.075 ;
        RECT 136.325 187.930 136.925 188.340 ;
        RECT 136.755 187.645 136.925 187.930 ;
        RECT 136.755 187.315 137.345 187.645 ;
        RECT 137.525 187.525 137.695 188.535 ;
        RECT 138.735 188.515 140.155 188.675 ;
        RECT 140.325 188.580 140.885 188.845 ;
        RECT 139.475 188.460 140.155 188.515 ;
        RECT 137.865 187.865 138.035 188.320 ;
        RECT 138.235 188.035 138.565 188.365 ;
        RECT 138.735 188.065 139.110 188.235 ;
        RECT 138.735 187.865 138.905 188.065 ;
        RECT 137.865 187.695 138.905 187.865 ;
        RECT 137.525 187.355 139.305 187.525 ;
        RECT 136.755 187.185 136.925 187.315 ;
        RECT 134.375 186.895 136.155 187.065 ;
        RECT 133.225 186.280 134.205 186.520 ;
        RECT 134.375 186.335 135.025 186.665 ;
        RECT 125.875 185.680 126.045 185.850 ;
        RECT 127.355 185.765 127.685 185.850 ;
        RECT 123.495 185.340 124.905 185.510 ;
        RECT 125.075 185.350 126.045 185.680 ;
        RECT 122.655 184.890 123.325 185.220 ;
        RECT 123.155 184.710 123.325 184.890 ;
        RECT 125.875 184.710 126.045 185.350 ;
        RECT 126.215 185.595 127.200 185.680 ;
        RECT 127.855 185.595 128.230 185.700 ;
        RECT 126.215 185.570 128.230 185.595 ;
        RECT 126.215 185.400 128.255 185.570 ;
        RECT 126.215 185.340 128.230 185.400 ;
        RECT 128.595 184.710 128.765 185.965 ;
        RECT 129.675 185.850 130.715 186.115 ;
        RECT 130.885 185.850 131.485 186.260 ;
        RECT 134.035 186.165 134.205 186.280 ;
        RECT 129.675 185.765 130.005 185.850 ;
        RECT 129.130 185.595 129.505 185.700 ;
        RECT 130.160 185.595 131.145 185.680 ;
        RECT 129.130 185.340 131.145 185.595 ;
        RECT 131.315 185.650 131.485 185.850 ;
        RECT 131.655 185.920 133.865 186.090 ;
        RECT 131.655 185.820 132.560 185.920 ;
        RECT 133.360 185.830 133.865 185.920 ;
        RECT 134.035 185.995 134.675 186.165 ;
        RECT 131.315 185.320 132.245 185.650 ;
        RECT 132.730 185.635 133.060 185.750 ;
        RECT 134.035 185.650 134.205 185.995 ;
        RECT 134.855 185.825 135.025 186.335 ;
        RECT 135.195 186.155 135.405 186.725 ;
        RECT 135.575 186.685 136.155 186.895 ;
        RECT 136.335 186.855 136.925 187.185 ;
        RECT 137.525 187.145 138.105 187.355 ;
        RECT 135.575 186.360 136.585 186.685 ;
        RECT 136.755 186.345 136.925 186.855 ;
        RECT 137.095 186.820 138.105 187.145 ;
        RECT 138.275 186.615 138.485 187.185 ;
        RECT 138.655 186.795 139.305 187.125 ;
        RECT 139.475 187.030 139.645 188.460 ;
        RECT 141.055 188.330 141.225 189.015 ;
        RECT 142.195 188.930 142.825 189.200 ;
        RECT 142.195 188.710 142.365 188.930 ;
        RECT 141.395 188.380 142.365 188.710 ;
        RECT 142.995 188.910 143.215 189.370 ;
        RECT 143.385 189.080 143.945 189.770 ;
        RECT 144.915 189.710 146.375 190.230 ;
        RECT 144.115 189.370 144.745 189.655 ;
        RECT 144.115 188.910 144.285 189.370 ;
        RECT 144.915 189.200 145.835 189.710 ;
        RECT 146.545 189.540 147.805 190.230 ;
        RECT 144.455 189.020 145.835 189.200 ;
        RECT 146.005 189.020 147.805 189.540 ;
        RECT 144.455 188.930 145.085 189.020 ;
        RECT 142.995 188.700 144.285 188.910 ;
        RECT 139.815 187.990 140.385 188.290 ;
        RECT 140.555 188.160 141.225 188.330 ;
        RECT 141.405 187.990 142.025 188.210 ;
        RECT 139.815 187.675 142.025 187.990 ;
        RECT 139.815 187.210 140.365 187.380 ;
        RECT 136.755 186.015 138.025 186.345 ;
        RECT 132.415 185.465 133.485 185.635 ;
        RECT 131.315 184.710 131.485 185.320 ;
        RECT 132.415 185.140 132.585 185.465 ;
        RECT 131.655 184.970 132.585 185.140 ;
        RECT 132.765 184.900 133.135 185.230 ;
        RECT 133.315 185.140 133.485 185.465 ;
        RECT 133.655 185.320 134.205 185.650 ;
        RECT 134.390 185.495 135.025 185.825 ;
        RECT 135.195 185.340 135.405 185.985 ;
        RECT 136.755 185.885 136.925 186.015 ;
        RECT 135.655 185.555 136.925 185.885 ;
        RECT 138.275 185.800 138.485 186.445 ;
        RECT 138.655 186.285 138.825 186.795 ;
        RECT 139.475 186.700 140.025 187.030 ;
        RECT 140.195 186.885 140.365 187.210 ;
        RECT 140.545 187.120 140.915 187.450 ;
        RECT 141.095 187.210 142.025 187.380 ;
        RECT 141.095 186.885 141.265 187.210 ;
        RECT 142.195 187.140 142.365 188.380 ;
        RECT 142.535 188.130 144.745 188.530 ;
        RECT 144.915 188.410 145.085 188.930 ;
        RECT 145.255 188.680 147.465 188.850 ;
        RECT 145.255 188.590 145.760 188.680 ;
        RECT 146.560 188.580 147.465 188.680 ;
        RECT 142.535 187.660 143.215 187.940 ;
        RECT 142.995 187.265 143.215 187.660 ;
        RECT 143.385 187.435 143.945 188.130 ;
        RECT 144.915 188.080 145.465 188.410 ;
        RECT 146.060 188.395 146.390 188.510 ;
        RECT 147.635 188.410 147.805 189.020 ;
        RECT 145.635 188.225 146.705 188.395 ;
        RECT 144.115 187.660 144.745 187.940 ;
        RECT 144.115 187.265 144.285 187.660 ;
        RECT 142.195 187.030 142.825 187.140 ;
        RECT 140.195 186.715 141.265 186.885 ;
        RECT 141.435 186.815 142.825 187.030 ;
        RECT 142.995 186.815 144.285 187.265 ;
        RECT 144.915 187.140 145.085 188.080 ;
        RECT 145.635 187.900 145.805 188.225 ;
        RECT 145.255 187.730 145.805 187.900 ;
        RECT 145.985 187.660 146.355 187.990 ;
        RECT 146.535 187.900 146.705 188.225 ;
        RECT 146.875 188.080 147.805 188.410 ;
        RECT 146.535 187.730 147.465 187.900 ;
        RECT 145.255 187.300 147.465 187.470 ;
        RECT 145.255 187.210 145.760 187.300 ;
        RECT 146.560 187.200 147.465 187.300 ;
        RECT 144.455 187.030 145.085 187.140 ;
        RECT 144.455 186.815 145.465 187.030 ;
        RECT 146.060 187.015 146.390 187.130 ;
        RECT 147.635 187.030 147.805 188.080 ;
        RECT 139.475 186.625 139.645 186.700 ;
        RECT 139.005 186.455 139.645 186.625 ;
        RECT 140.620 186.600 140.950 186.715 ;
        RECT 141.435 186.700 142.365 186.815 ;
        RECT 143.675 186.710 144.005 186.815 ;
        RECT 138.655 185.955 139.290 186.285 ;
        RECT 133.315 184.970 133.865 185.140 ;
        RECT 134.035 184.710 134.205 185.320 ;
        RECT 136.755 184.710 136.925 185.555 ;
        RECT 139.475 185.650 139.645 186.455 ;
        RECT 139.815 186.430 140.320 186.520 ;
        RECT 141.120 186.430 142.025 186.530 ;
        RECT 139.815 186.260 142.025 186.430 ;
        RECT 139.815 185.910 142.025 186.090 ;
        RECT 139.815 185.830 140.320 185.910 ;
        RECT 141.120 185.820 142.025 185.910 ;
        RECT 139.475 185.320 140.025 185.650 ;
        RECT 140.620 185.635 140.950 185.740 ;
        RECT 142.195 185.650 142.365 186.700 ;
        RECT 144.915 186.700 145.465 186.815 ;
        RECT 145.635 186.845 146.705 187.015 ;
        RECT 142.535 186.540 143.505 186.645 ;
        RECT 144.175 186.540 144.745 186.645 ;
        RECT 142.535 186.260 144.745 186.540 ;
        RECT 142.535 185.910 144.745 186.090 ;
        RECT 142.535 185.820 143.440 185.910 ;
        RECT 144.240 185.830 144.745 185.910 ;
        RECT 140.195 185.465 141.265 185.635 ;
        RECT 139.475 184.710 139.645 185.320 ;
        RECT 140.195 185.140 140.365 185.465 ;
        RECT 139.815 184.970 140.365 185.140 ;
        RECT 140.545 184.900 140.915 185.240 ;
        RECT 141.095 185.140 141.265 185.465 ;
        RECT 141.435 185.320 143.125 185.650 ;
        RECT 143.610 185.635 143.940 185.740 ;
        RECT 144.915 185.650 145.085 186.700 ;
        RECT 145.635 186.520 145.805 186.845 ;
        RECT 145.255 186.350 145.805 186.520 ;
        RECT 145.985 186.280 146.355 186.610 ;
        RECT 146.535 186.520 146.705 186.845 ;
        RECT 146.875 186.700 147.805 187.030 ;
        RECT 146.535 186.350 147.465 186.520 ;
        RECT 145.255 185.910 147.465 186.090 ;
        RECT 145.255 185.830 145.760 185.910 ;
        RECT 146.560 185.820 147.465 185.910 ;
        RECT 143.295 185.465 144.365 185.635 ;
        RECT 141.095 184.960 142.025 185.140 ;
        RECT 142.195 184.710 142.365 185.320 ;
        RECT 143.295 185.140 143.465 185.465 ;
        RECT 142.535 184.960 143.465 185.140 ;
        RECT 143.645 184.900 144.015 185.240 ;
        RECT 144.195 185.140 144.365 185.465 ;
        RECT 144.535 185.320 145.465 185.650 ;
        RECT 146.060 185.635 146.390 185.740 ;
        RECT 147.635 185.650 147.805 186.700 ;
        RECT 145.635 185.465 146.705 185.635 ;
        RECT 144.195 184.970 144.745 185.140 ;
        RECT 144.915 184.710 145.085 185.320 ;
        RECT 145.635 185.140 145.805 185.465 ;
        RECT 145.255 184.970 145.805 185.140 ;
        RECT 145.985 184.900 146.355 185.240 ;
        RECT 146.535 185.140 146.705 185.465 ;
        RECT 146.875 185.320 147.805 185.650 ;
        RECT 146.535 184.960 147.465 185.140 ;
        RECT 147.635 184.710 147.805 185.320 ;
        RECT 112.275 184.020 113.195 184.710 ;
        RECT 113.365 184.190 116.795 184.710 ;
        RECT 112.275 183.500 113.735 184.020 ;
        RECT 113.905 183.500 116.255 184.190 ;
        RECT 116.965 184.020 118.635 184.710 ;
        RECT 118.805 184.190 122.235 184.710 ;
        RECT 116.425 183.500 119.175 184.020 ;
        RECT 119.345 183.500 121.695 184.190 ;
        RECT 122.405 184.020 124.075 184.710 ;
        RECT 124.245 184.190 127.675 184.710 ;
        RECT 121.865 183.500 124.615 184.020 ;
        RECT 124.785 183.500 127.135 184.190 ;
        RECT 127.845 184.020 129.515 184.710 ;
        RECT 129.685 184.190 133.115 184.710 ;
        RECT 127.305 183.500 130.055 184.020 ;
        RECT 130.225 183.500 132.575 184.190 ;
        RECT 133.285 184.020 134.955 184.710 ;
        RECT 135.125 184.190 138.555 184.710 ;
        RECT 132.745 183.500 135.495 184.020 ;
        RECT 135.665 183.500 138.015 184.190 ;
        RECT 138.725 184.020 140.395 184.710 ;
        RECT 140.565 184.190 143.995 184.710 ;
        RECT 138.185 183.500 140.935 184.020 ;
        RECT 141.105 183.500 143.455 184.190 ;
        RECT 144.165 184.020 145.835 184.710 ;
        RECT 146.005 184.190 147.805 184.710 ;
        RECT 143.625 183.500 146.375 184.020 ;
        RECT 146.545 183.500 147.805 184.190 ;
        RECT 112.275 183.415 112.445 183.500 ;
        RECT 114.995 183.415 115.165 183.500 ;
        RECT 117.715 183.415 117.885 183.500 ;
        RECT 120.435 183.415 120.605 183.500 ;
        RECT 123.155 183.415 123.325 183.500 ;
        RECT 125.875 183.415 126.045 183.500 ;
        RECT 128.595 183.415 128.765 183.500 ;
        RECT 131.315 183.415 131.485 183.500 ;
        RECT 134.035 183.415 134.205 183.500 ;
        RECT 136.755 183.415 136.925 183.500 ;
        RECT 139.475 183.415 139.645 183.500 ;
        RECT 142.195 183.415 142.365 183.500 ;
        RECT 144.915 183.415 145.085 183.500 ;
        RECT 147.635 183.415 147.805 183.500 ;
        RECT 100.630 176.790 106.370 176.800 ;
        RECT 100.140 176.630 106.370 176.790 ;
        RECT 100.140 174.370 100.810 176.630 ;
        RECT 101.480 176.060 105.520 176.230 ;
        RECT 101.140 175.000 101.310 176.000 ;
        RECT 105.690 175.000 105.860 176.000 ;
        RECT 101.480 174.770 105.520 174.940 ;
        RECT 106.200 174.370 106.370 176.630 ;
        RECT 100.140 174.200 106.370 174.370 ;
        RECT 12.100 173.775 89.840 173.945 ;
        RECT 12.185 172.685 13.395 173.775 ;
        RECT 13.565 173.340 18.910 173.775 ;
        RECT 19.085 173.340 24.430 173.775 ;
        RECT 12.185 171.975 12.705 172.515 ;
        RECT 12.875 172.145 13.395 172.685 ;
        RECT 12.185 171.225 13.395 171.975 ;
        RECT 15.150 171.770 15.490 172.600 ;
        RECT 16.970 172.090 17.320 173.340 ;
        RECT 20.670 171.770 21.010 172.600 ;
        RECT 22.490 172.090 22.840 173.340 ;
        RECT 25.065 172.610 25.355 173.775 ;
        RECT 25.525 173.340 30.870 173.775 ;
        RECT 31.045 173.340 36.390 173.775 ;
        RECT 13.565 171.225 18.910 171.770 ;
        RECT 19.085 171.225 24.430 171.770 ;
        RECT 25.065 171.225 25.355 171.950 ;
        RECT 27.110 171.770 27.450 172.600 ;
        RECT 28.930 172.090 29.280 173.340 ;
        RECT 32.630 171.770 32.970 172.600 ;
        RECT 34.450 172.090 34.800 173.340 ;
        RECT 36.565 172.685 37.775 173.775 ;
        RECT 36.565 171.975 37.085 172.515 ;
        RECT 37.255 172.145 37.775 172.685 ;
        RECT 37.945 172.610 38.235 173.775 ;
        RECT 38.405 173.340 43.750 173.775 ;
        RECT 25.525 171.225 30.870 171.770 ;
        RECT 31.045 171.225 36.390 171.770 ;
        RECT 36.565 171.225 37.775 171.975 ;
        RECT 37.945 171.225 38.235 171.950 ;
        RECT 39.990 171.770 40.330 172.600 ;
        RECT 41.810 172.090 42.160 173.340 ;
        RECT 43.925 172.685 45.595 173.775 ;
        RECT 43.925 171.995 44.675 172.515 ;
        RECT 44.845 172.165 45.595 172.685 ;
        RECT 45.770 172.625 46.030 173.775 ;
        RECT 46.205 172.700 46.460 173.605 ;
        RECT 46.630 173.015 46.960 173.775 ;
        RECT 47.175 172.845 47.345 173.605 ;
        RECT 38.405 171.225 43.750 171.770 ;
        RECT 43.925 171.225 45.595 171.995 ;
        RECT 45.770 171.225 46.030 172.065 ;
        RECT 46.205 171.970 46.375 172.700 ;
        RECT 46.630 172.675 47.345 172.845 ;
        RECT 47.605 172.685 50.195 173.775 ;
        RECT 46.630 172.465 46.800 172.675 ;
        RECT 46.545 172.135 46.800 172.465 ;
        RECT 46.205 171.395 46.460 171.970 ;
        RECT 46.630 171.945 46.800 172.135 ;
        RECT 47.080 172.125 47.435 172.495 ;
        RECT 47.605 171.995 48.815 172.515 ;
        RECT 48.985 172.165 50.195 172.685 ;
        RECT 50.825 172.610 51.115 173.775 ;
        RECT 51.285 173.340 56.630 173.775 ;
        RECT 46.630 171.775 47.345 171.945 ;
        RECT 46.630 171.225 46.960 171.605 ;
        RECT 47.175 171.395 47.345 171.775 ;
        RECT 47.605 171.225 50.195 171.995 ;
        RECT 50.825 171.225 51.115 171.950 ;
        RECT 52.870 171.770 53.210 172.600 ;
        RECT 54.690 172.090 55.040 173.340 ;
        RECT 56.805 172.685 58.015 173.775 ;
        RECT 56.805 171.975 57.325 172.515 ;
        RECT 57.495 172.145 58.015 172.685 ;
        RECT 58.190 172.625 58.450 173.775 ;
        RECT 58.625 172.700 58.880 173.605 ;
        RECT 59.050 173.015 59.380 173.775 ;
        RECT 59.595 172.845 59.765 173.605 ;
        RECT 51.285 171.225 56.630 171.770 ;
        RECT 56.805 171.225 58.015 171.975 ;
        RECT 58.190 171.225 58.450 172.065 ;
        RECT 58.625 171.970 58.795 172.700 ;
        RECT 59.050 172.675 59.765 172.845 ;
        RECT 59.050 172.465 59.220 172.675 ;
        RECT 60.030 172.625 60.290 173.775 ;
        RECT 60.465 172.700 60.720 173.605 ;
        RECT 60.890 173.015 61.220 173.775 ;
        RECT 61.435 172.845 61.605 173.605 ;
        RECT 58.965 172.135 59.220 172.465 ;
        RECT 58.625 171.395 58.880 171.970 ;
        RECT 59.050 171.945 59.220 172.135 ;
        RECT 59.500 172.125 59.855 172.495 ;
        RECT 59.050 171.775 59.765 171.945 ;
        RECT 59.050 171.225 59.380 171.605 ;
        RECT 59.595 171.395 59.765 171.775 ;
        RECT 60.030 171.225 60.290 172.065 ;
        RECT 60.465 171.970 60.635 172.700 ;
        RECT 60.890 172.675 61.605 172.845 ;
        RECT 60.890 172.465 61.060 172.675 ;
        RECT 61.870 172.625 62.130 173.775 ;
        RECT 62.305 172.700 62.560 173.605 ;
        RECT 62.730 173.015 63.060 173.775 ;
        RECT 63.275 172.845 63.445 173.605 ;
        RECT 60.805 172.135 61.060 172.465 ;
        RECT 60.465 171.395 60.720 171.970 ;
        RECT 60.890 171.945 61.060 172.135 ;
        RECT 61.340 172.125 61.695 172.495 ;
        RECT 60.890 171.775 61.605 171.945 ;
        RECT 60.890 171.225 61.220 171.605 ;
        RECT 61.435 171.395 61.605 171.775 ;
        RECT 61.870 171.225 62.130 172.065 ;
        RECT 62.305 171.970 62.475 172.700 ;
        RECT 62.730 172.675 63.445 172.845 ;
        RECT 62.730 172.465 62.900 172.675 ;
        RECT 63.705 172.610 63.995 173.775 ;
        RECT 64.255 172.845 64.425 173.605 ;
        RECT 64.640 173.015 64.970 173.775 ;
        RECT 64.255 172.675 64.970 172.845 ;
        RECT 65.140 172.700 65.395 173.605 ;
        RECT 62.645 172.135 62.900 172.465 ;
        RECT 62.305 171.395 62.560 171.970 ;
        RECT 62.730 171.945 62.900 172.135 ;
        RECT 63.180 172.125 63.535 172.495 ;
        RECT 64.165 172.125 64.520 172.495 ;
        RECT 64.800 172.465 64.970 172.675 ;
        RECT 64.800 172.135 65.055 172.465 ;
        RECT 62.730 171.775 63.445 171.945 ;
        RECT 62.730 171.225 63.060 171.605 ;
        RECT 63.275 171.395 63.445 171.775 ;
        RECT 63.705 171.225 63.995 171.950 ;
        RECT 64.800 171.945 64.970 172.135 ;
        RECT 65.225 171.970 65.395 172.700 ;
        RECT 65.570 172.625 65.830 173.775 ;
        RECT 66.010 172.625 66.270 173.775 ;
        RECT 66.445 172.700 66.700 173.605 ;
        RECT 66.870 173.015 67.200 173.775 ;
        RECT 67.415 172.845 67.585 173.605 ;
        RECT 64.255 171.775 64.970 171.945 ;
        RECT 64.255 171.395 64.425 171.775 ;
        RECT 64.640 171.225 64.970 171.605 ;
        RECT 65.140 171.395 65.395 171.970 ;
        RECT 65.570 171.225 65.830 172.065 ;
        RECT 66.010 171.225 66.270 172.065 ;
        RECT 66.445 171.970 66.615 172.700 ;
        RECT 66.870 172.675 67.585 172.845 ;
        RECT 67.880 172.985 68.415 173.605 ;
        RECT 66.870 172.465 67.040 172.675 ;
        RECT 66.785 172.135 67.040 172.465 ;
        RECT 66.445 171.395 66.700 171.970 ;
        RECT 66.870 171.945 67.040 172.135 ;
        RECT 67.320 172.125 67.675 172.495 ;
        RECT 67.880 171.965 68.195 172.985 ;
        RECT 68.585 172.975 68.915 173.775 ;
        RECT 70.180 172.985 70.715 173.605 ;
        RECT 69.400 172.805 69.790 172.980 ;
        RECT 68.365 172.635 69.790 172.805 ;
        RECT 68.365 172.135 68.535 172.635 ;
        RECT 66.870 171.775 67.585 171.945 ;
        RECT 66.870 171.225 67.200 171.605 ;
        RECT 67.415 171.395 67.585 171.775 ;
        RECT 67.880 171.395 68.495 171.965 ;
        RECT 68.785 171.905 69.050 172.465 ;
        RECT 69.220 171.735 69.390 172.635 ;
        RECT 69.560 171.905 69.915 172.465 ;
        RECT 70.180 171.965 70.495 172.985 ;
        RECT 70.885 172.975 71.215 173.775 ;
        RECT 72.480 172.985 73.015 173.605 ;
        RECT 71.700 172.805 72.090 172.980 ;
        RECT 70.665 172.635 72.090 172.805 ;
        RECT 70.665 172.135 70.835 172.635 ;
        RECT 68.665 171.225 68.880 171.735 ;
        RECT 69.110 171.405 69.390 171.735 ;
        RECT 69.570 171.225 69.810 171.735 ;
        RECT 70.180 171.395 70.795 171.965 ;
        RECT 71.085 171.905 71.350 172.465 ;
        RECT 71.520 171.735 71.690 172.635 ;
        RECT 71.860 171.905 72.215 172.465 ;
        RECT 72.480 171.965 72.795 172.985 ;
        RECT 73.185 172.975 73.515 173.775 ;
        RECT 74.000 172.805 74.390 172.980 ;
        RECT 72.965 172.635 74.390 172.805 ;
        RECT 72.965 172.135 73.135 172.635 ;
        RECT 70.965 171.225 71.180 171.735 ;
        RECT 71.410 171.405 71.690 171.735 ;
        RECT 71.870 171.225 72.110 171.735 ;
        RECT 72.480 171.395 73.095 171.965 ;
        RECT 73.385 171.905 73.650 172.465 ;
        RECT 73.820 171.735 73.990 172.635 ;
        RECT 74.750 172.625 75.010 173.775 ;
        RECT 75.185 172.700 75.440 173.605 ;
        RECT 75.610 173.015 75.940 173.775 ;
        RECT 76.155 172.845 76.325 173.605 ;
        RECT 74.160 171.905 74.515 172.465 ;
        RECT 73.265 171.225 73.480 171.735 ;
        RECT 73.710 171.405 73.990 171.735 ;
        RECT 74.170 171.225 74.410 171.735 ;
        RECT 74.750 171.225 75.010 172.065 ;
        RECT 75.185 171.970 75.355 172.700 ;
        RECT 75.610 172.675 76.325 172.845 ;
        RECT 75.610 172.465 75.780 172.675 ;
        RECT 76.585 172.610 76.875 173.775 ;
        RECT 77.230 172.805 77.620 172.980 ;
        RECT 78.105 172.975 78.435 173.775 ;
        RECT 78.605 172.985 79.140 173.605 ;
        RECT 77.230 172.635 78.655 172.805 ;
        RECT 75.525 172.135 75.780 172.465 ;
        RECT 75.185 171.395 75.440 171.970 ;
        RECT 75.610 171.945 75.780 172.135 ;
        RECT 76.060 172.125 76.415 172.495 ;
        RECT 75.610 171.775 76.325 171.945 ;
        RECT 75.610 171.225 75.940 171.605 ;
        RECT 76.155 171.395 76.325 171.775 ;
        RECT 76.585 171.225 76.875 171.950 ;
        RECT 77.105 171.905 77.460 172.465 ;
        RECT 77.630 171.735 77.800 172.635 ;
        RECT 77.970 171.905 78.235 172.465 ;
        RECT 78.485 172.135 78.655 172.635 ;
        RECT 78.825 171.965 79.140 172.985 ;
        RECT 79.530 172.805 79.920 172.980 ;
        RECT 80.405 172.975 80.735 173.775 ;
        RECT 80.905 172.985 81.440 173.605 ;
        RECT 79.530 172.635 80.955 172.805 ;
        RECT 77.210 171.225 77.450 171.735 ;
        RECT 77.630 171.405 77.910 171.735 ;
        RECT 78.140 171.225 78.355 171.735 ;
        RECT 78.525 171.395 79.140 171.965 ;
        RECT 79.405 171.905 79.760 172.465 ;
        RECT 79.930 171.735 80.100 172.635 ;
        RECT 80.270 171.905 80.535 172.465 ;
        RECT 80.785 172.135 80.955 172.635 ;
        RECT 81.125 171.965 81.440 172.985 ;
        RECT 81.830 172.805 82.220 172.980 ;
        RECT 82.705 172.975 83.035 173.775 ;
        RECT 83.205 172.985 83.740 173.605 ;
        RECT 81.830 172.635 83.255 172.805 ;
        RECT 79.510 171.225 79.750 171.735 ;
        RECT 79.930 171.405 80.210 171.735 ;
        RECT 80.440 171.225 80.655 171.735 ;
        RECT 80.825 171.395 81.440 171.965 ;
        RECT 81.705 171.905 82.060 172.465 ;
        RECT 82.230 171.735 82.400 172.635 ;
        RECT 82.570 171.905 82.835 172.465 ;
        RECT 83.085 172.135 83.255 172.635 ;
        RECT 83.425 171.965 83.740 172.985 ;
        RECT 84.410 173.385 84.745 173.605 ;
        RECT 85.750 173.395 86.105 173.775 ;
        RECT 84.410 172.765 84.665 173.385 ;
        RECT 84.915 173.225 85.145 173.265 ;
        RECT 86.275 173.225 86.525 173.605 ;
        RECT 84.915 173.025 86.525 173.225 ;
        RECT 84.915 172.935 85.100 173.025 ;
        RECT 85.690 173.015 86.525 173.025 ;
        RECT 86.775 172.995 87.025 173.775 ;
        RECT 87.195 172.925 87.455 173.605 ;
        RECT 85.255 172.825 85.585 172.855 ;
        RECT 85.255 172.765 87.055 172.825 ;
        RECT 84.410 172.655 87.115 172.765 ;
        RECT 84.410 172.595 85.585 172.655 ;
        RECT 86.915 172.620 87.115 172.655 ;
        RECT 84.405 172.215 84.895 172.415 ;
        RECT 85.085 172.215 85.560 172.425 ;
        RECT 81.810 171.225 82.050 171.735 ;
        RECT 82.230 171.405 82.510 171.735 ;
        RECT 82.740 171.225 82.955 171.735 ;
        RECT 83.125 171.395 83.740 171.965 ;
        RECT 84.410 171.225 84.865 171.990 ;
        RECT 85.340 171.815 85.560 172.215 ;
        RECT 85.805 172.215 86.135 172.425 ;
        RECT 85.805 171.815 86.015 172.215 ;
        RECT 86.305 172.180 86.715 172.485 ;
        RECT 86.945 172.045 87.115 172.620 ;
        RECT 86.845 171.925 87.115 172.045 ;
        RECT 86.270 171.880 87.115 171.925 ;
        RECT 86.270 171.755 87.025 171.880 ;
        RECT 86.270 171.605 86.440 171.755 ;
        RECT 87.285 171.735 87.455 172.925 ;
        RECT 88.545 172.685 89.755 173.775 ;
        RECT 88.545 172.145 89.065 172.685 ;
        RECT 89.235 171.975 89.755 172.515 ;
        RECT 87.225 171.725 87.455 171.735 ;
        RECT 85.140 171.395 86.440 171.605 ;
        RECT 86.695 171.225 87.025 171.585 ;
        RECT 87.195 171.395 87.455 171.725 ;
        RECT 88.545 171.225 89.755 171.975 ;
        RECT 12.100 171.055 89.840 171.225 ;
        RECT 12.185 170.305 13.395 171.055 ;
        RECT 13.565 170.510 18.910 171.055 ;
        RECT 19.085 170.510 24.430 171.055 ;
        RECT 24.605 170.510 29.950 171.055 ;
        RECT 30.125 170.510 35.470 171.055 ;
        RECT 12.185 169.765 12.705 170.305 ;
        RECT 12.875 169.595 13.395 170.135 ;
        RECT 15.150 169.680 15.490 170.510 ;
        RECT 12.185 168.505 13.395 169.595 ;
        RECT 16.970 168.940 17.320 170.190 ;
        RECT 20.670 169.680 21.010 170.510 ;
        RECT 22.490 168.940 22.840 170.190 ;
        RECT 26.190 169.680 26.530 170.510 ;
        RECT 28.010 168.940 28.360 170.190 ;
        RECT 31.710 169.680 32.050 170.510 ;
        RECT 35.645 170.285 37.315 171.055 ;
        RECT 37.945 170.330 38.235 171.055 ;
        RECT 38.405 170.285 40.075 171.055 ;
        RECT 33.530 168.940 33.880 170.190 ;
        RECT 35.645 169.765 36.395 170.285 ;
        RECT 36.565 169.595 37.315 170.115 ;
        RECT 38.405 169.765 39.155 170.285 ;
        RECT 13.565 168.505 18.910 168.940 ;
        RECT 19.085 168.505 24.430 168.940 ;
        RECT 24.605 168.505 29.950 168.940 ;
        RECT 30.125 168.505 35.470 168.940 ;
        RECT 35.645 168.505 37.315 169.595 ;
        RECT 37.945 168.505 38.235 169.670 ;
        RECT 39.325 169.595 40.075 170.115 ;
        RECT 38.405 168.505 40.075 169.595 ;
        RECT 40.245 170.070 40.515 170.885 ;
        RECT 40.685 170.315 41.355 171.055 ;
        RECT 41.525 170.485 41.820 170.830 ;
        RECT 42.000 170.655 42.375 171.055 ;
        RECT 42.590 170.485 42.920 170.830 ;
        RECT 41.525 170.315 42.920 170.485 ;
        RECT 43.170 170.315 43.755 170.885 ;
        RECT 43.925 170.510 49.270 171.055 ;
        RECT 40.245 168.675 40.595 170.070 ;
        RECT 40.765 169.645 40.935 170.145 ;
        RECT 41.105 169.815 41.440 170.145 ;
        RECT 41.610 169.815 41.950 170.145 ;
        RECT 40.765 169.475 41.510 169.645 ;
        RECT 40.765 168.505 41.170 169.305 ;
        RECT 41.340 168.845 41.510 169.475 ;
        RECT 41.680 169.070 41.950 169.815 ;
        RECT 42.140 169.815 42.430 170.145 ;
        RECT 42.600 169.815 43.000 170.145 ;
        RECT 42.140 169.070 42.375 169.815 ;
        RECT 43.170 169.645 43.340 170.315 ;
        RECT 43.510 169.815 43.755 170.145 ;
        RECT 45.510 169.680 45.850 170.510 ;
        RECT 49.445 170.285 51.115 171.055 ;
        RECT 42.545 169.475 43.755 169.645 ;
        RECT 42.545 168.845 42.875 169.475 ;
        RECT 41.340 168.675 42.875 168.845 ;
        RECT 43.060 168.505 43.295 169.305 ;
        RECT 43.465 168.675 43.755 169.475 ;
        RECT 47.330 168.940 47.680 170.190 ;
        RECT 49.445 169.765 50.195 170.285 ;
        RECT 51.285 170.255 51.595 171.055 ;
        RECT 51.800 170.255 52.495 170.885 ;
        RECT 52.665 170.510 58.010 171.055 ;
        RECT 50.365 169.595 51.115 170.115 ;
        RECT 51.295 169.815 51.630 170.085 ;
        RECT 51.800 169.655 51.970 170.255 ;
        RECT 52.140 169.815 52.475 170.065 ;
        RECT 54.250 169.680 54.590 170.510 ;
        RECT 58.190 170.215 58.450 171.055 ;
        RECT 58.625 170.310 58.880 170.885 ;
        RECT 59.050 170.675 59.380 171.055 ;
        RECT 59.595 170.505 59.765 170.885 ;
        RECT 59.050 170.335 59.765 170.505 ;
        RECT 60.140 170.425 60.425 170.885 ;
        RECT 60.595 170.595 60.865 171.055 ;
        RECT 43.925 168.505 49.270 168.940 ;
        RECT 49.445 168.505 51.115 169.595 ;
        RECT 51.285 168.505 51.565 169.645 ;
        RECT 51.735 168.675 52.065 169.655 ;
        RECT 52.235 168.505 52.495 169.645 ;
        RECT 56.070 168.940 56.420 170.190 ;
        RECT 52.665 168.505 58.010 168.940 ;
        RECT 58.190 168.505 58.450 169.655 ;
        RECT 58.625 169.580 58.795 170.310 ;
        RECT 59.050 170.145 59.220 170.335 ;
        RECT 60.140 170.255 61.095 170.425 ;
        RECT 58.965 169.815 59.220 170.145 ;
        RECT 59.050 169.605 59.220 169.815 ;
        RECT 59.500 169.785 59.855 170.155 ;
        RECT 58.625 168.675 58.880 169.580 ;
        RECT 59.050 169.435 59.765 169.605 ;
        RECT 60.025 169.525 60.715 170.085 ;
        RECT 59.050 168.505 59.380 169.265 ;
        RECT 59.595 168.675 59.765 169.435 ;
        RECT 60.885 169.355 61.095 170.255 ;
        RECT 60.140 169.135 61.095 169.355 ;
        RECT 61.265 170.085 61.665 170.885 ;
        RECT 61.855 170.425 62.135 170.885 ;
        RECT 62.655 170.595 62.980 171.055 ;
        RECT 61.855 170.255 62.980 170.425 ;
        RECT 63.150 170.315 63.535 170.885 ;
        RECT 63.705 170.330 63.995 171.055 ;
        RECT 62.530 170.145 62.980 170.255 ;
        RECT 61.265 169.525 62.360 170.085 ;
        RECT 62.530 169.815 63.085 170.145 ;
        RECT 60.140 168.675 60.425 169.135 ;
        RECT 60.595 168.505 60.865 168.965 ;
        RECT 61.265 168.675 61.665 169.525 ;
        RECT 62.530 169.355 62.980 169.815 ;
        RECT 63.255 169.645 63.535 170.315 ;
        RECT 64.165 170.315 64.550 170.885 ;
        RECT 64.720 170.595 65.045 171.055 ;
        RECT 65.565 170.425 65.845 170.885 ;
        RECT 61.855 169.135 62.980 169.355 ;
        RECT 61.855 168.675 62.135 169.135 ;
        RECT 62.655 168.505 62.980 168.965 ;
        RECT 63.150 168.675 63.535 169.645 ;
        RECT 63.705 168.505 63.995 169.670 ;
        RECT 64.165 169.645 64.445 170.315 ;
        RECT 64.720 170.255 65.845 170.425 ;
        RECT 64.720 170.145 65.170 170.255 ;
        RECT 64.615 169.815 65.170 170.145 ;
        RECT 66.035 170.085 66.435 170.885 ;
        RECT 66.835 170.595 67.105 171.055 ;
        RECT 67.275 170.425 67.560 170.885 ;
        RECT 64.165 168.675 64.550 169.645 ;
        RECT 64.720 169.355 65.170 169.815 ;
        RECT 65.340 169.525 66.435 170.085 ;
        RECT 64.720 169.135 65.845 169.355 ;
        RECT 64.720 168.505 65.045 168.965 ;
        RECT 65.565 168.675 65.845 169.135 ;
        RECT 66.035 168.675 66.435 169.525 ;
        RECT 66.605 170.255 67.560 170.425 ;
        RECT 68.815 170.400 69.145 170.835 ;
        RECT 69.315 170.445 69.485 171.055 ;
        RECT 68.765 170.315 69.145 170.400 ;
        RECT 69.655 170.315 69.985 170.840 ;
        RECT 70.245 170.525 70.455 171.055 ;
        RECT 70.730 170.605 71.515 170.775 ;
        RECT 71.685 170.605 72.090 170.775 ;
        RECT 68.765 170.275 68.990 170.315 ;
        RECT 66.605 169.355 66.815 170.255 ;
        RECT 66.985 169.525 67.675 170.085 ;
        RECT 68.765 169.695 68.935 170.275 ;
        RECT 69.655 170.145 69.855 170.315 ;
        RECT 70.730 170.145 70.900 170.605 ;
        RECT 69.105 169.815 69.855 170.145 ;
        RECT 70.025 169.815 70.900 170.145 ;
        RECT 68.765 169.645 68.980 169.695 ;
        RECT 68.765 169.565 69.155 169.645 ;
        RECT 66.605 169.135 67.560 169.355 ;
        RECT 66.835 168.505 67.105 168.965 ;
        RECT 67.275 168.675 67.560 169.135 ;
        RECT 68.825 168.720 69.155 169.565 ;
        RECT 69.665 169.610 69.855 169.815 ;
        RECT 69.325 168.505 69.495 169.515 ;
        RECT 69.665 169.235 70.560 169.610 ;
        RECT 69.665 168.675 70.005 169.235 ;
        RECT 70.235 168.505 70.550 169.005 ;
        RECT 70.730 168.975 70.900 169.815 ;
        RECT 71.070 170.105 71.535 170.435 ;
        RECT 71.920 170.375 72.090 170.605 ;
        RECT 72.270 170.555 72.640 171.055 ;
        RECT 72.960 170.605 73.635 170.775 ;
        RECT 73.830 170.605 74.165 170.775 ;
        RECT 71.070 169.145 71.390 170.105 ;
        RECT 71.920 170.075 72.750 170.375 ;
        RECT 71.560 169.175 71.750 169.895 ;
        RECT 71.920 169.005 72.090 170.075 ;
        RECT 72.550 170.045 72.750 170.075 ;
        RECT 72.260 169.825 72.430 169.895 ;
        RECT 72.960 169.825 73.130 170.605 ;
        RECT 73.995 170.465 74.165 170.605 ;
        RECT 74.335 170.595 74.585 171.055 ;
        RECT 72.260 169.655 73.130 169.825 ;
        RECT 73.300 170.185 73.825 170.405 ;
        RECT 73.995 170.335 74.220 170.465 ;
        RECT 72.260 169.565 72.770 169.655 ;
        RECT 70.730 168.805 71.615 168.975 ;
        RECT 71.840 168.675 72.090 169.005 ;
        RECT 72.260 168.505 72.430 169.305 ;
        RECT 72.600 168.950 72.770 169.565 ;
        RECT 73.300 169.485 73.470 170.185 ;
        RECT 72.940 169.120 73.470 169.485 ;
        RECT 73.640 169.420 73.880 170.015 ;
        RECT 74.050 169.230 74.220 170.335 ;
        RECT 74.390 169.475 74.670 170.425 ;
        RECT 73.915 169.100 74.220 169.230 ;
        RECT 72.600 168.780 73.705 168.950 ;
        RECT 73.915 168.675 74.165 169.100 ;
        RECT 74.335 168.505 74.600 168.965 ;
        RECT 74.840 168.675 75.025 170.795 ;
        RECT 75.195 170.675 75.525 171.055 ;
        RECT 75.695 170.505 75.865 170.795 ;
        RECT 75.200 170.335 75.865 170.505 ;
        RECT 75.200 169.345 75.430 170.335 ;
        RECT 77.045 170.255 77.385 170.885 ;
        RECT 77.555 170.255 77.805 171.055 ;
        RECT 77.995 170.405 78.325 170.885 ;
        RECT 78.495 170.595 78.720 171.055 ;
        RECT 78.890 170.405 79.220 170.885 ;
        RECT 75.600 169.515 75.950 170.165 ;
        RECT 77.045 169.645 77.220 170.255 ;
        RECT 77.995 170.235 79.220 170.405 ;
        RECT 79.850 170.275 80.350 170.885 ;
        RECT 77.390 169.895 78.085 170.065 ;
        RECT 77.915 169.645 78.085 169.895 ;
        RECT 78.260 169.865 78.680 170.065 ;
        RECT 78.850 169.865 79.180 170.065 ;
        RECT 79.350 169.865 79.680 170.065 ;
        RECT 79.850 169.645 80.020 170.275 ;
        RECT 80.725 170.255 81.065 170.885 ;
        RECT 81.235 170.255 81.485 171.055 ;
        RECT 81.675 170.405 82.005 170.885 ;
        RECT 82.175 170.595 82.400 171.055 ;
        RECT 82.570 170.405 82.900 170.885 ;
        RECT 80.205 169.815 80.555 170.065 ;
        RECT 80.725 169.645 80.900 170.255 ;
        RECT 81.675 170.235 82.900 170.405 ;
        RECT 83.530 170.275 84.030 170.885 ;
        RECT 84.405 170.555 84.665 170.885 ;
        RECT 84.835 170.695 85.165 171.055 ;
        RECT 85.420 170.675 86.720 170.885 ;
        RECT 81.070 169.895 81.765 170.065 ;
        RECT 81.595 169.645 81.765 169.895 ;
        RECT 81.940 169.865 82.360 170.065 ;
        RECT 82.530 169.865 82.860 170.065 ;
        RECT 83.030 169.865 83.360 170.065 ;
        RECT 83.530 169.645 83.700 170.275 ;
        RECT 83.885 169.815 84.235 170.065 ;
        RECT 75.200 169.175 75.865 169.345 ;
        RECT 75.195 168.505 75.525 169.005 ;
        RECT 75.695 168.675 75.865 169.175 ;
        RECT 77.045 168.675 77.385 169.645 ;
        RECT 77.555 168.505 77.725 169.645 ;
        RECT 77.915 169.475 80.350 169.645 ;
        RECT 77.995 168.505 78.245 169.305 ;
        RECT 78.890 168.675 79.220 169.475 ;
        RECT 79.520 168.505 79.850 169.305 ;
        RECT 80.020 168.675 80.350 169.475 ;
        RECT 80.725 168.675 81.065 169.645 ;
        RECT 81.235 168.505 81.405 169.645 ;
        RECT 81.595 169.475 84.030 169.645 ;
        RECT 81.675 168.505 81.925 169.305 ;
        RECT 82.570 168.675 82.900 169.475 ;
        RECT 83.200 168.505 83.530 169.305 ;
        RECT 83.700 168.675 84.030 169.475 ;
        RECT 84.405 169.355 84.575 170.555 ;
        RECT 85.420 170.525 85.590 170.675 ;
        RECT 84.835 170.400 85.590 170.525 ;
        RECT 84.745 170.355 85.590 170.400 ;
        RECT 84.745 170.235 85.015 170.355 ;
        RECT 84.745 169.660 84.915 170.235 ;
        RECT 85.145 169.795 85.555 170.100 ;
        RECT 85.845 170.065 86.055 170.465 ;
        RECT 85.725 169.855 86.055 170.065 ;
        RECT 86.300 170.065 86.520 170.465 ;
        RECT 86.995 170.290 87.450 171.055 ;
        RECT 88.545 170.305 89.755 171.055 ;
        RECT 86.300 169.855 86.775 170.065 ;
        RECT 86.965 169.865 87.455 170.065 ;
        RECT 84.745 169.625 84.945 169.660 ;
        RECT 86.275 169.625 87.450 169.685 ;
        RECT 84.745 169.515 87.450 169.625 ;
        RECT 84.805 169.455 86.605 169.515 ;
        RECT 86.275 169.425 86.605 169.455 ;
        RECT 84.405 168.675 84.665 169.355 ;
        RECT 84.835 168.505 85.085 169.285 ;
        RECT 85.335 169.255 86.170 169.265 ;
        RECT 86.760 169.255 86.945 169.345 ;
        RECT 85.335 169.055 86.945 169.255 ;
        RECT 85.335 168.675 85.585 169.055 ;
        RECT 86.715 169.015 86.945 169.055 ;
        RECT 87.195 168.895 87.450 169.515 ;
        RECT 85.755 168.505 86.110 168.885 ;
        RECT 87.115 168.675 87.450 168.895 ;
        RECT 88.545 169.595 89.065 170.135 ;
        RECT 89.235 169.765 89.755 170.305 ;
        RECT 100.140 170.940 100.810 174.200 ;
        RECT 101.480 173.630 105.520 173.800 ;
        RECT 101.140 171.570 101.310 173.570 ;
        RECT 105.690 171.570 105.860 173.570 ;
        RECT 101.480 171.340 105.520 171.510 ;
        RECT 106.200 170.940 106.370 174.200 ;
        RECT 100.140 170.770 106.370 170.940 ;
        RECT 88.545 168.505 89.755 169.595 ;
        RECT 12.100 168.335 89.840 168.505 ;
        RECT 12.185 167.245 13.395 168.335 ;
        RECT 13.565 167.900 18.910 168.335 ;
        RECT 19.085 167.900 24.430 168.335 ;
        RECT 12.185 166.535 12.705 167.075 ;
        RECT 12.875 166.705 13.395 167.245 ;
        RECT 12.185 165.785 13.395 166.535 ;
        RECT 15.150 166.330 15.490 167.160 ;
        RECT 16.970 166.650 17.320 167.900 ;
        RECT 20.670 166.330 21.010 167.160 ;
        RECT 22.490 166.650 22.840 167.900 ;
        RECT 25.065 167.170 25.355 168.335 ;
        RECT 25.525 167.900 30.870 168.335 ;
        RECT 31.045 167.900 36.390 168.335 ;
        RECT 13.565 165.785 18.910 166.330 ;
        RECT 19.085 165.785 24.430 166.330 ;
        RECT 25.065 165.785 25.355 166.510 ;
        RECT 27.110 166.330 27.450 167.160 ;
        RECT 28.930 166.650 29.280 167.900 ;
        RECT 32.630 166.330 32.970 167.160 ;
        RECT 34.450 166.650 34.800 167.900 ;
        RECT 36.565 167.245 38.235 168.335 ;
        RECT 38.955 167.665 39.125 168.165 ;
        RECT 39.295 167.835 39.625 168.335 ;
        RECT 38.955 167.495 39.620 167.665 ;
        RECT 36.565 166.555 37.315 167.075 ;
        RECT 37.485 166.725 38.235 167.245 ;
        RECT 38.870 166.675 39.220 167.325 ;
        RECT 25.525 165.785 30.870 166.330 ;
        RECT 31.045 165.785 36.390 166.330 ;
        RECT 36.565 165.785 38.235 166.555 ;
        RECT 39.390 166.505 39.620 167.495 ;
        RECT 38.955 166.335 39.620 166.505 ;
        RECT 38.955 166.045 39.125 166.335 ;
        RECT 39.295 165.785 39.625 166.165 ;
        RECT 39.795 166.045 39.980 168.165 ;
        RECT 40.220 167.875 40.485 168.335 ;
        RECT 40.655 167.740 40.905 168.165 ;
        RECT 41.115 167.890 42.220 168.060 ;
        RECT 40.600 167.610 40.905 167.740 ;
        RECT 40.150 166.415 40.430 167.365 ;
        RECT 40.600 166.505 40.770 167.610 ;
        RECT 40.940 166.825 41.180 167.420 ;
        RECT 41.350 167.355 41.880 167.720 ;
        RECT 41.350 166.655 41.520 167.355 ;
        RECT 42.050 167.275 42.220 167.890 ;
        RECT 42.390 167.535 42.560 168.335 ;
        RECT 42.730 167.835 42.980 168.165 ;
        RECT 43.205 167.865 44.090 168.035 ;
        RECT 42.050 167.185 42.560 167.275 ;
        RECT 40.600 166.375 40.825 166.505 ;
        RECT 40.995 166.435 41.520 166.655 ;
        RECT 41.690 167.015 42.560 167.185 ;
        RECT 40.235 165.785 40.485 166.245 ;
        RECT 40.655 166.235 40.825 166.375 ;
        RECT 41.690 166.235 41.860 167.015 ;
        RECT 42.390 166.945 42.560 167.015 ;
        RECT 42.070 166.765 42.270 166.795 ;
        RECT 42.730 166.765 42.900 167.835 ;
        RECT 43.070 166.945 43.260 167.665 ;
        RECT 42.070 166.465 42.900 166.765 ;
        RECT 43.430 166.735 43.750 167.695 ;
        RECT 40.655 166.065 40.990 166.235 ;
        RECT 41.185 166.065 41.860 166.235 ;
        RECT 42.180 165.785 42.550 166.285 ;
        RECT 42.730 166.235 42.900 166.465 ;
        RECT 43.285 166.405 43.750 166.735 ;
        RECT 43.920 167.025 44.090 167.865 ;
        RECT 44.270 167.835 44.585 168.335 ;
        RECT 44.815 167.605 45.155 168.165 ;
        RECT 44.260 167.230 45.155 167.605 ;
        RECT 45.325 167.325 45.495 168.335 ;
        RECT 44.965 167.025 45.155 167.230 ;
        RECT 45.665 167.275 45.995 168.120 ;
        RECT 46.260 167.545 46.795 168.165 ;
        RECT 45.665 167.195 46.055 167.275 ;
        RECT 45.840 167.145 46.055 167.195 ;
        RECT 43.920 166.695 44.795 167.025 ;
        RECT 44.965 166.695 45.715 167.025 ;
        RECT 43.920 166.235 44.090 166.695 ;
        RECT 44.965 166.525 45.165 166.695 ;
        RECT 45.885 166.565 46.055 167.145 ;
        RECT 45.830 166.525 46.055 166.565 ;
        RECT 42.730 166.065 43.135 166.235 ;
        RECT 43.305 166.065 44.090 166.235 ;
        RECT 44.365 165.785 44.575 166.315 ;
        RECT 44.835 166.000 45.165 166.525 ;
        RECT 45.675 166.440 46.055 166.525 ;
        RECT 46.260 166.525 46.575 167.545 ;
        RECT 46.965 167.535 47.295 168.335 ;
        RECT 47.780 167.365 48.170 167.540 ;
        RECT 48.530 167.535 48.785 168.335 ;
        RECT 48.985 167.485 49.315 168.165 ;
        RECT 46.745 167.195 48.170 167.365 ;
        RECT 46.745 166.695 46.915 167.195 ;
        RECT 45.335 165.785 45.505 166.395 ;
        RECT 45.675 166.005 46.005 166.440 ;
        RECT 46.260 165.955 46.875 166.525 ;
        RECT 47.165 166.465 47.430 167.025 ;
        RECT 47.600 166.295 47.770 167.195 ;
        RECT 47.940 166.465 48.295 167.025 ;
        RECT 48.530 166.995 48.775 167.355 ;
        RECT 48.965 167.205 49.315 167.485 ;
        RECT 48.965 166.825 49.135 167.205 ;
        RECT 49.495 167.025 49.690 168.075 ;
        RECT 49.870 167.195 50.190 168.335 ;
        RECT 50.825 167.170 51.115 168.335 ;
        RECT 51.285 167.195 51.670 168.165 ;
        RECT 51.840 167.875 52.165 168.335 ;
        RECT 52.685 167.705 52.965 168.165 ;
        RECT 51.840 167.485 52.965 167.705 ;
        RECT 48.615 166.655 49.135 166.825 ;
        RECT 49.305 166.695 49.690 167.025 ;
        RECT 49.870 166.975 50.130 167.025 ;
        RECT 49.870 166.805 50.135 166.975 ;
        RECT 49.870 166.695 50.130 166.805 ;
        RECT 48.615 166.295 48.785 166.655 ;
        RECT 51.285 166.525 51.565 167.195 ;
        RECT 51.840 167.025 52.290 167.485 ;
        RECT 53.155 167.315 53.555 168.165 ;
        RECT 53.955 167.875 54.225 168.335 ;
        RECT 54.395 167.705 54.680 168.165 ;
        RECT 51.735 166.695 52.290 167.025 ;
        RECT 52.460 166.755 53.555 167.315 ;
        RECT 51.840 166.585 52.290 166.695 ;
        RECT 47.045 165.785 47.260 166.295 ;
        RECT 47.490 165.965 47.770 166.295 ;
        RECT 47.950 165.785 48.190 166.295 ;
        RECT 48.585 166.125 48.785 166.295 ;
        RECT 48.615 166.090 48.785 166.125 ;
        RECT 48.975 166.315 50.190 166.485 ;
        RECT 48.975 166.010 49.205 166.315 ;
        RECT 49.375 165.785 49.705 166.145 ;
        RECT 49.900 165.965 50.190 166.315 ;
        RECT 50.825 165.785 51.115 166.510 ;
        RECT 51.285 165.955 51.670 166.525 ;
        RECT 51.840 166.415 52.965 166.585 ;
        RECT 51.840 165.785 52.165 166.245 ;
        RECT 52.685 165.955 52.965 166.415 ;
        RECT 53.155 165.955 53.555 166.755 ;
        RECT 53.725 167.485 54.680 167.705 ;
        RECT 55.055 167.665 55.225 168.165 ;
        RECT 55.395 167.835 55.725 168.335 ;
        RECT 55.055 167.495 55.720 167.665 ;
        RECT 53.725 166.585 53.935 167.485 ;
        RECT 54.105 166.755 54.795 167.315 ;
        RECT 54.970 166.675 55.320 167.325 ;
        RECT 53.725 166.415 54.680 166.585 ;
        RECT 55.490 166.505 55.720 167.495 ;
        RECT 53.955 165.785 54.225 166.245 ;
        RECT 54.395 165.955 54.680 166.415 ;
        RECT 55.055 166.335 55.720 166.505 ;
        RECT 55.055 166.045 55.225 166.335 ;
        RECT 55.395 165.785 55.725 166.165 ;
        RECT 55.895 166.045 56.080 168.165 ;
        RECT 56.320 167.875 56.585 168.335 ;
        RECT 56.755 167.740 57.005 168.165 ;
        RECT 57.215 167.890 58.320 168.060 ;
        RECT 56.700 167.610 57.005 167.740 ;
        RECT 56.250 166.415 56.530 167.365 ;
        RECT 56.700 166.505 56.870 167.610 ;
        RECT 57.040 166.825 57.280 167.420 ;
        RECT 57.450 167.355 57.980 167.720 ;
        RECT 57.450 166.655 57.620 167.355 ;
        RECT 58.150 167.275 58.320 167.890 ;
        RECT 58.490 167.535 58.660 168.335 ;
        RECT 58.830 167.835 59.080 168.165 ;
        RECT 59.305 167.865 60.190 168.035 ;
        RECT 58.150 167.185 58.660 167.275 ;
        RECT 56.700 166.375 56.925 166.505 ;
        RECT 57.095 166.435 57.620 166.655 ;
        RECT 57.790 167.015 58.660 167.185 ;
        RECT 56.335 165.785 56.585 166.245 ;
        RECT 56.755 166.235 56.925 166.375 ;
        RECT 57.790 166.235 57.960 167.015 ;
        RECT 58.490 166.945 58.660 167.015 ;
        RECT 58.170 166.765 58.370 166.795 ;
        RECT 58.830 166.765 59.000 167.835 ;
        RECT 59.170 166.945 59.360 167.665 ;
        RECT 58.170 166.465 59.000 166.765 ;
        RECT 59.530 166.735 59.850 167.695 ;
        RECT 56.755 166.065 57.090 166.235 ;
        RECT 57.285 166.065 57.960 166.235 ;
        RECT 58.280 165.785 58.650 166.285 ;
        RECT 58.830 166.235 59.000 166.465 ;
        RECT 59.385 166.405 59.850 166.735 ;
        RECT 60.020 167.025 60.190 167.865 ;
        RECT 60.370 167.835 60.685 168.335 ;
        RECT 60.915 167.605 61.255 168.165 ;
        RECT 60.360 167.230 61.255 167.605 ;
        RECT 61.425 167.325 61.595 168.335 ;
        RECT 61.065 167.025 61.255 167.230 ;
        RECT 61.765 167.275 62.095 168.120 ;
        RECT 61.765 167.195 62.155 167.275 ;
        RECT 61.940 167.145 62.155 167.195 ;
        RECT 60.020 166.695 60.895 167.025 ;
        RECT 61.065 166.695 61.815 167.025 ;
        RECT 60.020 166.235 60.190 166.695 ;
        RECT 61.065 166.525 61.265 166.695 ;
        RECT 61.985 166.565 62.155 167.145 ;
        RECT 61.930 166.525 62.155 166.565 ;
        RECT 58.830 166.065 59.235 166.235 ;
        RECT 59.405 166.065 60.190 166.235 ;
        RECT 60.465 165.785 60.675 166.315 ;
        RECT 60.935 166.000 61.265 166.525 ;
        RECT 61.775 166.440 62.155 166.525 ;
        RECT 62.330 167.195 62.665 168.165 ;
        RECT 62.835 167.195 63.005 168.335 ;
        RECT 63.175 167.995 65.205 168.165 ;
        RECT 62.330 166.525 62.500 167.195 ;
        RECT 63.175 167.025 63.345 167.995 ;
        RECT 62.670 166.695 62.925 167.025 ;
        RECT 63.150 166.695 63.345 167.025 ;
        RECT 63.515 167.655 64.640 167.825 ;
        RECT 62.755 166.525 62.925 166.695 ;
        RECT 63.515 166.525 63.685 167.655 ;
        RECT 61.435 165.785 61.605 166.395 ;
        RECT 61.775 166.005 62.105 166.440 ;
        RECT 62.330 165.955 62.585 166.525 ;
        RECT 62.755 166.355 63.685 166.525 ;
        RECT 63.855 167.315 64.865 167.485 ;
        RECT 63.855 166.515 64.025 167.315 ;
        RECT 63.510 166.320 63.685 166.355 ;
        RECT 62.755 165.785 63.085 166.185 ;
        RECT 63.510 165.955 64.040 166.320 ;
        RECT 64.230 166.295 64.505 167.115 ;
        RECT 64.225 166.125 64.505 166.295 ;
        RECT 64.230 165.955 64.505 166.125 ;
        RECT 64.675 165.955 64.865 167.315 ;
        RECT 65.035 167.330 65.205 167.995 ;
        RECT 65.375 167.575 65.545 168.335 ;
        RECT 65.780 167.575 66.295 167.985 ;
        RECT 65.035 167.140 65.785 167.330 ;
        RECT 65.955 166.765 66.295 167.575 ;
        RECT 67.445 167.275 67.775 168.120 ;
        RECT 67.945 167.325 68.115 168.335 ;
        RECT 68.285 167.605 68.625 168.165 ;
        RECT 68.855 167.835 69.170 168.335 ;
        RECT 69.350 167.865 70.235 168.035 ;
        RECT 65.065 166.595 66.295 166.765 ;
        RECT 67.385 167.195 67.775 167.275 ;
        RECT 68.285 167.230 69.180 167.605 ;
        RECT 67.385 167.145 67.600 167.195 ;
        RECT 65.045 165.785 65.555 166.320 ;
        RECT 65.775 165.990 66.020 166.595 ;
        RECT 67.385 166.565 67.555 167.145 ;
        RECT 68.285 167.025 68.475 167.230 ;
        RECT 69.350 167.025 69.520 167.865 ;
        RECT 70.460 167.835 70.710 168.165 ;
        RECT 67.725 166.695 68.475 167.025 ;
        RECT 68.645 166.695 69.520 167.025 ;
        RECT 67.385 166.525 67.610 166.565 ;
        RECT 68.275 166.525 68.475 166.695 ;
        RECT 67.385 166.440 67.765 166.525 ;
        RECT 67.435 166.005 67.765 166.440 ;
        RECT 67.935 165.785 68.105 166.395 ;
        RECT 68.275 166.000 68.605 166.525 ;
        RECT 68.865 165.785 69.075 166.315 ;
        RECT 69.350 166.235 69.520 166.695 ;
        RECT 69.690 166.735 70.010 167.695 ;
        RECT 70.180 166.945 70.370 167.665 ;
        RECT 70.540 166.765 70.710 167.835 ;
        RECT 70.880 167.535 71.050 168.335 ;
        RECT 71.220 167.890 72.325 168.060 ;
        RECT 71.220 167.275 71.390 167.890 ;
        RECT 72.535 167.740 72.785 168.165 ;
        RECT 72.955 167.875 73.220 168.335 ;
        RECT 71.560 167.355 72.090 167.720 ;
        RECT 72.535 167.610 72.840 167.740 ;
        RECT 70.880 167.185 71.390 167.275 ;
        RECT 70.880 167.015 71.750 167.185 ;
        RECT 70.880 166.945 71.050 167.015 ;
        RECT 71.170 166.765 71.370 166.795 ;
        RECT 69.690 166.405 70.155 166.735 ;
        RECT 70.540 166.465 71.370 166.765 ;
        RECT 70.540 166.235 70.710 166.465 ;
        RECT 69.350 166.065 70.135 166.235 ;
        RECT 70.305 166.065 70.710 166.235 ;
        RECT 70.890 165.785 71.260 166.285 ;
        RECT 71.580 166.235 71.750 167.015 ;
        RECT 71.920 166.655 72.090 167.355 ;
        RECT 72.260 166.825 72.500 167.420 ;
        RECT 71.920 166.435 72.445 166.655 ;
        RECT 72.670 166.505 72.840 167.610 ;
        RECT 72.615 166.375 72.840 166.505 ;
        RECT 73.010 166.415 73.290 167.365 ;
        RECT 72.615 166.235 72.785 166.375 ;
        RECT 71.580 166.065 72.255 166.235 ;
        RECT 72.450 166.065 72.785 166.235 ;
        RECT 72.955 165.785 73.205 166.245 ;
        RECT 73.460 166.045 73.645 168.165 ;
        RECT 73.815 167.835 74.145 168.335 ;
        RECT 74.315 167.665 74.485 168.165 ;
        RECT 73.820 167.495 74.485 167.665 ;
        RECT 73.820 166.505 74.050 167.495 ;
        RECT 74.835 167.405 75.005 168.165 ;
        RECT 75.220 167.575 75.550 168.335 ;
        RECT 74.220 166.675 74.570 167.325 ;
        RECT 74.835 167.235 75.550 167.405 ;
        RECT 75.720 167.260 75.975 168.165 ;
        RECT 74.745 166.685 75.100 167.055 ;
        RECT 75.380 167.025 75.550 167.235 ;
        RECT 75.380 166.695 75.635 167.025 ;
        RECT 75.380 166.505 75.550 166.695 ;
        RECT 75.805 166.530 75.975 167.260 ;
        RECT 76.150 167.185 76.410 168.335 ;
        RECT 76.585 167.170 76.875 168.335 ;
        RECT 77.135 167.665 77.305 168.165 ;
        RECT 77.475 167.835 77.805 168.335 ;
        RECT 77.135 167.495 77.800 167.665 ;
        RECT 77.050 166.675 77.400 167.325 ;
        RECT 73.820 166.335 74.485 166.505 ;
        RECT 73.815 165.785 74.145 166.165 ;
        RECT 74.315 166.045 74.485 166.335 ;
        RECT 74.835 166.335 75.550 166.505 ;
        RECT 74.835 165.955 75.005 166.335 ;
        RECT 75.220 165.785 75.550 166.165 ;
        RECT 75.720 165.955 75.975 166.530 ;
        RECT 76.150 165.785 76.410 166.625 ;
        RECT 76.585 165.785 76.875 166.510 ;
        RECT 77.570 166.505 77.800 167.495 ;
        RECT 77.135 166.335 77.800 166.505 ;
        RECT 77.135 166.045 77.305 166.335 ;
        RECT 77.475 165.785 77.805 166.165 ;
        RECT 77.975 166.045 78.160 168.165 ;
        RECT 78.400 167.875 78.665 168.335 ;
        RECT 78.835 167.740 79.085 168.165 ;
        RECT 79.295 167.890 80.400 168.060 ;
        RECT 78.780 167.610 79.085 167.740 ;
        RECT 78.330 166.415 78.610 167.365 ;
        RECT 78.780 166.505 78.950 167.610 ;
        RECT 79.120 166.825 79.360 167.420 ;
        RECT 79.530 167.355 80.060 167.720 ;
        RECT 79.530 166.655 79.700 167.355 ;
        RECT 80.230 167.275 80.400 167.890 ;
        RECT 80.570 167.535 80.740 168.335 ;
        RECT 80.910 167.835 81.160 168.165 ;
        RECT 81.385 167.865 82.270 168.035 ;
        RECT 80.230 167.185 80.740 167.275 ;
        RECT 78.780 166.375 79.005 166.505 ;
        RECT 79.175 166.435 79.700 166.655 ;
        RECT 79.870 167.015 80.740 167.185 ;
        RECT 78.415 165.785 78.665 166.245 ;
        RECT 78.835 166.235 79.005 166.375 ;
        RECT 79.870 166.235 80.040 167.015 ;
        RECT 80.570 166.945 80.740 167.015 ;
        RECT 80.250 166.765 80.450 166.795 ;
        RECT 80.910 166.765 81.080 167.835 ;
        RECT 81.250 166.945 81.440 167.665 ;
        RECT 80.250 166.465 81.080 166.765 ;
        RECT 81.610 166.735 81.930 167.695 ;
        RECT 78.835 166.065 79.170 166.235 ;
        RECT 79.365 166.065 80.040 166.235 ;
        RECT 80.360 165.785 80.730 166.285 ;
        RECT 80.910 166.235 81.080 166.465 ;
        RECT 81.465 166.405 81.930 166.735 ;
        RECT 82.100 167.025 82.270 167.865 ;
        RECT 82.450 167.835 82.765 168.335 ;
        RECT 82.995 167.605 83.335 168.165 ;
        RECT 82.440 167.230 83.335 167.605 ;
        RECT 83.505 167.325 83.675 168.335 ;
        RECT 83.145 167.025 83.335 167.230 ;
        RECT 83.845 167.275 84.175 168.120 ;
        RECT 84.870 167.945 85.205 168.165 ;
        RECT 86.210 167.955 86.565 168.335 ;
        RECT 84.870 167.325 85.125 167.945 ;
        RECT 85.375 167.785 85.605 167.825 ;
        RECT 86.735 167.785 86.985 168.165 ;
        RECT 85.375 167.585 86.985 167.785 ;
        RECT 85.375 167.495 85.560 167.585 ;
        RECT 86.150 167.575 86.985 167.585 ;
        RECT 87.235 167.555 87.485 168.335 ;
        RECT 87.655 167.485 87.915 168.165 ;
        RECT 85.715 167.385 86.045 167.415 ;
        RECT 85.715 167.325 87.515 167.385 ;
        RECT 83.845 167.195 84.235 167.275 ;
        RECT 84.020 167.145 84.235 167.195 ;
        RECT 84.870 167.215 87.575 167.325 ;
        RECT 84.870 167.155 86.045 167.215 ;
        RECT 87.375 167.180 87.575 167.215 ;
        RECT 82.100 166.695 82.975 167.025 ;
        RECT 83.145 166.695 83.895 167.025 ;
        RECT 82.100 166.235 82.270 166.695 ;
        RECT 83.145 166.525 83.345 166.695 ;
        RECT 84.065 166.565 84.235 167.145 ;
        RECT 84.865 166.775 85.355 166.975 ;
        RECT 85.545 166.775 86.020 166.985 ;
        RECT 84.010 166.525 84.235 166.565 ;
        RECT 80.910 166.065 81.315 166.235 ;
        RECT 81.485 166.065 82.270 166.235 ;
        RECT 82.545 165.785 82.755 166.315 ;
        RECT 83.015 166.000 83.345 166.525 ;
        RECT 83.855 166.440 84.235 166.525 ;
        RECT 83.515 165.785 83.685 166.395 ;
        RECT 83.855 166.005 84.185 166.440 ;
        RECT 84.870 165.785 85.325 166.550 ;
        RECT 85.800 166.375 86.020 166.775 ;
        RECT 86.265 166.775 86.595 166.985 ;
        RECT 86.265 166.375 86.475 166.775 ;
        RECT 86.765 166.740 87.175 167.045 ;
        RECT 87.405 166.605 87.575 167.180 ;
        RECT 87.305 166.485 87.575 166.605 ;
        RECT 86.730 166.440 87.575 166.485 ;
        RECT 86.730 166.315 87.485 166.440 ;
        RECT 86.730 166.165 86.900 166.315 ;
        RECT 87.745 166.285 87.915 167.485 ;
        RECT 88.545 167.245 89.755 168.335 ;
        RECT 100.140 167.510 100.810 170.770 ;
        RECT 101.480 170.200 105.520 170.370 ;
        RECT 101.140 168.140 101.310 170.140 ;
        RECT 105.690 168.140 105.860 170.140 ;
        RECT 101.480 167.910 105.520 168.080 ;
        RECT 106.200 167.510 106.370 170.770 ;
        RECT 100.140 167.500 106.370 167.510 ;
        RECT 107.960 176.770 117.790 176.810 ;
        RECT 140.540 176.790 146.280 176.800 ;
        RECT 107.960 176.640 118.590 176.770 ;
        RECT 120.510 176.740 126.250 176.750 ;
        RECT 107.960 174.380 108.130 176.640 ;
        RECT 108.855 176.070 116.895 176.240 ;
        RECT 108.470 175.010 108.640 176.010 ;
        RECT 117.110 175.010 117.280 176.010 ;
        RECT 108.855 174.780 116.895 174.950 ;
        RECT 117.620 174.380 118.590 176.640 ;
        RECT 107.960 174.210 118.590 174.380 ;
        RECT 107.960 170.950 108.130 174.210 ;
        RECT 108.855 173.640 116.895 173.810 ;
        RECT 108.470 171.580 108.640 173.580 ;
        RECT 117.110 171.580 117.280 173.580 ;
        RECT 108.855 171.350 116.895 171.520 ;
        RECT 117.620 170.950 118.590 174.210 ;
        RECT 107.960 170.780 118.590 170.950 ;
        RECT 107.960 167.520 108.130 170.780 ;
        RECT 108.855 170.210 116.895 170.380 ;
        RECT 108.470 168.150 108.640 170.150 ;
        RECT 117.110 168.150 117.280 170.150 ;
        RECT 108.855 167.920 116.895 168.090 ;
        RECT 117.620 167.520 118.590 170.780 ;
        RECT 100.140 167.400 106.380 167.500 ;
        RECT 88.545 166.705 89.065 167.245 ;
        RECT 89.235 166.535 89.755 167.075 ;
        RECT 85.600 165.955 86.900 166.165 ;
        RECT 87.155 165.785 87.485 166.145 ;
        RECT 87.655 165.955 87.915 166.285 ;
        RECT 88.545 165.785 89.755 166.535 ;
        RECT 100.130 166.840 106.380 167.400 ;
        RECT 100.130 166.820 105.300 166.840 ;
        RECT 100.130 166.750 104.120 166.820 ;
        RECT 12.100 165.615 89.840 165.785 ;
        RECT 12.185 164.865 13.395 165.615 ;
        RECT 13.565 165.070 18.910 165.615 ;
        RECT 19.085 165.070 24.430 165.615 ;
        RECT 24.605 165.070 29.950 165.615 ;
        RECT 30.125 165.070 35.470 165.615 ;
        RECT 12.185 164.325 12.705 164.865 ;
        RECT 12.875 164.155 13.395 164.695 ;
        RECT 15.150 164.240 15.490 165.070 ;
        RECT 12.185 163.065 13.395 164.155 ;
        RECT 16.970 163.500 17.320 164.750 ;
        RECT 20.670 164.240 21.010 165.070 ;
        RECT 22.490 163.500 22.840 164.750 ;
        RECT 26.190 164.240 26.530 165.070 ;
        RECT 28.010 163.500 28.360 164.750 ;
        RECT 31.710 164.240 32.050 165.070 ;
        RECT 35.645 164.845 37.315 165.615 ;
        RECT 37.945 164.890 38.235 165.615 ;
        RECT 38.405 164.845 40.075 165.615 ;
        RECT 40.245 164.875 40.630 165.445 ;
        RECT 40.800 165.155 41.125 165.615 ;
        RECT 41.645 164.985 41.925 165.445 ;
        RECT 33.530 163.500 33.880 164.750 ;
        RECT 35.645 164.325 36.395 164.845 ;
        RECT 36.565 164.155 37.315 164.675 ;
        RECT 38.405 164.325 39.155 164.845 ;
        RECT 13.565 163.065 18.910 163.500 ;
        RECT 19.085 163.065 24.430 163.500 ;
        RECT 24.605 163.065 29.950 163.500 ;
        RECT 30.125 163.065 35.470 163.500 ;
        RECT 35.645 163.065 37.315 164.155 ;
        RECT 37.945 163.065 38.235 164.230 ;
        RECT 39.325 164.155 40.075 164.675 ;
        RECT 38.405 163.065 40.075 164.155 ;
        RECT 40.245 164.205 40.525 164.875 ;
        RECT 40.800 164.815 41.925 164.985 ;
        RECT 40.800 164.705 41.250 164.815 ;
        RECT 40.695 164.375 41.250 164.705 ;
        RECT 42.115 164.645 42.515 165.445 ;
        RECT 42.915 165.155 43.185 165.615 ;
        RECT 43.355 164.985 43.640 165.445 ;
        RECT 40.245 163.235 40.630 164.205 ;
        RECT 40.800 163.915 41.250 164.375 ;
        RECT 41.420 164.085 42.515 164.645 ;
        RECT 40.800 163.695 41.925 163.915 ;
        RECT 40.800 163.065 41.125 163.525 ;
        RECT 41.645 163.235 41.925 163.695 ;
        RECT 42.115 163.235 42.515 164.085 ;
        RECT 42.685 164.815 43.640 164.985 ;
        RECT 43.925 164.890 44.185 165.445 ;
        RECT 44.355 165.170 44.785 165.615 ;
        RECT 45.020 165.045 45.190 165.445 ;
        RECT 45.360 165.215 46.080 165.615 ;
        RECT 42.685 163.915 42.895 164.815 ;
        RECT 43.065 164.085 43.755 164.645 ;
        RECT 43.925 164.175 44.100 164.890 ;
        RECT 45.020 164.875 45.900 165.045 ;
        RECT 46.250 165.000 46.420 165.445 ;
        RECT 46.995 165.105 47.395 165.615 ;
        RECT 44.270 164.375 44.525 164.705 ;
        RECT 42.685 163.695 43.640 163.915 ;
        RECT 42.915 163.065 43.185 163.525 ;
        RECT 43.355 163.235 43.640 163.695 ;
        RECT 43.925 163.235 44.185 164.175 ;
        RECT 44.355 163.895 44.525 164.375 ;
        RECT 44.750 164.085 45.080 164.705 ;
        RECT 45.250 164.325 45.540 164.705 ;
        RECT 45.730 164.155 45.900 164.875 ;
        RECT 45.380 163.985 45.900 164.155 ;
        RECT 46.070 164.830 46.420 165.000 ;
        RECT 47.695 165.065 47.865 165.355 ;
        RECT 48.035 165.235 48.365 165.615 ;
        RECT 44.355 163.725 45.115 163.895 ;
        RECT 45.380 163.795 45.550 163.985 ;
        RECT 46.070 163.805 46.240 164.830 ;
        RECT 46.660 164.345 46.920 164.935 ;
        RECT 46.440 164.045 46.920 164.345 ;
        RECT 47.120 164.045 47.380 164.935 ;
        RECT 47.695 164.895 48.360 165.065 ;
        RECT 47.610 164.075 47.960 164.725 ;
        RECT 48.130 163.905 48.360 164.895 ;
        RECT 44.945 163.500 45.115 163.725 ;
        RECT 45.830 163.635 46.240 163.805 ;
        RECT 46.415 163.695 47.355 163.865 ;
        RECT 45.830 163.500 46.085 163.635 ;
        RECT 44.355 163.065 44.685 163.465 ;
        RECT 44.945 163.330 46.085 163.500 ;
        RECT 46.415 163.445 46.585 163.695 ;
        RECT 45.830 163.235 46.085 163.330 ;
        RECT 46.255 163.275 46.585 163.445 ;
        RECT 46.755 163.065 47.005 163.525 ;
        RECT 47.175 163.235 47.355 163.695 ;
        RECT 47.695 163.735 48.360 163.905 ;
        RECT 47.695 163.235 47.865 163.735 ;
        RECT 48.035 163.065 48.365 163.565 ;
        RECT 48.535 163.235 48.720 165.355 ;
        RECT 48.975 165.155 49.225 165.615 ;
        RECT 49.395 165.165 49.730 165.335 ;
        RECT 49.925 165.165 50.600 165.335 ;
        RECT 49.395 165.025 49.565 165.165 ;
        RECT 48.890 164.035 49.170 164.985 ;
        RECT 49.340 164.895 49.565 165.025 ;
        RECT 49.340 163.790 49.510 164.895 ;
        RECT 49.735 164.745 50.260 164.965 ;
        RECT 49.680 163.980 49.920 164.575 ;
        RECT 50.090 164.045 50.260 164.745 ;
        RECT 50.430 164.385 50.600 165.165 ;
        RECT 50.920 165.115 51.290 165.615 ;
        RECT 51.470 165.165 51.875 165.335 ;
        RECT 52.045 165.165 52.830 165.335 ;
        RECT 51.470 164.935 51.640 165.165 ;
        RECT 50.810 164.635 51.640 164.935 ;
        RECT 52.025 164.665 52.490 164.995 ;
        RECT 50.810 164.605 51.010 164.635 ;
        RECT 51.130 164.385 51.300 164.455 ;
        RECT 50.430 164.215 51.300 164.385 ;
        RECT 50.790 164.125 51.300 164.215 ;
        RECT 49.340 163.660 49.645 163.790 ;
        RECT 50.090 163.680 50.620 164.045 ;
        RECT 48.960 163.065 49.225 163.525 ;
        RECT 49.395 163.235 49.645 163.660 ;
        RECT 50.790 163.510 50.960 164.125 ;
        RECT 49.855 163.340 50.960 163.510 ;
        RECT 51.130 163.065 51.300 163.865 ;
        RECT 51.470 163.565 51.640 164.635 ;
        RECT 51.810 163.735 52.000 164.455 ;
        RECT 52.170 163.705 52.490 164.665 ;
        RECT 52.660 164.705 52.830 165.165 ;
        RECT 53.105 165.085 53.315 165.615 ;
        RECT 53.575 164.875 53.905 165.400 ;
        RECT 54.075 165.005 54.245 165.615 ;
        RECT 54.415 164.960 54.745 165.395 ;
        RECT 55.055 165.065 55.225 165.355 ;
        RECT 55.395 165.235 55.725 165.615 ;
        RECT 54.415 164.875 54.795 164.960 ;
        RECT 55.055 164.895 55.720 165.065 ;
        RECT 53.705 164.705 53.905 164.875 ;
        RECT 54.570 164.835 54.795 164.875 ;
        RECT 52.660 164.375 53.535 164.705 ;
        RECT 53.705 164.375 54.455 164.705 ;
        RECT 51.470 163.235 51.720 163.565 ;
        RECT 52.660 163.535 52.830 164.375 ;
        RECT 53.705 164.170 53.895 164.375 ;
        RECT 54.625 164.255 54.795 164.835 ;
        RECT 54.580 164.205 54.795 164.255 ;
        RECT 53.000 163.795 53.895 164.170 ;
        RECT 54.405 164.125 54.795 164.205 ;
        RECT 51.945 163.365 52.830 163.535 ;
        RECT 53.010 163.065 53.325 163.565 ;
        RECT 53.555 163.235 53.895 163.795 ;
        RECT 54.065 163.065 54.235 164.075 ;
        RECT 54.405 163.280 54.735 164.125 ;
        RECT 54.970 164.075 55.320 164.725 ;
        RECT 55.490 163.905 55.720 164.895 ;
        RECT 55.055 163.735 55.720 163.905 ;
        RECT 55.055 163.235 55.225 163.735 ;
        RECT 55.395 163.065 55.725 163.565 ;
        RECT 55.895 163.235 56.080 165.355 ;
        RECT 56.335 165.155 56.585 165.615 ;
        RECT 56.755 165.165 57.090 165.335 ;
        RECT 57.285 165.165 57.960 165.335 ;
        RECT 56.755 165.025 56.925 165.165 ;
        RECT 56.250 164.035 56.530 164.985 ;
        RECT 56.700 164.895 56.925 165.025 ;
        RECT 56.700 163.790 56.870 164.895 ;
        RECT 57.095 164.745 57.620 164.965 ;
        RECT 57.040 163.980 57.280 164.575 ;
        RECT 57.450 164.045 57.620 164.745 ;
        RECT 57.790 164.385 57.960 165.165 ;
        RECT 58.280 165.115 58.650 165.615 ;
        RECT 58.830 165.165 59.235 165.335 ;
        RECT 59.405 165.165 60.190 165.335 ;
        RECT 58.830 164.935 59.000 165.165 ;
        RECT 58.170 164.635 59.000 164.935 ;
        RECT 59.385 164.665 59.850 164.995 ;
        RECT 58.170 164.605 58.370 164.635 ;
        RECT 58.490 164.385 58.660 164.455 ;
        RECT 57.790 164.215 58.660 164.385 ;
        RECT 58.150 164.125 58.660 164.215 ;
        RECT 56.700 163.660 57.005 163.790 ;
        RECT 57.450 163.680 57.980 164.045 ;
        RECT 56.320 163.065 56.585 163.525 ;
        RECT 56.755 163.235 57.005 163.660 ;
        RECT 58.150 163.510 58.320 164.125 ;
        RECT 57.215 163.340 58.320 163.510 ;
        RECT 58.490 163.065 58.660 163.865 ;
        RECT 58.830 163.565 59.000 164.635 ;
        RECT 59.170 163.735 59.360 164.455 ;
        RECT 59.530 163.705 59.850 164.665 ;
        RECT 60.020 164.705 60.190 165.165 ;
        RECT 60.465 165.085 60.675 165.615 ;
        RECT 60.935 164.875 61.265 165.400 ;
        RECT 61.435 165.005 61.605 165.615 ;
        RECT 61.775 164.960 62.105 165.395 ;
        RECT 61.775 164.875 62.155 164.960 ;
        RECT 61.065 164.705 61.265 164.875 ;
        RECT 61.930 164.835 62.155 164.875 ;
        RECT 60.020 164.375 60.895 164.705 ;
        RECT 61.065 164.375 61.815 164.705 ;
        RECT 58.830 163.235 59.080 163.565 ;
        RECT 60.020 163.535 60.190 164.375 ;
        RECT 61.065 164.170 61.255 164.375 ;
        RECT 61.985 164.255 62.155 164.835 ;
        RECT 62.325 164.865 63.535 165.615 ;
        RECT 63.705 164.890 63.995 165.615 ;
        RECT 64.215 164.960 64.545 165.395 ;
        RECT 64.715 165.005 64.885 165.615 ;
        RECT 64.165 164.875 64.545 164.960 ;
        RECT 65.055 164.875 65.385 165.400 ;
        RECT 65.645 165.085 65.855 165.615 ;
        RECT 66.130 165.165 66.915 165.335 ;
        RECT 67.085 165.165 67.490 165.335 ;
        RECT 62.325 164.325 62.845 164.865 ;
        RECT 64.165 164.835 64.390 164.875 ;
        RECT 61.940 164.205 62.155 164.255 ;
        RECT 60.360 163.795 61.255 164.170 ;
        RECT 61.765 164.125 62.155 164.205 ;
        RECT 63.015 164.155 63.535 164.695 ;
        RECT 64.165 164.255 64.335 164.835 ;
        RECT 65.055 164.705 65.255 164.875 ;
        RECT 66.130 164.705 66.300 165.165 ;
        RECT 64.505 164.375 65.255 164.705 ;
        RECT 65.425 164.375 66.300 164.705 ;
        RECT 59.305 163.365 60.190 163.535 ;
        RECT 60.370 163.065 60.685 163.565 ;
        RECT 60.915 163.235 61.255 163.795 ;
        RECT 61.425 163.065 61.595 164.075 ;
        RECT 61.765 163.280 62.095 164.125 ;
        RECT 62.325 163.065 63.535 164.155 ;
        RECT 63.705 163.065 63.995 164.230 ;
        RECT 64.165 164.205 64.380 164.255 ;
        RECT 64.165 164.125 64.555 164.205 ;
        RECT 64.225 163.280 64.555 164.125 ;
        RECT 65.065 164.170 65.255 164.375 ;
        RECT 64.725 163.065 64.895 164.075 ;
        RECT 65.065 163.795 65.960 164.170 ;
        RECT 65.065 163.235 65.405 163.795 ;
        RECT 65.635 163.065 65.950 163.565 ;
        RECT 66.130 163.535 66.300 164.375 ;
        RECT 66.470 164.665 66.935 164.995 ;
        RECT 67.320 164.935 67.490 165.165 ;
        RECT 67.670 165.115 68.040 165.615 ;
        RECT 68.360 165.165 69.035 165.335 ;
        RECT 69.230 165.165 69.565 165.335 ;
        RECT 66.470 163.705 66.790 164.665 ;
        RECT 67.320 164.635 68.150 164.935 ;
        RECT 66.960 163.735 67.150 164.455 ;
        RECT 67.320 163.565 67.490 164.635 ;
        RECT 67.950 164.605 68.150 164.635 ;
        RECT 67.660 164.385 67.830 164.455 ;
        RECT 68.360 164.385 68.530 165.165 ;
        RECT 69.395 165.025 69.565 165.165 ;
        RECT 69.735 165.155 69.985 165.615 ;
        RECT 67.660 164.215 68.530 164.385 ;
        RECT 68.700 164.745 69.225 164.965 ;
        RECT 69.395 164.895 69.620 165.025 ;
        RECT 67.660 164.125 68.170 164.215 ;
        RECT 66.130 163.365 67.015 163.535 ;
        RECT 67.240 163.235 67.490 163.565 ;
        RECT 67.660 163.065 67.830 163.865 ;
        RECT 68.000 163.510 68.170 164.125 ;
        RECT 68.700 164.045 68.870 164.745 ;
        RECT 68.340 163.680 68.870 164.045 ;
        RECT 69.040 163.980 69.280 164.575 ;
        RECT 69.450 163.790 69.620 164.895 ;
        RECT 69.790 164.035 70.070 164.985 ;
        RECT 69.315 163.660 69.620 163.790 ;
        RECT 68.000 163.340 69.105 163.510 ;
        RECT 69.315 163.235 69.565 163.660 ;
        RECT 69.735 163.065 70.000 163.525 ;
        RECT 70.240 163.235 70.425 165.355 ;
        RECT 70.595 165.235 70.925 165.615 ;
        RECT 71.095 165.065 71.265 165.355 ;
        RECT 71.585 165.135 71.865 165.615 ;
        RECT 70.600 164.895 71.265 165.065 ;
        RECT 72.035 164.965 72.295 165.355 ;
        RECT 72.470 165.135 72.725 165.615 ;
        RECT 72.895 164.965 73.190 165.355 ;
        RECT 73.370 165.135 73.645 165.615 ;
        RECT 73.815 165.115 74.115 165.445 ;
        RECT 70.600 163.905 70.830 164.895 ;
        RECT 71.540 164.795 73.190 164.965 ;
        RECT 71.000 164.075 71.350 164.725 ;
        RECT 71.540 164.285 71.945 164.795 ;
        RECT 72.115 164.455 73.255 164.625 ;
        RECT 71.540 164.115 72.295 164.285 ;
        RECT 70.600 163.735 71.265 163.905 ;
        RECT 70.595 163.065 70.925 163.565 ;
        RECT 71.095 163.235 71.265 163.735 ;
        RECT 71.580 163.065 71.865 163.935 ;
        RECT 72.035 163.865 72.295 164.115 ;
        RECT 73.085 164.205 73.255 164.455 ;
        RECT 73.425 164.375 73.775 164.945 ;
        RECT 73.945 164.205 74.115 165.115 ;
        RECT 74.375 165.065 74.545 165.355 ;
        RECT 74.715 165.235 75.045 165.615 ;
        RECT 74.375 164.895 75.040 165.065 ;
        RECT 73.085 164.035 74.115 164.205 ;
        RECT 74.290 164.075 74.640 164.725 ;
        RECT 72.035 163.695 73.155 163.865 ;
        RECT 72.035 163.235 72.295 163.695 ;
        RECT 72.470 163.065 72.725 163.525 ;
        RECT 72.895 163.235 73.155 163.695 ;
        RECT 73.325 163.065 73.635 163.865 ;
        RECT 73.805 163.235 74.115 164.035 ;
        RECT 74.810 163.905 75.040 164.895 ;
        RECT 74.375 163.735 75.040 163.905 ;
        RECT 74.375 163.235 74.545 163.735 ;
        RECT 74.715 163.065 75.045 163.565 ;
        RECT 75.215 163.235 75.400 165.355 ;
        RECT 75.655 165.155 75.905 165.615 ;
        RECT 76.075 165.165 76.410 165.335 ;
        RECT 76.605 165.165 77.280 165.335 ;
        RECT 76.075 165.025 76.245 165.165 ;
        RECT 75.570 164.035 75.850 164.985 ;
        RECT 76.020 164.895 76.245 165.025 ;
        RECT 76.020 163.790 76.190 164.895 ;
        RECT 76.415 164.745 76.940 164.965 ;
        RECT 76.360 163.980 76.600 164.575 ;
        RECT 76.770 164.045 76.940 164.745 ;
        RECT 77.110 164.385 77.280 165.165 ;
        RECT 77.600 165.115 77.970 165.615 ;
        RECT 78.150 165.165 78.555 165.335 ;
        RECT 78.725 165.165 79.510 165.335 ;
        RECT 78.150 164.935 78.320 165.165 ;
        RECT 77.490 164.635 78.320 164.935 ;
        RECT 78.705 164.665 79.170 164.995 ;
        RECT 77.490 164.605 77.690 164.635 ;
        RECT 77.810 164.385 77.980 164.455 ;
        RECT 77.110 164.215 77.980 164.385 ;
        RECT 77.470 164.125 77.980 164.215 ;
        RECT 76.020 163.660 76.325 163.790 ;
        RECT 76.770 163.680 77.300 164.045 ;
        RECT 75.640 163.065 75.905 163.525 ;
        RECT 76.075 163.235 76.325 163.660 ;
        RECT 77.470 163.510 77.640 164.125 ;
        RECT 76.535 163.340 77.640 163.510 ;
        RECT 77.810 163.065 77.980 163.865 ;
        RECT 78.150 163.565 78.320 164.635 ;
        RECT 78.490 163.735 78.680 164.455 ;
        RECT 78.850 163.705 79.170 164.665 ;
        RECT 79.340 164.705 79.510 165.165 ;
        RECT 79.785 165.085 79.995 165.615 ;
        RECT 80.255 164.875 80.585 165.400 ;
        RECT 80.755 165.005 80.925 165.615 ;
        RECT 81.095 164.960 81.425 165.395 ;
        RECT 81.810 165.105 82.050 165.615 ;
        RECT 82.230 165.105 82.510 165.435 ;
        RECT 82.740 165.105 82.955 165.615 ;
        RECT 81.095 164.875 81.475 164.960 ;
        RECT 80.385 164.705 80.585 164.875 ;
        RECT 81.250 164.835 81.475 164.875 ;
        RECT 79.340 164.375 80.215 164.705 ;
        RECT 80.385 164.375 81.135 164.705 ;
        RECT 78.150 163.235 78.400 163.565 ;
        RECT 79.340 163.535 79.510 164.375 ;
        RECT 80.385 164.170 80.575 164.375 ;
        RECT 81.305 164.255 81.475 164.835 ;
        RECT 81.705 164.375 82.060 164.935 ;
        RECT 81.260 164.205 81.475 164.255 ;
        RECT 82.230 164.205 82.400 165.105 ;
        RECT 82.570 164.375 82.835 164.935 ;
        RECT 83.125 164.875 83.740 165.445 ;
        RECT 83.085 164.205 83.255 164.705 ;
        RECT 79.680 163.795 80.575 164.170 ;
        RECT 81.085 164.125 81.475 164.205 ;
        RECT 78.625 163.365 79.510 163.535 ;
        RECT 79.690 163.065 80.005 163.565 ;
        RECT 80.235 163.235 80.575 163.795 ;
        RECT 80.745 163.065 80.915 164.075 ;
        RECT 81.085 163.280 81.415 164.125 ;
        RECT 81.830 164.035 83.255 164.205 ;
        RECT 81.830 163.860 82.220 164.035 ;
        RECT 82.705 163.065 83.035 163.865 ;
        RECT 83.425 163.855 83.740 164.875 ;
        RECT 83.205 163.235 83.740 163.855 ;
        RECT 83.945 164.875 84.205 165.445 ;
        RECT 84.375 165.215 84.760 165.615 ;
        RECT 84.930 165.045 85.185 165.445 ;
        RECT 84.375 164.875 85.185 165.045 ;
        RECT 85.375 164.875 85.620 165.445 ;
        RECT 85.790 165.215 86.175 165.615 ;
        RECT 86.345 165.045 86.600 165.445 ;
        RECT 85.790 164.875 86.600 165.045 ;
        RECT 86.790 164.875 87.215 165.445 ;
        RECT 87.385 165.215 87.770 165.615 ;
        RECT 87.940 165.045 88.375 165.445 ;
        RECT 87.385 164.875 88.375 165.045 ;
        RECT 83.945 164.205 84.130 164.875 ;
        RECT 84.375 164.705 84.725 164.875 ;
        RECT 85.375 164.705 85.545 164.875 ;
        RECT 85.790 164.705 86.140 164.875 ;
        RECT 86.790 164.705 87.140 164.875 ;
        RECT 87.385 164.705 87.720 164.875 ;
        RECT 88.545 164.865 89.755 165.615 ;
        RECT 100.130 165.480 102.050 166.750 ;
        RECT 103.560 166.740 104.120 166.750 ;
        RECT 103.790 165.650 104.120 166.740 ;
        RECT 104.490 166.270 105.530 166.440 ;
        RECT 104.490 165.830 105.530 166.000 ;
        RECT 105.700 165.970 105.870 166.300 ;
        RECT 103.950 165.430 104.120 165.650 ;
        RECT 106.210 165.430 106.380 166.840 ;
        RECT 103.950 165.260 106.380 165.430 ;
        RECT 107.960 167.350 118.590 167.520 ;
        RECT 120.020 176.580 126.250 176.740 ;
        RECT 120.020 174.320 120.690 176.580 ;
        RECT 121.360 176.010 125.400 176.180 ;
        RECT 121.020 174.950 121.190 175.950 ;
        RECT 125.570 174.950 125.740 175.950 ;
        RECT 121.360 174.720 125.400 174.890 ;
        RECT 126.080 174.320 126.250 176.580 ;
        RECT 120.020 174.150 126.250 174.320 ;
        RECT 120.020 170.890 120.690 174.150 ;
        RECT 121.360 173.580 125.400 173.750 ;
        RECT 121.020 171.520 121.190 173.520 ;
        RECT 125.570 171.520 125.740 173.520 ;
        RECT 121.360 171.290 125.400 171.460 ;
        RECT 126.080 170.890 126.250 174.150 ;
        RECT 120.020 170.720 126.250 170.890 ;
        RECT 120.020 167.460 120.690 170.720 ;
        RECT 121.360 170.150 125.400 170.320 ;
        RECT 121.020 168.090 121.190 170.090 ;
        RECT 125.570 168.090 125.740 170.090 ;
        RECT 121.360 167.860 125.400 168.030 ;
        RECT 126.080 167.460 126.250 170.720 ;
        RECT 120.020 167.450 126.250 167.460 ;
        RECT 127.840 176.720 137.670 176.760 ;
        RECT 127.840 176.590 138.470 176.720 ;
        RECT 127.840 174.330 128.010 176.590 ;
        RECT 128.735 176.020 136.775 176.190 ;
        RECT 128.350 174.960 128.520 175.960 ;
        RECT 136.990 174.960 137.160 175.960 ;
        RECT 128.735 174.730 136.775 174.900 ;
        RECT 137.500 174.330 138.470 176.590 ;
        RECT 127.840 174.160 138.470 174.330 ;
        RECT 127.840 170.900 128.010 174.160 ;
        RECT 128.735 173.590 136.775 173.760 ;
        RECT 128.350 171.530 128.520 173.530 ;
        RECT 136.990 171.530 137.160 173.530 ;
        RECT 128.735 171.300 136.775 171.470 ;
        RECT 137.500 170.900 138.470 174.160 ;
        RECT 127.840 170.730 138.470 170.900 ;
        RECT 127.840 167.470 128.010 170.730 ;
        RECT 128.735 170.160 136.775 170.330 ;
        RECT 128.350 168.100 128.520 170.100 ;
        RECT 136.990 168.100 137.160 170.100 ;
        RECT 128.735 167.870 136.775 168.040 ;
        RECT 137.500 167.470 138.470 170.730 ;
        RECT 120.020 167.350 126.260 167.450 ;
        RECT 107.960 165.090 108.130 167.350 ;
        RECT 108.855 166.780 116.895 166.950 ;
        RECT 108.470 165.720 108.640 166.720 ;
        RECT 117.110 165.720 117.280 166.720 ;
        RECT 108.855 165.490 116.895 165.660 ;
        RECT 117.620 165.090 118.590 167.350 ;
        RECT 120.010 166.790 126.260 167.350 ;
        RECT 120.010 166.770 125.180 166.790 ;
        RECT 120.010 166.700 124.000 166.770 ;
        RECT 120.010 165.430 121.930 166.700 ;
        RECT 123.440 166.690 124.000 166.700 ;
        RECT 123.670 165.600 124.000 166.690 ;
        RECT 124.370 166.220 125.410 166.390 ;
        RECT 124.370 165.780 125.410 165.950 ;
        RECT 125.580 165.920 125.750 166.250 ;
        RECT 123.830 165.380 124.000 165.600 ;
        RECT 126.090 165.380 126.260 166.790 ;
        RECT 123.830 165.210 126.260 165.380 ;
        RECT 127.840 167.300 138.470 167.470 ;
        RECT 140.050 176.630 146.280 176.790 ;
        RECT 140.050 174.370 140.720 176.630 ;
        RECT 141.390 176.060 145.430 176.230 ;
        RECT 141.050 175.000 141.220 176.000 ;
        RECT 145.600 175.000 145.770 176.000 ;
        RECT 141.390 174.770 145.430 174.940 ;
        RECT 146.110 174.370 146.280 176.630 ;
        RECT 140.050 174.200 146.280 174.370 ;
        RECT 140.050 170.940 140.720 174.200 ;
        RECT 141.390 173.630 145.430 173.800 ;
        RECT 141.050 171.570 141.220 173.570 ;
        RECT 145.600 171.570 145.770 173.570 ;
        RECT 141.390 171.340 145.430 171.510 ;
        RECT 146.110 170.940 146.280 174.200 ;
        RECT 140.050 170.770 146.280 170.940 ;
        RECT 140.050 167.510 140.720 170.770 ;
        RECT 141.390 170.200 145.430 170.370 ;
        RECT 141.050 168.140 141.220 170.140 ;
        RECT 145.600 168.140 145.770 170.140 ;
        RECT 141.390 167.910 145.430 168.080 ;
        RECT 146.110 167.510 146.280 170.770 ;
        RECT 140.050 167.500 146.280 167.510 ;
        RECT 147.870 176.770 157.700 176.810 ;
        RECT 147.870 176.640 158.500 176.770 ;
        RECT 147.870 174.380 148.040 176.640 ;
        RECT 148.765 176.070 156.805 176.240 ;
        RECT 148.380 175.010 148.550 176.010 ;
        RECT 157.020 175.010 157.190 176.010 ;
        RECT 148.765 174.780 156.805 174.950 ;
        RECT 157.530 174.380 158.500 176.640 ;
        RECT 147.870 174.210 158.500 174.380 ;
        RECT 147.870 170.950 148.040 174.210 ;
        RECT 148.765 173.640 156.805 173.810 ;
        RECT 148.380 171.580 148.550 173.580 ;
        RECT 157.020 171.580 157.190 173.580 ;
        RECT 148.765 171.350 156.805 171.520 ;
        RECT 157.530 170.950 158.500 174.210 ;
        RECT 147.870 170.780 158.500 170.950 ;
        RECT 147.870 167.520 148.040 170.780 ;
        RECT 148.765 170.210 156.805 170.380 ;
        RECT 148.380 168.150 148.550 170.150 ;
        RECT 157.020 168.150 157.190 170.150 ;
        RECT 148.765 167.920 156.805 168.090 ;
        RECT 157.530 167.520 158.500 170.780 ;
        RECT 140.050 167.400 146.290 167.500 ;
        RECT 107.960 165.060 118.590 165.090 ;
        RECT 107.930 164.950 118.590 165.060 ;
        RECT 127.840 165.040 128.010 167.300 ;
        RECT 128.735 166.730 136.775 166.900 ;
        RECT 128.350 165.670 128.520 166.670 ;
        RECT 136.990 165.670 137.160 166.670 ;
        RECT 128.735 165.440 136.775 165.610 ;
        RECT 137.500 165.040 138.470 167.300 ;
        RECT 140.040 166.840 146.290 167.400 ;
        RECT 140.040 166.820 145.210 166.840 ;
        RECT 140.040 166.750 144.030 166.820 ;
        RECT 140.040 165.480 141.960 166.750 ;
        RECT 143.470 166.740 144.030 166.750 ;
        RECT 143.700 165.650 144.030 166.740 ;
        RECT 144.400 166.270 145.440 166.440 ;
        RECT 144.400 165.830 145.440 166.000 ;
        RECT 145.610 165.970 145.780 166.300 ;
        RECT 143.860 165.430 144.030 165.650 ;
        RECT 146.120 165.430 146.290 166.840 ;
        RECT 143.860 165.260 146.290 165.430 ;
        RECT 147.870 167.350 158.500 167.520 ;
        RECT 147.870 165.090 148.040 167.350 ;
        RECT 148.765 166.780 156.805 166.950 ;
        RECT 148.380 165.720 148.550 166.720 ;
        RECT 157.020 165.720 157.190 166.720 ;
        RECT 148.765 165.490 156.805 165.660 ;
        RECT 157.530 165.090 158.500 167.350 ;
        RECT 147.870 165.060 158.500 165.090 ;
        RECT 127.840 165.010 138.470 165.040 ;
        RECT 106.180 164.900 118.590 164.950 ;
        RECT 127.810 164.900 138.470 165.010 ;
        RECT 147.840 164.950 158.500 165.060 ;
        RECT 146.090 164.900 158.500 164.950 ;
        RECT 84.300 164.375 84.725 164.705 ;
        RECT 83.945 163.235 84.205 164.205 ;
        RECT 84.375 163.855 84.725 164.375 ;
        RECT 84.895 164.205 85.545 164.705 ;
        RECT 85.715 164.375 86.140 164.705 ;
        RECT 84.895 164.025 85.620 164.205 ;
        RECT 84.375 163.660 85.185 163.855 ;
        RECT 84.375 163.065 84.760 163.490 ;
        RECT 84.930 163.235 85.185 163.660 ;
        RECT 85.375 163.235 85.620 164.025 ;
        RECT 85.790 163.855 86.140 164.375 ;
        RECT 86.310 164.205 87.140 164.705 ;
        RECT 87.310 164.375 87.720 164.705 ;
        RECT 86.310 164.025 87.215 164.205 ;
        RECT 85.790 163.660 86.620 163.855 ;
        RECT 85.790 163.065 86.175 163.490 ;
        RECT 86.345 163.235 86.620 163.660 ;
        RECT 86.790 163.235 87.215 164.025 ;
        RECT 87.385 163.830 87.720 164.375 ;
        RECT 87.890 164.000 88.375 164.705 ;
        RECT 88.545 164.155 89.065 164.695 ;
        RECT 89.235 164.325 89.755 164.865 ;
        RECT 101.840 164.730 118.590 164.900 ;
        RECT 126.060 164.850 138.470 164.900 ;
        RECT 87.385 163.660 88.375 163.830 ;
        RECT 87.385 163.065 87.770 163.490 ;
        RECT 87.940 163.235 88.375 163.660 ;
        RECT 88.545 163.065 89.755 164.155 ;
        RECT 101.840 163.320 102.010 164.730 ;
        RECT 102.380 164.160 105.420 164.330 ;
        RECT 102.380 163.720 105.420 163.890 ;
        RECT 105.635 163.860 105.805 164.190 ;
        RECT 106.140 163.970 118.590 164.730 ;
        RECT 121.720 164.680 138.470 164.850 ;
        RECT 106.140 163.960 118.480 163.970 ;
        RECT 106.140 163.950 112.020 163.960 ;
        RECT 106.140 163.930 106.710 163.950 ;
        RECT 107.930 163.940 112.020 163.950 ;
        RECT 106.150 163.320 106.320 163.930 ;
        RECT 101.840 163.150 106.320 163.320 ;
        RECT 121.720 163.270 121.890 164.680 ;
        RECT 122.260 164.110 125.300 164.280 ;
        RECT 122.260 163.670 125.300 163.840 ;
        RECT 125.515 163.810 125.685 164.140 ;
        RECT 126.020 163.920 138.470 164.680 ;
        RECT 141.750 164.730 158.500 164.900 ;
        RECT 126.020 163.910 138.360 163.920 ;
        RECT 126.020 163.900 131.900 163.910 ;
        RECT 126.020 163.880 126.590 163.900 ;
        RECT 127.810 163.890 131.900 163.900 ;
        RECT 126.030 163.270 126.200 163.880 ;
        RECT 121.720 163.100 126.200 163.270 ;
        RECT 141.750 163.320 141.920 164.730 ;
        RECT 142.290 164.160 145.330 164.330 ;
        RECT 142.290 163.720 145.330 163.890 ;
        RECT 145.545 163.860 145.715 164.190 ;
        RECT 146.050 163.970 158.500 164.730 ;
        RECT 146.050 163.960 158.390 163.970 ;
        RECT 146.050 163.950 151.930 163.960 ;
        RECT 146.050 163.930 146.620 163.950 ;
        RECT 147.840 163.940 151.930 163.950 ;
        RECT 146.060 163.320 146.230 163.930 ;
        RECT 141.750 163.150 146.230 163.320 ;
        RECT 12.100 162.895 89.840 163.065 ;
        RECT 12.185 161.805 13.395 162.895 ;
        RECT 13.565 162.460 18.910 162.895 ;
        RECT 19.085 162.460 24.430 162.895 ;
        RECT 12.185 161.095 12.705 161.635 ;
        RECT 12.875 161.265 13.395 161.805 ;
        RECT 12.185 160.345 13.395 161.095 ;
        RECT 15.150 160.890 15.490 161.720 ;
        RECT 16.970 161.210 17.320 162.460 ;
        RECT 20.670 160.890 21.010 161.720 ;
        RECT 22.490 161.210 22.840 162.460 ;
        RECT 25.065 161.730 25.355 162.895 ;
        RECT 25.525 162.460 30.870 162.895 ;
        RECT 31.045 162.460 36.390 162.895 ;
        RECT 13.565 160.345 18.910 160.890 ;
        RECT 19.085 160.345 24.430 160.890 ;
        RECT 25.065 160.345 25.355 161.070 ;
        RECT 27.110 160.890 27.450 161.720 ;
        RECT 28.930 161.210 29.280 162.460 ;
        RECT 32.630 160.890 32.970 161.720 ;
        RECT 34.450 161.210 34.800 162.460 ;
        RECT 37.085 161.835 37.415 162.680 ;
        RECT 37.585 161.885 37.755 162.895 ;
        RECT 37.925 162.165 38.265 162.725 ;
        RECT 38.495 162.395 38.810 162.895 ;
        RECT 38.990 162.425 39.875 162.595 ;
        RECT 37.025 161.755 37.415 161.835 ;
        RECT 37.925 161.790 38.820 162.165 ;
        RECT 37.025 161.705 37.240 161.755 ;
        RECT 37.025 161.125 37.195 161.705 ;
        RECT 37.925 161.585 38.115 161.790 ;
        RECT 38.990 161.585 39.160 162.425 ;
        RECT 40.100 162.395 40.350 162.725 ;
        RECT 37.365 161.255 38.115 161.585 ;
        RECT 38.285 161.255 39.160 161.585 ;
        RECT 37.025 161.085 37.250 161.125 ;
        RECT 37.915 161.085 38.115 161.255 ;
        RECT 37.025 161.000 37.405 161.085 ;
        RECT 25.525 160.345 30.870 160.890 ;
        RECT 31.045 160.345 36.390 160.890 ;
        RECT 37.075 160.565 37.405 161.000 ;
        RECT 37.575 160.345 37.745 160.955 ;
        RECT 37.915 160.560 38.245 161.085 ;
        RECT 38.505 160.345 38.715 160.875 ;
        RECT 38.990 160.795 39.160 161.255 ;
        RECT 39.330 161.295 39.650 162.255 ;
        RECT 39.820 161.505 40.010 162.225 ;
        RECT 40.180 161.325 40.350 162.395 ;
        RECT 40.520 162.095 40.690 162.895 ;
        RECT 40.860 162.450 41.965 162.620 ;
        RECT 40.860 161.835 41.030 162.450 ;
        RECT 42.175 162.300 42.425 162.725 ;
        RECT 42.595 162.435 42.860 162.895 ;
        RECT 41.200 161.915 41.730 162.280 ;
        RECT 42.175 162.170 42.480 162.300 ;
        RECT 40.520 161.745 41.030 161.835 ;
        RECT 40.520 161.575 41.390 161.745 ;
        RECT 40.520 161.505 40.690 161.575 ;
        RECT 40.810 161.325 41.010 161.355 ;
        RECT 39.330 160.965 39.795 161.295 ;
        RECT 40.180 161.025 41.010 161.325 ;
        RECT 40.180 160.795 40.350 161.025 ;
        RECT 38.990 160.625 39.775 160.795 ;
        RECT 39.945 160.625 40.350 160.795 ;
        RECT 40.530 160.345 40.900 160.845 ;
        RECT 41.220 160.795 41.390 161.575 ;
        RECT 41.560 161.215 41.730 161.915 ;
        RECT 41.900 161.385 42.140 161.980 ;
        RECT 41.560 160.995 42.085 161.215 ;
        RECT 42.310 161.065 42.480 162.170 ;
        RECT 42.255 160.935 42.480 161.065 ;
        RECT 42.650 160.975 42.930 161.925 ;
        RECT 42.255 160.795 42.425 160.935 ;
        RECT 41.220 160.625 41.895 160.795 ;
        RECT 42.090 160.625 42.425 160.795 ;
        RECT 42.595 160.345 42.845 160.805 ;
        RECT 43.100 160.605 43.285 162.725 ;
        RECT 43.455 162.395 43.785 162.895 ;
        RECT 43.955 162.225 44.125 162.725 ;
        RECT 44.585 162.225 44.865 162.895 ;
        RECT 43.460 162.055 44.125 162.225 ;
        RECT 43.460 161.065 43.690 162.055 ;
        RECT 45.035 162.005 45.335 162.555 ;
        RECT 45.535 162.175 45.865 162.895 ;
        RECT 46.055 162.175 46.515 162.725 ;
        RECT 43.860 161.235 44.210 161.885 ;
        RECT 44.400 161.585 44.665 161.945 ;
        RECT 45.035 161.835 45.975 162.005 ;
        RECT 45.805 161.585 45.975 161.835 ;
        RECT 44.400 161.335 45.075 161.585 ;
        RECT 45.295 161.335 45.635 161.585 ;
        RECT 45.805 161.255 46.095 161.585 ;
        RECT 45.805 161.165 45.975 161.255 ;
        RECT 43.460 160.895 44.125 161.065 ;
        RECT 43.455 160.345 43.785 160.725 ;
        RECT 43.955 160.605 44.125 160.895 ;
        RECT 44.585 160.975 45.975 161.165 ;
        RECT 44.585 160.615 44.915 160.975 ;
        RECT 46.265 160.805 46.515 162.175 ;
        RECT 45.535 160.345 45.785 160.805 ;
        RECT 45.955 160.515 46.515 160.805 ;
        RECT 46.685 161.755 47.070 162.715 ;
        RECT 47.285 162.095 47.575 162.895 ;
        RECT 47.745 162.555 49.110 162.725 ;
        RECT 47.745 161.925 47.915 162.555 ;
        RECT 47.240 161.755 47.915 161.925 ;
        RECT 46.685 161.085 46.860 161.755 ;
        RECT 47.240 161.585 47.410 161.755 ;
        RECT 48.085 161.585 48.410 162.385 ;
        RECT 48.780 162.345 49.110 162.555 ;
        RECT 48.780 162.095 49.735 162.345 ;
        RECT 47.045 161.335 47.410 161.585 ;
        RECT 47.605 161.335 47.855 161.585 ;
        RECT 47.045 161.255 47.235 161.335 ;
        RECT 47.605 161.255 47.775 161.335 ;
        RECT 48.065 161.255 48.410 161.585 ;
        RECT 48.580 161.255 48.855 161.920 ;
        RECT 49.040 161.255 49.395 161.920 ;
        RECT 49.565 161.085 49.735 162.095 ;
        RECT 49.905 161.755 50.195 162.895 ;
        RECT 50.825 161.730 51.115 162.895 ;
        RECT 51.290 161.945 51.555 162.715 ;
        RECT 51.725 162.175 52.055 162.895 ;
        RECT 52.245 162.355 52.505 162.715 ;
        RECT 52.675 162.525 53.005 162.895 ;
        RECT 53.175 162.355 53.435 162.715 ;
        RECT 52.245 162.125 53.435 162.355 ;
        RECT 54.005 161.945 54.295 162.715 ;
        RECT 49.920 161.255 50.195 161.585 ;
        RECT 46.685 160.515 47.195 161.085 ;
        RECT 47.740 160.915 49.140 161.085 ;
        RECT 47.365 160.345 47.535 160.905 ;
        RECT 47.740 160.515 48.070 160.915 ;
        RECT 48.245 160.345 48.575 160.745 ;
        RECT 48.810 160.725 49.140 160.915 ;
        RECT 49.310 160.895 49.735 161.085 ;
        RECT 49.905 160.725 50.195 160.995 ;
        RECT 48.810 160.515 50.195 160.725 ;
        RECT 50.825 160.345 51.115 161.070 ;
        RECT 51.290 160.525 51.625 161.945 ;
        RECT 51.800 161.765 54.295 161.945 ;
        RECT 51.800 161.075 52.025 161.765 ;
        RECT 54.505 161.755 54.775 162.725 ;
        RECT 54.985 162.095 55.265 162.895 ;
        RECT 55.435 162.385 57.090 162.675 ;
        RECT 55.500 162.045 57.090 162.215 ;
        RECT 55.500 161.925 55.670 162.045 ;
        RECT 54.945 161.755 55.670 161.925 ;
        RECT 52.225 161.255 52.505 161.585 ;
        RECT 52.685 161.255 53.260 161.585 ;
        RECT 53.440 161.255 53.875 161.585 ;
        RECT 54.055 161.255 54.325 161.585 ;
        RECT 51.800 160.885 54.285 161.075 ;
        RECT 51.805 160.345 52.550 160.715 ;
        RECT 53.115 160.525 53.370 160.885 ;
        RECT 53.550 160.345 53.880 160.715 ;
        RECT 54.060 160.525 54.285 160.885 ;
        RECT 54.505 161.020 54.675 161.755 ;
        RECT 54.945 161.585 55.115 161.755 ;
        RECT 55.860 161.705 56.575 161.875 ;
        RECT 56.770 161.755 57.090 162.045 ;
        RECT 57.270 161.755 57.605 162.725 ;
        RECT 57.775 161.755 57.945 162.895 ;
        RECT 58.115 162.555 60.145 162.725 ;
        RECT 54.845 161.255 55.115 161.585 ;
        RECT 55.285 161.255 55.690 161.585 ;
        RECT 55.860 161.255 56.570 161.705 ;
        RECT 54.945 161.085 55.115 161.255 ;
        RECT 54.505 160.675 54.775 161.020 ;
        RECT 54.945 160.915 56.555 161.085 ;
        RECT 56.740 161.015 57.090 161.585 ;
        RECT 57.270 161.085 57.440 161.755 ;
        RECT 58.115 161.585 58.285 162.555 ;
        RECT 57.610 161.255 57.865 161.585 ;
        RECT 58.090 161.255 58.285 161.585 ;
        RECT 58.455 162.215 59.580 162.385 ;
        RECT 57.695 161.085 57.865 161.255 ;
        RECT 58.455 161.085 58.625 162.215 ;
        RECT 54.965 160.345 55.345 160.745 ;
        RECT 55.515 160.565 55.685 160.915 ;
        RECT 55.855 160.345 56.185 160.745 ;
        RECT 56.385 160.565 56.555 160.915 ;
        RECT 56.755 160.345 57.085 160.845 ;
        RECT 57.270 160.515 57.525 161.085 ;
        RECT 57.695 160.915 58.625 161.085 ;
        RECT 58.795 161.875 59.805 162.045 ;
        RECT 58.795 161.075 58.965 161.875 ;
        RECT 59.170 161.535 59.445 161.675 ;
        RECT 59.165 161.365 59.445 161.535 ;
        RECT 58.450 160.880 58.625 160.915 ;
        RECT 57.695 160.345 58.025 160.745 ;
        RECT 58.450 160.515 58.980 160.880 ;
        RECT 59.170 160.515 59.445 161.365 ;
        RECT 59.615 160.515 59.805 161.875 ;
        RECT 59.975 161.890 60.145 162.555 ;
        RECT 60.315 162.135 60.485 162.895 ;
        RECT 60.720 162.135 61.235 162.545 ;
        RECT 59.975 161.700 60.725 161.890 ;
        RECT 60.895 161.325 61.235 162.135 ;
        RECT 61.495 162.225 61.665 162.725 ;
        RECT 61.835 162.395 62.165 162.895 ;
        RECT 61.495 162.055 62.160 162.225 ;
        RECT 60.005 161.155 61.235 161.325 ;
        RECT 61.410 161.235 61.760 161.885 ;
        RECT 59.985 160.345 60.495 160.880 ;
        RECT 60.715 160.550 60.960 161.155 ;
        RECT 61.930 161.065 62.160 162.055 ;
        RECT 61.495 160.895 62.160 161.065 ;
        RECT 61.495 160.605 61.665 160.895 ;
        RECT 61.835 160.345 62.165 160.725 ;
        RECT 62.335 160.605 62.520 162.725 ;
        RECT 62.760 162.435 63.025 162.895 ;
        RECT 63.195 162.300 63.445 162.725 ;
        RECT 63.655 162.450 64.760 162.620 ;
        RECT 63.140 162.170 63.445 162.300 ;
        RECT 62.690 160.975 62.970 161.925 ;
        RECT 63.140 161.065 63.310 162.170 ;
        RECT 63.480 161.385 63.720 161.980 ;
        RECT 63.890 161.915 64.420 162.280 ;
        RECT 63.890 161.215 64.060 161.915 ;
        RECT 64.590 161.835 64.760 162.450 ;
        RECT 64.930 162.095 65.100 162.895 ;
        RECT 65.270 162.395 65.520 162.725 ;
        RECT 65.745 162.425 66.630 162.595 ;
        RECT 64.590 161.745 65.100 161.835 ;
        RECT 63.140 160.935 63.365 161.065 ;
        RECT 63.535 160.995 64.060 161.215 ;
        RECT 64.230 161.575 65.100 161.745 ;
        RECT 62.775 160.345 63.025 160.805 ;
        RECT 63.195 160.795 63.365 160.935 ;
        RECT 64.230 160.795 64.400 161.575 ;
        RECT 64.930 161.505 65.100 161.575 ;
        RECT 64.610 161.325 64.810 161.355 ;
        RECT 65.270 161.325 65.440 162.395 ;
        RECT 65.610 161.505 65.800 162.225 ;
        RECT 64.610 161.025 65.440 161.325 ;
        RECT 65.970 161.295 66.290 162.255 ;
        RECT 63.195 160.625 63.530 160.795 ;
        RECT 63.725 160.625 64.400 160.795 ;
        RECT 64.720 160.345 65.090 160.845 ;
        RECT 65.270 160.795 65.440 161.025 ;
        RECT 65.825 160.965 66.290 161.295 ;
        RECT 66.460 161.585 66.630 162.425 ;
        RECT 66.810 162.395 67.125 162.895 ;
        RECT 67.355 162.165 67.695 162.725 ;
        RECT 66.800 161.790 67.695 162.165 ;
        RECT 67.865 161.885 68.035 162.895 ;
        RECT 67.505 161.585 67.695 161.790 ;
        RECT 68.205 161.835 68.535 162.680 ;
        RECT 68.205 161.755 68.595 161.835 ;
        RECT 68.380 161.705 68.595 161.755 ;
        RECT 66.460 161.255 67.335 161.585 ;
        RECT 67.505 161.255 68.255 161.585 ;
        RECT 66.460 160.795 66.630 161.255 ;
        RECT 67.505 161.085 67.705 161.255 ;
        RECT 68.425 161.125 68.595 161.705 ;
        RECT 68.370 161.085 68.595 161.125 ;
        RECT 65.270 160.625 65.675 160.795 ;
        RECT 65.845 160.625 66.630 160.795 ;
        RECT 66.905 160.345 67.115 160.875 ;
        RECT 67.375 160.560 67.705 161.085 ;
        RECT 68.215 161.000 68.595 161.085 ;
        RECT 68.770 161.755 69.105 162.725 ;
        RECT 69.275 161.755 69.445 162.895 ;
        RECT 69.615 162.555 71.645 162.725 ;
        RECT 68.770 161.085 68.940 161.755 ;
        RECT 69.615 161.585 69.785 162.555 ;
        RECT 69.110 161.255 69.365 161.585 ;
        RECT 69.590 161.255 69.785 161.585 ;
        RECT 69.955 162.215 71.080 162.385 ;
        RECT 69.195 161.085 69.365 161.255 ;
        RECT 69.955 161.085 70.125 162.215 ;
        RECT 67.875 160.345 68.045 160.955 ;
        RECT 68.215 160.565 68.545 161.000 ;
        RECT 68.770 160.515 69.025 161.085 ;
        RECT 69.195 160.915 70.125 161.085 ;
        RECT 70.295 161.875 71.305 162.045 ;
        RECT 70.295 161.075 70.465 161.875 ;
        RECT 70.670 161.195 70.945 161.675 ;
        RECT 70.665 161.025 70.945 161.195 ;
        RECT 69.950 160.880 70.125 160.915 ;
        RECT 69.195 160.345 69.525 160.745 ;
        RECT 69.950 160.515 70.480 160.880 ;
        RECT 70.670 160.515 70.945 161.025 ;
        RECT 71.115 160.515 71.305 161.875 ;
        RECT 71.475 161.890 71.645 162.555 ;
        RECT 71.815 162.135 71.985 162.895 ;
        RECT 72.220 162.135 72.735 162.545 ;
        RECT 71.475 161.700 72.225 161.890 ;
        RECT 72.395 161.325 72.735 162.135 ;
        RECT 71.505 161.155 72.735 161.325 ;
        RECT 72.905 161.755 73.290 162.725 ;
        RECT 73.460 162.435 73.785 162.895 ;
        RECT 74.305 162.265 74.585 162.725 ;
        RECT 73.460 162.045 74.585 162.265 ;
        RECT 71.485 160.345 71.995 160.880 ;
        RECT 72.215 160.550 72.460 161.155 ;
        RECT 72.905 161.085 73.185 161.755 ;
        RECT 73.460 161.585 73.910 162.045 ;
        RECT 74.775 161.875 75.175 162.725 ;
        RECT 75.575 162.435 75.845 162.895 ;
        RECT 76.015 162.265 76.300 162.725 ;
        RECT 73.355 161.255 73.910 161.585 ;
        RECT 74.080 161.315 75.175 161.875 ;
        RECT 73.460 161.145 73.910 161.255 ;
        RECT 72.905 160.515 73.290 161.085 ;
        RECT 73.460 160.975 74.585 161.145 ;
        RECT 73.460 160.345 73.785 160.805 ;
        RECT 74.305 160.515 74.585 160.975 ;
        RECT 74.775 160.515 75.175 161.315 ;
        RECT 75.345 162.045 76.300 162.265 ;
        RECT 75.345 161.145 75.555 162.045 ;
        RECT 75.725 161.315 76.415 161.875 ;
        RECT 76.585 161.730 76.875 162.895 ;
        RECT 77.045 161.755 77.385 162.725 ;
        RECT 77.555 161.755 77.725 162.895 ;
        RECT 77.995 162.095 78.245 162.895 ;
        RECT 78.890 161.925 79.220 162.725 ;
        RECT 79.520 162.095 79.850 162.895 ;
        RECT 80.020 161.925 80.350 162.725 ;
        RECT 81.275 162.225 81.445 162.725 ;
        RECT 81.615 162.395 81.945 162.895 ;
        RECT 81.275 162.055 81.940 162.225 ;
        RECT 77.915 161.755 80.350 161.925 ;
        RECT 77.045 161.195 77.220 161.755 ;
        RECT 77.915 161.505 78.085 161.755 ;
        RECT 77.390 161.335 78.085 161.505 ;
        RECT 78.260 161.335 78.680 161.535 ;
        RECT 78.850 161.335 79.180 161.535 ;
        RECT 79.350 161.335 79.680 161.535 ;
        RECT 77.045 161.145 77.275 161.195 ;
        RECT 75.345 160.975 76.300 161.145 ;
        RECT 75.575 160.345 75.845 160.805 ;
        RECT 76.015 160.515 76.300 160.975 ;
        RECT 76.585 160.345 76.875 161.070 ;
        RECT 77.045 160.515 77.385 161.145 ;
        RECT 77.555 160.345 77.805 161.145 ;
        RECT 77.995 160.995 79.220 161.165 ;
        RECT 77.995 160.515 78.325 160.995 ;
        RECT 78.495 160.345 78.720 160.805 ;
        RECT 78.890 160.515 79.220 160.995 ;
        RECT 79.850 161.125 80.020 161.755 ;
        RECT 80.205 161.335 80.555 161.585 ;
        RECT 81.190 161.235 81.540 161.885 ;
        RECT 79.850 160.515 80.350 161.125 ;
        RECT 81.710 161.065 81.940 162.055 ;
        RECT 81.275 160.895 81.940 161.065 ;
        RECT 81.275 160.605 81.445 160.895 ;
        RECT 81.615 160.345 81.945 160.725 ;
        RECT 82.115 160.605 82.300 162.725 ;
        RECT 82.540 162.435 82.805 162.895 ;
        RECT 82.975 162.300 83.225 162.725 ;
        RECT 83.435 162.450 84.540 162.620 ;
        RECT 82.920 162.170 83.225 162.300 ;
        RECT 82.470 160.975 82.750 161.925 ;
        RECT 82.920 161.065 83.090 162.170 ;
        RECT 83.260 161.385 83.500 161.980 ;
        RECT 83.670 161.915 84.200 162.280 ;
        RECT 83.670 161.215 83.840 161.915 ;
        RECT 84.370 161.835 84.540 162.450 ;
        RECT 84.710 162.095 84.880 162.895 ;
        RECT 85.050 162.395 85.300 162.725 ;
        RECT 85.525 162.425 86.410 162.595 ;
        RECT 84.370 161.745 84.880 161.835 ;
        RECT 82.920 160.935 83.145 161.065 ;
        RECT 83.315 160.995 83.840 161.215 ;
        RECT 84.010 161.575 84.880 161.745 ;
        RECT 82.555 160.345 82.805 160.805 ;
        RECT 82.975 160.795 83.145 160.935 ;
        RECT 84.010 160.795 84.180 161.575 ;
        RECT 84.710 161.505 84.880 161.575 ;
        RECT 84.390 161.325 84.590 161.355 ;
        RECT 85.050 161.325 85.220 162.395 ;
        RECT 85.390 161.505 85.580 162.225 ;
        RECT 84.390 161.025 85.220 161.325 ;
        RECT 85.750 161.295 86.070 162.255 ;
        RECT 82.975 160.625 83.310 160.795 ;
        RECT 83.505 160.625 84.180 160.795 ;
        RECT 84.500 160.345 84.870 160.845 ;
        RECT 85.050 160.795 85.220 161.025 ;
        RECT 85.605 160.965 86.070 161.295 ;
        RECT 86.240 161.585 86.410 162.425 ;
        RECT 86.590 162.395 86.905 162.895 ;
        RECT 87.135 162.165 87.475 162.725 ;
        RECT 86.580 161.790 87.475 162.165 ;
        RECT 87.645 161.885 87.815 162.895 ;
        RECT 87.285 161.585 87.475 161.790 ;
        RECT 87.985 161.835 88.315 162.680 ;
        RECT 87.985 161.755 88.375 161.835 ;
        RECT 88.160 161.705 88.375 161.755 ;
        RECT 86.240 161.255 87.115 161.585 ;
        RECT 87.285 161.255 88.035 161.585 ;
        RECT 86.240 160.795 86.410 161.255 ;
        RECT 87.285 161.085 87.485 161.255 ;
        RECT 88.205 161.125 88.375 161.705 ;
        RECT 88.545 161.805 89.755 162.895 ;
        RECT 88.545 161.265 89.065 161.805 ;
        RECT 100.630 161.790 106.370 161.800 ;
        RECT 88.150 161.085 88.375 161.125 ;
        RECT 89.235 161.095 89.755 161.635 ;
        RECT 85.050 160.625 85.455 160.795 ;
        RECT 85.625 160.625 86.410 160.795 ;
        RECT 86.685 160.345 86.895 160.875 ;
        RECT 87.155 160.560 87.485 161.085 ;
        RECT 87.995 161.000 88.375 161.085 ;
        RECT 87.655 160.345 87.825 160.955 ;
        RECT 87.995 160.565 88.325 161.000 ;
        RECT 88.545 160.345 89.755 161.095 ;
        RECT 100.140 161.630 106.370 161.790 ;
        RECT 12.100 160.175 89.840 160.345 ;
        RECT 12.185 159.425 13.395 160.175 ;
        RECT 13.565 159.630 18.910 160.175 ;
        RECT 19.085 159.630 24.430 160.175 ;
        RECT 24.605 159.630 29.950 160.175 ;
        RECT 12.185 158.885 12.705 159.425 ;
        RECT 12.875 158.715 13.395 159.255 ;
        RECT 15.150 158.800 15.490 159.630 ;
        RECT 12.185 157.625 13.395 158.715 ;
        RECT 16.970 158.060 17.320 159.310 ;
        RECT 20.670 158.800 21.010 159.630 ;
        RECT 22.490 158.060 22.840 159.310 ;
        RECT 26.190 158.800 26.530 159.630 ;
        RECT 30.125 159.405 33.635 160.175 ;
        RECT 28.010 158.060 28.360 159.310 ;
        RECT 30.125 158.885 31.775 159.405 ;
        RECT 33.805 159.375 34.115 160.175 ;
        RECT 34.320 159.375 35.015 160.005 ;
        RECT 31.945 158.715 33.635 159.235 ;
        RECT 33.815 158.935 34.150 159.205 ;
        RECT 34.320 158.775 34.490 159.375 ;
        RECT 34.660 158.935 34.995 159.185 ;
        RECT 13.565 157.625 18.910 158.060 ;
        RECT 19.085 157.625 24.430 158.060 ;
        RECT 24.605 157.625 29.950 158.060 ;
        RECT 30.125 157.625 33.635 158.715 ;
        RECT 33.805 157.625 34.085 158.765 ;
        RECT 34.255 157.795 34.585 158.775 ;
        RECT 34.755 157.625 35.015 158.765 ;
        RECT 35.195 157.805 35.455 159.995 ;
        RECT 35.715 159.805 36.385 160.175 ;
        RECT 36.565 159.625 36.875 159.995 ;
        RECT 35.645 159.425 36.875 159.625 ;
        RECT 35.645 158.755 35.935 159.425 ;
        RECT 37.055 159.245 37.285 159.885 ;
        RECT 37.465 159.445 37.755 160.175 ;
        RECT 37.945 159.450 38.235 160.175 ;
        RECT 38.495 159.625 38.665 159.915 ;
        RECT 38.835 159.795 39.165 160.175 ;
        RECT 38.495 159.455 39.160 159.625 ;
        RECT 36.115 158.935 36.580 159.245 ;
        RECT 36.760 158.935 37.285 159.245 ;
        RECT 37.465 158.935 37.765 159.265 ;
        RECT 35.645 158.535 36.415 158.755 ;
        RECT 35.625 157.625 35.965 158.355 ;
        RECT 36.145 157.805 36.415 158.535 ;
        RECT 36.595 158.515 37.755 158.755 ;
        RECT 36.595 157.805 36.825 158.515 ;
        RECT 36.995 157.625 37.325 158.335 ;
        RECT 37.495 157.805 37.755 158.515 ;
        RECT 37.945 157.625 38.235 158.790 ;
        RECT 38.410 158.635 38.760 159.285 ;
        RECT 38.930 158.465 39.160 159.455 ;
        RECT 38.495 158.295 39.160 158.465 ;
        RECT 38.495 157.795 38.665 158.295 ;
        RECT 38.835 157.625 39.165 158.125 ;
        RECT 39.335 157.795 39.520 159.915 ;
        RECT 39.775 159.715 40.025 160.175 ;
        RECT 40.195 159.725 40.530 159.895 ;
        RECT 40.725 159.725 41.400 159.895 ;
        RECT 40.195 159.585 40.365 159.725 ;
        RECT 39.690 158.595 39.970 159.545 ;
        RECT 40.140 159.455 40.365 159.585 ;
        RECT 40.140 158.350 40.310 159.455 ;
        RECT 40.535 159.305 41.060 159.525 ;
        RECT 40.480 158.540 40.720 159.135 ;
        RECT 40.890 158.605 41.060 159.305 ;
        RECT 41.230 158.945 41.400 159.725 ;
        RECT 41.720 159.675 42.090 160.175 ;
        RECT 42.270 159.725 42.675 159.895 ;
        RECT 42.845 159.725 43.630 159.895 ;
        RECT 42.270 159.495 42.440 159.725 ;
        RECT 41.610 159.195 42.440 159.495 ;
        RECT 42.825 159.225 43.290 159.555 ;
        RECT 41.610 159.165 41.810 159.195 ;
        RECT 41.930 158.945 42.100 159.015 ;
        RECT 41.230 158.775 42.100 158.945 ;
        RECT 41.590 158.685 42.100 158.775 ;
        RECT 40.140 158.220 40.445 158.350 ;
        RECT 40.890 158.240 41.420 158.605 ;
        RECT 39.760 157.625 40.025 158.085 ;
        RECT 40.195 157.795 40.445 158.220 ;
        RECT 41.590 158.070 41.760 158.685 ;
        RECT 40.655 157.900 41.760 158.070 ;
        RECT 41.930 157.625 42.100 158.425 ;
        RECT 42.270 158.125 42.440 159.195 ;
        RECT 42.610 158.295 42.800 159.015 ;
        RECT 42.970 158.265 43.290 159.225 ;
        RECT 43.460 159.265 43.630 159.725 ;
        RECT 43.905 159.645 44.115 160.175 ;
        RECT 44.375 159.435 44.705 159.960 ;
        RECT 44.875 159.565 45.045 160.175 ;
        RECT 45.215 159.520 45.545 159.955 ;
        RECT 46.315 159.625 46.485 159.915 ;
        RECT 46.655 159.795 46.985 160.175 ;
        RECT 45.215 159.435 45.595 159.520 ;
        RECT 46.315 159.455 46.980 159.625 ;
        RECT 44.505 159.265 44.705 159.435 ;
        RECT 45.370 159.395 45.595 159.435 ;
        RECT 43.460 158.935 44.335 159.265 ;
        RECT 44.505 158.935 45.255 159.265 ;
        RECT 42.270 157.795 42.520 158.125 ;
        RECT 43.460 158.095 43.630 158.935 ;
        RECT 44.505 158.730 44.695 158.935 ;
        RECT 45.425 158.815 45.595 159.395 ;
        RECT 45.380 158.765 45.595 158.815 ;
        RECT 43.800 158.355 44.695 158.730 ;
        RECT 45.205 158.685 45.595 158.765 ;
        RECT 42.745 157.925 43.630 158.095 ;
        RECT 43.810 157.625 44.125 158.125 ;
        RECT 44.355 157.795 44.695 158.355 ;
        RECT 44.865 157.625 45.035 158.635 ;
        RECT 45.205 157.840 45.535 158.685 ;
        RECT 46.230 158.635 46.580 159.285 ;
        RECT 46.750 158.465 46.980 159.455 ;
        RECT 46.315 158.295 46.980 158.465 ;
        RECT 46.315 157.795 46.485 158.295 ;
        RECT 46.655 157.625 46.985 158.125 ;
        RECT 47.155 157.795 47.340 159.915 ;
        RECT 47.595 159.715 47.845 160.175 ;
        RECT 48.015 159.725 48.350 159.895 ;
        RECT 48.545 159.725 49.220 159.895 ;
        RECT 48.015 159.585 48.185 159.725 ;
        RECT 47.510 158.595 47.790 159.545 ;
        RECT 47.960 159.455 48.185 159.585 ;
        RECT 47.960 158.350 48.130 159.455 ;
        RECT 48.355 159.305 48.880 159.525 ;
        RECT 48.300 158.540 48.540 159.135 ;
        RECT 48.710 158.605 48.880 159.305 ;
        RECT 49.050 158.945 49.220 159.725 ;
        RECT 49.540 159.675 49.910 160.175 ;
        RECT 50.090 159.725 50.495 159.895 ;
        RECT 50.665 159.725 51.450 159.895 ;
        RECT 50.090 159.495 50.260 159.725 ;
        RECT 49.430 159.195 50.260 159.495 ;
        RECT 50.645 159.225 51.110 159.555 ;
        RECT 49.430 159.165 49.630 159.195 ;
        RECT 49.750 158.945 49.920 159.015 ;
        RECT 49.050 158.775 49.920 158.945 ;
        RECT 49.410 158.685 49.920 158.775 ;
        RECT 47.960 158.220 48.265 158.350 ;
        RECT 48.710 158.240 49.240 158.605 ;
        RECT 47.580 157.625 47.845 158.085 ;
        RECT 48.015 157.795 48.265 158.220 ;
        RECT 49.410 158.070 49.580 158.685 ;
        RECT 48.475 157.900 49.580 158.070 ;
        RECT 49.750 157.625 49.920 158.425 ;
        RECT 50.090 158.125 50.260 159.195 ;
        RECT 50.430 158.295 50.620 159.015 ;
        RECT 50.790 158.265 51.110 159.225 ;
        RECT 51.280 159.265 51.450 159.725 ;
        RECT 51.725 159.645 51.935 160.175 ;
        RECT 52.195 159.435 52.525 159.960 ;
        RECT 52.695 159.565 52.865 160.175 ;
        RECT 53.035 159.520 53.365 159.955 ;
        RECT 53.585 159.675 53.925 160.175 ;
        RECT 53.035 159.435 53.415 159.520 ;
        RECT 52.325 159.265 52.525 159.435 ;
        RECT 53.190 159.395 53.415 159.435 ;
        RECT 51.280 158.935 52.155 159.265 ;
        RECT 52.325 158.935 53.075 159.265 ;
        RECT 50.090 157.795 50.340 158.125 ;
        RECT 51.280 158.095 51.450 158.935 ;
        RECT 52.325 158.730 52.515 158.935 ;
        RECT 53.245 158.815 53.415 159.395 ;
        RECT 53.585 158.935 53.925 159.505 ;
        RECT 54.095 159.265 54.340 159.955 ;
        RECT 54.535 159.675 54.865 160.175 ;
        RECT 55.065 159.605 55.235 159.955 ;
        RECT 55.410 159.775 55.740 160.175 ;
        RECT 55.910 159.605 56.080 159.955 ;
        RECT 56.250 159.775 56.630 160.175 ;
        RECT 55.065 159.435 56.650 159.605 ;
        RECT 56.820 159.500 57.095 159.845 ;
        RECT 56.480 159.265 56.650 159.435 ;
        RECT 54.095 158.935 54.750 159.265 ;
        RECT 53.200 158.765 53.415 158.815 ;
        RECT 51.620 158.355 52.515 158.730 ;
        RECT 53.025 158.685 53.415 158.765 ;
        RECT 50.565 157.925 51.450 158.095 ;
        RECT 51.630 157.625 51.945 158.125 ;
        RECT 52.175 157.795 52.515 158.355 ;
        RECT 52.685 157.625 52.855 158.635 ;
        RECT 53.025 157.840 53.355 158.685 ;
        RECT 53.585 157.625 53.925 158.700 ;
        RECT 54.095 158.340 54.335 158.935 ;
        RECT 54.530 158.475 54.850 158.765 ;
        RECT 55.020 158.645 55.760 159.265 ;
        RECT 55.930 158.935 56.310 159.265 ;
        RECT 56.480 158.935 56.755 159.265 ;
        RECT 56.480 158.765 56.650 158.935 ;
        RECT 56.925 158.765 57.095 159.500 ;
        RECT 55.990 158.595 56.650 158.765 ;
        RECT 55.990 158.475 56.160 158.595 ;
        RECT 54.530 158.305 56.160 158.475 ;
        RECT 54.110 157.845 56.160 158.135 ;
        RECT 56.330 157.625 56.610 158.425 ;
        RECT 56.820 157.795 57.095 158.765 ;
        RECT 57.265 159.525 57.525 160.005 ;
        RECT 57.695 159.715 58.025 160.175 ;
        RECT 58.215 159.535 58.415 159.955 ;
        RECT 57.265 158.495 57.435 159.525 ;
        RECT 57.605 158.835 57.835 159.265 ;
        RECT 58.005 159.015 58.415 159.535 ;
        RECT 58.585 159.690 59.375 159.955 ;
        RECT 58.585 158.835 58.840 159.690 ;
        RECT 59.555 159.355 59.885 159.775 ;
        RECT 60.055 159.355 60.315 160.175 ;
        RECT 60.505 159.485 60.745 160.005 ;
        RECT 60.915 159.680 61.310 160.175 ;
        RECT 61.875 159.845 62.045 159.990 ;
        RECT 61.670 159.650 62.045 159.845 ;
        RECT 59.555 159.265 59.805 159.355 ;
        RECT 59.010 159.015 59.805 159.265 ;
        RECT 57.605 158.665 59.395 158.835 ;
        RECT 57.265 157.795 57.540 158.495 ;
        RECT 57.710 158.370 58.425 158.665 ;
        RECT 58.645 158.305 58.975 158.495 ;
        RECT 57.750 157.625 57.965 158.170 ;
        RECT 58.135 157.795 58.610 158.135 ;
        RECT 58.780 158.130 58.975 158.305 ;
        RECT 59.145 158.300 59.395 158.665 ;
        RECT 58.780 157.625 59.395 158.130 ;
        RECT 59.635 157.795 59.805 159.015 ;
        RECT 59.975 158.305 60.315 159.185 ;
        RECT 60.505 158.815 60.680 159.485 ;
        RECT 61.670 159.315 61.840 159.650 ;
        RECT 62.325 159.605 62.565 159.980 ;
        RECT 62.735 159.670 63.070 160.175 ;
        RECT 62.325 159.455 62.545 159.605 ;
        RECT 60.855 158.955 61.840 159.315 ;
        RECT 62.010 159.125 62.545 159.455 ;
        RECT 60.855 158.935 62.140 158.955 ;
        RECT 60.505 158.680 60.715 158.815 ;
        RECT 61.280 158.785 62.140 158.935 ;
        RECT 60.055 157.625 60.315 158.135 ;
        RECT 60.505 157.895 60.810 158.680 ;
        RECT 60.985 158.305 61.680 158.615 ;
        RECT 60.990 157.625 61.675 158.095 ;
        RECT 61.855 157.840 62.140 158.785 ;
        RECT 62.310 158.475 62.545 159.125 ;
        RECT 62.715 158.645 63.015 159.495 ;
        RECT 63.705 159.450 63.995 160.175 ;
        RECT 64.170 159.435 64.425 160.005 ;
        RECT 64.595 159.775 64.925 160.175 ;
        RECT 65.350 159.640 65.880 160.005 ;
        RECT 66.070 159.835 66.345 160.005 ;
        RECT 66.065 159.665 66.345 159.835 ;
        RECT 65.350 159.605 65.525 159.640 ;
        RECT 64.595 159.435 65.525 159.605 ;
        RECT 62.310 158.245 62.985 158.475 ;
        RECT 62.315 157.625 62.645 158.075 ;
        RECT 62.815 157.815 62.985 158.245 ;
        RECT 63.705 157.625 63.995 158.790 ;
        RECT 64.170 158.765 64.340 159.435 ;
        RECT 64.595 159.265 64.765 159.435 ;
        RECT 64.510 158.935 64.765 159.265 ;
        RECT 64.990 158.935 65.185 159.265 ;
        RECT 64.170 157.795 64.505 158.765 ;
        RECT 64.675 157.625 64.845 158.765 ;
        RECT 65.015 157.965 65.185 158.935 ;
        RECT 65.355 158.305 65.525 159.435 ;
        RECT 65.695 158.645 65.865 159.445 ;
        RECT 66.070 158.845 66.345 159.665 ;
        RECT 66.515 158.645 66.705 160.005 ;
        RECT 66.885 159.640 67.395 160.175 ;
        RECT 67.615 159.365 67.860 159.970 ;
        RECT 68.310 159.435 68.565 160.005 ;
        RECT 68.735 159.775 69.065 160.175 ;
        RECT 69.490 159.640 70.020 160.005 ;
        RECT 70.210 159.835 70.485 160.005 ;
        RECT 70.205 159.665 70.485 159.835 ;
        RECT 69.490 159.605 69.665 159.640 ;
        RECT 68.735 159.435 69.665 159.605 ;
        RECT 66.905 159.195 68.135 159.365 ;
        RECT 65.695 158.475 66.705 158.645 ;
        RECT 66.875 158.630 67.625 158.820 ;
        RECT 65.355 158.135 66.480 158.305 ;
        RECT 66.875 157.965 67.045 158.630 ;
        RECT 67.795 158.385 68.135 159.195 ;
        RECT 65.015 157.795 67.045 157.965 ;
        RECT 67.215 157.625 67.385 158.385 ;
        RECT 67.620 157.975 68.135 158.385 ;
        RECT 68.310 158.765 68.480 159.435 ;
        RECT 68.735 159.265 68.905 159.435 ;
        RECT 68.650 158.935 68.905 159.265 ;
        RECT 69.130 158.935 69.325 159.265 ;
        RECT 68.310 157.795 68.645 158.765 ;
        RECT 68.815 157.625 68.985 158.765 ;
        RECT 69.155 157.965 69.325 158.935 ;
        RECT 69.495 158.305 69.665 159.435 ;
        RECT 69.835 158.645 70.005 159.445 ;
        RECT 70.210 158.845 70.485 159.665 ;
        RECT 70.655 158.645 70.845 160.005 ;
        RECT 71.025 159.640 71.535 160.175 ;
        RECT 71.755 159.365 72.000 159.970 ;
        RECT 72.445 159.435 72.830 160.005 ;
        RECT 73.000 159.715 73.325 160.175 ;
        RECT 73.845 159.545 74.125 160.005 ;
        RECT 71.045 159.195 72.275 159.365 ;
        RECT 69.835 158.475 70.845 158.645 ;
        RECT 71.015 158.630 71.765 158.820 ;
        RECT 69.495 158.135 70.620 158.305 ;
        RECT 71.015 157.965 71.185 158.630 ;
        RECT 71.935 158.385 72.275 159.195 ;
        RECT 69.155 157.795 71.185 157.965 ;
        RECT 71.355 157.625 71.525 158.385 ;
        RECT 71.760 157.975 72.275 158.385 ;
        RECT 72.445 158.765 72.725 159.435 ;
        RECT 73.000 159.375 74.125 159.545 ;
        RECT 73.000 159.265 73.450 159.375 ;
        RECT 72.895 158.935 73.450 159.265 ;
        RECT 74.315 159.205 74.715 160.005 ;
        RECT 75.115 159.715 75.385 160.175 ;
        RECT 75.555 159.545 75.840 160.005 ;
        RECT 72.445 157.795 72.830 158.765 ;
        RECT 73.000 158.475 73.450 158.935 ;
        RECT 73.620 158.645 74.715 159.205 ;
        RECT 73.000 158.255 74.125 158.475 ;
        RECT 73.000 157.625 73.325 158.085 ;
        RECT 73.845 157.795 74.125 158.255 ;
        RECT 74.315 157.795 74.715 158.645 ;
        RECT 74.885 159.375 75.840 159.545 ;
        RECT 76.125 159.375 76.465 160.005 ;
        RECT 76.635 159.375 76.885 160.175 ;
        RECT 77.075 159.525 77.405 160.005 ;
        RECT 77.575 159.715 77.800 160.175 ;
        RECT 77.970 159.525 78.300 160.005 ;
        RECT 74.885 158.475 75.095 159.375 ;
        RECT 76.125 159.325 76.355 159.375 ;
        RECT 77.075 159.355 78.300 159.525 ;
        RECT 78.930 159.395 79.430 160.005 ;
        RECT 79.805 159.500 80.065 160.005 ;
        RECT 80.245 159.795 80.575 160.175 ;
        RECT 80.755 159.625 80.925 160.005 ;
        RECT 75.265 158.645 75.955 159.205 ;
        RECT 76.125 158.765 76.300 159.325 ;
        RECT 76.470 159.015 77.165 159.185 ;
        RECT 76.995 158.765 77.165 159.015 ;
        RECT 77.340 158.985 77.760 159.185 ;
        RECT 77.930 158.985 78.260 159.185 ;
        RECT 78.430 158.985 78.760 159.185 ;
        RECT 78.930 158.765 79.100 159.395 ;
        RECT 79.285 158.935 79.635 159.185 ;
        RECT 74.885 158.255 75.840 158.475 ;
        RECT 75.115 157.625 75.385 158.085 ;
        RECT 75.555 157.795 75.840 158.255 ;
        RECT 76.125 157.795 76.465 158.765 ;
        RECT 76.635 157.625 76.805 158.765 ;
        RECT 76.995 158.595 79.430 158.765 ;
        RECT 77.075 157.625 77.325 158.425 ;
        RECT 77.970 157.795 78.300 158.595 ;
        RECT 78.600 157.625 78.930 158.425 ;
        RECT 79.100 157.795 79.430 158.595 ;
        RECT 79.805 158.700 79.975 159.500 ;
        RECT 80.260 159.455 80.925 159.625 ;
        RECT 81.275 159.625 81.445 159.915 ;
        RECT 81.615 159.795 81.945 160.175 ;
        RECT 81.275 159.455 81.940 159.625 ;
        RECT 80.260 159.200 80.430 159.455 ;
        RECT 80.145 158.870 80.430 159.200 ;
        RECT 80.665 158.905 80.995 159.275 ;
        RECT 80.260 158.725 80.430 158.870 ;
        RECT 79.805 157.795 80.075 158.700 ;
        RECT 80.260 158.555 80.925 158.725 ;
        RECT 81.190 158.635 81.540 159.285 ;
        RECT 80.245 157.625 80.575 158.385 ;
        RECT 80.755 157.795 80.925 158.555 ;
        RECT 81.710 158.465 81.940 159.455 ;
        RECT 81.275 158.295 81.940 158.465 ;
        RECT 81.275 157.795 81.445 158.295 ;
        RECT 81.615 157.625 81.945 158.125 ;
        RECT 82.115 157.795 82.300 159.915 ;
        RECT 82.555 159.715 82.805 160.175 ;
        RECT 82.975 159.725 83.310 159.895 ;
        RECT 83.505 159.725 84.180 159.895 ;
        RECT 82.975 159.585 83.145 159.725 ;
        RECT 82.470 158.595 82.750 159.545 ;
        RECT 82.920 159.455 83.145 159.585 ;
        RECT 82.920 158.350 83.090 159.455 ;
        RECT 83.315 159.305 83.840 159.525 ;
        RECT 83.260 158.540 83.500 159.135 ;
        RECT 83.670 158.605 83.840 159.305 ;
        RECT 84.010 158.945 84.180 159.725 ;
        RECT 84.500 159.675 84.870 160.175 ;
        RECT 85.050 159.725 85.455 159.895 ;
        RECT 85.625 159.725 86.410 159.895 ;
        RECT 85.050 159.495 85.220 159.725 ;
        RECT 84.390 159.195 85.220 159.495 ;
        RECT 85.605 159.225 86.070 159.555 ;
        RECT 84.390 159.165 84.590 159.195 ;
        RECT 84.710 158.945 84.880 159.015 ;
        RECT 84.010 158.775 84.880 158.945 ;
        RECT 84.370 158.685 84.880 158.775 ;
        RECT 82.920 158.220 83.225 158.350 ;
        RECT 83.670 158.240 84.200 158.605 ;
        RECT 82.540 157.625 82.805 158.085 ;
        RECT 82.975 157.795 83.225 158.220 ;
        RECT 84.370 158.070 84.540 158.685 ;
        RECT 83.435 157.900 84.540 158.070 ;
        RECT 84.710 157.625 84.880 158.425 ;
        RECT 85.050 158.125 85.220 159.195 ;
        RECT 85.390 158.295 85.580 159.015 ;
        RECT 85.750 158.265 86.070 159.225 ;
        RECT 86.240 159.265 86.410 159.725 ;
        RECT 86.685 159.645 86.895 160.175 ;
        RECT 87.155 159.435 87.485 159.960 ;
        RECT 87.655 159.565 87.825 160.175 ;
        RECT 87.995 159.520 88.325 159.955 ;
        RECT 87.995 159.435 88.375 159.520 ;
        RECT 87.285 159.265 87.485 159.435 ;
        RECT 88.150 159.395 88.375 159.435 ;
        RECT 88.545 159.425 89.755 160.175 ;
        RECT 86.240 158.935 87.115 159.265 ;
        RECT 87.285 158.935 88.035 159.265 ;
        RECT 85.050 157.795 85.300 158.125 ;
        RECT 86.240 158.095 86.410 158.935 ;
        RECT 87.285 158.730 87.475 158.935 ;
        RECT 88.205 158.815 88.375 159.395 ;
        RECT 88.160 158.765 88.375 158.815 ;
        RECT 86.580 158.355 87.475 158.730 ;
        RECT 87.985 158.685 88.375 158.765 ;
        RECT 88.545 158.715 89.065 159.255 ;
        RECT 89.235 158.885 89.755 159.425 ;
        RECT 100.140 159.370 100.810 161.630 ;
        RECT 101.480 161.060 105.520 161.230 ;
        RECT 101.140 160.000 101.310 161.000 ;
        RECT 105.690 160.000 105.860 161.000 ;
        RECT 101.480 159.770 105.520 159.940 ;
        RECT 106.200 159.370 106.370 161.630 ;
        RECT 100.140 159.200 106.370 159.370 ;
        RECT 85.525 157.925 86.410 158.095 ;
        RECT 86.590 157.625 86.905 158.125 ;
        RECT 87.135 157.795 87.475 158.355 ;
        RECT 87.645 157.625 87.815 158.635 ;
        RECT 87.985 157.840 88.315 158.685 ;
        RECT 88.545 157.625 89.755 158.715 ;
        RECT 12.100 157.455 89.840 157.625 ;
        RECT 12.185 156.365 13.395 157.455 ;
        RECT 13.565 157.020 18.910 157.455 ;
        RECT 19.085 157.020 24.430 157.455 ;
        RECT 12.185 155.655 12.705 156.195 ;
        RECT 12.875 155.825 13.395 156.365 ;
        RECT 12.185 154.905 13.395 155.655 ;
        RECT 15.150 155.450 15.490 156.280 ;
        RECT 16.970 155.770 17.320 157.020 ;
        RECT 20.670 155.450 21.010 156.280 ;
        RECT 22.490 155.770 22.840 157.020 ;
        RECT 25.065 156.290 25.355 157.455 ;
        RECT 25.525 157.020 30.870 157.455 ;
        RECT 13.565 154.905 18.910 155.450 ;
        RECT 19.085 154.905 24.430 155.450 ;
        RECT 25.065 154.905 25.355 155.630 ;
        RECT 27.110 155.450 27.450 156.280 ;
        RECT 28.930 155.770 29.280 157.020 ;
        RECT 31.045 156.365 34.555 157.455 ;
        RECT 31.045 155.675 32.695 156.195 ;
        RECT 32.865 155.845 34.555 156.365 ;
        RECT 35.190 156.315 35.465 157.285 ;
        RECT 35.675 156.655 35.955 157.455 ;
        RECT 36.125 156.945 37.315 157.235 ;
        RECT 36.125 156.605 37.295 156.775 ;
        RECT 36.125 156.485 36.295 156.605 ;
        RECT 35.635 156.315 36.295 156.485 ;
        RECT 25.525 154.905 30.870 155.450 ;
        RECT 31.045 154.905 34.555 155.675 ;
        RECT 35.190 155.580 35.360 156.315 ;
        RECT 35.635 156.145 35.805 156.315 ;
        RECT 36.605 156.145 36.800 156.435 ;
        RECT 36.970 156.315 37.295 156.605 ;
        RECT 37.670 156.485 38.060 156.660 ;
        RECT 38.545 156.655 38.875 157.455 ;
        RECT 39.045 156.665 39.580 157.285 ;
        RECT 37.670 156.315 39.095 156.485 ;
        RECT 35.530 155.815 35.805 156.145 ;
        RECT 35.975 155.815 36.800 156.145 ;
        RECT 36.970 155.815 37.315 156.145 ;
        RECT 35.635 155.645 35.805 155.815 ;
        RECT 35.190 155.235 35.465 155.580 ;
        RECT 35.635 155.475 37.300 155.645 ;
        RECT 37.545 155.585 37.900 156.145 ;
        RECT 35.655 154.905 36.035 155.305 ;
        RECT 36.205 155.125 36.375 155.475 ;
        RECT 36.545 154.905 36.875 155.305 ;
        RECT 37.045 155.125 37.300 155.475 ;
        RECT 38.070 155.415 38.240 156.315 ;
        RECT 38.410 155.585 38.675 156.145 ;
        RECT 38.925 155.815 39.095 156.315 ;
        RECT 39.265 155.645 39.580 156.665 ;
        RECT 37.650 154.905 37.890 155.415 ;
        RECT 38.070 155.085 38.350 155.415 ;
        RECT 38.580 154.905 38.795 155.415 ;
        RECT 38.965 155.075 39.580 155.645 ;
        RECT 39.785 156.315 40.060 157.285 ;
        RECT 40.270 156.655 40.550 157.455 ;
        RECT 40.720 156.945 42.335 157.275 ;
        RECT 40.720 156.605 41.895 156.775 ;
        RECT 40.720 156.485 40.890 156.605 ;
        RECT 40.230 156.315 40.890 156.485 ;
        RECT 39.785 155.580 39.955 156.315 ;
        RECT 40.230 156.145 40.400 156.315 ;
        RECT 41.150 156.145 41.395 156.435 ;
        RECT 41.565 156.315 41.895 156.605 ;
        RECT 42.155 156.145 42.325 156.705 ;
        RECT 42.575 156.315 42.835 157.455 ;
        RECT 43.005 156.315 43.390 157.285 ;
        RECT 43.560 156.995 43.885 157.455 ;
        RECT 44.405 156.825 44.685 157.285 ;
        RECT 43.560 156.605 44.685 156.825 ;
        RECT 40.125 155.815 40.400 156.145 ;
        RECT 40.570 155.815 41.395 156.145 ;
        RECT 41.610 155.815 42.325 156.145 ;
        RECT 42.495 155.895 42.830 156.145 ;
        RECT 40.230 155.645 40.400 155.815 ;
        RECT 42.075 155.725 42.325 155.815 ;
        RECT 39.785 155.235 40.060 155.580 ;
        RECT 40.230 155.475 41.895 155.645 ;
        RECT 40.250 154.905 40.625 155.305 ;
        RECT 40.795 155.125 40.965 155.475 ;
        RECT 41.135 154.905 41.465 155.305 ;
        RECT 41.635 155.075 41.895 155.475 ;
        RECT 42.075 155.305 42.405 155.725 ;
        RECT 42.575 154.905 42.835 155.725 ;
        RECT 43.005 155.645 43.285 156.315 ;
        RECT 43.560 156.145 44.010 156.605 ;
        RECT 44.875 156.435 45.275 157.285 ;
        RECT 45.675 156.995 45.945 157.455 ;
        RECT 46.115 156.825 46.400 157.285 ;
        RECT 43.455 155.815 44.010 156.145 ;
        RECT 44.180 155.875 45.275 156.435 ;
        RECT 43.560 155.705 44.010 155.815 ;
        RECT 43.005 155.075 43.390 155.645 ;
        RECT 43.560 155.535 44.685 155.705 ;
        RECT 43.560 154.905 43.885 155.365 ;
        RECT 44.405 155.075 44.685 155.535 ;
        RECT 44.875 155.075 45.275 155.875 ;
        RECT 45.445 156.605 46.400 156.825 ;
        RECT 46.800 156.825 47.085 157.285 ;
        RECT 47.255 156.995 47.525 157.455 ;
        RECT 46.800 156.605 47.755 156.825 ;
        RECT 45.445 155.705 45.655 156.605 ;
        RECT 45.825 155.875 46.515 156.435 ;
        RECT 46.685 155.875 47.375 156.435 ;
        RECT 47.545 155.705 47.755 156.605 ;
        RECT 45.445 155.535 46.400 155.705 ;
        RECT 45.675 154.905 45.945 155.365 ;
        RECT 46.115 155.075 46.400 155.535 ;
        RECT 46.800 155.535 47.755 155.705 ;
        RECT 47.925 156.435 48.325 157.285 ;
        RECT 48.515 156.825 48.795 157.285 ;
        RECT 49.315 156.995 49.640 157.455 ;
        RECT 48.515 156.605 49.640 156.825 ;
        RECT 47.925 155.875 49.020 156.435 ;
        RECT 49.190 156.145 49.640 156.605 ;
        RECT 49.810 156.315 50.195 157.285 ;
        RECT 46.800 155.075 47.085 155.535 ;
        RECT 47.255 154.905 47.525 155.365 ;
        RECT 47.925 155.075 48.325 155.875 ;
        RECT 49.190 155.815 49.745 156.145 ;
        RECT 49.190 155.705 49.640 155.815 ;
        RECT 48.515 155.535 49.640 155.705 ;
        RECT 49.915 155.645 50.195 156.315 ;
        RECT 50.825 156.290 51.115 157.455 ;
        RECT 51.285 156.315 51.545 157.455 ;
        RECT 51.715 156.305 52.045 157.285 ;
        RECT 52.215 156.315 52.495 157.455 ;
        RECT 52.665 156.315 53.005 157.285 ;
        RECT 53.175 156.315 53.345 157.455 ;
        RECT 53.615 156.655 53.865 157.455 ;
        RECT 54.510 156.485 54.840 157.285 ;
        RECT 55.140 156.655 55.470 157.455 ;
        RECT 55.640 156.485 55.970 157.285 ;
        RECT 53.535 156.315 55.970 156.485 ;
        RECT 56.345 156.585 56.620 157.285 ;
        RECT 56.830 156.910 57.045 157.455 ;
        RECT 57.215 156.945 57.690 157.285 ;
        RECT 57.860 156.950 58.475 157.455 ;
        RECT 57.860 156.775 58.055 156.950 ;
        RECT 51.305 155.895 51.640 156.145 ;
        RECT 51.810 155.705 51.980 156.305 ;
        RECT 52.150 155.875 52.485 156.145 ;
        RECT 52.665 155.705 52.840 156.315 ;
        RECT 53.535 156.065 53.705 156.315 ;
        RECT 53.010 155.895 53.705 156.065 ;
        RECT 53.880 155.895 54.300 156.095 ;
        RECT 54.470 155.895 54.800 156.095 ;
        RECT 54.970 155.895 55.300 156.095 ;
        RECT 48.515 155.075 48.795 155.535 ;
        RECT 49.315 154.905 49.640 155.365 ;
        RECT 49.810 155.075 50.195 155.645 ;
        RECT 50.825 154.905 51.115 155.630 ;
        RECT 51.285 155.075 51.980 155.705 ;
        RECT 52.185 154.905 52.495 155.705 ;
        RECT 52.665 155.075 53.005 155.705 ;
        RECT 53.175 154.905 53.425 155.705 ;
        RECT 53.615 155.555 54.840 155.725 ;
        RECT 53.615 155.075 53.945 155.555 ;
        RECT 54.115 154.905 54.340 155.365 ;
        RECT 54.510 155.075 54.840 155.555 ;
        RECT 55.470 155.685 55.640 156.315 ;
        RECT 55.825 155.895 56.175 156.145 ;
        RECT 55.470 155.075 55.970 155.685 ;
        RECT 56.345 155.555 56.515 156.585 ;
        RECT 56.790 156.415 57.505 156.710 ;
        RECT 57.725 156.585 58.055 156.775 ;
        RECT 58.225 156.415 58.475 156.780 ;
        RECT 56.685 156.245 58.475 156.415 ;
        RECT 56.685 155.815 56.915 156.245 ;
        RECT 56.345 155.075 56.605 155.555 ;
        RECT 57.085 155.545 57.495 156.065 ;
        RECT 56.775 154.905 57.105 155.365 ;
        RECT 57.295 155.125 57.495 155.545 ;
        RECT 57.665 155.390 57.920 156.245 ;
        RECT 58.715 156.065 58.885 157.285 ;
        RECT 59.135 156.945 59.395 157.455 ;
        RECT 58.090 155.815 58.885 156.065 ;
        RECT 59.055 155.895 59.395 156.775 ;
        RECT 59.585 156.400 59.890 157.185 ;
        RECT 60.070 156.985 60.755 157.455 ;
        RECT 60.065 156.465 60.760 156.775 ;
        RECT 58.635 155.725 58.885 155.815 ;
        RECT 57.665 155.125 58.455 155.390 ;
        RECT 58.635 155.305 58.965 155.725 ;
        RECT 59.135 154.905 59.395 155.725 ;
        RECT 59.585 155.595 59.760 156.400 ;
        RECT 60.935 156.295 61.220 157.240 ;
        RECT 61.395 157.005 61.725 157.455 ;
        RECT 61.895 156.835 62.065 157.265 ;
        RECT 60.360 156.145 61.220 156.295 ;
        RECT 59.935 156.125 61.220 156.145 ;
        RECT 61.390 156.605 62.065 156.835 ;
        RECT 59.935 155.765 60.920 156.125 ;
        RECT 61.390 155.955 61.625 156.605 ;
        RECT 62.330 156.505 62.595 157.275 ;
        RECT 62.765 156.735 63.095 157.455 ;
        RECT 63.285 156.915 63.545 157.275 ;
        RECT 63.715 157.085 64.045 157.455 ;
        RECT 64.215 156.915 64.475 157.275 ;
        RECT 63.285 156.685 64.475 156.915 ;
        RECT 65.045 156.505 65.335 157.275 ;
        RECT 59.585 155.075 59.825 155.595 ;
        RECT 60.750 155.430 60.920 155.765 ;
        RECT 61.090 155.625 61.625 155.955 ;
        RECT 61.405 155.475 61.625 155.625 ;
        RECT 61.795 155.585 62.095 156.435 ;
        RECT 59.995 154.905 60.390 155.400 ;
        RECT 60.750 155.235 61.125 155.430 ;
        RECT 60.955 155.090 61.125 155.235 ;
        RECT 61.405 155.100 61.645 155.475 ;
        RECT 61.815 154.905 62.150 155.410 ;
        RECT 62.330 155.085 62.665 156.505 ;
        RECT 62.840 156.325 65.335 156.505 ;
        RECT 62.840 155.635 63.065 156.325 ;
        RECT 65.550 156.315 65.885 157.285 ;
        RECT 66.055 156.315 66.225 157.455 ;
        RECT 66.395 157.115 68.425 157.285 ;
        RECT 63.265 155.815 63.545 156.145 ;
        RECT 63.725 155.815 64.300 156.145 ;
        RECT 64.480 155.815 64.915 156.145 ;
        RECT 65.095 155.815 65.365 156.145 ;
        RECT 65.550 155.645 65.720 156.315 ;
        RECT 66.395 156.145 66.565 157.115 ;
        RECT 65.890 155.815 66.145 156.145 ;
        RECT 66.370 155.815 66.565 156.145 ;
        RECT 66.735 156.775 67.860 156.945 ;
        RECT 65.975 155.645 66.145 155.815 ;
        RECT 66.735 155.645 66.905 156.775 ;
        RECT 62.840 155.445 65.325 155.635 ;
        RECT 62.845 154.905 63.590 155.275 ;
        RECT 64.155 155.085 64.410 155.445 ;
        RECT 64.590 154.905 64.920 155.275 ;
        RECT 65.100 155.085 65.325 155.445 ;
        RECT 65.550 155.075 65.805 155.645 ;
        RECT 65.975 155.475 66.905 155.645 ;
        RECT 67.075 156.435 68.085 156.605 ;
        RECT 67.075 155.635 67.245 156.435 ;
        RECT 67.450 156.095 67.725 156.235 ;
        RECT 67.445 155.925 67.725 156.095 ;
        RECT 66.730 155.440 66.905 155.475 ;
        RECT 65.975 154.905 66.305 155.305 ;
        RECT 66.730 155.075 67.260 155.440 ;
        RECT 67.450 155.075 67.725 155.925 ;
        RECT 67.895 155.075 68.085 156.435 ;
        RECT 68.255 156.450 68.425 157.115 ;
        RECT 68.595 156.695 68.765 157.455 ;
        RECT 69.000 156.695 69.515 157.105 ;
        RECT 68.255 156.260 69.005 156.450 ;
        RECT 69.175 155.885 69.515 156.695 ;
        RECT 68.285 155.715 69.515 155.885 ;
        RECT 69.690 156.315 70.025 157.285 ;
        RECT 70.195 156.315 70.365 157.455 ;
        RECT 70.535 157.115 72.565 157.285 ;
        RECT 68.265 154.905 68.775 155.440 ;
        RECT 68.995 155.110 69.240 155.715 ;
        RECT 69.690 155.645 69.860 156.315 ;
        RECT 70.535 156.145 70.705 157.115 ;
        RECT 70.030 155.815 70.285 156.145 ;
        RECT 70.510 155.815 70.705 156.145 ;
        RECT 70.875 156.775 72.000 156.945 ;
        RECT 70.115 155.645 70.285 155.815 ;
        RECT 70.875 155.645 71.045 156.775 ;
        RECT 69.690 155.075 69.945 155.645 ;
        RECT 70.115 155.475 71.045 155.645 ;
        RECT 71.215 156.435 72.225 156.605 ;
        RECT 71.215 155.635 71.385 156.435 ;
        RECT 71.590 156.095 71.865 156.235 ;
        RECT 71.585 155.925 71.865 156.095 ;
        RECT 70.870 155.440 71.045 155.475 ;
        RECT 70.115 154.905 70.445 155.305 ;
        RECT 70.870 155.075 71.400 155.440 ;
        RECT 71.590 155.075 71.865 155.925 ;
        RECT 72.035 155.075 72.225 156.435 ;
        RECT 72.395 156.450 72.565 157.115 ;
        RECT 72.735 156.695 72.905 157.455 ;
        RECT 73.140 156.695 73.655 157.105 ;
        RECT 72.395 156.260 73.145 156.450 ;
        RECT 73.315 155.885 73.655 156.695 ;
        RECT 74.470 156.485 74.860 156.660 ;
        RECT 75.345 156.655 75.675 157.455 ;
        RECT 75.845 156.665 76.380 157.285 ;
        RECT 74.470 156.315 75.895 156.485 ;
        RECT 72.425 155.715 73.655 155.885 ;
        RECT 72.405 154.905 72.915 155.440 ;
        RECT 73.135 155.110 73.380 155.715 ;
        RECT 74.345 155.585 74.700 156.145 ;
        RECT 74.870 155.415 75.040 156.315 ;
        RECT 75.210 155.585 75.475 156.145 ;
        RECT 75.725 155.815 75.895 156.315 ;
        RECT 76.065 155.645 76.380 156.665 ;
        RECT 76.585 156.290 76.875 157.455 ;
        RECT 77.045 156.315 77.430 157.285 ;
        RECT 77.600 156.995 77.925 157.455 ;
        RECT 78.445 156.825 78.725 157.285 ;
        RECT 77.600 156.605 78.725 156.825 ;
        RECT 74.450 154.905 74.690 155.415 ;
        RECT 74.870 155.085 75.150 155.415 ;
        RECT 75.380 154.905 75.595 155.415 ;
        RECT 75.765 155.075 76.380 155.645 ;
        RECT 77.045 155.645 77.325 156.315 ;
        RECT 77.600 156.145 78.050 156.605 ;
        RECT 78.915 156.435 79.315 157.285 ;
        RECT 79.715 156.995 79.985 157.455 ;
        RECT 80.155 156.825 80.440 157.285 ;
        RECT 77.495 155.815 78.050 156.145 ;
        RECT 78.220 155.875 79.315 156.435 ;
        RECT 77.600 155.705 78.050 155.815 ;
        RECT 76.585 154.905 76.875 155.630 ;
        RECT 77.045 155.075 77.430 155.645 ;
        RECT 77.600 155.535 78.725 155.705 ;
        RECT 77.600 154.905 77.925 155.365 ;
        RECT 78.445 155.075 78.725 155.535 ;
        RECT 78.915 155.075 79.315 155.875 ;
        RECT 79.485 156.605 80.440 156.825 ;
        RECT 79.485 155.705 79.695 156.605 ;
        RECT 79.865 155.875 80.555 156.435 ;
        RECT 80.725 156.315 81.065 157.285 ;
        RECT 81.235 156.315 81.405 157.455 ;
        RECT 81.675 156.655 81.925 157.455 ;
        RECT 82.570 156.485 82.900 157.285 ;
        RECT 83.200 156.655 83.530 157.455 ;
        RECT 83.700 156.485 84.030 157.285 ;
        RECT 81.595 156.315 84.030 156.485 ;
        RECT 84.405 156.315 84.745 157.285 ;
        RECT 84.915 156.315 85.085 157.455 ;
        RECT 85.355 156.655 85.605 157.455 ;
        RECT 86.250 156.485 86.580 157.285 ;
        RECT 86.880 156.655 87.210 157.455 ;
        RECT 87.380 156.485 87.710 157.285 ;
        RECT 85.275 156.315 87.710 156.485 ;
        RECT 88.545 156.365 89.755 157.455 ;
        RECT 80.725 155.705 80.900 156.315 ;
        RECT 81.595 156.065 81.765 156.315 ;
        RECT 81.070 155.895 81.765 156.065 ;
        RECT 81.940 155.895 82.360 156.095 ;
        RECT 82.530 155.895 82.860 156.095 ;
        RECT 83.030 155.895 83.360 156.095 ;
        RECT 79.485 155.535 80.440 155.705 ;
        RECT 79.715 154.905 79.985 155.365 ;
        RECT 80.155 155.075 80.440 155.535 ;
        RECT 80.725 155.075 81.065 155.705 ;
        RECT 81.235 154.905 81.485 155.705 ;
        RECT 81.675 155.555 82.900 155.725 ;
        RECT 81.675 155.075 82.005 155.555 ;
        RECT 82.175 154.905 82.400 155.365 ;
        RECT 82.570 155.075 82.900 155.555 ;
        RECT 83.530 155.685 83.700 156.315 ;
        RECT 83.885 155.895 84.235 156.145 ;
        RECT 84.405 155.705 84.580 156.315 ;
        RECT 85.275 156.065 85.445 156.315 ;
        RECT 84.750 155.895 85.445 156.065 ;
        RECT 85.620 155.895 86.040 156.095 ;
        RECT 86.210 155.895 86.540 156.095 ;
        RECT 86.710 155.895 87.040 156.095 ;
        RECT 83.530 155.075 84.030 155.685 ;
        RECT 84.405 155.075 84.745 155.705 ;
        RECT 84.915 154.905 85.165 155.705 ;
        RECT 85.355 155.555 86.580 155.725 ;
        RECT 85.355 155.075 85.685 155.555 ;
        RECT 85.855 154.905 86.080 155.365 ;
        RECT 86.250 155.075 86.580 155.555 ;
        RECT 87.210 155.685 87.380 156.315 ;
        RECT 87.565 155.895 87.915 156.145 ;
        RECT 88.545 155.825 89.065 156.365 ;
        RECT 87.210 155.075 87.710 155.685 ;
        RECT 89.235 155.655 89.755 156.195 ;
        RECT 88.545 154.905 89.755 155.655 ;
        RECT 100.140 155.940 100.810 159.200 ;
        RECT 101.480 158.630 105.520 158.800 ;
        RECT 101.140 156.570 101.310 158.570 ;
        RECT 105.690 156.570 105.860 158.570 ;
        RECT 101.480 156.340 105.520 156.510 ;
        RECT 106.200 155.940 106.370 159.200 ;
        RECT 100.140 155.770 106.370 155.940 ;
        RECT 12.100 154.735 89.840 154.905 ;
        RECT 12.185 153.985 13.395 154.735 ;
        RECT 13.565 154.190 18.910 154.735 ;
        RECT 19.085 154.190 24.430 154.735 ;
        RECT 24.605 154.190 29.950 154.735 ;
        RECT 30.125 154.190 35.470 154.735 ;
        RECT 12.185 153.445 12.705 153.985 ;
        RECT 12.875 153.275 13.395 153.815 ;
        RECT 15.150 153.360 15.490 154.190 ;
        RECT 12.185 152.185 13.395 153.275 ;
        RECT 16.970 152.620 17.320 153.870 ;
        RECT 20.670 153.360 21.010 154.190 ;
        RECT 22.490 152.620 22.840 153.870 ;
        RECT 26.190 153.360 26.530 154.190 ;
        RECT 28.010 152.620 28.360 153.870 ;
        RECT 31.710 153.360 32.050 154.190 ;
        RECT 35.645 153.965 37.315 154.735 ;
        RECT 37.945 154.010 38.235 154.735 ;
        RECT 39.335 154.010 39.665 154.520 ;
        RECT 39.835 154.335 40.165 154.735 ;
        RECT 41.215 154.165 41.545 154.505 ;
        RECT 41.715 154.335 42.045 154.735 ;
        RECT 33.530 152.620 33.880 153.870 ;
        RECT 35.645 153.445 36.395 153.965 ;
        RECT 36.565 153.275 37.315 153.795 ;
        RECT 13.565 152.185 18.910 152.620 ;
        RECT 19.085 152.185 24.430 152.620 ;
        RECT 24.605 152.185 29.950 152.620 ;
        RECT 30.125 152.185 35.470 152.620 ;
        RECT 35.645 152.185 37.315 153.275 ;
        RECT 37.945 152.185 38.235 153.350 ;
        RECT 39.335 153.245 39.525 154.010 ;
        RECT 39.835 153.995 42.200 154.165 ;
        RECT 43.055 154.080 43.385 154.515 ;
        RECT 43.555 154.125 43.725 154.735 ;
        RECT 39.835 153.825 40.005 153.995 ;
        RECT 39.695 153.495 40.005 153.825 ;
        RECT 40.175 153.495 40.480 153.825 ;
        RECT 39.335 152.395 39.665 153.245 ;
        RECT 39.835 152.185 40.085 153.325 ;
        RECT 40.265 153.165 40.480 153.495 ;
        RECT 40.655 153.165 40.940 153.825 ;
        RECT 41.135 153.165 41.400 153.825 ;
        RECT 41.615 153.165 41.860 153.825 ;
        RECT 42.030 152.995 42.200 153.995 ;
        RECT 43.005 153.995 43.385 154.080 ;
        RECT 43.895 153.995 44.225 154.520 ;
        RECT 44.485 154.205 44.695 154.735 ;
        RECT 44.970 154.285 45.755 154.455 ;
        RECT 45.925 154.285 46.330 154.455 ;
        RECT 43.005 153.955 43.230 153.995 ;
        RECT 43.005 153.375 43.175 153.955 ;
        RECT 43.895 153.825 44.095 153.995 ;
        RECT 44.970 153.825 45.140 154.285 ;
        RECT 43.345 153.495 44.095 153.825 ;
        RECT 44.265 153.495 45.140 153.825 ;
        RECT 43.005 153.325 43.220 153.375 ;
        RECT 43.005 153.245 43.395 153.325 ;
        RECT 40.275 152.825 41.565 152.995 ;
        RECT 40.275 152.405 40.525 152.825 ;
        RECT 40.755 152.185 41.085 152.655 ;
        RECT 41.315 152.405 41.565 152.825 ;
        RECT 41.745 152.825 42.200 152.995 ;
        RECT 41.745 152.395 42.075 152.825 ;
        RECT 43.065 152.400 43.395 153.245 ;
        RECT 43.905 153.290 44.095 153.495 ;
        RECT 43.565 152.185 43.735 153.195 ;
        RECT 43.905 152.915 44.800 153.290 ;
        RECT 43.905 152.355 44.245 152.915 ;
        RECT 44.475 152.185 44.790 152.685 ;
        RECT 44.970 152.655 45.140 153.495 ;
        RECT 45.310 153.785 45.775 154.115 ;
        RECT 46.160 154.055 46.330 154.285 ;
        RECT 46.510 154.235 46.880 154.735 ;
        RECT 47.200 154.285 47.875 154.455 ;
        RECT 48.070 154.285 48.405 154.455 ;
        RECT 45.310 152.825 45.630 153.785 ;
        RECT 46.160 153.755 46.990 154.055 ;
        RECT 45.800 152.855 45.990 153.575 ;
        RECT 46.160 152.685 46.330 153.755 ;
        RECT 46.790 153.725 46.990 153.755 ;
        RECT 46.500 153.505 46.670 153.575 ;
        RECT 47.200 153.505 47.370 154.285 ;
        RECT 48.235 154.145 48.405 154.285 ;
        RECT 48.575 154.275 48.825 154.735 ;
        RECT 46.500 153.335 47.370 153.505 ;
        RECT 47.540 153.865 48.065 154.085 ;
        RECT 48.235 154.015 48.460 154.145 ;
        RECT 46.500 153.245 47.010 153.335 ;
        RECT 44.970 152.485 45.855 152.655 ;
        RECT 46.080 152.355 46.330 152.685 ;
        RECT 46.500 152.185 46.670 152.985 ;
        RECT 46.840 152.630 47.010 153.245 ;
        RECT 47.540 153.165 47.710 153.865 ;
        RECT 47.180 152.800 47.710 153.165 ;
        RECT 47.880 153.100 48.120 153.695 ;
        RECT 48.290 152.910 48.460 154.015 ;
        RECT 48.630 153.155 48.910 154.105 ;
        RECT 48.155 152.780 48.460 152.910 ;
        RECT 46.840 152.460 47.945 152.630 ;
        RECT 48.155 152.355 48.405 152.780 ;
        RECT 48.575 152.185 48.840 152.645 ;
        RECT 49.080 152.355 49.265 154.475 ;
        RECT 49.435 154.355 49.765 154.735 ;
        RECT 49.935 154.185 50.105 154.475 ;
        RECT 49.440 154.015 50.105 154.185 ;
        RECT 49.440 153.025 49.670 154.015 ;
        RECT 49.840 153.195 50.190 153.845 ;
        RECT 49.440 152.855 50.105 153.025 ;
        RECT 49.435 152.185 49.765 152.685 ;
        RECT 49.935 152.355 50.105 152.855 ;
        RECT 50.375 152.365 50.635 154.555 ;
        RECT 50.895 154.365 51.565 154.735 ;
        RECT 51.745 154.185 52.055 154.555 ;
        RECT 50.825 153.985 52.055 154.185 ;
        RECT 50.825 153.315 51.115 153.985 ;
        RECT 52.235 153.805 52.465 154.445 ;
        RECT 52.645 154.005 52.935 154.735 ;
        RECT 54.135 154.185 54.305 154.475 ;
        RECT 54.475 154.355 54.805 154.735 ;
        RECT 54.135 154.015 54.800 154.185 ;
        RECT 51.295 153.495 51.760 153.805 ;
        RECT 51.940 153.495 52.465 153.805 ;
        RECT 52.645 153.495 52.945 153.825 ;
        RECT 50.825 153.095 51.595 153.315 ;
        RECT 50.805 152.185 51.145 152.915 ;
        RECT 51.325 152.365 51.595 153.095 ;
        RECT 51.775 153.075 52.935 153.315 ;
        RECT 54.050 153.195 54.400 153.845 ;
        RECT 51.775 152.365 52.005 153.075 ;
        RECT 52.175 152.185 52.505 152.895 ;
        RECT 52.675 152.365 52.935 153.075 ;
        RECT 54.570 153.025 54.800 154.015 ;
        RECT 54.135 152.855 54.800 153.025 ;
        RECT 54.135 152.355 54.305 152.855 ;
        RECT 54.475 152.185 54.805 152.685 ;
        RECT 54.975 152.355 55.160 154.475 ;
        RECT 55.415 154.275 55.665 154.735 ;
        RECT 55.835 154.285 56.170 154.455 ;
        RECT 56.365 154.285 57.040 154.455 ;
        RECT 55.835 154.145 56.005 154.285 ;
        RECT 55.330 153.155 55.610 154.105 ;
        RECT 55.780 154.015 56.005 154.145 ;
        RECT 55.780 152.910 55.950 154.015 ;
        RECT 56.175 153.865 56.700 154.085 ;
        RECT 56.120 153.100 56.360 153.695 ;
        RECT 56.530 153.165 56.700 153.865 ;
        RECT 56.870 153.505 57.040 154.285 ;
        RECT 57.360 154.235 57.730 154.735 ;
        RECT 57.910 154.285 58.315 154.455 ;
        RECT 58.485 154.285 59.270 154.455 ;
        RECT 57.910 154.055 58.080 154.285 ;
        RECT 57.250 153.755 58.080 154.055 ;
        RECT 58.465 153.785 58.930 154.115 ;
        RECT 57.250 153.725 57.450 153.755 ;
        RECT 57.570 153.505 57.740 153.575 ;
        RECT 56.870 153.335 57.740 153.505 ;
        RECT 57.230 153.245 57.740 153.335 ;
        RECT 55.780 152.780 56.085 152.910 ;
        RECT 56.530 152.800 57.060 153.165 ;
        RECT 55.400 152.185 55.665 152.645 ;
        RECT 55.835 152.355 56.085 152.780 ;
        RECT 57.230 152.630 57.400 153.245 ;
        RECT 56.295 152.460 57.400 152.630 ;
        RECT 57.570 152.185 57.740 152.985 ;
        RECT 57.910 152.685 58.080 153.755 ;
        RECT 58.250 152.855 58.440 153.575 ;
        RECT 58.610 152.825 58.930 153.785 ;
        RECT 59.100 153.825 59.270 154.285 ;
        RECT 59.545 154.205 59.755 154.735 ;
        RECT 60.015 153.995 60.345 154.520 ;
        RECT 60.515 154.125 60.685 154.735 ;
        RECT 60.855 154.080 61.185 154.515 ;
        RECT 61.405 154.085 61.665 154.565 ;
        RECT 61.835 154.195 62.085 154.735 ;
        RECT 60.855 153.995 61.235 154.080 ;
        RECT 60.145 153.825 60.345 153.995 ;
        RECT 61.010 153.955 61.235 153.995 ;
        RECT 59.100 153.495 59.975 153.825 ;
        RECT 60.145 153.495 60.895 153.825 ;
        RECT 57.910 152.355 58.160 152.685 ;
        RECT 59.100 152.655 59.270 153.495 ;
        RECT 60.145 153.290 60.335 153.495 ;
        RECT 61.065 153.375 61.235 153.955 ;
        RECT 61.020 153.325 61.235 153.375 ;
        RECT 59.440 152.915 60.335 153.290 ;
        RECT 60.845 153.245 61.235 153.325 ;
        RECT 58.385 152.485 59.270 152.655 ;
        RECT 59.450 152.185 59.765 152.685 ;
        RECT 59.995 152.355 60.335 152.915 ;
        RECT 60.505 152.185 60.675 153.195 ;
        RECT 60.845 152.400 61.175 153.245 ;
        RECT 61.405 153.055 61.575 154.085 ;
        RECT 62.255 154.030 62.475 154.515 ;
        RECT 61.745 153.435 61.975 153.830 ;
        RECT 62.145 153.605 62.475 154.030 ;
        RECT 62.645 154.355 63.535 154.525 ;
        RECT 62.645 153.630 62.815 154.355 ;
        RECT 62.985 153.800 63.535 154.185 ;
        RECT 63.705 154.010 63.995 154.735 ;
        RECT 64.165 153.995 64.550 154.565 ;
        RECT 64.720 154.275 65.045 154.735 ;
        RECT 65.565 154.105 65.845 154.565 ;
        RECT 62.645 153.560 63.535 153.630 ;
        RECT 62.640 153.535 63.535 153.560 ;
        RECT 62.630 153.520 63.535 153.535 ;
        RECT 62.625 153.505 63.535 153.520 ;
        RECT 62.615 153.500 63.535 153.505 ;
        RECT 62.610 153.490 63.535 153.500 ;
        RECT 62.605 153.480 63.535 153.490 ;
        RECT 62.595 153.475 63.535 153.480 ;
        RECT 62.585 153.465 63.535 153.475 ;
        RECT 62.575 153.460 63.535 153.465 ;
        RECT 62.575 153.455 62.910 153.460 ;
        RECT 62.560 153.450 62.910 153.455 ;
        RECT 62.545 153.440 62.910 153.450 ;
        RECT 62.520 153.435 62.910 153.440 ;
        RECT 61.745 153.430 62.910 153.435 ;
        RECT 61.745 153.395 62.880 153.430 ;
        RECT 61.745 153.370 62.845 153.395 ;
        RECT 61.745 153.340 62.815 153.370 ;
        RECT 61.745 153.310 62.795 153.340 ;
        RECT 61.745 153.280 62.775 153.310 ;
        RECT 61.745 153.270 62.705 153.280 ;
        RECT 61.745 153.260 62.680 153.270 ;
        RECT 61.745 153.245 62.660 153.260 ;
        RECT 61.745 153.230 62.640 153.245 ;
        RECT 61.850 153.220 62.635 153.230 ;
        RECT 61.850 153.185 62.620 153.220 ;
        RECT 61.405 152.355 61.680 153.055 ;
        RECT 61.850 152.935 62.605 153.185 ;
        RECT 62.775 152.865 63.105 153.110 ;
        RECT 63.275 153.010 63.535 153.460 ;
        RECT 62.920 152.840 63.105 152.865 ;
        RECT 62.920 152.740 63.535 152.840 ;
        RECT 61.850 152.185 62.105 152.730 ;
        RECT 62.275 152.355 62.755 152.695 ;
        RECT 62.930 152.185 63.535 152.740 ;
        RECT 63.705 152.185 63.995 153.350 ;
        RECT 64.165 153.325 64.445 153.995 ;
        RECT 64.720 153.935 65.845 154.105 ;
        RECT 64.720 153.825 65.170 153.935 ;
        RECT 64.615 153.495 65.170 153.825 ;
        RECT 66.035 153.765 66.435 154.565 ;
        RECT 66.835 154.275 67.105 154.735 ;
        RECT 67.275 154.105 67.560 154.565 ;
        RECT 64.165 152.355 64.550 153.325 ;
        RECT 64.720 153.035 65.170 153.495 ;
        RECT 65.340 153.205 66.435 153.765 ;
        RECT 64.720 152.815 65.845 153.035 ;
        RECT 64.720 152.185 65.045 152.645 ;
        RECT 65.565 152.355 65.845 152.815 ;
        RECT 66.035 152.355 66.435 153.205 ;
        RECT 66.605 153.935 67.560 154.105 ;
        RECT 67.935 154.185 68.105 154.475 ;
        RECT 68.275 154.355 68.605 154.735 ;
        RECT 67.935 154.015 68.600 154.185 ;
        RECT 66.605 153.035 66.815 153.935 ;
        RECT 66.985 153.205 67.675 153.765 ;
        RECT 67.850 153.195 68.200 153.845 ;
        RECT 66.605 152.815 67.560 153.035 ;
        RECT 68.370 153.025 68.600 154.015 ;
        RECT 66.835 152.185 67.105 152.645 ;
        RECT 67.275 152.355 67.560 152.815 ;
        RECT 67.935 152.855 68.600 153.025 ;
        RECT 67.935 152.355 68.105 152.855 ;
        RECT 68.275 152.185 68.605 152.685 ;
        RECT 68.775 152.355 68.960 154.475 ;
        RECT 69.215 154.275 69.465 154.735 ;
        RECT 69.635 154.285 69.970 154.455 ;
        RECT 70.165 154.285 70.840 154.455 ;
        RECT 69.635 154.145 69.805 154.285 ;
        RECT 69.130 153.155 69.410 154.105 ;
        RECT 69.580 154.015 69.805 154.145 ;
        RECT 69.580 152.910 69.750 154.015 ;
        RECT 69.975 153.865 70.500 154.085 ;
        RECT 69.920 153.100 70.160 153.695 ;
        RECT 70.330 153.165 70.500 153.865 ;
        RECT 70.670 153.505 70.840 154.285 ;
        RECT 71.160 154.235 71.530 154.735 ;
        RECT 71.710 154.285 72.115 154.455 ;
        RECT 72.285 154.285 73.070 154.455 ;
        RECT 71.710 154.055 71.880 154.285 ;
        RECT 71.050 153.755 71.880 154.055 ;
        RECT 72.265 153.785 72.730 154.115 ;
        RECT 71.050 153.725 71.250 153.755 ;
        RECT 71.370 153.505 71.540 153.575 ;
        RECT 70.670 153.335 71.540 153.505 ;
        RECT 71.030 153.245 71.540 153.335 ;
        RECT 69.580 152.780 69.885 152.910 ;
        RECT 70.330 152.800 70.860 153.165 ;
        RECT 69.200 152.185 69.465 152.645 ;
        RECT 69.635 152.355 69.885 152.780 ;
        RECT 71.030 152.630 71.200 153.245 ;
        RECT 70.095 152.460 71.200 152.630 ;
        RECT 71.370 152.185 71.540 152.985 ;
        RECT 71.710 152.685 71.880 153.755 ;
        RECT 72.050 152.855 72.240 153.575 ;
        RECT 72.410 152.825 72.730 153.785 ;
        RECT 72.900 153.825 73.070 154.285 ;
        RECT 73.345 154.205 73.555 154.735 ;
        RECT 73.815 153.995 74.145 154.520 ;
        RECT 74.315 154.125 74.485 154.735 ;
        RECT 74.655 154.080 74.985 154.515 ;
        RECT 74.655 153.995 75.035 154.080 ;
        RECT 73.945 153.825 74.145 153.995 ;
        RECT 74.810 153.955 75.035 153.995 ;
        RECT 72.900 153.495 73.775 153.825 ;
        RECT 73.945 153.495 74.695 153.825 ;
        RECT 71.710 152.355 71.960 152.685 ;
        RECT 72.900 152.655 73.070 153.495 ;
        RECT 73.945 153.290 74.135 153.495 ;
        RECT 74.865 153.375 75.035 153.955 ;
        RECT 74.820 153.325 75.035 153.375 ;
        RECT 73.240 152.915 74.135 153.290 ;
        RECT 74.645 153.245 75.035 153.325 ;
        RECT 75.205 153.995 75.590 154.565 ;
        RECT 75.760 154.275 76.085 154.735 ;
        RECT 76.605 154.105 76.885 154.565 ;
        RECT 75.205 153.325 75.485 153.995 ;
        RECT 75.760 153.935 76.885 154.105 ;
        RECT 75.760 153.825 76.210 153.935 ;
        RECT 75.655 153.495 76.210 153.825 ;
        RECT 77.075 153.765 77.475 154.565 ;
        RECT 77.875 154.275 78.145 154.735 ;
        RECT 78.315 154.105 78.600 154.565 ;
        RECT 72.185 152.485 73.070 152.655 ;
        RECT 73.250 152.185 73.565 152.685 ;
        RECT 73.795 152.355 74.135 152.915 ;
        RECT 74.305 152.185 74.475 153.195 ;
        RECT 74.645 152.400 74.975 153.245 ;
        RECT 75.205 152.355 75.590 153.325 ;
        RECT 75.760 153.035 76.210 153.495 ;
        RECT 76.380 153.205 77.475 153.765 ;
        RECT 75.760 152.815 76.885 153.035 ;
        RECT 75.760 152.185 76.085 152.645 ;
        RECT 76.605 152.355 76.885 152.815 ;
        RECT 77.075 152.355 77.475 153.205 ;
        RECT 77.645 153.935 78.600 154.105 ;
        RECT 77.645 153.035 77.855 153.935 ;
        RECT 78.025 153.205 78.715 153.765 ;
        RECT 78.890 153.135 79.225 154.555 ;
        RECT 79.405 154.365 80.150 154.735 ;
        RECT 80.715 154.195 80.970 154.555 ;
        RECT 81.150 154.365 81.480 154.735 ;
        RECT 81.660 154.195 81.885 154.555 ;
        RECT 79.400 154.005 81.885 154.195 ;
        RECT 82.195 154.185 82.365 154.565 ;
        RECT 82.580 154.355 82.910 154.735 ;
        RECT 82.195 154.015 82.910 154.185 ;
        RECT 79.400 153.315 79.625 154.005 ;
        RECT 79.825 153.495 80.105 153.825 ;
        RECT 80.285 153.495 80.860 153.825 ;
        RECT 81.040 153.495 81.475 153.825 ;
        RECT 81.655 153.495 81.925 153.825 ;
        RECT 82.105 153.465 82.460 153.835 ;
        RECT 82.740 153.825 82.910 154.015 ;
        RECT 83.080 153.990 83.335 154.565 ;
        RECT 82.740 153.495 82.995 153.825 ;
        RECT 79.400 153.135 81.895 153.315 ;
        RECT 82.740 153.285 82.910 153.495 ;
        RECT 77.645 152.815 78.600 153.035 ;
        RECT 77.875 152.185 78.145 152.645 ;
        RECT 78.315 152.355 78.600 152.815 ;
        RECT 78.890 152.365 79.155 153.135 ;
        RECT 79.325 152.185 79.655 152.905 ;
        RECT 79.845 152.725 81.035 152.955 ;
        RECT 79.845 152.365 80.105 152.725 ;
        RECT 80.275 152.185 80.605 152.555 ;
        RECT 80.775 152.365 81.035 152.725 ;
        RECT 81.605 152.365 81.895 153.135 ;
        RECT 82.195 153.115 82.910 153.285 ;
        RECT 83.165 153.260 83.335 153.990 ;
        RECT 83.510 153.895 83.770 154.735 ;
        RECT 82.195 152.355 82.365 153.115 ;
        RECT 82.580 152.185 82.910 152.945 ;
        RECT 83.080 152.355 83.335 153.260 ;
        RECT 83.510 152.185 83.770 153.335 ;
        RECT 83.950 153.135 84.285 154.555 ;
        RECT 84.465 154.365 85.210 154.735 ;
        RECT 85.775 154.195 86.030 154.555 ;
        RECT 86.210 154.365 86.540 154.735 ;
        RECT 86.720 154.195 86.945 154.555 ;
        RECT 84.460 154.005 86.945 154.195 ;
        RECT 87.165 154.060 87.425 154.565 ;
        RECT 87.605 154.355 87.935 154.735 ;
        RECT 88.115 154.185 88.285 154.565 ;
        RECT 84.460 153.315 84.685 154.005 ;
        RECT 84.885 153.495 85.165 153.825 ;
        RECT 85.345 153.495 85.920 153.825 ;
        RECT 86.100 153.495 86.535 153.825 ;
        RECT 86.715 153.495 86.985 153.825 ;
        RECT 84.460 153.135 86.955 153.315 ;
        RECT 83.950 152.365 84.215 153.135 ;
        RECT 84.385 152.185 84.715 152.905 ;
        RECT 84.905 152.725 86.095 152.955 ;
        RECT 84.905 152.365 85.165 152.725 ;
        RECT 85.335 152.185 85.665 152.555 ;
        RECT 85.835 152.365 86.095 152.725 ;
        RECT 86.665 152.365 86.955 153.135 ;
        RECT 87.165 153.260 87.345 154.060 ;
        RECT 87.620 154.015 88.285 154.185 ;
        RECT 87.620 153.760 87.790 154.015 ;
        RECT 88.545 153.985 89.755 154.735 ;
        RECT 87.515 153.430 87.790 153.760 ;
        RECT 88.015 153.465 88.355 153.835 ;
        RECT 87.620 153.285 87.790 153.430 ;
        RECT 87.165 152.355 87.435 153.260 ;
        RECT 87.620 153.115 88.295 153.285 ;
        RECT 87.605 152.185 87.935 152.945 ;
        RECT 88.115 152.355 88.295 153.115 ;
        RECT 88.545 153.275 89.065 153.815 ;
        RECT 89.235 153.445 89.755 153.985 ;
        RECT 88.545 152.185 89.755 153.275 ;
        RECT 100.140 152.510 100.810 155.770 ;
        RECT 101.480 155.200 105.520 155.370 ;
        RECT 101.140 153.140 101.310 155.140 ;
        RECT 105.690 153.140 105.860 155.140 ;
        RECT 101.480 152.910 105.520 153.080 ;
        RECT 106.200 152.510 106.370 155.770 ;
        RECT 100.140 152.500 106.370 152.510 ;
        RECT 107.960 161.770 117.790 161.810 ;
        RECT 120.510 161.790 126.250 161.800 ;
        RECT 107.960 161.640 118.590 161.770 ;
        RECT 107.960 159.380 108.130 161.640 ;
        RECT 108.855 161.070 116.895 161.240 ;
        RECT 108.470 160.010 108.640 161.010 ;
        RECT 117.110 160.010 117.280 161.010 ;
        RECT 108.855 159.780 116.895 159.950 ;
        RECT 117.620 159.380 118.590 161.640 ;
        RECT 107.960 159.210 118.590 159.380 ;
        RECT 107.960 155.950 108.130 159.210 ;
        RECT 108.855 158.640 116.895 158.810 ;
        RECT 108.470 156.580 108.640 158.580 ;
        RECT 117.110 156.580 117.280 158.580 ;
        RECT 108.855 156.350 116.895 156.520 ;
        RECT 117.620 155.950 118.590 159.210 ;
        RECT 107.960 155.780 118.590 155.950 ;
        RECT 107.960 152.520 108.130 155.780 ;
        RECT 108.855 155.210 116.895 155.380 ;
        RECT 108.470 153.150 108.640 155.150 ;
        RECT 117.110 153.150 117.280 155.150 ;
        RECT 108.855 152.920 116.895 153.090 ;
        RECT 117.620 152.520 118.590 155.780 ;
        RECT 100.140 152.400 106.380 152.500 ;
        RECT 12.100 152.015 89.840 152.185 ;
        RECT 12.185 150.925 13.395 152.015 ;
        RECT 13.565 151.580 18.910 152.015 ;
        RECT 12.185 150.215 12.705 150.755 ;
        RECT 12.875 150.385 13.395 150.925 ;
        RECT 12.185 149.465 13.395 150.215 ;
        RECT 15.150 150.010 15.490 150.840 ;
        RECT 16.970 150.330 17.320 151.580 ;
        RECT 19.085 150.925 22.595 152.015 ;
        RECT 23.230 151.590 23.565 152.015 ;
        RECT 23.735 151.410 23.920 151.815 ;
        RECT 19.085 150.235 20.735 150.755 ;
        RECT 20.905 150.405 22.595 150.925 ;
        RECT 23.255 151.235 23.920 151.410 ;
        RECT 24.125 151.235 24.455 152.015 ;
        RECT 13.565 149.465 18.910 150.010 ;
        RECT 19.085 149.465 22.595 150.235 ;
        RECT 23.255 150.205 23.595 151.235 ;
        RECT 24.625 151.045 24.895 151.815 ;
        RECT 23.765 150.875 24.895 151.045 ;
        RECT 23.765 150.375 24.015 150.875 ;
        RECT 23.255 150.035 23.940 150.205 ;
        RECT 24.195 150.125 24.555 150.705 ;
        RECT 23.230 149.465 23.565 149.865 ;
        RECT 23.735 149.635 23.940 150.035 ;
        RECT 24.725 149.965 24.895 150.875 ;
        RECT 25.065 150.850 25.355 152.015 ;
        RECT 25.525 151.580 30.870 152.015 ;
        RECT 31.045 151.580 36.390 152.015 ;
        RECT 24.150 149.465 24.425 149.945 ;
        RECT 24.635 149.635 24.895 149.965 ;
        RECT 25.065 149.465 25.355 150.190 ;
        RECT 27.110 150.010 27.450 150.840 ;
        RECT 28.930 150.330 29.280 151.580 ;
        RECT 32.630 150.010 32.970 150.840 ;
        RECT 34.450 150.330 34.800 151.580 ;
        RECT 36.565 150.925 40.075 152.015 ;
        RECT 36.565 150.235 38.215 150.755 ;
        RECT 38.385 150.405 40.075 150.925 ;
        RECT 40.285 150.875 40.515 152.015 ;
        RECT 40.685 150.865 41.015 151.845 ;
        RECT 41.185 150.875 41.395 152.015 ;
        RECT 41.625 150.875 41.885 152.015 ;
        RECT 42.055 150.865 42.385 151.845 ;
        RECT 42.555 150.875 42.835 152.015 ;
        RECT 43.005 150.925 44.215 152.015 ;
        RECT 40.265 150.455 40.595 150.705 ;
        RECT 25.525 149.465 30.870 150.010 ;
        RECT 31.045 149.465 36.390 150.010 ;
        RECT 36.565 149.465 40.075 150.235 ;
        RECT 40.285 149.465 40.515 150.285 ;
        RECT 40.765 150.265 41.015 150.865 ;
        RECT 41.645 150.455 41.980 150.705 ;
        RECT 40.685 149.635 41.015 150.265 ;
        RECT 41.185 149.465 41.395 150.285 ;
        RECT 42.150 150.265 42.320 150.865 ;
        RECT 42.490 150.435 42.825 150.705 ;
        RECT 41.625 149.635 42.320 150.265 ;
        RECT 42.525 149.465 42.835 150.265 ;
        RECT 43.005 150.215 43.525 150.755 ;
        RECT 43.695 150.385 44.215 150.925 ;
        RECT 44.385 150.875 44.770 151.845 ;
        RECT 44.940 151.555 45.265 152.015 ;
        RECT 45.785 151.385 46.065 151.845 ;
        RECT 44.940 151.165 46.065 151.385 ;
        RECT 43.005 149.465 44.215 150.215 ;
        RECT 44.385 150.205 44.665 150.875 ;
        RECT 44.940 150.705 45.390 151.165 ;
        RECT 46.255 150.995 46.655 151.845 ;
        RECT 47.055 151.555 47.325 152.015 ;
        RECT 47.495 151.385 47.780 151.845 ;
        RECT 44.835 150.375 45.390 150.705 ;
        RECT 45.560 150.435 46.655 150.995 ;
        RECT 44.940 150.265 45.390 150.375 ;
        RECT 44.385 149.635 44.770 150.205 ;
        RECT 44.940 150.095 46.065 150.265 ;
        RECT 44.940 149.465 45.265 149.925 ;
        RECT 45.785 149.635 46.065 150.095 ;
        RECT 46.255 149.635 46.655 150.435 ;
        RECT 46.825 151.165 47.780 151.385 ;
        RECT 46.825 150.265 47.035 151.165 ;
        RECT 47.205 150.435 47.895 150.995 ;
        RECT 48.065 150.925 49.275 152.015 ;
        RECT 46.825 150.095 47.780 150.265 ;
        RECT 47.055 149.465 47.325 149.925 ;
        RECT 47.495 149.635 47.780 150.095 ;
        RECT 48.065 150.215 48.585 150.755 ;
        RECT 48.755 150.385 49.275 150.925 ;
        RECT 49.455 150.875 49.785 152.015 ;
        RECT 50.315 151.045 50.645 151.830 ;
        RECT 49.965 150.875 50.645 151.045 ;
        RECT 49.445 150.455 49.795 150.705 ;
        RECT 49.965 150.275 50.135 150.875 ;
        RECT 50.825 150.850 51.115 152.015 ;
        RECT 51.285 151.460 51.890 152.015 ;
        RECT 52.065 151.505 52.545 151.845 ;
        RECT 52.715 151.470 52.970 152.015 ;
        RECT 51.285 151.360 51.900 151.460 ;
        RECT 51.715 151.335 51.900 151.360 ;
        RECT 51.285 150.740 51.545 151.190 ;
        RECT 51.715 151.090 52.045 151.335 ;
        RECT 52.215 151.015 52.970 151.265 ;
        RECT 53.140 151.145 53.415 151.845 ;
        RECT 52.200 150.980 52.970 151.015 ;
        RECT 52.185 150.970 52.970 150.980 ;
        RECT 52.180 150.955 53.075 150.970 ;
        RECT 52.160 150.940 53.075 150.955 ;
        RECT 52.140 150.930 53.075 150.940 ;
        RECT 52.115 150.920 53.075 150.930 ;
        RECT 52.045 150.890 53.075 150.920 ;
        RECT 52.025 150.860 53.075 150.890 ;
        RECT 52.005 150.830 53.075 150.860 ;
        RECT 51.975 150.805 53.075 150.830 ;
        RECT 51.940 150.770 53.075 150.805 ;
        RECT 51.910 150.765 53.075 150.770 ;
        RECT 51.910 150.760 52.300 150.765 ;
        RECT 51.910 150.750 52.275 150.760 ;
        RECT 51.910 150.745 52.260 150.750 ;
        RECT 51.910 150.740 52.245 150.745 ;
        RECT 51.285 150.735 52.245 150.740 ;
        RECT 51.285 150.725 52.235 150.735 ;
        RECT 51.285 150.720 52.225 150.725 ;
        RECT 51.285 150.710 52.215 150.720 ;
        RECT 50.305 150.455 50.655 150.705 ;
        RECT 51.285 150.700 52.210 150.710 ;
        RECT 51.285 150.695 52.205 150.700 ;
        RECT 51.285 150.680 52.195 150.695 ;
        RECT 51.285 150.665 52.190 150.680 ;
        RECT 51.285 150.640 52.180 150.665 ;
        RECT 51.285 150.570 52.175 150.640 ;
        RECT 48.065 149.465 49.275 150.215 ;
        RECT 49.455 149.465 49.725 150.275 ;
        RECT 49.895 149.635 50.225 150.275 ;
        RECT 50.395 149.465 50.635 150.275 ;
        RECT 50.825 149.465 51.115 150.190 ;
        RECT 51.285 150.015 51.835 150.400 ;
        RECT 52.005 149.845 52.175 150.570 ;
        RECT 51.285 149.675 52.175 149.845 ;
        RECT 52.345 150.170 52.675 150.595 ;
        RECT 52.845 150.370 53.075 150.765 ;
        RECT 52.345 149.685 52.565 150.170 ;
        RECT 53.245 150.115 53.415 151.145 ;
        RECT 53.585 150.925 55.255 152.015 ;
        RECT 52.735 149.465 52.985 150.005 ;
        RECT 53.155 149.635 53.415 150.115 ;
        RECT 53.585 150.235 54.335 150.755 ;
        RECT 54.505 150.405 55.255 150.925 ;
        RECT 55.430 150.865 55.690 152.015 ;
        RECT 55.865 150.940 56.120 151.845 ;
        RECT 56.290 151.255 56.620 152.015 ;
        RECT 56.835 151.085 57.005 151.845 ;
        RECT 53.585 149.465 55.255 150.235 ;
        RECT 55.430 149.465 55.690 150.305 ;
        RECT 55.865 150.210 56.035 150.940 ;
        RECT 56.290 150.915 57.005 151.085 ;
        RECT 56.290 150.705 56.460 150.915 ;
        RECT 57.270 150.875 57.605 151.845 ;
        RECT 57.775 150.875 57.945 152.015 ;
        RECT 58.115 151.675 60.145 151.845 ;
        RECT 56.205 150.375 56.460 150.705 ;
        RECT 55.865 149.635 56.120 150.210 ;
        RECT 56.290 150.185 56.460 150.375 ;
        RECT 56.740 150.365 57.095 150.735 ;
        RECT 57.270 150.205 57.440 150.875 ;
        RECT 58.115 150.705 58.285 151.675 ;
        RECT 57.610 150.375 57.865 150.705 ;
        RECT 58.090 150.375 58.285 150.705 ;
        RECT 58.455 151.335 59.580 151.505 ;
        RECT 57.695 150.205 57.865 150.375 ;
        RECT 58.455 150.205 58.625 151.335 ;
        RECT 56.290 150.015 57.005 150.185 ;
        RECT 56.290 149.465 56.620 149.845 ;
        RECT 56.835 149.635 57.005 150.015 ;
        RECT 57.270 149.635 57.525 150.205 ;
        RECT 57.695 150.035 58.625 150.205 ;
        RECT 58.795 150.995 59.805 151.165 ;
        RECT 58.795 150.195 58.965 150.995 ;
        RECT 58.450 150.000 58.625 150.035 ;
        RECT 57.695 149.465 58.025 149.865 ;
        RECT 58.450 149.635 58.980 150.000 ;
        RECT 59.170 149.975 59.445 150.795 ;
        RECT 59.165 149.805 59.445 149.975 ;
        RECT 59.170 149.635 59.445 149.805 ;
        RECT 59.615 149.635 59.805 150.995 ;
        RECT 59.975 151.010 60.145 151.675 ;
        RECT 60.315 151.255 60.485 152.015 ;
        RECT 60.720 151.255 61.235 151.665 ;
        RECT 59.975 150.820 60.725 151.010 ;
        RECT 60.895 150.445 61.235 151.255 ;
        RECT 61.415 150.875 61.745 152.015 ;
        RECT 60.005 150.275 61.235 150.445 ;
        RECT 59.985 149.465 60.495 150.000 ;
        RECT 60.715 149.670 60.960 150.275 ;
        RECT 61.405 150.125 61.745 150.705 ;
        RECT 61.915 150.675 62.275 151.845 ;
        RECT 62.475 150.845 62.805 152.015 ;
        RECT 63.005 150.675 63.335 151.845 ;
        RECT 63.535 150.845 63.865 152.015 ;
        RECT 64.740 151.385 65.025 151.845 ;
        RECT 65.195 151.555 65.465 152.015 ;
        RECT 64.740 151.165 65.695 151.385 ;
        RECT 61.915 150.395 63.335 150.675 ;
        RECT 64.625 150.435 65.315 150.995 ;
        RECT 61.915 150.060 62.275 150.395 ;
        RECT 65.485 150.265 65.695 151.165 ;
        RECT 61.415 149.465 61.745 149.955 ;
        RECT 61.915 149.635 62.535 150.060 ;
        RECT 62.995 149.465 63.325 150.155 ;
        RECT 64.740 150.095 65.695 150.265 ;
        RECT 65.865 150.995 66.265 151.845 ;
        RECT 66.455 151.385 66.735 151.845 ;
        RECT 67.255 151.555 67.580 152.015 ;
        RECT 66.455 151.165 67.580 151.385 ;
        RECT 65.865 150.435 66.960 150.995 ;
        RECT 67.130 150.705 67.580 151.165 ;
        RECT 67.750 150.875 68.135 151.845 ;
        RECT 68.395 151.345 68.565 151.845 ;
        RECT 68.735 151.515 69.065 152.015 ;
        RECT 68.395 151.175 69.060 151.345 ;
        RECT 64.740 149.635 65.025 150.095 ;
        RECT 65.195 149.465 65.465 149.925 ;
        RECT 65.865 149.635 66.265 150.435 ;
        RECT 67.130 150.375 67.685 150.705 ;
        RECT 67.130 150.265 67.580 150.375 ;
        RECT 66.455 150.095 67.580 150.265 ;
        RECT 67.855 150.205 68.135 150.875 ;
        RECT 68.310 150.355 68.660 151.005 ;
        RECT 66.455 149.635 66.735 150.095 ;
        RECT 67.255 149.465 67.580 149.925 ;
        RECT 67.750 149.635 68.135 150.205 ;
        RECT 68.830 150.185 69.060 151.175 ;
        RECT 68.395 150.015 69.060 150.185 ;
        RECT 68.395 149.725 68.565 150.015 ;
        RECT 68.735 149.465 69.065 149.845 ;
        RECT 69.235 149.725 69.420 151.845 ;
        RECT 69.660 151.555 69.925 152.015 ;
        RECT 70.095 151.420 70.345 151.845 ;
        RECT 70.555 151.570 71.660 151.740 ;
        RECT 70.040 151.290 70.345 151.420 ;
        RECT 69.590 150.095 69.870 151.045 ;
        RECT 70.040 150.185 70.210 151.290 ;
        RECT 70.380 150.505 70.620 151.100 ;
        RECT 70.790 151.035 71.320 151.400 ;
        RECT 70.790 150.335 70.960 151.035 ;
        RECT 71.490 150.955 71.660 151.570 ;
        RECT 71.830 151.215 72.000 152.015 ;
        RECT 72.170 151.515 72.420 151.845 ;
        RECT 72.645 151.545 73.530 151.715 ;
        RECT 71.490 150.865 72.000 150.955 ;
        RECT 70.040 150.055 70.265 150.185 ;
        RECT 70.435 150.115 70.960 150.335 ;
        RECT 71.130 150.695 72.000 150.865 ;
        RECT 69.675 149.465 69.925 149.925 ;
        RECT 70.095 149.915 70.265 150.055 ;
        RECT 71.130 149.915 71.300 150.695 ;
        RECT 71.830 150.625 72.000 150.695 ;
        RECT 71.510 150.445 71.710 150.475 ;
        RECT 72.170 150.445 72.340 151.515 ;
        RECT 72.510 150.625 72.700 151.345 ;
        RECT 71.510 150.145 72.340 150.445 ;
        RECT 72.870 150.415 73.190 151.375 ;
        RECT 70.095 149.745 70.430 149.915 ;
        RECT 70.625 149.745 71.300 149.915 ;
        RECT 71.620 149.465 71.990 149.965 ;
        RECT 72.170 149.915 72.340 150.145 ;
        RECT 72.725 150.085 73.190 150.415 ;
        RECT 73.360 150.705 73.530 151.545 ;
        RECT 73.710 151.515 74.025 152.015 ;
        RECT 74.255 151.285 74.595 151.845 ;
        RECT 73.700 150.910 74.595 151.285 ;
        RECT 74.765 151.005 74.935 152.015 ;
        RECT 74.405 150.705 74.595 150.910 ;
        RECT 75.105 150.955 75.435 151.800 ;
        RECT 75.105 150.875 75.495 150.955 ;
        RECT 75.280 150.825 75.495 150.875 ;
        RECT 76.585 150.850 76.875 152.015 ;
        RECT 77.250 151.045 77.580 151.845 ;
        RECT 77.750 151.215 78.080 152.015 ;
        RECT 78.380 151.045 78.710 151.845 ;
        RECT 79.355 151.215 79.605 152.015 ;
        RECT 77.250 150.875 79.685 151.045 ;
        RECT 79.875 150.875 80.045 152.015 ;
        RECT 80.215 150.875 80.555 151.845 ;
        RECT 81.275 151.345 81.445 151.845 ;
        RECT 81.615 151.515 81.945 152.015 ;
        RECT 81.275 151.175 81.940 151.345 ;
        RECT 73.360 150.375 74.235 150.705 ;
        RECT 74.405 150.375 75.155 150.705 ;
        RECT 73.360 149.915 73.530 150.375 ;
        RECT 74.405 150.205 74.605 150.375 ;
        RECT 75.325 150.245 75.495 150.825 ;
        RECT 77.045 150.455 77.395 150.705 ;
        RECT 77.580 150.245 77.750 150.875 ;
        RECT 77.920 150.455 78.250 150.655 ;
        RECT 78.420 150.455 78.750 150.655 ;
        RECT 78.920 150.455 79.340 150.655 ;
        RECT 79.515 150.625 79.685 150.875 ;
        RECT 79.515 150.455 80.210 150.625 ;
        RECT 75.270 150.205 75.495 150.245 ;
        RECT 72.170 149.745 72.575 149.915 ;
        RECT 72.745 149.745 73.530 149.915 ;
        RECT 73.805 149.465 74.015 149.995 ;
        RECT 74.275 149.680 74.605 150.205 ;
        RECT 75.115 150.120 75.495 150.205 ;
        RECT 74.775 149.465 74.945 150.075 ;
        RECT 75.115 149.685 75.445 150.120 ;
        RECT 76.585 149.465 76.875 150.190 ;
        RECT 77.250 149.635 77.750 150.245 ;
        RECT 78.380 150.115 79.605 150.285 ;
        RECT 80.380 150.265 80.555 150.875 ;
        RECT 81.190 150.355 81.540 151.005 ;
        RECT 78.380 149.635 78.710 150.115 ;
        RECT 78.880 149.465 79.105 149.925 ;
        RECT 79.275 149.635 79.605 150.115 ;
        RECT 79.795 149.465 80.045 150.265 ;
        RECT 80.215 149.635 80.555 150.265 ;
        RECT 81.710 150.185 81.940 151.175 ;
        RECT 81.275 150.015 81.940 150.185 ;
        RECT 81.275 149.725 81.445 150.015 ;
        RECT 81.615 149.465 81.945 149.845 ;
        RECT 82.115 149.725 82.300 151.845 ;
        RECT 82.540 151.555 82.805 152.015 ;
        RECT 82.975 151.420 83.225 151.845 ;
        RECT 83.435 151.570 84.540 151.740 ;
        RECT 82.920 151.290 83.225 151.420 ;
        RECT 82.470 150.095 82.750 151.045 ;
        RECT 82.920 150.185 83.090 151.290 ;
        RECT 83.260 150.505 83.500 151.100 ;
        RECT 83.670 151.035 84.200 151.400 ;
        RECT 83.670 150.335 83.840 151.035 ;
        RECT 84.370 150.955 84.540 151.570 ;
        RECT 84.710 151.215 84.880 152.015 ;
        RECT 85.050 151.515 85.300 151.845 ;
        RECT 85.525 151.545 86.410 151.715 ;
        RECT 84.370 150.865 84.880 150.955 ;
        RECT 82.920 150.055 83.145 150.185 ;
        RECT 83.315 150.115 83.840 150.335 ;
        RECT 84.010 150.695 84.880 150.865 ;
        RECT 82.555 149.465 82.805 149.925 ;
        RECT 82.975 149.915 83.145 150.055 ;
        RECT 84.010 149.915 84.180 150.695 ;
        RECT 84.710 150.625 84.880 150.695 ;
        RECT 84.390 150.445 84.590 150.475 ;
        RECT 85.050 150.445 85.220 151.515 ;
        RECT 85.390 150.625 85.580 151.345 ;
        RECT 84.390 150.145 85.220 150.445 ;
        RECT 85.750 150.415 86.070 151.375 ;
        RECT 82.975 149.745 83.310 149.915 ;
        RECT 83.505 149.745 84.180 149.915 ;
        RECT 84.500 149.465 84.870 149.965 ;
        RECT 85.050 149.915 85.220 150.145 ;
        RECT 85.605 150.085 86.070 150.415 ;
        RECT 86.240 150.705 86.410 151.545 ;
        RECT 86.590 151.515 86.905 152.015 ;
        RECT 87.135 151.285 87.475 151.845 ;
        RECT 86.580 150.910 87.475 151.285 ;
        RECT 87.645 151.005 87.815 152.015 ;
        RECT 87.285 150.705 87.475 150.910 ;
        RECT 87.985 150.955 88.315 151.800 ;
        RECT 87.985 150.875 88.375 150.955 ;
        RECT 88.160 150.825 88.375 150.875 ;
        RECT 86.240 150.375 87.115 150.705 ;
        RECT 87.285 150.375 88.035 150.705 ;
        RECT 86.240 149.915 86.410 150.375 ;
        RECT 87.285 150.205 87.485 150.375 ;
        RECT 88.205 150.245 88.375 150.825 ;
        RECT 88.545 150.925 89.755 152.015 ;
        RECT 100.130 151.840 106.380 152.400 ;
        RECT 100.130 151.820 105.300 151.840 ;
        RECT 100.130 151.750 104.120 151.820 ;
        RECT 88.545 150.385 89.065 150.925 ;
        RECT 88.150 150.205 88.375 150.245 ;
        RECT 89.235 150.215 89.755 150.755 ;
        RECT 100.130 150.480 102.050 151.750 ;
        RECT 103.560 151.740 104.120 151.750 ;
        RECT 103.790 150.650 104.120 151.740 ;
        RECT 104.490 151.270 105.530 151.440 ;
        RECT 104.490 150.830 105.530 151.000 ;
        RECT 105.700 150.970 105.870 151.300 ;
        RECT 103.950 150.430 104.120 150.650 ;
        RECT 106.210 150.430 106.380 151.840 ;
        RECT 103.950 150.260 106.380 150.430 ;
        RECT 107.960 152.350 118.590 152.520 ;
        RECT 120.020 161.630 126.250 161.790 ;
        RECT 120.020 159.370 120.690 161.630 ;
        RECT 121.360 161.060 125.400 161.230 ;
        RECT 121.020 160.000 121.190 161.000 ;
        RECT 125.570 160.000 125.740 161.000 ;
        RECT 121.360 159.770 125.400 159.940 ;
        RECT 126.080 159.370 126.250 161.630 ;
        RECT 120.020 159.200 126.250 159.370 ;
        RECT 120.020 155.940 120.690 159.200 ;
        RECT 121.360 158.630 125.400 158.800 ;
        RECT 121.020 156.570 121.190 158.570 ;
        RECT 125.570 156.570 125.740 158.570 ;
        RECT 121.360 156.340 125.400 156.510 ;
        RECT 126.080 155.940 126.250 159.200 ;
        RECT 120.020 155.770 126.250 155.940 ;
        RECT 120.020 152.510 120.690 155.770 ;
        RECT 121.360 155.200 125.400 155.370 ;
        RECT 121.020 153.140 121.190 155.140 ;
        RECT 125.570 153.140 125.740 155.140 ;
        RECT 121.360 152.910 125.400 153.080 ;
        RECT 126.080 152.510 126.250 155.770 ;
        RECT 120.020 152.500 126.250 152.510 ;
        RECT 127.840 161.770 137.670 161.810 ;
        RECT 127.840 161.640 138.470 161.770 ;
        RECT 140.590 161.740 146.330 161.750 ;
        RECT 127.840 159.380 128.010 161.640 ;
        RECT 128.735 161.070 136.775 161.240 ;
        RECT 128.350 160.010 128.520 161.010 ;
        RECT 136.990 160.010 137.160 161.010 ;
        RECT 128.735 159.780 136.775 159.950 ;
        RECT 137.500 159.380 138.470 161.640 ;
        RECT 127.840 159.210 138.470 159.380 ;
        RECT 127.840 155.950 128.010 159.210 ;
        RECT 128.735 158.640 136.775 158.810 ;
        RECT 128.350 156.580 128.520 158.580 ;
        RECT 136.990 156.580 137.160 158.580 ;
        RECT 128.735 156.350 136.775 156.520 ;
        RECT 137.500 155.950 138.470 159.210 ;
        RECT 127.840 155.780 138.470 155.950 ;
        RECT 127.840 152.520 128.010 155.780 ;
        RECT 128.735 155.210 136.775 155.380 ;
        RECT 128.350 153.150 128.520 155.150 ;
        RECT 136.990 153.150 137.160 155.150 ;
        RECT 128.735 152.920 136.775 153.090 ;
        RECT 137.500 152.520 138.470 155.780 ;
        RECT 120.020 152.400 126.260 152.500 ;
        RECT 85.050 149.745 85.455 149.915 ;
        RECT 85.625 149.745 86.410 149.915 ;
        RECT 86.685 149.465 86.895 149.995 ;
        RECT 87.155 149.680 87.485 150.205 ;
        RECT 87.995 150.120 88.375 150.205 ;
        RECT 87.655 149.465 87.825 150.075 ;
        RECT 87.995 149.685 88.325 150.120 ;
        RECT 88.545 149.465 89.755 150.215 ;
        RECT 107.960 150.090 108.130 152.350 ;
        RECT 108.855 151.780 116.895 151.950 ;
        RECT 108.470 150.720 108.640 151.720 ;
        RECT 117.110 150.720 117.280 151.720 ;
        RECT 108.855 150.490 116.895 150.660 ;
        RECT 117.620 150.090 118.590 152.350 ;
        RECT 120.010 151.840 126.260 152.400 ;
        RECT 120.010 151.820 125.180 151.840 ;
        RECT 120.010 151.750 124.000 151.820 ;
        RECT 120.010 150.480 121.930 151.750 ;
        RECT 123.440 151.740 124.000 151.750 ;
        RECT 123.670 150.650 124.000 151.740 ;
        RECT 124.370 151.270 125.410 151.440 ;
        RECT 124.370 150.830 125.410 151.000 ;
        RECT 125.580 150.970 125.750 151.300 ;
        RECT 123.830 150.430 124.000 150.650 ;
        RECT 126.090 150.430 126.260 151.840 ;
        RECT 123.830 150.260 126.260 150.430 ;
        RECT 127.840 152.350 138.470 152.520 ;
        RECT 140.100 161.580 146.330 161.740 ;
        RECT 140.100 159.320 140.770 161.580 ;
        RECT 141.440 161.010 145.480 161.180 ;
        RECT 141.100 159.950 141.270 160.950 ;
        RECT 145.650 159.950 145.820 160.950 ;
        RECT 141.440 159.720 145.480 159.890 ;
        RECT 146.160 159.320 146.330 161.580 ;
        RECT 140.100 159.150 146.330 159.320 ;
        RECT 140.100 155.890 140.770 159.150 ;
        RECT 141.440 158.580 145.480 158.750 ;
        RECT 141.100 156.520 141.270 158.520 ;
        RECT 145.650 156.520 145.820 158.520 ;
        RECT 141.440 156.290 145.480 156.460 ;
        RECT 146.160 155.890 146.330 159.150 ;
        RECT 140.100 155.720 146.330 155.890 ;
        RECT 140.100 152.460 140.770 155.720 ;
        RECT 141.440 155.150 145.480 155.320 ;
        RECT 141.100 153.090 141.270 155.090 ;
        RECT 145.650 153.090 145.820 155.090 ;
        RECT 141.440 152.860 145.480 153.030 ;
        RECT 146.160 152.460 146.330 155.720 ;
        RECT 140.100 152.450 146.330 152.460 ;
        RECT 147.920 161.720 157.750 161.760 ;
        RECT 147.920 161.590 158.550 161.720 ;
        RECT 147.920 159.330 148.090 161.590 ;
        RECT 148.815 161.020 156.855 161.190 ;
        RECT 148.430 159.960 148.600 160.960 ;
        RECT 157.070 159.960 157.240 160.960 ;
        RECT 148.815 159.730 156.855 159.900 ;
        RECT 157.580 159.330 158.550 161.590 ;
        RECT 147.920 159.160 158.550 159.330 ;
        RECT 147.920 155.900 148.090 159.160 ;
        RECT 148.815 158.590 156.855 158.760 ;
        RECT 148.430 156.530 148.600 158.530 ;
        RECT 157.070 156.530 157.240 158.530 ;
        RECT 148.815 156.300 156.855 156.470 ;
        RECT 157.580 155.900 158.550 159.160 ;
        RECT 147.920 155.730 158.550 155.900 ;
        RECT 147.920 152.470 148.090 155.730 ;
        RECT 148.815 155.160 156.855 155.330 ;
        RECT 148.430 153.100 148.600 155.100 ;
        RECT 157.070 153.100 157.240 155.100 ;
        RECT 148.815 152.870 156.855 153.040 ;
        RECT 157.580 152.470 158.550 155.730 ;
        RECT 140.100 152.350 146.340 152.450 ;
        RECT 107.960 150.060 118.590 150.090 ;
        RECT 127.840 150.090 128.010 152.350 ;
        RECT 128.735 151.780 136.775 151.950 ;
        RECT 128.350 150.720 128.520 151.720 ;
        RECT 136.990 150.720 137.160 151.720 ;
        RECT 128.735 150.490 136.775 150.660 ;
        RECT 137.500 150.090 138.470 152.350 ;
        RECT 140.090 151.790 146.340 152.350 ;
        RECT 140.090 151.770 145.260 151.790 ;
        RECT 140.090 151.700 144.080 151.770 ;
        RECT 140.090 150.430 142.010 151.700 ;
        RECT 143.520 151.690 144.080 151.700 ;
        RECT 143.750 150.600 144.080 151.690 ;
        RECT 144.450 151.220 145.490 151.390 ;
        RECT 144.450 150.780 145.490 150.950 ;
        RECT 145.660 150.920 145.830 151.250 ;
        RECT 143.910 150.380 144.080 150.600 ;
        RECT 146.170 150.380 146.340 151.790 ;
        RECT 143.910 150.210 146.340 150.380 ;
        RECT 147.920 152.300 158.550 152.470 ;
        RECT 127.840 150.060 138.470 150.090 ;
        RECT 107.930 149.950 118.590 150.060 ;
        RECT 127.810 149.950 138.470 150.060 ;
        RECT 147.920 150.040 148.090 152.300 ;
        RECT 148.815 151.730 156.855 151.900 ;
        RECT 148.430 150.670 148.600 151.670 ;
        RECT 157.070 150.670 157.240 151.670 ;
        RECT 148.815 150.440 156.855 150.610 ;
        RECT 157.580 150.040 158.550 152.300 ;
        RECT 147.920 150.010 158.550 150.040 ;
        RECT 106.180 149.900 118.590 149.950 ;
        RECT 126.060 149.900 138.470 149.950 ;
        RECT 147.890 149.900 158.550 150.010 ;
        RECT 101.840 149.730 118.590 149.900 ;
        RECT 12.100 149.295 89.840 149.465 ;
        RECT 12.185 148.545 13.395 149.295 ;
        RECT 13.565 148.750 18.910 149.295 ;
        RECT 12.185 148.005 12.705 148.545 ;
        RECT 12.875 147.835 13.395 148.375 ;
        RECT 15.150 147.920 15.490 148.750 ;
        RECT 19.085 148.545 20.295 149.295 ;
        RECT 20.555 148.745 20.725 149.035 ;
        RECT 20.895 148.915 21.225 149.295 ;
        RECT 20.555 148.575 21.220 148.745 ;
        RECT 12.185 146.745 13.395 147.835 ;
        RECT 16.970 147.180 17.320 148.430 ;
        RECT 19.085 148.005 19.605 148.545 ;
        RECT 19.775 147.835 20.295 148.375 ;
        RECT 13.565 146.745 18.910 147.180 ;
        RECT 19.085 146.745 20.295 147.835 ;
        RECT 20.470 147.755 20.820 148.405 ;
        RECT 20.990 147.585 21.220 148.575 ;
        RECT 20.555 147.415 21.220 147.585 ;
        RECT 20.555 146.915 20.725 147.415 ;
        RECT 20.895 146.745 21.225 147.245 ;
        RECT 21.395 146.915 21.580 149.035 ;
        RECT 21.835 148.835 22.085 149.295 ;
        RECT 22.255 148.845 22.590 149.015 ;
        RECT 22.785 148.845 23.460 149.015 ;
        RECT 22.255 148.705 22.425 148.845 ;
        RECT 21.750 147.715 22.030 148.665 ;
        RECT 22.200 148.575 22.425 148.705 ;
        RECT 22.200 147.470 22.370 148.575 ;
        RECT 22.595 148.425 23.120 148.645 ;
        RECT 22.540 147.660 22.780 148.255 ;
        RECT 22.950 147.725 23.120 148.425 ;
        RECT 23.290 148.065 23.460 148.845 ;
        RECT 23.780 148.795 24.150 149.295 ;
        RECT 24.330 148.845 24.735 149.015 ;
        RECT 24.905 148.845 25.690 149.015 ;
        RECT 24.330 148.615 24.500 148.845 ;
        RECT 23.670 148.315 24.500 148.615 ;
        RECT 24.885 148.345 25.350 148.675 ;
        RECT 23.670 148.285 23.870 148.315 ;
        RECT 23.990 148.065 24.160 148.135 ;
        RECT 23.290 147.895 24.160 148.065 ;
        RECT 23.650 147.805 24.160 147.895 ;
        RECT 22.200 147.340 22.505 147.470 ;
        RECT 22.950 147.360 23.480 147.725 ;
        RECT 21.820 146.745 22.085 147.205 ;
        RECT 22.255 146.915 22.505 147.340 ;
        RECT 23.650 147.190 23.820 147.805 ;
        RECT 22.715 147.020 23.820 147.190 ;
        RECT 23.990 146.745 24.160 147.545 ;
        RECT 24.330 147.245 24.500 148.315 ;
        RECT 24.670 147.415 24.860 148.135 ;
        RECT 25.030 147.385 25.350 148.345 ;
        RECT 25.520 148.385 25.690 148.845 ;
        RECT 25.965 148.765 26.175 149.295 ;
        RECT 26.435 148.555 26.765 149.080 ;
        RECT 26.935 148.685 27.105 149.295 ;
        RECT 27.275 148.640 27.605 149.075 ;
        RECT 27.275 148.555 27.655 148.640 ;
        RECT 26.565 148.385 26.765 148.555 ;
        RECT 27.430 148.515 27.655 148.555 ;
        RECT 25.520 148.055 26.395 148.385 ;
        RECT 26.565 148.055 27.315 148.385 ;
        RECT 24.330 146.915 24.580 147.245 ;
        RECT 25.520 147.215 25.690 148.055 ;
        RECT 26.565 147.850 26.755 148.055 ;
        RECT 27.485 147.935 27.655 148.515 ;
        RECT 27.845 148.485 28.085 149.295 ;
        RECT 28.255 148.485 28.585 149.125 ;
        RECT 28.755 148.485 29.025 149.295 ;
        RECT 29.205 148.750 34.550 149.295 ;
        RECT 27.825 148.055 28.175 148.305 ;
        RECT 27.440 147.885 27.655 147.935 ;
        RECT 28.345 147.885 28.515 148.485 ;
        RECT 28.685 148.055 29.035 148.305 ;
        RECT 30.790 147.920 31.130 148.750 ;
        RECT 34.725 148.525 37.315 149.295 ;
        RECT 37.945 148.570 38.235 149.295 ;
        RECT 38.405 148.525 40.075 149.295 ;
        RECT 25.860 147.475 26.755 147.850 ;
        RECT 27.265 147.805 27.655 147.885 ;
        RECT 24.805 147.045 25.690 147.215 ;
        RECT 25.870 146.745 26.185 147.245 ;
        RECT 26.415 146.915 26.755 147.475 ;
        RECT 26.925 146.745 27.095 147.755 ;
        RECT 27.265 146.960 27.595 147.805 ;
        RECT 27.835 147.715 28.515 147.885 ;
        RECT 27.835 146.930 28.165 147.715 ;
        RECT 28.695 146.745 29.025 147.885 ;
        RECT 32.610 147.180 32.960 148.430 ;
        RECT 34.725 148.005 35.935 148.525 ;
        RECT 36.105 147.835 37.315 148.355 ;
        RECT 38.405 148.005 39.155 148.525 ;
        RECT 40.245 148.495 40.555 149.295 ;
        RECT 40.760 148.495 41.455 149.125 ;
        RECT 41.625 148.570 41.885 149.125 ;
        RECT 42.055 148.850 42.485 149.295 ;
        RECT 42.720 148.725 42.890 149.125 ;
        RECT 43.060 148.895 43.780 149.295 ;
        RECT 40.760 148.445 40.935 148.495 ;
        RECT 29.205 146.745 34.550 147.180 ;
        RECT 34.725 146.745 37.315 147.835 ;
        RECT 37.945 146.745 38.235 147.910 ;
        RECT 39.325 147.835 40.075 148.355 ;
        RECT 40.255 148.055 40.590 148.325 ;
        RECT 40.760 147.895 40.930 148.445 ;
        RECT 41.100 148.055 41.435 148.305 ;
        RECT 38.405 146.745 40.075 147.835 ;
        RECT 40.245 146.745 40.525 147.885 ;
        RECT 40.695 146.915 41.025 147.895 ;
        RECT 41.195 146.745 41.455 147.885 ;
        RECT 41.625 147.855 41.800 148.570 ;
        RECT 42.720 148.555 43.600 148.725 ;
        RECT 43.950 148.680 44.120 149.125 ;
        RECT 44.695 148.785 45.095 149.295 ;
        RECT 41.970 148.055 42.225 148.385 ;
        RECT 41.625 146.915 41.885 147.855 ;
        RECT 42.055 147.575 42.225 148.055 ;
        RECT 42.450 147.765 42.780 148.385 ;
        RECT 42.950 148.005 43.240 148.385 ;
        RECT 43.430 147.835 43.600 148.555 ;
        RECT 43.080 147.665 43.600 147.835 ;
        RECT 43.770 148.510 44.120 148.680 ;
        RECT 42.055 147.405 42.815 147.575 ;
        RECT 43.080 147.475 43.250 147.665 ;
        RECT 43.770 147.485 43.940 148.510 ;
        RECT 44.360 148.025 44.620 148.615 ;
        RECT 44.140 147.725 44.620 148.025 ;
        RECT 44.820 147.725 45.080 148.615 ;
        RECT 45.340 148.555 45.955 149.125 ;
        RECT 46.125 148.785 46.340 149.295 ;
        RECT 46.570 148.785 46.850 149.115 ;
        RECT 47.030 148.785 47.270 149.295 ;
        RECT 42.645 147.180 42.815 147.405 ;
        RECT 43.530 147.315 43.940 147.485 ;
        RECT 44.115 147.375 45.055 147.545 ;
        RECT 43.530 147.180 43.785 147.315 ;
        RECT 42.055 146.745 42.385 147.145 ;
        RECT 42.645 147.010 43.785 147.180 ;
        RECT 44.115 147.125 44.285 147.375 ;
        RECT 43.530 146.915 43.785 147.010 ;
        RECT 43.955 146.955 44.285 147.125 ;
        RECT 44.455 146.745 44.705 147.205 ;
        RECT 44.875 146.915 45.055 147.375 ;
        RECT 45.340 147.535 45.655 148.555 ;
        RECT 45.825 147.885 45.995 148.385 ;
        RECT 46.245 148.055 46.510 148.615 ;
        RECT 46.680 147.885 46.850 148.785 ;
        RECT 47.605 148.620 47.865 149.125 ;
        RECT 48.045 148.915 48.375 149.295 ;
        RECT 48.555 148.745 48.725 149.125 ;
        RECT 47.020 148.055 47.375 148.615 ;
        RECT 45.825 147.715 47.250 147.885 ;
        RECT 45.340 146.915 45.875 147.535 ;
        RECT 46.045 146.745 46.375 147.545 ;
        RECT 46.860 147.540 47.250 147.715 ;
        RECT 47.605 147.820 47.785 148.620 ;
        RECT 48.060 148.575 48.725 148.745 ;
        RECT 48.060 148.320 48.230 148.575 ;
        RECT 48.985 148.545 50.195 149.295 ;
        RECT 50.370 148.555 50.625 149.125 ;
        RECT 50.795 148.895 51.125 149.295 ;
        RECT 51.550 148.760 52.080 149.125 ;
        RECT 51.550 148.725 51.725 148.760 ;
        RECT 50.795 148.555 51.725 148.725 ;
        RECT 47.955 147.990 48.230 148.320 ;
        RECT 48.455 148.025 48.795 148.395 ;
        RECT 48.985 148.005 49.505 148.545 ;
        RECT 48.060 147.845 48.230 147.990 ;
        RECT 47.605 146.915 47.875 147.820 ;
        RECT 48.060 147.675 48.735 147.845 ;
        RECT 49.675 147.835 50.195 148.375 ;
        RECT 48.045 146.745 48.375 147.505 ;
        RECT 48.555 146.915 48.735 147.675 ;
        RECT 48.985 146.745 50.195 147.835 ;
        RECT 50.370 147.885 50.540 148.555 ;
        RECT 50.795 148.385 50.965 148.555 ;
        RECT 50.710 148.055 50.965 148.385 ;
        RECT 51.190 148.055 51.385 148.385 ;
        RECT 50.370 146.915 50.705 147.885 ;
        RECT 50.875 146.745 51.045 147.885 ;
        RECT 51.215 147.085 51.385 148.055 ;
        RECT 51.555 147.425 51.725 148.555 ;
        RECT 51.895 147.765 52.065 148.565 ;
        RECT 52.270 148.275 52.545 149.125 ;
        RECT 52.265 148.105 52.545 148.275 ;
        RECT 52.270 147.965 52.545 148.105 ;
        RECT 52.715 147.765 52.905 149.125 ;
        RECT 53.085 148.760 53.595 149.295 ;
        RECT 53.815 148.485 54.060 149.090 ;
        RECT 54.505 148.525 58.015 149.295 ;
        RECT 58.185 148.545 59.395 149.295 ;
        RECT 59.570 148.555 59.825 149.125 ;
        RECT 59.995 148.895 60.325 149.295 ;
        RECT 60.750 148.760 61.280 149.125 ;
        RECT 61.470 148.955 61.745 149.125 ;
        RECT 61.465 148.785 61.745 148.955 ;
        RECT 60.750 148.725 60.925 148.760 ;
        RECT 59.995 148.555 60.925 148.725 ;
        RECT 53.105 148.315 54.335 148.485 ;
        RECT 51.895 147.595 52.905 147.765 ;
        RECT 53.075 147.750 53.825 147.940 ;
        RECT 51.555 147.255 52.680 147.425 ;
        RECT 53.075 147.085 53.245 147.750 ;
        RECT 53.995 147.505 54.335 148.315 ;
        RECT 54.505 148.005 56.155 148.525 ;
        RECT 56.325 147.835 58.015 148.355 ;
        RECT 58.185 148.005 58.705 148.545 ;
        RECT 58.875 147.835 59.395 148.375 ;
        RECT 51.215 146.915 53.245 147.085 ;
        RECT 53.415 146.745 53.585 147.505 ;
        RECT 53.820 147.095 54.335 147.505 ;
        RECT 54.505 146.745 58.015 147.835 ;
        RECT 58.185 146.745 59.395 147.835 ;
        RECT 59.570 147.885 59.740 148.555 ;
        RECT 59.995 148.385 60.165 148.555 ;
        RECT 59.910 148.055 60.165 148.385 ;
        RECT 60.390 148.055 60.585 148.385 ;
        RECT 59.570 146.915 59.905 147.885 ;
        RECT 60.075 146.745 60.245 147.885 ;
        RECT 60.415 147.085 60.585 148.055 ;
        RECT 60.755 147.425 60.925 148.555 ;
        RECT 61.095 147.765 61.265 148.565 ;
        RECT 61.470 147.965 61.745 148.785 ;
        RECT 61.915 147.765 62.105 149.125 ;
        RECT 62.285 148.760 62.795 149.295 ;
        RECT 63.015 148.485 63.260 149.090 ;
        RECT 63.705 148.570 63.995 149.295 ;
        RECT 64.215 148.640 64.545 149.075 ;
        RECT 64.715 148.685 64.885 149.295 ;
        RECT 64.165 148.555 64.545 148.640 ;
        RECT 65.055 148.555 65.385 149.080 ;
        RECT 65.645 148.765 65.855 149.295 ;
        RECT 66.130 148.845 66.915 149.015 ;
        RECT 67.085 148.845 67.490 149.015 ;
        RECT 64.165 148.515 64.390 148.555 ;
        RECT 62.305 148.315 63.535 148.485 ;
        RECT 61.095 147.595 62.105 147.765 ;
        RECT 62.275 147.750 63.025 147.940 ;
        RECT 60.755 147.255 61.880 147.425 ;
        RECT 62.275 147.085 62.445 147.750 ;
        RECT 63.195 147.505 63.535 148.315 ;
        RECT 64.165 147.935 64.335 148.515 ;
        RECT 65.055 148.385 65.255 148.555 ;
        RECT 66.130 148.385 66.300 148.845 ;
        RECT 64.505 148.055 65.255 148.385 ;
        RECT 65.425 148.055 66.300 148.385 ;
        RECT 60.415 146.915 62.445 147.085 ;
        RECT 62.615 146.745 62.785 147.505 ;
        RECT 63.020 147.095 63.535 147.505 ;
        RECT 63.705 146.745 63.995 147.910 ;
        RECT 64.165 147.885 64.380 147.935 ;
        RECT 64.165 147.805 64.555 147.885 ;
        RECT 64.225 146.960 64.555 147.805 ;
        RECT 65.065 147.850 65.255 148.055 ;
        RECT 64.725 146.745 64.895 147.755 ;
        RECT 65.065 147.475 65.960 147.850 ;
        RECT 65.065 146.915 65.405 147.475 ;
        RECT 65.635 146.745 65.950 147.245 ;
        RECT 66.130 147.215 66.300 148.055 ;
        RECT 66.470 148.345 66.935 148.675 ;
        RECT 67.320 148.615 67.490 148.845 ;
        RECT 67.670 148.795 68.040 149.295 ;
        RECT 68.360 148.845 69.035 149.015 ;
        RECT 69.230 148.845 69.565 149.015 ;
        RECT 66.470 147.385 66.790 148.345 ;
        RECT 67.320 148.315 68.150 148.615 ;
        RECT 66.960 147.415 67.150 148.135 ;
        RECT 67.320 147.245 67.490 148.315 ;
        RECT 67.950 148.285 68.150 148.315 ;
        RECT 67.660 148.065 67.830 148.135 ;
        RECT 68.360 148.065 68.530 148.845 ;
        RECT 69.395 148.705 69.565 148.845 ;
        RECT 69.735 148.835 69.985 149.295 ;
        RECT 67.660 147.895 68.530 148.065 ;
        RECT 68.700 148.425 69.225 148.645 ;
        RECT 69.395 148.575 69.620 148.705 ;
        RECT 67.660 147.805 68.170 147.895 ;
        RECT 66.130 147.045 67.015 147.215 ;
        RECT 67.240 146.915 67.490 147.245 ;
        RECT 67.660 146.745 67.830 147.545 ;
        RECT 68.000 147.190 68.170 147.805 ;
        RECT 68.700 147.725 68.870 148.425 ;
        RECT 68.340 147.360 68.870 147.725 ;
        RECT 69.040 147.660 69.280 148.255 ;
        RECT 69.450 147.470 69.620 148.575 ;
        RECT 69.790 147.715 70.070 148.665 ;
        RECT 69.315 147.340 69.620 147.470 ;
        RECT 68.000 147.020 69.105 147.190 ;
        RECT 69.315 146.915 69.565 147.340 ;
        RECT 69.735 146.745 70.000 147.205 ;
        RECT 70.240 146.915 70.425 149.035 ;
        RECT 70.595 148.915 70.925 149.295 ;
        RECT 71.095 148.745 71.265 149.035 ;
        RECT 70.600 148.575 71.265 148.745 ;
        RECT 70.600 147.585 70.830 148.575 ;
        RECT 71.530 148.555 71.785 149.125 ;
        RECT 71.955 148.895 72.285 149.295 ;
        RECT 72.710 148.760 73.240 149.125 ;
        RECT 73.430 148.955 73.705 149.125 ;
        RECT 73.425 148.785 73.705 148.955 ;
        RECT 72.710 148.725 72.885 148.760 ;
        RECT 71.955 148.555 72.885 148.725 ;
        RECT 71.000 147.755 71.350 148.405 ;
        RECT 71.530 147.885 71.700 148.555 ;
        RECT 71.955 148.385 72.125 148.555 ;
        RECT 71.870 148.055 72.125 148.385 ;
        RECT 72.350 148.055 72.545 148.385 ;
        RECT 70.600 147.415 71.265 147.585 ;
        RECT 70.595 146.745 70.925 147.245 ;
        RECT 71.095 146.915 71.265 147.415 ;
        RECT 71.530 146.915 71.865 147.885 ;
        RECT 72.035 146.745 72.205 147.885 ;
        RECT 72.375 147.085 72.545 148.055 ;
        RECT 72.715 147.425 72.885 148.555 ;
        RECT 73.055 147.765 73.225 148.565 ;
        RECT 73.430 147.965 73.705 148.785 ;
        RECT 73.875 147.765 74.065 149.125 ;
        RECT 74.245 148.760 74.755 149.295 ;
        RECT 74.975 148.485 75.220 149.090 ;
        RECT 75.665 148.555 76.050 149.125 ;
        RECT 76.220 148.835 76.545 149.295 ;
        RECT 77.065 148.665 77.345 149.125 ;
        RECT 74.265 148.315 75.495 148.485 ;
        RECT 73.055 147.595 74.065 147.765 ;
        RECT 74.235 147.750 74.985 147.940 ;
        RECT 72.715 147.255 73.840 147.425 ;
        RECT 74.235 147.085 74.405 147.750 ;
        RECT 75.155 147.505 75.495 148.315 ;
        RECT 72.375 146.915 74.405 147.085 ;
        RECT 74.575 146.745 74.745 147.505 ;
        RECT 74.980 147.095 75.495 147.505 ;
        RECT 75.665 147.885 75.945 148.555 ;
        RECT 76.220 148.495 77.345 148.665 ;
        RECT 76.220 148.385 76.670 148.495 ;
        RECT 76.115 148.055 76.670 148.385 ;
        RECT 77.535 148.325 77.935 149.125 ;
        RECT 78.335 148.835 78.605 149.295 ;
        RECT 78.775 148.665 79.060 149.125 ;
        RECT 75.665 146.915 76.050 147.885 ;
        RECT 76.220 147.595 76.670 148.055 ;
        RECT 76.840 147.765 77.935 148.325 ;
        RECT 76.220 147.375 77.345 147.595 ;
        RECT 76.220 146.745 76.545 147.205 ;
        RECT 77.065 146.915 77.345 147.375 ;
        RECT 77.535 146.915 77.935 147.765 ;
        RECT 78.105 148.495 79.060 148.665 ;
        RECT 79.345 148.555 79.730 149.125 ;
        RECT 79.900 148.835 80.225 149.295 ;
        RECT 80.745 148.665 81.025 149.125 ;
        RECT 78.105 147.595 78.315 148.495 ;
        RECT 78.485 147.765 79.175 148.325 ;
        RECT 79.345 147.885 79.625 148.555 ;
        RECT 79.900 148.495 81.025 148.665 ;
        RECT 79.900 148.385 80.350 148.495 ;
        RECT 79.795 148.055 80.350 148.385 ;
        RECT 81.215 148.325 81.615 149.125 ;
        RECT 82.015 148.835 82.285 149.295 ;
        RECT 82.455 148.665 82.740 149.125 ;
        RECT 78.105 147.375 79.060 147.595 ;
        RECT 78.335 146.745 78.605 147.205 ;
        RECT 78.775 146.915 79.060 147.375 ;
        RECT 79.345 146.915 79.730 147.885 ;
        RECT 79.900 147.595 80.350 148.055 ;
        RECT 80.520 147.765 81.615 148.325 ;
        RECT 79.900 147.375 81.025 147.595 ;
        RECT 79.900 146.745 80.225 147.205 ;
        RECT 80.745 146.915 81.025 147.375 ;
        RECT 81.215 146.915 81.615 147.765 ;
        RECT 81.785 148.495 82.740 148.665 ;
        RECT 83.025 148.495 83.365 149.125 ;
        RECT 83.535 148.495 83.785 149.295 ;
        RECT 83.975 148.645 84.305 149.125 ;
        RECT 84.475 148.835 84.700 149.295 ;
        RECT 84.870 148.645 85.200 149.125 ;
        RECT 81.785 147.595 81.995 148.495 ;
        RECT 82.165 147.765 82.855 148.325 ;
        RECT 83.025 147.885 83.200 148.495 ;
        RECT 83.975 148.475 85.200 148.645 ;
        RECT 85.830 148.515 86.330 149.125 ;
        RECT 86.795 148.745 86.965 149.125 ;
        RECT 87.180 148.915 87.510 149.295 ;
        RECT 86.795 148.575 87.510 148.745 ;
        RECT 83.370 148.135 84.065 148.305 ;
        RECT 83.895 147.885 84.065 148.135 ;
        RECT 84.240 148.105 84.660 148.305 ;
        RECT 84.830 148.105 85.160 148.305 ;
        RECT 85.330 148.105 85.660 148.305 ;
        RECT 85.830 147.885 86.000 148.515 ;
        RECT 86.185 148.055 86.535 148.305 ;
        RECT 86.705 148.025 87.060 148.395 ;
        RECT 87.340 148.385 87.510 148.575 ;
        RECT 87.680 148.550 87.935 149.125 ;
        RECT 87.340 148.055 87.595 148.385 ;
        RECT 81.785 147.375 82.740 147.595 ;
        RECT 82.015 146.745 82.285 147.205 ;
        RECT 82.455 146.915 82.740 147.375 ;
        RECT 83.025 146.915 83.365 147.885 ;
        RECT 83.535 146.745 83.705 147.885 ;
        RECT 83.895 147.715 86.330 147.885 ;
        RECT 87.340 147.845 87.510 148.055 ;
        RECT 83.975 146.745 84.225 147.545 ;
        RECT 84.870 146.915 85.200 147.715 ;
        RECT 85.500 146.745 85.830 147.545 ;
        RECT 86.000 146.915 86.330 147.715 ;
        RECT 86.795 147.675 87.510 147.845 ;
        RECT 87.765 147.820 87.935 148.550 ;
        RECT 88.110 148.455 88.370 149.295 ;
        RECT 88.545 148.545 89.755 149.295 ;
        RECT 86.795 146.915 86.965 147.675 ;
        RECT 87.180 146.745 87.510 147.505 ;
        RECT 87.680 146.915 87.935 147.820 ;
        RECT 88.110 146.745 88.370 147.895 ;
        RECT 88.545 147.835 89.065 148.375 ;
        RECT 89.235 148.005 89.755 148.545 ;
        RECT 101.840 148.320 102.010 149.730 ;
        RECT 102.380 149.160 105.420 149.330 ;
        RECT 102.380 148.720 105.420 148.890 ;
        RECT 105.635 148.860 105.805 149.190 ;
        RECT 106.140 148.970 118.590 149.730 ;
        RECT 121.720 149.730 138.470 149.900 ;
        RECT 146.140 149.850 158.550 149.900 ;
        RECT 106.140 148.960 118.480 148.970 ;
        RECT 106.140 148.950 112.020 148.960 ;
        RECT 106.140 148.930 106.710 148.950 ;
        RECT 107.930 148.940 112.020 148.950 ;
        RECT 106.150 148.320 106.320 148.930 ;
        RECT 101.840 148.150 106.320 148.320 ;
        RECT 121.720 148.320 121.890 149.730 ;
        RECT 122.260 149.160 125.300 149.330 ;
        RECT 122.260 148.720 125.300 148.890 ;
        RECT 125.515 148.860 125.685 149.190 ;
        RECT 126.020 148.970 138.470 149.730 ;
        RECT 141.800 149.680 158.550 149.850 ;
        RECT 126.020 148.960 138.360 148.970 ;
        RECT 126.020 148.950 131.900 148.960 ;
        RECT 126.020 148.930 126.590 148.950 ;
        RECT 127.810 148.940 131.900 148.950 ;
        RECT 126.030 148.320 126.200 148.930 ;
        RECT 121.720 148.150 126.200 148.320 ;
        RECT 141.800 148.270 141.970 149.680 ;
        RECT 142.340 149.110 145.380 149.280 ;
        RECT 142.340 148.670 145.380 148.840 ;
        RECT 145.595 148.810 145.765 149.140 ;
        RECT 146.100 148.920 158.550 149.680 ;
        RECT 146.100 148.910 158.440 148.920 ;
        RECT 146.100 148.900 151.980 148.910 ;
        RECT 146.100 148.880 146.670 148.900 ;
        RECT 147.890 148.890 151.980 148.900 ;
        RECT 146.110 148.270 146.280 148.880 ;
        RECT 141.800 148.100 146.280 148.270 ;
        RECT 88.545 146.745 89.755 147.835 ;
        RECT 12.100 146.575 89.840 146.745 ;
        RECT 100.630 146.740 106.370 146.750 ;
        RECT 100.140 146.580 106.370 146.740 ;
        RECT 12.185 145.485 13.395 146.575 ;
        RECT 13.565 145.485 16.155 146.575 ;
        RECT 16.875 145.905 17.045 146.405 ;
        RECT 17.215 146.075 17.545 146.575 ;
        RECT 16.875 145.735 17.540 145.905 ;
        RECT 12.185 144.775 12.705 145.315 ;
        RECT 12.875 144.945 13.395 145.485 ;
        RECT 13.565 144.795 14.775 145.315 ;
        RECT 14.945 144.965 16.155 145.485 ;
        RECT 16.790 144.915 17.140 145.565 ;
        RECT 12.185 144.025 13.395 144.775 ;
        RECT 13.565 144.025 16.155 144.795 ;
        RECT 17.310 144.745 17.540 145.735 ;
        RECT 16.875 144.575 17.540 144.745 ;
        RECT 16.875 144.285 17.045 144.575 ;
        RECT 17.215 144.025 17.545 144.405 ;
        RECT 17.715 144.285 17.900 146.405 ;
        RECT 18.140 146.115 18.405 146.575 ;
        RECT 18.575 145.980 18.825 146.405 ;
        RECT 19.035 146.130 20.140 146.300 ;
        RECT 18.520 145.850 18.825 145.980 ;
        RECT 18.070 144.655 18.350 145.605 ;
        RECT 18.520 144.745 18.690 145.850 ;
        RECT 18.860 145.065 19.100 145.660 ;
        RECT 19.270 145.595 19.800 145.960 ;
        RECT 19.270 144.895 19.440 145.595 ;
        RECT 19.970 145.515 20.140 146.130 ;
        RECT 20.310 145.775 20.480 146.575 ;
        RECT 20.650 146.075 20.900 146.405 ;
        RECT 21.125 146.105 22.010 146.275 ;
        RECT 19.970 145.425 20.480 145.515 ;
        RECT 18.520 144.615 18.745 144.745 ;
        RECT 18.915 144.675 19.440 144.895 ;
        RECT 19.610 145.255 20.480 145.425 ;
        RECT 18.155 144.025 18.405 144.485 ;
        RECT 18.575 144.475 18.745 144.615 ;
        RECT 19.610 144.475 19.780 145.255 ;
        RECT 20.310 145.185 20.480 145.255 ;
        RECT 19.990 145.005 20.190 145.035 ;
        RECT 20.650 145.005 20.820 146.075 ;
        RECT 20.990 145.185 21.180 145.905 ;
        RECT 19.990 144.705 20.820 145.005 ;
        RECT 21.350 144.975 21.670 145.935 ;
        RECT 18.575 144.305 18.910 144.475 ;
        RECT 19.105 144.305 19.780 144.475 ;
        RECT 20.100 144.025 20.470 144.525 ;
        RECT 20.650 144.475 20.820 144.705 ;
        RECT 21.205 144.645 21.670 144.975 ;
        RECT 21.840 145.265 22.010 146.105 ;
        RECT 22.190 146.075 22.505 146.575 ;
        RECT 22.735 145.845 23.075 146.405 ;
        RECT 22.180 145.470 23.075 145.845 ;
        RECT 23.245 145.565 23.415 146.575 ;
        RECT 22.885 145.265 23.075 145.470 ;
        RECT 23.585 145.515 23.915 146.360 ;
        RECT 23.585 145.435 23.975 145.515 ;
        RECT 23.760 145.385 23.975 145.435 ;
        RECT 25.065 145.410 25.355 146.575 ;
        RECT 25.535 145.605 25.865 146.390 ;
        RECT 25.535 145.435 26.215 145.605 ;
        RECT 26.395 145.435 26.725 146.575 ;
        RECT 26.995 145.905 27.165 146.405 ;
        RECT 27.335 146.075 27.665 146.575 ;
        RECT 26.995 145.735 27.660 145.905 ;
        RECT 21.840 144.935 22.715 145.265 ;
        RECT 22.885 144.935 23.635 145.265 ;
        RECT 21.840 144.475 22.010 144.935 ;
        RECT 22.885 144.765 23.085 144.935 ;
        RECT 23.805 144.805 23.975 145.385 ;
        RECT 25.525 145.015 25.875 145.265 ;
        RECT 26.045 144.835 26.215 145.435 ;
        RECT 26.385 145.015 26.735 145.265 ;
        RECT 26.910 144.915 27.260 145.565 ;
        RECT 23.750 144.765 23.975 144.805 ;
        RECT 20.650 144.305 21.055 144.475 ;
        RECT 21.225 144.305 22.010 144.475 ;
        RECT 22.285 144.025 22.495 144.555 ;
        RECT 22.755 144.240 23.085 144.765 ;
        RECT 23.595 144.680 23.975 144.765 ;
        RECT 23.255 144.025 23.425 144.635 ;
        RECT 23.595 144.245 23.925 144.680 ;
        RECT 25.065 144.025 25.355 144.750 ;
        RECT 25.545 144.025 25.785 144.835 ;
        RECT 25.955 144.195 26.285 144.835 ;
        RECT 26.455 144.025 26.725 144.835 ;
        RECT 27.430 144.745 27.660 145.735 ;
        RECT 26.995 144.575 27.660 144.745 ;
        RECT 26.995 144.285 27.165 144.575 ;
        RECT 27.335 144.025 27.665 144.405 ;
        RECT 27.835 144.285 28.020 146.405 ;
        RECT 28.260 146.115 28.525 146.575 ;
        RECT 28.695 145.980 28.945 146.405 ;
        RECT 29.155 146.130 30.260 146.300 ;
        RECT 28.640 145.850 28.945 145.980 ;
        RECT 28.190 144.655 28.470 145.605 ;
        RECT 28.640 144.745 28.810 145.850 ;
        RECT 28.980 145.065 29.220 145.660 ;
        RECT 29.390 145.595 29.920 145.960 ;
        RECT 29.390 144.895 29.560 145.595 ;
        RECT 30.090 145.515 30.260 146.130 ;
        RECT 30.430 145.775 30.600 146.575 ;
        RECT 30.770 146.075 31.020 146.405 ;
        RECT 31.245 146.105 32.130 146.275 ;
        RECT 30.090 145.425 30.600 145.515 ;
        RECT 28.640 144.615 28.865 144.745 ;
        RECT 29.035 144.675 29.560 144.895 ;
        RECT 29.730 145.255 30.600 145.425 ;
        RECT 28.275 144.025 28.525 144.485 ;
        RECT 28.695 144.475 28.865 144.615 ;
        RECT 29.730 144.475 29.900 145.255 ;
        RECT 30.430 145.185 30.600 145.255 ;
        RECT 30.110 145.005 30.310 145.035 ;
        RECT 30.770 145.005 30.940 146.075 ;
        RECT 31.110 145.185 31.300 145.905 ;
        RECT 30.110 144.705 30.940 145.005 ;
        RECT 31.470 144.975 31.790 145.935 ;
        RECT 28.695 144.305 29.030 144.475 ;
        RECT 29.225 144.305 29.900 144.475 ;
        RECT 30.220 144.025 30.590 144.525 ;
        RECT 30.770 144.475 30.940 144.705 ;
        RECT 31.325 144.645 31.790 144.975 ;
        RECT 31.960 145.265 32.130 146.105 ;
        RECT 32.310 146.075 32.625 146.575 ;
        RECT 32.855 145.845 33.195 146.405 ;
        RECT 32.300 145.470 33.195 145.845 ;
        RECT 33.365 145.565 33.535 146.575 ;
        RECT 33.005 145.265 33.195 145.470 ;
        RECT 33.705 145.515 34.035 146.360 ;
        RECT 34.355 145.905 34.525 146.405 ;
        RECT 34.695 146.075 35.025 146.575 ;
        RECT 34.355 145.735 35.020 145.905 ;
        RECT 33.705 145.435 34.095 145.515 ;
        RECT 33.880 145.385 34.095 145.435 ;
        RECT 31.960 144.935 32.835 145.265 ;
        RECT 33.005 144.935 33.755 145.265 ;
        RECT 31.960 144.475 32.130 144.935 ;
        RECT 33.005 144.765 33.205 144.935 ;
        RECT 33.925 144.805 34.095 145.385 ;
        RECT 34.270 144.915 34.620 145.565 ;
        RECT 33.870 144.765 34.095 144.805 ;
        RECT 30.770 144.305 31.175 144.475 ;
        RECT 31.345 144.305 32.130 144.475 ;
        RECT 32.405 144.025 32.615 144.555 ;
        RECT 32.875 144.240 33.205 144.765 ;
        RECT 33.715 144.680 34.095 144.765 ;
        RECT 34.790 144.745 35.020 145.735 ;
        RECT 33.375 144.025 33.545 144.635 ;
        RECT 33.715 144.245 34.045 144.680 ;
        RECT 34.355 144.575 35.020 144.745 ;
        RECT 34.355 144.285 34.525 144.575 ;
        RECT 34.695 144.025 35.025 144.405 ;
        RECT 35.195 144.285 35.380 146.405 ;
        RECT 35.620 146.115 35.885 146.575 ;
        RECT 36.055 145.980 36.305 146.405 ;
        RECT 36.515 146.130 37.620 146.300 ;
        RECT 36.000 145.850 36.305 145.980 ;
        RECT 35.550 144.655 35.830 145.605 ;
        RECT 36.000 144.745 36.170 145.850 ;
        RECT 36.340 145.065 36.580 145.660 ;
        RECT 36.750 145.595 37.280 145.960 ;
        RECT 36.750 144.895 36.920 145.595 ;
        RECT 37.450 145.515 37.620 146.130 ;
        RECT 37.790 145.775 37.960 146.575 ;
        RECT 38.130 146.075 38.380 146.405 ;
        RECT 38.605 146.105 39.490 146.275 ;
        RECT 37.450 145.425 37.960 145.515 ;
        RECT 36.000 144.615 36.225 144.745 ;
        RECT 36.395 144.675 36.920 144.895 ;
        RECT 37.090 145.255 37.960 145.425 ;
        RECT 35.635 144.025 35.885 144.485 ;
        RECT 36.055 144.475 36.225 144.615 ;
        RECT 37.090 144.475 37.260 145.255 ;
        RECT 37.790 145.185 37.960 145.255 ;
        RECT 37.470 145.005 37.670 145.035 ;
        RECT 38.130 145.005 38.300 146.075 ;
        RECT 38.470 145.185 38.660 145.905 ;
        RECT 37.470 144.705 38.300 145.005 ;
        RECT 38.830 144.975 39.150 145.935 ;
        RECT 36.055 144.305 36.390 144.475 ;
        RECT 36.585 144.305 37.260 144.475 ;
        RECT 37.580 144.025 37.950 144.525 ;
        RECT 38.130 144.475 38.300 144.705 ;
        RECT 38.685 144.645 39.150 144.975 ;
        RECT 39.320 145.265 39.490 146.105 ;
        RECT 39.670 146.075 39.985 146.575 ;
        RECT 40.215 145.845 40.555 146.405 ;
        RECT 39.660 145.470 40.555 145.845 ;
        RECT 40.725 145.565 40.895 146.575 ;
        RECT 40.365 145.265 40.555 145.470 ;
        RECT 41.065 145.515 41.395 146.360 ;
        RECT 41.065 145.435 41.455 145.515 ;
        RECT 41.240 145.385 41.455 145.435 ;
        RECT 39.320 144.935 40.195 145.265 ;
        RECT 40.365 144.935 41.115 145.265 ;
        RECT 39.320 144.475 39.490 144.935 ;
        RECT 40.365 144.765 40.565 144.935 ;
        RECT 41.285 144.805 41.455 145.385 ;
        RECT 41.230 144.765 41.455 144.805 ;
        RECT 38.130 144.305 38.535 144.475 ;
        RECT 38.705 144.305 39.490 144.475 ;
        RECT 39.765 144.025 39.975 144.555 ;
        RECT 40.235 144.240 40.565 144.765 ;
        RECT 41.075 144.680 41.455 144.765 ;
        RECT 41.625 145.435 42.010 146.405 ;
        RECT 42.180 146.115 42.505 146.575 ;
        RECT 43.025 145.945 43.305 146.405 ;
        RECT 42.180 145.725 43.305 145.945 ;
        RECT 41.625 144.765 41.905 145.435 ;
        RECT 42.180 145.265 42.630 145.725 ;
        RECT 43.495 145.555 43.895 146.405 ;
        RECT 44.295 146.115 44.565 146.575 ;
        RECT 44.735 145.945 45.020 146.405 ;
        RECT 42.075 144.935 42.630 145.265 ;
        RECT 42.800 144.995 43.895 145.555 ;
        RECT 42.180 144.825 42.630 144.935 ;
        RECT 40.735 144.025 40.905 144.635 ;
        RECT 41.075 144.245 41.405 144.680 ;
        RECT 41.625 144.195 42.010 144.765 ;
        RECT 42.180 144.655 43.305 144.825 ;
        RECT 42.180 144.025 42.505 144.485 ;
        RECT 43.025 144.195 43.305 144.655 ;
        RECT 43.495 144.195 43.895 144.995 ;
        RECT 44.065 145.725 45.020 145.945 ;
        RECT 44.065 144.825 44.275 145.725 ;
        RECT 44.445 144.995 45.135 145.555 ;
        RECT 45.305 145.485 46.975 146.575 ;
        RECT 44.065 144.655 45.020 144.825 ;
        RECT 44.295 144.025 44.565 144.485 ;
        RECT 44.735 144.195 45.020 144.655 ;
        RECT 45.305 144.795 46.055 145.315 ;
        RECT 46.225 144.965 46.975 145.485 ;
        RECT 47.145 145.435 47.530 146.405 ;
        RECT 47.700 146.115 48.025 146.575 ;
        RECT 48.545 145.945 48.825 146.405 ;
        RECT 47.700 145.725 48.825 145.945 ;
        RECT 45.305 144.025 46.975 144.795 ;
        RECT 47.145 144.765 47.425 145.435 ;
        RECT 47.700 145.265 48.150 145.725 ;
        RECT 49.015 145.555 49.415 146.405 ;
        RECT 49.815 146.115 50.085 146.575 ;
        RECT 50.255 145.945 50.540 146.405 ;
        RECT 47.595 144.935 48.150 145.265 ;
        RECT 48.320 144.995 49.415 145.555 ;
        RECT 47.700 144.825 48.150 144.935 ;
        RECT 47.145 144.195 47.530 144.765 ;
        RECT 47.700 144.655 48.825 144.825 ;
        RECT 47.700 144.025 48.025 144.485 ;
        RECT 48.545 144.195 48.825 144.655 ;
        RECT 49.015 144.195 49.415 144.995 ;
        RECT 49.585 145.725 50.540 145.945 ;
        RECT 49.585 144.825 49.795 145.725 ;
        RECT 49.965 144.995 50.655 145.555 ;
        RECT 50.825 145.410 51.115 146.575 ;
        RECT 51.295 145.605 51.625 146.390 ;
        RECT 51.295 145.435 51.975 145.605 ;
        RECT 52.155 145.435 52.485 146.575 ;
        RECT 52.665 145.485 54.335 146.575 ;
        RECT 54.595 145.905 54.765 146.405 ;
        RECT 54.935 146.075 55.265 146.575 ;
        RECT 54.595 145.735 55.260 145.905 ;
        RECT 51.285 145.015 51.635 145.265 ;
        RECT 51.805 144.835 51.975 145.435 ;
        RECT 52.145 145.015 52.495 145.265 ;
        RECT 49.585 144.655 50.540 144.825 ;
        RECT 49.815 144.025 50.085 144.485 ;
        RECT 50.255 144.195 50.540 144.655 ;
        RECT 50.825 144.025 51.115 144.750 ;
        RECT 51.305 144.025 51.545 144.835 ;
        RECT 51.715 144.195 52.045 144.835 ;
        RECT 52.215 144.025 52.485 144.835 ;
        RECT 52.665 144.795 53.415 145.315 ;
        RECT 53.585 144.965 54.335 145.485 ;
        RECT 54.510 144.915 54.860 145.565 ;
        RECT 52.665 144.025 54.335 144.795 ;
        RECT 55.030 144.745 55.260 145.735 ;
        RECT 54.595 144.575 55.260 144.745 ;
        RECT 54.595 144.285 54.765 144.575 ;
        RECT 54.935 144.025 55.265 144.405 ;
        RECT 55.435 144.285 55.620 146.405 ;
        RECT 55.860 146.115 56.125 146.575 ;
        RECT 56.295 145.980 56.545 146.405 ;
        RECT 56.755 146.130 57.860 146.300 ;
        RECT 56.240 145.850 56.545 145.980 ;
        RECT 55.790 144.655 56.070 145.605 ;
        RECT 56.240 144.745 56.410 145.850 ;
        RECT 56.580 145.065 56.820 145.660 ;
        RECT 56.990 145.595 57.520 145.960 ;
        RECT 56.990 144.895 57.160 145.595 ;
        RECT 57.690 145.515 57.860 146.130 ;
        RECT 58.030 145.775 58.200 146.575 ;
        RECT 58.370 146.075 58.620 146.405 ;
        RECT 58.845 146.105 59.730 146.275 ;
        RECT 57.690 145.425 58.200 145.515 ;
        RECT 56.240 144.615 56.465 144.745 ;
        RECT 56.635 144.675 57.160 144.895 ;
        RECT 57.330 145.255 58.200 145.425 ;
        RECT 55.875 144.025 56.125 144.485 ;
        RECT 56.295 144.475 56.465 144.615 ;
        RECT 57.330 144.475 57.500 145.255 ;
        RECT 58.030 145.185 58.200 145.255 ;
        RECT 57.710 145.005 57.910 145.035 ;
        RECT 58.370 145.005 58.540 146.075 ;
        RECT 58.710 145.185 58.900 145.905 ;
        RECT 57.710 144.705 58.540 145.005 ;
        RECT 59.070 144.975 59.390 145.935 ;
        RECT 56.295 144.305 56.630 144.475 ;
        RECT 56.825 144.305 57.500 144.475 ;
        RECT 57.820 144.025 58.190 144.525 ;
        RECT 58.370 144.475 58.540 144.705 ;
        RECT 58.925 144.645 59.390 144.975 ;
        RECT 59.560 145.265 59.730 146.105 ;
        RECT 59.910 146.075 60.225 146.575 ;
        RECT 60.455 145.845 60.795 146.405 ;
        RECT 59.900 145.470 60.795 145.845 ;
        RECT 60.965 145.565 61.135 146.575 ;
        RECT 60.605 145.265 60.795 145.470 ;
        RECT 61.305 145.515 61.635 146.360 ;
        RECT 61.305 145.435 61.695 145.515 ;
        RECT 61.480 145.385 61.695 145.435 ;
        RECT 62.330 145.425 62.590 146.575 ;
        RECT 62.765 145.500 63.020 146.405 ;
        RECT 63.190 145.815 63.520 146.575 ;
        RECT 63.735 145.645 63.905 146.405 ;
        RECT 59.560 144.935 60.435 145.265 ;
        RECT 60.605 144.935 61.355 145.265 ;
        RECT 59.560 144.475 59.730 144.935 ;
        RECT 60.605 144.765 60.805 144.935 ;
        RECT 61.525 144.805 61.695 145.385 ;
        RECT 61.470 144.765 61.695 144.805 ;
        RECT 58.370 144.305 58.775 144.475 ;
        RECT 58.945 144.305 59.730 144.475 ;
        RECT 60.005 144.025 60.215 144.555 ;
        RECT 60.475 144.240 60.805 144.765 ;
        RECT 61.315 144.680 61.695 144.765 ;
        RECT 60.975 144.025 61.145 144.635 ;
        RECT 61.315 144.245 61.645 144.680 ;
        RECT 62.330 144.025 62.590 144.865 ;
        RECT 62.765 144.770 62.935 145.500 ;
        RECT 63.190 145.475 63.905 145.645 ;
        RECT 64.165 145.815 64.680 146.225 ;
        RECT 64.915 145.815 65.085 146.575 ;
        RECT 65.255 146.235 67.285 146.405 ;
        RECT 63.190 145.265 63.360 145.475 ;
        RECT 63.105 144.935 63.360 145.265 ;
        RECT 62.765 144.195 63.020 144.770 ;
        RECT 63.190 144.745 63.360 144.935 ;
        RECT 63.640 144.925 63.995 145.295 ;
        RECT 64.165 145.005 64.505 145.815 ;
        RECT 65.255 145.570 65.425 146.235 ;
        RECT 65.820 145.895 66.945 146.065 ;
        RECT 64.675 145.380 65.425 145.570 ;
        RECT 65.595 145.555 66.605 145.725 ;
        RECT 64.165 144.835 65.395 145.005 ;
        RECT 63.190 144.575 63.905 144.745 ;
        RECT 63.190 144.025 63.520 144.405 ;
        RECT 63.735 144.195 63.905 144.575 ;
        RECT 64.440 144.230 64.685 144.835 ;
        RECT 64.905 144.025 65.415 144.560 ;
        RECT 65.595 144.195 65.785 145.555 ;
        RECT 65.955 144.535 66.230 145.355 ;
        RECT 66.435 144.755 66.605 145.555 ;
        RECT 66.775 144.765 66.945 145.895 ;
        RECT 67.115 145.265 67.285 146.235 ;
        RECT 67.455 145.435 67.625 146.575 ;
        RECT 67.795 145.435 68.130 146.405 ;
        RECT 67.115 144.935 67.310 145.265 ;
        RECT 67.535 144.935 67.790 145.265 ;
        RECT 67.535 144.765 67.705 144.935 ;
        RECT 67.960 144.765 68.130 145.435 ;
        RECT 66.775 144.595 67.705 144.765 ;
        RECT 66.775 144.560 66.950 144.595 ;
        RECT 65.955 144.365 66.235 144.535 ;
        RECT 65.955 144.195 66.230 144.365 ;
        RECT 66.420 144.195 66.950 144.560 ;
        RECT 67.375 144.025 67.705 144.425 ;
        RECT 67.875 144.195 68.130 144.765 ;
        RECT 68.310 145.435 68.645 146.405 ;
        RECT 68.815 145.435 68.985 146.575 ;
        RECT 69.155 146.235 71.185 146.405 ;
        RECT 68.310 144.765 68.480 145.435 ;
        RECT 69.155 145.265 69.325 146.235 ;
        RECT 68.650 144.935 68.905 145.265 ;
        RECT 69.130 144.935 69.325 145.265 ;
        RECT 69.495 145.895 70.620 146.065 ;
        RECT 68.735 144.765 68.905 144.935 ;
        RECT 69.495 144.765 69.665 145.895 ;
        RECT 68.310 144.195 68.565 144.765 ;
        RECT 68.735 144.595 69.665 144.765 ;
        RECT 69.835 145.555 70.845 145.725 ;
        RECT 69.835 144.755 70.005 145.555 ;
        RECT 70.210 144.875 70.485 145.355 ;
        RECT 70.205 144.705 70.485 144.875 ;
        RECT 69.490 144.560 69.665 144.595 ;
        RECT 68.735 144.025 69.065 144.425 ;
        RECT 69.490 144.195 70.020 144.560 ;
        RECT 70.210 144.195 70.485 144.705 ;
        RECT 70.655 144.195 70.845 145.555 ;
        RECT 71.015 145.570 71.185 146.235 ;
        RECT 71.355 145.815 71.525 146.575 ;
        RECT 71.760 145.815 72.275 146.225 ;
        RECT 71.015 145.380 71.765 145.570 ;
        RECT 71.935 145.005 72.275 145.815 ;
        RECT 71.045 144.835 72.275 145.005 ;
        RECT 72.450 145.435 72.785 146.405 ;
        RECT 72.955 145.435 73.125 146.575 ;
        RECT 73.295 146.235 75.325 146.405 ;
        RECT 71.025 144.025 71.535 144.560 ;
        RECT 71.755 144.230 72.000 144.835 ;
        RECT 72.450 144.765 72.620 145.435 ;
        RECT 73.295 145.265 73.465 146.235 ;
        RECT 72.790 144.935 73.045 145.265 ;
        RECT 73.270 144.935 73.465 145.265 ;
        RECT 73.635 145.895 74.760 146.065 ;
        RECT 72.875 144.765 73.045 144.935 ;
        RECT 73.635 144.765 73.805 145.895 ;
        RECT 72.450 144.195 72.705 144.765 ;
        RECT 72.875 144.595 73.805 144.765 ;
        RECT 73.975 145.555 74.985 145.725 ;
        RECT 73.975 144.755 74.145 145.555 ;
        RECT 74.350 145.215 74.625 145.355 ;
        RECT 74.345 145.045 74.625 145.215 ;
        RECT 73.630 144.560 73.805 144.595 ;
        RECT 72.875 144.025 73.205 144.425 ;
        RECT 73.630 144.195 74.160 144.560 ;
        RECT 74.350 144.195 74.625 145.045 ;
        RECT 74.795 144.195 74.985 145.555 ;
        RECT 75.155 145.570 75.325 146.235 ;
        RECT 75.495 145.815 75.665 146.575 ;
        RECT 75.900 145.815 76.415 146.225 ;
        RECT 75.155 145.380 75.905 145.570 ;
        RECT 76.075 145.005 76.415 145.815 ;
        RECT 76.585 145.410 76.875 146.575 ;
        RECT 77.135 145.905 77.305 146.405 ;
        RECT 77.475 146.075 77.805 146.575 ;
        RECT 77.135 145.735 77.800 145.905 ;
        RECT 75.185 144.835 76.415 145.005 ;
        RECT 77.050 144.915 77.400 145.565 ;
        RECT 75.165 144.025 75.675 144.560 ;
        RECT 75.895 144.230 76.140 144.835 ;
        RECT 76.585 144.025 76.875 144.750 ;
        RECT 77.570 144.745 77.800 145.735 ;
        RECT 77.135 144.575 77.800 144.745 ;
        RECT 77.135 144.285 77.305 144.575 ;
        RECT 77.475 144.025 77.805 144.405 ;
        RECT 77.975 144.285 78.160 146.405 ;
        RECT 78.400 146.115 78.665 146.575 ;
        RECT 78.835 145.980 79.085 146.405 ;
        RECT 79.295 146.130 80.400 146.300 ;
        RECT 78.780 145.850 79.085 145.980 ;
        RECT 78.330 144.655 78.610 145.605 ;
        RECT 78.780 144.745 78.950 145.850 ;
        RECT 79.120 145.065 79.360 145.660 ;
        RECT 79.530 145.595 80.060 145.960 ;
        RECT 79.530 144.895 79.700 145.595 ;
        RECT 80.230 145.515 80.400 146.130 ;
        RECT 80.570 145.775 80.740 146.575 ;
        RECT 80.910 146.075 81.160 146.405 ;
        RECT 81.385 146.105 82.270 146.275 ;
        RECT 80.230 145.425 80.740 145.515 ;
        RECT 78.780 144.615 79.005 144.745 ;
        RECT 79.175 144.675 79.700 144.895 ;
        RECT 79.870 145.255 80.740 145.425 ;
        RECT 78.415 144.025 78.665 144.485 ;
        RECT 78.835 144.475 79.005 144.615 ;
        RECT 79.870 144.475 80.040 145.255 ;
        RECT 80.570 145.185 80.740 145.255 ;
        RECT 80.250 145.005 80.450 145.035 ;
        RECT 80.910 145.005 81.080 146.075 ;
        RECT 81.250 145.185 81.440 145.905 ;
        RECT 80.250 144.705 81.080 145.005 ;
        RECT 81.610 144.975 81.930 145.935 ;
        RECT 78.835 144.305 79.170 144.475 ;
        RECT 79.365 144.305 80.040 144.475 ;
        RECT 80.360 144.025 80.730 144.525 ;
        RECT 80.910 144.475 81.080 144.705 ;
        RECT 81.465 144.645 81.930 144.975 ;
        RECT 82.100 145.265 82.270 146.105 ;
        RECT 82.450 146.075 82.765 146.575 ;
        RECT 82.995 145.845 83.335 146.405 ;
        RECT 82.440 145.470 83.335 145.845 ;
        RECT 83.505 145.565 83.675 146.575 ;
        RECT 83.145 145.265 83.335 145.470 ;
        RECT 83.845 145.515 84.175 146.360 ;
        RECT 83.845 145.435 84.235 145.515 ;
        RECT 84.020 145.385 84.235 145.435 ;
        RECT 82.100 144.935 82.975 145.265 ;
        RECT 83.145 144.935 83.895 145.265 ;
        RECT 82.100 144.475 82.270 144.935 ;
        RECT 83.145 144.765 83.345 144.935 ;
        RECT 84.065 144.805 84.235 145.385 ;
        RECT 84.010 144.765 84.235 144.805 ;
        RECT 80.910 144.305 81.315 144.475 ;
        RECT 81.485 144.305 82.270 144.475 ;
        RECT 82.545 144.025 82.755 144.555 ;
        RECT 83.015 144.240 83.345 144.765 ;
        RECT 83.855 144.680 84.235 144.765 ;
        RECT 84.405 145.435 84.745 146.405 ;
        RECT 84.915 145.435 85.085 146.575 ;
        RECT 85.355 145.775 85.605 146.575 ;
        RECT 86.250 145.605 86.580 146.405 ;
        RECT 86.880 145.775 87.210 146.575 ;
        RECT 87.380 145.605 87.710 146.405 ;
        RECT 85.275 145.435 87.710 145.605 ;
        RECT 88.545 145.485 89.755 146.575 ;
        RECT 84.405 144.825 84.580 145.435 ;
        RECT 85.275 145.185 85.445 145.435 ;
        RECT 84.750 145.015 85.445 145.185 ;
        RECT 85.620 145.015 86.040 145.215 ;
        RECT 86.210 145.015 86.540 145.215 ;
        RECT 86.710 145.015 87.040 145.215 ;
        RECT 83.515 144.025 83.685 144.635 ;
        RECT 83.855 144.245 84.185 144.680 ;
        RECT 84.405 144.195 84.745 144.825 ;
        RECT 84.915 144.025 85.165 144.825 ;
        RECT 85.355 144.675 86.580 144.845 ;
        RECT 85.355 144.195 85.685 144.675 ;
        RECT 85.855 144.025 86.080 144.485 ;
        RECT 86.250 144.195 86.580 144.675 ;
        RECT 87.210 144.805 87.380 145.435 ;
        RECT 87.565 145.015 87.915 145.265 ;
        RECT 88.545 144.945 89.065 145.485 ;
        RECT 87.210 144.195 87.710 144.805 ;
        RECT 89.235 144.775 89.755 145.315 ;
        RECT 88.545 144.025 89.755 144.775 ;
        RECT 100.140 144.320 100.810 146.580 ;
        RECT 101.480 146.010 105.520 146.180 ;
        RECT 101.140 144.950 101.310 145.950 ;
        RECT 105.690 144.950 105.860 145.950 ;
        RECT 101.480 144.720 105.520 144.890 ;
        RECT 106.200 144.320 106.370 146.580 ;
        RECT 100.140 144.150 106.370 144.320 ;
        RECT 12.100 143.855 89.840 144.025 ;
        RECT 12.185 143.105 13.395 143.855 ;
        RECT 12.185 142.565 12.705 143.105 ;
        RECT 14.035 143.045 14.305 143.855 ;
        RECT 14.475 143.045 14.805 143.685 ;
        RECT 14.975 143.045 15.215 143.855 ;
        RECT 15.490 143.285 15.665 143.685 ;
        RECT 15.835 143.475 16.165 143.855 ;
        RECT 16.410 143.355 16.640 143.685 ;
        RECT 15.490 143.115 16.120 143.285 ;
        RECT 12.875 142.395 13.395 142.935 ;
        RECT 14.025 142.615 14.375 142.865 ;
        RECT 14.545 142.445 14.715 143.045 ;
        RECT 15.950 142.945 16.120 143.115 ;
        RECT 14.885 142.615 15.235 142.865 ;
        RECT 12.185 141.305 13.395 142.395 ;
        RECT 14.035 141.305 14.365 142.445 ;
        RECT 14.545 142.275 15.225 142.445 ;
        RECT 14.895 141.490 15.225 142.275 ;
        RECT 15.405 142.265 15.770 142.945 ;
        RECT 15.950 142.615 16.300 142.945 ;
        RECT 15.950 142.095 16.120 142.615 ;
        RECT 15.490 141.925 16.120 142.095 ;
        RECT 16.470 142.065 16.640 143.355 ;
        RECT 16.840 142.245 17.120 143.520 ;
        RECT 17.345 143.515 17.615 143.520 ;
        RECT 17.305 143.345 17.615 143.515 ;
        RECT 18.075 143.475 18.405 143.855 ;
        RECT 18.575 143.600 18.910 143.645 ;
        RECT 17.345 142.245 17.615 143.345 ;
        RECT 17.805 142.245 18.145 143.275 ;
        RECT 18.575 143.135 18.915 143.600 ;
        RECT 18.315 142.615 18.575 142.945 ;
        RECT 18.315 142.065 18.485 142.615 ;
        RECT 18.745 142.445 18.915 143.135 ;
        RECT 19.170 143.285 19.345 143.685 ;
        RECT 19.515 143.475 19.845 143.855 ;
        RECT 20.090 143.355 20.320 143.685 ;
        RECT 19.170 143.115 19.800 143.285 ;
        RECT 19.630 142.945 19.800 143.115 ;
        RECT 15.490 141.475 15.665 141.925 ;
        RECT 16.470 141.895 18.485 142.065 ;
        RECT 15.835 141.305 16.165 141.745 ;
        RECT 16.470 141.475 16.640 141.895 ;
        RECT 16.875 141.305 17.545 141.715 ;
        RECT 17.760 141.475 17.930 141.895 ;
        RECT 18.130 141.305 18.460 141.715 ;
        RECT 18.655 141.475 18.915 142.445 ;
        RECT 19.085 142.265 19.450 142.945 ;
        RECT 19.630 142.615 19.980 142.945 ;
        RECT 19.630 142.095 19.800 142.615 ;
        RECT 19.170 141.925 19.800 142.095 ;
        RECT 20.150 142.065 20.320 143.355 ;
        RECT 20.520 142.245 20.800 143.520 ;
        RECT 21.025 143.515 21.295 143.520 ;
        RECT 20.985 143.345 21.295 143.515 ;
        RECT 21.755 143.475 22.085 143.855 ;
        RECT 22.255 143.600 22.590 143.645 ;
        RECT 21.025 142.245 21.295 143.345 ;
        RECT 21.485 142.245 21.825 143.275 ;
        RECT 22.255 143.135 22.595 143.600 ;
        RECT 22.855 143.305 23.025 143.595 ;
        RECT 23.195 143.475 23.525 143.855 ;
        RECT 22.855 143.135 23.520 143.305 ;
        RECT 21.995 142.615 22.255 142.945 ;
        RECT 21.995 142.065 22.165 142.615 ;
        RECT 22.425 142.445 22.595 143.135 ;
        RECT 19.170 141.475 19.345 141.925 ;
        RECT 20.150 141.895 22.165 142.065 ;
        RECT 19.515 141.305 19.845 141.745 ;
        RECT 20.150 141.475 20.320 141.895 ;
        RECT 20.555 141.305 21.225 141.715 ;
        RECT 21.440 141.475 21.610 141.895 ;
        RECT 21.810 141.305 22.140 141.715 ;
        RECT 22.335 141.475 22.595 142.445 ;
        RECT 22.770 142.315 23.120 142.965 ;
        RECT 23.290 142.145 23.520 143.135 ;
        RECT 22.855 141.975 23.520 142.145 ;
        RECT 22.855 141.475 23.025 141.975 ;
        RECT 23.195 141.305 23.525 141.805 ;
        RECT 23.695 141.475 23.880 143.595 ;
        RECT 24.135 143.395 24.385 143.855 ;
        RECT 24.555 143.405 24.890 143.575 ;
        RECT 25.085 143.405 25.760 143.575 ;
        RECT 24.555 143.265 24.725 143.405 ;
        RECT 24.050 142.275 24.330 143.225 ;
        RECT 24.500 143.135 24.725 143.265 ;
        RECT 24.500 142.030 24.670 143.135 ;
        RECT 24.895 142.985 25.420 143.205 ;
        RECT 24.840 142.220 25.080 142.815 ;
        RECT 25.250 142.285 25.420 142.985 ;
        RECT 25.590 142.625 25.760 143.405 ;
        RECT 26.080 143.355 26.450 143.855 ;
        RECT 26.630 143.405 27.035 143.575 ;
        RECT 27.205 143.405 27.990 143.575 ;
        RECT 26.630 143.175 26.800 143.405 ;
        RECT 25.970 142.875 26.800 143.175 ;
        RECT 27.185 142.905 27.650 143.235 ;
        RECT 25.970 142.845 26.170 142.875 ;
        RECT 26.290 142.625 26.460 142.695 ;
        RECT 25.590 142.455 26.460 142.625 ;
        RECT 25.950 142.365 26.460 142.455 ;
        RECT 24.500 141.900 24.805 142.030 ;
        RECT 25.250 141.920 25.780 142.285 ;
        RECT 24.120 141.305 24.385 141.765 ;
        RECT 24.555 141.475 24.805 141.900 ;
        RECT 25.950 141.750 26.120 142.365 ;
        RECT 25.015 141.580 26.120 141.750 ;
        RECT 26.290 141.305 26.460 142.105 ;
        RECT 26.630 141.805 26.800 142.875 ;
        RECT 26.970 141.975 27.160 142.695 ;
        RECT 27.330 141.945 27.650 142.905 ;
        RECT 27.820 142.945 27.990 143.405 ;
        RECT 28.265 143.325 28.475 143.855 ;
        RECT 28.735 143.115 29.065 143.640 ;
        RECT 29.235 143.245 29.405 143.855 ;
        RECT 29.575 143.200 29.905 143.635 ;
        RECT 30.215 143.305 30.385 143.595 ;
        RECT 30.555 143.475 30.885 143.855 ;
        RECT 29.575 143.115 29.955 143.200 ;
        RECT 30.215 143.135 30.880 143.305 ;
        RECT 28.865 142.945 29.065 143.115 ;
        RECT 29.730 143.075 29.955 143.115 ;
        RECT 27.820 142.615 28.695 142.945 ;
        RECT 28.865 142.615 29.615 142.945 ;
        RECT 26.630 141.475 26.880 141.805 ;
        RECT 27.820 141.775 27.990 142.615 ;
        RECT 28.865 142.410 29.055 142.615 ;
        RECT 29.785 142.495 29.955 143.075 ;
        RECT 29.740 142.445 29.955 142.495 ;
        RECT 28.160 142.035 29.055 142.410 ;
        RECT 29.565 142.365 29.955 142.445 ;
        RECT 27.105 141.605 27.990 141.775 ;
        RECT 28.170 141.305 28.485 141.805 ;
        RECT 28.715 141.475 29.055 142.035 ;
        RECT 29.225 141.305 29.395 142.315 ;
        RECT 29.565 141.520 29.895 142.365 ;
        RECT 30.130 142.315 30.480 142.965 ;
        RECT 30.650 142.145 30.880 143.135 ;
        RECT 30.215 141.975 30.880 142.145 ;
        RECT 30.215 141.475 30.385 141.975 ;
        RECT 30.555 141.305 30.885 141.805 ;
        RECT 31.055 141.475 31.240 143.595 ;
        RECT 31.495 143.395 31.745 143.855 ;
        RECT 31.915 143.405 32.250 143.575 ;
        RECT 32.445 143.405 33.120 143.575 ;
        RECT 31.915 143.265 32.085 143.405 ;
        RECT 31.410 142.275 31.690 143.225 ;
        RECT 31.860 143.135 32.085 143.265 ;
        RECT 31.860 142.030 32.030 143.135 ;
        RECT 32.255 142.985 32.780 143.205 ;
        RECT 32.200 142.220 32.440 142.815 ;
        RECT 32.610 142.285 32.780 142.985 ;
        RECT 32.950 142.625 33.120 143.405 ;
        RECT 33.440 143.355 33.810 143.855 ;
        RECT 33.990 143.405 34.395 143.575 ;
        RECT 34.565 143.405 35.350 143.575 ;
        RECT 33.990 143.175 34.160 143.405 ;
        RECT 33.330 142.875 34.160 143.175 ;
        RECT 34.545 142.905 35.010 143.235 ;
        RECT 33.330 142.845 33.530 142.875 ;
        RECT 33.650 142.625 33.820 142.695 ;
        RECT 32.950 142.455 33.820 142.625 ;
        RECT 33.310 142.365 33.820 142.455 ;
        RECT 31.860 141.900 32.165 142.030 ;
        RECT 32.610 141.920 33.140 142.285 ;
        RECT 31.480 141.305 31.745 141.765 ;
        RECT 31.915 141.475 32.165 141.900 ;
        RECT 33.310 141.750 33.480 142.365 ;
        RECT 32.375 141.580 33.480 141.750 ;
        RECT 33.650 141.305 33.820 142.105 ;
        RECT 33.990 141.805 34.160 142.875 ;
        RECT 34.330 141.975 34.520 142.695 ;
        RECT 34.690 141.945 35.010 142.905 ;
        RECT 35.180 142.945 35.350 143.405 ;
        RECT 35.625 143.325 35.835 143.855 ;
        RECT 36.095 143.115 36.425 143.640 ;
        RECT 36.595 143.245 36.765 143.855 ;
        RECT 36.935 143.200 37.265 143.635 ;
        RECT 37.435 143.340 37.605 143.855 ;
        RECT 36.935 143.115 37.315 143.200 ;
        RECT 37.945 143.130 38.235 143.855 ;
        RECT 38.495 143.305 38.665 143.595 ;
        RECT 38.835 143.475 39.165 143.855 ;
        RECT 38.495 143.135 39.160 143.305 ;
        RECT 36.225 142.945 36.425 143.115 ;
        RECT 37.090 143.075 37.315 143.115 ;
        RECT 35.180 142.615 36.055 142.945 ;
        RECT 36.225 142.615 36.975 142.945 ;
        RECT 33.990 141.475 34.240 141.805 ;
        RECT 35.180 141.775 35.350 142.615 ;
        RECT 36.225 142.410 36.415 142.615 ;
        RECT 37.145 142.495 37.315 143.075 ;
        RECT 37.100 142.445 37.315 142.495 ;
        RECT 35.520 142.035 36.415 142.410 ;
        RECT 36.925 142.365 37.315 142.445 ;
        RECT 34.465 141.605 35.350 141.775 ;
        RECT 35.530 141.305 35.845 141.805 ;
        RECT 36.075 141.475 36.415 142.035 ;
        RECT 36.585 141.305 36.755 142.315 ;
        RECT 36.925 141.520 37.255 142.365 ;
        RECT 37.425 141.305 37.595 142.220 ;
        RECT 37.945 141.305 38.235 142.470 ;
        RECT 38.410 142.315 38.760 142.965 ;
        RECT 38.930 142.145 39.160 143.135 ;
        RECT 38.495 141.975 39.160 142.145 ;
        RECT 38.495 141.475 38.665 141.975 ;
        RECT 38.835 141.305 39.165 141.805 ;
        RECT 39.335 141.475 39.520 143.595 ;
        RECT 39.775 143.395 40.025 143.855 ;
        RECT 40.195 143.405 40.530 143.575 ;
        RECT 40.725 143.405 41.400 143.575 ;
        RECT 40.195 143.265 40.365 143.405 ;
        RECT 39.690 142.275 39.970 143.225 ;
        RECT 40.140 143.135 40.365 143.265 ;
        RECT 40.140 142.030 40.310 143.135 ;
        RECT 40.535 142.985 41.060 143.205 ;
        RECT 40.480 142.220 40.720 142.815 ;
        RECT 40.890 142.285 41.060 142.985 ;
        RECT 41.230 142.625 41.400 143.405 ;
        RECT 41.720 143.355 42.090 143.855 ;
        RECT 42.270 143.405 42.675 143.575 ;
        RECT 42.845 143.405 43.630 143.575 ;
        RECT 42.270 143.175 42.440 143.405 ;
        RECT 41.610 142.875 42.440 143.175 ;
        RECT 42.825 142.905 43.290 143.235 ;
        RECT 41.610 142.845 41.810 142.875 ;
        RECT 41.930 142.625 42.100 142.695 ;
        RECT 41.230 142.455 42.100 142.625 ;
        RECT 41.590 142.365 42.100 142.455 ;
        RECT 40.140 141.900 40.445 142.030 ;
        RECT 40.890 141.920 41.420 142.285 ;
        RECT 39.760 141.305 40.025 141.765 ;
        RECT 40.195 141.475 40.445 141.900 ;
        RECT 41.590 141.750 41.760 142.365 ;
        RECT 40.655 141.580 41.760 141.750 ;
        RECT 41.930 141.305 42.100 142.105 ;
        RECT 42.270 141.805 42.440 142.875 ;
        RECT 42.610 141.975 42.800 142.695 ;
        RECT 42.970 141.945 43.290 142.905 ;
        RECT 43.460 142.945 43.630 143.405 ;
        RECT 43.905 143.325 44.115 143.855 ;
        RECT 44.375 143.115 44.705 143.640 ;
        RECT 44.875 143.245 45.045 143.855 ;
        RECT 45.215 143.200 45.545 143.635 ;
        RECT 46.775 143.305 46.945 143.595 ;
        RECT 47.115 143.475 47.445 143.855 ;
        RECT 45.215 143.115 45.595 143.200 ;
        RECT 46.775 143.135 47.440 143.305 ;
        RECT 44.505 142.945 44.705 143.115 ;
        RECT 45.370 143.075 45.595 143.115 ;
        RECT 43.460 142.615 44.335 142.945 ;
        RECT 44.505 142.615 45.255 142.945 ;
        RECT 42.270 141.475 42.520 141.805 ;
        RECT 43.460 141.775 43.630 142.615 ;
        RECT 44.505 142.410 44.695 142.615 ;
        RECT 45.425 142.495 45.595 143.075 ;
        RECT 45.380 142.445 45.595 142.495 ;
        RECT 43.800 142.035 44.695 142.410 ;
        RECT 45.205 142.365 45.595 142.445 ;
        RECT 42.745 141.605 43.630 141.775 ;
        RECT 43.810 141.305 44.125 141.805 ;
        RECT 44.355 141.475 44.695 142.035 ;
        RECT 44.865 141.305 45.035 142.315 ;
        RECT 45.205 141.520 45.535 142.365 ;
        RECT 46.690 142.315 47.040 142.965 ;
        RECT 47.210 142.145 47.440 143.135 ;
        RECT 46.775 141.975 47.440 142.145 ;
        RECT 46.775 141.475 46.945 141.975 ;
        RECT 47.115 141.305 47.445 141.805 ;
        RECT 47.615 141.475 47.800 143.595 ;
        RECT 48.055 143.395 48.305 143.855 ;
        RECT 48.475 143.405 48.810 143.575 ;
        RECT 49.005 143.405 49.680 143.575 ;
        RECT 48.475 143.265 48.645 143.405 ;
        RECT 47.970 142.275 48.250 143.225 ;
        RECT 48.420 143.135 48.645 143.265 ;
        RECT 48.420 142.030 48.590 143.135 ;
        RECT 48.815 142.985 49.340 143.205 ;
        RECT 48.760 142.220 49.000 142.815 ;
        RECT 49.170 142.285 49.340 142.985 ;
        RECT 49.510 142.625 49.680 143.405 ;
        RECT 50.000 143.355 50.370 143.855 ;
        RECT 50.550 143.405 50.955 143.575 ;
        RECT 51.125 143.405 51.910 143.575 ;
        RECT 50.550 143.175 50.720 143.405 ;
        RECT 49.890 142.875 50.720 143.175 ;
        RECT 51.105 142.905 51.570 143.235 ;
        RECT 49.890 142.845 50.090 142.875 ;
        RECT 50.210 142.625 50.380 142.695 ;
        RECT 49.510 142.455 50.380 142.625 ;
        RECT 49.870 142.365 50.380 142.455 ;
        RECT 48.420 141.900 48.725 142.030 ;
        RECT 49.170 141.920 49.700 142.285 ;
        RECT 48.040 141.305 48.305 141.765 ;
        RECT 48.475 141.475 48.725 141.900 ;
        RECT 49.870 141.750 50.040 142.365 ;
        RECT 48.935 141.580 50.040 141.750 ;
        RECT 50.210 141.305 50.380 142.105 ;
        RECT 50.550 141.805 50.720 142.875 ;
        RECT 50.890 141.975 51.080 142.695 ;
        RECT 51.250 141.945 51.570 142.905 ;
        RECT 51.740 142.945 51.910 143.405 ;
        RECT 52.185 143.325 52.395 143.855 ;
        RECT 52.655 143.115 52.985 143.640 ;
        RECT 53.155 143.245 53.325 143.855 ;
        RECT 53.495 143.200 53.825 143.635 ;
        RECT 53.495 143.115 53.875 143.200 ;
        RECT 52.785 142.945 52.985 143.115 ;
        RECT 53.650 143.075 53.875 143.115 ;
        RECT 51.740 142.615 52.615 142.945 ;
        RECT 52.785 142.615 53.535 142.945 ;
        RECT 50.550 141.475 50.800 141.805 ;
        RECT 51.740 141.775 51.910 142.615 ;
        RECT 52.785 142.410 52.975 142.615 ;
        RECT 53.705 142.495 53.875 143.075 ;
        RECT 53.660 142.445 53.875 142.495 ;
        RECT 52.080 142.035 52.975 142.410 ;
        RECT 53.485 142.365 53.875 142.445 ;
        RECT 54.510 143.115 54.765 143.685 ;
        RECT 54.935 143.455 55.265 143.855 ;
        RECT 55.690 143.320 56.220 143.685 ;
        RECT 55.690 143.285 55.865 143.320 ;
        RECT 54.935 143.115 55.865 143.285 ;
        RECT 54.510 142.445 54.680 143.115 ;
        RECT 54.935 142.945 55.105 143.115 ;
        RECT 54.850 142.615 55.105 142.945 ;
        RECT 55.330 142.615 55.525 142.945 ;
        RECT 51.025 141.605 51.910 141.775 ;
        RECT 52.090 141.305 52.405 141.805 ;
        RECT 52.635 141.475 52.975 142.035 ;
        RECT 53.145 141.305 53.315 142.315 ;
        RECT 53.485 141.520 53.815 142.365 ;
        RECT 54.510 141.475 54.845 142.445 ;
        RECT 55.015 141.305 55.185 142.445 ;
        RECT 55.355 141.645 55.525 142.615 ;
        RECT 55.695 141.985 55.865 143.115 ;
        RECT 56.035 142.325 56.205 143.125 ;
        RECT 56.410 142.835 56.685 143.685 ;
        RECT 56.405 142.665 56.685 142.835 ;
        RECT 56.410 142.525 56.685 142.665 ;
        RECT 56.855 142.325 57.045 143.685 ;
        RECT 57.225 143.320 57.735 143.855 ;
        RECT 57.955 143.045 58.200 143.650 ;
        RECT 58.645 143.115 59.030 143.685 ;
        RECT 59.200 143.395 59.525 143.855 ;
        RECT 60.045 143.225 60.325 143.685 ;
        RECT 57.245 142.875 58.475 143.045 ;
        RECT 56.035 142.155 57.045 142.325 ;
        RECT 57.215 142.310 57.965 142.500 ;
        RECT 55.695 141.815 56.820 141.985 ;
        RECT 57.215 141.645 57.385 142.310 ;
        RECT 58.135 142.065 58.475 142.875 ;
        RECT 55.355 141.475 57.385 141.645 ;
        RECT 57.555 141.305 57.725 142.065 ;
        RECT 57.960 141.655 58.475 142.065 ;
        RECT 58.645 142.445 58.925 143.115 ;
        RECT 59.200 143.055 60.325 143.225 ;
        RECT 59.200 142.945 59.650 143.055 ;
        RECT 59.095 142.615 59.650 142.945 ;
        RECT 60.515 142.885 60.915 143.685 ;
        RECT 61.315 143.395 61.585 143.855 ;
        RECT 61.755 143.225 62.040 143.685 ;
        RECT 58.645 141.475 59.030 142.445 ;
        RECT 59.200 142.155 59.650 142.615 ;
        RECT 59.820 142.325 60.915 142.885 ;
        RECT 59.200 141.935 60.325 142.155 ;
        RECT 59.200 141.305 59.525 141.765 ;
        RECT 60.045 141.475 60.325 141.935 ;
        RECT 60.515 141.475 60.915 142.325 ;
        RECT 61.085 143.055 62.040 143.225 ;
        RECT 62.325 143.105 63.535 143.855 ;
        RECT 63.705 143.130 63.995 143.855 ;
        RECT 64.410 143.375 64.710 143.855 ;
        RECT 64.880 143.205 65.140 143.660 ;
        RECT 65.310 143.375 65.570 143.855 ;
        RECT 65.740 143.205 66.000 143.660 ;
        RECT 66.170 143.375 66.430 143.855 ;
        RECT 66.600 143.205 66.860 143.660 ;
        RECT 67.030 143.375 67.290 143.855 ;
        RECT 67.460 143.205 67.720 143.660 ;
        RECT 67.890 143.330 68.150 143.855 ;
        RECT 61.085 142.155 61.295 143.055 ;
        RECT 61.465 142.325 62.155 142.885 ;
        RECT 62.325 142.565 62.845 143.105 ;
        RECT 64.410 143.035 67.720 143.205 ;
        RECT 63.015 142.395 63.535 142.935 ;
        RECT 61.085 141.935 62.040 142.155 ;
        RECT 61.315 141.305 61.585 141.765 ;
        RECT 61.755 141.475 62.040 141.935 ;
        RECT 62.325 141.305 63.535 142.395 ;
        RECT 63.705 141.305 63.995 142.470 ;
        RECT 64.410 142.445 65.380 143.035 ;
        RECT 68.320 142.865 68.570 143.675 ;
        RECT 68.750 143.395 68.995 143.855 ;
        RECT 65.550 142.615 68.570 142.865 ;
        RECT 68.740 142.615 69.055 143.225 ;
        RECT 69.230 143.115 69.485 143.685 ;
        RECT 69.655 143.455 69.985 143.855 ;
        RECT 70.410 143.320 70.940 143.685 ;
        RECT 71.130 143.515 71.405 143.685 ;
        RECT 71.125 143.345 71.405 143.515 ;
        RECT 70.410 143.285 70.585 143.320 ;
        RECT 69.655 143.115 70.585 143.285 ;
        RECT 64.410 142.205 67.720 142.445 ;
        RECT 64.415 141.305 64.710 142.035 ;
        RECT 64.880 141.480 65.140 142.205 ;
        RECT 65.310 141.305 65.570 142.035 ;
        RECT 65.740 141.480 66.000 142.205 ;
        RECT 66.170 141.305 66.430 142.035 ;
        RECT 66.600 141.480 66.860 142.205 ;
        RECT 67.030 141.305 67.290 142.035 ;
        RECT 67.460 141.480 67.720 142.205 ;
        RECT 67.890 141.305 68.150 142.415 ;
        RECT 68.320 141.480 68.570 142.615 ;
        RECT 69.230 142.445 69.400 143.115 ;
        RECT 69.655 142.945 69.825 143.115 ;
        RECT 69.570 142.615 69.825 142.945 ;
        RECT 70.050 142.615 70.245 142.945 ;
        RECT 68.750 141.305 69.045 142.415 ;
        RECT 69.230 141.475 69.565 142.445 ;
        RECT 69.735 141.305 69.905 142.445 ;
        RECT 70.075 141.645 70.245 142.615 ;
        RECT 70.415 141.985 70.585 143.115 ;
        RECT 70.755 142.325 70.925 143.125 ;
        RECT 71.130 142.525 71.405 143.345 ;
        RECT 71.575 142.325 71.765 143.685 ;
        RECT 71.945 143.320 72.455 143.855 ;
        RECT 72.675 143.045 72.920 143.650 ;
        RECT 73.875 143.200 74.205 143.635 ;
        RECT 74.375 143.245 74.545 143.855 ;
        RECT 73.825 143.115 74.205 143.200 ;
        RECT 74.715 143.115 75.045 143.640 ;
        RECT 75.305 143.325 75.515 143.855 ;
        RECT 75.790 143.405 76.575 143.575 ;
        RECT 76.745 143.405 77.150 143.575 ;
        RECT 73.825 143.075 74.050 143.115 ;
        RECT 71.965 142.875 73.195 143.045 ;
        RECT 70.755 142.155 71.765 142.325 ;
        RECT 71.935 142.310 72.685 142.500 ;
        RECT 70.415 141.815 71.540 141.985 ;
        RECT 71.935 141.645 72.105 142.310 ;
        RECT 72.855 142.065 73.195 142.875 ;
        RECT 73.825 142.495 73.995 143.075 ;
        RECT 74.715 142.945 74.915 143.115 ;
        RECT 75.790 142.945 75.960 143.405 ;
        RECT 74.165 142.615 74.915 142.945 ;
        RECT 75.085 142.615 75.960 142.945 ;
        RECT 73.825 142.445 74.040 142.495 ;
        RECT 73.825 142.365 74.215 142.445 ;
        RECT 70.075 141.475 72.105 141.645 ;
        RECT 72.275 141.305 72.445 142.065 ;
        RECT 72.680 141.655 73.195 142.065 ;
        RECT 73.885 141.520 74.215 142.365 ;
        RECT 74.725 142.410 74.915 142.615 ;
        RECT 74.385 141.305 74.555 142.315 ;
        RECT 74.725 142.035 75.620 142.410 ;
        RECT 74.725 141.475 75.065 142.035 ;
        RECT 75.295 141.305 75.610 141.805 ;
        RECT 75.790 141.775 75.960 142.615 ;
        RECT 76.130 142.905 76.595 143.235 ;
        RECT 76.980 143.175 77.150 143.405 ;
        RECT 77.330 143.355 77.700 143.855 ;
        RECT 78.020 143.405 78.695 143.575 ;
        RECT 78.890 143.405 79.225 143.575 ;
        RECT 76.130 141.945 76.450 142.905 ;
        RECT 76.980 142.875 77.810 143.175 ;
        RECT 76.620 141.975 76.810 142.695 ;
        RECT 76.980 141.805 77.150 142.875 ;
        RECT 77.610 142.845 77.810 142.875 ;
        RECT 77.320 142.625 77.490 142.695 ;
        RECT 78.020 142.625 78.190 143.405 ;
        RECT 79.055 143.265 79.225 143.405 ;
        RECT 79.395 143.395 79.645 143.855 ;
        RECT 77.320 142.455 78.190 142.625 ;
        RECT 78.360 142.985 78.885 143.205 ;
        RECT 79.055 143.135 79.280 143.265 ;
        RECT 77.320 142.365 77.830 142.455 ;
        RECT 75.790 141.605 76.675 141.775 ;
        RECT 76.900 141.475 77.150 141.805 ;
        RECT 77.320 141.305 77.490 142.105 ;
        RECT 77.660 141.750 77.830 142.365 ;
        RECT 78.360 142.285 78.530 142.985 ;
        RECT 78.000 141.920 78.530 142.285 ;
        RECT 78.700 142.220 78.940 142.815 ;
        RECT 79.110 142.030 79.280 143.135 ;
        RECT 79.450 142.275 79.730 143.225 ;
        RECT 78.975 141.900 79.280 142.030 ;
        RECT 77.660 141.580 78.765 141.750 ;
        RECT 78.975 141.475 79.225 141.900 ;
        RECT 79.395 141.305 79.660 141.765 ;
        RECT 79.900 141.475 80.085 143.595 ;
        RECT 80.255 143.475 80.585 143.855 ;
        RECT 80.755 143.305 80.925 143.595 ;
        RECT 80.260 143.135 80.925 143.305 ;
        RECT 81.275 143.305 81.445 143.595 ;
        RECT 81.615 143.475 81.945 143.855 ;
        RECT 81.275 143.135 81.940 143.305 ;
        RECT 80.260 142.145 80.490 143.135 ;
        RECT 80.660 142.315 81.010 142.965 ;
        RECT 81.190 142.315 81.540 142.965 ;
        RECT 81.710 142.145 81.940 143.135 ;
        RECT 80.260 141.975 80.925 142.145 ;
        RECT 80.255 141.305 80.585 141.805 ;
        RECT 80.755 141.475 80.925 141.975 ;
        RECT 81.275 141.975 81.940 142.145 ;
        RECT 81.275 141.475 81.445 141.975 ;
        RECT 81.615 141.305 81.945 141.805 ;
        RECT 82.115 141.475 82.300 143.595 ;
        RECT 82.555 143.395 82.805 143.855 ;
        RECT 82.975 143.405 83.310 143.575 ;
        RECT 83.505 143.405 84.180 143.575 ;
        RECT 82.975 143.265 83.145 143.405 ;
        RECT 82.470 142.275 82.750 143.225 ;
        RECT 82.920 143.135 83.145 143.265 ;
        RECT 82.920 142.030 83.090 143.135 ;
        RECT 83.315 142.985 83.840 143.205 ;
        RECT 83.260 142.220 83.500 142.815 ;
        RECT 83.670 142.285 83.840 142.985 ;
        RECT 84.010 142.625 84.180 143.405 ;
        RECT 84.500 143.355 84.870 143.855 ;
        RECT 85.050 143.405 85.455 143.575 ;
        RECT 85.625 143.405 86.410 143.575 ;
        RECT 85.050 143.175 85.220 143.405 ;
        RECT 84.390 142.875 85.220 143.175 ;
        RECT 85.605 142.905 86.070 143.235 ;
        RECT 84.390 142.845 84.590 142.875 ;
        RECT 84.710 142.625 84.880 142.695 ;
        RECT 84.010 142.455 84.880 142.625 ;
        RECT 84.370 142.365 84.880 142.455 ;
        RECT 82.920 141.900 83.225 142.030 ;
        RECT 83.670 141.920 84.200 142.285 ;
        RECT 82.540 141.305 82.805 141.765 ;
        RECT 82.975 141.475 83.225 141.900 ;
        RECT 84.370 141.750 84.540 142.365 ;
        RECT 83.435 141.580 84.540 141.750 ;
        RECT 84.710 141.305 84.880 142.105 ;
        RECT 85.050 141.805 85.220 142.875 ;
        RECT 85.390 141.975 85.580 142.695 ;
        RECT 85.750 141.945 86.070 142.905 ;
        RECT 86.240 142.945 86.410 143.405 ;
        RECT 86.685 143.325 86.895 143.855 ;
        RECT 87.155 143.115 87.485 143.640 ;
        RECT 87.655 143.245 87.825 143.855 ;
        RECT 87.995 143.200 88.325 143.635 ;
        RECT 87.995 143.115 88.375 143.200 ;
        RECT 87.285 142.945 87.485 143.115 ;
        RECT 88.150 143.075 88.375 143.115 ;
        RECT 88.545 143.105 89.755 143.855 ;
        RECT 86.240 142.615 87.115 142.945 ;
        RECT 87.285 142.615 88.035 142.945 ;
        RECT 85.050 141.475 85.300 141.805 ;
        RECT 86.240 141.775 86.410 142.615 ;
        RECT 87.285 142.410 87.475 142.615 ;
        RECT 88.205 142.495 88.375 143.075 ;
        RECT 88.160 142.445 88.375 142.495 ;
        RECT 86.580 142.035 87.475 142.410 ;
        RECT 87.985 142.365 88.375 142.445 ;
        RECT 88.545 142.395 89.065 142.935 ;
        RECT 89.235 142.565 89.755 143.105 ;
        RECT 85.525 141.605 86.410 141.775 ;
        RECT 86.590 141.305 86.905 141.805 ;
        RECT 87.135 141.475 87.475 142.035 ;
        RECT 87.645 141.305 87.815 142.315 ;
        RECT 87.985 141.520 88.315 142.365 ;
        RECT 88.545 141.305 89.755 142.395 ;
        RECT 12.100 141.135 89.840 141.305 ;
        RECT 12.185 140.045 13.395 141.135 ;
        RECT 13.565 140.045 16.155 141.135 ;
        RECT 12.185 139.335 12.705 139.875 ;
        RECT 12.875 139.505 13.395 140.045 ;
        RECT 13.565 139.355 14.775 139.875 ;
        RECT 14.945 139.525 16.155 140.045 ;
        RECT 16.325 140.035 16.645 140.965 ;
        RECT 16.825 140.455 17.225 140.965 ;
        RECT 17.395 140.625 17.565 141.135 ;
        RECT 17.735 140.455 18.065 140.965 ;
        RECT 16.825 140.285 18.065 140.455 ;
        RECT 18.235 140.285 18.405 141.135 ;
        RECT 18.995 140.285 19.375 140.965 ;
        RECT 16.325 139.865 16.955 140.035 ;
        RECT 12.185 138.585 13.395 139.335 ;
        RECT 13.565 138.585 16.155 139.355 ;
        RECT 16.325 138.585 16.615 139.420 ;
        RECT 16.785 138.985 16.955 139.865 ;
        RECT 17.730 139.945 19.035 140.115 ;
        RECT 17.125 139.325 17.355 139.825 ;
        RECT 17.730 139.745 17.900 139.945 ;
        RECT 17.525 139.575 17.900 139.745 ;
        RECT 18.070 139.575 18.620 139.775 ;
        RECT 18.790 139.495 19.035 139.945 ;
        RECT 19.205 139.325 19.375 140.285 ;
        RECT 17.125 139.155 19.375 139.325 ;
        RECT 19.545 139.995 19.805 140.965 ;
        RECT 20.000 140.725 20.330 141.135 ;
        RECT 20.530 140.545 20.700 140.965 ;
        RECT 20.915 140.725 21.585 141.135 ;
        RECT 21.820 140.545 21.990 140.965 ;
        RECT 22.295 140.695 22.625 141.135 ;
        RECT 19.975 140.375 21.990 140.545 ;
        RECT 22.795 140.515 22.970 140.965 ;
        RECT 19.545 139.305 19.715 139.995 ;
        RECT 19.975 139.825 20.145 140.375 ;
        RECT 19.885 139.495 20.145 139.825 ;
        RECT 16.785 138.815 17.740 138.985 ;
        RECT 18.155 138.585 18.485 138.975 ;
        RECT 18.655 138.835 18.825 139.155 ;
        RECT 18.995 138.585 19.325 138.975 ;
        RECT 19.545 138.840 19.885 139.305 ;
        RECT 20.315 139.165 20.655 140.195 ;
        RECT 20.845 139.095 21.115 140.195 ;
        RECT 19.550 138.795 19.885 138.840 ;
        RECT 20.055 138.585 20.385 138.965 ;
        RECT 20.845 138.925 21.155 139.095 ;
        RECT 20.845 138.920 21.115 138.925 ;
        RECT 21.340 138.920 21.620 140.195 ;
        RECT 21.820 139.085 21.990 140.375 ;
        RECT 22.340 140.345 22.970 140.515 ;
        RECT 23.235 140.525 23.565 140.955 ;
        RECT 23.745 140.695 23.940 141.135 ;
        RECT 24.110 140.525 24.440 140.955 ;
        RECT 23.235 140.355 24.440 140.525 ;
        RECT 22.340 139.825 22.510 140.345 ;
        RECT 22.160 139.495 22.510 139.825 ;
        RECT 22.690 139.495 23.055 140.175 ;
        RECT 23.235 140.025 24.130 140.355 ;
        RECT 24.610 140.185 24.885 140.955 ;
        RECT 24.300 139.995 24.885 140.185 ;
        RECT 23.240 139.495 23.535 139.825 ;
        RECT 23.715 139.495 24.130 139.825 ;
        RECT 22.340 139.325 22.510 139.495 ;
        RECT 22.340 139.155 22.970 139.325 ;
        RECT 21.820 138.755 22.050 139.085 ;
        RECT 22.295 138.585 22.625 138.965 ;
        RECT 22.795 138.755 22.970 139.155 ;
        RECT 23.235 138.585 23.535 139.315 ;
        RECT 23.715 138.875 23.945 139.495 ;
        RECT 24.300 139.325 24.475 139.995 ;
        RECT 25.065 139.970 25.355 141.135 ;
        RECT 26.530 140.515 26.705 140.965 ;
        RECT 26.875 140.695 27.205 141.135 ;
        RECT 27.510 140.545 27.680 140.965 ;
        RECT 27.915 140.725 28.585 141.135 ;
        RECT 28.800 140.545 28.970 140.965 ;
        RECT 29.170 140.725 29.500 141.135 ;
        RECT 26.530 140.345 27.160 140.515 ;
        RECT 24.145 139.145 24.475 139.325 ;
        RECT 24.645 139.175 24.885 139.825 ;
        RECT 26.445 139.495 26.810 140.175 ;
        RECT 26.990 139.825 27.160 140.345 ;
        RECT 27.510 140.375 29.525 140.545 ;
        RECT 26.990 139.495 27.340 139.825 ;
        RECT 26.990 139.325 27.160 139.495 ;
        RECT 24.145 138.765 24.370 139.145 ;
        RECT 24.540 138.585 24.870 138.975 ;
        RECT 25.065 138.585 25.355 139.310 ;
        RECT 26.530 139.155 27.160 139.325 ;
        RECT 26.530 138.755 26.705 139.155 ;
        RECT 27.510 139.085 27.680 140.375 ;
        RECT 26.875 138.585 27.205 138.965 ;
        RECT 27.450 138.755 27.680 139.085 ;
        RECT 27.880 138.920 28.160 140.195 ;
        RECT 28.385 139.435 28.655 140.195 ;
        RECT 28.345 139.265 28.655 139.435 ;
        RECT 28.385 138.920 28.655 139.265 ;
        RECT 28.845 139.165 29.185 140.195 ;
        RECT 29.355 139.825 29.525 140.375 ;
        RECT 29.695 139.995 29.955 140.965 ;
        RECT 30.210 140.515 30.385 140.965 ;
        RECT 30.555 140.695 30.885 141.135 ;
        RECT 31.190 140.545 31.360 140.965 ;
        RECT 31.595 140.725 32.265 141.135 ;
        RECT 32.480 140.545 32.650 140.965 ;
        RECT 32.850 140.725 33.180 141.135 ;
        RECT 30.210 140.345 30.840 140.515 ;
        RECT 29.355 139.495 29.615 139.825 ;
        RECT 29.785 139.305 29.955 139.995 ;
        RECT 30.125 139.495 30.490 140.175 ;
        RECT 30.670 139.825 30.840 140.345 ;
        RECT 31.190 140.375 33.205 140.545 ;
        RECT 30.670 139.495 31.020 139.825 ;
        RECT 30.670 139.325 30.840 139.495 ;
        RECT 29.115 138.585 29.445 138.965 ;
        RECT 29.615 138.840 29.955 139.305 ;
        RECT 30.210 139.155 30.840 139.325 ;
        RECT 29.615 138.795 29.950 138.840 ;
        RECT 30.210 138.755 30.385 139.155 ;
        RECT 31.190 139.085 31.360 140.375 ;
        RECT 30.555 138.585 30.885 138.965 ;
        RECT 31.130 138.755 31.360 139.085 ;
        RECT 31.560 138.920 31.840 140.195 ;
        RECT 32.065 140.115 32.335 140.195 ;
        RECT 32.025 139.945 32.335 140.115 ;
        RECT 32.065 138.920 32.335 139.945 ;
        RECT 32.525 139.165 32.865 140.195 ;
        RECT 33.035 139.825 33.205 140.375 ;
        RECT 33.375 139.995 33.635 140.965 ;
        RECT 33.815 140.525 34.145 140.955 ;
        RECT 34.325 140.695 34.520 141.135 ;
        RECT 34.690 140.525 35.020 140.955 ;
        RECT 33.815 140.355 35.020 140.525 ;
        RECT 33.815 140.025 34.710 140.355 ;
        RECT 35.190 140.185 35.465 140.955 ;
        RECT 33.035 139.495 33.295 139.825 ;
        RECT 33.465 139.305 33.635 139.995 ;
        RECT 34.880 139.995 35.465 140.185 ;
        RECT 35.655 140.185 35.930 140.955 ;
        RECT 36.100 140.525 36.430 140.955 ;
        RECT 36.600 140.695 36.795 141.135 ;
        RECT 36.975 140.525 37.305 140.955 ;
        RECT 36.100 140.355 37.305 140.525 ;
        RECT 35.655 139.995 36.240 140.185 ;
        RECT 36.410 140.025 37.305 140.355 ;
        RECT 37.945 139.995 38.225 141.135 ;
        RECT 33.820 139.495 34.115 139.825 ;
        RECT 34.295 139.495 34.710 139.825 ;
        RECT 32.795 138.585 33.125 138.965 ;
        RECT 33.295 138.840 33.635 139.305 ;
        RECT 33.295 138.795 33.630 138.840 ;
        RECT 33.815 138.585 34.115 139.315 ;
        RECT 34.295 138.875 34.525 139.495 ;
        RECT 34.880 139.325 35.055 139.995 ;
        RECT 34.725 139.145 35.055 139.325 ;
        RECT 35.225 139.175 35.465 139.825 ;
        RECT 35.655 139.175 35.895 139.825 ;
        RECT 36.065 139.325 36.240 139.995 ;
        RECT 38.395 139.985 38.725 140.965 ;
        RECT 38.895 139.995 39.155 141.135 ;
        RECT 39.415 140.465 39.585 140.965 ;
        RECT 39.755 140.635 40.085 141.135 ;
        RECT 39.415 140.295 40.080 140.465 ;
        RECT 36.410 139.495 36.825 139.825 ;
        RECT 37.005 139.495 37.300 139.825 ;
        RECT 37.955 139.555 38.290 139.825 ;
        RECT 36.065 139.145 36.395 139.325 ;
        RECT 34.725 138.765 34.950 139.145 ;
        RECT 35.120 138.585 35.450 138.975 ;
        RECT 35.670 138.585 36.000 138.975 ;
        RECT 36.170 138.765 36.395 139.145 ;
        RECT 36.595 138.875 36.825 139.495 ;
        RECT 38.460 139.385 38.630 139.985 ;
        RECT 38.800 139.575 39.135 139.825 ;
        RECT 39.330 139.475 39.680 140.125 ;
        RECT 37.005 138.585 37.305 139.315 ;
        RECT 37.945 138.585 38.255 139.385 ;
        RECT 38.460 138.755 39.155 139.385 ;
        RECT 39.850 139.305 40.080 140.295 ;
        RECT 39.415 139.135 40.080 139.305 ;
        RECT 39.415 138.845 39.585 139.135 ;
        RECT 39.755 138.585 40.085 138.965 ;
        RECT 40.255 138.845 40.440 140.965 ;
        RECT 40.680 140.675 40.945 141.135 ;
        RECT 41.115 140.540 41.365 140.965 ;
        RECT 41.575 140.690 42.680 140.860 ;
        RECT 41.060 140.410 41.365 140.540 ;
        RECT 40.610 139.215 40.890 140.165 ;
        RECT 41.060 139.305 41.230 140.410 ;
        RECT 41.400 139.625 41.640 140.220 ;
        RECT 41.810 140.155 42.340 140.520 ;
        RECT 41.810 139.455 41.980 140.155 ;
        RECT 42.510 140.075 42.680 140.690 ;
        RECT 42.850 140.335 43.020 141.135 ;
        RECT 43.190 140.635 43.440 140.965 ;
        RECT 43.665 140.665 44.550 140.835 ;
        RECT 42.510 139.985 43.020 140.075 ;
        RECT 41.060 139.175 41.285 139.305 ;
        RECT 41.455 139.235 41.980 139.455 ;
        RECT 42.150 139.815 43.020 139.985 ;
        RECT 40.695 138.585 40.945 139.045 ;
        RECT 41.115 139.035 41.285 139.175 ;
        RECT 42.150 139.035 42.320 139.815 ;
        RECT 42.850 139.745 43.020 139.815 ;
        RECT 42.530 139.565 42.730 139.595 ;
        RECT 43.190 139.565 43.360 140.635 ;
        RECT 43.530 139.745 43.720 140.465 ;
        RECT 42.530 139.265 43.360 139.565 ;
        RECT 43.890 139.535 44.210 140.495 ;
        RECT 41.115 138.865 41.450 139.035 ;
        RECT 41.645 138.865 42.320 139.035 ;
        RECT 42.640 138.585 43.010 139.085 ;
        RECT 43.190 139.035 43.360 139.265 ;
        RECT 43.745 139.205 44.210 139.535 ;
        RECT 44.380 139.825 44.550 140.665 ;
        RECT 44.730 140.635 45.045 141.135 ;
        RECT 45.275 140.405 45.615 140.965 ;
        RECT 44.720 140.030 45.615 140.405 ;
        RECT 45.785 140.125 45.955 141.135 ;
        RECT 45.425 139.825 45.615 140.030 ;
        RECT 46.125 140.075 46.455 140.920 ;
        RECT 46.125 139.995 46.515 140.075 ;
        RECT 46.300 139.945 46.515 139.995 ;
        RECT 44.380 139.495 45.255 139.825 ;
        RECT 45.425 139.495 46.175 139.825 ;
        RECT 44.380 139.035 44.550 139.495 ;
        RECT 45.425 139.325 45.625 139.495 ;
        RECT 46.345 139.365 46.515 139.945 ;
        RECT 46.290 139.325 46.515 139.365 ;
        RECT 43.190 138.865 43.595 139.035 ;
        RECT 43.765 138.865 44.550 139.035 ;
        RECT 44.825 138.585 45.035 139.115 ;
        RECT 45.295 138.800 45.625 139.325 ;
        RECT 46.135 139.240 46.515 139.325 ;
        RECT 46.690 139.995 47.025 140.965 ;
        RECT 47.195 139.995 47.365 141.135 ;
        RECT 47.535 140.795 49.565 140.965 ;
        RECT 46.690 139.325 46.860 139.995 ;
        RECT 47.535 139.825 47.705 140.795 ;
        RECT 47.030 139.495 47.285 139.825 ;
        RECT 47.510 139.495 47.705 139.825 ;
        RECT 47.875 140.455 49.000 140.625 ;
        RECT 47.115 139.325 47.285 139.495 ;
        RECT 47.875 139.325 48.045 140.455 ;
        RECT 45.795 138.585 45.965 139.195 ;
        RECT 46.135 138.805 46.465 139.240 ;
        RECT 46.690 138.755 46.945 139.325 ;
        RECT 47.115 139.155 48.045 139.325 ;
        RECT 48.215 140.115 49.225 140.285 ;
        RECT 48.215 139.315 48.385 140.115 ;
        RECT 48.590 139.435 48.865 139.915 ;
        RECT 48.585 139.265 48.865 139.435 ;
        RECT 47.870 139.120 48.045 139.155 ;
        RECT 47.115 138.585 47.445 138.985 ;
        RECT 47.870 138.755 48.400 139.120 ;
        RECT 48.590 138.755 48.865 139.265 ;
        RECT 49.035 138.755 49.225 140.115 ;
        RECT 49.395 140.130 49.565 140.795 ;
        RECT 49.735 140.375 49.905 141.135 ;
        RECT 50.140 140.375 50.655 140.785 ;
        RECT 49.395 139.940 50.145 140.130 ;
        RECT 50.315 139.565 50.655 140.375 ;
        RECT 50.825 139.970 51.115 141.135 ;
        RECT 51.375 140.465 51.545 140.965 ;
        RECT 51.715 140.635 52.045 141.135 ;
        RECT 51.375 140.295 52.040 140.465 ;
        RECT 49.425 139.395 50.655 139.565 ;
        RECT 51.290 139.475 51.640 140.125 ;
        RECT 49.405 138.585 49.915 139.120 ;
        RECT 50.135 138.790 50.380 139.395 ;
        RECT 50.825 138.585 51.115 139.310 ;
        RECT 51.810 139.305 52.040 140.295 ;
        RECT 51.375 139.135 52.040 139.305 ;
        RECT 51.375 138.845 51.545 139.135 ;
        RECT 51.715 138.585 52.045 138.965 ;
        RECT 52.215 138.845 52.400 140.965 ;
        RECT 52.640 140.675 52.905 141.135 ;
        RECT 53.075 140.540 53.325 140.965 ;
        RECT 53.535 140.690 54.640 140.860 ;
        RECT 53.020 140.410 53.325 140.540 ;
        RECT 52.570 139.215 52.850 140.165 ;
        RECT 53.020 139.305 53.190 140.410 ;
        RECT 53.360 139.625 53.600 140.220 ;
        RECT 53.770 140.155 54.300 140.520 ;
        RECT 53.770 139.455 53.940 140.155 ;
        RECT 54.470 140.075 54.640 140.690 ;
        RECT 54.810 140.335 54.980 141.135 ;
        RECT 55.150 140.635 55.400 140.965 ;
        RECT 55.625 140.665 56.510 140.835 ;
        RECT 54.470 139.985 54.980 140.075 ;
        RECT 53.020 139.175 53.245 139.305 ;
        RECT 53.415 139.235 53.940 139.455 ;
        RECT 54.110 139.815 54.980 139.985 ;
        RECT 52.655 138.585 52.905 139.045 ;
        RECT 53.075 139.035 53.245 139.175 ;
        RECT 54.110 139.035 54.280 139.815 ;
        RECT 54.810 139.745 54.980 139.815 ;
        RECT 54.490 139.565 54.690 139.595 ;
        RECT 55.150 139.565 55.320 140.635 ;
        RECT 55.490 139.745 55.680 140.465 ;
        RECT 54.490 139.265 55.320 139.565 ;
        RECT 55.850 139.535 56.170 140.495 ;
        RECT 53.075 138.865 53.410 139.035 ;
        RECT 53.605 138.865 54.280 139.035 ;
        RECT 54.600 138.585 54.970 139.085 ;
        RECT 55.150 139.035 55.320 139.265 ;
        RECT 55.705 139.205 56.170 139.535 ;
        RECT 56.340 139.825 56.510 140.665 ;
        RECT 56.690 140.635 57.005 141.135 ;
        RECT 57.235 140.405 57.575 140.965 ;
        RECT 56.680 140.030 57.575 140.405 ;
        RECT 57.745 140.125 57.915 141.135 ;
        RECT 57.385 139.825 57.575 140.030 ;
        RECT 58.085 140.075 58.415 140.920 ;
        RECT 58.735 140.465 58.905 140.965 ;
        RECT 59.075 140.635 59.405 141.135 ;
        RECT 58.735 140.295 59.400 140.465 ;
        RECT 58.085 139.995 58.475 140.075 ;
        RECT 58.260 139.945 58.475 139.995 ;
        RECT 56.340 139.495 57.215 139.825 ;
        RECT 57.385 139.495 58.135 139.825 ;
        RECT 56.340 139.035 56.510 139.495 ;
        RECT 57.385 139.325 57.585 139.495 ;
        RECT 58.305 139.365 58.475 139.945 ;
        RECT 58.650 139.475 59.000 140.125 ;
        RECT 58.250 139.325 58.475 139.365 ;
        RECT 55.150 138.865 55.555 139.035 ;
        RECT 55.725 138.865 56.510 139.035 ;
        RECT 56.785 138.585 56.995 139.115 ;
        RECT 57.255 138.800 57.585 139.325 ;
        RECT 58.095 139.240 58.475 139.325 ;
        RECT 59.170 139.305 59.400 140.295 ;
        RECT 57.755 138.585 57.925 139.195 ;
        RECT 58.095 138.805 58.425 139.240 ;
        RECT 58.735 139.135 59.400 139.305 ;
        RECT 58.735 138.845 58.905 139.135 ;
        RECT 59.075 138.585 59.405 138.965 ;
        RECT 59.575 138.845 59.760 140.965 ;
        RECT 60.000 140.675 60.265 141.135 ;
        RECT 60.435 140.540 60.685 140.965 ;
        RECT 60.895 140.690 62.000 140.860 ;
        RECT 60.380 140.410 60.685 140.540 ;
        RECT 59.930 139.215 60.210 140.165 ;
        RECT 60.380 139.305 60.550 140.410 ;
        RECT 60.720 139.625 60.960 140.220 ;
        RECT 61.130 140.155 61.660 140.520 ;
        RECT 61.130 139.455 61.300 140.155 ;
        RECT 61.830 140.075 62.000 140.690 ;
        RECT 62.170 140.335 62.340 141.135 ;
        RECT 62.510 140.635 62.760 140.965 ;
        RECT 62.985 140.665 63.870 140.835 ;
        RECT 61.830 139.985 62.340 140.075 ;
        RECT 60.380 139.175 60.605 139.305 ;
        RECT 60.775 139.235 61.300 139.455 ;
        RECT 61.470 139.815 62.340 139.985 ;
        RECT 60.015 138.585 60.265 139.045 ;
        RECT 60.435 139.035 60.605 139.175 ;
        RECT 61.470 139.035 61.640 139.815 ;
        RECT 62.170 139.745 62.340 139.815 ;
        RECT 61.850 139.565 62.050 139.595 ;
        RECT 62.510 139.565 62.680 140.635 ;
        RECT 62.850 139.745 63.040 140.465 ;
        RECT 61.850 139.265 62.680 139.565 ;
        RECT 63.210 139.535 63.530 140.495 ;
        RECT 60.435 138.865 60.770 139.035 ;
        RECT 60.965 138.865 61.640 139.035 ;
        RECT 61.960 138.585 62.330 139.085 ;
        RECT 62.510 139.035 62.680 139.265 ;
        RECT 63.065 139.205 63.530 139.535 ;
        RECT 63.700 139.825 63.870 140.665 ;
        RECT 64.050 140.635 64.365 141.135 ;
        RECT 64.595 140.405 64.935 140.965 ;
        RECT 64.040 140.030 64.935 140.405 ;
        RECT 65.105 140.125 65.275 141.135 ;
        RECT 64.745 139.825 64.935 140.030 ;
        RECT 65.445 140.075 65.775 140.920 ;
        RECT 66.065 140.075 66.395 140.920 ;
        RECT 66.565 140.125 66.735 141.135 ;
        RECT 66.905 140.405 67.245 140.965 ;
        RECT 67.475 140.635 67.790 141.135 ;
        RECT 67.970 140.665 68.855 140.835 ;
        RECT 65.445 139.995 65.835 140.075 ;
        RECT 65.620 139.945 65.835 139.995 ;
        RECT 63.700 139.495 64.575 139.825 ;
        RECT 64.745 139.495 65.495 139.825 ;
        RECT 63.700 139.035 63.870 139.495 ;
        RECT 64.745 139.325 64.945 139.495 ;
        RECT 65.665 139.365 65.835 139.945 ;
        RECT 65.610 139.325 65.835 139.365 ;
        RECT 62.510 138.865 62.915 139.035 ;
        RECT 63.085 138.865 63.870 139.035 ;
        RECT 64.145 138.585 64.355 139.115 ;
        RECT 64.615 138.800 64.945 139.325 ;
        RECT 65.455 139.240 65.835 139.325 ;
        RECT 66.005 139.995 66.395 140.075 ;
        RECT 66.905 140.030 67.800 140.405 ;
        RECT 66.005 139.945 66.220 139.995 ;
        RECT 66.005 139.365 66.175 139.945 ;
        RECT 66.905 139.825 67.095 140.030 ;
        RECT 67.970 139.825 68.140 140.665 ;
        RECT 69.080 140.635 69.330 140.965 ;
        RECT 66.345 139.495 67.095 139.825 ;
        RECT 67.265 139.495 68.140 139.825 ;
        RECT 66.005 139.325 66.230 139.365 ;
        RECT 66.895 139.325 67.095 139.495 ;
        RECT 66.005 139.240 66.385 139.325 ;
        RECT 65.115 138.585 65.285 139.195 ;
        RECT 65.455 138.805 65.785 139.240 ;
        RECT 66.055 138.805 66.385 139.240 ;
        RECT 66.555 138.585 66.725 139.195 ;
        RECT 66.895 138.800 67.225 139.325 ;
        RECT 67.485 138.585 67.695 139.115 ;
        RECT 67.970 139.035 68.140 139.495 ;
        RECT 68.310 139.535 68.630 140.495 ;
        RECT 68.800 139.745 68.990 140.465 ;
        RECT 69.160 139.565 69.330 140.635 ;
        RECT 69.500 140.335 69.670 141.135 ;
        RECT 69.840 140.690 70.945 140.860 ;
        RECT 69.840 140.075 70.010 140.690 ;
        RECT 71.155 140.540 71.405 140.965 ;
        RECT 71.575 140.675 71.840 141.135 ;
        RECT 70.180 140.155 70.710 140.520 ;
        RECT 71.155 140.410 71.460 140.540 ;
        RECT 69.500 139.985 70.010 140.075 ;
        RECT 69.500 139.815 70.370 139.985 ;
        RECT 69.500 139.745 69.670 139.815 ;
        RECT 69.790 139.565 69.990 139.595 ;
        RECT 68.310 139.205 68.775 139.535 ;
        RECT 69.160 139.265 69.990 139.565 ;
        RECT 69.160 139.035 69.330 139.265 ;
        RECT 67.970 138.865 68.755 139.035 ;
        RECT 68.925 138.865 69.330 139.035 ;
        RECT 69.510 138.585 69.880 139.085 ;
        RECT 70.200 139.035 70.370 139.815 ;
        RECT 70.540 139.455 70.710 140.155 ;
        RECT 70.880 139.625 71.120 140.220 ;
        RECT 70.540 139.235 71.065 139.455 ;
        RECT 71.290 139.305 71.460 140.410 ;
        RECT 71.235 139.175 71.460 139.305 ;
        RECT 71.630 139.215 71.910 140.165 ;
        RECT 71.235 139.035 71.405 139.175 ;
        RECT 70.200 138.865 70.875 139.035 ;
        RECT 71.070 138.865 71.405 139.035 ;
        RECT 71.575 138.585 71.825 139.045 ;
        RECT 72.080 138.845 72.265 140.965 ;
        RECT 72.435 140.635 72.765 141.135 ;
        RECT 72.935 140.465 73.105 140.965 ;
        RECT 72.440 140.295 73.105 140.465 ;
        RECT 72.440 139.305 72.670 140.295 ;
        RECT 74.470 140.165 74.860 140.340 ;
        RECT 75.345 140.335 75.675 141.135 ;
        RECT 75.845 140.345 76.380 140.965 ;
        RECT 72.840 139.475 73.190 140.125 ;
        RECT 74.470 139.995 75.895 140.165 ;
        RECT 72.440 139.135 73.105 139.305 ;
        RECT 74.345 139.265 74.700 139.825 ;
        RECT 72.435 138.585 72.765 138.965 ;
        RECT 72.935 138.845 73.105 139.135 ;
        RECT 74.870 139.095 75.040 139.995 ;
        RECT 75.210 139.265 75.475 139.825 ;
        RECT 75.725 139.495 75.895 139.995 ;
        RECT 76.065 139.325 76.380 140.345 ;
        RECT 76.585 139.970 76.875 141.135 ;
        RECT 77.045 139.995 77.430 140.965 ;
        RECT 77.600 140.675 77.925 141.135 ;
        RECT 78.445 140.505 78.725 140.965 ;
        RECT 77.600 140.285 78.725 140.505 ;
        RECT 74.450 138.585 74.690 139.095 ;
        RECT 74.870 138.765 75.150 139.095 ;
        RECT 75.380 138.585 75.595 139.095 ;
        RECT 75.765 138.755 76.380 139.325 ;
        RECT 77.045 139.325 77.325 139.995 ;
        RECT 77.600 139.825 78.050 140.285 ;
        RECT 78.915 140.115 79.315 140.965 ;
        RECT 79.715 140.675 79.985 141.135 ;
        RECT 80.155 140.505 80.440 140.965 ;
        RECT 77.495 139.495 78.050 139.825 ;
        RECT 78.220 139.555 79.315 140.115 ;
        RECT 77.600 139.385 78.050 139.495 ;
        RECT 76.585 138.585 76.875 139.310 ;
        RECT 77.045 138.755 77.430 139.325 ;
        RECT 77.600 139.215 78.725 139.385 ;
        RECT 77.600 138.585 77.925 139.045 ;
        RECT 78.445 138.755 78.725 139.215 ;
        RECT 78.915 138.755 79.315 139.555 ;
        RECT 79.485 140.285 80.440 140.505 ;
        RECT 79.485 139.385 79.695 140.285 ;
        RECT 79.865 139.555 80.555 140.115 ;
        RECT 80.725 139.995 81.110 140.965 ;
        RECT 81.280 140.675 81.605 141.135 ;
        RECT 82.125 140.505 82.405 140.965 ;
        RECT 81.280 140.285 82.405 140.505 ;
        RECT 79.485 139.215 80.440 139.385 ;
        RECT 79.715 138.585 79.985 139.045 ;
        RECT 80.155 138.755 80.440 139.215 ;
        RECT 80.725 139.325 81.005 139.995 ;
        RECT 81.280 139.825 81.730 140.285 ;
        RECT 82.595 140.115 82.995 140.965 ;
        RECT 83.395 140.675 83.665 141.135 ;
        RECT 83.835 140.505 84.120 140.965 ;
        RECT 81.175 139.495 81.730 139.825 ;
        RECT 81.900 139.555 82.995 140.115 ;
        RECT 81.280 139.385 81.730 139.495 ;
        RECT 80.725 138.755 81.110 139.325 ;
        RECT 81.280 139.215 82.405 139.385 ;
        RECT 81.280 138.585 81.605 139.045 ;
        RECT 82.125 138.755 82.405 139.215 ;
        RECT 82.595 138.755 82.995 139.555 ;
        RECT 83.165 140.285 84.120 140.505 ;
        RECT 83.165 139.385 83.375 140.285 ;
        RECT 83.545 139.555 84.235 140.115 ;
        RECT 84.405 139.995 84.745 140.965 ;
        RECT 84.915 139.995 85.085 141.135 ;
        RECT 85.355 140.335 85.605 141.135 ;
        RECT 86.250 140.165 86.580 140.965 ;
        RECT 86.880 140.335 87.210 141.135 ;
        RECT 87.380 140.165 87.710 140.965 ;
        RECT 85.275 139.995 87.710 140.165 ;
        RECT 88.545 140.045 89.755 141.135 ;
        RECT 100.140 140.890 100.810 144.150 ;
        RECT 101.480 143.580 105.520 143.750 ;
        RECT 101.140 141.520 101.310 143.520 ;
        RECT 105.690 141.520 105.860 143.520 ;
        RECT 101.480 141.290 105.520 141.460 ;
        RECT 106.200 140.890 106.370 144.150 ;
        RECT 100.140 140.720 106.370 140.890 ;
        RECT 84.405 139.385 84.580 139.995 ;
        RECT 85.275 139.745 85.445 139.995 ;
        RECT 84.750 139.575 85.445 139.745 ;
        RECT 85.620 139.575 86.040 139.775 ;
        RECT 86.210 139.575 86.540 139.775 ;
        RECT 86.710 139.575 87.040 139.775 ;
        RECT 83.165 139.215 84.120 139.385 ;
        RECT 83.395 138.585 83.665 139.045 ;
        RECT 83.835 138.755 84.120 139.215 ;
        RECT 84.405 138.755 84.745 139.385 ;
        RECT 84.915 138.585 85.165 139.385 ;
        RECT 85.355 139.235 86.580 139.405 ;
        RECT 85.355 138.755 85.685 139.235 ;
        RECT 85.855 138.585 86.080 139.045 ;
        RECT 86.250 138.755 86.580 139.235 ;
        RECT 87.210 139.365 87.380 139.995 ;
        RECT 87.565 139.575 87.915 139.825 ;
        RECT 88.545 139.505 89.065 140.045 ;
        RECT 87.210 138.755 87.710 139.365 ;
        RECT 89.235 139.335 89.755 139.875 ;
        RECT 88.545 138.585 89.755 139.335 ;
        RECT 12.100 138.415 89.840 138.585 ;
        RECT 12.185 137.665 13.395 138.415 ;
        RECT 13.565 137.870 18.910 138.415 ;
        RECT 12.185 137.125 12.705 137.665 ;
        RECT 12.875 136.955 13.395 137.495 ;
        RECT 15.150 137.040 15.490 137.870 ;
        RECT 19.085 137.645 21.675 138.415 ;
        RECT 22.305 137.765 22.565 138.245 ;
        RECT 22.735 137.875 22.985 138.415 ;
        RECT 12.185 135.865 13.395 136.955 ;
        RECT 16.970 136.300 17.320 137.550 ;
        RECT 19.085 137.125 20.295 137.645 ;
        RECT 20.465 136.955 21.675 137.475 ;
        RECT 13.565 135.865 18.910 136.300 ;
        RECT 19.085 135.865 21.675 136.955 ;
        RECT 22.305 136.735 22.475 137.765 ;
        RECT 23.155 137.735 23.375 138.195 ;
        RECT 23.125 137.710 23.375 137.735 ;
        RECT 22.645 137.115 22.875 137.510 ;
        RECT 23.045 137.285 23.375 137.710 ;
        RECT 23.545 138.035 24.435 138.205 ;
        RECT 23.545 137.310 23.715 138.035 ;
        RECT 23.885 137.480 24.435 137.865 ;
        RECT 24.605 137.695 24.945 138.205 ;
        RECT 23.545 137.240 24.435 137.310 ;
        RECT 23.540 137.215 24.435 137.240 ;
        RECT 23.530 137.200 24.435 137.215 ;
        RECT 23.525 137.185 24.435 137.200 ;
        RECT 23.515 137.180 24.435 137.185 ;
        RECT 23.510 137.170 24.435 137.180 ;
        RECT 23.505 137.160 24.435 137.170 ;
        RECT 23.495 137.155 24.435 137.160 ;
        RECT 23.485 137.145 24.435 137.155 ;
        RECT 23.475 137.140 24.435 137.145 ;
        RECT 23.475 137.135 23.810 137.140 ;
        RECT 23.460 137.130 23.810 137.135 ;
        RECT 23.445 137.120 23.810 137.130 ;
        RECT 23.420 137.115 23.810 137.120 ;
        RECT 22.645 137.110 23.810 137.115 ;
        RECT 22.645 137.075 23.780 137.110 ;
        RECT 22.645 137.050 23.745 137.075 ;
        RECT 22.645 137.020 23.715 137.050 ;
        RECT 22.645 136.990 23.695 137.020 ;
        RECT 22.645 136.960 23.675 136.990 ;
        RECT 22.645 136.950 23.605 136.960 ;
        RECT 22.645 136.940 23.580 136.950 ;
        RECT 22.645 136.925 23.560 136.940 ;
        RECT 22.645 136.910 23.540 136.925 ;
        RECT 22.750 136.900 23.535 136.910 ;
        RECT 22.750 136.865 23.520 136.900 ;
        RECT 22.305 136.035 22.580 136.735 ;
        RECT 22.750 136.615 23.505 136.865 ;
        RECT 23.675 136.545 24.005 136.790 ;
        RECT 24.175 136.690 24.435 137.140 ;
        RECT 23.820 136.520 24.005 136.545 ;
        RECT 23.820 136.420 24.435 136.520 ;
        RECT 22.750 135.865 23.005 136.410 ;
        RECT 23.175 136.035 23.655 136.375 ;
        RECT 23.830 135.865 24.435 136.420 ;
        RECT 24.605 136.295 24.865 137.695 ;
        RECT 25.115 137.615 25.385 138.415 ;
        RECT 25.040 137.175 25.370 137.425 ;
        RECT 25.565 137.175 25.845 138.145 ;
        RECT 26.025 137.175 26.325 138.145 ;
        RECT 26.505 137.175 26.855 138.140 ;
        RECT 27.075 137.915 27.570 138.245 ;
        RECT 25.055 137.005 25.370 137.175 ;
        RECT 27.075 137.005 27.245 137.915 ;
        RECT 25.055 136.835 27.245 137.005 ;
        RECT 24.605 136.035 24.945 136.295 ;
        RECT 25.115 135.865 25.445 136.665 ;
        RECT 25.910 136.035 26.160 136.835 ;
        RECT 26.345 135.865 26.675 136.585 ;
        RECT 26.895 136.035 27.145 136.835 ;
        RECT 27.415 136.425 27.655 137.735 ;
        RECT 27.825 137.580 28.115 138.415 ;
        RECT 28.285 138.015 29.240 138.185 ;
        RECT 29.655 138.025 29.985 138.415 ;
        RECT 28.285 137.135 28.455 138.015 ;
        RECT 30.155 137.845 30.325 138.165 ;
        RECT 30.495 138.025 30.825 138.415 ;
        RECT 28.625 137.675 30.875 137.845 ;
        RECT 28.625 137.175 28.855 137.675 ;
        RECT 29.025 137.255 29.400 137.425 ;
        RECT 27.825 136.965 28.455 137.135 ;
        RECT 29.230 137.055 29.400 137.255 ;
        RECT 29.570 137.225 30.120 137.425 ;
        RECT 30.290 137.055 30.535 137.505 ;
        RECT 27.315 135.865 27.650 136.245 ;
        RECT 27.825 136.035 28.145 136.965 ;
        RECT 29.230 136.885 30.535 137.055 ;
        RECT 30.705 136.715 30.875 137.675 ;
        RECT 31.045 137.665 32.255 138.415 ;
        RECT 32.425 138.035 33.315 138.205 ;
        RECT 31.045 137.125 31.565 137.665 ;
        RECT 31.735 136.955 32.255 137.495 ;
        RECT 32.425 137.480 32.975 137.865 ;
        RECT 33.145 137.310 33.315 138.035 ;
        RECT 28.325 136.545 29.565 136.715 ;
        RECT 28.325 136.035 28.725 136.545 ;
        RECT 28.895 135.865 29.065 136.375 ;
        RECT 29.235 136.035 29.565 136.545 ;
        RECT 29.735 135.865 29.905 136.715 ;
        RECT 30.495 136.035 30.875 136.715 ;
        RECT 31.045 135.865 32.255 136.955 ;
        RECT 32.425 137.240 33.315 137.310 ;
        RECT 33.485 137.710 33.705 138.195 ;
        RECT 33.875 137.875 34.125 138.415 ;
        RECT 34.295 137.765 34.555 138.245 ;
        RECT 33.485 137.285 33.815 137.710 ;
        RECT 32.425 137.215 33.320 137.240 ;
        RECT 32.425 137.200 33.330 137.215 ;
        RECT 32.425 137.185 33.335 137.200 ;
        RECT 32.425 137.180 33.345 137.185 ;
        RECT 32.425 137.170 33.350 137.180 ;
        RECT 32.425 137.160 33.355 137.170 ;
        RECT 32.425 137.155 33.365 137.160 ;
        RECT 32.425 137.145 33.375 137.155 ;
        RECT 32.425 137.140 33.385 137.145 ;
        RECT 32.425 136.690 32.685 137.140 ;
        RECT 33.050 137.135 33.385 137.140 ;
        RECT 33.050 137.130 33.400 137.135 ;
        RECT 33.050 137.120 33.415 137.130 ;
        RECT 33.050 137.115 33.440 137.120 ;
        RECT 33.985 137.115 34.215 137.510 ;
        RECT 33.050 137.110 34.215 137.115 ;
        RECT 33.080 137.075 34.215 137.110 ;
        RECT 33.115 137.050 34.215 137.075 ;
        RECT 33.145 137.020 34.215 137.050 ;
        RECT 33.165 136.990 34.215 137.020 ;
        RECT 33.185 136.960 34.215 136.990 ;
        RECT 33.255 136.950 34.215 136.960 ;
        RECT 33.280 136.940 34.215 136.950 ;
        RECT 33.300 136.925 34.215 136.940 ;
        RECT 33.320 136.910 34.215 136.925 ;
        RECT 33.325 136.900 34.110 136.910 ;
        RECT 33.340 136.865 34.110 136.900 ;
        RECT 32.855 136.545 33.185 136.790 ;
        RECT 33.355 136.615 34.110 136.865 ;
        RECT 34.385 136.735 34.555 137.765 ;
        RECT 34.745 137.605 34.985 138.415 ;
        RECT 35.155 137.605 35.485 138.245 ;
        RECT 35.655 137.605 35.925 138.415 ;
        RECT 34.725 137.175 35.075 137.425 ;
        RECT 35.245 137.005 35.415 137.605 ;
        RECT 36.625 137.595 36.835 138.415 ;
        RECT 37.005 137.615 37.335 138.245 ;
        RECT 35.585 137.175 35.935 137.425 ;
        RECT 37.005 137.015 37.255 137.615 ;
        RECT 37.505 137.595 37.735 138.415 ;
        RECT 37.945 137.690 38.235 138.415 ;
        RECT 38.980 137.785 39.265 138.245 ;
        RECT 39.435 137.955 39.705 138.415 ;
        RECT 38.980 137.615 39.935 137.785 ;
        RECT 37.425 137.175 37.755 137.425 ;
        RECT 32.855 136.520 33.040 136.545 ;
        RECT 32.425 136.420 33.040 136.520 ;
        RECT 32.425 135.865 33.030 136.420 ;
        RECT 33.205 136.035 33.685 136.375 ;
        RECT 33.855 135.865 34.110 136.410 ;
        RECT 34.280 136.035 34.555 136.735 ;
        RECT 34.735 136.835 35.415 137.005 ;
        RECT 34.735 136.050 35.065 136.835 ;
        RECT 35.595 135.865 35.925 137.005 ;
        RECT 36.625 135.865 36.835 137.005 ;
        RECT 37.005 136.035 37.335 137.015 ;
        RECT 37.505 135.865 37.735 137.005 ;
        RECT 37.945 135.865 38.235 137.030 ;
        RECT 38.865 136.885 39.555 137.445 ;
        RECT 39.725 136.715 39.935 137.615 ;
        RECT 38.980 136.495 39.935 136.715 ;
        RECT 40.105 137.445 40.505 138.245 ;
        RECT 40.695 137.785 40.975 138.245 ;
        RECT 41.495 137.955 41.820 138.415 ;
        RECT 40.695 137.615 41.820 137.785 ;
        RECT 41.990 137.675 42.375 138.245 ;
        RECT 42.605 137.955 42.850 138.415 ;
        RECT 41.370 137.505 41.820 137.615 ;
        RECT 40.105 136.885 41.200 137.445 ;
        RECT 41.370 137.175 41.925 137.505 ;
        RECT 38.980 136.035 39.265 136.495 ;
        RECT 39.435 135.865 39.705 136.325 ;
        RECT 40.105 136.035 40.505 136.885 ;
        RECT 41.370 136.715 41.820 137.175 ;
        RECT 42.095 137.005 42.375 137.675 ;
        RECT 42.545 137.175 42.860 137.785 ;
        RECT 43.030 137.425 43.280 138.235 ;
        RECT 43.450 137.890 43.710 138.415 ;
        RECT 43.880 137.765 44.140 138.220 ;
        RECT 44.310 137.935 44.570 138.415 ;
        RECT 44.740 137.765 45.000 138.220 ;
        RECT 45.170 137.935 45.430 138.415 ;
        RECT 45.600 137.765 45.860 138.220 ;
        RECT 46.030 137.935 46.290 138.415 ;
        RECT 46.460 137.765 46.720 138.220 ;
        RECT 46.890 137.935 47.190 138.415 ;
        RECT 47.695 137.865 47.865 138.155 ;
        RECT 48.035 138.035 48.365 138.415 ;
        RECT 43.880 137.595 47.190 137.765 ;
        RECT 47.695 137.695 48.360 137.865 ;
        RECT 43.030 137.175 46.050 137.425 ;
        RECT 40.695 136.495 41.820 136.715 ;
        RECT 40.695 136.035 40.975 136.495 ;
        RECT 41.495 135.865 41.820 136.325 ;
        RECT 41.990 136.035 42.375 137.005 ;
        RECT 42.555 135.865 42.850 136.975 ;
        RECT 43.030 136.040 43.280 137.175 ;
        RECT 46.220 137.005 47.190 137.595 ;
        RECT 43.450 135.865 43.710 136.975 ;
        RECT 43.880 136.765 47.190 137.005 ;
        RECT 47.610 136.875 47.960 137.525 ;
        RECT 43.880 136.040 44.140 136.765 ;
        RECT 44.310 135.865 44.570 136.595 ;
        RECT 44.740 136.040 45.000 136.765 ;
        RECT 45.170 135.865 45.430 136.595 ;
        RECT 45.600 136.040 45.860 136.765 ;
        RECT 46.030 135.865 46.290 136.595 ;
        RECT 46.460 136.040 46.720 136.765 ;
        RECT 48.130 136.705 48.360 137.695 ;
        RECT 46.890 135.865 47.185 136.595 ;
        RECT 47.695 136.535 48.360 136.705 ;
        RECT 47.695 136.035 47.865 136.535 ;
        RECT 48.035 135.865 48.365 136.365 ;
        RECT 48.535 136.035 48.720 138.155 ;
        RECT 48.975 137.955 49.225 138.415 ;
        RECT 49.395 137.965 49.730 138.135 ;
        RECT 49.925 137.965 50.600 138.135 ;
        RECT 49.395 137.825 49.565 137.965 ;
        RECT 48.890 136.835 49.170 137.785 ;
        RECT 49.340 137.695 49.565 137.825 ;
        RECT 49.340 136.590 49.510 137.695 ;
        RECT 49.735 137.545 50.260 137.765 ;
        RECT 49.680 136.780 49.920 137.375 ;
        RECT 50.090 136.845 50.260 137.545 ;
        RECT 50.430 137.185 50.600 137.965 ;
        RECT 50.920 137.915 51.290 138.415 ;
        RECT 51.470 137.965 51.875 138.135 ;
        RECT 52.045 137.965 52.830 138.135 ;
        RECT 51.470 137.735 51.640 137.965 ;
        RECT 50.810 137.435 51.640 137.735 ;
        RECT 52.025 137.465 52.490 137.795 ;
        RECT 50.810 137.405 51.010 137.435 ;
        RECT 51.130 137.185 51.300 137.255 ;
        RECT 50.430 137.015 51.300 137.185 ;
        RECT 50.790 136.925 51.300 137.015 ;
        RECT 49.340 136.460 49.645 136.590 ;
        RECT 50.090 136.480 50.620 136.845 ;
        RECT 48.960 135.865 49.225 136.325 ;
        RECT 49.395 136.035 49.645 136.460 ;
        RECT 50.790 136.310 50.960 136.925 ;
        RECT 49.855 136.140 50.960 136.310 ;
        RECT 51.130 135.865 51.300 136.665 ;
        RECT 51.470 136.365 51.640 137.435 ;
        RECT 51.810 136.535 52.000 137.255 ;
        RECT 52.170 136.505 52.490 137.465 ;
        RECT 52.660 137.505 52.830 137.965 ;
        RECT 53.105 137.885 53.315 138.415 ;
        RECT 53.575 137.675 53.905 138.200 ;
        RECT 54.075 137.805 54.245 138.415 ;
        RECT 54.415 137.760 54.745 138.195 ;
        RECT 54.415 137.675 54.795 137.760 ;
        RECT 53.705 137.505 53.905 137.675 ;
        RECT 54.570 137.635 54.795 137.675 ;
        RECT 52.660 137.175 53.535 137.505 ;
        RECT 53.705 137.175 54.455 137.505 ;
        RECT 51.470 136.035 51.720 136.365 ;
        RECT 52.660 136.335 52.830 137.175 ;
        RECT 53.705 136.970 53.895 137.175 ;
        RECT 54.625 137.055 54.795 137.635 ;
        RECT 54.580 137.005 54.795 137.055 ;
        RECT 53.000 136.595 53.895 136.970 ;
        RECT 54.405 136.925 54.795 137.005 ;
        RECT 54.970 137.675 55.225 138.245 ;
        RECT 55.395 138.015 55.725 138.415 ;
        RECT 56.150 137.880 56.680 138.245 ;
        RECT 56.150 137.845 56.325 137.880 ;
        RECT 55.395 137.675 56.325 137.845 ;
        RECT 56.870 137.735 57.145 138.245 ;
        RECT 54.970 137.005 55.140 137.675 ;
        RECT 55.395 137.505 55.565 137.675 ;
        RECT 55.310 137.175 55.565 137.505 ;
        RECT 55.790 137.175 55.985 137.505 ;
        RECT 51.945 136.165 52.830 136.335 ;
        RECT 53.010 135.865 53.325 136.365 ;
        RECT 53.555 136.035 53.895 136.595 ;
        RECT 54.065 135.865 54.235 136.875 ;
        RECT 54.405 136.080 54.735 136.925 ;
        RECT 54.970 136.035 55.305 137.005 ;
        RECT 55.475 135.865 55.645 137.005 ;
        RECT 55.815 136.205 55.985 137.175 ;
        RECT 56.155 136.545 56.325 137.675 ;
        RECT 56.495 136.885 56.665 137.685 ;
        RECT 56.865 137.565 57.145 137.735 ;
        RECT 56.870 137.085 57.145 137.565 ;
        RECT 57.315 136.885 57.505 138.245 ;
        RECT 57.685 137.880 58.195 138.415 ;
        RECT 58.415 137.605 58.660 138.210 ;
        RECT 59.570 137.675 59.825 138.245 ;
        RECT 59.995 138.015 60.325 138.415 ;
        RECT 60.750 137.880 61.280 138.245 ;
        RECT 61.470 138.075 61.745 138.245 ;
        RECT 61.465 137.905 61.745 138.075 ;
        RECT 60.750 137.845 60.925 137.880 ;
        RECT 59.995 137.675 60.925 137.845 ;
        RECT 57.705 137.435 58.935 137.605 ;
        RECT 56.495 136.715 57.505 136.885 ;
        RECT 57.675 136.870 58.425 137.060 ;
        RECT 56.155 136.375 57.280 136.545 ;
        RECT 57.675 136.205 57.845 136.870 ;
        RECT 58.595 136.625 58.935 137.435 ;
        RECT 55.815 136.035 57.845 136.205 ;
        RECT 58.015 135.865 58.185 136.625 ;
        RECT 58.420 136.215 58.935 136.625 ;
        RECT 59.570 137.005 59.740 137.675 ;
        RECT 59.995 137.505 60.165 137.675 ;
        RECT 59.910 137.175 60.165 137.505 ;
        RECT 60.390 137.175 60.585 137.505 ;
        RECT 59.570 136.035 59.905 137.005 ;
        RECT 60.075 135.865 60.245 137.005 ;
        RECT 60.415 136.205 60.585 137.175 ;
        RECT 60.755 136.545 60.925 137.675 ;
        RECT 61.095 136.885 61.265 137.685 ;
        RECT 61.470 137.085 61.745 137.905 ;
        RECT 61.915 136.885 62.105 138.245 ;
        RECT 62.285 137.880 62.795 138.415 ;
        RECT 63.015 137.605 63.260 138.210 ;
        RECT 63.705 137.690 63.995 138.415 ;
        RECT 64.165 137.665 65.375 138.415 ;
        RECT 65.595 137.760 65.925 138.195 ;
        RECT 66.095 137.805 66.265 138.415 ;
        RECT 65.545 137.675 65.925 137.760 ;
        RECT 66.435 137.675 66.765 138.200 ;
        RECT 67.025 137.885 67.235 138.415 ;
        RECT 67.510 137.965 68.295 138.135 ;
        RECT 68.465 137.965 68.870 138.135 ;
        RECT 62.305 137.435 63.535 137.605 ;
        RECT 61.095 136.715 62.105 136.885 ;
        RECT 62.275 136.870 63.025 137.060 ;
        RECT 60.755 136.375 61.880 136.545 ;
        RECT 62.275 136.205 62.445 136.870 ;
        RECT 63.195 136.625 63.535 137.435 ;
        RECT 64.165 137.125 64.685 137.665 ;
        RECT 65.545 137.635 65.770 137.675 ;
        RECT 60.415 136.035 62.445 136.205 ;
        RECT 62.615 135.865 62.785 136.625 ;
        RECT 63.020 136.215 63.535 136.625 ;
        RECT 63.705 135.865 63.995 137.030 ;
        RECT 64.855 136.955 65.375 137.495 ;
        RECT 64.165 135.865 65.375 136.955 ;
        RECT 65.545 137.055 65.715 137.635 ;
        RECT 66.435 137.505 66.635 137.675 ;
        RECT 67.510 137.505 67.680 137.965 ;
        RECT 65.885 137.175 66.635 137.505 ;
        RECT 66.805 137.175 67.680 137.505 ;
        RECT 65.545 137.005 65.760 137.055 ;
        RECT 65.545 136.925 65.935 137.005 ;
        RECT 65.605 136.080 65.935 136.925 ;
        RECT 66.445 136.970 66.635 137.175 ;
        RECT 66.105 135.865 66.275 136.875 ;
        RECT 66.445 136.595 67.340 136.970 ;
        RECT 66.445 136.035 66.785 136.595 ;
        RECT 67.015 135.865 67.330 136.365 ;
        RECT 67.510 136.335 67.680 137.175 ;
        RECT 67.850 137.465 68.315 137.795 ;
        RECT 68.700 137.735 68.870 137.965 ;
        RECT 69.050 137.915 69.420 138.415 ;
        RECT 69.740 137.965 70.415 138.135 ;
        RECT 70.610 137.965 70.945 138.135 ;
        RECT 67.850 136.505 68.170 137.465 ;
        RECT 68.700 137.435 69.530 137.735 ;
        RECT 68.340 136.535 68.530 137.255 ;
        RECT 68.700 136.365 68.870 137.435 ;
        RECT 69.330 137.405 69.530 137.435 ;
        RECT 69.040 137.185 69.210 137.255 ;
        RECT 69.740 137.185 69.910 137.965 ;
        RECT 70.775 137.825 70.945 137.965 ;
        RECT 71.115 137.955 71.365 138.415 ;
        RECT 69.040 137.015 69.910 137.185 ;
        RECT 70.080 137.545 70.605 137.765 ;
        RECT 70.775 137.695 71.000 137.825 ;
        RECT 69.040 136.925 69.550 137.015 ;
        RECT 67.510 136.165 68.395 136.335 ;
        RECT 68.620 136.035 68.870 136.365 ;
        RECT 69.040 135.865 69.210 136.665 ;
        RECT 69.380 136.310 69.550 136.925 ;
        RECT 70.080 136.845 70.250 137.545 ;
        RECT 69.720 136.480 70.250 136.845 ;
        RECT 70.420 136.780 70.660 137.375 ;
        RECT 70.830 136.590 71.000 137.695 ;
        RECT 71.170 136.835 71.450 137.785 ;
        RECT 70.695 136.460 71.000 136.590 ;
        RECT 69.380 136.140 70.485 136.310 ;
        RECT 70.695 136.035 70.945 136.460 ;
        RECT 71.115 135.865 71.380 136.325 ;
        RECT 71.620 136.035 71.805 138.155 ;
        RECT 71.975 138.035 72.305 138.415 ;
        RECT 72.475 137.865 72.645 138.155 ;
        RECT 72.965 137.955 73.210 138.415 ;
        RECT 71.980 137.695 72.645 137.865 ;
        RECT 71.980 136.705 72.210 137.695 ;
        RECT 72.380 136.875 72.730 137.525 ;
        RECT 72.905 137.175 73.220 137.785 ;
        RECT 73.390 137.425 73.640 138.235 ;
        RECT 73.810 137.890 74.070 138.415 ;
        RECT 74.240 137.765 74.500 138.220 ;
        RECT 74.670 137.935 74.930 138.415 ;
        RECT 75.100 137.765 75.360 138.220 ;
        RECT 75.530 137.935 75.790 138.415 ;
        RECT 75.960 137.765 76.220 138.220 ;
        RECT 76.390 137.935 76.650 138.415 ;
        RECT 76.820 137.765 77.080 138.220 ;
        RECT 77.250 137.935 77.550 138.415 ;
        RECT 74.240 137.595 77.550 137.765 ;
        RECT 73.390 137.175 76.410 137.425 ;
        RECT 71.980 136.535 72.645 136.705 ;
        RECT 71.975 135.865 72.305 136.365 ;
        RECT 72.475 136.035 72.645 136.535 ;
        RECT 72.915 135.865 73.210 136.975 ;
        RECT 73.390 136.040 73.640 137.175 ;
        RECT 76.580 137.005 77.550 137.595 ;
        RECT 73.810 135.865 74.070 136.975 ;
        RECT 74.240 136.765 77.550 137.005 ;
        RECT 77.970 137.675 78.225 138.245 ;
        RECT 78.395 138.015 78.725 138.415 ;
        RECT 79.150 137.880 79.680 138.245 ;
        RECT 79.870 138.075 80.145 138.245 ;
        RECT 79.865 137.905 80.145 138.075 ;
        RECT 79.150 137.845 79.325 137.880 ;
        RECT 78.395 137.675 79.325 137.845 ;
        RECT 77.970 137.005 78.140 137.675 ;
        RECT 78.395 137.505 78.565 137.675 ;
        RECT 78.310 137.175 78.565 137.505 ;
        RECT 78.790 137.175 78.985 137.505 ;
        RECT 74.240 136.040 74.500 136.765 ;
        RECT 74.670 135.865 74.930 136.595 ;
        RECT 75.100 136.040 75.360 136.765 ;
        RECT 75.530 135.865 75.790 136.595 ;
        RECT 75.960 136.040 76.220 136.765 ;
        RECT 76.390 135.865 76.650 136.595 ;
        RECT 76.820 136.040 77.080 136.765 ;
        RECT 77.250 135.865 77.545 136.595 ;
        RECT 77.970 136.035 78.305 137.005 ;
        RECT 78.475 135.865 78.645 137.005 ;
        RECT 78.815 136.205 78.985 137.175 ;
        RECT 79.155 136.545 79.325 137.675 ;
        RECT 79.495 136.885 79.665 137.685 ;
        RECT 79.870 137.085 80.145 137.905 ;
        RECT 80.315 136.885 80.505 138.245 ;
        RECT 80.685 137.880 81.195 138.415 ;
        RECT 81.415 137.605 81.660 138.210 ;
        RECT 80.705 137.435 81.935 137.605 ;
        RECT 79.495 136.715 80.505 136.885 ;
        RECT 80.675 136.870 81.425 137.060 ;
        RECT 79.155 136.375 80.280 136.545 ;
        RECT 80.675 136.205 80.845 136.870 ;
        RECT 81.595 136.625 81.935 137.435 ;
        RECT 78.815 136.035 80.845 136.205 ;
        RECT 81.015 135.865 81.185 136.625 ;
        RECT 81.420 136.215 81.935 136.625 ;
        RECT 82.110 136.815 82.445 138.235 ;
        RECT 82.625 138.045 83.370 138.415 ;
        RECT 83.935 137.875 84.190 138.235 ;
        RECT 84.370 138.045 84.700 138.415 ;
        RECT 84.880 137.875 85.105 138.235 ;
        RECT 82.620 137.685 85.105 137.875 ;
        RECT 82.620 136.995 82.845 137.685 ;
        RECT 85.360 137.675 85.975 138.245 ;
        RECT 86.145 137.905 86.360 138.415 ;
        RECT 86.590 137.905 86.870 138.235 ;
        RECT 87.050 137.905 87.290 138.415 ;
        RECT 83.045 137.175 83.325 137.505 ;
        RECT 83.505 137.175 84.080 137.505 ;
        RECT 84.260 137.175 84.695 137.505 ;
        RECT 84.875 137.175 85.145 137.505 ;
        RECT 82.620 136.815 85.115 136.995 ;
        RECT 82.110 136.045 82.375 136.815 ;
        RECT 82.545 135.865 82.875 136.585 ;
        RECT 83.065 136.405 84.255 136.635 ;
        RECT 83.065 136.045 83.325 136.405 ;
        RECT 83.495 135.865 83.825 136.235 ;
        RECT 83.995 136.045 84.255 136.405 ;
        RECT 84.825 136.045 85.115 136.815 ;
        RECT 85.360 136.655 85.675 137.675 ;
        RECT 85.845 137.005 86.015 137.505 ;
        RECT 86.265 137.175 86.530 137.735 ;
        RECT 86.700 137.005 86.870 137.905 ;
        RECT 87.040 137.175 87.395 137.735 ;
        RECT 88.545 137.665 89.755 138.415 ;
        RECT 85.845 136.835 87.270 137.005 ;
        RECT 85.360 136.035 85.895 136.655 ;
        RECT 86.065 135.865 86.395 136.665 ;
        RECT 86.880 136.660 87.270 136.835 ;
        RECT 88.545 136.955 89.065 137.495 ;
        RECT 89.235 137.125 89.755 137.665 ;
        RECT 100.140 137.460 100.810 140.720 ;
        RECT 101.480 140.150 105.520 140.320 ;
        RECT 101.140 138.090 101.310 140.090 ;
        RECT 105.690 138.090 105.860 140.090 ;
        RECT 101.480 137.860 105.520 138.030 ;
        RECT 106.200 137.460 106.370 140.720 ;
        RECT 100.140 137.450 106.370 137.460 ;
        RECT 107.960 146.720 117.790 146.760 ;
        RECT 120.510 146.740 126.250 146.750 ;
        RECT 107.960 146.590 118.590 146.720 ;
        RECT 107.960 144.330 108.130 146.590 ;
        RECT 108.855 146.020 116.895 146.190 ;
        RECT 108.470 144.960 108.640 145.960 ;
        RECT 117.110 144.960 117.280 145.960 ;
        RECT 108.855 144.730 116.895 144.900 ;
        RECT 117.620 144.330 118.590 146.590 ;
        RECT 107.960 144.160 118.590 144.330 ;
        RECT 107.960 140.900 108.130 144.160 ;
        RECT 108.855 143.590 116.895 143.760 ;
        RECT 108.470 141.530 108.640 143.530 ;
        RECT 117.110 141.530 117.280 143.530 ;
        RECT 108.855 141.300 116.895 141.470 ;
        RECT 117.620 140.900 118.590 144.160 ;
        RECT 107.960 140.730 118.590 140.900 ;
        RECT 107.960 137.470 108.130 140.730 ;
        RECT 108.855 140.160 116.895 140.330 ;
        RECT 108.470 138.100 108.640 140.100 ;
        RECT 117.110 138.100 117.280 140.100 ;
        RECT 108.855 137.870 116.895 138.040 ;
        RECT 117.620 137.470 118.590 140.730 ;
        RECT 100.140 137.350 106.380 137.450 ;
        RECT 88.545 135.865 89.755 136.955 ;
        RECT 100.130 136.790 106.380 137.350 ;
        RECT 100.130 136.770 105.300 136.790 ;
        RECT 100.130 136.700 104.120 136.770 ;
        RECT 12.100 135.695 89.840 135.865 ;
        RECT 12.185 134.605 13.395 135.695 ;
        RECT 12.185 133.895 12.705 134.435 ;
        RECT 12.875 134.065 13.395 134.605 ;
        RECT 13.655 134.765 13.825 135.525 ;
        RECT 14.005 134.935 14.335 135.695 ;
        RECT 13.655 134.595 14.320 134.765 ;
        RECT 14.505 134.620 14.775 135.525 ;
        RECT 14.945 135.260 20.290 135.695 ;
        RECT 14.150 134.450 14.320 134.595 ;
        RECT 13.585 134.045 13.915 134.415 ;
        RECT 14.150 134.120 14.435 134.450 ;
        RECT 12.185 133.145 13.395 133.895 ;
        RECT 14.150 133.865 14.320 134.120 ;
        RECT 13.655 133.695 14.320 133.865 ;
        RECT 14.605 133.820 14.775 134.620 ;
        RECT 13.655 133.315 13.825 133.695 ;
        RECT 14.005 133.145 14.335 133.525 ;
        RECT 14.515 133.315 14.775 133.820 ;
        RECT 16.530 133.690 16.870 134.520 ;
        RECT 18.350 134.010 18.700 135.260 ;
        RECT 20.465 134.605 23.975 135.695 ;
        RECT 20.465 133.915 22.115 134.435 ;
        RECT 22.285 134.085 23.975 134.605 ;
        RECT 25.065 134.530 25.355 135.695 ;
        RECT 25.525 135.260 30.870 135.695 ;
        RECT 14.945 133.145 20.290 133.690 ;
        RECT 20.465 133.145 23.975 133.915 ;
        RECT 25.065 133.145 25.355 133.870 ;
        RECT 27.110 133.690 27.450 134.520 ;
        RECT 28.930 134.010 29.280 135.260 ;
        RECT 31.045 134.605 33.635 135.695 ;
        RECT 34.515 134.965 34.810 135.695 ;
        RECT 34.980 134.795 35.240 135.520 ;
        RECT 35.410 134.965 35.670 135.695 ;
        RECT 35.840 134.795 36.100 135.520 ;
        RECT 36.270 134.965 36.530 135.695 ;
        RECT 36.700 134.795 36.960 135.520 ;
        RECT 37.130 134.965 37.390 135.695 ;
        RECT 37.560 134.795 37.820 135.520 ;
        RECT 31.045 133.915 32.255 134.435 ;
        RECT 32.425 134.085 33.635 134.605 ;
        RECT 34.510 134.555 37.820 134.795 ;
        RECT 37.990 134.585 38.250 135.695 ;
        RECT 34.510 133.965 35.480 134.555 ;
        RECT 38.420 134.385 38.670 135.520 ;
        RECT 38.850 134.585 39.145 135.695 ;
        RECT 39.785 135.105 40.485 135.525 ;
        RECT 40.685 135.335 41.015 135.695 ;
        RECT 41.185 135.105 41.515 135.505 ;
        RECT 39.785 134.875 41.515 135.105 ;
        RECT 35.650 134.135 38.670 134.385 ;
        RECT 25.525 133.145 30.870 133.690 ;
        RECT 31.045 133.145 33.635 133.915 ;
        RECT 34.510 133.795 37.820 133.965 ;
        RECT 34.510 133.145 34.810 133.625 ;
        RECT 34.980 133.340 35.240 133.795 ;
        RECT 35.410 133.145 35.670 133.625 ;
        RECT 35.840 133.340 36.100 133.795 ;
        RECT 36.270 133.145 36.530 133.625 ;
        RECT 36.700 133.340 36.960 133.795 ;
        RECT 37.130 133.145 37.390 133.625 ;
        RECT 37.560 133.340 37.820 133.795 ;
        RECT 37.990 133.145 38.250 133.670 ;
        RECT 38.420 133.325 38.670 134.135 ;
        RECT 38.840 133.775 39.155 134.385 ;
        RECT 39.785 133.905 39.990 134.875 ;
        RECT 40.160 134.135 40.490 134.675 ;
        RECT 40.665 134.385 40.990 134.675 ;
        RECT 41.185 134.655 41.515 134.875 ;
        RECT 41.685 134.385 41.855 135.355 ;
        RECT 42.035 134.635 42.365 135.695 ;
        RECT 43.075 134.690 43.330 135.495 ;
        RECT 43.500 134.860 43.760 135.695 ;
        RECT 43.930 134.690 44.190 135.495 ;
        RECT 44.360 134.860 44.615 135.695 ;
        RECT 43.075 134.520 44.675 134.690 ;
        RECT 40.665 134.055 41.160 134.385 ;
        RECT 41.480 134.055 41.855 134.385 ;
        RECT 42.065 134.055 42.375 134.385 ;
        RECT 43.005 134.125 44.225 134.350 ;
        RECT 44.395 133.955 44.675 134.520 ;
        RECT 38.850 133.145 39.095 133.605 ;
        RECT 39.785 133.315 40.495 133.905 ;
        RECT 41.005 133.675 42.365 133.885 ;
        RECT 41.005 133.315 41.335 133.675 ;
        RECT 41.535 133.145 41.865 133.505 ;
        RECT 42.035 133.315 42.365 133.675 ;
        RECT 43.945 133.785 44.675 133.955 ;
        RECT 44.850 134.555 45.125 135.525 ;
        RECT 45.335 134.895 45.615 135.695 ;
        RECT 45.785 135.185 46.975 135.475 ;
        RECT 45.785 134.845 46.955 135.015 ;
        RECT 45.785 134.725 45.955 134.845 ;
        RECT 45.295 134.555 45.955 134.725 ;
        RECT 44.850 133.820 45.020 134.555 ;
        RECT 45.295 134.385 45.465 134.555 ;
        RECT 46.265 134.385 46.460 134.675 ;
        RECT 46.630 134.555 46.955 134.845 ;
        RECT 47.145 134.555 47.530 135.525 ;
        RECT 47.700 135.235 48.025 135.695 ;
        RECT 48.545 135.065 48.825 135.525 ;
        RECT 47.700 134.845 48.825 135.065 ;
        RECT 45.190 134.055 45.465 134.385 ;
        RECT 45.635 134.055 46.460 134.385 ;
        RECT 46.630 134.055 46.975 134.385 ;
        RECT 45.295 133.885 45.465 134.055 ;
        RECT 47.145 133.885 47.425 134.555 ;
        RECT 47.700 134.385 48.150 134.845 ;
        RECT 49.015 134.675 49.415 135.525 ;
        RECT 49.815 135.235 50.085 135.695 ;
        RECT 50.255 135.065 50.540 135.525 ;
        RECT 47.595 134.055 48.150 134.385 ;
        RECT 48.320 134.115 49.415 134.675 ;
        RECT 47.700 133.945 48.150 134.055 ;
        RECT 43.480 133.145 43.775 133.670 ;
        RECT 43.945 133.340 44.170 133.785 ;
        RECT 44.340 133.145 44.670 133.615 ;
        RECT 44.850 133.475 45.125 133.820 ;
        RECT 45.295 133.715 46.960 133.885 ;
        RECT 45.315 133.145 45.695 133.545 ;
        RECT 45.865 133.365 46.035 133.715 ;
        RECT 46.205 133.145 46.535 133.545 ;
        RECT 46.705 133.365 46.960 133.715 ;
        RECT 47.145 133.315 47.530 133.885 ;
        RECT 47.700 133.775 48.825 133.945 ;
        RECT 47.700 133.145 48.025 133.605 ;
        RECT 48.545 133.315 48.825 133.775 ;
        RECT 49.015 133.315 49.415 134.115 ;
        RECT 49.585 134.845 50.540 135.065 ;
        RECT 49.585 133.945 49.795 134.845 ;
        RECT 49.965 134.115 50.655 134.675 ;
        RECT 50.825 134.530 51.115 135.695 ;
        RECT 51.750 134.555 52.085 135.525 ;
        RECT 52.255 134.555 52.425 135.695 ;
        RECT 52.595 135.355 54.625 135.525 ;
        RECT 49.585 133.775 50.540 133.945 ;
        RECT 51.750 133.885 51.920 134.555 ;
        RECT 52.595 134.385 52.765 135.355 ;
        RECT 52.090 134.055 52.345 134.385 ;
        RECT 52.570 134.055 52.765 134.385 ;
        RECT 52.935 135.015 54.060 135.185 ;
        RECT 52.175 133.885 52.345 134.055 ;
        RECT 52.935 133.885 53.105 135.015 ;
        RECT 49.815 133.145 50.085 133.605 ;
        RECT 50.255 133.315 50.540 133.775 ;
        RECT 50.825 133.145 51.115 133.870 ;
        RECT 51.750 133.315 52.005 133.885 ;
        RECT 52.175 133.715 53.105 133.885 ;
        RECT 53.275 134.675 54.285 134.845 ;
        RECT 53.275 133.875 53.445 134.675 ;
        RECT 53.650 133.995 53.925 134.475 ;
        RECT 53.645 133.825 53.925 133.995 ;
        RECT 52.930 133.680 53.105 133.715 ;
        RECT 52.175 133.145 52.505 133.545 ;
        RECT 52.930 133.315 53.460 133.680 ;
        RECT 53.650 133.315 53.925 133.825 ;
        RECT 54.095 133.315 54.285 134.675 ;
        RECT 54.455 134.690 54.625 135.355 ;
        RECT 54.795 134.935 54.965 135.695 ;
        RECT 55.200 134.935 55.715 135.345 ;
        RECT 54.455 134.500 55.205 134.690 ;
        RECT 55.375 134.125 55.715 134.935 ;
        RECT 54.485 133.955 55.715 134.125 ;
        RECT 55.885 134.555 56.270 135.525 ;
        RECT 56.440 135.235 56.765 135.695 ;
        RECT 57.285 135.065 57.565 135.525 ;
        RECT 56.440 134.845 57.565 135.065 ;
        RECT 54.465 133.145 54.975 133.680 ;
        RECT 55.195 133.350 55.440 133.955 ;
        RECT 55.885 133.885 56.165 134.555 ;
        RECT 56.440 134.385 56.890 134.845 ;
        RECT 57.755 134.675 58.155 135.525 ;
        RECT 58.555 135.235 58.825 135.695 ;
        RECT 58.995 135.065 59.280 135.525 ;
        RECT 56.335 134.055 56.890 134.385 ;
        RECT 57.060 134.115 58.155 134.675 ;
        RECT 56.440 133.945 56.890 134.055 ;
        RECT 55.885 133.315 56.270 133.885 ;
        RECT 56.440 133.775 57.565 133.945 ;
        RECT 56.440 133.145 56.765 133.605 ;
        RECT 57.285 133.315 57.565 133.775 ;
        RECT 57.755 133.315 58.155 134.115 ;
        RECT 58.325 134.845 59.280 135.065 ;
        RECT 58.325 133.945 58.535 134.845 ;
        RECT 58.705 134.115 59.395 134.675 ;
        RECT 59.565 134.605 61.235 135.695 ;
        RECT 58.325 133.775 59.280 133.945 ;
        RECT 58.555 133.145 58.825 133.605 ;
        RECT 58.995 133.315 59.280 133.775 ;
        RECT 59.565 133.915 60.315 134.435 ;
        RECT 60.485 134.085 61.235 134.605 ;
        RECT 61.410 134.545 61.670 135.695 ;
        RECT 61.845 134.620 62.100 135.525 ;
        RECT 62.270 134.935 62.600 135.695 ;
        RECT 62.815 134.765 62.985 135.525 ;
        RECT 63.360 135.065 63.645 135.525 ;
        RECT 63.815 135.235 64.085 135.695 ;
        RECT 63.360 134.845 64.315 135.065 ;
        RECT 59.565 133.145 61.235 133.915 ;
        RECT 61.410 133.145 61.670 133.985 ;
        RECT 61.845 133.890 62.015 134.620 ;
        RECT 62.270 134.595 62.985 134.765 ;
        RECT 62.270 134.385 62.440 134.595 ;
        RECT 62.185 134.055 62.440 134.385 ;
        RECT 61.845 133.315 62.100 133.890 ;
        RECT 62.270 133.865 62.440 134.055 ;
        RECT 62.720 134.045 63.075 134.415 ;
        RECT 63.245 134.115 63.935 134.675 ;
        RECT 64.105 133.945 64.315 134.845 ;
        RECT 62.270 133.695 62.985 133.865 ;
        RECT 62.270 133.145 62.600 133.525 ;
        RECT 62.815 133.315 62.985 133.695 ;
        RECT 63.360 133.775 64.315 133.945 ;
        RECT 64.485 134.675 64.885 135.525 ;
        RECT 65.075 135.065 65.355 135.525 ;
        RECT 65.875 135.235 66.200 135.695 ;
        RECT 65.075 134.845 66.200 135.065 ;
        RECT 64.485 134.115 65.580 134.675 ;
        RECT 65.750 134.385 66.200 134.845 ;
        RECT 66.370 134.555 66.755 135.525 ;
        RECT 63.360 133.315 63.645 133.775 ;
        RECT 63.815 133.145 64.085 133.605 ;
        RECT 64.485 133.315 64.885 134.115 ;
        RECT 65.750 134.055 66.305 134.385 ;
        RECT 65.750 133.945 66.200 134.055 ;
        RECT 65.075 133.775 66.200 133.945 ;
        RECT 66.475 133.885 66.755 134.555 ;
        RECT 66.930 134.545 67.190 135.695 ;
        RECT 67.365 134.620 67.620 135.525 ;
        RECT 67.790 134.935 68.120 135.695 ;
        RECT 68.335 134.765 68.505 135.525 ;
        RECT 65.075 133.315 65.355 133.775 ;
        RECT 65.875 133.145 66.200 133.605 ;
        RECT 66.370 133.315 66.755 133.885 ;
        RECT 66.930 133.145 67.190 133.985 ;
        RECT 67.365 133.890 67.535 134.620 ;
        RECT 67.790 134.595 68.505 134.765 ;
        RECT 67.790 134.385 67.960 134.595 ;
        RECT 68.765 134.555 69.150 135.525 ;
        RECT 69.320 135.235 69.645 135.695 ;
        RECT 70.165 135.065 70.445 135.525 ;
        RECT 69.320 134.845 70.445 135.065 ;
        RECT 67.705 134.055 67.960 134.385 ;
        RECT 67.365 133.315 67.620 133.890 ;
        RECT 67.790 133.865 67.960 134.055 ;
        RECT 68.240 134.045 68.595 134.415 ;
        RECT 68.765 133.885 69.045 134.555 ;
        RECT 69.320 134.385 69.770 134.845 ;
        RECT 70.635 134.675 71.035 135.525 ;
        RECT 71.435 135.235 71.705 135.695 ;
        RECT 71.875 135.065 72.160 135.525 ;
        RECT 69.215 134.055 69.770 134.385 ;
        RECT 69.940 134.115 71.035 134.675 ;
        RECT 69.320 133.945 69.770 134.055 ;
        RECT 67.790 133.695 68.505 133.865 ;
        RECT 67.790 133.145 68.120 133.525 ;
        RECT 68.335 133.315 68.505 133.695 ;
        RECT 68.765 133.315 69.150 133.885 ;
        RECT 69.320 133.775 70.445 133.945 ;
        RECT 69.320 133.145 69.645 133.605 ;
        RECT 70.165 133.315 70.445 133.775 ;
        RECT 70.635 133.315 71.035 134.115 ;
        RECT 71.205 134.845 72.160 135.065 ;
        RECT 72.560 135.065 72.845 135.525 ;
        RECT 73.015 135.235 73.285 135.695 ;
        RECT 72.560 134.845 73.515 135.065 ;
        RECT 71.205 133.945 71.415 134.845 ;
        RECT 71.585 134.115 72.275 134.675 ;
        RECT 72.445 134.115 73.135 134.675 ;
        RECT 73.305 133.945 73.515 134.845 ;
        RECT 71.205 133.775 72.160 133.945 ;
        RECT 71.435 133.145 71.705 133.605 ;
        RECT 71.875 133.315 72.160 133.775 ;
        RECT 72.560 133.775 73.515 133.945 ;
        RECT 73.685 134.675 74.085 135.525 ;
        RECT 74.275 135.065 74.555 135.525 ;
        RECT 75.075 135.235 75.400 135.695 ;
        RECT 74.275 134.845 75.400 135.065 ;
        RECT 73.685 134.115 74.780 134.675 ;
        RECT 74.950 134.385 75.400 134.845 ;
        RECT 75.570 134.555 75.955 135.525 ;
        RECT 72.560 133.315 72.845 133.775 ;
        RECT 73.015 133.145 73.285 133.605 ;
        RECT 73.685 133.315 74.085 134.115 ;
        RECT 74.950 134.055 75.505 134.385 ;
        RECT 74.950 133.945 75.400 134.055 ;
        RECT 74.275 133.775 75.400 133.945 ;
        RECT 75.675 133.885 75.955 134.555 ;
        RECT 76.585 134.530 76.875 135.695 ;
        RECT 77.050 134.745 77.315 135.515 ;
        RECT 77.485 134.975 77.815 135.695 ;
        RECT 78.005 135.155 78.265 135.515 ;
        RECT 78.435 135.325 78.765 135.695 ;
        RECT 78.935 135.155 79.195 135.515 ;
        RECT 78.005 134.925 79.195 135.155 ;
        RECT 79.765 134.745 80.055 135.515 ;
        RECT 81.275 135.025 81.445 135.525 ;
        RECT 81.615 135.195 81.945 135.695 ;
        RECT 81.275 134.855 81.940 135.025 ;
        RECT 74.275 133.315 74.555 133.775 ;
        RECT 75.075 133.145 75.400 133.605 ;
        RECT 75.570 133.315 75.955 133.885 ;
        RECT 76.585 133.145 76.875 133.870 ;
        RECT 77.050 133.325 77.385 134.745 ;
        RECT 77.560 134.565 80.055 134.745 ;
        RECT 77.560 133.875 77.785 134.565 ;
        RECT 77.985 134.055 78.265 134.385 ;
        RECT 78.445 134.055 79.020 134.385 ;
        RECT 79.200 134.055 79.635 134.385 ;
        RECT 79.815 134.055 80.085 134.385 ;
        RECT 81.190 134.035 81.540 134.685 ;
        RECT 77.560 133.685 80.045 133.875 ;
        RECT 81.710 133.865 81.940 134.855 ;
        RECT 77.565 133.145 78.310 133.515 ;
        RECT 78.875 133.325 79.130 133.685 ;
        RECT 79.310 133.145 79.640 133.515 ;
        RECT 79.820 133.325 80.045 133.685 ;
        RECT 81.275 133.695 81.940 133.865 ;
        RECT 81.275 133.405 81.445 133.695 ;
        RECT 81.615 133.145 81.945 133.525 ;
        RECT 82.115 133.405 82.300 135.525 ;
        RECT 82.540 135.235 82.805 135.695 ;
        RECT 82.975 135.100 83.225 135.525 ;
        RECT 83.435 135.250 84.540 135.420 ;
        RECT 82.920 134.970 83.225 135.100 ;
        RECT 82.470 133.775 82.750 134.725 ;
        RECT 82.920 133.865 83.090 134.970 ;
        RECT 83.260 134.185 83.500 134.780 ;
        RECT 83.670 134.715 84.200 135.080 ;
        RECT 83.670 134.015 83.840 134.715 ;
        RECT 84.370 134.635 84.540 135.250 ;
        RECT 84.710 134.895 84.880 135.695 ;
        RECT 85.050 135.195 85.300 135.525 ;
        RECT 85.525 135.225 86.410 135.395 ;
        RECT 84.370 134.545 84.880 134.635 ;
        RECT 82.920 133.735 83.145 133.865 ;
        RECT 83.315 133.795 83.840 134.015 ;
        RECT 84.010 134.375 84.880 134.545 ;
        RECT 82.555 133.145 82.805 133.605 ;
        RECT 82.975 133.595 83.145 133.735 ;
        RECT 84.010 133.595 84.180 134.375 ;
        RECT 84.710 134.305 84.880 134.375 ;
        RECT 84.390 134.125 84.590 134.155 ;
        RECT 85.050 134.125 85.220 135.195 ;
        RECT 85.390 134.305 85.580 135.025 ;
        RECT 84.390 133.825 85.220 134.125 ;
        RECT 85.750 134.095 86.070 135.055 ;
        RECT 82.975 133.425 83.310 133.595 ;
        RECT 83.505 133.425 84.180 133.595 ;
        RECT 84.500 133.145 84.870 133.645 ;
        RECT 85.050 133.595 85.220 133.825 ;
        RECT 85.605 133.765 86.070 134.095 ;
        RECT 86.240 134.385 86.410 135.225 ;
        RECT 86.590 135.195 86.905 135.695 ;
        RECT 87.135 134.965 87.475 135.525 ;
        RECT 86.580 134.590 87.475 134.965 ;
        RECT 87.645 134.685 87.815 135.695 ;
        RECT 87.285 134.385 87.475 134.590 ;
        RECT 87.985 134.635 88.315 135.480 ;
        RECT 87.985 134.555 88.375 134.635 ;
        RECT 88.160 134.505 88.375 134.555 ;
        RECT 86.240 134.055 87.115 134.385 ;
        RECT 87.285 134.055 88.035 134.385 ;
        RECT 86.240 133.595 86.410 134.055 ;
        RECT 87.285 133.885 87.485 134.055 ;
        RECT 88.205 133.925 88.375 134.505 ;
        RECT 88.545 134.605 89.755 135.695 ;
        RECT 100.130 135.430 102.050 136.700 ;
        RECT 103.560 136.690 104.120 136.700 ;
        RECT 103.790 135.600 104.120 136.690 ;
        RECT 104.490 136.220 105.530 136.390 ;
        RECT 104.490 135.780 105.530 135.950 ;
        RECT 105.700 135.920 105.870 136.250 ;
        RECT 103.950 135.380 104.120 135.600 ;
        RECT 106.210 135.380 106.380 136.790 ;
        RECT 103.950 135.210 106.380 135.380 ;
        RECT 107.960 137.300 118.590 137.470 ;
        RECT 120.020 146.580 126.250 146.740 ;
        RECT 120.020 144.320 120.690 146.580 ;
        RECT 121.360 146.010 125.400 146.180 ;
        RECT 121.020 144.950 121.190 145.950 ;
        RECT 125.570 144.950 125.740 145.950 ;
        RECT 121.360 144.720 125.400 144.890 ;
        RECT 126.080 144.320 126.250 146.580 ;
        RECT 120.020 144.150 126.250 144.320 ;
        RECT 120.020 140.890 120.690 144.150 ;
        RECT 121.360 143.580 125.400 143.750 ;
        RECT 121.020 141.520 121.190 143.520 ;
        RECT 125.570 141.520 125.740 143.520 ;
        RECT 121.360 141.290 125.400 141.460 ;
        RECT 126.080 140.890 126.250 144.150 ;
        RECT 120.020 140.720 126.250 140.890 ;
        RECT 120.020 137.460 120.690 140.720 ;
        RECT 121.360 140.150 125.400 140.320 ;
        RECT 121.020 138.090 121.190 140.090 ;
        RECT 125.570 138.090 125.740 140.090 ;
        RECT 121.360 137.860 125.400 138.030 ;
        RECT 126.080 137.460 126.250 140.720 ;
        RECT 120.020 137.450 126.250 137.460 ;
        RECT 127.840 146.720 137.670 146.760 ;
        RECT 140.540 146.740 146.280 146.750 ;
        RECT 127.840 146.590 138.470 146.720 ;
        RECT 127.840 144.330 128.010 146.590 ;
        RECT 128.735 146.020 136.775 146.190 ;
        RECT 128.350 144.960 128.520 145.960 ;
        RECT 136.990 144.960 137.160 145.960 ;
        RECT 128.735 144.730 136.775 144.900 ;
        RECT 137.500 144.330 138.470 146.590 ;
        RECT 127.840 144.160 138.470 144.330 ;
        RECT 127.840 140.900 128.010 144.160 ;
        RECT 128.735 143.590 136.775 143.760 ;
        RECT 128.350 141.530 128.520 143.530 ;
        RECT 136.990 141.530 137.160 143.530 ;
        RECT 128.735 141.300 136.775 141.470 ;
        RECT 137.500 140.900 138.470 144.160 ;
        RECT 127.840 140.730 138.470 140.900 ;
        RECT 127.840 137.470 128.010 140.730 ;
        RECT 128.735 140.160 136.775 140.330 ;
        RECT 128.350 138.100 128.520 140.100 ;
        RECT 136.990 138.100 137.160 140.100 ;
        RECT 128.735 137.870 136.775 138.040 ;
        RECT 137.500 137.470 138.470 140.730 ;
        RECT 120.020 137.350 126.260 137.450 ;
        RECT 107.960 135.040 108.130 137.300 ;
        RECT 108.855 136.730 116.895 136.900 ;
        RECT 108.470 135.670 108.640 136.670 ;
        RECT 117.110 135.670 117.280 136.670 ;
        RECT 108.855 135.440 116.895 135.610 ;
        RECT 117.620 135.040 118.590 137.300 ;
        RECT 120.010 136.790 126.260 137.350 ;
        RECT 120.010 136.770 125.180 136.790 ;
        RECT 120.010 136.700 124.000 136.770 ;
        RECT 120.010 135.430 121.930 136.700 ;
        RECT 123.440 136.690 124.000 136.700 ;
        RECT 123.670 135.600 124.000 136.690 ;
        RECT 124.370 136.220 125.410 136.390 ;
        RECT 124.370 135.780 125.410 135.950 ;
        RECT 125.580 135.920 125.750 136.250 ;
        RECT 123.830 135.380 124.000 135.600 ;
        RECT 126.090 135.380 126.260 136.790 ;
        RECT 123.830 135.210 126.260 135.380 ;
        RECT 127.840 137.300 138.470 137.470 ;
        RECT 140.050 146.580 146.280 146.740 ;
        RECT 140.050 144.320 140.720 146.580 ;
        RECT 141.390 146.010 145.430 146.180 ;
        RECT 141.050 144.950 141.220 145.950 ;
        RECT 145.600 144.950 145.770 145.950 ;
        RECT 141.390 144.720 145.430 144.890 ;
        RECT 146.110 144.320 146.280 146.580 ;
        RECT 140.050 144.150 146.280 144.320 ;
        RECT 140.050 140.890 140.720 144.150 ;
        RECT 141.390 143.580 145.430 143.750 ;
        RECT 141.050 141.520 141.220 143.520 ;
        RECT 145.600 141.520 145.770 143.520 ;
        RECT 141.390 141.290 145.430 141.460 ;
        RECT 146.110 140.890 146.280 144.150 ;
        RECT 140.050 140.720 146.280 140.890 ;
        RECT 140.050 137.460 140.720 140.720 ;
        RECT 141.390 140.150 145.430 140.320 ;
        RECT 141.050 138.090 141.220 140.090 ;
        RECT 145.600 138.090 145.770 140.090 ;
        RECT 141.390 137.860 145.430 138.030 ;
        RECT 146.110 137.460 146.280 140.720 ;
        RECT 140.050 137.450 146.280 137.460 ;
        RECT 147.870 146.720 157.700 146.760 ;
        RECT 147.870 146.590 158.500 146.720 ;
        RECT 147.870 144.330 148.040 146.590 ;
        RECT 148.765 146.020 156.805 146.190 ;
        RECT 148.380 144.960 148.550 145.960 ;
        RECT 157.020 144.960 157.190 145.960 ;
        RECT 148.765 144.730 156.805 144.900 ;
        RECT 157.530 144.330 158.500 146.590 ;
        RECT 147.870 144.160 158.500 144.330 ;
        RECT 147.870 140.900 148.040 144.160 ;
        RECT 148.765 143.590 156.805 143.760 ;
        RECT 148.380 141.530 148.550 143.530 ;
        RECT 157.020 141.530 157.190 143.530 ;
        RECT 148.765 141.300 156.805 141.470 ;
        RECT 157.530 140.900 158.500 144.160 ;
        RECT 147.870 140.730 158.500 140.900 ;
        RECT 147.870 137.470 148.040 140.730 ;
        RECT 148.765 140.160 156.805 140.330 ;
        RECT 148.380 138.100 148.550 140.100 ;
        RECT 157.020 138.100 157.190 140.100 ;
        RECT 148.765 137.870 156.805 138.040 ;
        RECT 157.530 137.470 158.500 140.730 ;
        RECT 140.050 137.350 146.290 137.450 ;
        RECT 107.960 135.010 118.590 135.040 ;
        RECT 127.840 135.040 128.010 137.300 ;
        RECT 128.735 136.730 136.775 136.900 ;
        RECT 128.350 135.670 128.520 136.670 ;
        RECT 136.990 135.670 137.160 136.670 ;
        RECT 128.735 135.440 136.775 135.610 ;
        RECT 137.500 135.040 138.470 137.300 ;
        RECT 140.040 136.790 146.290 137.350 ;
        RECT 140.040 136.770 145.210 136.790 ;
        RECT 140.040 136.700 144.030 136.770 ;
        RECT 140.040 135.430 141.960 136.700 ;
        RECT 143.470 136.690 144.030 136.700 ;
        RECT 143.700 135.600 144.030 136.690 ;
        RECT 144.400 136.220 145.440 136.390 ;
        RECT 144.400 135.780 145.440 135.950 ;
        RECT 145.610 135.920 145.780 136.250 ;
        RECT 143.860 135.380 144.030 135.600 ;
        RECT 146.120 135.380 146.290 136.790 ;
        RECT 143.860 135.210 146.290 135.380 ;
        RECT 147.870 137.300 158.500 137.470 ;
        RECT 127.840 135.010 138.470 135.040 ;
        RECT 147.870 135.040 148.040 137.300 ;
        RECT 148.765 136.730 156.805 136.900 ;
        RECT 148.380 135.670 148.550 136.670 ;
        RECT 157.020 135.670 157.190 136.670 ;
        RECT 148.765 135.440 156.805 135.610 ;
        RECT 157.530 135.040 158.500 137.300 ;
        RECT 147.870 135.010 158.500 135.040 ;
        RECT 107.930 134.900 118.590 135.010 ;
        RECT 127.810 134.900 138.470 135.010 ;
        RECT 147.840 134.900 158.500 135.010 ;
        RECT 106.180 134.850 118.590 134.900 ;
        RECT 126.060 134.850 138.470 134.900 ;
        RECT 146.090 134.850 158.500 134.900 ;
        RECT 101.840 134.680 118.590 134.850 ;
        RECT 88.545 134.065 89.065 134.605 ;
        RECT 88.150 133.885 88.375 133.925 ;
        RECT 89.235 133.895 89.755 134.435 ;
        RECT 85.050 133.425 85.455 133.595 ;
        RECT 85.625 133.425 86.410 133.595 ;
        RECT 86.685 133.145 86.895 133.675 ;
        RECT 87.155 133.360 87.485 133.885 ;
        RECT 87.995 133.800 88.375 133.885 ;
        RECT 87.655 133.145 87.825 133.755 ;
        RECT 87.995 133.365 88.325 133.800 ;
        RECT 88.545 133.145 89.755 133.895 ;
        RECT 101.840 133.270 102.010 134.680 ;
        RECT 102.380 134.110 105.420 134.280 ;
        RECT 102.380 133.670 105.420 133.840 ;
        RECT 105.635 133.810 105.805 134.140 ;
        RECT 106.140 133.920 118.590 134.680 ;
        RECT 121.720 134.680 138.470 134.850 ;
        RECT 106.140 133.910 118.480 133.920 ;
        RECT 106.140 133.900 112.020 133.910 ;
        RECT 106.140 133.880 106.710 133.900 ;
        RECT 107.930 133.890 112.020 133.900 ;
        RECT 106.150 133.270 106.320 133.880 ;
        RECT 12.100 132.975 89.840 133.145 ;
        RECT 101.840 133.100 106.320 133.270 ;
        RECT 121.720 133.270 121.890 134.680 ;
        RECT 122.260 134.110 125.300 134.280 ;
        RECT 122.260 133.670 125.300 133.840 ;
        RECT 125.515 133.810 125.685 134.140 ;
        RECT 126.020 133.920 138.470 134.680 ;
        RECT 141.750 134.680 158.500 134.850 ;
        RECT 126.020 133.910 138.360 133.920 ;
        RECT 126.020 133.900 131.900 133.910 ;
        RECT 126.020 133.880 126.590 133.900 ;
        RECT 127.810 133.890 131.900 133.900 ;
        RECT 126.030 133.270 126.200 133.880 ;
        RECT 121.720 133.100 126.200 133.270 ;
        RECT 141.750 133.270 141.920 134.680 ;
        RECT 142.290 134.110 145.330 134.280 ;
        RECT 142.290 133.670 145.330 133.840 ;
        RECT 145.545 133.810 145.715 134.140 ;
        RECT 146.050 133.920 158.500 134.680 ;
        RECT 146.050 133.910 158.390 133.920 ;
        RECT 146.050 133.900 151.930 133.910 ;
        RECT 146.050 133.880 146.620 133.900 ;
        RECT 147.840 133.890 151.930 133.900 ;
        RECT 146.060 133.270 146.230 133.880 ;
        RECT 141.750 133.100 146.230 133.270 ;
        RECT 12.185 132.225 13.395 132.975 ;
        RECT 13.565 132.225 14.775 132.975 ;
        RECT 14.950 132.720 15.285 132.765 ;
        RECT 14.945 132.255 15.285 132.720 ;
        RECT 15.455 132.595 15.785 132.975 ;
        RECT 12.185 131.685 12.705 132.225 ;
        RECT 12.875 131.515 13.395 132.055 ;
        RECT 13.565 131.685 14.085 132.225 ;
        RECT 14.255 131.515 14.775 132.055 ;
        RECT 12.185 130.425 13.395 131.515 ;
        RECT 13.565 130.425 14.775 131.515 ;
        RECT 14.945 131.565 15.115 132.255 ;
        RECT 15.285 131.735 15.545 132.065 ;
        RECT 14.945 130.595 15.205 131.565 ;
        RECT 15.375 131.185 15.545 131.735 ;
        RECT 15.715 131.365 16.055 132.395 ;
        RECT 16.245 131.955 16.515 132.640 ;
        RECT 16.245 131.785 16.555 131.955 ;
        RECT 16.245 131.365 16.515 131.785 ;
        RECT 16.740 131.365 17.020 132.640 ;
        RECT 17.220 132.475 17.450 132.805 ;
        RECT 17.695 132.595 18.025 132.975 ;
        RECT 17.220 131.185 17.390 132.475 ;
        RECT 18.195 132.405 18.370 132.805 ;
        RECT 18.625 132.430 23.970 132.975 ;
        RECT 17.740 132.235 18.370 132.405 ;
        RECT 17.740 132.065 17.910 132.235 ;
        RECT 17.560 131.735 17.910 132.065 ;
        RECT 15.375 131.015 17.390 131.185 ;
        RECT 17.740 131.215 17.910 131.735 ;
        RECT 18.090 131.385 18.455 132.065 ;
        RECT 20.210 131.600 20.550 132.430 ;
        RECT 24.235 132.425 24.405 132.805 ;
        RECT 24.620 132.595 24.950 132.975 ;
        RECT 24.235 132.255 24.950 132.425 ;
        RECT 17.740 131.045 18.370 131.215 ;
        RECT 15.400 130.425 15.730 130.835 ;
        RECT 15.930 130.595 16.100 131.015 ;
        RECT 16.315 130.425 16.985 130.835 ;
        RECT 17.220 130.595 17.390 131.015 ;
        RECT 17.695 130.425 18.025 130.865 ;
        RECT 18.195 130.595 18.370 131.045 ;
        RECT 22.030 130.860 22.380 132.110 ;
        RECT 24.145 131.705 24.500 132.075 ;
        RECT 24.780 132.065 24.950 132.255 ;
        RECT 25.120 132.230 25.375 132.805 ;
        RECT 24.780 131.735 25.035 132.065 ;
        RECT 24.780 131.525 24.950 131.735 ;
        RECT 24.235 131.355 24.950 131.525 ;
        RECT 25.205 131.500 25.375 132.230 ;
        RECT 25.550 132.135 25.810 132.975 ;
        RECT 25.985 132.345 26.325 132.805 ;
        RECT 26.495 132.515 26.665 132.975 ;
        RECT 27.295 132.540 27.655 132.805 ;
        RECT 27.300 132.535 27.655 132.540 ;
        RECT 27.305 132.525 27.655 132.535 ;
        RECT 27.310 132.520 27.655 132.525 ;
        RECT 27.315 132.510 27.655 132.520 ;
        RECT 27.895 132.515 28.065 132.975 ;
        RECT 27.320 132.505 27.655 132.510 ;
        RECT 27.330 132.495 27.655 132.505 ;
        RECT 27.340 132.485 27.655 132.495 ;
        RECT 26.835 132.345 27.165 132.425 ;
        RECT 25.985 132.155 27.165 132.345 ;
        RECT 27.355 132.345 27.655 132.485 ;
        RECT 27.355 132.155 28.065 132.345 ;
        RECT 25.985 131.785 26.315 131.985 ;
        RECT 26.625 131.965 26.955 131.985 ;
        RECT 26.505 131.785 26.955 131.965 ;
        RECT 18.625 130.425 23.970 130.860 ;
        RECT 24.235 130.595 24.405 131.355 ;
        RECT 24.620 130.425 24.950 131.185 ;
        RECT 25.120 130.595 25.375 131.500 ;
        RECT 25.550 130.425 25.810 131.575 ;
        RECT 25.985 131.445 26.215 131.785 ;
        RECT 25.995 130.425 26.325 131.145 ;
        RECT 26.505 130.670 26.720 131.785 ;
        RECT 27.125 131.755 27.595 131.985 ;
        RECT 27.780 131.585 28.065 132.155 ;
        RECT 28.235 132.030 28.575 132.805 ;
        RECT 26.915 131.370 28.065 131.585 ;
        RECT 26.915 130.595 27.245 131.370 ;
        RECT 27.415 130.425 28.125 131.200 ;
        RECT 28.295 130.595 28.575 132.030 ;
        RECT 28.745 132.515 29.305 132.805 ;
        RECT 29.475 132.515 29.725 132.975 ;
        RECT 28.745 131.145 28.995 132.515 ;
        RECT 30.345 132.345 30.675 132.705 ;
        RECT 29.285 132.155 30.675 132.345 ;
        RECT 31.045 132.205 32.715 132.975 ;
        RECT 29.285 132.065 29.455 132.155 ;
        RECT 29.165 131.735 29.455 132.065 ;
        RECT 29.625 131.735 29.965 131.985 ;
        RECT 30.185 131.735 30.860 131.985 ;
        RECT 29.285 131.485 29.455 131.735 ;
        RECT 29.285 131.315 30.225 131.485 ;
        RECT 30.595 131.375 30.860 131.735 ;
        RECT 31.045 131.685 31.795 132.205 ;
        RECT 32.895 132.165 33.165 132.975 ;
        RECT 33.335 132.165 33.665 132.805 ;
        RECT 33.835 132.165 34.075 132.975 ;
        RECT 34.745 132.505 35.040 132.975 ;
        RECT 35.210 132.335 35.470 132.780 ;
        RECT 35.640 132.505 35.900 132.975 ;
        RECT 36.070 132.335 36.325 132.780 ;
        RECT 36.495 132.505 36.795 132.975 ;
        RECT 34.285 132.165 37.315 132.335 ;
        RECT 37.945 132.250 38.235 132.975 ;
        RECT 38.425 132.165 38.665 132.975 ;
        RECT 38.835 132.165 39.165 132.805 ;
        RECT 39.335 132.165 39.605 132.975 ;
        RECT 40.795 132.425 40.965 132.715 ;
        RECT 41.135 132.595 41.465 132.975 ;
        RECT 40.795 132.255 41.460 132.425 ;
        RECT 31.965 131.515 32.715 132.035 ;
        RECT 32.885 131.735 33.235 131.985 ;
        RECT 33.405 131.565 33.575 132.165 ;
        RECT 33.745 131.735 34.095 131.985 ;
        RECT 34.285 131.600 34.455 132.165 ;
        RECT 34.625 131.770 36.840 131.995 ;
        RECT 37.015 131.600 37.315 132.165 ;
        RECT 38.405 131.735 38.755 131.985 ;
        RECT 28.745 130.595 29.205 131.145 ;
        RECT 29.395 130.425 29.725 131.145 ;
        RECT 29.925 130.765 30.225 131.315 ;
        RECT 30.395 130.425 30.675 131.095 ;
        RECT 31.045 130.425 32.715 131.515 ;
        RECT 32.895 130.425 33.225 131.565 ;
        RECT 33.405 131.395 34.085 131.565 ;
        RECT 34.285 131.430 37.315 131.600 ;
        RECT 33.755 130.610 34.085 131.395 ;
        RECT 34.265 130.425 34.610 131.260 ;
        RECT 34.785 130.625 35.040 131.430 ;
        RECT 35.210 130.425 35.470 131.260 ;
        RECT 35.645 130.625 35.900 131.430 ;
        RECT 36.070 130.425 36.330 131.260 ;
        RECT 36.500 130.625 36.760 131.430 ;
        RECT 36.930 130.425 37.315 131.260 ;
        RECT 37.945 130.425 38.235 131.590 ;
        RECT 38.925 131.565 39.095 132.165 ;
        RECT 39.265 131.735 39.615 131.985 ;
        RECT 38.415 131.395 39.095 131.565 ;
        RECT 38.415 130.610 38.745 131.395 ;
        RECT 39.275 130.425 39.605 131.565 ;
        RECT 40.710 131.435 41.060 132.085 ;
        RECT 41.230 131.265 41.460 132.255 ;
        RECT 40.795 131.095 41.460 131.265 ;
        RECT 40.795 130.595 40.965 131.095 ;
        RECT 41.135 130.425 41.465 130.925 ;
        RECT 41.635 130.595 41.820 132.715 ;
        RECT 42.075 132.515 42.325 132.975 ;
        RECT 42.495 132.525 42.830 132.695 ;
        RECT 43.025 132.525 43.700 132.695 ;
        RECT 42.495 132.385 42.665 132.525 ;
        RECT 41.990 131.395 42.270 132.345 ;
        RECT 42.440 132.255 42.665 132.385 ;
        RECT 42.440 131.150 42.610 132.255 ;
        RECT 42.835 132.105 43.360 132.325 ;
        RECT 42.780 131.340 43.020 131.935 ;
        RECT 43.190 131.405 43.360 132.105 ;
        RECT 43.530 131.745 43.700 132.525 ;
        RECT 44.020 132.475 44.390 132.975 ;
        RECT 44.570 132.525 44.975 132.695 ;
        RECT 45.145 132.525 45.930 132.695 ;
        RECT 44.570 132.295 44.740 132.525 ;
        RECT 43.910 131.995 44.740 132.295 ;
        RECT 45.125 132.025 45.590 132.355 ;
        RECT 43.910 131.965 44.110 131.995 ;
        RECT 44.230 131.745 44.400 131.815 ;
        RECT 43.530 131.575 44.400 131.745 ;
        RECT 43.890 131.485 44.400 131.575 ;
        RECT 42.440 131.020 42.745 131.150 ;
        RECT 43.190 131.040 43.720 131.405 ;
        RECT 42.060 130.425 42.325 130.885 ;
        RECT 42.495 130.595 42.745 131.020 ;
        RECT 43.890 130.870 44.060 131.485 ;
        RECT 42.955 130.700 44.060 130.870 ;
        RECT 44.230 130.425 44.400 131.225 ;
        RECT 44.570 130.925 44.740 131.995 ;
        RECT 44.910 131.095 45.100 131.815 ;
        RECT 45.270 131.065 45.590 132.025 ;
        RECT 45.760 132.065 45.930 132.525 ;
        RECT 46.205 132.445 46.415 132.975 ;
        RECT 46.675 132.235 47.005 132.760 ;
        RECT 47.175 132.365 47.345 132.975 ;
        RECT 47.515 132.320 47.845 132.755 ;
        RECT 47.515 132.235 47.895 132.320 ;
        RECT 46.805 132.065 47.005 132.235 ;
        RECT 47.670 132.195 47.895 132.235 ;
        RECT 45.760 131.735 46.635 132.065 ;
        RECT 46.805 131.735 47.555 132.065 ;
        RECT 44.570 130.595 44.820 130.925 ;
        RECT 45.760 130.895 45.930 131.735 ;
        RECT 46.805 131.530 46.995 131.735 ;
        RECT 47.725 131.615 47.895 132.195 ;
        RECT 47.680 131.565 47.895 131.615 ;
        RECT 46.100 131.155 46.995 131.530 ;
        RECT 47.505 131.485 47.895 131.565 ;
        RECT 48.070 132.235 48.325 132.805 ;
        RECT 48.495 132.575 48.825 132.975 ;
        RECT 49.250 132.440 49.780 132.805 ;
        RECT 49.250 132.405 49.425 132.440 ;
        RECT 48.495 132.235 49.425 132.405 ;
        RECT 49.970 132.295 50.245 132.805 ;
        RECT 48.070 131.565 48.240 132.235 ;
        RECT 48.495 132.065 48.665 132.235 ;
        RECT 48.410 131.735 48.665 132.065 ;
        RECT 48.890 131.735 49.085 132.065 ;
        RECT 45.045 130.725 45.930 130.895 ;
        RECT 46.110 130.425 46.425 130.925 ;
        RECT 46.655 130.595 46.995 131.155 ;
        RECT 47.165 130.425 47.335 131.435 ;
        RECT 47.505 130.640 47.835 131.485 ;
        RECT 48.070 130.595 48.405 131.565 ;
        RECT 48.575 130.425 48.745 131.565 ;
        RECT 48.915 130.765 49.085 131.735 ;
        RECT 49.255 131.105 49.425 132.235 ;
        RECT 49.595 131.445 49.765 132.245 ;
        RECT 49.965 132.125 50.245 132.295 ;
        RECT 49.970 131.645 50.245 132.125 ;
        RECT 50.415 131.445 50.605 132.805 ;
        RECT 50.785 132.440 51.295 132.975 ;
        RECT 51.515 132.165 51.760 132.770 ;
        RECT 52.205 132.475 52.505 132.805 ;
        RECT 52.675 132.495 52.950 132.975 ;
        RECT 50.805 131.995 52.035 132.165 ;
        RECT 49.595 131.275 50.605 131.445 ;
        RECT 50.775 131.430 51.525 131.620 ;
        RECT 49.255 130.935 50.380 131.105 ;
        RECT 50.775 130.765 50.945 131.430 ;
        RECT 51.695 131.185 52.035 131.995 ;
        RECT 48.915 130.595 50.945 130.765 ;
        RECT 51.115 130.425 51.285 131.185 ;
        RECT 51.520 130.775 52.035 131.185 ;
        RECT 52.205 131.565 52.375 132.475 ;
        RECT 53.130 132.325 53.425 132.715 ;
        RECT 53.595 132.495 53.850 132.975 ;
        RECT 54.025 132.325 54.285 132.715 ;
        RECT 54.455 132.495 54.735 132.975 ;
        RECT 52.545 131.735 52.895 132.305 ;
        RECT 53.130 132.155 54.780 132.325 ;
        RECT 53.065 131.815 54.205 131.985 ;
        RECT 53.065 131.565 53.235 131.815 ;
        RECT 54.375 131.645 54.780 132.155 ;
        RECT 54.965 132.225 56.175 132.975 ;
        RECT 56.435 132.425 56.605 132.715 ;
        RECT 56.775 132.595 57.105 132.975 ;
        RECT 56.435 132.255 57.100 132.425 ;
        RECT 54.965 131.685 55.485 132.225 ;
        RECT 52.205 131.395 53.235 131.565 ;
        RECT 54.025 131.475 54.780 131.645 ;
        RECT 55.655 131.515 56.175 132.055 ;
        RECT 52.205 130.595 52.515 131.395 ;
        RECT 54.025 131.225 54.285 131.475 ;
        RECT 52.685 130.425 52.995 131.225 ;
        RECT 53.165 131.055 54.285 131.225 ;
        RECT 53.165 130.595 53.425 131.055 ;
        RECT 53.595 130.425 53.850 130.885 ;
        RECT 54.025 130.595 54.285 131.055 ;
        RECT 54.455 130.425 54.740 131.295 ;
        RECT 54.965 130.425 56.175 131.515 ;
        RECT 56.350 131.435 56.700 132.085 ;
        RECT 56.870 131.265 57.100 132.255 ;
        RECT 56.435 131.095 57.100 131.265 ;
        RECT 56.435 130.595 56.605 131.095 ;
        RECT 56.775 130.425 57.105 130.925 ;
        RECT 57.275 130.595 57.460 132.715 ;
        RECT 57.715 132.515 57.965 132.975 ;
        RECT 58.135 132.525 58.470 132.695 ;
        RECT 58.665 132.525 59.340 132.695 ;
        RECT 58.135 132.385 58.305 132.525 ;
        RECT 57.630 131.395 57.910 132.345 ;
        RECT 58.080 132.255 58.305 132.385 ;
        RECT 58.080 131.150 58.250 132.255 ;
        RECT 58.475 132.105 59.000 132.325 ;
        RECT 58.420 131.340 58.660 131.935 ;
        RECT 58.830 131.405 59.000 132.105 ;
        RECT 59.170 131.745 59.340 132.525 ;
        RECT 59.660 132.475 60.030 132.975 ;
        RECT 60.210 132.525 60.615 132.695 ;
        RECT 60.785 132.525 61.570 132.695 ;
        RECT 60.210 132.295 60.380 132.525 ;
        RECT 59.550 131.995 60.380 132.295 ;
        RECT 60.765 132.025 61.230 132.355 ;
        RECT 59.550 131.965 59.750 131.995 ;
        RECT 59.870 131.745 60.040 131.815 ;
        RECT 59.170 131.575 60.040 131.745 ;
        RECT 59.530 131.485 60.040 131.575 ;
        RECT 58.080 131.020 58.385 131.150 ;
        RECT 58.830 131.040 59.360 131.405 ;
        RECT 57.700 130.425 57.965 130.885 ;
        RECT 58.135 130.595 58.385 131.020 ;
        RECT 59.530 130.870 59.700 131.485 ;
        RECT 58.595 130.700 59.700 130.870 ;
        RECT 59.870 130.425 60.040 131.225 ;
        RECT 60.210 130.925 60.380 131.995 ;
        RECT 60.550 131.095 60.740 131.815 ;
        RECT 60.910 131.065 61.230 132.025 ;
        RECT 61.400 132.065 61.570 132.525 ;
        RECT 61.845 132.445 62.055 132.975 ;
        RECT 62.315 132.235 62.645 132.760 ;
        RECT 62.815 132.365 62.985 132.975 ;
        RECT 63.155 132.320 63.485 132.755 ;
        RECT 63.155 132.235 63.535 132.320 ;
        RECT 63.705 132.250 63.995 132.975 ;
        RECT 64.255 132.425 64.425 132.715 ;
        RECT 64.595 132.595 64.925 132.975 ;
        RECT 64.255 132.255 64.920 132.425 ;
        RECT 62.445 132.065 62.645 132.235 ;
        RECT 63.310 132.195 63.535 132.235 ;
        RECT 61.400 131.735 62.275 132.065 ;
        RECT 62.445 131.735 63.195 132.065 ;
        RECT 60.210 130.595 60.460 130.925 ;
        RECT 61.400 130.895 61.570 131.735 ;
        RECT 62.445 131.530 62.635 131.735 ;
        RECT 63.365 131.615 63.535 132.195 ;
        RECT 63.320 131.565 63.535 131.615 ;
        RECT 61.740 131.155 62.635 131.530 ;
        RECT 63.145 131.485 63.535 131.565 ;
        RECT 60.685 130.725 61.570 130.895 ;
        RECT 61.750 130.425 62.065 130.925 ;
        RECT 62.295 130.595 62.635 131.155 ;
        RECT 62.805 130.425 62.975 131.435 ;
        RECT 63.145 130.640 63.475 131.485 ;
        RECT 63.705 130.425 63.995 131.590 ;
        RECT 64.170 131.435 64.520 132.085 ;
        RECT 64.690 131.265 64.920 132.255 ;
        RECT 64.255 131.095 64.920 131.265 ;
        RECT 64.255 130.595 64.425 131.095 ;
        RECT 64.595 130.425 64.925 130.925 ;
        RECT 65.095 130.595 65.280 132.715 ;
        RECT 65.535 132.515 65.785 132.975 ;
        RECT 65.955 132.525 66.290 132.695 ;
        RECT 66.485 132.525 67.160 132.695 ;
        RECT 65.955 132.385 66.125 132.525 ;
        RECT 65.450 131.395 65.730 132.345 ;
        RECT 65.900 132.255 66.125 132.385 ;
        RECT 65.900 131.150 66.070 132.255 ;
        RECT 66.295 132.105 66.820 132.325 ;
        RECT 66.240 131.340 66.480 131.935 ;
        RECT 66.650 131.405 66.820 132.105 ;
        RECT 66.990 131.745 67.160 132.525 ;
        RECT 67.480 132.475 67.850 132.975 ;
        RECT 68.030 132.525 68.435 132.695 ;
        RECT 68.605 132.525 69.390 132.695 ;
        RECT 68.030 132.295 68.200 132.525 ;
        RECT 67.370 131.995 68.200 132.295 ;
        RECT 68.585 132.025 69.050 132.355 ;
        RECT 67.370 131.965 67.570 131.995 ;
        RECT 67.690 131.745 67.860 131.815 ;
        RECT 66.990 131.575 67.860 131.745 ;
        RECT 67.350 131.485 67.860 131.575 ;
        RECT 65.900 131.020 66.205 131.150 ;
        RECT 66.650 131.040 67.180 131.405 ;
        RECT 65.520 130.425 65.785 130.885 ;
        RECT 65.955 130.595 66.205 131.020 ;
        RECT 67.350 130.870 67.520 131.485 ;
        RECT 66.415 130.700 67.520 130.870 ;
        RECT 67.690 130.425 67.860 131.225 ;
        RECT 68.030 130.925 68.200 131.995 ;
        RECT 68.370 131.095 68.560 131.815 ;
        RECT 68.730 131.065 69.050 132.025 ;
        RECT 69.220 132.065 69.390 132.525 ;
        RECT 69.665 132.445 69.875 132.975 ;
        RECT 70.135 132.235 70.465 132.760 ;
        RECT 70.635 132.365 70.805 132.975 ;
        RECT 70.975 132.320 71.305 132.755 ;
        RECT 70.975 132.235 71.355 132.320 ;
        RECT 70.265 132.065 70.465 132.235 ;
        RECT 71.130 132.195 71.355 132.235 ;
        RECT 69.220 131.735 70.095 132.065 ;
        RECT 70.265 131.735 71.015 132.065 ;
        RECT 68.030 130.595 68.280 130.925 ;
        RECT 69.220 130.895 69.390 131.735 ;
        RECT 70.265 131.530 70.455 131.735 ;
        RECT 71.185 131.615 71.355 132.195 ;
        RECT 71.140 131.565 71.355 131.615 ;
        RECT 69.560 131.155 70.455 131.530 ;
        RECT 70.965 131.485 71.355 131.565 ;
        RECT 71.530 132.235 71.785 132.805 ;
        RECT 71.955 132.575 72.285 132.975 ;
        RECT 72.710 132.440 73.240 132.805 ;
        RECT 73.430 132.635 73.705 132.805 ;
        RECT 73.425 132.465 73.705 132.635 ;
        RECT 72.710 132.405 72.885 132.440 ;
        RECT 71.955 132.235 72.885 132.405 ;
        RECT 71.530 131.565 71.700 132.235 ;
        RECT 71.955 132.065 72.125 132.235 ;
        RECT 71.870 131.735 72.125 132.065 ;
        RECT 72.350 131.735 72.545 132.065 ;
        RECT 68.505 130.725 69.390 130.895 ;
        RECT 69.570 130.425 69.885 130.925 ;
        RECT 70.115 130.595 70.455 131.155 ;
        RECT 70.625 130.425 70.795 131.435 ;
        RECT 70.965 130.640 71.295 131.485 ;
        RECT 71.530 130.595 71.865 131.565 ;
        RECT 72.035 130.425 72.205 131.565 ;
        RECT 72.375 130.765 72.545 131.735 ;
        RECT 72.715 131.105 72.885 132.235 ;
        RECT 73.055 131.445 73.225 132.245 ;
        RECT 73.430 131.645 73.705 132.465 ;
        RECT 73.875 131.445 74.065 132.805 ;
        RECT 74.245 132.440 74.755 132.975 ;
        RECT 74.975 132.165 75.220 132.770 ;
        RECT 74.265 131.995 75.495 132.165 ;
        RECT 75.670 132.135 75.930 132.975 ;
        RECT 76.105 132.230 76.360 132.805 ;
        RECT 76.530 132.595 76.860 132.975 ;
        RECT 77.075 132.425 77.245 132.805 ;
        RECT 76.530 132.255 77.245 132.425 ;
        RECT 73.055 131.275 74.065 131.445 ;
        RECT 74.235 131.430 74.985 131.620 ;
        RECT 72.715 130.935 73.840 131.105 ;
        RECT 74.235 130.765 74.405 131.430 ;
        RECT 75.155 131.185 75.495 131.995 ;
        RECT 72.375 130.595 74.405 130.765 ;
        RECT 74.575 130.425 74.745 131.185 ;
        RECT 74.980 130.775 75.495 131.185 ;
        RECT 75.670 130.425 75.930 131.575 ;
        RECT 76.105 131.500 76.275 132.230 ;
        RECT 76.530 132.065 76.700 132.255 ;
        RECT 77.710 132.195 78.210 132.805 ;
        RECT 76.445 131.735 76.700 132.065 ;
        RECT 76.530 131.525 76.700 131.735 ;
        RECT 76.980 131.705 77.335 132.075 ;
        RECT 77.505 131.735 77.855 131.985 ;
        RECT 78.040 131.565 78.210 132.195 ;
        RECT 78.840 132.325 79.170 132.805 ;
        RECT 79.340 132.515 79.565 132.975 ;
        RECT 79.735 132.325 80.065 132.805 ;
        RECT 78.840 132.155 80.065 132.325 ;
        RECT 80.255 132.175 80.505 132.975 ;
        RECT 80.675 132.175 81.015 132.805 ;
        RECT 81.275 132.425 81.445 132.715 ;
        RECT 81.615 132.595 81.945 132.975 ;
        RECT 81.275 132.255 81.940 132.425 ;
        RECT 78.380 131.785 78.710 131.985 ;
        RECT 78.880 131.785 79.210 131.985 ;
        RECT 79.380 131.785 79.800 131.985 ;
        RECT 79.975 131.815 80.670 131.985 ;
        RECT 79.975 131.565 80.145 131.815 ;
        RECT 80.840 131.565 81.015 132.175 ;
        RECT 76.105 130.595 76.360 131.500 ;
        RECT 76.530 131.355 77.245 131.525 ;
        RECT 76.530 130.425 76.860 131.185 ;
        RECT 77.075 130.595 77.245 131.355 ;
        RECT 77.710 131.395 80.145 131.565 ;
        RECT 77.710 130.595 78.040 131.395 ;
        RECT 78.210 130.425 78.540 131.225 ;
        RECT 78.840 130.595 79.170 131.395 ;
        RECT 79.815 130.425 80.065 131.225 ;
        RECT 80.335 130.425 80.505 131.565 ;
        RECT 80.675 130.595 81.015 131.565 ;
        RECT 81.190 131.435 81.540 132.085 ;
        RECT 81.710 131.265 81.940 132.255 ;
        RECT 81.275 131.095 81.940 131.265 ;
        RECT 81.275 130.595 81.445 131.095 ;
        RECT 81.615 130.425 81.945 130.925 ;
        RECT 82.115 130.595 82.300 132.715 ;
        RECT 82.555 132.515 82.805 132.975 ;
        RECT 82.975 132.525 83.310 132.695 ;
        RECT 83.505 132.525 84.180 132.695 ;
        RECT 82.975 132.385 83.145 132.525 ;
        RECT 82.470 131.395 82.750 132.345 ;
        RECT 82.920 132.255 83.145 132.385 ;
        RECT 82.920 131.150 83.090 132.255 ;
        RECT 83.315 132.105 83.840 132.325 ;
        RECT 83.260 131.340 83.500 131.935 ;
        RECT 83.670 131.405 83.840 132.105 ;
        RECT 84.010 131.745 84.180 132.525 ;
        RECT 84.500 132.475 84.870 132.975 ;
        RECT 85.050 132.525 85.455 132.695 ;
        RECT 85.625 132.525 86.410 132.695 ;
        RECT 85.050 132.295 85.220 132.525 ;
        RECT 84.390 131.995 85.220 132.295 ;
        RECT 85.605 132.025 86.070 132.355 ;
        RECT 84.390 131.965 84.590 131.995 ;
        RECT 84.710 131.745 84.880 131.815 ;
        RECT 84.010 131.575 84.880 131.745 ;
        RECT 84.370 131.485 84.880 131.575 ;
        RECT 82.920 131.020 83.225 131.150 ;
        RECT 83.670 131.040 84.200 131.405 ;
        RECT 82.540 130.425 82.805 130.885 ;
        RECT 82.975 130.595 83.225 131.020 ;
        RECT 84.370 130.870 84.540 131.485 ;
        RECT 83.435 130.700 84.540 130.870 ;
        RECT 84.710 130.425 84.880 131.225 ;
        RECT 85.050 130.925 85.220 131.995 ;
        RECT 85.390 131.095 85.580 131.815 ;
        RECT 85.750 131.065 86.070 132.025 ;
        RECT 86.240 132.065 86.410 132.525 ;
        RECT 86.685 132.445 86.895 132.975 ;
        RECT 87.155 132.235 87.485 132.760 ;
        RECT 87.655 132.365 87.825 132.975 ;
        RECT 87.995 132.320 88.325 132.755 ;
        RECT 87.995 132.235 88.375 132.320 ;
        RECT 87.285 132.065 87.485 132.235 ;
        RECT 88.150 132.195 88.375 132.235 ;
        RECT 88.545 132.225 89.755 132.975 ;
        RECT 86.240 131.735 87.115 132.065 ;
        RECT 87.285 131.735 88.035 132.065 ;
        RECT 85.050 130.595 85.300 130.925 ;
        RECT 86.240 130.895 86.410 131.735 ;
        RECT 87.285 131.530 87.475 131.735 ;
        RECT 88.205 131.615 88.375 132.195 ;
        RECT 88.160 131.565 88.375 131.615 ;
        RECT 86.580 131.155 87.475 131.530 ;
        RECT 87.985 131.485 88.375 131.565 ;
        RECT 88.545 131.515 89.065 132.055 ;
        RECT 89.235 131.685 89.755 132.225 ;
        RECT 120.510 131.800 126.250 131.810 ;
        RECT 100.630 131.740 106.370 131.750 ;
        RECT 100.140 131.580 106.370 131.740 ;
        RECT 85.525 130.725 86.410 130.895 ;
        RECT 86.590 130.425 86.905 130.925 ;
        RECT 87.135 130.595 87.475 131.155 ;
        RECT 87.645 130.425 87.815 131.435 ;
        RECT 87.985 130.640 88.315 131.485 ;
        RECT 88.545 130.425 89.755 131.515 ;
        RECT 12.100 130.255 89.840 130.425 ;
        RECT 12.185 129.165 13.395 130.255 ;
        RECT 14.115 129.585 14.285 130.085 ;
        RECT 14.455 129.755 14.785 130.255 ;
        RECT 14.115 129.415 14.780 129.585 ;
        RECT 12.185 128.455 12.705 128.995 ;
        RECT 12.875 128.625 13.395 129.165 ;
        RECT 14.030 128.595 14.380 129.245 ;
        RECT 12.185 127.705 13.395 128.455 ;
        RECT 14.550 128.425 14.780 129.415 ;
        RECT 14.115 128.255 14.780 128.425 ;
        RECT 14.115 127.965 14.285 128.255 ;
        RECT 14.455 127.705 14.785 128.085 ;
        RECT 14.955 127.965 15.140 130.085 ;
        RECT 15.380 129.795 15.645 130.255 ;
        RECT 15.815 129.660 16.065 130.085 ;
        RECT 16.275 129.810 17.380 129.980 ;
        RECT 15.760 129.530 16.065 129.660 ;
        RECT 15.310 128.335 15.590 129.285 ;
        RECT 15.760 128.425 15.930 129.530 ;
        RECT 16.100 128.745 16.340 129.340 ;
        RECT 16.510 129.275 17.040 129.640 ;
        RECT 16.510 128.575 16.680 129.275 ;
        RECT 17.210 129.195 17.380 129.810 ;
        RECT 17.550 129.455 17.720 130.255 ;
        RECT 17.890 129.755 18.140 130.085 ;
        RECT 18.365 129.785 19.250 129.955 ;
        RECT 17.210 129.105 17.720 129.195 ;
        RECT 15.760 128.295 15.985 128.425 ;
        RECT 16.155 128.355 16.680 128.575 ;
        RECT 16.850 128.935 17.720 129.105 ;
        RECT 15.395 127.705 15.645 128.165 ;
        RECT 15.815 128.155 15.985 128.295 ;
        RECT 16.850 128.155 17.020 128.935 ;
        RECT 17.550 128.865 17.720 128.935 ;
        RECT 17.230 128.685 17.430 128.715 ;
        RECT 17.890 128.685 18.060 129.755 ;
        RECT 18.230 128.865 18.420 129.585 ;
        RECT 17.230 128.385 18.060 128.685 ;
        RECT 18.590 128.655 18.910 129.615 ;
        RECT 15.815 127.985 16.150 128.155 ;
        RECT 16.345 127.985 17.020 128.155 ;
        RECT 17.340 127.705 17.710 128.205 ;
        RECT 17.890 128.155 18.060 128.385 ;
        RECT 18.445 128.325 18.910 128.655 ;
        RECT 19.080 128.945 19.250 129.785 ;
        RECT 19.430 129.755 19.745 130.255 ;
        RECT 19.975 129.525 20.315 130.085 ;
        RECT 19.420 129.150 20.315 129.525 ;
        RECT 20.485 129.245 20.655 130.255 ;
        RECT 20.125 128.945 20.315 129.150 ;
        RECT 20.825 129.195 21.155 130.040 ;
        RECT 21.395 129.285 21.725 130.070 ;
        RECT 20.825 129.115 21.215 129.195 ;
        RECT 21.395 129.115 22.075 129.285 ;
        RECT 22.255 129.115 22.585 130.255 ;
        RECT 23.265 129.795 23.480 130.255 ;
        RECT 23.650 129.625 23.980 130.085 ;
        RECT 22.810 129.455 23.980 129.625 ;
        RECT 24.150 129.455 24.400 130.255 ;
        RECT 21.000 129.065 21.215 129.115 ;
        RECT 19.080 128.615 19.955 128.945 ;
        RECT 20.125 128.615 20.875 128.945 ;
        RECT 19.080 128.155 19.250 128.615 ;
        RECT 20.125 128.445 20.325 128.615 ;
        RECT 21.045 128.485 21.215 129.065 ;
        RECT 21.385 128.695 21.735 128.945 ;
        RECT 21.905 128.515 22.075 129.115 ;
        RECT 22.245 128.695 22.595 128.945 ;
        RECT 20.990 128.445 21.215 128.485 ;
        RECT 17.890 127.985 18.295 128.155 ;
        RECT 18.465 127.985 19.250 128.155 ;
        RECT 19.525 127.705 19.735 128.235 ;
        RECT 19.995 127.920 20.325 128.445 ;
        RECT 20.835 128.360 21.215 128.445 ;
        RECT 20.495 127.705 20.665 128.315 ;
        RECT 20.835 127.925 21.165 128.360 ;
        RECT 21.405 127.705 21.645 128.515 ;
        RECT 21.815 127.875 22.145 128.515 ;
        RECT 22.315 127.705 22.585 128.515 ;
        RECT 22.810 128.165 23.180 129.455 ;
        RECT 24.610 129.285 24.890 129.445 ;
        RECT 23.555 129.115 24.890 129.285 ;
        RECT 23.555 128.945 23.725 129.115 ;
        RECT 25.065 129.090 25.355 130.255 ;
        RECT 25.525 129.115 25.805 130.255 ;
        RECT 25.975 129.105 26.305 130.085 ;
        RECT 26.475 129.115 26.735 130.255 ;
        RECT 26.905 129.285 27.215 130.085 ;
        RECT 27.385 129.455 27.695 130.255 ;
        RECT 27.865 129.625 28.125 130.085 ;
        RECT 28.295 129.795 28.550 130.255 ;
        RECT 28.725 129.625 28.985 130.085 ;
        RECT 27.865 129.455 28.985 129.625 ;
        RECT 26.905 129.115 27.935 129.285 ;
        RECT 23.350 128.695 23.725 128.945 ;
        RECT 23.895 128.695 24.370 128.935 ;
        RECT 24.540 128.695 24.890 128.935 ;
        RECT 23.555 128.525 23.725 128.695 ;
        RECT 25.535 128.675 25.870 128.945 ;
        RECT 23.555 128.355 24.890 128.525 ;
        RECT 26.040 128.505 26.210 129.105 ;
        RECT 26.380 128.695 26.715 128.945 ;
        RECT 22.810 127.875 23.560 128.165 ;
        RECT 24.070 127.705 24.400 128.165 ;
        RECT 24.620 128.145 24.890 128.355 ;
        RECT 25.065 127.705 25.355 128.430 ;
        RECT 25.525 127.705 25.835 128.505 ;
        RECT 26.040 127.875 26.735 128.505 ;
        RECT 26.905 128.205 27.075 129.115 ;
        RECT 27.245 128.375 27.595 128.945 ;
        RECT 27.765 128.865 27.935 129.115 ;
        RECT 28.725 129.205 28.985 129.455 ;
        RECT 29.155 129.385 29.440 130.255 ;
        RECT 29.750 129.635 29.925 130.085 ;
        RECT 30.095 129.815 30.425 130.255 ;
        RECT 30.730 129.665 30.900 130.085 ;
        RECT 31.135 129.845 31.805 130.255 ;
        RECT 32.020 129.665 32.190 130.085 ;
        RECT 32.390 129.845 32.720 130.255 ;
        RECT 29.750 129.465 30.380 129.635 ;
        RECT 28.725 129.035 29.480 129.205 ;
        RECT 27.765 128.695 28.905 128.865 ;
        RECT 29.075 128.525 29.480 129.035 ;
        RECT 29.665 128.615 30.030 129.295 ;
        RECT 30.210 128.945 30.380 129.465 ;
        RECT 30.730 129.495 32.745 129.665 ;
        RECT 30.210 128.615 30.560 128.945 ;
        RECT 27.830 128.355 29.480 128.525 ;
        RECT 30.210 128.445 30.380 128.615 ;
        RECT 26.905 127.875 27.205 128.205 ;
        RECT 27.375 127.705 27.650 128.185 ;
        RECT 27.830 127.965 28.125 128.355 ;
        RECT 28.295 127.705 28.550 128.185 ;
        RECT 28.725 127.965 28.985 128.355 ;
        RECT 29.750 128.275 30.380 128.445 ;
        RECT 29.155 127.705 29.435 128.185 ;
        RECT 29.750 127.875 29.925 128.275 ;
        RECT 30.730 128.205 30.900 129.495 ;
        RECT 30.095 127.705 30.425 128.085 ;
        RECT 30.670 127.875 30.900 128.205 ;
        RECT 31.100 128.040 31.380 129.315 ;
        RECT 31.605 129.235 31.875 129.315 ;
        RECT 31.565 129.065 31.875 129.235 ;
        RECT 31.605 128.040 31.875 129.065 ;
        RECT 32.065 128.285 32.405 129.315 ;
        RECT 32.575 128.945 32.745 129.495 ;
        RECT 32.915 129.115 33.175 130.085 ;
        RECT 33.430 129.635 33.605 130.085 ;
        RECT 33.775 129.815 34.105 130.255 ;
        RECT 34.410 129.665 34.580 130.085 ;
        RECT 34.815 129.845 35.485 130.255 ;
        RECT 35.700 129.665 35.870 130.085 ;
        RECT 36.070 129.845 36.400 130.255 ;
        RECT 33.430 129.465 34.060 129.635 ;
        RECT 32.575 128.615 32.835 128.945 ;
        RECT 33.005 128.425 33.175 129.115 ;
        RECT 33.345 128.615 33.710 129.295 ;
        RECT 33.890 128.945 34.060 129.465 ;
        RECT 34.410 129.495 36.425 129.665 ;
        RECT 33.890 128.615 34.240 128.945 ;
        RECT 33.890 128.445 34.060 128.615 ;
        RECT 32.335 127.705 32.665 128.085 ;
        RECT 32.835 127.960 33.175 128.425 ;
        RECT 33.430 128.275 34.060 128.445 ;
        RECT 32.835 127.915 33.170 127.960 ;
        RECT 33.430 127.875 33.605 128.275 ;
        RECT 34.410 128.205 34.580 129.495 ;
        RECT 33.775 127.705 34.105 128.085 ;
        RECT 34.350 127.875 34.580 128.205 ;
        RECT 34.780 128.040 35.060 129.315 ;
        RECT 35.285 128.215 35.555 129.315 ;
        RECT 35.745 128.285 36.085 129.315 ;
        RECT 36.255 128.945 36.425 129.495 ;
        RECT 36.595 129.115 36.855 130.085 ;
        RECT 37.030 129.875 37.365 130.255 ;
        RECT 36.255 128.615 36.515 128.945 ;
        RECT 36.685 128.425 36.855 129.115 ;
        RECT 35.245 128.045 35.555 128.215 ;
        RECT 35.285 128.040 35.555 128.045 ;
        RECT 36.015 127.705 36.345 128.085 ;
        RECT 36.515 127.960 36.855 128.425 ;
        RECT 37.025 128.385 37.265 129.695 ;
        RECT 37.535 129.285 37.785 130.085 ;
        RECT 38.005 129.535 38.335 130.255 ;
        RECT 38.520 129.285 38.770 130.085 ;
        RECT 39.235 129.455 39.565 130.255 ;
        RECT 39.735 129.825 40.075 130.085 ;
        RECT 37.435 129.115 39.625 129.285 ;
        RECT 37.435 128.205 37.605 129.115 ;
        RECT 39.310 128.945 39.625 129.115 ;
        RECT 36.515 127.915 36.850 127.960 ;
        RECT 37.110 127.875 37.605 128.205 ;
        RECT 37.825 127.980 38.175 128.945 ;
        RECT 38.355 127.975 38.655 128.945 ;
        RECT 38.835 127.975 39.115 128.945 ;
        RECT 39.310 128.695 39.640 128.945 ;
        RECT 39.295 127.705 39.565 128.505 ;
        RECT 39.815 128.425 40.075 129.825 ;
        RECT 40.245 129.745 40.545 130.255 ;
        RECT 40.715 129.575 41.045 130.085 ;
        RECT 41.215 129.745 41.845 130.255 ;
        RECT 42.425 129.745 42.805 129.915 ;
        RECT 42.975 129.745 43.275 130.255 ;
        RECT 42.635 129.575 42.805 129.745 ;
        RECT 39.735 127.915 40.075 128.425 ;
        RECT 40.245 129.405 42.465 129.575 ;
        RECT 40.245 128.445 40.415 129.405 ;
        RECT 40.585 129.065 42.125 129.235 ;
        RECT 40.585 128.615 40.830 129.065 ;
        RECT 41.090 128.695 41.785 128.895 ;
        RECT 41.955 128.865 42.125 129.065 ;
        RECT 42.295 129.205 42.465 129.405 ;
        RECT 42.635 129.375 43.295 129.575 ;
        RECT 42.295 129.035 42.955 129.205 ;
        RECT 41.955 128.695 42.555 128.865 ;
        RECT 42.785 128.615 42.955 129.035 ;
        RECT 40.245 127.900 40.710 128.445 ;
        RECT 41.215 127.705 41.385 128.525 ;
        RECT 41.555 128.445 42.465 128.525 ;
        RECT 43.125 128.445 43.295 129.375 ;
        RECT 43.525 129.195 43.855 130.040 ;
        RECT 44.025 129.245 44.195 130.255 ;
        RECT 44.365 129.525 44.705 130.085 ;
        RECT 44.935 129.755 45.250 130.255 ;
        RECT 45.430 129.785 46.315 129.955 ;
        RECT 41.555 128.355 42.805 128.445 ;
        RECT 41.555 127.875 41.885 128.355 ;
        RECT 42.295 128.275 42.805 128.355 ;
        RECT 42.055 127.705 42.405 128.095 ;
        RECT 42.575 127.875 42.805 128.275 ;
        RECT 42.975 127.965 43.295 128.445 ;
        RECT 43.465 129.115 43.855 129.195 ;
        RECT 44.365 129.150 45.260 129.525 ;
        RECT 43.465 129.065 43.680 129.115 ;
        RECT 43.465 128.485 43.635 129.065 ;
        RECT 44.365 128.945 44.555 129.150 ;
        RECT 45.430 128.945 45.600 129.785 ;
        RECT 46.540 129.755 46.790 130.085 ;
        RECT 43.805 128.615 44.555 128.945 ;
        RECT 44.725 128.615 45.600 128.945 ;
        RECT 43.465 128.445 43.690 128.485 ;
        RECT 44.355 128.445 44.555 128.615 ;
        RECT 43.465 128.360 43.845 128.445 ;
        RECT 43.515 127.925 43.845 128.360 ;
        RECT 44.015 127.705 44.185 128.315 ;
        RECT 44.355 127.920 44.685 128.445 ;
        RECT 44.945 127.705 45.155 128.235 ;
        RECT 45.430 128.155 45.600 128.615 ;
        RECT 45.770 128.655 46.090 129.615 ;
        RECT 46.260 128.865 46.450 129.585 ;
        RECT 46.620 128.685 46.790 129.755 ;
        RECT 46.960 129.455 47.130 130.255 ;
        RECT 47.300 129.810 48.405 129.980 ;
        RECT 47.300 129.195 47.470 129.810 ;
        RECT 48.615 129.660 48.865 130.085 ;
        RECT 49.035 129.795 49.300 130.255 ;
        RECT 47.640 129.275 48.170 129.640 ;
        RECT 48.615 129.530 48.920 129.660 ;
        RECT 46.960 129.105 47.470 129.195 ;
        RECT 46.960 128.935 47.830 129.105 ;
        RECT 46.960 128.865 47.130 128.935 ;
        RECT 47.250 128.685 47.450 128.715 ;
        RECT 45.770 128.325 46.235 128.655 ;
        RECT 46.620 128.385 47.450 128.685 ;
        RECT 46.620 128.155 46.790 128.385 ;
        RECT 45.430 127.985 46.215 128.155 ;
        RECT 46.385 127.985 46.790 128.155 ;
        RECT 46.970 127.705 47.340 128.205 ;
        RECT 47.660 128.155 47.830 128.935 ;
        RECT 48.000 128.575 48.170 129.275 ;
        RECT 48.340 128.745 48.580 129.340 ;
        RECT 48.000 128.355 48.525 128.575 ;
        RECT 48.750 128.425 48.920 129.530 ;
        RECT 48.695 128.295 48.920 128.425 ;
        RECT 49.090 128.335 49.370 129.285 ;
        RECT 48.695 128.155 48.865 128.295 ;
        RECT 47.660 127.985 48.335 128.155 ;
        RECT 48.530 127.985 48.865 128.155 ;
        RECT 49.035 127.705 49.285 128.165 ;
        RECT 49.540 127.965 49.725 130.085 ;
        RECT 49.895 129.755 50.225 130.255 ;
        RECT 50.395 129.585 50.565 130.085 ;
        RECT 49.900 129.415 50.565 129.585 ;
        RECT 49.900 128.425 50.130 129.415 ;
        RECT 50.300 128.595 50.650 129.245 ;
        RECT 50.825 129.090 51.115 130.255 ;
        RECT 51.285 129.165 53.875 130.255 ;
        RECT 51.285 128.475 52.495 128.995 ;
        RECT 52.665 128.645 53.875 129.165 ;
        RECT 54.565 129.115 54.775 130.255 ;
        RECT 54.945 129.105 55.275 130.085 ;
        RECT 55.445 129.115 55.675 130.255 ;
        RECT 55.885 129.115 56.165 130.255 ;
        RECT 56.335 129.105 56.665 130.085 ;
        RECT 56.835 129.115 57.095 130.255 ;
        RECT 57.270 129.115 57.605 130.085 ;
        RECT 57.775 129.115 57.945 130.255 ;
        RECT 58.115 129.915 60.145 130.085 ;
        RECT 49.900 128.255 50.565 128.425 ;
        RECT 49.895 127.705 50.225 128.085 ;
        RECT 50.395 127.965 50.565 128.255 ;
        RECT 50.825 127.705 51.115 128.430 ;
        RECT 51.285 127.705 53.875 128.475 ;
        RECT 54.565 127.705 54.775 128.525 ;
        RECT 54.945 128.505 55.195 129.105 ;
        RECT 55.365 128.695 55.695 128.945 ;
        RECT 55.895 128.675 56.230 128.945 ;
        RECT 56.400 128.555 56.570 129.105 ;
        RECT 56.740 128.695 57.075 128.945 ;
        RECT 54.945 127.875 55.275 128.505 ;
        RECT 55.445 127.705 55.675 128.525 ;
        RECT 56.400 128.505 56.575 128.555 ;
        RECT 55.885 127.705 56.195 128.505 ;
        RECT 56.400 127.875 57.095 128.505 ;
        RECT 57.270 128.445 57.440 129.115 ;
        RECT 58.115 128.945 58.285 129.915 ;
        RECT 57.610 128.615 57.865 128.945 ;
        RECT 58.090 128.615 58.285 128.945 ;
        RECT 58.455 129.575 59.580 129.745 ;
        RECT 57.695 128.445 57.865 128.615 ;
        RECT 58.455 128.445 58.625 129.575 ;
        RECT 57.270 127.875 57.525 128.445 ;
        RECT 57.695 128.275 58.625 128.445 ;
        RECT 58.795 129.235 59.805 129.405 ;
        RECT 58.795 128.435 58.965 129.235 ;
        RECT 58.450 128.240 58.625 128.275 ;
        RECT 57.695 127.705 58.025 128.105 ;
        RECT 58.450 127.875 58.980 128.240 ;
        RECT 59.170 128.215 59.445 129.035 ;
        RECT 59.165 128.045 59.445 128.215 ;
        RECT 59.170 127.875 59.445 128.045 ;
        RECT 59.615 127.875 59.805 129.235 ;
        RECT 59.975 129.250 60.145 129.915 ;
        RECT 60.315 129.495 60.485 130.255 ;
        RECT 60.720 129.495 61.235 129.905 ;
        RECT 59.975 129.060 60.725 129.250 ;
        RECT 60.895 128.685 61.235 129.495 ;
        RECT 61.410 129.105 61.670 130.255 ;
        RECT 61.845 129.180 62.100 130.085 ;
        RECT 62.270 129.495 62.600 130.255 ;
        RECT 62.815 129.325 62.985 130.085 ;
        RECT 60.005 128.515 61.235 128.685 ;
        RECT 59.985 127.705 60.495 128.240 ;
        RECT 60.715 127.910 60.960 128.515 ;
        RECT 61.410 127.705 61.670 128.545 ;
        RECT 61.845 128.450 62.015 129.180 ;
        RECT 62.270 129.155 62.985 129.325 ;
        RECT 62.270 128.945 62.440 129.155 ;
        RECT 63.245 129.115 63.505 130.255 ;
        RECT 63.675 129.105 64.005 130.085 ;
        RECT 64.175 129.115 64.455 130.255 ;
        RECT 64.625 129.115 64.885 130.255 ;
        RECT 65.055 129.105 65.385 130.085 ;
        RECT 65.555 129.115 65.835 130.255 ;
        RECT 66.525 129.195 66.855 130.040 ;
        RECT 67.025 129.245 67.195 130.255 ;
        RECT 67.365 129.525 67.705 130.085 ;
        RECT 67.935 129.755 68.250 130.255 ;
        RECT 68.430 129.785 69.315 129.955 ;
        RECT 66.465 129.115 66.855 129.195 ;
        RECT 67.365 129.150 68.260 129.525 ;
        RECT 62.185 128.615 62.440 128.945 ;
        RECT 61.845 127.875 62.100 128.450 ;
        RECT 62.270 128.425 62.440 128.615 ;
        RECT 62.720 128.605 63.075 128.975 ;
        RECT 63.265 128.695 63.600 128.945 ;
        RECT 63.770 128.505 63.940 129.105 ;
        RECT 64.110 128.675 64.445 128.945 ;
        RECT 64.645 128.695 64.980 128.945 ;
        RECT 65.150 128.505 65.320 129.105 ;
        RECT 66.465 129.065 66.680 129.115 ;
        RECT 65.490 128.675 65.825 128.945 ;
        RECT 62.270 128.255 62.985 128.425 ;
        RECT 62.270 127.705 62.600 128.085 ;
        RECT 62.815 127.875 62.985 128.255 ;
        RECT 63.245 127.875 63.940 128.505 ;
        RECT 64.145 127.705 64.455 128.505 ;
        RECT 64.625 127.875 65.320 128.505 ;
        RECT 65.525 127.705 65.835 128.505 ;
        RECT 66.465 128.485 66.635 129.065 ;
        RECT 67.365 128.945 67.555 129.150 ;
        RECT 68.430 128.945 68.600 129.785 ;
        RECT 69.540 129.755 69.790 130.085 ;
        RECT 66.805 128.615 67.555 128.945 ;
        RECT 67.725 128.615 68.600 128.945 ;
        RECT 66.465 128.445 66.690 128.485 ;
        RECT 67.355 128.445 67.555 128.615 ;
        RECT 66.465 128.360 66.845 128.445 ;
        RECT 66.515 127.925 66.845 128.360 ;
        RECT 67.015 127.705 67.185 128.315 ;
        RECT 67.355 127.920 67.685 128.445 ;
        RECT 67.945 127.705 68.155 128.235 ;
        RECT 68.430 128.155 68.600 128.615 ;
        RECT 68.770 128.655 69.090 129.615 ;
        RECT 69.260 128.865 69.450 129.585 ;
        RECT 69.620 128.685 69.790 129.755 ;
        RECT 69.960 129.455 70.130 130.255 ;
        RECT 70.300 129.810 71.405 129.980 ;
        RECT 70.300 129.195 70.470 129.810 ;
        RECT 71.615 129.660 71.865 130.085 ;
        RECT 72.035 129.795 72.300 130.255 ;
        RECT 70.640 129.275 71.170 129.640 ;
        RECT 71.615 129.530 71.920 129.660 ;
        RECT 69.960 129.105 70.470 129.195 ;
        RECT 69.960 128.935 70.830 129.105 ;
        RECT 69.960 128.865 70.130 128.935 ;
        RECT 70.250 128.685 70.450 128.715 ;
        RECT 68.770 128.325 69.235 128.655 ;
        RECT 69.620 128.385 70.450 128.685 ;
        RECT 69.620 128.155 69.790 128.385 ;
        RECT 68.430 127.985 69.215 128.155 ;
        RECT 69.385 127.985 69.790 128.155 ;
        RECT 69.970 127.705 70.340 128.205 ;
        RECT 70.660 128.155 70.830 128.935 ;
        RECT 71.000 128.575 71.170 129.275 ;
        RECT 71.340 128.745 71.580 129.340 ;
        RECT 71.000 128.355 71.525 128.575 ;
        RECT 71.750 128.425 71.920 129.530 ;
        RECT 71.695 128.295 71.920 128.425 ;
        RECT 72.090 128.335 72.370 129.285 ;
        RECT 71.695 128.155 71.865 128.295 ;
        RECT 70.660 127.985 71.335 128.155 ;
        RECT 71.530 127.985 71.865 128.155 ;
        RECT 72.035 127.705 72.285 128.165 ;
        RECT 72.540 127.965 72.725 130.085 ;
        RECT 72.895 129.755 73.225 130.255 ;
        RECT 73.395 129.585 73.565 130.085 ;
        RECT 72.900 129.415 73.565 129.585 ;
        RECT 72.900 128.425 73.130 129.415 ;
        RECT 74.470 129.285 74.860 129.460 ;
        RECT 75.345 129.455 75.675 130.255 ;
        RECT 75.845 129.465 76.380 130.085 ;
        RECT 73.300 128.595 73.650 129.245 ;
        RECT 74.470 129.115 75.895 129.285 ;
        RECT 72.900 128.255 73.565 128.425 ;
        RECT 74.345 128.385 74.700 128.945 ;
        RECT 72.895 127.705 73.225 128.085 ;
        RECT 73.395 127.965 73.565 128.255 ;
        RECT 74.870 128.215 75.040 129.115 ;
        RECT 75.210 128.385 75.475 128.945 ;
        RECT 75.725 128.615 75.895 129.115 ;
        RECT 76.065 128.445 76.380 129.465 ;
        RECT 76.585 129.090 76.875 130.255 ;
        RECT 77.045 129.115 77.385 130.085 ;
        RECT 77.555 129.115 77.725 130.255 ;
        RECT 77.995 129.455 78.245 130.255 ;
        RECT 78.890 129.285 79.220 130.085 ;
        RECT 79.520 129.455 79.850 130.255 ;
        RECT 80.020 129.285 80.350 130.085 ;
        RECT 77.915 129.115 80.350 129.285 ;
        RECT 80.930 129.285 81.260 130.085 ;
        RECT 81.430 129.455 81.760 130.255 ;
        RECT 82.060 129.285 82.390 130.085 ;
        RECT 83.035 129.455 83.285 130.255 ;
        RECT 80.930 129.115 83.365 129.285 ;
        RECT 83.555 129.115 83.725 130.255 ;
        RECT 83.895 129.115 84.235 130.085 ;
        RECT 74.450 127.705 74.690 128.215 ;
        RECT 74.870 127.885 75.150 128.215 ;
        RECT 75.380 127.705 75.595 128.215 ;
        RECT 75.765 127.875 76.380 128.445 ;
        RECT 77.045 128.505 77.220 129.115 ;
        RECT 77.915 128.865 78.085 129.115 ;
        RECT 77.390 128.695 78.085 128.865 ;
        RECT 78.260 128.695 78.680 128.895 ;
        RECT 78.850 128.695 79.180 128.895 ;
        RECT 79.350 128.695 79.680 128.895 ;
        RECT 76.585 127.705 76.875 128.430 ;
        RECT 77.045 127.875 77.385 128.505 ;
        RECT 77.555 127.705 77.805 128.505 ;
        RECT 77.995 128.355 79.220 128.525 ;
        RECT 77.995 127.875 78.325 128.355 ;
        RECT 78.495 127.705 78.720 128.165 ;
        RECT 78.890 127.875 79.220 128.355 ;
        RECT 79.850 128.485 80.020 129.115 ;
        RECT 80.205 128.695 80.555 128.945 ;
        RECT 80.725 128.695 81.075 128.945 ;
        RECT 81.260 128.485 81.430 129.115 ;
        RECT 81.600 128.695 81.930 128.895 ;
        RECT 82.100 128.695 82.430 128.895 ;
        RECT 82.600 128.695 83.020 128.895 ;
        RECT 83.195 128.865 83.365 129.115 ;
        RECT 83.195 128.695 83.890 128.865 ;
        RECT 79.850 127.875 80.350 128.485 ;
        RECT 80.930 127.875 81.430 128.485 ;
        RECT 82.060 128.355 83.285 128.525 ;
        RECT 84.060 128.505 84.235 129.115 ;
        RECT 82.060 127.875 82.390 128.355 ;
        RECT 82.560 127.705 82.785 128.165 ;
        RECT 82.955 127.875 83.285 128.355 ;
        RECT 83.475 127.705 83.725 128.505 ;
        RECT 83.895 127.875 84.235 128.505 ;
        RECT 84.405 129.405 84.665 130.085 ;
        RECT 84.835 129.475 85.085 130.255 ;
        RECT 85.335 129.705 85.585 130.085 ;
        RECT 85.755 129.875 86.110 130.255 ;
        RECT 87.115 129.865 87.450 130.085 ;
        RECT 86.715 129.705 86.945 129.745 ;
        RECT 85.335 129.505 86.945 129.705 ;
        RECT 85.335 129.495 86.170 129.505 ;
        RECT 86.760 129.415 86.945 129.505 ;
        RECT 84.405 128.205 84.575 129.405 ;
        RECT 86.275 129.305 86.605 129.335 ;
        RECT 84.805 129.245 86.605 129.305 ;
        RECT 87.195 129.245 87.450 129.865 ;
        RECT 84.745 129.135 87.450 129.245 ;
        RECT 84.745 129.100 84.945 129.135 ;
        RECT 84.745 128.525 84.915 129.100 ;
        RECT 86.275 129.075 87.450 129.135 ;
        RECT 88.545 129.165 89.755 130.255 ;
        RECT 100.140 129.320 100.810 131.580 ;
        RECT 101.480 131.010 105.520 131.180 ;
        RECT 101.140 129.950 101.310 130.950 ;
        RECT 105.690 129.950 105.860 130.950 ;
        RECT 101.480 129.720 105.520 129.890 ;
        RECT 106.200 129.320 106.370 131.580 ;
        RECT 85.145 128.660 85.555 128.965 ;
        RECT 85.725 128.695 86.055 128.905 ;
        RECT 84.745 128.405 85.015 128.525 ;
        RECT 84.745 128.360 85.590 128.405 ;
        RECT 84.835 128.235 85.590 128.360 ;
        RECT 85.845 128.295 86.055 128.695 ;
        RECT 86.300 128.695 86.775 128.905 ;
        RECT 86.965 128.695 87.455 128.895 ;
        RECT 86.300 128.295 86.520 128.695 ;
        RECT 88.545 128.625 89.065 129.165 ;
        RECT 100.140 129.150 106.370 129.320 ;
        RECT 84.405 127.875 84.665 128.205 ;
        RECT 85.420 128.085 85.590 128.235 ;
        RECT 84.835 127.705 85.165 128.065 ;
        RECT 85.420 127.875 86.720 128.085 ;
        RECT 86.995 127.705 87.450 128.470 ;
        RECT 89.235 128.455 89.755 128.995 ;
        RECT 88.545 127.705 89.755 128.455 ;
        RECT 12.100 127.535 89.840 127.705 ;
        RECT 12.185 126.785 13.395 127.535 ;
        RECT 13.655 126.985 13.825 127.275 ;
        RECT 13.995 127.155 14.325 127.535 ;
        RECT 13.655 126.815 14.320 126.985 ;
        RECT 12.185 126.245 12.705 126.785 ;
        RECT 12.875 126.075 13.395 126.615 ;
        RECT 12.185 124.985 13.395 126.075 ;
        RECT 13.570 125.995 13.920 126.645 ;
        RECT 14.090 125.825 14.320 126.815 ;
        RECT 13.655 125.655 14.320 125.825 ;
        RECT 13.655 125.155 13.825 125.655 ;
        RECT 13.995 124.985 14.325 125.485 ;
        RECT 14.495 125.155 14.680 127.275 ;
        RECT 14.935 127.075 15.185 127.535 ;
        RECT 15.355 127.085 15.690 127.255 ;
        RECT 15.885 127.085 16.560 127.255 ;
        RECT 15.355 126.945 15.525 127.085 ;
        RECT 14.850 125.955 15.130 126.905 ;
        RECT 15.300 126.815 15.525 126.945 ;
        RECT 15.300 125.710 15.470 126.815 ;
        RECT 15.695 126.665 16.220 126.885 ;
        RECT 15.640 125.900 15.880 126.495 ;
        RECT 16.050 125.965 16.220 126.665 ;
        RECT 16.390 126.305 16.560 127.085 ;
        RECT 16.880 127.035 17.250 127.535 ;
        RECT 17.430 127.085 17.835 127.255 ;
        RECT 18.005 127.085 18.790 127.255 ;
        RECT 17.430 126.855 17.600 127.085 ;
        RECT 16.770 126.555 17.600 126.855 ;
        RECT 17.985 126.585 18.450 126.915 ;
        RECT 16.770 126.525 16.970 126.555 ;
        RECT 17.090 126.305 17.260 126.375 ;
        RECT 16.390 126.135 17.260 126.305 ;
        RECT 16.750 126.045 17.260 126.135 ;
        RECT 15.300 125.580 15.605 125.710 ;
        RECT 16.050 125.600 16.580 125.965 ;
        RECT 14.920 124.985 15.185 125.445 ;
        RECT 15.355 125.155 15.605 125.580 ;
        RECT 16.750 125.430 16.920 126.045 ;
        RECT 15.815 125.260 16.920 125.430 ;
        RECT 17.090 124.985 17.260 125.785 ;
        RECT 17.430 125.485 17.600 126.555 ;
        RECT 17.770 125.655 17.960 126.375 ;
        RECT 18.130 125.625 18.450 126.585 ;
        RECT 18.620 126.625 18.790 127.085 ;
        RECT 19.065 127.005 19.275 127.535 ;
        RECT 19.535 126.795 19.865 127.320 ;
        RECT 20.035 126.925 20.205 127.535 ;
        RECT 20.375 126.880 20.705 127.315 ;
        RECT 20.375 126.795 20.755 126.880 ;
        RECT 19.665 126.625 19.865 126.795 ;
        RECT 20.530 126.755 20.755 126.795 ;
        RECT 18.620 126.295 19.495 126.625 ;
        RECT 19.665 126.295 20.415 126.625 ;
        RECT 17.430 125.155 17.680 125.485 ;
        RECT 18.620 125.455 18.790 126.295 ;
        RECT 19.665 126.090 19.855 126.295 ;
        RECT 20.585 126.175 20.755 126.755 ;
        RECT 20.945 126.725 21.185 127.535 ;
        RECT 21.355 126.725 21.685 127.365 ;
        RECT 21.855 126.725 22.125 127.535 ;
        RECT 22.510 126.755 23.010 127.365 ;
        RECT 20.925 126.295 21.275 126.545 ;
        RECT 20.540 126.125 20.755 126.175 ;
        RECT 21.445 126.125 21.615 126.725 ;
        RECT 21.785 126.295 22.135 126.545 ;
        RECT 22.305 126.295 22.655 126.545 ;
        RECT 22.840 126.125 23.010 126.755 ;
        RECT 23.640 126.885 23.970 127.365 ;
        RECT 24.140 127.075 24.365 127.535 ;
        RECT 24.535 126.885 24.865 127.365 ;
        RECT 23.640 126.715 24.865 126.885 ;
        RECT 25.055 126.735 25.305 127.535 ;
        RECT 25.475 126.735 25.815 127.365 ;
        RECT 23.180 126.345 23.510 126.545 ;
        RECT 23.680 126.345 24.010 126.545 ;
        RECT 24.180 126.345 24.600 126.545 ;
        RECT 24.775 126.375 25.470 126.545 ;
        RECT 24.775 126.125 24.945 126.375 ;
        RECT 25.640 126.125 25.815 126.735 ;
        RECT 18.960 125.715 19.855 126.090 ;
        RECT 20.365 126.045 20.755 126.125 ;
        RECT 17.905 125.285 18.790 125.455 ;
        RECT 18.970 124.985 19.285 125.485 ;
        RECT 19.515 125.155 19.855 125.715 ;
        RECT 20.025 124.985 20.195 125.995 ;
        RECT 20.365 125.200 20.695 126.045 ;
        RECT 20.935 125.955 21.615 126.125 ;
        RECT 20.935 125.170 21.265 125.955 ;
        RECT 21.795 124.985 22.125 126.125 ;
        RECT 22.510 125.955 24.945 126.125 ;
        RECT 22.510 125.155 22.840 125.955 ;
        RECT 23.010 124.985 23.340 125.785 ;
        RECT 23.640 125.155 23.970 125.955 ;
        RECT 24.615 124.985 24.865 125.785 ;
        RECT 25.135 124.985 25.305 126.125 ;
        RECT 25.475 125.155 25.815 126.125 ;
        RECT 26.445 125.155 26.725 127.255 ;
        RECT 26.955 127.075 27.125 127.535 ;
        RECT 27.395 127.145 28.645 127.325 ;
        RECT 27.780 126.905 28.145 126.975 ;
        RECT 26.895 126.725 28.145 126.905 ;
        RECT 28.315 126.925 28.645 127.145 ;
        RECT 28.815 127.095 28.985 127.535 ;
        RECT 29.155 126.925 29.495 127.340 ;
        RECT 28.315 126.755 29.495 126.925 ;
        RECT 30.675 126.985 30.845 127.275 ;
        RECT 31.015 127.155 31.345 127.535 ;
        RECT 30.675 126.815 31.340 126.985 ;
        RECT 26.895 126.125 27.170 126.725 ;
        RECT 27.340 126.295 27.695 126.545 ;
        RECT 27.890 126.515 28.355 126.545 ;
        RECT 27.885 126.345 28.355 126.515 ;
        RECT 27.890 126.295 28.355 126.345 ;
        RECT 28.525 126.295 28.855 126.545 ;
        RECT 29.030 126.345 29.495 126.545 ;
        RECT 28.675 126.175 28.855 126.295 ;
        RECT 26.895 125.915 28.505 126.125 ;
        RECT 28.675 126.005 29.005 126.175 ;
        RECT 28.095 125.815 28.505 125.915 ;
        RECT 26.915 124.985 27.700 125.745 ;
        RECT 28.095 125.155 28.480 125.815 ;
        RECT 28.805 125.215 29.005 126.005 ;
        RECT 29.175 124.985 29.495 126.165 ;
        RECT 30.590 125.995 30.940 126.645 ;
        RECT 31.110 125.825 31.340 126.815 ;
        RECT 30.675 125.655 31.340 125.825 ;
        RECT 30.675 125.155 30.845 125.655 ;
        RECT 31.015 124.985 31.345 125.485 ;
        RECT 31.515 125.155 31.700 127.275 ;
        RECT 31.955 127.075 32.205 127.535 ;
        RECT 32.375 127.085 32.710 127.255 ;
        RECT 32.905 127.085 33.580 127.255 ;
        RECT 32.375 126.945 32.545 127.085 ;
        RECT 31.870 125.955 32.150 126.905 ;
        RECT 32.320 126.815 32.545 126.945 ;
        RECT 32.320 125.710 32.490 126.815 ;
        RECT 32.715 126.665 33.240 126.885 ;
        RECT 32.660 125.900 32.900 126.495 ;
        RECT 33.070 125.965 33.240 126.665 ;
        RECT 33.410 126.305 33.580 127.085 ;
        RECT 33.900 127.035 34.270 127.535 ;
        RECT 34.450 127.085 34.855 127.255 ;
        RECT 35.025 127.085 35.810 127.255 ;
        RECT 34.450 126.855 34.620 127.085 ;
        RECT 33.790 126.555 34.620 126.855 ;
        RECT 35.005 126.585 35.470 126.915 ;
        RECT 33.790 126.525 33.990 126.555 ;
        RECT 34.110 126.305 34.280 126.375 ;
        RECT 33.410 126.135 34.280 126.305 ;
        RECT 33.770 126.045 34.280 126.135 ;
        RECT 32.320 125.580 32.625 125.710 ;
        RECT 33.070 125.600 33.600 125.965 ;
        RECT 31.940 124.985 32.205 125.445 ;
        RECT 32.375 125.155 32.625 125.580 ;
        RECT 33.770 125.430 33.940 126.045 ;
        RECT 32.835 125.260 33.940 125.430 ;
        RECT 34.110 124.985 34.280 125.785 ;
        RECT 34.450 125.485 34.620 126.555 ;
        RECT 34.790 125.655 34.980 126.375 ;
        RECT 35.150 125.625 35.470 126.585 ;
        RECT 35.640 126.625 35.810 127.085 ;
        RECT 36.085 127.005 36.295 127.535 ;
        RECT 36.555 126.795 36.885 127.320 ;
        RECT 37.055 126.925 37.225 127.535 ;
        RECT 37.395 126.880 37.725 127.315 ;
        RECT 37.395 126.795 37.775 126.880 ;
        RECT 37.945 126.810 38.235 127.535 ;
        RECT 38.405 126.990 43.750 127.535 ;
        RECT 43.925 126.990 49.270 127.535 ;
        RECT 36.685 126.625 36.885 126.795 ;
        RECT 37.550 126.755 37.775 126.795 ;
        RECT 35.640 126.295 36.515 126.625 ;
        RECT 36.685 126.295 37.435 126.625 ;
        RECT 34.450 125.155 34.700 125.485 ;
        RECT 35.640 125.455 35.810 126.295 ;
        RECT 36.685 126.090 36.875 126.295 ;
        RECT 37.605 126.175 37.775 126.755 ;
        RECT 37.560 126.125 37.775 126.175 ;
        RECT 39.990 126.160 40.330 126.990 ;
        RECT 35.980 125.715 36.875 126.090 ;
        RECT 37.385 126.045 37.775 126.125 ;
        RECT 34.925 125.285 35.810 125.455 ;
        RECT 35.990 124.985 36.305 125.485 ;
        RECT 36.535 125.155 36.875 125.715 ;
        RECT 37.045 124.985 37.215 125.995 ;
        RECT 37.385 125.200 37.715 126.045 ;
        RECT 37.945 124.985 38.235 126.150 ;
        RECT 41.810 125.420 42.160 126.670 ;
        RECT 45.510 126.160 45.850 126.990 ;
        RECT 49.445 126.765 52.035 127.535 ;
        RECT 52.755 126.985 52.925 127.275 ;
        RECT 53.095 127.155 53.425 127.535 ;
        RECT 52.755 126.815 53.420 126.985 ;
        RECT 47.330 125.420 47.680 126.670 ;
        RECT 49.445 126.245 50.655 126.765 ;
        RECT 50.825 126.075 52.035 126.595 ;
        RECT 38.405 124.985 43.750 125.420 ;
        RECT 43.925 124.985 49.270 125.420 ;
        RECT 49.445 124.985 52.035 126.075 ;
        RECT 52.670 125.995 53.020 126.645 ;
        RECT 53.190 125.825 53.420 126.815 ;
        RECT 52.755 125.655 53.420 125.825 ;
        RECT 52.755 125.155 52.925 125.655 ;
        RECT 53.095 124.985 53.425 125.485 ;
        RECT 53.595 125.155 53.780 127.275 ;
        RECT 54.035 127.075 54.285 127.535 ;
        RECT 54.455 127.085 54.790 127.255 ;
        RECT 54.985 127.085 55.660 127.255 ;
        RECT 54.455 126.945 54.625 127.085 ;
        RECT 53.950 125.955 54.230 126.905 ;
        RECT 54.400 126.815 54.625 126.945 ;
        RECT 54.400 125.710 54.570 126.815 ;
        RECT 54.795 126.665 55.320 126.885 ;
        RECT 54.740 125.900 54.980 126.495 ;
        RECT 55.150 125.965 55.320 126.665 ;
        RECT 55.490 126.305 55.660 127.085 ;
        RECT 55.980 127.035 56.350 127.535 ;
        RECT 56.530 127.085 56.935 127.255 ;
        RECT 57.105 127.085 57.890 127.255 ;
        RECT 56.530 126.855 56.700 127.085 ;
        RECT 55.870 126.555 56.700 126.855 ;
        RECT 57.085 126.585 57.550 126.915 ;
        RECT 55.870 126.525 56.070 126.555 ;
        RECT 56.190 126.305 56.360 126.375 ;
        RECT 55.490 126.135 56.360 126.305 ;
        RECT 55.850 126.045 56.360 126.135 ;
        RECT 54.400 125.580 54.705 125.710 ;
        RECT 55.150 125.600 55.680 125.965 ;
        RECT 54.020 124.985 54.285 125.445 ;
        RECT 54.455 125.155 54.705 125.580 ;
        RECT 55.850 125.430 56.020 126.045 ;
        RECT 54.915 125.260 56.020 125.430 ;
        RECT 56.190 124.985 56.360 125.785 ;
        RECT 56.530 125.485 56.700 126.555 ;
        RECT 56.870 125.655 57.060 126.375 ;
        RECT 57.230 125.625 57.550 126.585 ;
        RECT 57.720 126.625 57.890 127.085 ;
        RECT 58.165 127.005 58.375 127.535 ;
        RECT 58.635 126.795 58.965 127.320 ;
        RECT 59.135 126.925 59.305 127.535 ;
        RECT 59.475 126.880 59.805 127.315 ;
        RECT 60.140 126.905 60.425 127.365 ;
        RECT 60.595 127.075 60.865 127.535 ;
        RECT 59.475 126.795 59.855 126.880 ;
        RECT 58.765 126.625 58.965 126.795 ;
        RECT 59.630 126.755 59.855 126.795 ;
        RECT 57.720 126.295 58.595 126.625 ;
        RECT 58.765 126.295 59.515 126.625 ;
        RECT 56.530 125.155 56.780 125.485 ;
        RECT 57.720 125.455 57.890 126.295 ;
        RECT 58.765 126.090 58.955 126.295 ;
        RECT 59.685 126.175 59.855 126.755 ;
        RECT 60.140 126.735 61.095 126.905 ;
        RECT 59.640 126.125 59.855 126.175 ;
        RECT 58.060 125.715 58.955 126.090 ;
        RECT 59.465 126.045 59.855 126.125 ;
        RECT 57.005 125.285 57.890 125.455 ;
        RECT 58.070 124.985 58.385 125.485 ;
        RECT 58.615 125.155 58.955 125.715 ;
        RECT 59.125 124.985 59.295 125.995 ;
        RECT 59.465 125.200 59.795 126.045 ;
        RECT 60.025 126.005 60.715 126.565 ;
        RECT 60.885 125.835 61.095 126.735 ;
        RECT 60.140 125.615 61.095 125.835 ;
        RECT 61.265 126.565 61.665 127.365 ;
        RECT 61.855 126.905 62.135 127.365 ;
        RECT 62.655 127.075 62.980 127.535 ;
        RECT 61.855 126.735 62.980 126.905 ;
        RECT 63.150 126.795 63.535 127.365 ;
        RECT 63.705 126.810 63.995 127.535 ;
        RECT 64.165 127.035 64.425 127.365 ;
        RECT 64.595 127.175 64.925 127.535 ;
        RECT 65.180 127.155 66.480 127.365 ;
        RECT 62.530 126.625 62.980 126.735 ;
        RECT 61.265 126.005 62.360 126.565 ;
        RECT 62.530 126.295 63.085 126.625 ;
        RECT 60.140 125.155 60.425 125.615 ;
        RECT 60.595 124.985 60.865 125.445 ;
        RECT 61.265 125.155 61.665 126.005 ;
        RECT 62.530 125.835 62.980 126.295 ;
        RECT 63.255 126.125 63.535 126.795 ;
        RECT 61.855 125.615 62.980 125.835 ;
        RECT 61.855 125.155 62.135 125.615 ;
        RECT 62.655 124.985 62.980 125.445 ;
        RECT 63.150 125.155 63.535 126.125 ;
        RECT 63.705 124.985 63.995 126.150 ;
        RECT 64.165 125.835 64.335 127.035 ;
        RECT 65.180 127.005 65.350 127.155 ;
        RECT 64.595 126.880 65.350 127.005 ;
        RECT 64.505 126.835 65.350 126.880 ;
        RECT 64.505 126.715 64.775 126.835 ;
        RECT 64.505 126.140 64.675 126.715 ;
        RECT 64.905 126.275 65.315 126.580 ;
        RECT 65.605 126.545 65.815 126.945 ;
        RECT 65.485 126.335 65.815 126.545 ;
        RECT 66.060 126.545 66.280 126.945 ;
        RECT 66.755 126.770 67.210 127.535 ;
        RECT 67.390 126.695 67.650 127.535 ;
        RECT 67.825 126.790 68.080 127.365 ;
        RECT 68.250 127.155 68.580 127.535 ;
        RECT 68.795 126.985 68.965 127.365 ;
        RECT 68.250 126.815 68.965 126.985 ;
        RECT 66.060 126.335 66.535 126.545 ;
        RECT 66.725 126.345 67.215 126.545 ;
        RECT 64.505 126.105 64.705 126.140 ;
        RECT 66.035 126.105 67.210 126.165 ;
        RECT 64.505 125.995 67.210 126.105 ;
        RECT 64.565 125.935 66.365 125.995 ;
        RECT 66.035 125.905 66.365 125.935 ;
        RECT 64.165 125.155 64.425 125.835 ;
        RECT 64.595 124.985 64.845 125.765 ;
        RECT 65.095 125.735 65.930 125.745 ;
        RECT 66.520 125.735 66.705 125.825 ;
        RECT 65.095 125.535 66.705 125.735 ;
        RECT 65.095 125.155 65.345 125.535 ;
        RECT 66.475 125.495 66.705 125.535 ;
        RECT 66.955 125.375 67.210 125.995 ;
        RECT 65.515 124.985 65.870 125.365 ;
        RECT 66.875 125.155 67.210 125.375 ;
        RECT 67.390 124.985 67.650 126.135 ;
        RECT 67.825 126.060 67.995 126.790 ;
        RECT 68.250 126.625 68.420 126.815 ;
        RECT 69.230 126.770 69.685 127.535 ;
        RECT 69.960 127.155 71.260 127.365 ;
        RECT 71.515 127.175 71.845 127.535 ;
        RECT 71.090 127.005 71.260 127.155 ;
        RECT 72.015 127.035 72.275 127.365 ;
        RECT 72.045 127.025 72.275 127.035 ;
        RECT 68.165 126.295 68.420 126.625 ;
        RECT 68.250 126.085 68.420 126.295 ;
        RECT 68.700 126.265 69.055 126.635 ;
        RECT 70.160 126.545 70.380 126.945 ;
        RECT 69.225 126.345 69.715 126.545 ;
        RECT 69.905 126.335 70.380 126.545 ;
        RECT 70.625 126.545 70.835 126.945 ;
        RECT 71.090 126.880 71.845 127.005 ;
        RECT 71.090 126.835 71.935 126.880 ;
        RECT 71.665 126.715 71.935 126.835 ;
        RECT 70.625 126.335 70.955 126.545 ;
        RECT 71.125 126.275 71.535 126.580 ;
        RECT 69.230 126.105 70.405 126.165 ;
        RECT 71.765 126.140 71.935 126.715 ;
        RECT 71.735 126.105 71.935 126.140 ;
        RECT 67.825 125.155 68.080 126.060 ;
        RECT 68.250 125.915 68.965 126.085 ;
        RECT 68.250 124.985 68.580 125.745 ;
        RECT 68.795 125.155 68.965 125.915 ;
        RECT 69.230 125.995 71.935 126.105 ;
        RECT 69.230 125.375 69.485 125.995 ;
        RECT 70.075 125.935 71.875 125.995 ;
        RECT 70.075 125.905 70.405 125.935 ;
        RECT 72.105 125.835 72.275 127.025 ;
        RECT 72.535 126.985 72.705 127.275 ;
        RECT 72.875 127.155 73.205 127.535 ;
        RECT 72.535 126.815 73.200 126.985 ;
        RECT 72.450 125.995 72.800 126.645 ;
        RECT 69.735 125.735 69.920 125.825 ;
        RECT 70.510 125.735 71.345 125.745 ;
        RECT 69.735 125.535 71.345 125.735 ;
        RECT 69.735 125.495 69.965 125.535 ;
        RECT 69.230 125.155 69.565 125.375 ;
        RECT 70.570 124.985 70.925 125.365 ;
        RECT 71.095 125.155 71.345 125.535 ;
        RECT 71.595 124.985 71.845 125.765 ;
        RECT 72.015 125.155 72.275 125.835 ;
        RECT 72.970 125.825 73.200 126.815 ;
        RECT 72.535 125.655 73.200 125.825 ;
        RECT 72.535 125.155 72.705 125.655 ;
        RECT 72.875 124.985 73.205 125.485 ;
        RECT 73.375 125.155 73.560 127.275 ;
        RECT 73.815 127.075 74.065 127.535 ;
        RECT 74.235 127.085 74.570 127.255 ;
        RECT 74.765 127.085 75.440 127.255 ;
        RECT 74.235 126.945 74.405 127.085 ;
        RECT 73.730 125.955 74.010 126.905 ;
        RECT 74.180 126.815 74.405 126.945 ;
        RECT 74.180 125.710 74.350 126.815 ;
        RECT 74.575 126.665 75.100 126.885 ;
        RECT 74.520 125.900 74.760 126.495 ;
        RECT 74.930 125.965 75.100 126.665 ;
        RECT 75.270 126.305 75.440 127.085 ;
        RECT 75.760 127.035 76.130 127.535 ;
        RECT 76.310 127.085 76.715 127.255 ;
        RECT 76.885 127.085 77.670 127.255 ;
        RECT 76.310 126.855 76.480 127.085 ;
        RECT 75.650 126.555 76.480 126.855 ;
        RECT 76.865 126.585 77.330 126.915 ;
        RECT 75.650 126.525 75.850 126.555 ;
        RECT 75.970 126.305 76.140 126.375 ;
        RECT 75.270 126.135 76.140 126.305 ;
        RECT 75.630 126.045 76.140 126.135 ;
        RECT 74.180 125.580 74.485 125.710 ;
        RECT 74.930 125.600 75.460 125.965 ;
        RECT 73.800 124.985 74.065 125.445 ;
        RECT 74.235 125.155 74.485 125.580 ;
        RECT 75.630 125.430 75.800 126.045 ;
        RECT 74.695 125.260 75.800 125.430 ;
        RECT 75.970 124.985 76.140 125.785 ;
        RECT 76.310 125.485 76.480 126.555 ;
        RECT 76.650 125.655 76.840 126.375 ;
        RECT 77.010 125.625 77.330 126.585 ;
        RECT 77.500 126.625 77.670 127.085 ;
        RECT 77.945 127.005 78.155 127.535 ;
        RECT 78.415 126.795 78.745 127.320 ;
        RECT 78.915 126.925 79.085 127.535 ;
        RECT 79.255 126.880 79.585 127.315 ;
        RECT 79.970 127.025 80.210 127.535 ;
        RECT 80.390 127.025 80.670 127.355 ;
        RECT 80.900 127.025 81.115 127.535 ;
        RECT 79.255 126.795 79.635 126.880 ;
        RECT 78.545 126.625 78.745 126.795 ;
        RECT 79.410 126.755 79.635 126.795 ;
        RECT 77.500 126.295 78.375 126.625 ;
        RECT 78.545 126.295 79.295 126.625 ;
        RECT 76.310 125.155 76.560 125.485 ;
        RECT 77.500 125.455 77.670 126.295 ;
        RECT 78.545 126.090 78.735 126.295 ;
        RECT 79.465 126.175 79.635 126.755 ;
        RECT 79.865 126.295 80.220 126.855 ;
        RECT 79.420 126.125 79.635 126.175 ;
        RECT 80.390 126.125 80.560 127.025 ;
        RECT 80.730 126.295 80.995 126.855 ;
        RECT 81.285 126.795 81.900 127.365 ;
        RECT 81.245 126.125 81.415 126.625 ;
        RECT 77.840 125.715 78.735 126.090 ;
        RECT 79.245 126.045 79.635 126.125 ;
        RECT 76.785 125.285 77.670 125.455 ;
        RECT 77.850 124.985 78.165 125.485 ;
        RECT 78.395 125.155 78.735 125.715 ;
        RECT 78.905 124.985 79.075 125.995 ;
        RECT 79.245 125.200 79.575 126.045 ;
        RECT 79.990 125.955 81.415 126.125 ;
        RECT 79.990 125.780 80.380 125.955 ;
        RECT 80.865 124.985 81.195 125.785 ;
        RECT 81.585 125.775 81.900 126.795 ;
        RECT 82.110 126.770 82.565 127.535 ;
        RECT 82.840 127.155 84.140 127.365 ;
        RECT 84.395 127.175 84.725 127.535 ;
        RECT 83.970 127.005 84.140 127.155 ;
        RECT 84.895 127.035 85.155 127.365 ;
        RECT 83.040 126.545 83.260 126.945 ;
        RECT 82.105 126.345 82.595 126.545 ;
        RECT 82.785 126.335 83.260 126.545 ;
        RECT 83.505 126.545 83.715 126.945 ;
        RECT 83.970 126.880 84.725 127.005 ;
        RECT 83.970 126.835 84.815 126.880 ;
        RECT 84.545 126.715 84.815 126.835 ;
        RECT 83.505 126.335 83.835 126.545 ;
        RECT 84.005 126.275 84.415 126.580 ;
        RECT 81.365 125.155 81.900 125.775 ;
        RECT 82.110 126.105 83.285 126.165 ;
        RECT 84.645 126.140 84.815 126.715 ;
        RECT 84.615 126.105 84.815 126.140 ;
        RECT 82.110 125.995 84.815 126.105 ;
        RECT 82.110 125.375 82.365 125.995 ;
        RECT 82.955 125.935 84.755 125.995 ;
        RECT 82.955 125.905 83.285 125.935 ;
        RECT 84.985 125.835 85.155 127.035 ;
        RECT 82.615 125.735 82.800 125.825 ;
        RECT 83.390 125.735 84.225 125.745 ;
        RECT 82.615 125.535 84.225 125.735 ;
        RECT 82.615 125.495 82.845 125.535 ;
        RECT 82.110 125.155 82.445 125.375 ;
        RECT 83.450 124.985 83.805 125.365 ;
        RECT 83.975 125.155 84.225 125.535 ;
        RECT 84.475 124.985 84.725 125.765 ;
        RECT 84.895 125.155 85.155 125.835 ;
        RECT 85.360 126.795 85.975 127.365 ;
        RECT 86.145 127.025 86.360 127.535 ;
        RECT 86.590 127.025 86.870 127.355 ;
        RECT 87.050 127.025 87.290 127.535 ;
        RECT 85.360 125.775 85.675 126.795 ;
        RECT 85.845 126.125 86.015 126.625 ;
        RECT 86.265 126.295 86.530 126.855 ;
        RECT 86.700 126.125 86.870 127.025 ;
        RECT 87.040 126.295 87.395 126.855 ;
        RECT 88.545 126.785 89.755 127.535 ;
        RECT 85.845 125.955 87.270 126.125 ;
        RECT 85.360 125.155 85.895 125.775 ;
        RECT 86.065 124.985 86.395 125.785 ;
        RECT 86.880 125.780 87.270 125.955 ;
        RECT 88.545 126.075 89.065 126.615 ;
        RECT 89.235 126.245 89.755 126.785 ;
        RECT 88.545 124.985 89.755 126.075 ;
        RECT 100.140 125.890 100.810 129.150 ;
        RECT 101.480 128.580 105.520 128.750 ;
        RECT 101.140 126.520 101.310 128.520 ;
        RECT 105.690 126.520 105.860 128.520 ;
        RECT 101.480 126.290 105.520 126.460 ;
        RECT 106.200 125.890 106.370 129.150 ;
        RECT 100.140 125.720 106.370 125.890 ;
        RECT 12.100 124.815 89.840 124.985 ;
        RECT 12.185 123.725 13.395 124.815 ;
        RECT 12.185 123.015 12.705 123.555 ;
        RECT 12.875 123.185 13.395 123.725 ;
        RECT 14.485 123.675 14.745 124.645 ;
        RECT 14.940 124.405 15.270 124.815 ;
        RECT 15.470 124.225 15.640 124.645 ;
        RECT 15.855 124.405 16.525 124.815 ;
        RECT 16.760 124.225 16.930 124.645 ;
        RECT 17.235 124.375 17.565 124.815 ;
        RECT 14.915 124.055 16.930 124.225 ;
        RECT 17.735 124.195 17.910 124.645 ;
        RECT 12.185 122.265 13.395 123.015 ;
        RECT 14.485 122.985 14.655 123.675 ;
        RECT 14.915 123.505 15.085 124.055 ;
        RECT 14.825 123.175 15.085 123.505 ;
        RECT 14.485 122.520 14.825 122.985 ;
        RECT 15.255 122.845 15.595 123.875 ;
        RECT 15.785 123.455 16.055 123.875 ;
        RECT 15.785 123.285 16.095 123.455 ;
        RECT 14.490 122.475 14.825 122.520 ;
        RECT 14.995 122.265 15.325 122.645 ;
        RECT 15.785 122.600 16.055 123.285 ;
        RECT 16.280 122.600 16.560 123.875 ;
        RECT 16.760 122.765 16.930 124.055 ;
        RECT 17.280 124.025 17.910 124.195 ;
        RECT 17.280 123.505 17.450 124.025 ;
        RECT 17.100 123.175 17.450 123.505 ;
        RECT 17.630 123.175 17.995 123.855 ;
        RECT 18.175 123.845 18.505 124.630 ;
        RECT 18.175 123.675 18.855 123.845 ;
        RECT 19.035 123.675 19.365 124.815 ;
        RECT 19.545 124.385 19.885 124.645 ;
        RECT 18.165 123.255 18.515 123.505 ;
        RECT 17.280 123.005 17.450 123.175 ;
        RECT 18.685 123.075 18.855 123.675 ;
        RECT 19.025 123.255 19.375 123.505 ;
        RECT 17.280 122.835 17.910 123.005 ;
        RECT 16.760 122.435 16.990 122.765 ;
        RECT 17.235 122.265 17.565 122.645 ;
        RECT 17.735 122.435 17.910 122.835 ;
        RECT 18.185 122.265 18.425 123.075 ;
        RECT 18.595 122.435 18.925 123.075 ;
        RECT 19.095 122.265 19.365 123.075 ;
        RECT 19.545 122.985 19.805 124.385 ;
        RECT 20.055 124.015 20.385 124.815 ;
        RECT 20.850 123.845 21.100 124.645 ;
        RECT 21.285 124.095 21.615 124.815 ;
        RECT 21.835 123.845 22.085 124.645 ;
        RECT 22.255 124.435 22.590 124.815 ;
        RECT 22.765 124.305 23.955 124.595 ;
        RECT 19.995 123.675 22.185 123.845 ;
        RECT 19.995 123.505 20.310 123.675 ;
        RECT 19.980 123.255 20.310 123.505 ;
        RECT 19.545 122.475 19.885 122.985 ;
        RECT 20.055 122.265 20.325 123.065 ;
        RECT 20.505 122.535 20.785 123.505 ;
        RECT 20.965 122.535 21.265 123.505 ;
        RECT 21.445 122.540 21.795 123.505 ;
        RECT 22.015 122.765 22.185 123.675 ;
        RECT 22.355 122.945 22.595 124.255 ;
        RECT 22.785 123.965 23.955 124.135 ;
        RECT 24.125 124.015 24.405 124.815 ;
        RECT 22.785 123.675 23.110 123.965 ;
        RECT 23.785 123.845 23.955 123.965 ;
        RECT 23.280 123.505 23.475 123.795 ;
        RECT 23.785 123.675 24.445 123.845 ;
        RECT 24.615 123.675 24.890 124.645 ;
        RECT 24.275 123.505 24.445 123.675 ;
        RECT 22.765 123.175 23.110 123.505 ;
        RECT 23.280 123.175 24.105 123.505 ;
        RECT 24.275 123.175 24.550 123.505 ;
        RECT 24.275 123.005 24.445 123.175 ;
        RECT 22.780 122.835 24.445 123.005 ;
        RECT 24.720 122.940 24.890 123.675 ;
        RECT 25.065 123.650 25.355 124.815 ;
        RECT 25.730 123.845 26.060 124.645 ;
        RECT 26.230 124.015 26.560 124.815 ;
        RECT 26.860 123.845 27.190 124.645 ;
        RECT 27.835 124.015 28.085 124.815 ;
        RECT 25.730 123.675 28.165 123.845 ;
        RECT 28.355 123.675 28.525 124.815 ;
        RECT 28.695 123.675 29.035 124.645 ;
        RECT 29.390 123.845 29.780 124.020 ;
        RECT 30.265 124.015 30.595 124.815 ;
        RECT 30.765 124.025 31.300 124.645 ;
        RECT 29.390 123.675 30.815 123.845 ;
        RECT 25.525 123.255 25.875 123.505 ;
        RECT 26.060 123.045 26.230 123.675 ;
        RECT 26.400 123.255 26.730 123.455 ;
        RECT 26.900 123.255 27.230 123.455 ;
        RECT 27.400 123.255 27.820 123.455 ;
        RECT 27.995 123.425 28.165 123.675 ;
        RECT 27.995 123.255 28.690 123.425 ;
        RECT 22.015 122.435 22.510 122.765 ;
        RECT 22.780 122.485 23.035 122.835 ;
        RECT 23.205 122.265 23.535 122.665 ;
        RECT 23.705 122.485 23.875 122.835 ;
        RECT 24.045 122.265 24.425 122.665 ;
        RECT 24.615 122.595 24.890 122.940 ;
        RECT 25.065 122.265 25.355 122.990 ;
        RECT 25.730 122.435 26.230 123.045 ;
        RECT 26.860 122.915 28.085 123.085 ;
        RECT 28.860 123.065 29.035 123.675 ;
        RECT 26.860 122.435 27.190 122.915 ;
        RECT 27.360 122.265 27.585 122.725 ;
        RECT 27.755 122.435 28.085 122.915 ;
        RECT 28.275 122.265 28.525 123.065 ;
        RECT 28.695 122.435 29.035 123.065 ;
        RECT 29.265 122.945 29.620 123.505 ;
        RECT 29.790 122.775 29.960 123.675 ;
        RECT 30.130 122.945 30.395 123.505 ;
        RECT 30.645 123.175 30.815 123.675 ;
        RECT 30.985 123.005 31.300 124.025 ;
        RECT 32.025 123.755 32.355 124.600 ;
        RECT 32.525 123.805 32.695 124.815 ;
        RECT 32.865 124.085 33.205 124.645 ;
        RECT 33.435 124.315 33.750 124.815 ;
        RECT 33.930 124.345 34.815 124.515 ;
        RECT 29.370 122.265 29.610 122.775 ;
        RECT 29.790 122.445 30.070 122.775 ;
        RECT 30.300 122.265 30.515 122.775 ;
        RECT 30.685 122.435 31.300 123.005 ;
        RECT 31.965 123.675 32.355 123.755 ;
        RECT 32.865 123.710 33.760 124.085 ;
        RECT 31.965 123.625 32.180 123.675 ;
        RECT 31.965 123.045 32.135 123.625 ;
        RECT 32.865 123.505 33.055 123.710 ;
        RECT 33.930 123.505 34.100 124.345 ;
        RECT 35.040 124.315 35.290 124.645 ;
        RECT 32.305 123.175 33.055 123.505 ;
        RECT 33.225 123.175 34.100 123.505 ;
        RECT 31.965 123.005 32.190 123.045 ;
        RECT 32.855 123.005 33.055 123.175 ;
        RECT 31.965 122.920 32.345 123.005 ;
        RECT 32.015 122.485 32.345 122.920 ;
        RECT 32.515 122.265 32.685 122.875 ;
        RECT 32.855 122.480 33.185 123.005 ;
        RECT 33.445 122.265 33.655 122.795 ;
        RECT 33.930 122.715 34.100 123.175 ;
        RECT 34.270 123.215 34.590 124.175 ;
        RECT 34.760 123.425 34.950 124.145 ;
        RECT 35.120 123.245 35.290 124.315 ;
        RECT 35.460 124.015 35.630 124.815 ;
        RECT 35.800 124.370 36.905 124.540 ;
        RECT 35.800 123.755 35.970 124.370 ;
        RECT 37.115 124.220 37.365 124.645 ;
        RECT 37.535 124.355 37.800 124.815 ;
        RECT 36.140 123.835 36.670 124.200 ;
        RECT 37.115 124.090 37.420 124.220 ;
        RECT 35.460 123.665 35.970 123.755 ;
        RECT 35.460 123.495 36.330 123.665 ;
        RECT 35.460 123.425 35.630 123.495 ;
        RECT 35.750 123.245 35.950 123.275 ;
        RECT 34.270 122.885 34.735 123.215 ;
        RECT 35.120 122.945 35.950 123.245 ;
        RECT 35.120 122.715 35.290 122.945 ;
        RECT 33.930 122.545 34.715 122.715 ;
        RECT 34.885 122.545 35.290 122.715 ;
        RECT 35.470 122.265 35.840 122.765 ;
        RECT 36.160 122.715 36.330 123.495 ;
        RECT 36.500 123.135 36.670 123.835 ;
        RECT 36.840 123.305 37.080 123.900 ;
        RECT 36.500 122.915 37.025 123.135 ;
        RECT 37.250 122.985 37.420 124.090 ;
        RECT 37.195 122.855 37.420 122.985 ;
        RECT 37.590 122.895 37.870 123.845 ;
        RECT 37.195 122.715 37.365 122.855 ;
        RECT 36.160 122.545 36.835 122.715 ;
        RECT 37.030 122.545 37.365 122.715 ;
        RECT 37.535 122.265 37.785 122.725 ;
        RECT 38.040 122.525 38.225 124.645 ;
        RECT 38.395 124.315 38.725 124.815 ;
        RECT 38.895 124.145 39.065 124.645 ;
        RECT 38.400 123.975 39.065 124.145 ;
        RECT 38.400 122.985 38.630 123.975 ;
        RECT 38.800 123.155 39.150 123.805 ;
        RECT 39.385 123.755 39.715 124.600 ;
        RECT 39.885 123.805 40.055 124.815 ;
        RECT 40.225 124.085 40.565 124.645 ;
        RECT 40.795 124.315 41.110 124.815 ;
        RECT 41.290 124.345 42.175 124.515 ;
        RECT 39.325 123.675 39.715 123.755 ;
        RECT 40.225 123.710 41.120 124.085 ;
        RECT 39.325 123.625 39.540 123.675 ;
        RECT 39.325 123.045 39.495 123.625 ;
        RECT 40.225 123.505 40.415 123.710 ;
        RECT 41.290 123.505 41.460 124.345 ;
        RECT 42.400 124.315 42.650 124.645 ;
        RECT 39.665 123.175 40.415 123.505 ;
        RECT 40.585 123.175 41.460 123.505 ;
        RECT 39.325 123.005 39.550 123.045 ;
        RECT 40.215 123.005 40.415 123.175 ;
        RECT 38.400 122.815 39.065 122.985 ;
        RECT 39.325 122.920 39.705 123.005 ;
        RECT 38.395 122.265 38.725 122.645 ;
        RECT 38.895 122.525 39.065 122.815 ;
        RECT 39.375 122.485 39.705 122.920 ;
        RECT 39.875 122.265 40.045 122.875 ;
        RECT 40.215 122.480 40.545 123.005 ;
        RECT 40.805 122.265 41.015 122.795 ;
        RECT 41.290 122.715 41.460 123.175 ;
        RECT 41.630 123.215 41.950 124.175 ;
        RECT 42.120 123.425 42.310 124.145 ;
        RECT 42.480 123.245 42.650 124.315 ;
        RECT 42.820 124.015 42.990 124.815 ;
        RECT 43.160 124.370 44.265 124.540 ;
        RECT 43.160 123.755 43.330 124.370 ;
        RECT 44.475 124.220 44.725 124.645 ;
        RECT 44.895 124.355 45.160 124.815 ;
        RECT 43.500 123.835 44.030 124.200 ;
        RECT 44.475 124.090 44.780 124.220 ;
        RECT 42.820 123.665 43.330 123.755 ;
        RECT 42.820 123.495 43.690 123.665 ;
        RECT 42.820 123.425 42.990 123.495 ;
        RECT 43.110 123.245 43.310 123.275 ;
        RECT 41.630 122.885 42.095 123.215 ;
        RECT 42.480 122.945 43.310 123.245 ;
        RECT 42.480 122.715 42.650 122.945 ;
        RECT 41.290 122.545 42.075 122.715 ;
        RECT 42.245 122.545 42.650 122.715 ;
        RECT 42.830 122.265 43.200 122.765 ;
        RECT 43.520 122.715 43.690 123.495 ;
        RECT 43.860 123.135 44.030 123.835 ;
        RECT 44.200 123.305 44.440 123.900 ;
        RECT 43.860 122.915 44.385 123.135 ;
        RECT 44.610 122.985 44.780 124.090 ;
        RECT 44.555 122.855 44.780 122.985 ;
        RECT 44.950 122.895 45.230 123.845 ;
        RECT 44.555 122.715 44.725 122.855 ;
        RECT 43.520 122.545 44.195 122.715 ;
        RECT 44.390 122.545 44.725 122.715 ;
        RECT 44.895 122.265 45.145 122.725 ;
        RECT 45.400 122.525 45.585 124.645 ;
        RECT 45.755 124.315 46.085 124.815 ;
        RECT 46.255 124.145 46.425 124.645 ;
        RECT 45.760 123.975 46.425 124.145 ;
        RECT 45.760 122.985 45.990 123.975 ;
        RECT 46.695 123.845 47.025 124.630 ;
        RECT 46.160 123.155 46.510 123.805 ;
        RECT 46.695 123.675 47.375 123.845 ;
        RECT 47.555 123.675 47.885 124.815 ;
        RECT 48.065 123.725 50.655 124.815 ;
        RECT 46.685 123.255 47.035 123.505 ;
        RECT 47.205 123.075 47.375 123.675 ;
        RECT 47.545 123.255 47.895 123.505 ;
        RECT 45.760 122.815 46.425 122.985 ;
        RECT 45.755 122.265 46.085 122.645 ;
        RECT 46.255 122.525 46.425 122.815 ;
        RECT 46.705 122.265 46.945 123.075 ;
        RECT 47.115 122.435 47.445 123.075 ;
        RECT 47.615 122.265 47.885 123.075 ;
        RECT 48.065 123.035 49.275 123.555 ;
        RECT 49.445 123.205 50.655 123.725 ;
        RECT 50.825 123.650 51.115 124.815 ;
        RECT 52.210 123.675 52.545 124.645 ;
        RECT 52.715 123.675 52.885 124.815 ;
        RECT 53.055 124.475 55.085 124.645 ;
        RECT 48.065 122.265 50.655 123.035 ;
        RECT 52.210 123.005 52.380 123.675 ;
        RECT 53.055 123.505 53.225 124.475 ;
        RECT 52.550 123.175 52.805 123.505 ;
        RECT 53.030 123.175 53.225 123.505 ;
        RECT 53.395 124.135 54.520 124.305 ;
        RECT 52.635 123.005 52.805 123.175 ;
        RECT 53.395 123.005 53.565 124.135 ;
        RECT 50.825 122.265 51.115 122.990 ;
        RECT 52.210 122.435 52.465 123.005 ;
        RECT 52.635 122.835 53.565 123.005 ;
        RECT 53.735 123.795 54.745 123.965 ;
        RECT 53.735 122.995 53.905 123.795 ;
        RECT 53.390 122.800 53.565 122.835 ;
        RECT 52.635 122.265 52.965 122.665 ;
        RECT 53.390 122.435 53.920 122.800 ;
        RECT 54.110 122.775 54.385 123.595 ;
        RECT 54.105 122.605 54.385 122.775 ;
        RECT 54.110 122.435 54.385 122.605 ;
        RECT 54.555 122.435 54.745 123.795 ;
        RECT 54.915 123.810 55.085 124.475 ;
        RECT 55.255 124.055 55.425 124.815 ;
        RECT 55.660 124.055 56.175 124.465 ;
        RECT 54.915 123.620 55.665 123.810 ;
        RECT 55.835 123.245 56.175 124.055 ;
        RECT 56.460 124.185 56.745 124.645 ;
        RECT 56.915 124.355 57.185 124.815 ;
        RECT 56.460 123.965 57.415 124.185 ;
        RECT 54.945 123.075 56.175 123.245 ;
        RECT 56.345 123.235 57.035 123.795 ;
        RECT 54.925 122.265 55.435 122.800 ;
        RECT 55.655 122.470 55.900 123.075 ;
        RECT 57.205 123.065 57.415 123.965 ;
        RECT 56.460 122.895 57.415 123.065 ;
        RECT 57.585 123.795 57.985 124.645 ;
        RECT 58.175 124.185 58.455 124.645 ;
        RECT 58.975 124.355 59.300 124.815 ;
        RECT 58.175 123.965 59.300 124.185 ;
        RECT 57.585 123.235 58.680 123.795 ;
        RECT 58.850 123.505 59.300 123.965 ;
        RECT 59.470 123.675 59.855 124.645 ;
        RECT 56.460 122.435 56.745 122.895 ;
        RECT 56.915 122.265 57.185 122.725 ;
        RECT 57.585 122.435 57.985 123.235 ;
        RECT 58.850 123.175 59.405 123.505 ;
        RECT 58.850 123.065 59.300 123.175 ;
        RECT 58.175 122.895 59.300 123.065 ;
        RECT 59.575 123.005 59.855 123.675 ;
        RECT 58.175 122.435 58.455 122.895 ;
        RECT 58.975 122.265 59.300 122.725 ;
        RECT 59.470 122.435 59.855 123.005 ;
        RECT 60.025 122.545 60.305 124.645 ;
        RECT 60.495 124.055 61.280 124.815 ;
        RECT 61.675 123.985 62.060 124.645 ;
        RECT 61.675 123.885 62.085 123.985 ;
        RECT 60.475 123.675 62.085 123.885 ;
        RECT 62.385 123.795 62.585 124.585 ;
        RECT 60.475 123.075 60.750 123.675 ;
        RECT 62.255 123.625 62.585 123.795 ;
        RECT 62.755 123.635 63.075 124.815 ;
        RECT 63.250 123.675 63.570 124.815 ;
        RECT 62.255 123.505 62.435 123.625 ;
        RECT 63.750 123.505 63.945 124.555 ;
        RECT 64.125 123.965 64.455 124.645 ;
        RECT 64.655 124.015 64.910 124.815 ;
        RECT 65.090 124.015 65.345 124.815 ;
        RECT 65.545 123.965 65.875 124.645 ;
        RECT 64.125 123.685 64.475 123.965 ;
        RECT 60.920 123.255 61.275 123.505 ;
        RECT 61.470 123.455 61.935 123.505 ;
        RECT 61.465 123.285 61.935 123.455 ;
        RECT 61.470 123.255 61.935 123.285 ;
        RECT 62.105 123.255 62.435 123.505 ;
        RECT 63.310 123.455 63.570 123.505 ;
        RECT 62.610 123.255 63.075 123.455 ;
        RECT 63.305 123.285 63.570 123.455 ;
        RECT 63.310 123.175 63.570 123.285 ;
        RECT 63.750 123.175 64.135 123.505 ;
        RECT 64.305 123.305 64.475 123.685 ;
        RECT 64.665 123.475 64.910 123.835 ;
        RECT 65.090 123.475 65.335 123.835 ;
        RECT 65.525 123.685 65.875 123.965 ;
        RECT 65.525 123.305 65.695 123.685 ;
        RECT 66.055 123.505 66.250 124.555 ;
        RECT 66.430 123.675 66.750 124.815 ;
        RECT 66.925 123.965 67.185 124.645 ;
        RECT 67.355 124.035 67.605 124.815 ;
        RECT 67.855 124.265 68.105 124.645 ;
        RECT 68.275 124.435 68.630 124.815 ;
        RECT 69.635 124.425 69.970 124.645 ;
        RECT 69.235 124.265 69.465 124.305 ;
        RECT 67.855 124.065 69.465 124.265 ;
        RECT 67.855 124.055 68.690 124.065 ;
        RECT 69.280 123.975 69.465 124.065 ;
        RECT 64.305 123.135 64.825 123.305 ;
        RECT 60.475 122.895 61.725 123.075 ;
        RECT 61.360 122.825 61.725 122.895 ;
        RECT 61.895 122.875 63.075 123.045 ;
        RECT 60.535 122.265 60.705 122.725 ;
        RECT 61.895 122.655 62.225 122.875 ;
        RECT 60.975 122.475 62.225 122.655 ;
        RECT 62.395 122.265 62.565 122.705 ;
        RECT 62.735 122.460 63.075 122.875 ;
        RECT 63.250 122.795 64.465 122.965 ;
        RECT 63.250 122.445 63.540 122.795 ;
        RECT 63.735 122.265 64.065 122.625 ;
        RECT 64.235 122.490 64.465 122.795 ;
        RECT 64.655 122.570 64.825 123.135 ;
        RECT 65.175 123.135 65.695 123.305 ;
        RECT 65.865 123.175 66.250 123.505 ;
        RECT 66.430 123.455 66.690 123.505 ;
        RECT 66.430 123.285 66.695 123.455 ;
        RECT 66.430 123.175 66.690 123.285 ;
        RECT 65.175 122.570 65.345 123.135 ;
        RECT 65.535 122.795 66.750 122.965 ;
        RECT 65.535 122.490 65.765 122.795 ;
        RECT 65.935 122.265 66.265 122.625 ;
        RECT 66.460 122.445 66.750 122.795 ;
        RECT 66.925 122.775 67.095 123.965 ;
        RECT 68.795 123.865 69.125 123.895 ;
        RECT 67.325 123.805 69.125 123.865 ;
        RECT 69.715 123.805 69.970 124.425 ;
        RECT 70.260 124.185 70.545 124.645 ;
        RECT 70.715 124.355 70.985 124.815 ;
        RECT 70.260 123.965 71.215 124.185 ;
        RECT 67.265 123.695 69.970 123.805 ;
        RECT 67.265 123.660 67.465 123.695 ;
        RECT 67.265 123.085 67.435 123.660 ;
        RECT 68.795 123.635 69.970 123.695 ;
        RECT 67.665 123.220 68.075 123.525 ;
        RECT 68.245 123.255 68.575 123.465 ;
        RECT 67.265 122.965 67.535 123.085 ;
        RECT 67.265 122.920 68.110 122.965 ;
        RECT 67.355 122.795 68.110 122.920 ;
        RECT 68.365 122.855 68.575 123.255 ;
        RECT 68.820 123.255 69.295 123.465 ;
        RECT 69.485 123.255 69.975 123.455 ;
        RECT 68.820 122.855 69.040 123.255 ;
        RECT 70.145 123.235 70.835 123.795 ;
        RECT 71.005 123.065 71.215 123.965 ;
        RECT 66.925 122.765 67.155 122.775 ;
        RECT 66.925 122.435 67.185 122.765 ;
        RECT 67.940 122.645 68.110 122.795 ;
        RECT 67.355 122.265 67.685 122.625 ;
        RECT 67.940 122.435 69.240 122.645 ;
        RECT 69.515 122.265 69.970 123.030 ;
        RECT 70.260 122.895 71.215 123.065 ;
        RECT 71.385 123.795 71.785 124.645 ;
        RECT 71.975 124.185 72.255 124.645 ;
        RECT 72.775 124.355 73.100 124.815 ;
        RECT 71.975 123.965 73.100 124.185 ;
        RECT 71.385 123.235 72.480 123.795 ;
        RECT 72.650 123.505 73.100 123.965 ;
        RECT 73.270 123.675 73.655 124.645 ;
        RECT 73.835 123.675 74.165 124.815 ;
        RECT 70.260 122.435 70.545 122.895 ;
        RECT 70.715 122.265 70.985 122.725 ;
        RECT 71.385 122.435 71.785 123.235 ;
        RECT 72.650 123.175 73.205 123.505 ;
        RECT 72.650 123.065 73.100 123.175 ;
        RECT 71.975 122.895 73.100 123.065 ;
        RECT 73.375 123.005 73.655 123.675 ;
        RECT 71.975 122.435 72.255 122.895 ;
        RECT 72.775 122.265 73.100 122.725 ;
        RECT 73.270 122.435 73.655 123.005 ;
        RECT 73.825 122.925 74.165 123.505 ;
        RECT 74.335 123.475 74.695 124.645 ;
        RECT 74.895 123.645 75.225 124.815 ;
        RECT 75.425 123.475 75.755 124.645 ;
        RECT 75.955 123.645 76.285 124.815 ;
        RECT 76.585 123.650 76.875 124.815 ;
        RECT 77.250 123.845 77.580 124.645 ;
        RECT 77.750 124.015 78.080 124.815 ;
        RECT 78.380 123.845 78.710 124.645 ;
        RECT 79.355 124.015 79.605 124.815 ;
        RECT 77.250 123.675 79.685 123.845 ;
        RECT 79.875 123.675 80.045 124.815 ;
        RECT 80.215 123.675 80.555 124.645 ;
        RECT 80.815 124.145 80.985 124.645 ;
        RECT 81.155 124.315 81.485 124.815 ;
        RECT 80.815 123.975 81.480 124.145 ;
        RECT 74.335 123.195 75.755 123.475 ;
        RECT 77.045 123.255 77.395 123.505 ;
        RECT 74.335 122.860 74.695 123.195 ;
        RECT 77.580 123.045 77.750 123.675 ;
        RECT 77.920 123.255 78.250 123.455 ;
        RECT 78.420 123.255 78.750 123.455 ;
        RECT 78.920 123.255 79.340 123.455 ;
        RECT 79.515 123.425 79.685 123.675 ;
        RECT 79.515 123.255 80.210 123.425 ;
        RECT 80.380 123.115 80.555 123.675 ;
        RECT 80.730 123.155 81.080 123.805 ;
        RECT 73.835 122.265 74.165 122.755 ;
        RECT 74.335 122.435 74.955 122.860 ;
        RECT 75.415 122.265 75.745 122.955 ;
        RECT 76.585 122.265 76.875 122.990 ;
        RECT 77.250 122.435 77.750 123.045 ;
        RECT 78.380 122.915 79.605 123.085 ;
        RECT 80.325 123.065 80.555 123.115 ;
        RECT 78.380 122.435 78.710 122.915 ;
        RECT 78.880 122.265 79.105 122.725 ;
        RECT 79.275 122.435 79.605 122.915 ;
        RECT 79.795 122.265 80.045 123.065 ;
        RECT 80.215 122.435 80.555 123.065 ;
        RECT 81.250 122.985 81.480 123.975 ;
        RECT 80.815 122.815 81.480 122.985 ;
        RECT 80.815 122.525 80.985 122.815 ;
        RECT 81.155 122.265 81.485 122.645 ;
        RECT 81.655 122.525 81.840 124.645 ;
        RECT 82.080 124.355 82.345 124.815 ;
        RECT 82.515 124.220 82.765 124.645 ;
        RECT 82.975 124.370 84.080 124.540 ;
        RECT 82.460 124.090 82.765 124.220 ;
        RECT 82.010 122.895 82.290 123.845 ;
        RECT 82.460 122.985 82.630 124.090 ;
        RECT 82.800 123.305 83.040 123.900 ;
        RECT 83.210 123.835 83.740 124.200 ;
        RECT 83.210 123.135 83.380 123.835 ;
        RECT 83.910 123.755 84.080 124.370 ;
        RECT 84.250 124.015 84.420 124.815 ;
        RECT 84.590 124.315 84.840 124.645 ;
        RECT 85.065 124.345 85.950 124.515 ;
        RECT 83.910 123.665 84.420 123.755 ;
        RECT 82.460 122.855 82.685 122.985 ;
        RECT 82.855 122.915 83.380 123.135 ;
        RECT 83.550 123.495 84.420 123.665 ;
        RECT 82.095 122.265 82.345 122.725 ;
        RECT 82.515 122.715 82.685 122.855 ;
        RECT 83.550 122.715 83.720 123.495 ;
        RECT 84.250 123.425 84.420 123.495 ;
        RECT 83.930 123.245 84.130 123.275 ;
        RECT 84.590 123.245 84.760 124.315 ;
        RECT 84.930 123.425 85.120 124.145 ;
        RECT 83.930 122.945 84.760 123.245 ;
        RECT 85.290 123.215 85.610 124.175 ;
        RECT 82.515 122.545 82.850 122.715 ;
        RECT 83.045 122.545 83.720 122.715 ;
        RECT 84.040 122.265 84.410 122.765 ;
        RECT 84.590 122.715 84.760 122.945 ;
        RECT 85.145 122.885 85.610 123.215 ;
        RECT 85.780 123.505 85.950 124.345 ;
        RECT 86.130 124.315 86.445 124.815 ;
        RECT 86.675 124.085 87.015 124.645 ;
        RECT 86.120 123.710 87.015 124.085 ;
        RECT 87.185 123.805 87.355 124.815 ;
        RECT 86.825 123.505 87.015 123.710 ;
        RECT 87.525 123.755 87.855 124.600 ;
        RECT 87.525 123.675 87.915 123.755 ;
        RECT 87.700 123.625 87.915 123.675 ;
        RECT 85.780 123.175 86.655 123.505 ;
        RECT 86.825 123.175 87.575 123.505 ;
        RECT 85.780 122.715 85.950 123.175 ;
        RECT 86.825 123.005 87.025 123.175 ;
        RECT 87.745 123.045 87.915 123.625 ;
        RECT 88.545 123.725 89.755 124.815 ;
        RECT 88.545 123.185 89.065 123.725 ;
        RECT 87.690 123.005 87.915 123.045 ;
        RECT 89.235 123.015 89.755 123.555 ;
        RECT 84.590 122.545 84.995 122.715 ;
        RECT 85.165 122.545 85.950 122.715 ;
        RECT 86.225 122.265 86.435 122.795 ;
        RECT 86.695 122.480 87.025 123.005 ;
        RECT 87.535 122.920 87.915 123.005 ;
        RECT 87.195 122.265 87.365 122.875 ;
        RECT 87.535 122.485 87.865 122.920 ;
        RECT 88.545 122.265 89.755 123.015 ;
        RECT 100.140 122.460 100.810 125.720 ;
        RECT 101.480 125.150 105.520 125.320 ;
        RECT 101.140 123.090 101.310 125.090 ;
        RECT 105.690 123.090 105.860 125.090 ;
        RECT 101.480 122.860 105.520 123.030 ;
        RECT 106.200 122.460 106.370 125.720 ;
        RECT 100.140 122.450 106.370 122.460 ;
        RECT 107.960 131.720 117.790 131.760 ;
        RECT 107.960 131.590 118.590 131.720 ;
        RECT 107.960 129.330 108.130 131.590 ;
        RECT 108.855 131.020 116.895 131.190 ;
        RECT 108.470 129.960 108.640 130.960 ;
        RECT 117.110 129.960 117.280 130.960 ;
        RECT 108.855 129.730 116.895 129.900 ;
        RECT 117.620 129.330 118.590 131.590 ;
        RECT 107.960 129.160 118.590 129.330 ;
        RECT 107.960 125.900 108.130 129.160 ;
        RECT 108.855 128.590 116.895 128.760 ;
        RECT 108.470 126.530 108.640 128.530 ;
        RECT 117.110 126.530 117.280 128.530 ;
        RECT 108.855 126.300 116.895 126.470 ;
        RECT 117.620 125.900 118.590 129.160 ;
        RECT 107.960 125.730 118.590 125.900 ;
        RECT 107.960 122.470 108.130 125.730 ;
        RECT 108.855 125.160 116.895 125.330 ;
        RECT 108.470 123.100 108.640 125.100 ;
        RECT 117.110 123.100 117.280 125.100 ;
        RECT 108.855 122.870 116.895 123.040 ;
        RECT 117.620 122.470 118.590 125.730 ;
        RECT 100.140 122.350 106.380 122.450 ;
        RECT 12.100 122.095 89.840 122.265 ;
        RECT 12.185 121.345 13.395 122.095 ;
        RECT 12.185 120.805 12.705 121.345 ;
        RECT 13.565 121.325 16.155 122.095 ;
        RECT 16.335 121.365 16.635 122.095 ;
        RECT 12.875 120.635 13.395 121.175 ;
        RECT 13.565 120.805 14.775 121.325 ;
        RECT 16.815 121.185 17.045 121.805 ;
        RECT 17.245 121.535 17.470 121.915 ;
        RECT 17.640 121.705 17.970 122.095 ;
        RECT 18.165 121.715 19.055 121.885 ;
        RECT 17.245 121.355 17.575 121.535 ;
        RECT 14.945 120.635 16.155 121.155 ;
        RECT 16.340 120.855 16.635 121.185 ;
        RECT 16.815 120.855 17.230 121.185 ;
        RECT 17.400 120.685 17.575 121.355 ;
        RECT 17.745 120.855 17.985 121.505 ;
        RECT 18.165 121.160 18.715 121.545 ;
        RECT 18.885 120.990 19.055 121.715 ;
        RECT 18.165 120.920 19.055 120.990 ;
        RECT 19.225 121.390 19.445 121.875 ;
        RECT 19.615 121.555 19.865 122.095 ;
        RECT 20.035 121.445 20.295 121.925 ;
        RECT 19.225 120.965 19.555 121.390 ;
        RECT 18.165 120.895 19.060 120.920 ;
        RECT 18.165 120.880 19.070 120.895 ;
        RECT 18.165 120.865 19.075 120.880 ;
        RECT 18.165 120.860 19.085 120.865 ;
        RECT 18.165 120.850 19.090 120.860 ;
        RECT 18.165 120.840 19.095 120.850 ;
        RECT 18.165 120.835 19.105 120.840 ;
        RECT 18.165 120.825 19.115 120.835 ;
        RECT 18.165 120.820 19.125 120.825 ;
        RECT 12.185 119.545 13.395 120.635 ;
        RECT 13.565 119.545 16.155 120.635 ;
        RECT 16.335 120.325 17.230 120.655 ;
        RECT 17.400 120.495 17.985 120.685 ;
        RECT 16.335 120.155 17.540 120.325 ;
        RECT 16.335 119.725 16.665 120.155 ;
        RECT 16.845 119.545 17.040 119.985 ;
        RECT 17.210 119.725 17.540 120.155 ;
        RECT 17.710 119.725 17.985 120.495 ;
        RECT 18.165 120.370 18.425 120.820 ;
        RECT 18.790 120.815 19.125 120.820 ;
        RECT 18.790 120.810 19.140 120.815 ;
        RECT 18.790 120.800 19.155 120.810 ;
        RECT 18.790 120.795 19.180 120.800 ;
        RECT 19.725 120.795 19.955 121.190 ;
        RECT 18.790 120.790 19.955 120.795 ;
        RECT 18.820 120.755 19.955 120.790 ;
        RECT 18.855 120.730 19.955 120.755 ;
        RECT 18.885 120.700 19.955 120.730 ;
        RECT 18.905 120.670 19.955 120.700 ;
        RECT 18.925 120.640 19.955 120.670 ;
        RECT 18.995 120.630 19.955 120.640 ;
        RECT 19.020 120.620 19.955 120.630 ;
        RECT 19.040 120.605 19.955 120.620 ;
        RECT 19.060 120.590 19.955 120.605 ;
        RECT 19.065 120.580 19.850 120.590 ;
        RECT 19.080 120.545 19.850 120.580 ;
        RECT 18.595 120.225 18.925 120.470 ;
        RECT 19.095 120.295 19.850 120.545 ;
        RECT 20.125 120.415 20.295 121.445 ;
        RECT 18.595 120.200 18.780 120.225 ;
        RECT 18.165 120.100 18.780 120.200 ;
        RECT 18.165 119.545 18.770 120.100 ;
        RECT 18.945 119.715 19.425 120.055 ;
        RECT 19.595 119.545 19.850 120.090 ;
        RECT 20.020 119.715 20.295 120.415 ;
        RECT 20.925 121.355 21.390 121.900 ;
        RECT 20.925 120.395 21.095 121.355 ;
        RECT 21.895 121.275 22.065 122.095 ;
        RECT 22.235 121.445 22.565 121.925 ;
        RECT 22.735 121.705 23.085 122.095 ;
        RECT 23.255 121.525 23.485 121.925 ;
        RECT 22.975 121.445 23.485 121.525 ;
        RECT 22.235 121.355 23.485 121.445 ;
        RECT 23.655 121.355 23.975 121.835 ;
        RECT 22.235 121.275 23.145 121.355 ;
        RECT 21.265 120.735 21.510 121.185 ;
        RECT 21.770 120.905 22.465 121.105 ;
        RECT 22.635 120.935 23.235 121.105 ;
        RECT 22.635 120.735 22.805 120.935 ;
        RECT 23.465 120.765 23.635 121.185 ;
        RECT 21.265 120.565 22.805 120.735 ;
        RECT 22.975 120.595 23.635 120.765 ;
        RECT 22.975 120.395 23.145 120.595 ;
        RECT 23.805 120.425 23.975 121.355 ;
        RECT 24.145 121.325 25.815 122.095 ;
        RECT 24.145 120.805 24.895 121.325 ;
        RECT 25.985 121.275 26.245 122.095 ;
        RECT 26.415 121.275 26.745 121.695 ;
        RECT 26.925 121.525 27.185 121.925 ;
        RECT 27.355 121.695 27.685 122.095 ;
        RECT 27.855 121.525 28.025 121.875 ;
        RECT 28.195 121.695 28.570 122.095 ;
        RECT 26.925 121.355 28.590 121.525 ;
        RECT 28.760 121.420 29.035 121.765 ;
        RECT 26.495 121.185 26.745 121.275 ;
        RECT 28.420 121.185 28.590 121.355 ;
        RECT 25.065 120.635 25.815 121.155 ;
        RECT 25.990 120.855 26.325 121.105 ;
        RECT 26.495 120.855 27.210 121.185 ;
        RECT 27.425 120.855 28.250 121.185 ;
        RECT 28.420 120.855 28.695 121.185 ;
        RECT 20.925 120.225 23.145 120.395 ;
        RECT 23.315 120.225 23.975 120.425 ;
        RECT 20.925 119.545 21.225 120.055 ;
        RECT 21.395 119.715 21.725 120.225 ;
        RECT 23.315 120.055 23.485 120.225 ;
        RECT 21.895 119.545 22.525 120.055 ;
        RECT 23.105 119.885 23.485 120.055 ;
        RECT 23.655 119.545 23.955 120.055 ;
        RECT 24.145 119.545 25.815 120.635 ;
        RECT 25.985 119.545 26.245 120.685 ;
        RECT 26.495 120.295 26.665 120.855 ;
        RECT 26.925 120.395 27.255 120.685 ;
        RECT 27.425 120.565 27.670 120.855 ;
        RECT 28.420 120.685 28.590 120.855 ;
        RECT 28.865 120.685 29.035 121.420 ;
        RECT 29.220 121.525 29.475 121.875 ;
        RECT 29.645 121.695 29.975 122.095 ;
        RECT 30.145 121.525 30.315 121.875 ;
        RECT 30.485 121.695 30.865 122.095 ;
        RECT 29.220 121.355 30.885 121.525 ;
        RECT 31.055 121.420 31.330 121.765 ;
        RECT 31.555 121.705 31.885 122.095 ;
        RECT 32.055 121.525 32.225 121.845 ;
        RECT 32.395 121.705 32.725 122.095 ;
        RECT 33.140 121.695 34.095 121.865 ;
        RECT 30.715 121.185 30.885 121.355 ;
        RECT 29.205 120.855 29.550 121.185 ;
        RECT 29.720 120.855 30.545 121.185 ;
        RECT 30.715 120.855 30.990 121.185 ;
        RECT 27.930 120.515 28.590 120.685 ;
        RECT 27.930 120.395 28.100 120.515 ;
        RECT 26.925 120.225 28.100 120.395 ;
        RECT 26.485 119.725 28.100 120.055 ;
        RECT 28.270 119.545 28.550 120.345 ;
        RECT 28.760 119.715 29.035 120.685 ;
        RECT 29.225 120.395 29.550 120.685 ;
        RECT 29.720 120.565 29.915 120.855 ;
        RECT 30.715 120.685 30.885 120.855 ;
        RECT 31.160 120.685 31.330 121.420 ;
        RECT 30.225 120.515 30.885 120.685 ;
        RECT 30.225 120.395 30.395 120.515 ;
        RECT 29.225 120.225 30.395 120.395 ;
        RECT 29.205 119.765 30.395 120.055 ;
        RECT 30.565 119.545 30.845 120.345 ;
        RECT 31.055 119.715 31.330 120.685 ;
        RECT 31.505 121.355 33.755 121.525 ;
        RECT 31.505 120.395 31.675 121.355 ;
        RECT 31.845 120.735 32.090 121.185 ;
        RECT 32.260 120.905 32.810 121.105 ;
        RECT 32.980 120.935 33.355 121.105 ;
        RECT 32.980 120.735 33.150 120.935 ;
        RECT 33.525 120.855 33.755 121.355 ;
        RECT 31.845 120.565 33.150 120.735 ;
        RECT 33.925 120.815 34.095 121.695 ;
        RECT 34.265 121.260 34.555 122.095 ;
        RECT 34.735 121.370 35.065 121.880 ;
        RECT 35.235 121.695 35.565 122.095 ;
        RECT 36.615 121.525 36.945 121.865 ;
        RECT 37.115 121.695 37.445 122.095 ;
        RECT 33.925 120.645 34.555 120.815 ;
        RECT 31.505 119.715 31.885 120.395 ;
        RECT 32.475 119.545 32.645 120.395 ;
        RECT 32.815 120.225 34.055 120.395 ;
        RECT 32.815 119.715 33.145 120.225 ;
        RECT 33.315 119.545 33.485 120.055 ;
        RECT 33.655 119.715 34.055 120.225 ;
        RECT 34.235 119.715 34.555 120.645 ;
        RECT 34.735 120.605 34.925 121.370 ;
        RECT 35.235 121.355 37.600 121.525 ;
        RECT 37.945 121.370 38.235 122.095 ;
        RECT 38.410 121.695 38.745 122.095 ;
        RECT 38.915 121.525 39.120 121.925 ;
        RECT 39.330 121.615 39.605 122.095 ;
        RECT 39.815 121.595 40.075 121.925 ;
        RECT 35.235 121.185 35.405 121.355 ;
        RECT 35.095 120.855 35.405 121.185 ;
        RECT 35.575 120.855 35.880 121.185 ;
        RECT 34.735 119.755 35.065 120.605 ;
        RECT 35.235 119.545 35.485 120.685 ;
        RECT 35.665 120.525 35.880 120.855 ;
        RECT 36.055 120.525 36.340 121.185 ;
        RECT 36.535 120.525 36.800 121.185 ;
        RECT 37.015 120.525 37.260 121.185 ;
        RECT 37.430 120.355 37.600 121.355 ;
        RECT 38.435 121.355 39.120 121.525 ;
        RECT 35.675 120.185 36.965 120.355 ;
        RECT 35.675 119.765 35.925 120.185 ;
        RECT 36.155 119.545 36.485 120.015 ;
        RECT 36.715 119.765 36.965 120.185 ;
        RECT 37.145 120.185 37.600 120.355 ;
        RECT 37.145 119.755 37.475 120.185 ;
        RECT 37.945 119.545 38.235 120.710 ;
        RECT 38.435 120.325 38.775 121.355 ;
        RECT 38.945 120.685 39.195 121.185 ;
        RECT 39.375 120.855 39.735 121.435 ;
        RECT 39.905 120.685 40.075 121.595 ;
        RECT 41.255 121.545 41.425 121.835 ;
        RECT 41.595 121.715 41.925 122.095 ;
        RECT 41.255 121.375 41.920 121.545 ;
        RECT 38.945 120.515 40.075 120.685 ;
        RECT 41.170 120.555 41.520 121.205 ;
        RECT 38.435 120.150 39.100 120.325 ;
        RECT 38.410 119.545 38.745 119.970 ;
        RECT 38.915 119.745 39.100 120.150 ;
        RECT 39.305 119.545 39.635 120.325 ;
        RECT 39.805 119.745 40.075 120.515 ;
        RECT 41.690 120.385 41.920 121.375 ;
        RECT 41.255 120.215 41.920 120.385 ;
        RECT 41.255 119.715 41.425 120.215 ;
        RECT 41.595 119.545 41.925 120.045 ;
        RECT 42.095 119.715 42.280 121.835 ;
        RECT 42.535 121.635 42.785 122.095 ;
        RECT 42.955 121.645 43.290 121.815 ;
        RECT 43.485 121.645 44.160 121.815 ;
        RECT 42.955 121.505 43.125 121.645 ;
        RECT 42.450 120.515 42.730 121.465 ;
        RECT 42.900 121.375 43.125 121.505 ;
        RECT 42.900 120.270 43.070 121.375 ;
        RECT 43.295 121.225 43.820 121.445 ;
        RECT 43.240 120.460 43.480 121.055 ;
        RECT 43.650 120.525 43.820 121.225 ;
        RECT 43.990 120.865 44.160 121.645 ;
        RECT 44.480 121.595 44.850 122.095 ;
        RECT 45.030 121.645 45.435 121.815 ;
        RECT 45.605 121.645 46.390 121.815 ;
        RECT 45.030 121.415 45.200 121.645 ;
        RECT 44.370 121.115 45.200 121.415 ;
        RECT 45.585 121.145 46.050 121.475 ;
        RECT 44.370 121.085 44.570 121.115 ;
        RECT 44.690 120.865 44.860 120.935 ;
        RECT 43.990 120.695 44.860 120.865 ;
        RECT 44.350 120.605 44.860 120.695 ;
        RECT 42.900 120.140 43.205 120.270 ;
        RECT 43.650 120.160 44.180 120.525 ;
        RECT 42.520 119.545 42.785 120.005 ;
        RECT 42.955 119.715 43.205 120.140 ;
        RECT 44.350 119.990 44.520 120.605 ;
        RECT 43.415 119.820 44.520 119.990 ;
        RECT 44.690 119.545 44.860 120.345 ;
        RECT 45.030 120.045 45.200 121.115 ;
        RECT 45.370 120.215 45.560 120.935 ;
        RECT 45.730 120.185 46.050 121.145 ;
        RECT 46.220 121.185 46.390 121.645 ;
        RECT 46.665 121.565 46.875 122.095 ;
        RECT 47.135 121.355 47.465 121.880 ;
        RECT 47.635 121.485 47.805 122.095 ;
        RECT 47.975 121.440 48.305 121.875 ;
        RECT 48.615 121.545 48.785 121.835 ;
        RECT 48.955 121.715 49.285 122.095 ;
        RECT 47.975 121.355 48.355 121.440 ;
        RECT 48.615 121.375 49.280 121.545 ;
        RECT 47.265 121.185 47.465 121.355 ;
        RECT 48.130 121.315 48.355 121.355 ;
        RECT 46.220 120.855 47.095 121.185 ;
        RECT 47.265 120.855 48.015 121.185 ;
        RECT 45.030 119.715 45.280 120.045 ;
        RECT 46.220 120.015 46.390 120.855 ;
        RECT 47.265 120.650 47.455 120.855 ;
        RECT 48.185 120.735 48.355 121.315 ;
        RECT 48.140 120.685 48.355 120.735 ;
        RECT 46.560 120.275 47.455 120.650 ;
        RECT 47.965 120.605 48.355 120.685 ;
        RECT 45.505 119.845 46.390 120.015 ;
        RECT 46.570 119.545 46.885 120.045 ;
        RECT 47.115 119.715 47.455 120.275 ;
        RECT 47.625 119.545 47.795 120.555 ;
        RECT 47.965 119.760 48.295 120.605 ;
        RECT 48.530 120.555 48.880 121.205 ;
        RECT 49.050 120.385 49.280 121.375 ;
        RECT 48.615 120.215 49.280 120.385 ;
        RECT 48.615 119.715 48.785 120.215 ;
        RECT 48.955 119.545 49.285 120.045 ;
        RECT 49.455 119.715 49.640 121.835 ;
        RECT 49.895 121.635 50.145 122.095 ;
        RECT 50.315 121.645 50.650 121.815 ;
        RECT 50.845 121.645 51.520 121.815 ;
        RECT 50.315 121.505 50.485 121.645 ;
        RECT 49.810 120.515 50.090 121.465 ;
        RECT 50.260 121.375 50.485 121.505 ;
        RECT 50.260 120.270 50.430 121.375 ;
        RECT 50.655 121.225 51.180 121.445 ;
        RECT 50.600 120.460 50.840 121.055 ;
        RECT 51.010 120.525 51.180 121.225 ;
        RECT 51.350 120.865 51.520 121.645 ;
        RECT 51.840 121.595 52.210 122.095 ;
        RECT 52.390 121.645 52.795 121.815 ;
        RECT 52.965 121.645 53.750 121.815 ;
        RECT 52.390 121.415 52.560 121.645 ;
        RECT 51.730 121.115 52.560 121.415 ;
        RECT 52.945 121.145 53.410 121.475 ;
        RECT 51.730 121.085 51.930 121.115 ;
        RECT 52.050 120.865 52.220 120.935 ;
        RECT 51.350 120.695 52.220 120.865 ;
        RECT 51.710 120.605 52.220 120.695 ;
        RECT 50.260 120.140 50.565 120.270 ;
        RECT 51.010 120.160 51.540 120.525 ;
        RECT 49.880 119.545 50.145 120.005 ;
        RECT 50.315 119.715 50.565 120.140 ;
        RECT 51.710 119.990 51.880 120.605 ;
        RECT 50.775 119.820 51.880 119.990 ;
        RECT 52.050 119.545 52.220 120.345 ;
        RECT 52.390 120.045 52.560 121.115 ;
        RECT 52.730 120.215 52.920 120.935 ;
        RECT 53.090 120.185 53.410 121.145 ;
        RECT 53.580 121.185 53.750 121.645 ;
        RECT 54.025 121.565 54.235 122.095 ;
        RECT 54.495 121.355 54.825 121.880 ;
        RECT 54.995 121.485 55.165 122.095 ;
        RECT 55.335 121.440 55.665 121.875 ;
        RECT 55.335 121.355 55.715 121.440 ;
        RECT 54.625 121.185 54.825 121.355 ;
        RECT 55.490 121.315 55.715 121.355 ;
        RECT 53.580 120.855 54.455 121.185 ;
        RECT 54.625 120.855 55.375 121.185 ;
        RECT 52.390 119.715 52.640 120.045 ;
        RECT 53.580 120.015 53.750 120.855 ;
        RECT 54.625 120.650 54.815 120.855 ;
        RECT 55.545 120.735 55.715 121.315 ;
        RECT 55.500 120.685 55.715 120.735 ;
        RECT 53.920 120.275 54.815 120.650 ;
        RECT 55.325 120.605 55.715 120.685 ;
        RECT 55.885 121.355 56.270 121.925 ;
        RECT 56.440 121.635 56.765 122.095 ;
        RECT 57.285 121.465 57.565 121.925 ;
        RECT 55.885 120.685 56.165 121.355 ;
        RECT 56.440 121.295 57.565 121.465 ;
        RECT 56.440 121.185 56.890 121.295 ;
        RECT 56.335 120.855 56.890 121.185 ;
        RECT 57.755 121.125 58.155 121.925 ;
        RECT 58.555 121.635 58.825 122.095 ;
        RECT 58.995 121.465 59.280 121.925 ;
        RECT 52.865 119.845 53.750 120.015 ;
        RECT 53.930 119.545 54.245 120.045 ;
        RECT 54.475 119.715 54.815 120.275 ;
        RECT 54.985 119.545 55.155 120.555 ;
        RECT 55.325 119.760 55.655 120.605 ;
        RECT 55.885 119.715 56.270 120.685 ;
        RECT 56.440 120.395 56.890 120.855 ;
        RECT 57.060 120.565 58.155 121.125 ;
        RECT 56.440 120.175 57.565 120.395 ;
        RECT 56.440 119.545 56.765 120.005 ;
        RECT 57.285 119.715 57.565 120.175 ;
        RECT 57.755 119.715 58.155 120.565 ;
        RECT 58.325 121.295 59.280 121.465 ;
        RECT 59.570 121.330 60.025 122.095 ;
        RECT 60.300 121.715 61.600 121.925 ;
        RECT 61.855 121.735 62.185 122.095 ;
        RECT 61.430 121.565 61.600 121.715 ;
        RECT 62.355 121.595 62.615 121.925 ;
        RECT 62.385 121.585 62.615 121.595 ;
        RECT 58.325 120.395 58.535 121.295 ;
        RECT 58.705 120.565 59.395 121.125 ;
        RECT 60.500 121.105 60.720 121.505 ;
        RECT 59.565 120.905 60.055 121.105 ;
        RECT 60.245 120.895 60.720 121.105 ;
        RECT 60.965 121.105 61.175 121.505 ;
        RECT 61.430 121.440 62.185 121.565 ;
        RECT 61.430 121.395 62.275 121.440 ;
        RECT 62.005 121.275 62.275 121.395 ;
        RECT 60.965 120.895 61.295 121.105 ;
        RECT 61.465 120.835 61.875 121.140 ;
        RECT 59.570 120.665 60.745 120.725 ;
        RECT 62.105 120.700 62.275 121.275 ;
        RECT 62.075 120.665 62.275 120.700 ;
        RECT 59.570 120.555 62.275 120.665 ;
        RECT 58.325 120.175 59.280 120.395 ;
        RECT 58.555 119.545 58.825 120.005 ;
        RECT 58.995 119.715 59.280 120.175 ;
        RECT 59.570 119.935 59.825 120.555 ;
        RECT 60.415 120.495 62.215 120.555 ;
        RECT 60.415 120.465 60.745 120.495 ;
        RECT 62.445 120.395 62.615 121.585 ;
        RECT 63.705 121.370 63.995 122.095 ;
        RECT 64.210 121.635 64.475 122.095 ;
        RECT 64.845 121.455 65.015 121.925 ;
        RECT 65.265 121.635 65.435 122.095 ;
        RECT 65.685 121.455 65.855 121.925 ;
        RECT 66.105 121.635 66.275 122.095 ;
        RECT 66.525 121.455 66.695 121.925 ;
        RECT 66.865 121.630 67.115 122.095 ;
        RECT 64.845 121.275 67.215 121.455 ;
        RECT 67.435 121.440 67.765 121.875 ;
        RECT 67.935 121.485 68.105 122.095 ;
        RECT 64.185 120.855 66.695 121.105 ;
        RECT 60.075 120.295 60.260 120.385 ;
        RECT 60.850 120.295 61.685 120.305 ;
        RECT 60.075 120.095 61.685 120.295 ;
        RECT 60.075 120.055 60.305 120.095 ;
        RECT 59.570 119.715 59.905 119.935 ;
        RECT 60.910 119.545 61.265 119.925 ;
        RECT 61.435 119.715 61.685 120.095 ;
        RECT 61.935 119.545 62.185 120.325 ;
        RECT 62.355 119.715 62.615 120.395 ;
        RECT 63.705 119.545 63.995 120.710 ;
        RECT 66.865 120.685 67.215 121.275 ;
        RECT 64.210 119.545 64.505 120.685 ;
        RECT 64.765 120.515 67.215 120.685 ;
        RECT 67.385 121.355 67.765 121.440 ;
        RECT 68.275 121.355 68.605 121.880 ;
        RECT 68.865 121.565 69.075 122.095 ;
        RECT 69.350 121.645 70.135 121.815 ;
        RECT 70.305 121.645 70.710 121.815 ;
        RECT 67.385 121.315 67.610 121.355 ;
        RECT 67.385 120.735 67.555 121.315 ;
        RECT 68.275 121.185 68.475 121.355 ;
        RECT 69.350 121.185 69.520 121.645 ;
        RECT 67.725 120.855 68.475 121.185 ;
        RECT 68.645 120.855 69.520 121.185 ;
        RECT 67.385 120.685 67.600 120.735 ;
        RECT 67.385 120.605 67.775 120.685 ;
        RECT 64.765 119.715 65.095 120.515 ;
        RECT 65.265 119.545 65.435 120.345 ;
        RECT 65.605 119.715 65.935 120.515 ;
        RECT 66.445 120.495 67.215 120.515 ;
        RECT 66.105 119.545 66.275 120.345 ;
        RECT 66.445 119.715 66.775 120.495 ;
        RECT 66.945 119.545 67.115 120.005 ;
        RECT 67.445 119.760 67.775 120.605 ;
        RECT 68.285 120.650 68.475 120.855 ;
        RECT 67.945 119.545 68.115 120.555 ;
        RECT 68.285 120.275 69.180 120.650 ;
        RECT 68.285 119.715 68.625 120.275 ;
        RECT 68.855 119.545 69.170 120.045 ;
        RECT 69.350 120.015 69.520 120.855 ;
        RECT 69.690 121.145 70.155 121.475 ;
        RECT 70.540 121.415 70.710 121.645 ;
        RECT 70.890 121.595 71.260 122.095 ;
        RECT 71.580 121.645 72.255 121.815 ;
        RECT 72.450 121.645 72.785 121.815 ;
        RECT 69.690 120.185 70.010 121.145 ;
        RECT 70.540 121.115 71.370 121.415 ;
        RECT 70.180 120.215 70.370 120.935 ;
        RECT 70.540 120.045 70.710 121.115 ;
        RECT 71.170 121.085 71.370 121.115 ;
        RECT 70.880 120.865 71.050 120.935 ;
        RECT 71.580 120.865 71.750 121.645 ;
        RECT 72.615 121.505 72.785 121.645 ;
        RECT 72.955 121.635 73.205 122.095 ;
        RECT 70.880 120.695 71.750 120.865 ;
        RECT 71.920 121.225 72.445 121.445 ;
        RECT 72.615 121.375 72.840 121.505 ;
        RECT 70.880 120.605 71.390 120.695 ;
        RECT 69.350 119.845 70.235 120.015 ;
        RECT 70.460 119.715 70.710 120.045 ;
        RECT 70.880 119.545 71.050 120.345 ;
        RECT 71.220 119.990 71.390 120.605 ;
        RECT 71.920 120.525 72.090 121.225 ;
        RECT 71.560 120.160 72.090 120.525 ;
        RECT 72.260 120.460 72.500 121.055 ;
        RECT 72.670 120.270 72.840 121.375 ;
        RECT 73.010 120.515 73.290 121.465 ;
        RECT 72.535 120.140 72.840 120.270 ;
        RECT 71.220 119.820 72.325 119.990 ;
        RECT 72.535 119.715 72.785 120.140 ;
        RECT 72.955 119.545 73.220 120.005 ;
        RECT 73.460 119.715 73.645 121.835 ;
        RECT 73.815 121.715 74.145 122.095 ;
        RECT 74.315 121.545 74.485 121.835 ;
        RECT 73.820 121.375 74.485 121.545 ;
        RECT 73.820 120.385 74.050 121.375 ;
        RECT 74.745 121.295 75.440 121.925 ;
        RECT 75.645 121.295 75.955 122.095 ;
        RECT 76.215 121.545 76.385 121.835 ;
        RECT 76.555 121.715 76.885 122.095 ;
        RECT 76.215 121.375 76.880 121.545 ;
        RECT 75.265 121.245 75.440 121.295 ;
        RECT 74.220 120.555 74.570 121.205 ;
        RECT 74.765 120.855 75.100 121.105 ;
        RECT 75.270 120.695 75.440 121.245 ;
        RECT 75.610 120.855 75.945 121.125 ;
        RECT 73.820 120.215 74.485 120.385 ;
        RECT 73.815 119.545 74.145 120.045 ;
        RECT 74.315 119.715 74.485 120.215 ;
        RECT 74.745 119.545 75.005 120.685 ;
        RECT 75.175 119.715 75.505 120.695 ;
        RECT 75.675 119.545 75.955 120.685 ;
        RECT 76.130 120.555 76.480 121.205 ;
        RECT 76.650 120.385 76.880 121.375 ;
        RECT 76.215 120.215 76.880 120.385 ;
        RECT 76.215 119.715 76.385 120.215 ;
        RECT 76.555 119.545 76.885 120.045 ;
        RECT 77.055 119.715 77.240 121.835 ;
        RECT 77.495 121.635 77.745 122.095 ;
        RECT 77.915 121.645 78.250 121.815 ;
        RECT 78.445 121.645 79.120 121.815 ;
        RECT 77.915 121.505 78.085 121.645 ;
        RECT 77.410 120.515 77.690 121.465 ;
        RECT 77.860 121.375 78.085 121.505 ;
        RECT 77.860 120.270 78.030 121.375 ;
        RECT 78.255 121.225 78.780 121.445 ;
        RECT 78.200 120.460 78.440 121.055 ;
        RECT 78.610 120.525 78.780 121.225 ;
        RECT 78.950 120.865 79.120 121.645 ;
        RECT 79.440 121.595 79.810 122.095 ;
        RECT 79.990 121.645 80.395 121.815 ;
        RECT 80.565 121.645 81.350 121.815 ;
        RECT 79.990 121.415 80.160 121.645 ;
        RECT 79.330 121.115 80.160 121.415 ;
        RECT 80.545 121.145 81.010 121.475 ;
        RECT 79.330 121.085 79.530 121.115 ;
        RECT 79.650 120.865 79.820 120.935 ;
        RECT 78.950 120.695 79.820 120.865 ;
        RECT 79.310 120.605 79.820 120.695 ;
        RECT 77.860 120.140 78.165 120.270 ;
        RECT 78.610 120.160 79.140 120.525 ;
        RECT 77.480 119.545 77.745 120.005 ;
        RECT 77.915 119.715 78.165 120.140 ;
        RECT 79.310 119.990 79.480 120.605 ;
        RECT 78.375 119.820 79.480 119.990 ;
        RECT 79.650 119.545 79.820 120.345 ;
        RECT 79.990 120.045 80.160 121.115 ;
        RECT 80.330 120.215 80.520 120.935 ;
        RECT 80.690 120.185 81.010 121.145 ;
        RECT 81.180 121.185 81.350 121.645 ;
        RECT 81.625 121.565 81.835 122.095 ;
        RECT 82.095 121.355 82.425 121.880 ;
        RECT 82.595 121.485 82.765 122.095 ;
        RECT 82.935 121.440 83.265 121.875 ;
        RECT 82.935 121.355 83.315 121.440 ;
        RECT 82.225 121.185 82.425 121.355 ;
        RECT 83.090 121.315 83.315 121.355 ;
        RECT 81.180 120.855 82.055 121.185 ;
        RECT 82.225 120.855 82.975 121.185 ;
        RECT 79.990 119.715 80.240 120.045 ;
        RECT 81.180 120.015 81.350 120.855 ;
        RECT 82.225 120.650 82.415 120.855 ;
        RECT 83.145 120.735 83.315 121.315 ;
        RECT 83.100 120.685 83.315 120.735 ;
        RECT 81.520 120.275 82.415 120.650 ;
        RECT 82.925 120.605 83.315 120.685 ;
        RECT 83.520 121.355 84.135 121.925 ;
        RECT 84.305 121.585 84.520 122.095 ;
        RECT 84.750 121.585 85.030 121.915 ;
        RECT 85.210 121.585 85.450 122.095 ;
        RECT 85.950 121.585 86.190 122.095 ;
        RECT 86.370 121.585 86.650 121.915 ;
        RECT 86.880 121.585 87.095 122.095 ;
        RECT 80.465 119.845 81.350 120.015 ;
        RECT 81.530 119.545 81.845 120.045 ;
        RECT 82.075 119.715 82.415 120.275 ;
        RECT 82.585 119.545 82.755 120.555 ;
        RECT 82.925 119.760 83.255 120.605 ;
        RECT 83.520 120.335 83.835 121.355 ;
        RECT 84.005 120.685 84.175 121.185 ;
        RECT 84.425 120.855 84.690 121.415 ;
        RECT 84.860 120.685 85.030 121.585 ;
        RECT 85.200 120.855 85.555 121.415 ;
        RECT 85.845 120.855 86.200 121.415 ;
        RECT 86.370 120.685 86.540 121.585 ;
        RECT 86.710 120.855 86.975 121.415 ;
        RECT 87.265 121.355 87.880 121.925 ;
        RECT 87.225 120.685 87.395 121.185 ;
        RECT 84.005 120.515 85.430 120.685 ;
        RECT 83.520 119.715 84.055 120.335 ;
        RECT 84.225 119.545 84.555 120.345 ;
        RECT 85.040 120.340 85.430 120.515 ;
        RECT 85.970 120.515 87.395 120.685 ;
        RECT 85.970 120.340 86.360 120.515 ;
        RECT 86.845 119.545 87.175 120.345 ;
        RECT 87.565 120.335 87.880 121.355 ;
        RECT 88.545 121.345 89.755 122.095 ;
        RECT 87.345 119.715 87.880 120.335 ;
        RECT 88.545 120.635 89.065 121.175 ;
        RECT 89.235 120.805 89.755 121.345 ;
        RECT 100.130 121.790 106.380 122.350 ;
        RECT 100.130 121.770 105.300 121.790 ;
        RECT 100.130 121.700 104.120 121.770 ;
        RECT 88.545 119.545 89.755 120.635 ;
        RECT 100.130 120.430 102.050 121.700 ;
        RECT 103.560 121.690 104.120 121.700 ;
        RECT 103.790 120.600 104.120 121.690 ;
        RECT 104.490 121.220 105.530 121.390 ;
        RECT 104.490 120.780 105.530 120.950 ;
        RECT 105.700 120.920 105.870 121.250 ;
        RECT 103.950 120.380 104.120 120.600 ;
        RECT 106.210 120.380 106.380 121.790 ;
        RECT 103.950 120.210 106.380 120.380 ;
        RECT 107.960 122.300 118.590 122.470 ;
        RECT 120.020 131.640 126.250 131.800 ;
        RECT 120.020 129.380 120.690 131.640 ;
        RECT 121.360 131.070 125.400 131.240 ;
        RECT 121.020 130.010 121.190 131.010 ;
        RECT 125.570 130.010 125.740 131.010 ;
        RECT 121.360 129.780 125.400 129.950 ;
        RECT 126.080 129.380 126.250 131.640 ;
        RECT 120.020 129.210 126.250 129.380 ;
        RECT 120.020 125.950 120.690 129.210 ;
        RECT 121.360 128.640 125.400 128.810 ;
        RECT 121.020 126.580 121.190 128.580 ;
        RECT 125.570 126.580 125.740 128.580 ;
        RECT 121.360 126.350 125.400 126.520 ;
        RECT 126.080 125.950 126.250 129.210 ;
        RECT 120.020 125.780 126.250 125.950 ;
        RECT 120.020 122.520 120.690 125.780 ;
        RECT 121.360 125.210 125.400 125.380 ;
        RECT 121.020 123.150 121.190 125.150 ;
        RECT 125.570 123.150 125.740 125.150 ;
        RECT 121.360 122.920 125.400 123.090 ;
        RECT 126.080 122.520 126.250 125.780 ;
        RECT 120.020 122.510 126.250 122.520 ;
        RECT 127.840 131.780 137.670 131.820 ;
        RECT 140.540 131.800 146.280 131.810 ;
        RECT 127.840 131.650 138.470 131.780 ;
        RECT 127.840 129.390 128.010 131.650 ;
        RECT 128.735 131.080 136.775 131.250 ;
        RECT 128.350 130.020 128.520 131.020 ;
        RECT 136.990 130.020 137.160 131.020 ;
        RECT 128.735 129.790 136.775 129.960 ;
        RECT 137.500 129.390 138.470 131.650 ;
        RECT 127.840 129.220 138.470 129.390 ;
        RECT 127.840 125.960 128.010 129.220 ;
        RECT 128.735 128.650 136.775 128.820 ;
        RECT 128.350 126.590 128.520 128.590 ;
        RECT 136.990 126.590 137.160 128.590 ;
        RECT 128.735 126.360 136.775 126.530 ;
        RECT 137.500 125.960 138.470 129.220 ;
        RECT 127.840 125.790 138.470 125.960 ;
        RECT 127.840 122.530 128.010 125.790 ;
        RECT 128.735 125.220 136.775 125.390 ;
        RECT 128.350 123.160 128.520 125.160 ;
        RECT 136.990 123.160 137.160 125.160 ;
        RECT 128.735 122.930 136.775 123.100 ;
        RECT 137.500 122.530 138.470 125.790 ;
        RECT 120.020 122.410 126.260 122.510 ;
        RECT 107.960 120.040 108.130 122.300 ;
        RECT 108.855 121.730 116.895 121.900 ;
        RECT 108.470 120.670 108.640 121.670 ;
        RECT 117.110 120.670 117.280 121.670 ;
        RECT 108.855 120.440 116.895 120.610 ;
        RECT 117.620 120.040 118.590 122.300 ;
        RECT 120.010 121.850 126.260 122.410 ;
        RECT 120.010 121.830 125.180 121.850 ;
        RECT 120.010 121.760 124.000 121.830 ;
        RECT 120.010 120.490 121.930 121.760 ;
        RECT 123.440 121.750 124.000 121.760 ;
        RECT 123.670 120.660 124.000 121.750 ;
        RECT 124.370 121.280 125.410 121.450 ;
        RECT 124.370 120.840 125.410 121.010 ;
        RECT 125.580 120.980 125.750 121.310 ;
        RECT 123.830 120.440 124.000 120.660 ;
        RECT 126.090 120.440 126.260 121.850 ;
        RECT 123.830 120.270 126.260 120.440 ;
        RECT 127.840 122.360 138.470 122.530 ;
        RECT 140.050 131.640 146.280 131.800 ;
        RECT 140.050 129.380 140.720 131.640 ;
        RECT 141.390 131.070 145.430 131.240 ;
        RECT 141.050 130.010 141.220 131.010 ;
        RECT 145.600 130.010 145.770 131.010 ;
        RECT 141.390 129.780 145.430 129.950 ;
        RECT 146.110 129.380 146.280 131.640 ;
        RECT 140.050 129.210 146.280 129.380 ;
        RECT 140.050 125.950 140.720 129.210 ;
        RECT 141.390 128.640 145.430 128.810 ;
        RECT 141.050 126.580 141.220 128.580 ;
        RECT 145.600 126.580 145.770 128.580 ;
        RECT 141.390 126.350 145.430 126.520 ;
        RECT 146.110 125.950 146.280 129.210 ;
        RECT 140.050 125.780 146.280 125.950 ;
        RECT 140.050 122.520 140.720 125.780 ;
        RECT 141.390 125.210 145.430 125.380 ;
        RECT 141.050 123.150 141.220 125.150 ;
        RECT 145.600 123.150 145.770 125.150 ;
        RECT 141.390 122.920 145.430 123.090 ;
        RECT 146.110 122.520 146.280 125.780 ;
        RECT 140.050 122.510 146.280 122.520 ;
        RECT 147.870 131.780 157.700 131.820 ;
        RECT 147.870 131.650 158.500 131.780 ;
        RECT 147.870 129.390 148.040 131.650 ;
        RECT 148.765 131.080 156.805 131.250 ;
        RECT 148.380 130.020 148.550 131.020 ;
        RECT 157.020 130.020 157.190 131.020 ;
        RECT 148.765 129.790 156.805 129.960 ;
        RECT 157.530 129.390 158.500 131.650 ;
        RECT 147.870 129.220 158.500 129.390 ;
        RECT 147.870 125.960 148.040 129.220 ;
        RECT 148.765 128.650 156.805 128.820 ;
        RECT 148.380 126.590 148.550 128.590 ;
        RECT 157.020 126.590 157.190 128.590 ;
        RECT 148.765 126.360 156.805 126.530 ;
        RECT 157.530 125.960 158.500 129.220 ;
        RECT 147.870 125.790 158.500 125.960 ;
        RECT 147.870 122.530 148.040 125.790 ;
        RECT 148.765 125.220 156.805 125.390 ;
        RECT 148.380 123.160 148.550 125.160 ;
        RECT 157.020 123.160 157.190 125.160 ;
        RECT 148.765 122.930 156.805 123.100 ;
        RECT 157.530 122.530 158.500 125.790 ;
        RECT 140.050 122.410 146.290 122.510 ;
        RECT 127.840 120.100 128.010 122.360 ;
        RECT 128.735 121.790 136.775 121.960 ;
        RECT 128.350 120.730 128.520 121.730 ;
        RECT 136.990 120.730 137.160 121.730 ;
        RECT 128.735 120.500 136.775 120.670 ;
        RECT 137.500 120.100 138.470 122.360 ;
        RECT 140.040 121.850 146.290 122.410 ;
        RECT 140.040 121.830 145.210 121.850 ;
        RECT 140.040 121.760 144.030 121.830 ;
        RECT 140.040 120.490 141.960 121.760 ;
        RECT 143.470 121.750 144.030 121.760 ;
        RECT 143.700 120.660 144.030 121.750 ;
        RECT 144.400 121.280 145.440 121.450 ;
        RECT 144.400 120.840 145.440 121.010 ;
        RECT 145.610 120.980 145.780 121.310 ;
        RECT 143.860 120.440 144.030 120.660 ;
        RECT 146.120 120.440 146.290 121.850 ;
        RECT 143.860 120.270 146.290 120.440 ;
        RECT 147.870 122.360 158.500 122.530 ;
        RECT 127.840 120.070 138.470 120.100 ;
        RECT 147.870 120.100 148.040 122.360 ;
        RECT 148.765 121.790 156.805 121.960 ;
        RECT 148.380 120.730 148.550 121.730 ;
        RECT 157.020 120.730 157.190 121.730 ;
        RECT 148.765 120.500 156.805 120.670 ;
        RECT 157.530 120.100 158.500 122.360 ;
        RECT 147.870 120.070 158.500 120.100 ;
        RECT 107.960 120.010 118.590 120.040 ;
        RECT 107.930 119.900 118.590 120.010 ;
        RECT 127.810 119.960 138.470 120.070 ;
        RECT 147.840 119.960 158.500 120.070 ;
        RECT 126.060 119.910 138.470 119.960 ;
        RECT 146.090 119.910 158.500 119.960 ;
        RECT 106.180 119.850 118.590 119.900 ;
        RECT 101.840 119.680 118.590 119.850 ;
        RECT 12.100 119.375 89.840 119.545 ;
        RECT 12.185 118.285 13.395 119.375 ;
        RECT 13.565 118.940 18.910 119.375 ;
        RECT 12.185 117.575 12.705 118.115 ;
        RECT 12.875 117.745 13.395 118.285 ;
        RECT 12.185 116.825 13.395 117.575 ;
        RECT 15.150 117.370 15.490 118.200 ;
        RECT 16.970 117.690 17.320 118.940 ;
        RECT 19.085 118.285 21.675 119.375 ;
        RECT 21.845 118.865 22.145 119.375 ;
        RECT 22.315 118.695 22.645 119.205 ;
        RECT 22.815 118.865 23.445 119.375 ;
        RECT 24.025 118.865 24.405 119.035 ;
        RECT 24.575 118.865 24.875 119.375 ;
        RECT 24.235 118.695 24.405 118.865 ;
        RECT 19.085 117.595 20.295 118.115 ;
        RECT 20.465 117.765 21.675 118.285 ;
        RECT 21.845 118.525 24.065 118.695 ;
        RECT 13.565 116.825 18.910 117.370 ;
        RECT 19.085 116.825 21.675 117.595 ;
        RECT 21.845 117.565 22.015 118.525 ;
        RECT 22.185 118.185 23.725 118.355 ;
        RECT 22.185 117.735 22.430 118.185 ;
        RECT 22.690 117.815 23.385 118.015 ;
        RECT 23.555 117.985 23.725 118.185 ;
        RECT 23.895 118.325 24.065 118.525 ;
        RECT 24.235 118.495 24.895 118.695 ;
        RECT 23.895 118.155 24.555 118.325 ;
        RECT 23.555 117.815 24.155 117.985 ;
        RECT 24.385 117.735 24.555 118.155 ;
        RECT 21.845 117.020 22.310 117.565 ;
        RECT 22.815 116.825 22.985 117.645 ;
        RECT 23.155 117.565 24.065 117.645 ;
        RECT 24.725 117.565 24.895 118.495 ;
        RECT 25.065 118.210 25.355 119.375 ;
        RECT 26.535 118.365 26.705 119.205 ;
        RECT 26.875 119.035 28.045 119.205 ;
        RECT 26.875 118.535 27.205 119.035 ;
        RECT 27.715 118.995 28.045 119.035 ;
        RECT 28.235 118.955 28.590 119.375 ;
        RECT 27.375 118.775 27.605 118.865 ;
        RECT 28.760 118.775 29.010 119.205 ;
        RECT 27.375 118.535 29.010 118.775 ;
        RECT 29.180 118.615 29.510 119.375 ;
        RECT 29.680 118.535 29.935 119.205 ;
        RECT 30.755 118.575 31.010 119.375 ;
        RECT 26.535 118.195 29.595 118.365 ;
        RECT 26.450 117.815 26.800 118.025 ;
        RECT 26.970 117.815 27.415 118.015 ;
        RECT 27.585 117.815 28.060 118.015 ;
        RECT 23.155 117.475 24.405 117.565 ;
        RECT 23.155 116.995 23.485 117.475 ;
        RECT 23.895 117.395 24.405 117.475 ;
        RECT 23.655 116.825 24.005 117.215 ;
        RECT 24.175 116.995 24.405 117.395 ;
        RECT 24.575 117.085 24.895 117.565 ;
        RECT 25.065 116.825 25.355 117.550 ;
        RECT 26.535 117.475 27.600 117.645 ;
        RECT 26.535 116.995 26.705 117.475 ;
        RECT 26.875 116.825 27.205 117.305 ;
        RECT 27.430 117.245 27.600 117.475 ;
        RECT 27.780 117.415 28.060 117.815 ;
        RECT 28.330 117.815 28.660 118.015 ;
        RECT 28.830 117.845 29.205 118.015 ;
        RECT 28.830 117.815 29.195 117.845 ;
        RECT 28.330 117.415 28.615 117.815 ;
        RECT 29.425 117.645 29.595 118.195 ;
        RECT 28.795 117.475 29.595 117.645 ;
        RECT 28.795 117.245 28.965 117.475 ;
        RECT 29.765 117.405 29.935 118.535 ;
        RECT 31.180 118.405 31.510 119.205 ;
        RECT 31.680 118.575 31.850 119.375 ;
        RECT 32.020 118.405 32.350 119.205 ;
        RECT 32.520 118.575 32.690 119.375 ;
        RECT 32.860 118.405 33.190 119.205 ;
        RECT 33.360 118.575 33.530 119.375 ;
        RECT 33.700 118.405 34.030 119.205 ;
        RECT 34.200 118.575 34.500 119.375 ;
        RECT 30.585 118.235 34.555 118.405 ;
        RECT 34.735 118.265 35.030 119.375 ;
        RECT 30.585 117.645 30.930 118.235 ;
        RECT 31.180 117.815 34.035 118.065 ;
        RECT 34.235 117.645 34.555 118.235 ;
        RECT 35.210 118.065 35.460 119.200 ;
        RECT 35.630 118.265 35.890 119.375 ;
        RECT 36.060 118.475 36.320 119.200 ;
        RECT 36.490 118.645 36.750 119.375 ;
        RECT 36.920 118.475 37.180 119.200 ;
        RECT 37.350 118.645 37.610 119.375 ;
        RECT 37.780 118.475 38.040 119.200 ;
        RECT 38.210 118.645 38.470 119.375 ;
        RECT 38.640 118.475 38.900 119.200 ;
        RECT 39.070 118.645 39.365 119.375 ;
        RECT 36.060 118.235 39.370 118.475 ;
        RECT 39.785 118.235 40.065 119.375 ;
        RECT 30.585 117.455 34.555 117.645 ;
        RECT 34.725 117.455 35.040 118.065 ;
        RECT 35.210 117.815 38.230 118.065 ;
        RECT 29.750 117.335 29.935 117.405 ;
        RECT 29.725 117.325 29.935 117.335 ;
        RECT 27.430 116.995 28.965 117.245 ;
        RECT 29.135 116.825 29.465 117.305 ;
        RECT 29.680 116.995 29.935 117.325 ;
        RECT 30.755 116.825 31.010 117.285 ;
        RECT 31.180 116.995 31.510 117.455 ;
        RECT 31.680 116.825 31.850 117.285 ;
        RECT 32.020 116.995 32.350 117.455 ;
        RECT 32.520 116.825 32.690 117.285 ;
        RECT 32.860 116.995 33.190 117.455 ;
        RECT 33.360 116.825 33.530 117.285 ;
        RECT 33.700 116.995 34.030 117.455 ;
        RECT 34.200 116.825 34.505 117.285 ;
        RECT 34.785 116.825 35.030 117.285 ;
        RECT 35.210 117.005 35.460 117.815 ;
        RECT 38.400 117.645 39.370 118.235 ;
        RECT 40.235 118.225 40.565 119.205 ;
        RECT 40.735 118.235 40.995 119.375 ;
        RECT 41.255 118.705 41.425 119.205 ;
        RECT 41.595 118.875 41.925 119.375 ;
        RECT 41.255 118.535 41.920 118.705 ;
        RECT 39.795 117.795 40.130 118.065 ;
        RECT 36.060 117.475 39.370 117.645 ;
        RECT 40.300 117.625 40.470 118.225 ;
        RECT 40.640 117.815 40.975 118.065 ;
        RECT 41.170 117.715 41.520 118.365 ;
        RECT 35.630 116.825 35.890 117.350 ;
        RECT 36.060 117.020 36.320 117.475 ;
        RECT 36.490 116.825 36.750 117.305 ;
        RECT 36.920 117.020 37.180 117.475 ;
        RECT 37.350 116.825 37.610 117.305 ;
        RECT 37.780 117.020 38.040 117.475 ;
        RECT 38.210 116.825 38.470 117.305 ;
        RECT 38.640 117.020 38.900 117.475 ;
        RECT 39.070 116.825 39.370 117.305 ;
        RECT 39.785 116.825 40.095 117.625 ;
        RECT 40.300 116.995 40.995 117.625 ;
        RECT 41.690 117.545 41.920 118.535 ;
        RECT 41.255 117.375 41.920 117.545 ;
        RECT 41.255 117.085 41.425 117.375 ;
        RECT 41.595 116.825 41.925 117.205 ;
        RECT 42.095 117.085 42.280 119.205 ;
        RECT 42.520 118.915 42.785 119.375 ;
        RECT 42.955 118.780 43.205 119.205 ;
        RECT 43.415 118.930 44.520 119.100 ;
        RECT 42.900 118.650 43.205 118.780 ;
        RECT 42.450 117.455 42.730 118.405 ;
        RECT 42.900 117.545 43.070 118.650 ;
        RECT 43.240 117.865 43.480 118.460 ;
        RECT 43.650 118.395 44.180 118.760 ;
        RECT 43.650 117.695 43.820 118.395 ;
        RECT 44.350 118.315 44.520 118.930 ;
        RECT 44.690 118.575 44.860 119.375 ;
        RECT 45.030 118.875 45.280 119.205 ;
        RECT 45.505 118.905 46.390 119.075 ;
        RECT 44.350 118.225 44.860 118.315 ;
        RECT 42.900 117.415 43.125 117.545 ;
        RECT 43.295 117.475 43.820 117.695 ;
        RECT 43.990 118.055 44.860 118.225 ;
        RECT 42.535 116.825 42.785 117.285 ;
        RECT 42.955 117.275 43.125 117.415 ;
        RECT 43.990 117.275 44.160 118.055 ;
        RECT 44.690 117.985 44.860 118.055 ;
        RECT 44.370 117.805 44.570 117.835 ;
        RECT 45.030 117.805 45.200 118.875 ;
        RECT 45.370 117.985 45.560 118.705 ;
        RECT 44.370 117.505 45.200 117.805 ;
        RECT 45.730 117.775 46.050 118.735 ;
        RECT 42.955 117.105 43.290 117.275 ;
        RECT 43.485 117.105 44.160 117.275 ;
        RECT 44.480 116.825 44.850 117.325 ;
        RECT 45.030 117.275 45.200 117.505 ;
        RECT 45.585 117.445 46.050 117.775 ;
        RECT 46.220 118.065 46.390 118.905 ;
        RECT 46.570 118.875 46.885 119.375 ;
        RECT 47.115 118.645 47.455 119.205 ;
        RECT 46.560 118.270 47.455 118.645 ;
        RECT 47.625 118.365 47.795 119.375 ;
        RECT 47.265 118.065 47.455 118.270 ;
        RECT 47.965 118.315 48.295 119.160 ;
        RECT 47.965 118.235 48.355 118.315 ;
        RECT 48.525 118.285 50.195 119.375 ;
        RECT 48.140 118.185 48.355 118.235 ;
        RECT 46.220 117.735 47.095 118.065 ;
        RECT 47.265 117.735 48.015 118.065 ;
        RECT 46.220 117.275 46.390 117.735 ;
        RECT 47.265 117.565 47.465 117.735 ;
        RECT 48.185 117.605 48.355 118.185 ;
        RECT 48.130 117.565 48.355 117.605 ;
        RECT 45.030 117.105 45.435 117.275 ;
        RECT 45.605 117.105 46.390 117.275 ;
        RECT 46.665 116.825 46.875 117.355 ;
        RECT 47.135 117.040 47.465 117.565 ;
        RECT 47.975 117.480 48.355 117.565 ;
        RECT 48.525 117.595 49.275 118.115 ;
        RECT 49.445 117.765 50.195 118.285 ;
        RECT 50.825 118.210 51.115 119.375 ;
        RECT 51.290 118.235 51.625 119.205 ;
        RECT 51.795 118.235 51.965 119.375 ;
        RECT 52.135 119.035 54.165 119.205 ;
        RECT 47.635 116.825 47.805 117.435 ;
        RECT 47.975 117.045 48.305 117.480 ;
        RECT 48.525 116.825 50.195 117.595 ;
        RECT 51.290 117.565 51.460 118.235 ;
        RECT 52.135 118.065 52.305 119.035 ;
        RECT 51.630 117.735 51.885 118.065 ;
        RECT 52.110 117.735 52.305 118.065 ;
        RECT 52.475 118.695 53.600 118.865 ;
        RECT 51.715 117.565 51.885 117.735 ;
        RECT 52.475 117.565 52.645 118.695 ;
        RECT 50.825 116.825 51.115 117.550 ;
        RECT 51.290 116.995 51.545 117.565 ;
        RECT 51.715 117.395 52.645 117.565 ;
        RECT 52.815 118.355 53.825 118.525 ;
        RECT 52.815 117.555 52.985 118.355 ;
        RECT 52.470 117.360 52.645 117.395 ;
        RECT 51.715 116.825 52.045 117.225 ;
        RECT 52.470 116.995 53.000 117.360 ;
        RECT 53.190 117.335 53.465 118.155 ;
        RECT 53.185 117.165 53.465 117.335 ;
        RECT 53.190 116.995 53.465 117.165 ;
        RECT 53.635 116.995 53.825 118.355 ;
        RECT 53.995 118.370 54.165 119.035 ;
        RECT 54.335 118.615 54.505 119.375 ;
        RECT 54.740 118.615 55.255 119.025 ;
        RECT 53.995 118.180 54.745 118.370 ;
        RECT 54.915 117.805 55.255 118.615 ;
        RECT 55.465 118.425 55.755 119.195 ;
        RECT 56.325 118.835 56.585 119.195 ;
        RECT 56.755 119.005 57.085 119.375 ;
        RECT 57.255 118.835 57.515 119.195 ;
        RECT 56.325 118.605 57.515 118.835 ;
        RECT 57.705 118.655 58.035 119.375 ;
        RECT 58.205 118.425 58.470 119.195 ;
        RECT 59.305 118.705 59.585 119.375 ;
        RECT 59.755 118.485 60.055 119.035 ;
        RECT 60.255 118.655 60.585 119.375 ;
        RECT 60.775 118.655 61.235 119.205 ;
        RECT 55.465 118.245 57.960 118.425 ;
        RECT 54.025 117.635 55.255 117.805 ;
        RECT 55.435 117.735 55.705 118.065 ;
        RECT 55.885 117.735 56.320 118.065 ;
        RECT 56.500 117.735 57.075 118.065 ;
        RECT 57.255 117.735 57.535 118.065 ;
        RECT 54.005 116.825 54.515 117.360 ;
        RECT 54.735 117.030 54.980 117.635 ;
        RECT 57.735 117.555 57.960 118.245 ;
        RECT 55.475 117.365 57.960 117.555 ;
        RECT 55.475 117.005 55.700 117.365 ;
        RECT 55.880 116.825 56.210 117.195 ;
        RECT 56.390 117.005 56.645 117.365 ;
        RECT 57.210 116.825 57.955 117.195 ;
        RECT 58.135 117.005 58.470 118.425 ;
        RECT 59.120 118.065 59.385 118.425 ;
        RECT 59.755 118.315 60.695 118.485 ;
        RECT 60.525 118.065 60.695 118.315 ;
        RECT 59.120 117.815 59.795 118.065 ;
        RECT 60.015 117.815 60.355 118.065 ;
        RECT 60.525 117.735 60.815 118.065 ;
        RECT 60.525 117.645 60.695 117.735 ;
        RECT 59.305 117.455 60.695 117.645 ;
        RECT 59.305 117.095 59.635 117.455 ;
        RECT 60.985 117.285 61.235 118.655 ;
        RECT 61.415 118.265 61.710 119.375 ;
        RECT 61.890 118.065 62.140 119.200 ;
        RECT 62.310 118.265 62.570 119.375 ;
        RECT 62.740 118.475 63.000 119.200 ;
        RECT 63.170 118.645 63.430 119.375 ;
        RECT 63.600 118.475 63.860 119.200 ;
        RECT 64.030 118.645 64.290 119.375 ;
        RECT 64.460 118.475 64.720 119.200 ;
        RECT 64.890 118.645 65.150 119.375 ;
        RECT 65.320 118.475 65.580 119.200 ;
        RECT 65.750 118.645 66.045 119.375 ;
        RECT 62.740 118.235 66.050 118.475 ;
        RECT 61.405 117.455 61.720 118.065 ;
        RECT 61.890 117.815 64.910 118.065 ;
        RECT 60.255 116.825 60.505 117.285 ;
        RECT 60.675 116.995 61.235 117.285 ;
        RECT 61.465 116.825 61.710 117.285 ;
        RECT 61.890 117.005 62.140 117.815 ;
        RECT 65.080 117.645 66.050 118.235 ;
        RECT 62.740 117.475 66.050 117.645 ;
        RECT 66.475 118.315 66.805 119.165 ;
        RECT 66.475 117.550 66.665 118.315 ;
        RECT 66.975 118.235 67.225 119.375 ;
        RECT 67.415 118.735 67.665 119.155 ;
        RECT 67.895 118.905 68.225 119.375 ;
        RECT 68.455 118.735 68.705 119.155 ;
        RECT 67.415 118.565 68.705 118.735 ;
        RECT 68.885 118.735 69.215 119.165 ;
        RECT 68.885 118.565 69.340 118.735 ;
        RECT 67.405 118.065 67.620 118.395 ;
        RECT 66.835 117.735 67.145 118.065 ;
        RECT 67.315 117.735 67.620 118.065 ;
        RECT 67.795 117.735 68.080 118.395 ;
        RECT 68.275 117.735 68.540 118.395 ;
        RECT 68.755 117.735 69.000 118.395 ;
        RECT 66.975 117.565 67.145 117.735 ;
        RECT 69.170 117.565 69.340 118.565 ;
        RECT 70.605 118.615 71.120 119.025 ;
        RECT 71.355 118.615 71.525 119.375 ;
        RECT 71.695 119.035 73.725 119.205 ;
        RECT 70.605 117.805 70.945 118.615 ;
        RECT 71.695 118.370 71.865 119.035 ;
        RECT 72.260 118.695 73.385 118.865 ;
        RECT 71.115 118.180 71.865 118.370 ;
        RECT 72.035 118.355 73.045 118.525 ;
        RECT 70.605 117.635 71.835 117.805 ;
        RECT 62.310 116.825 62.570 117.350 ;
        RECT 62.740 117.020 63.000 117.475 ;
        RECT 63.170 116.825 63.430 117.305 ;
        RECT 63.600 117.020 63.860 117.475 ;
        RECT 64.030 116.825 64.290 117.305 ;
        RECT 64.460 117.020 64.720 117.475 ;
        RECT 64.890 116.825 65.150 117.305 ;
        RECT 65.320 117.020 65.580 117.475 ;
        RECT 65.750 116.825 66.050 117.305 ;
        RECT 66.475 117.040 66.805 117.550 ;
        RECT 66.975 117.395 69.340 117.565 ;
        RECT 66.975 116.825 67.305 117.225 ;
        RECT 68.355 117.055 68.685 117.395 ;
        RECT 68.855 116.825 69.185 117.225 ;
        RECT 70.880 117.030 71.125 117.635 ;
        RECT 71.345 116.825 71.855 117.360 ;
        RECT 72.035 116.995 72.225 118.355 ;
        RECT 72.395 118.015 72.670 118.155 ;
        RECT 72.395 117.845 72.675 118.015 ;
        RECT 72.395 116.995 72.670 117.845 ;
        RECT 72.875 117.555 73.045 118.355 ;
        RECT 73.215 117.565 73.385 118.695 ;
        RECT 73.555 118.065 73.725 119.035 ;
        RECT 73.895 118.235 74.065 119.375 ;
        RECT 74.235 118.235 74.570 119.205 ;
        RECT 73.555 117.735 73.750 118.065 ;
        RECT 73.975 117.735 74.230 118.065 ;
        RECT 73.975 117.565 74.145 117.735 ;
        RECT 74.400 117.565 74.570 118.235 ;
        RECT 74.750 118.225 75.010 119.375 ;
        RECT 75.185 118.300 75.440 119.205 ;
        RECT 75.610 118.615 75.940 119.375 ;
        RECT 76.155 118.445 76.325 119.205 ;
        RECT 73.215 117.395 74.145 117.565 ;
        RECT 73.215 117.360 73.390 117.395 ;
        RECT 72.860 116.995 73.390 117.360 ;
        RECT 73.815 116.825 74.145 117.225 ;
        RECT 74.315 116.995 74.570 117.565 ;
        RECT 74.750 116.825 75.010 117.665 ;
        RECT 75.185 117.570 75.355 118.300 ;
        RECT 75.610 118.275 76.325 118.445 ;
        RECT 75.610 118.065 75.780 118.275 ;
        RECT 76.585 118.210 76.875 119.375 ;
        RECT 77.055 118.265 77.350 119.375 ;
        RECT 75.525 117.735 75.780 118.065 ;
        RECT 75.185 116.995 75.440 117.570 ;
        RECT 75.610 117.545 75.780 117.735 ;
        RECT 76.060 117.725 76.415 118.095 ;
        RECT 77.530 118.065 77.780 119.200 ;
        RECT 77.950 118.265 78.210 119.375 ;
        RECT 78.380 118.475 78.640 119.200 ;
        RECT 78.810 118.645 79.070 119.375 ;
        RECT 79.240 118.475 79.500 119.200 ;
        RECT 79.670 118.645 79.930 119.375 ;
        RECT 80.100 118.475 80.360 119.200 ;
        RECT 80.530 118.645 80.790 119.375 ;
        RECT 80.960 118.475 81.220 119.200 ;
        RECT 81.390 118.645 81.685 119.375 ;
        RECT 78.380 118.235 81.690 118.475 ;
        RECT 75.610 117.375 76.325 117.545 ;
        RECT 75.610 116.825 75.940 117.205 ;
        RECT 76.155 116.995 76.325 117.375 ;
        RECT 76.585 116.825 76.875 117.550 ;
        RECT 77.045 117.455 77.360 118.065 ;
        RECT 77.530 117.815 80.550 118.065 ;
        RECT 77.105 116.825 77.350 117.285 ;
        RECT 77.530 117.005 77.780 117.815 ;
        RECT 80.720 117.645 81.690 118.235 ;
        RECT 82.110 118.225 82.370 119.375 ;
        RECT 82.545 118.300 82.800 119.205 ;
        RECT 82.970 118.615 83.300 119.375 ;
        RECT 83.515 118.445 83.685 119.205 ;
        RECT 78.380 117.475 81.690 117.645 ;
        RECT 77.950 116.825 78.210 117.350 ;
        RECT 78.380 117.020 78.640 117.475 ;
        RECT 78.810 116.825 79.070 117.305 ;
        RECT 79.240 117.020 79.500 117.475 ;
        RECT 79.670 116.825 79.930 117.305 ;
        RECT 80.100 117.020 80.360 117.475 ;
        RECT 80.530 116.825 80.790 117.305 ;
        RECT 80.960 117.020 81.220 117.475 ;
        RECT 81.390 116.825 81.690 117.305 ;
        RECT 82.110 116.825 82.370 117.665 ;
        RECT 82.545 117.570 82.715 118.300 ;
        RECT 82.970 118.275 83.685 118.445 ;
        RECT 84.955 118.445 85.125 119.205 ;
        RECT 85.340 118.615 85.670 119.375 ;
        RECT 84.955 118.275 85.670 118.445 ;
        RECT 85.840 118.300 86.095 119.205 ;
        RECT 82.970 118.065 83.140 118.275 ;
        RECT 82.885 117.735 83.140 118.065 ;
        RECT 82.545 116.995 82.800 117.570 ;
        RECT 82.970 117.545 83.140 117.735 ;
        RECT 83.420 117.725 83.775 118.095 ;
        RECT 84.865 117.725 85.220 118.095 ;
        RECT 85.500 118.065 85.670 118.275 ;
        RECT 85.500 117.735 85.755 118.065 ;
        RECT 85.500 117.545 85.670 117.735 ;
        RECT 85.925 117.570 86.095 118.300 ;
        RECT 86.270 118.225 86.530 119.375 ;
        RECT 86.795 118.445 86.965 119.205 ;
        RECT 87.180 118.615 87.510 119.375 ;
        RECT 86.795 118.275 87.510 118.445 ;
        RECT 87.680 118.300 87.935 119.205 ;
        RECT 86.705 117.725 87.060 118.095 ;
        RECT 87.340 118.065 87.510 118.275 ;
        RECT 87.340 117.735 87.595 118.065 ;
        RECT 82.970 117.375 83.685 117.545 ;
        RECT 82.970 116.825 83.300 117.205 ;
        RECT 83.515 116.995 83.685 117.375 ;
        RECT 84.955 117.375 85.670 117.545 ;
        RECT 84.955 116.995 85.125 117.375 ;
        RECT 85.340 116.825 85.670 117.205 ;
        RECT 85.840 116.995 86.095 117.570 ;
        RECT 86.270 116.825 86.530 117.665 ;
        RECT 87.340 117.545 87.510 117.735 ;
        RECT 87.765 117.570 87.935 118.300 ;
        RECT 88.110 118.225 88.370 119.375 ;
        RECT 88.545 118.285 89.755 119.375 ;
        RECT 88.545 117.745 89.065 118.285 ;
        RECT 101.840 118.270 102.010 119.680 ;
        RECT 102.380 119.110 105.420 119.280 ;
        RECT 102.380 118.670 105.420 118.840 ;
        RECT 105.635 118.810 105.805 119.140 ;
        RECT 106.140 118.920 118.590 119.680 ;
        RECT 121.720 119.740 138.470 119.910 ;
        RECT 106.140 118.910 118.480 118.920 ;
        RECT 106.140 118.900 112.020 118.910 ;
        RECT 106.140 118.880 106.710 118.900 ;
        RECT 107.930 118.890 112.020 118.900 ;
        RECT 106.150 118.270 106.320 118.880 ;
        RECT 86.795 117.375 87.510 117.545 ;
        RECT 86.795 116.995 86.965 117.375 ;
        RECT 87.180 116.825 87.510 117.205 ;
        RECT 87.680 116.995 87.935 117.570 ;
        RECT 88.110 116.825 88.370 117.665 ;
        RECT 89.235 117.575 89.755 118.115 ;
        RECT 101.840 118.100 106.320 118.270 ;
        RECT 121.720 118.330 121.890 119.740 ;
        RECT 122.260 119.170 125.300 119.340 ;
        RECT 122.260 118.730 125.300 118.900 ;
        RECT 125.515 118.870 125.685 119.200 ;
        RECT 126.020 118.980 138.470 119.740 ;
        RECT 141.750 119.740 158.500 119.910 ;
        RECT 126.020 118.970 138.360 118.980 ;
        RECT 126.020 118.960 131.900 118.970 ;
        RECT 126.020 118.940 126.590 118.960 ;
        RECT 127.810 118.950 131.900 118.960 ;
        RECT 126.030 118.330 126.200 118.940 ;
        RECT 121.720 118.160 126.200 118.330 ;
        RECT 141.750 118.330 141.920 119.740 ;
        RECT 142.290 119.170 145.330 119.340 ;
        RECT 142.290 118.730 145.330 118.900 ;
        RECT 145.545 118.870 145.715 119.200 ;
        RECT 146.050 118.980 158.500 119.740 ;
        RECT 146.050 118.970 158.390 118.980 ;
        RECT 146.050 118.960 151.930 118.970 ;
        RECT 146.050 118.940 146.620 118.960 ;
        RECT 147.840 118.950 151.930 118.960 ;
        RECT 146.060 118.330 146.230 118.940 ;
        RECT 141.750 118.160 146.230 118.330 ;
        RECT 88.545 116.825 89.755 117.575 ;
        RECT 12.100 116.655 89.840 116.825 ;
        RECT 100.580 116.800 106.320 116.810 ;
        RECT 12.185 115.905 13.395 116.655 ;
        RECT 13.655 116.105 13.825 116.485 ;
        RECT 14.005 116.275 14.335 116.655 ;
        RECT 13.655 115.935 14.320 116.105 ;
        RECT 14.515 115.980 14.775 116.485 ;
        RECT 14.945 116.110 20.290 116.655 ;
        RECT 12.185 115.365 12.705 115.905 ;
        RECT 12.875 115.195 13.395 115.735 ;
        RECT 13.585 115.385 13.925 115.755 ;
        RECT 14.150 115.680 14.320 115.935 ;
        RECT 14.150 115.350 14.425 115.680 ;
        RECT 14.150 115.205 14.320 115.350 ;
        RECT 12.185 114.105 13.395 115.195 ;
        RECT 13.645 115.035 14.320 115.205 ;
        RECT 14.595 115.180 14.775 115.980 ;
        RECT 16.530 115.280 16.870 116.110 ;
        RECT 20.935 115.845 21.205 116.655 ;
        RECT 21.375 115.845 21.705 116.485 ;
        RECT 21.875 115.845 22.115 116.655 ;
        RECT 22.770 115.890 23.225 116.655 ;
        RECT 23.500 116.275 24.800 116.485 ;
        RECT 25.055 116.295 25.385 116.655 ;
        RECT 24.630 116.125 24.800 116.275 ;
        RECT 25.555 116.155 25.815 116.485 ;
        RECT 13.645 114.275 13.825 115.035 ;
        RECT 14.005 114.105 14.335 114.865 ;
        RECT 14.505 114.275 14.775 115.180 ;
        RECT 18.350 114.540 18.700 115.790 ;
        RECT 20.925 115.415 21.275 115.665 ;
        RECT 21.445 115.245 21.615 115.845 ;
        RECT 23.700 115.665 23.920 116.065 ;
        RECT 21.785 115.415 22.135 115.665 ;
        RECT 22.765 115.465 23.255 115.665 ;
        RECT 23.445 115.455 23.920 115.665 ;
        RECT 24.165 115.665 24.375 116.065 ;
        RECT 24.630 116.000 25.385 116.125 ;
        RECT 24.630 115.955 25.475 116.000 ;
        RECT 25.205 115.835 25.475 115.955 ;
        RECT 24.165 115.455 24.495 115.665 ;
        RECT 24.665 115.395 25.075 115.700 ;
        RECT 14.945 114.105 20.290 114.540 ;
        RECT 20.935 114.105 21.265 115.245 ;
        RECT 21.445 115.075 22.125 115.245 ;
        RECT 21.795 114.290 22.125 115.075 ;
        RECT 22.770 115.225 23.945 115.285 ;
        RECT 25.305 115.260 25.475 115.835 ;
        RECT 25.275 115.225 25.475 115.260 ;
        RECT 22.770 115.115 25.475 115.225 ;
        RECT 22.770 114.495 23.025 115.115 ;
        RECT 23.615 115.055 25.415 115.115 ;
        RECT 23.615 115.025 23.945 115.055 ;
        RECT 25.645 114.955 25.815 116.155 ;
        RECT 23.275 114.855 23.460 114.945 ;
        RECT 24.050 114.855 24.885 114.865 ;
        RECT 23.275 114.655 24.885 114.855 ;
        RECT 23.275 114.615 23.505 114.655 ;
        RECT 22.770 114.275 23.105 114.495 ;
        RECT 24.110 114.105 24.465 114.485 ;
        RECT 24.635 114.275 24.885 114.655 ;
        RECT 25.135 114.105 25.385 114.885 ;
        RECT 25.555 114.275 25.815 114.955 ;
        RECT 25.990 115.055 26.325 116.475 ;
        RECT 26.505 116.285 27.250 116.655 ;
        RECT 27.815 116.115 28.070 116.475 ;
        RECT 28.250 116.285 28.580 116.655 ;
        RECT 28.760 116.115 28.985 116.475 ;
        RECT 26.500 115.925 28.985 116.115 ;
        RECT 26.500 115.235 26.725 115.925 ;
        RECT 29.240 115.915 29.855 116.485 ;
        RECT 30.025 116.145 30.240 116.655 ;
        RECT 30.470 116.145 30.750 116.475 ;
        RECT 30.930 116.145 31.170 116.655 ;
        RECT 26.925 115.415 27.205 115.745 ;
        RECT 27.385 115.415 27.960 115.745 ;
        RECT 28.140 115.415 28.575 115.745 ;
        RECT 28.755 115.415 29.025 115.745 ;
        RECT 26.500 115.055 28.995 115.235 ;
        RECT 25.990 114.285 26.255 115.055 ;
        RECT 26.425 114.105 26.755 114.825 ;
        RECT 26.945 114.645 28.135 114.875 ;
        RECT 26.945 114.285 27.205 114.645 ;
        RECT 27.375 114.105 27.705 114.475 ;
        RECT 27.875 114.285 28.135 114.645 ;
        RECT 28.705 114.285 28.995 115.055 ;
        RECT 29.240 114.895 29.555 115.915 ;
        RECT 29.725 115.245 29.895 115.745 ;
        RECT 30.145 115.415 30.410 115.975 ;
        RECT 30.580 115.245 30.750 116.145 ;
        RECT 31.590 116.085 31.765 116.485 ;
        RECT 31.935 116.275 32.265 116.655 ;
        RECT 32.510 116.155 32.740 116.485 ;
        RECT 30.920 115.415 31.275 115.975 ;
        RECT 31.590 115.915 32.220 116.085 ;
        RECT 32.050 115.745 32.220 115.915 ;
        RECT 29.725 115.075 31.150 115.245 ;
        RECT 29.240 114.275 29.775 114.895 ;
        RECT 29.945 114.105 30.275 114.905 ;
        RECT 30.760 114.900 31.150 115.075 ;
        RECT 31.505 115.065 31.870 115.745 ;
        RECT 32.050 115.415 32.400 115.745 ;
        RECT 32.050 114.895 32.220 115.415 ;
        RECT 31.590 114.725 32.220 114.895 ;
        RECT 32.570 114.865 32.740 116.155 ;
        RECT 32.940 115.045 33.220 116.320 ;
        RECT 33.445 116.315 33.715 116.320 ;
        RECT 33.405 116.145 33.715 116.315 ;
        RECT 34.175 116.275 34.505 116.655 ;
        RECT 34.675 116.400 35.010 116.445 ;
        RECT 33.445 115.045 33.715 116.145 ;
        RECT 33.905 115.045 34.245 116.075 ;
        RECT 34.675 115.935 35.015 116.400 ;
        RECT 34.415 115.415 34.675 115.745 ;
        RECT 34.415 114.865 34.585 115.415 ;
        RECT 34.845 115.245 35.015 115.935 ;
        RECT 31.590 114.275 31.765 114.725 ;
        RECT 32.570 114.695 34.585 114.865 ;
        RECT 31.935 114.105 32.265 114.545 ;
        RECT 32.570 114.275 32.740 114.695 ;
        RECT 32.975 114.105 33.645 114.515 ;
        RECT 33.860 114.275 34.030 114.695 ;
        RECT 34.230 114.105 34.560 114.515 ;
        RECT 34.755 114.275 35.015 115.245 ;
        RECT 35.195 114.285 35.455 116.475 ;
        RECT 35.715 116.285 36.385 116.655 ;
        RECT 36.565 116.105 36.875 116.475 ;
        RECT 35.645 115.905 36.875 116.105 ;
        RECT 35.645 115.235 35.935 115.905 ;
        RECT 37.055 115.725 37.285 116.365 ;
        RECT 37.465 115.925 37.755 116.655 ;
        RECT 37.945 115.930 38.235 116.655 ;
        RECT 38.410 116.255 38.745 116.655 ;
        RECT 38.915 116.085 39.120 116.485 ;
        RECT 39.330 116.175 39.605 116.655 ;
        RECT 39.815 116.155 40.075 116.485 ;
        RECT 38.435 115.915 39.120 116.085 ;
        RECT 36.115 115.415 36.580 115.725 ;
        RECT 36.760 115.415 37.285 115.725 ;
        RECT 37.465 115.415 37.765 115.745 ;
        RECT 35.645 115.015 36.415 115.235 ;
        RECT 35.625 114.105 35.965 114.835 ;
        RECT 36.145 114.285 36.415 115.015 ;
        RECT 36.595 114.995 37.755 115.235 ;
        RECT 36.595 114.285 36.825 114.995 ;
        RECT 36.995 114.105 37.325 114.815 ;
        RECT 37.495 114.285 37.755 114.995 ;
        RECT 37.945 114.105 38.235 115.270 ;
        RECT 38.435 114.885 38.775 115.915 ;
        RECT 38.945 115.245 39.195 115.745 ;
        RECT 39.375 115.415 39.735 115.995 ;
        RECT 39.905 115.245 40.075 116.155 ;
        RECT 41.280 116.025 41.565 116.485 ;
        RECT 41.735 116.195 42.005 116.655 ;
        RECT 41.280 115.855 42.235 116.025 ;
        RECT 38.945 115.075 40.075 115.245 ;
        RECT 41.165 115.125 41.855 115.685 ;
        RECT 38.435 114.710 39.100 114.885 ;
        RECT 38.410 114.105 38.745 114.530 ;
        RECT 38.915 114.305 39.100 114.710 ;
        RECT 39.305 114.105 39.635 114.885 ;
        RECT 39.805 114.305 40.075 115.075 ;
        RECT 42.025 114.955 42.235 115.855 ;
        RECT 41.280 114.735 42.235 114.955 ;
        RECT 42.405 115.685 42.805 116.485 ;
        RECT 42.995 116.025 43.275 116.485 ;
        RECT 43.795 116.195 44.120 116.655 ;
        RECT 42.995 115.855 44.120 116.025 ;
        RECT 44.290 115.915 44.675 116.485 ;
        RECT 43.670 115.745 44.120 115.855 ;
        RECT 42.405 115.125 43.500 115.685 ;
        RECT 43.670 115.415 44.225 115.745 ;
        RECT 41.280 114.275 41.565 114.735 ;
        RECT 41.735 114.105 42.005 114.565 ;
        RECT 42.405 114.275 42.805 115.125 ;
        RECT 43.670 114.955 44.120 115.415 ;
        RECT 44.395 115.245 44.675 115.915 ;
        RECT 44.865 115.845 45.105 116.655 ;
        RECT 45.275 115.845 45.605 116.485 ;
        RECT 45.775 115.845 46.045 116.655 ;
        RECT 46.225 115.905 47.435 116.655 ;
        RECT 47.665 116.195 47.910 116.655 ;
        RECT 44.845 115.415 45.195 115.665 ;
        RECT 45.365 115.245 45.535 115.845 ;
        RECT 45.705 115.415 46.055 115.665 ;
        RECT 46.225 115.365 46.745 115.905 ;
        RECT 42.995 114.735 44.120 114.955 ;
        RECT 42.995 114.275 43.275 114.735 ;
        RECT 43.795 114.105 44.120 114.565 ;
        RECT 44.290 114.275 44.675 115.245 ;
        RECT 44.855 115.075 45.535 115.245 ;
        RECT 44.855 114.290 45.185 115.075 ;
        RECT 45.715 114.105 46.045 115.245 ;
        RECT 46.915 115.195 47.435 115.735 ;
        RECT 47.605 115.415 47.920 116.025 ;
        RECT 48.090 115.665 48.340 116.475 ;
        RECT 48.510 116.130 48.770 116.655 ;
        RECT 48.940 116.005 49.200 116.460 ;
        RECT 49.370 116.175 49.630 116.655 ;
        RECT 49.800 116.005 50.060 116.460 ;
        RECT 50.230 116.175 50.490 116.655 ;
        RECT 50.660 116.005 50.920 116.460 ;
        RECT 51.090 116.175 51.350 116.655 ;
        RECT 51.520 116.005 51.780 116.460 ;
        RECT 51.950 116.175 52.250 116.655 ;
        RECT 48.940 115.835 52.250 116.005 ;
        RECT 48.090 115.415 51.110 115.665 ;
        RECT 46.225 114.105 47.435 115.195 ;
        RECT 47.615 114.105 47.910 115.215 ;
        RECT 48.090 114.280 48.340 115.415 ;
        RECT 51.280 115.245 52.250 115.835 ;
        RECT 52.665 115.905 53.875 116.655 ;
        RECT 54.135 116.105 54.305 116.395 ;
        RECT 54.475 116.275 54.805 116.655 ;
        RECT 54.135 115.935 54.800 116.105 ;
        RECT 52.665 115.365 53.185 115.905 ;
        RECT 48.510 114.105 48.770 115.215 ;
        RECT 48.940 115.005 52.250 115.245 ;
        RECT 53.355 115.195 53.875 115.735 ;
        RECT 48.940 114.280 49.200 115.005 ;
        RECT 49.370 114.105 49.630 114.835 ;
        RECT 49.800 114.280 50.060 115.005 ;
        RECT 50.230 114.105 50.490 114.835 ;
        RECT 50.660 114.280 50.920 115.005 ;
        RECT 51.090 114.105 51.350 114.835 ;
        RECT 51.520 114.280 51.780 115.005 ;
        RECT 51.950 114.105 52.245 114.835 ;
        RECT 52.665 114.105 53.875 115.195 ;
        RECT 54.050 115.115 54.400 115.765 ;
        RECT 54.570 114.945 54.800 115.935 ;
        RECT 54.135 114.775 54.800 114.945 ;
        RECT 54.135 114.275 54.305 114.775 ;
        RECT 54.475 114.105 54.805 114.605 ;
        RECT 54.975 114.275 55.160 116.395 ;
        RECT 55.415 116.195 55.665 116.655 ;
        RECT 55.835 116.205 56.170 116.375 ;
        RECT 56.365 116.205 57.040 116.375 ;
        RECT 55.835 116.065 56.005 116.205 ;
        RECT 55.330 115.075 55.610 116.025 ;
        RECT 55.780 115.935 56.005 116.065 ;
        RECT 55.780 114.830 55.950 115.935 ;
        RECT 56.175 115.785 56.700 116.005 ;
        RECT 56.120 115.020 56.360 115.615 ;
        RECT 56.530 115.085 56.700 115.785 ;
        RECT 56.870 115.425 57.040 116.205 ;
        RECT 57.360 116.155 57.730 116.655 ;
        RECT 57.910 116.205 58.315 116.375 ;
        RECT 58.485 116.205 59.270 116.375 ;
        RECT 57.910 115.975 58.080 116.205 ;
        RECT 57.250 115.675 58.080 115.975 ;
        RECT 58.465 115.705 58.930 116.035 ;
        RECT 57.250 115.645 57.450 115.675 ;
        RECT 57.570 115.425 57.740 115.495 ;
        RECT 56.870 115.255 57.740 115.425 ;
        RECT 57.230 115.165 57.740 115.255 ;
        RECT 55.780 114.700 56.085 114.830 ;
        RECT 56.530 114.720 57.060 115.085 ;
        RECT 55.400 114.105 55.665 114.565 ;
        RECT 55.835 114.275 56.085 114.700 ;
        RECT 57.230 114.550 57.400 115.165 ;
        RECT 56.295 114.380 57.400 114.550 ;
        RECT 57.570 114.105 57.740 114.905 ;
        RECT 57.910 114.605 58.080 115.675 ;
        RECT 58.250 114.775 58.440 115.495 ;
        RECT 58.610 114.745 58.930 115.705 ;
        RECT 59.100 115.745 59.270 116.205 ;
        RECT 59.545 116.125 59.755 116.655 ;
        RECT 60.015 115.915 60.345 116.440 ;
        RECT 60.515 116.045 60.685 116.655 ;
        RECT 60.855 116.000 61.185 116.435 ;
        RECT 61.420 116.085 61.675 116.435 ;
        RECT 61.845 116.255 62.175 116.655 ;
        RECT 62.345 116.085 62.515 116.435 ;
        RECT 62.685 116.255 63.065 116.655 ;
        RECT 60.855 115.915 61.235 116.000 ;
        RECT 61.420 115.915 63.085 116.085 ;
        RECT 63.255 115.980 63.530 116.325 ;
        RECT 60.145 115.745 60.345 115.915 ;
        RECT 61.010 115.875 61.235 115.915 ;
        RECT 59.100 115.415 59.975 115.745 ;
        RECT 60.145 115.415 60.895 115.745 ;
        RECT 57.910 114.275 58.160 114.605 ;
        RECT 59.100 114.575 59.270 115.415 ;
        RECT 60.145 115.210 60.335 115.415 ;
        RECT 61.065 115.295 61.235 115.875 ;
        RECT 62.915 115.745 63.085 115.915 ;
        RECT 61.405 115.415 61.750 115.745 ;
        RECT 61.920 115.415 62.745 115.745 ;
        RECT 62.915 115.415 63.190 115.745 ;
        RECT 61.020 115.245 61.235 115.295 ;
        RECT 59.440 114.835 60.335 115.210 ;
        RECT 60.845 115.165 61.235 115.245 ;
        RECT 58.385 114.405 59.270 114.575 ;
        RECT 59.450 114.105 59.765 114.605 ;
        RECT 59.995 114.275 60.335 114.835 ;
        RECT 60.505 114.105 60.675 115.115 ;
        RECT 60.845 114.320 61.175 115.165 ;
        RECT 61.425 114.955 61.750 115.245 ;
        RECT 61.920 115.125 62.115 115.415 ;
        RECT 62.915 115.245 63.085 115.415 ;
        RECT 63.360 115.245 63.530 115.980 ;
        RECT 63.705 115.930 63.995 116.655 ;
        RECT 64.325 116.095 64.655 116.485 ;
        RECT 64.825 116.265 66.010 116.435 ;
        RECT 66.270 116.185 66.440 116.655 ;
        RECT 64.325 115.915 64.835 116.095 ;
        RECT 64.165 115.455 64.495 115.745 ;
        RECT 64.665 115.285 64.835 115.915 ;
        RECT 65.240 116.005 65.625 116.095 ;
        RECT 66.610 116.005 66.940 116.470 ;
        RECT 65.240 115.835 66.940 116.005 ;
        RECT 67.110 115.835 67.280 116.655 ;
        RECT 67.450 115.835 68.135 116.475 ;
        RECT 68.395 116.105 68.565 116.395 ;
        RECT 68.735 116.275 69.065 116.655 ;
        RECT 68.395 115.935 69.060 116.105 ;
        RECT 65.005 115.455 65.335 115.665 ;
        RECT 65.515 115.415 65.895 115.665 ;
        RECT 62.425 115.075 63.085 115.245 ;
        RECT 62.425 114.955 62.595 115.075 ;
        RECT 61.425 114.785 62.595 114.955 ;
        RECT 61.405 114.325 62.595 114.615 ;
        RECT 62.765 114.105 63.045 114.905 ;
        RECT 63.255 114.275 63.530 115.245 ;
        RECT 63.705 114.105 63.995 115.270 ;
        RECT 64.320 115.115 65.405 115.285 ;
        RECT 64.320 114.275 64.620 115.115 ;
        RECT 64.815 114.105 65.065 114.945 ;
        RECT 65.235 114.865 65.405 115.115 ;
        RECT 65.575 115.035 65.895 115.415 ;
        RECT 66.085 115.455 66.570 115.665 ;
        RECT 66.760 115.455 67.210 115.665 ;
        RECT 67.380 115.455 67.715 115.665 ;
        RECT 66.085 115.295 66.460 115.455 ;
        RECT 66.065 115.125 66.460 115.295 ;
        RECT 67.380 115.285 67.550 115.455 ;
        RECT 66.085 115.035 66.460 115.125 ;
        RECT 66.630 115.115 67.550 115.285 ;
        RECT 66.630 114.865 66.800 115.115 ;
        RECT 65.235 114.695 66.800 114.865 ;
        RECT 65.655 114.275 66.460 114.695 ;
        RECT 66.970 114.105 67.300 114.945 ;
        RECT 67.885 114.865 68.135 115.835 ;
        RECT 68.310 115.115 68.660 115.765 ;
        RECT 68.830 114.945 69.060 115.935 ;
        RECT 67.470 114.275 68.135 114.865 ;
        RECT 68.395 114.775 69.060 114.945 ;
        RECT 68.395 114.275 68.565 114.775 ;
        RECT 68.735 114.105 69.065 114.605 ;
        RECT 69.235 114.275 69.420 116.395 ;
        RECT 69.675 116.195 69.925 116.655 ;
        RECT 70.095 116.205 70.430 116.375 ;
        RECT 70.625 116.205 71.300 116.375 ;
        RECT 70.095 116.065 70.265 116.205 ;
        RECT 69.590 115.075 69.870 116.025 ;
        RECT 70.040 115.935 70.265 116.065 ;
        RECT 70.040 114.830 70.210 115.935 ;
        RECT 70.435 115.785 70.960 116.005 ;
        RECT 70.380 115.020 70.620 115.615 ;
        RECT 70.790 115.085 70.960 115.785 ;
        RECT 71.130 115.425 71.300 116.205 ;
        RECT 71.620 116.155 71.990 116.655 ;
        RECT 72.170 116.205 72.575 116.375 ;
        RECT 72.745 116.205 73.530 116.375 ;
        RECT 72.170 115.975 72.340 116.205 ;
        RECT 71.510 115.675 72.340 115.975 ;
        RECT 72.725 115.705 73.190 116.035 ;
        RECT 71.510 115.645 71.710 115.675 ;
        RECT 71.830 115.425 72.000 115.495 ;
        RECT 71.130 115.255 72.000 115.425 ;
        RECT 71.490 115.165 72.000 115.255 ;
        RECT 70.040 114.700 70.345 114.830 ;
        RECT 70.790 114.720 71.320 115.085 ;
        RECT 69.660 114.105 69.925 114.565 ;
        RECT 70.095 114.275 70.345 114.700 ;
        RECT 71.490 114.550 71.660 115.165 ;
        RECT 70.555 114.380 71.660 114.550 ;
        RECT 71.830 114.105 72.000 114.905 ;
        RECT 72.170 114.605 72.340 115.675 ;
        RECT 72.510 114.775 72.700 115.495 ;
        RECT 72.870 114.745 73.190 115.705 ;
        RECT 73.360 115.745 73.530 116.205 ;
        RECT 73.805 116.125 74.015 116.655 ;
        RECT 74.275 115.915 74.605 116.440 ;
        RECT 74.775 116.045 74.945 116.655 ;
        RECT 75.115 116.000 75.445 116.435 ;
        RECT 75.115 115.915 75.495 116.000 ;
        RECT 74.405 115.745 74.605 115.915 ;
        RECT 75.270 115.875 75.495 115.915 ;
        RECT 73.360 115.415 74.235 115.745 ;
        RECT 74.405 115.415 75.155 115.745 ;
        RECT 72.170 114.275 72.420 114.605 ;
        RECT 73.360 114.575 73.530 115.415 ;
        RECT 74.405 115.210 74.595 115.415 ;
        RECT 75.325 115.295 75.495 115.875 ;
        RECT 75.280 115.245 75.495 115.295 ;
        RECT 73.700 114.835 74.595 115.210 ;
        RECT 75.105 115.165 75.495 115.245 ;
        RECT 75.665 115.915 76.050 116.485 ;
        RECT 76.220 116.195 76.545 116.655 ;
        RECT 77.065 116.025 77.345 116.485 ;
        RECT 75.665 115.245 75.945 115.915 ;
        RECT 76.220 115.855 77.345 116.025 ;
        RECT 76.220 115.745 76.670 115.855 ;
        RECT 76.115 115.415 76.670 115.745 ;
        RECT 77.535 115.685 77.935 116.485 ;
        RECT 78.335 116.195 78.605 116.655 ;
        RECT 78.775 116.025 79.060 116.485 ;
        RECT 72.645 114.405 73.530 114.575 ;
        RECT 73.710 114.105 74.025 114.605 ;
        RECT 74.255 114.275 74.595 114.835 ;
        RECT 74.765 114.105 74.935 115.115 ;
        RECT 75.105 114.320 75.435 115.165 ;
        RECT 75.665 114.275 76.050 115.245 ;
        RECT 76.220 114.955 76.670 115.415 ;
        RECT 76.840 115.125 77.935 115.685 ;
        RECT 76.220 114.735 77.345 114.955 ;
        RECT 76.220 114.105 76.545 114.565 ;
        RECT 77.065 114.275 77.345 114.735 ;
        RECT 77.535 114.275 77.935 115.125 ;
        RECT 78.105 115.855 79.060 116.025 ;
        RECT 79.345 115.855 79.685 116.485 ;
        RECT 79.855 115.855 80.105 116.655 ;
        RECT 80.295 116.005 80.625 116.485 ;
        RECT 80.795 116.195 81.020 116.655 ;
        RECT 81.190 116.005 81.520 116.485 ;
        RECT 78.105 114.955 78.315 115.855 ;
        RECT 78.485 115.125 79.175 115.685 ;
        RECT 79.345 115.245 79.520 115.855 ;
        RECT 80.295 115.835 81.520 116.005 ;
        RECT 82.150 115.875 82.650 116.485 ;
        RECT 83.115 116.105 83.285 116.485 ;
        RECT 83.465 116.275 83.795 116.655 ;
        RECT 83.115 115.935 83.780 116.105 ;
        RECT 83.975 115.980 84.235 116.485 ;
        RECT 79.690 115.495 80.385 115.665 ;
        RECT 80.215 115.245 80.385 115.495 ;
        RECT 80.560 115.465 80.980 115.665 ;
        RECT 81.150 115.465 81.480 115.665 ;
        RECT 81.650 115.465 81.980 115.665 ;
        RECT 82.150 115.245 82.320 115.875 ;
        RECT 82.505 115.415 82.855 115.665 ;
        RECT 83.045 115.385 83.375 115.755 ;
        RECT 83.610 115.680 83.780 115.935 ;
        RECT 83.610 115.350 83.895 115.680 ;
        RECT 78.105 114.735 79.060 114.955 ;
        RECT 78.335 114.105 78.605 114.565 ;
        RECT 78.775 114.275 79.060 114.735 ;
        RECT 79.345 114.275 79.685 115.245 ;
        RECT 79.855 114.105 80.025 115.245 ;
        RECT 80.215 115.075 82.650 115.245 ;
        RECT 83.610 115.205 83.780 115.350 ;
        RECT 80.295 114.105 80.545 114.905 ;
        RECT 81.190 114.275 81.520 115.075 ;
        RECT 81.820 114.105 82.150 114.905 ;
        RECT 82.320 114.275 82.650 115.075 ;
        RECT 83.115 115.035 83.780 115.205 ;
        RECT 84.065 115.180 84.235 115.980 ;
        RECT 83.115 114.275 83.285 115.035 ;
        RECT 83.465 114.105 83.795 114.865 ;
        RECT 83.965 114.275 84.235 115.180 ;
        RECT 84.440 115.915 85.055 116.485 ;
        RECT 85.225 116.145 85.440 116.655 ;
        RECT 85.670 116.145 85.950 116.475 ;
        RECT 86.130 116.145 86.370 116.655 ;
        RECT 84.440 114.895 84.755 115.915 ;
        RECT 84.925 115.245 85.095 115.745 ;
        RECT 85.345 115.415 85.610 115.975 ;
        RECT 85.780 115.245 85.950 116.145 ;
        RECT 86.795 116.105 86.965 116.485 ;
        RECT 87.180 116.275 87.510 116.655 ;
        RECT 86.120 115.415 86.475 115.975 ;
        RECT 86.795 115.935 87.510 116.105 ;
        RECT 86.705 115.385 87.060 115.755 ;
        RECT 87.340 115.745 87.510 115.935 ;
        RECT 87.680 115.910 87.935 116.485 ;
        RECT 87.340 115.415 87.595 115.745 ;
        RECT 84.925 115.075 86.350 115.245 ;
        RECT 87.340 115.205 87.510 115.415 ;
        RECT 84.440 114.275 84.975 114.895 ;
        RECT 85.145 114.105 85.475 114.905 ;
        RECT 85.960 114.900 86.350 115.075 ;
        RECT 86.795 115.035 87.510 115.205 ;
        RECT 87.765 115.180 87.935 115.910 ;
        RECT 88.110 115.815 88.370 116.655 ;
        RECT 88.545 115.905 89.755 116.655 ;
        RECT 86.795 114.275 86.965 115.035 ;
        RECT 87.180 114.105 87.510 114.865 ;
        RECT 87.680 114.275 87.935 115.180 ;
        RECT 88.110 114.105 88.370 115.255 ;
        RECT 88.545 115.195 89.065 115.735 ;
        RECT 89.235 115.365 89.755 115.905 ;
        RECT 100.090 116.640 106.320 116.800 ;
        RECT 88.545 114.105 89.755 115.195 ;
        RECT 100.090 114.380 100.760 116.640 ;
        RECT 101.430 116.070 105.470 116.240 ;
        RECT 101.090 115.010 101.260 116.010 ;
        RECT 105.640 115.010 105.810 116.010 ;
        RECT 101.430 114.780 105.470 114.950 ;
        RECT 106.150 114.380 106.320 116.640 ;
        RECT 100.090 114.210 106.320 114.380 ;
        RECT 12.100 113.935 89.840 114.105 ;
        RECT 12.185 112.845 13.395 113.935 ;
        RECT 12.185 112.135 12.705 112.675 ;
        RECT 12.875 112.305 13.395 112.845 ;
        RECT 12.185 111.385 13.395 112.135 ;
        RECT 14.025 111.555 14.285 113.765 ;
        RECT 14.455 113.555 14.785 113.935 ;
        RECT 15.210 113.385 15.380 113.765 ;
        RECT 15.640 113.555 15.970 113.935 ;
        RECT 16.165 113.385 16.335 113.765 ;
        RECT 16.545 113.555 16.875 113.935 ;
        RECT 17.125 113.385 17.315 113.765 ;
        RECT 17.555 113.555 17.885 113.935 ;
        RECT 18.195 113.435 18.455 113.765 ;
        RECT 14.455 113.215 16.405 113.385 ;
        RECT 14.455 112.295 14.625 113.215 ;
        RECT 14.995 112.625 15.190 112.935 ;
        RECT 15.460 112.625 15.645 112.935 ;
        RECT 14.935 112.295 15.190 112.625 ;
        RECT 15.415 112.295 15.645 112.625 ;
        RECT 14.455 111.385 14.785 111.765 ;
        RECT 14.995 111.720 15.190 112.295 ;
        RECT 15.460 111.715 15.645 112.295 ;
        RECT 15.895 111.725 16.065 112.625 ;
        RECT 16.235 112.225 16.405 113.215 ;
        RECT 16.575 113.215 17.315 113.385 ;
        RECT 16.575 112.705 16.745 113.215 ;
        RECT 16.915 112.875 17.495 113.045 ;
        RECT 17.765 112.925 18.115 113.255 ;
        RECT 17.325 112.755 17.495 112.875 ;
        RECT 18.285 112.755 18.455 113.435 ;
        RECT 16.575 112.535 17.145 112.705 ;
        RECT 17.325 112.585 18.455 112.755 ;
        RECT 16.235 111.895 16.785 112.225 ;
        RECT 16.975 112.055 17.145 112.535 ;
        RECT 17.315 112.245 17.935 112.415 ;
        RECT 17.725 112.065 17.935 112.245 ;
        RECT 16.975 111.725 17.375 112.055 ;
        RECT 18.285 111.885 18.455 112.585 ;
        RECT 15.895 111.555 17.375 111.725 ;
        RECT 17.555 111.385 17.885 111.765 ;
        RECT 18.195 111.555 18.455 111.885 ;
        RECT 18.625 112.795 18.885 113.765 ;
        RECT 19.080 113.525 19.410 113.935 ;
        RECT 19.610 113.345 19.780 113.765 ;
        RECT 19.995 113.525 20.665 113.935 ;
        RECT 20.900 113.345 21.070 113.765 ;
        RECT 21.375 113.495 21.705 113.935 ;
        RECT 19.055 113.175 21.070 113.345 ;
        RECT 21.875 113.315 22.050 113.765 ;
        RECT 18.625 112.105 18.795 112.795 ;
        RECT 19.055 112.625 19.225 113.175 ;
        RECT 18.965 112.295 19.225 112.625 ;
        RECT 18.625 111.640 18.965 112.105 ;
        RECT 19.395 111.965 19.735 112.995 ;
        RECT 19.925 112.915 20.195 112.995 ;
        RECT 19.925 112.745 20.235 112.915 ;
        RECT 18.630 111.595 18.965 111.640 ;
        RECT 19.135 111.385 19.465 111.765 ;
        RECT 19.925 111.720 20.195 112.745 ;
        RECT 20.420 111.720 20.700 112.995 ;
        RECT 20.900 111.885 21.070 113.175 ;
        RECT 21.420 113.145 22.050 113.315 ;
        RECT 21.420 112.625 21.590 113.145 ;
        RECT 22.800 113.135 23.050 113.935 ;
        RECT 23.220 113.305 23.550 113.765 ;
        RECT 23.720 113.475 23.935 113.935 ;
        RECT 23.220 113.135 24.390 113.305 ;
        RECT 21.240 112.295 21.590 112.625 ;
        RECT 21.770 112.295 22.135 112.975 ;
        RECT 22.310 112.965 22.590 113.125 ;
        RECT 22.310 112.795 23.645 112.965 ;
        RECT 23.475 112.625 23.645 112.795 ;
        RECT 22.310 112.375 22.660 112.615 ;
        RECT 22.830 112.375 23.305 112.615 ;
        RECT 23.475 112.375 23.850 112.625 ;
        RECT 21.420 112.125 21.590 112.295 ;
        RECT 23.475 112.205 23.645 112.375 ;
        RECT 21.420 111.955 22.050 112.125 ;
        RECT 20.900 111.555 21.130 111.885 ;
        RECT 21.375 111.385 21.705 111.765 ;
        RECT 21.875 111.555 22.050 111.955 ;
        RECT 22.310 112.035 23.645 112.205 ;
        RECT 22.310 111.825 22.580 112.035 ;
        RECT 24.020 111.845 24.390 113.135 ;
        RECT 25.065 112.770 25.355 113.935 ;
        RECT 25.525 113.095 25.785 113.765 ;
        RECT 25.955 113.535 26.285 113.935 ;
        RECT 27.155 113.535 27.555 113.935 ;
        RECT 27.845 113.355 28.175 113.590 ;
        RECT 26.095 113.185 28.175 113.355 ;
        RECT 25.525 112.125 25.700 113.095 ;
        RECT 26.095 112.915 26.265 113.185 ;
        RECT 25.870 112.745 26.265 112.915 ;
        RECT 26.435 112.795 27.450 113.015 ;
        RECT 25.870 112.295 26.040 112.745 ;
        RECT 27.175 112.655 27.450 112.795 ;
        RECT 27.620 112.795 28.175 113.185 ;
        RECT 26.210 112.375 26.660 112.575 ;
        RECT 26.830 112.205 27.005 112.400 ;
        RECT 22.800 111.385 23.130 111.845 ;
        RECT 23.640 111.555 24.390 111.845 ;
        RECT 25.065 111.385 25.355 112.110 ;
        RECT 25.525 111.555 25.865 112.125 ;
        RECT 26.060 111.385 26.230 112.050 ;
        RECT 26.510 112.035 27.005 112.205 ;
        RECT 26.510 111.895 26.730 112.035 ;
        RECT 26.505 111.725 26.730 111.895 ;
        RECT 27.175 111.865 27.345 112.655 ;
        RECT 27.620 112.545 27.790 112.795 ;
        RECT 28.345 112.625 28.520 113.725 ;
        RECT 28.690 113.115 29.035 113.935 ;
        RECT 29.205 113.340 29.640 113.765 ;
        RECT 29.810 113.510 30.195 113.935 ;
        RECT 29.205 113.170 30.195 113.340 ;
        RECT 27.595 112.375 27.790 112.545 ;
        RECT 27.960 112.375 28.520 112.625 ;
        RECT 28.690 112.375 29.035 112.945 ;
        RECT 27.595 111.990 27.765 112.375 ;
        RECT 29.205 112.295 29.690 113.000 ;
        RECT 29.860 112.625 30.195 113.170 ;
        RECT 30.365 112.975 30.790 113.765 ;
        RECT 30.960 113.340 31.235 113.765 ;
        RECT 31.405 113.510 31.790 113.935 ;
        RECT 30.960 113.145 31.790 113.340 ;
        RECT 30.365 112.795 31.270 112.975 ;
        RECT 29.860 112.295 30.270 112.625 ;
        RECT 30.440 112.295 31.270 112.795 ;
        RECT 31.440 112.625 31.790 113.145 ;
        RECT 31.960 112.975 32.205 113.765 ;
        RECT 32.395 113.340 32.650 113.765 ;
        RECT 32.820 113.510 33.205 113.935 ;
        RECT 32.395 113.145 33.205 113.340 ;
        RECT 31.960 112.795 32.685 112.975 ;
        RECT 31.440 112.295 31.865 112.625 ;
        RECT 32.035 112.295 32.685 112.795 ;
        RECT 32.855 112.625 33.205 113.145 ;
        RECT 33.375 112.795 33.635 113.765 ;
        RECT 34.350 113.315 34.525 113.765 ;
        RECT 34.695 113.495 35.025 113.935 ;
        RECT 35.330 113.345 35.500 113.765 ;
        RECT 35.735 113.525 36.405 113.935 ;
        RECT 36.620 113.345 36.790 113.765 ;
        RECT 36.990 113.525 37.320 113.935 ;
        RECT 34.350 113.145 34.980 113.315 ;
        RECT 32.855 112.295 33.280 112.625 ;
        RECT 26.510 111.680 26.730 111.725 ;
        RECT 26.900 111.695 27.345 111.865 ;
        RECT 27.515 111.620 27.765 111.990 ;
        RECT 27.935 112.025 29.035 112.205 ;
        RECT 29.860 112.125 30.195 112.295 ;
        RECT 30.440 112.125 30.790 112.295 ;
        RECT 31.440 112.125 31.790 112.295 ;
        RECT 32.035 112.125 32.205 112.295 ;
        RECT 32.855 112.125 33.205 112.295 ;
        RECT 33.450 112.125 33.635 112.795 ;
        RECT 34.265 112.295 34.630 112.975 ;
        RECT 34.810 112.625 34.980 113.145 ;
        RECT 35.330 113.175 37.345 113.345 ;
        RECT 34.810 112.295 35.160 112.625 ;
        RECT 34.810 112.125 34.980 112.295 ;
        RECT 27.935 111.620 28.185 112.025 ;
        RECT 28.355 111.385 28.525 111.855 ;
        RECT 28.695 111.620 29.035 112.025 ;
        RECT 29.205 111.955 30.195 112.125 ;
        RECT 29.205 111.555 29.640 111.955 ;
        RECT 29.810 111.385 30.195 111.785 ;
        RECT 30.365 111.555 30.790 112.125 ;
        RECT 30.980 111.955 31.790 112.125 ;
        RECT 30.980 111.555 31.235 111.955 ;
        RECT 31.405 111.385 31.790 111.785 ;
        RECT 31.960 111.555 32.205 112.125 ;
        RECT 32.395 111.955 33.205 112.125 ;
        RECT 32.395 111.555 32.650 111.955 ;
        RECT 32.820 111.385 33.205 111.785 ;
        RECT 33.375 111.555 33.635 112.125 ;
        RECT 34.350 111.955 34.980 112.125 ;
        RECT 34.350 111.555 34.525 111.955 ;
        RECT 35.330 111.885 35.500 113.175 ;
        RECT 34.695 111.385 35.025 111.765 ;
        RECT 35.270 111.555 35.500 111.885 ;
        RECT 35.700 111.720 35.980 112.995 ;
        RECT 36.205 112.235 36.475 112.995 ;
        RECT 36.165 112.065 36.475 112.235 ;
        RECT 36.205 111.720 36.475 112.065 ;
        RECT 36.665 111.965 37.005 112.995 ;
        RECT 37.175 112.625 37.345 113.175 ;
        RECT 37.515 112.795 37.775 113.765 ;
        RECT 37.965 113.425 38.265 113.935 ;
        RECT 38.435 113.425 38.815 113.595 ;
        RECT 39.395 113.425 40.025 113.935 ;
        RECT 38.435 113.255 38.605 113.425 ;
        RECT 40.195 113.255 40.525 113.765 ;
        RECT 40.695 113.425 40.995 113.935 ;
        RECT 41.255 113.265 41.425 113.765 ;
        RECT 41.595 113.435 41.925 113.935 ;
        RECT 37.175 112.295 37.435 112.625 ;
        RECT 37.605 112.105 37.775 112.795 ;
        RECT 36.935 111.385 37.265 111.765 ;
        RECT 37.435 111.640 37.775 112.105 ;
        RECT 37.945 113.055 38.605 113.255 ;
        RECT 38.775 113.085 40.995 113.255 ;
        RECT 41.255 113.095 41.920 113.265 ;
        RECT 37.945 112.125 38.115 113.055 ;
        RECT 38.775 112.885 38.945 113.085 ;
        RECT 38.285 112.715 38.945 112.885 ;
        RECT 39.115 112.745 40.655 112.915 ;
        RECT 38.285 112.295 38.455 112.715 ;
        RECT 39.115 112.545 39.285 112.745 ;
        RECT 38.685 112.375 39.285 112.545 ;
        RECT 39.455 112.375 40.150 112.575 ;
        RECT 40.410 112.295 40.655 112.745 ;
        RECT 38.775 112.125 39.685 112.205 ;
        RECT 37.945 111.645 38.265 112.125 ;
        RECT 38.435 112.035 39.685 112.125 ;
        RECT 38.435 111.955 38.945 112.035 ;
        RECT 37.435 111.595 37.770 111.640 ;
        RECT 38.435 111.555 38.665 111.955 ;
        RECT 38.835 111.385 39.185 111.775 ;
        RECT 39.355 111.555 39.685 112.035 ;
        RECT 39.855 111.385 40.025 112.205 ;
        RECT 40.825 112.125 40.995 113.085 ;
        RECT 41.170 112.275 41.520 112.925 ;
        RECT 40.530 111.580 40.995 112.125 ;
        RECT 41.690 112.105 41.920 113.095 ;
        RECT 41.255 111.935 41.920 112.105 ;
        RECT 41.255 111.645 41.425 111.935 ;
        RECT 41.595 111.385 41.925 111.765 ;
        RECT 42.095 111.645 42.280 113.765 ;
        RECT 42.520 113.475 42.785 113.935 ;
        RECT 42.955 113.340 43.205 113.765 ;
        RECT 43.415 113.490 44.520 113.660 ;
        RECT 42.900 113.210 43.205 113.340 ;
        RECT 42.450 112.015 42.730 112.965 ;
        RECT 42.900 112.105 43.070 113.210 ;
        RECT 43.240 112.425 43.480 113.020 ;
        RECT 43.650 112.955 44.180 113.320 ;
        RECT 43.650 112.255 43.820 112.955 ;
        RECT 44.350 112.875 44.520 113.490 ;
        RECT 44.690 113.135 44.860 113.935 ;
        RECT 45.030 113.435 45.280 113.765 ;
        RECT 45.505 113.465 46.390 113.635 ;
        RECT 44.350 112.785 44.860 112.875 ;
        RECT 42.900 111.975 43.125 112.105 ;
        RECT 43.295 112.035 43.820 112.255 ;
        RECT 43.990 112.615 44.860 112.785 ;
        RECT 42.535 111.385 42.785 111.845 ;
        RECT 42.955 111.835 43.125 111.975 ;
        RECT 43.990 111.835 44.160 112.615 ;
        RECT 44.690 112.545 44.860 112.615 ;
        RECT 44.370 112.365 44.570 112.395 ;
        RECT 45.030 112.365 45.200 113.435 ;
        RECT 45.370 112.545 45.560 113.265 ;
        RECT 44.370 112.065 45.200 112.365 ;
        RECT 45.730 112.335 46.050 113.295 ;
        RECT 42.955 111.665 43.290 111.835 ;
        RECT 43.485 111.665 44.160 111.835 ;
        RECT 44.480 111.385 44.850 111.885 ;
        RECT 45.030 111.835 45.200 112.065 ;
        RECT 45.585 112.005 46.050 112.335 ;
        RECT 46.220 112.625 46.390 113.465 ;
        RECT 46.570 113.435 46.885 113.935 ;
        RECT 47.115 113.205 47.455 113.765 ;
        RECT 46.560 112.830 47.455 113.205 ;
        RECT 47.625 112.925 47.795 113.935 ;
        RECT 47.265 112.625 47.455 112.830 ;
        RECT 47.965 112.875 48.295 113.720 ;
        RECT 47.965 112.795 48.355 112.875 ;
        RECT 48.525 112.845 50.195 113.935 ;
        RECT 48.140 112.745 48.355 112.795 ;
        RECT 46.220 112.295 47.095 112.625 ;
        RECT 47.265 112.295 48.015 112.625 ;
        RECT 46.220 111.835 46.390 112.295 ;
        RECT 47.265 112.125 47.465 112.295 ;
        RECT 48.185 112.165 48.355 112.745 ;
        RECT 48.130 112.125 48.355 112.165 ;
        RECT 45.030 111.665 45.435 111.835 ;
        RECT 45.605 111.665 46.390 111.835 ;
        RECT 46.665 111.385 46.875 111.915 ;
        RECT 47.135 111.600 47.465 112.125 ;
        RECT 47.975 112.040 48.355 112.125 ;
        RECT 48.525 112.155 49.275 112.675 ;
        RECT 49.445 112.325 50.195 112.845 ;
        RECT 50.825 112.770 51.115 113.935 ;
        RECT 51.330 112.795 51.625 113.935 ;
        RECT 51.885 112.965 52.215 113.765 ;
        RECT 52.385 113.135 52.555 113.935 ;
        RECT 52.725 112.965 53.055 113.765 ;
        RECT 53.225 113.135 53.395 113.935 ;
        RECT 53.565 112.985 53.895 113.765 ;
        RECT 54.065 113.475 54.235 113.935 ;
        RECT 55.425 113.135 55.865 113.765 ;
        RECT 53.565 112.965 54.335 112.985 ;
        RECT 51.885 112.795 54.335 112.965 ;
        RECT 51.305 112.375 53.815 112.625 ;
        RECT 53.985 112.205 54.335 112.795 ;
        RECT 47.635 111.385 47.805 111.995 ;
        RECT 47.975 111.605 48.305 112.040 ;
        RECT 48.525 111.385 50.195 112.155 ;
        RECT 50.825 111.385 51.115 112.110 ;
        RECT 51.965 112.025 54.335 112.205 ;
        RECT 55.425 112.125 55.735 113.135 ;
        RECT 56.040 113.085 56.355 113.935 ;
        RECT 56.525 113.595 57.955 113.765 ;
        RECT 56.525 112.915 56.695 113.595 ;
        RECT 55.905 112.745 56.695 112.915 ;
        RECT 55.905 112.295 56.075 112.745 ;
        RECT 56.865 112.625 57.065 113.425 ;
        RECT 56.245 112.295 56.635 112.575 ;
        RECT 56.820 112.295 57.065 112.625 ;
        RECT 57.265 112.295 57.515 113.425 ;
        RECT 57.705 112.965 57.955 113.595 ;
        RECT 58.135 113.135 58.465 113.935 ;
        RECT 58.655 112.965 58.985 113.750 ;
        RECT 57.705 112.795 58.475 112.965 ;
        RECT 58.655 112.795 59.335 112.965 ;
        RECT 59.515 112.795 59.845 113.935 ;
        RECT 60.025 112.795 60.285 113.935 ;
        RECT 57.730 112.295 58.135 112.625 ;
        RECT 58.305 112.125 58.475 112.795 ;
        RECT 58.645 112.375 58.995 112.625 ;
        RECT 59.165 112.195 59.335 112.795 ;
        RECT 60.455 112.785 60.785 113.765 ;
        RECT 60.955 112.795 61.235 113.935 ;
        RECT 61.520 113.305 61.805 113.765 ;
        RECT 61.975 113.475 62.245 113.935 ;
        RECT 61.520 113.085 62.475 113.305 ;
        RECT 59.505 112.375 59.855 112.625 ;
        RECT 60.045 112.375 60.380 112.625 ;
        RECT 51.330 111.385 51.595 111.845 ;
        RECT 51.965 111.555 52.135 112.025 ;
        RECT 52.385 111.385 52.555 111.845 ;
        RECT 52.805 111.555 52.975 112.025 ;
        RECT 53.225 111.385 53.395 111.845 ;
        RECT 53.645 111.555 53.815 112.025 ;
        RECT 53.985 111.385 54.235 111.850 ;
        RECT 55.425 111.565 55.865 112.125 ;
        RECT 56.035 111.385 56.485 112.125 ;
        RECT 56.655 111.955 57.815 112.125 ;
        RECT 56.655 111.555 56.825 111.955 ;
        RECT 56.995 111.385 57.415 111.785 ;
        RECT 57.585 111.555 57.815 111.955 ;
        RECT 57.985 111.555 58.475 112.125 ;
        RECT 58.665 111.385 58.905 112.195 ;
        RECT 59.075 111.555 59.405 112.195 ;
        RECT 59.575 111.385 59.845 112.195 ;
        RECT 60.550 112.185 60.720 112.785 ;
        RECT 60.890 112.355 61.225 112.625 ;
        RECT 61.405 112.355 62.095 112.915 ;
        RECT 62.265 112.185 62.475 113.085 ;
        RECT 60.025 111.555 60.720 112.185 ;
        RECT 60.925 111.385 61.235 112.185 ;
        RECT 61.520 112.015 62.475 112.185 ;
        RECT 62.645 112.915 63.045 113.765 ;
        RECT 63.235 113.305 63.515 113.765 ;
        RECT 64.035 113.475 64.360 113.935 ;
        RECT 63.235 113.085 64.360 113.305 ;
        RECT 62.645 112.355 63.740 112.915 ;
        RECT 63.910 112.625 64.360 113.085 ;
        RECT 64.530 112.795 64.915 113.765 ;
        RECT 65.290 112.965 65.620 113.765 ;
        RECT 65.790 113.135 66.120 113.935 ;
        RECT 66.420 112.965 66.750 113.765 ;
        RECT 67.395 113.135 67.645 113.935 ;
        RECT 65.290 112.795 67.725 112.965 ;
        RECT 67.915 112.795 68.085 113.935 ;
        RECT 68.255 112.795 68.595 113.765 ;
        RECT 68.765 112.795 69.045 113.935 ;
        RECT 61.520 111.555 61.805 112.015 ;
        RECT 61.975 111.385 62.245 111.845 ;
        RECT 62.645 111.555 63.045 112.355 ;
        RECT 63.910 112.295 64.465 112.625 ;
        RECT 63.910 112.185 64.360 112.295 ;
        RECT 63.235 112.015 64.360 112.185 ;
        RECT 64.635 112.125 64.915 112.795 ;
        RECT 65.085 112.375 65.435 112.625 ;
        RECT 65.620 112.165 65.790 112.795 ;
        RECT 65.960 112.375 66.290 112.575 ;
        RECT 66.460 112.375 66.790 112.575 ;
        RECT 66.960 112.375 67.380 112.575 ;
        RECT 67.555 112.545 67.725 112.795 ;
        RECT 67.555 112.375 68.250 112.545 ;
        RECT 63.235 111.555 63.515 112.015 ;
        RECT 64.035 111.385 64.360 111.845 ;
        RECT 64.530 111.555 64.915 112.125 ;
        RECT 65.290 111.555 65.790 112.165 ;
        RECT 66.420 112.035 67.645 112.205 ;
        RECT 68.420 112.185 68.595 112.795 ;
        RECT 69.215 112.785 69.545 113.765 ;
        RECT 69.715 112.795 69.975 113.935 ;
        RECT 70.150 112.795 70.485 113.765 ;
        RECT 70.655 112.795 70.825 113.935 ;
        RECT 70.995 113.595 73.025 113.765 ;
        RECT 68.775 112.355 69.110 112.625 ;
        RECT 69.280 112.185 69.450 112.785 ;
        RECT 69.620 112.375 69.955 112.625 ;
        RECT 66.420 111.555 66.750 112.035 ;
        RECT 66.920 111.385 67.145 111.845 ;
        RECT 67.315 111.555 67.645 112.035 ;
        RECT 67.835 111.385 68.085 112.185 ;
        RECT 68.255 111.555 68.595 112.185 ;
        RECT 68.765 111.385 69.075 112.185 ;
        RECT 69.280 111.555 69.975 112.185 ;
        RECT 70.150 112.125 70.320 112.795 ;
        RECT 70.995 112.625 71.165 113.595 ;
        RECT 70.490 112.295 70.745 112.625 ;
        RECT 70.970 112.295 71.165 112.625 ;
        RECT 71.335 113.255 72.460 113.425 ;
        RECT 70.575 112.125 70.745 112.295 ;
        RECT 71.335 112.125 71.505 113.255 ;
        RECT 70.150 111.555 70.405 112.125 ;
        RECT 70.575 111.955 71.505 112.125 ;
        RECT 71.675 112.915 72.685 113.085 ;
        RECT 71.675 112.115 71.845 112.915 ;
        RECT 72.050 112.575 72.325 112.715 ;
        RECT 72.045 112.405 72.325 112.575 ;
        RECT 71.330 111.920 71.505 111.955 ;
        RECT 70.575 111.385 70.905 111.785 ;
        RECT 71.330 111.555 71.860 111.920 ;
        RECT 72.050 111.555 72.325 112.405 ;
        RECT 72.495 111.555 72.685 112.915 ;
        RECT 72.855 112.930 73.025 113.595 ;
        RECT 73.195 113.175 73.365 113.935 ;
        RECT 73.600 113.175 74.115 113.585 ;
        RECT 72.855 112.740 73.605 112.930 ;
        RECT 73.775 112.365 74.115 113.175 ;
        RECT 74.285 112.845 75.955 113.935 ;
        RECT 72.885 112.195 74.115 112.365 ;
        RECT 72.865 111.385 73.375 111.920 ;
        RECT 73.595 111.590 73.840 112.195 ;
        RECT 74.285 112.155 75.035 112.675 ;
        RECT 75.205 112.325 75.955 112.845 ;
        RECT 76.585 112.770 76.875 113.935 ;
        RECT 77.540 113.145 78.075 113.765 ;
        RECT 74.285 111.385 75.955 112.155 ;
        RECT 77.540 112.125 77.855 113.145 ;
        RECT 78.245 113.135 78.575 113.935 ;
        RECT 79.060 112.965 79.450 113.140 ;
        RECT 78.025 112.795 79.450 112.965 ;
        RECT 79.805 112.845 81.015 113.935 ;
        RECT 81.275 113.265 81.445 113.765 ;
        RECT 81.615 113.435 81.945 113.935 ;
        RECT 81.275 113.095 81.940 113.265 ;
        RECT 78.025 112.295 78.195 112.795 ;
        RECT 76.585 111.385 76.875 112.110 ;
        RECT 77.540 111.555 78.155 112.125 ;
        RECT 78.445 112.065 78.710 112.625 ;
        RECT 78.880 111.895 79.050 112.795 ;
        RECT 79.220 112.065 79.575 112.625 ;
        RECT 79.805 112.135 80.325 112.675 ;
        RECT 80.495 112.305 81.015 112.845 ;
        RECT 81.190 112.275 81.540 112.925 ;
        RECT 78.325 111.385 78.540 111.895 ;
        RECT 78.770 111.565 79.050 111.895 ;
        RECT 79.230 111.385 79.470 111.895 ;
        RECT 79.805 111.385 81.015 112.135 ;
        RECT 81.710 112.105 81.940 113.095 ;
        RECT 81.275 111.935 81.940 112.105 ;
        RECT 81.275 111.645 81.445 111.935 ;
        RECT 81.615 111.385 81.945 111.765 ;
        RECT 82.115 111.645 82.300 113.765 ;
        RECT 82.540 113.475 82.805 113.935 ;
        RECT 82.975 113.340 83.225 113.765 ;
        RECT 83.435 113.490 84.540 113.660 ;
        RECT 82.920 113.210 83.225 113.340 ;
        RECT 82.470 112.015 82.750 112.965 ;
        RECT 82.920 112.105 83.090 113.210 ;
        RECT 83.260 112.425 83.500 113.020 ;
        RECT 83.670 112.955 84.200 113.320 ;
        RECT 83.670 112.255 83.840 112.955 ;
        RECT 84.370 112.875 84.540 113.490 ;
        RECT 84.710 113.135 84.880 113.935 ;
        RECT 85.050 113.435 85.300 113.765 ;
        RECT 85.525 113.465 86.410 113.635 ;
        RECT 84.370 112.785 84.880 112.875 ;
        RECT 82.920 111.975 83.145 112.105 ;
        RECT 83.315 112.035 83.840 112.255 ;
        RECT 84.010 112.615 84.880 112.785 ;
        RECT 82.555 111.385 82.805 111.845 ;
        RECT 82.975 111.835 83.145 111.975 ;
        RECT 84.010 111.835 84.180 112.615 ;
        RECT 84.710 112.545 84.880 112.615 ;
        RECT 84.390 112.365 84.590 112.395 ;
        RECT 85.050 112.365 85.220 113.435 ;
        RECT 85.390 112.545 85.580 113.265 ;
        RECT 84.390 112.065 85.220 112.365 ;
        RECT 85.750 112.335 86.070 113.295 ;
        RECT 82.975 111.665 83.310 111.835 ;
        RECT 83.505 111.665 84.180 111.835 ;
        RECT 84.500 111.385 84.870 111.885 ;
        RECT 85.050 111.835 85.220 112.065 ;
        RECT 85.605 112.005 86.070 112.335 ;
        RECT 86.240 112.625 86.410 113.465 ;
        RECT 86.590 113.435 86.905 113.935 ;
        RECT 87.135 113.205 87.475 113.765 ;
        RECT 86.580 112.830 87.475 113.205 ;
        RECT 87.645 112.925 87.815 113.935 ;
        RECT 87.285 112.625 87.475 112.830 ;
        RECT 87.985 112.875 88.315 113.720 ;
        RECT 87.985 112.795 88.375 112.875 ;
        RECT 88.160 112.745 88.375 112.795 ;
        RECT 86.240 112.295 87.115 112.625 ;
        RECT 87.285 112.295 88.035 112.625 ;
        RECT 86.240 111.835 86.410 112.295 ;
        RECT 87.285 112.125 87.485 112.295 ;
        RECT 88.205 112.165 88.375 112.745 ;
        RECT 88.545 112.845 89.755 113.935 ;
        RECT 88.545 112.305 89.065 112.845 ;
        RECT 88.150 112.125 88.375 112.165 ;
        RECT 89.235 112.135 89.755 112.675 ;
        RECT 85.050 111.665 85.455 111.835 ;
        RECT 85.625 111.665 86.410 111.835 ;
        RECT 86.685 111.385 86.895 111.915 ;
        RECT 87.155 111.600 87.485 112.125 ;
        RECT 87.995 112.040 88.375 112.125 ;
        RECT 87.655 111.385 87.825 111.995 ;
        RECT 87.995 111.605 88.325 112.040 ;
        RECT 88.545 111.385 89.755 112.135 ;
        RECT 12.100 111.215 89.840 111.385 ;
        RECT 12.185 110.465 13.395 111.215 ;
        RECT 14.115 110.665 14.285 110.955 ;
        RECT 14.455 110.835 14.785 111.215 ;
        RECT 14.115 110.495 14.780 110.665 ;
        RECT 12.185 109.925 12.705 110.465 ;
        RECT 12.875 109.755 13.395 110.295 ;
        RECT 12.185 108.665 13.395 109.755 ;
        RECT 14.030 109.675 14.380 110.325 ;
        RECT 14.550 109.505 14.780 110.495 ;
        RECT 14.115 109.335 14.780 109.505 ;
        RECT 14.115 108.835 14.285 109.335 ;
        RECT 14.455 108.665 14.785 109.165 ;
        RECT 14.955 108.835 15.140 110.955 ;
        RECT 15.395 110.755 15.645 111.215 ;
        RECT 15.815 110.765 16.150 110.935 ;
        RECT 16.345 110.765 17.020 110.935 ;
        RECT 15.815 110.625 15.985 110.765 ;
        RECT 15.310 109.635 15.590 110.585 ;
        RECT 15.760 110.495 15.985 110.625 ;
        RECT 15.760 109.390 15.930 110.495 ;
        RECT 16.155 110.345 16.680 110.565 ;
        RECT 16.100 109.580 16.340 110.175 ;
        RECT 16.510 109.645 16.680 110.345 ;
        RECT 16.850 109.985 17.020 110.765 ;
        RECT 17.340 110.715 17.710 111.215 ;
        RECT 17.890 110.765 18.295 110.935 ;
        RECT 18.465 110.765 19.250 110.935 ;
        RECT 17.890 110.535 18.060 110.765 ;
        RECT 17.230 110.235 18.060 110.535 ;
        RECT 18.445 110.265 18.910 110.595 ;
        RECT 17.230 110.205 17.430 110.235 ;
        RECT 17.550 109.985 17.720 110.055 ;
        RECT 16.850 109.815 17.720 109.985 ;
        RECT 17.210 109.725 17.720 109.815 ;
        RECT 15.760 109.260 16.065 109.390 ;
        RECT 16.510 109.280 17.040 109.645 ;
        RECT 15.380 108.665 15.645 109.125 ;
        RECT 15.815 108.835 16.065 109.260 ;
        RECT 17.210 109.110 17.380 109.725 ;
        RECT 16.275 108.940 17.380 109.110 ;
        RECT 17.550 108.665 17.720 109.465 ;
        RECT 17.890 109.165 18.060 110.235 ;
        RECT 18.230 109.335 18.420 110.055 ;
        RECT 18.590 109.305 18.910 110.265 ;
        RECT 19.080 110.305 19.250 110.765 ;
        RECT 19.525 110.685 19.735 111.215 ;
        RECT 19.995 110.475 20.325 111.000 ;
        RECT 20.495 110.605 20.665 111.215 ;
        RECT 20.835 110.560 21.165 110.995 ;
        RECT 20.835 110.475 21.215 110.560 ;
        RECT 20.125 110.305 20.325 110.475 ;
        RECT 20.990 110.435 21.215 110.475 ;
        RECT 19.080 109.975 19.955 110.305 ;
        RECT 20.125 109.975 20.875 110.305 ;
        RECT 17.890 108.835 18.140 109.165 ;
        RECT 19.080 109.135 19.250 109.975 ;
        RECT 20.125 109.770 20.315 109.975 ;
        RECT 21.045 109.855 21.215 110.435 ;
        RECT 21.385 110.380 21.675 111.215 ;
        RECT 21.845 110.815 22.800 110.985 ;
        RECT 23.215 110.825 23.545 111.215 ;
        RECT 21.845 109.935 22.015 110.815 ;
        RECT 23.715 110.645 23.885 110.965 ;
        RECT 24.055 110.825 24.385 111.215 ;
        RECT 25.525 110.715 25.865 111.215 ;
        RECT 22.185 110.475 24.435 110.645 ;
        RECT 22.185 109.975 22.415 110.475 ;
        RECT 22.585 110.055 22.960 110.225 ;
        RECT 21.000 109.805 21.215 109.855 ;
        RECT 19.420 109.395 20.315 109.770 ;
        RECT 20.825 109.725 21.215 109.805 ;
        RECT 21.385 109.765 22.015 109.935 ;
        RECT 22.790 109.855 22.960 110.055 ;
        RECT 23.130 110.025 23.680 110.225 ;
        RECT 23.850 109.855 24.095 110.305 ;
        RECT 18.365 108.965 19.250 109.135 ;
        RECT 19.430 108.665 19.745 109.165 ;
        RECT 19.975 108.835 20.315 109.395 ;
        RECT 20.485 108.665 20.655 109.675 ;
        RECT 20.825 108.880 21.155 109.725 ;
        RECT 21.385 108.835 21.705 109.765 ;
        RECT 22.790 109.685 24.095 109.855 ;
        RECT 24.265 109.515 24.435 110.475 ;
        RECT 25.525 109.975 25.865 110.545 ;
        RECT 26.035 110.305 26.280 110.995 ;
        RECT 26.475 110.715 26.805 111.215 ;
        RECT 27.005 110.645 27.175 110.995 ;
        RECT 27.350 110.815 27.680 111.215 ;
        RECT 27.850 110.645 28.020 110.995 ;
        RECT 28.190 110.815 28.570 111.215 ;
        RECT 27.005 110.475 28.590 110.645 ;
        RECT 28.760 110.540 29.035 110.885 ;
        RECT 30.180 110.820 30.880 110.990 ;
        RECT 31.125 110.850 32.580 111.030 ;
        RECT 30.180 110.705 30.350 110.820 ;
        RECT 31.125 110.645 31.295 110.850 ;
        RECT 32.940 110.845 34.255 111.045 ;
        RECT 34.425 110.855 34.755 111.215 ;
        RECT 35.285 110.855 35.615 111.215 ;
        RECT 34.025 110.675 34.255 110.845 ;
        RECT 36.225 110.775 36.395 111.215 ;
        RECT 36.620 110.675 36.835 110.875 ;
        RECT 37.005 110.855 37.335 111.215 ;
        RECT 37.505 110.675 37.705 110.765 ;
        RECT 28.420 110.305 28.590 110.475 ;
        RECT 26.035 109.975 26.690 110.305 ;
        RECT 21.885 109.345 23.125 109.515 ;
        RECT 21.885 108.835 22.285 109.345 ;
        RECT 22.455 108.665 22.625 109.175 ;
        RECT 22.795 108.835 23.125 109.345 ;
        RECT 23.295 108.665 23.465 109.515 ;
        RECT 24.055 108.835 24.435 109.515 ;
        RECT 25.525 108.665 25.865 109.740 ;
        RECT 26.035 109.380 26.275 109.975 ;
        RECT 26.470 109.515 26.790 109.805 ;
        RECT 26.960 109.685 27.700 110.305 ;
        RECT 27.870 109.975 28.250 110.305 ;
        RECT 28.420 109.975 28.695 110.305 ;
        RECT 28.420 109.805 28.590 109.975 ;
        RECT 28.865 109.805 29.035 110.540 ;
        RECT 30.510 110.475 31.295 110.645 ;
        RECT 31.690 110.485 33.855 110.665 ;
        RECT 34.025 110.605 36.085 110.675 ;
        RECT 36.620 110.605 37.705 110.675 ;
        RECT 34.025 110.505 37.705 110.605 ;
        RECT 30.510 109.960 30.690 110.475 ;
        RECT 34.730 110.435 37.705 110.505 ;
        RECT 37.945 110.490 38.235 111.215 ;
        RECT 38.455 110.560 38.785 110.995 ;
        RECT 38.955 110.605 39.125 111.215 ;
        RECT 36.065 110.395 37.705 110.435 ;
        RECT 38.405 110.475 38.785 110.560 ;
        RECT 39.295 110.475 39.625 111.000 ;
        RECT 39.885 110.685 40.095 111.215 ;
        RECT 40.370 110.765 41.155 110.935 ;
        RECT 41.325 110.765 41.730 110.935 ;
        RECT 38.405 110.435 38.630 110.475 ;
        RECT 27.930 109.635 28.590 109.805 ;
        RECT 27.930 109.515 28.100 109.635 ;
        RECT 26.470 109.345 28.100 109.515 ;
        RECT 26.045 109.005 28.100 109.175 ;
        RECT 26.050 108.885 28.100 109.005 ;
        RECT 28.270 108.665 28.550 109.465 ;
        RECT 28.760 108.835 29.035 109.805 ;
        RECT 30.180 109.445 30.690 109.960 ;
        RECT 30.860 109.785 31.030 110.305 ;
        RECT 31.420 109.955 32.490 110.225 ;
        RECT 32.885 109.890 34.060 110.305 ;
        RECT 32.885 109.785 33.600 109.890 ;
        RECT 30.860 109.615 33.600 109.785 ;
        RECT 34.230 109.785 34.510 110.305 ;
        RECT 34.680 109.955 36.155 110.225 ;
        RECT 36.450 109.970 37.460 110.225 ;
        RECT 36.450 109.785 36.895 109.970 ;
        RECT 38.405 109.855 38.575 110.435 ;
        RECT 39.295 110.305 39.495 110.475 ;
        RECT 40.370 110.305 40.540 110.765 ;
        RECT 38.745 109.975 39.495 110.305 ;
        RECT 39.665 109.975 40.540 110.305 ;
        RECT 34.230 109.615 36.895 109.785 ;
        RECT 33.865 109.445 34.035 109.515 ;
        RECT 30.180 109.275 36.055 109.445 ;
        RECT 37.085 109.365 37.305 109.440 ;
        RECT 30.180 109.195 33.815 109.275 ;
        RECT 34.390 109.195 36.055 109.275 ;
        RECT 36.225 109.195 37.305 109.365 ;
        RECT 30.175 108.665 30.505 109.025 ;
        RECT 31.405 108.665 31.740 109.025 ;
        RECT 32.250 108.665 32.580 109.025 ;
        RECT 33.095 108.665 33.425 109.025 ;
        RECT 33.975 108.665 34.245 109.105 ;
        RECT 36.225 109.025 36.405 109.195 ;
        RECT 37.085 109.110 37.305 109.195 ;
        RECT 34.425 108.835 36.405 109.025 ;
        RECT 36.575 108.665 36.905 109.025 ;
        RECT 37.475 108.665 37.770 109.635 ;
        RECT 37.945 108.665 38.235 109.830 ;
        RECT 38.405 109.805 38.620 109.855 ;
        RECT 38.405 109.725 38.795 109.805 ;
        RECT 38.465 108.880 38.795 109.725 ;
        RECT 39.305 109.770 39.495 109.975 ;
        RECT 38.965 108.665 39.135 109.675 ;
        RECT 39.305 109.395 40.200 109.770 ;
        RECT 39.305 108.835 39.645 109.395 ;
        RECT 39.875 108.665 40.190 109.165 ;
        RECT 40.370 109.135 40.540 109.975 ;
        RECT 40.710 110.265 41.175 110.595 ;
        RECT 41.560 110.535 41.730 110.765 ;
        RECT 41.910 110.715 42.280 111.215 ;
        RECT 42.600 110.765 43.275 110.935 ;
        RECT 43.470 110.765 43.805 110.935 ;
        RECT 40.710 109.305 41.030 110.265 ;
        RECT 41.560 110.235 42.390 110.535 ;
        RECT 41.200 109.335 41.390 110.055 ;
        RECT 41.560 109.165 41.730 110.235 ;
        RECT 42.190 110.205 42.390 110.235 ;
        RECT 41.900 109.985 42.070 110.055 ;
        RECT 42.600 109.985 42.770 110.765 ;
        RECT 43.635 110.625 43.805 110.765 ;
        RECT 43.975 110.755 44.225 111.215 ;
        RECT 41.900 109.815 42.770 109.985 ;
        RECT 42.940 110.345 43.465 110.565 ;
        RECT 43.635 110.495 43.860 110.625 ;
        RECT 41.900 109.725 42.410 109.815 ;
        RECT 40.370 108.965 41.255 109.135 ;
        RECT 41.480 108.835 41.730 109.165 ;
        RECT 41.900 108.665 42.070 109.465 ;
        RECT 42.240 109.110 42.410 109.725 ;
        RECT 42.940 109.645 43.110 110.345 ;
        RECT 42.580 109.280 43.110 109.645 ;
        RECT 43.280 109.580 43.520 110.175 ;
        RECT 43.690 109.390 43.860 110.495 ;
        RECT 44.030 109.635 44.310 110.585 ;
        RECT 43.555 109.260 43.860 109.390 ;
        RECT 42.240 108.940 43.345 109.110 ;
        RECT 43.555 108.835 43.805 109.260 ;
        RECT 43.975 108.665 44.240 109.125 ;
        RECT 44.480 108.835 44.665 110.955 ;
        RECT 44.835 110.835 45.165 111.215 ;
        RECT 45.335 110.665 45.505 110.955 ;
        RECT 44.840 110.495 45.505 110.665 ;
        RECT 44.840 109.505 45.070 110.495 ;
        RECT 45.765 110.465 46.975 111.215 ;
        RECT 47.145 110.475 47.530 111.045 ;
        RECT 47.700 110.755 48.025 111.215 ;
        RECT 48.545 110.585 48.825 111.045 ;
        RECT 45.240 109.675 45.590 110.325 ;
        RECT 45.765 109.925 46.285 110.465 ;
        RECT 46.455 109.755 46.975 110.295 ;
        RECT 44.840 109.335 45.505 109.505 ;
        RECT 44.835 108.665 45.165 109.165 ;
        RECT 45.335 108.835 45.505 109.335 ;
        RECT 45.765 108.665 46.975 109.755 ;
        RECT 47.145 109.805 47.425 110.475 ;
        RECT 47.700 110.415 48.825 110.585 ;
        RECT 47.700 110.305 48.150 110.415 ;
        RECT 47.595 109.975 48.150 110.305 ;
        RECT 49.015 110.245 49.415 111.045 ;
        RECT 49.815 110.755 50.085 111.215 ;
        RECT 50.255 110.585 50.540 111.045 ;
        RECT 47.145 108.835 47.530 109.805 ;
        RECT 47.700 109.515 48.150 109.975 ;
        RECT 48.320 109.685 49.415 110.245 ;
        RECT 47.700 109.295 48.825 109.515 ;
        RECT 47.700 108.665 48.025 109.125 ;
        RECT 48.545 108.835 48.825 109.295 ;
        RECT 49.015 108.835 49.415 109.685 ;
        RECT 49.585 110.415 50.540 110.585 ;
        RECT 50.825 110.475 51.210 111.045 ;
        RECT 51.380 110.755 51.705 111.215 ;
        RECT 52.225 110.585 52.505 111.045 ;
        RECT 49.585 109.515 49.795 110.415 ;
        RECT 49.965 109.685 50.655 110.245 ;
        RECT 50.825 109.805 51.105 110.475 ;
        RECT 51.380 110.415 52.505 110.585 ;
        RECT 51.380 110.305 51.830 110.415 ;
        RECT 51.275 109.975 51.830 110.305 ;
        RECT 52.695 110.245 53.095 111.045 ;
        RECT 53.495 110.755 53.765 111.215 ;
        RECT 53.935 110.585 54.220 111.045 ;
        RECT 49.585 109.295 50.540 109.515 ;
        RECT 49.815 108.665 50.085 109.125 ;
        RECT 50.255 108.835 50.540 109.295 ;
        RECT 50.825 108.835 51.210 109.805 ;
        RECT 51.380 109.515 51.830 109.975 ;
        RECT 52.000 109.685 53.095 110.245 ;
        RECT 51.380 109.295 52.505 109.515 ;
        RECT 51.380 108.665 51.705 109.125 ;
        RECT 52.225 108.835 52.505 109.295 ;
        RECT 52.695 108.835 53.095 109.685 ;
        RECT 53.265 110.415 54.220 110.585 ;
        RECT 54.505 110.445 58.015 111.215 ;
        RECT 58.185 110.465 59.395 111.215 ;
        RECT 59.575 110.490 59.905 111.000 ;
        RECT 60.075 110.815 60.405 111.215 ;
        RECT 61.455 110.645 61.785 110.985 ;
        RECT 61.955 110.815 62.285 111.215 ;
        RECT 53.265 109.515 53.475 110.415 ;
        RECT 53.645 109.685 54.335 110.245 ;
        RECT 54.505 109.925 56.155 110.445 ;
        RECT 56.325 109.755 58.015 110.275 ;
        RECT 58.185 109.925 58.705 110.465 ;
        RECT 58.875 109.755 59.395 110.295 ;
        RECT 53.265 109.295 54.220 109.515 ;
        RECT 53.495 108.665 53.765 109.125 ;
        RECT 53.935 108.835 54.220 109.295 ;
        RECT 54.505 108.665 58.015 109.755 ;
        RECT 58.185 108.665 59.395 109.755 ;
        RECT 59.575 109.725 59.765 110.490 ;
        RECT 60.075 110.475 62.440 110.645 ;
        RECT 63.705 110.490 63.995 111.215 ;
        RECT 60.075 110.305 60.245 110.475 ;
        RECT 59.935 109.975 60.245 110.305 ;
        RECT 60.415 109.975 60.720 110.305 ;
        RECT 59.575 108.875 59.905 109.725 ;
        RECT 60.075 108.665 60.325 109.805 ;
        RECT 60.505 109.645 60.720 109.975 ;
        RECT 60.895 109.645 61.180 110.305 ;
        RECT 61.375 109.645 61.640 110.305 ;
        RECT 61.855 109.645 62.100 110.305 ;
        RECT 62.270 109.475 62.440 110.475 ;
        RECT 64.205 110.395 64.435 111.215 ;
        RECT 64.605 110.415 64.935 111.045 ;
        RECT 64.185 109.975 64.515 110.225 ;
        RECT 60.515 109.305 61.805 109.475 ;
        RECT 60.515 108.885 60.765 109.305 ;
        RECT 60.995 108.665 61.325 109.135 ;
        RECT 61.555 108.885 61.805 109.305 ;
        RECT 61.985 109.305 62.440 109.475 ;
        RECT 61.985 108.875 62.315 109.305 ;
        RECT 63.705 108.665 63.995 109.830 ;
        RECT 64.685 109.815 64.935 110.415 ;
        RECT 65.105 110.395 65.315 111.215 ;
        RECT 65.545 110.445 69.055 111.215 ;
        RECT 65.545 109.925 67.195 110.445 ;
        RECT 70.350 110.435 70.850 111.045 ;
        RECT 64.205 108.665 64.435 109.805 ;
        RECT 64.605 108.835 64.935 109.815 ;
        RECT 65.105 108.665 65.315 109.805 ;
        RECT 67.365 109.755 69.055 110.275 ;
        RECT 70.145 109.975 70.495 110.225 ;
        RECT 70.680 109.805 70.850 110.435 ;
        RECT 71.480 110.565 71.810 111.045 ;
        RECT 71.980 110.755 72.205 111.215 ;
        RECT 72.375 110.565 72.705 111.045 ;
        RECT 71.480 110.395 72.705 110.565 ;
        RECT 72.895 110.415 73.145 111.215 ;
        RECT 73.315 110.415 73.655 111.045 ;
        RECT 73.915 110.665 74.085 110.955 ;
        RECT 74.255 110.835 74.585 111.215 ;
        RECT 73.915 110.495 74.580 110.665 ;
        RECT 73.425 110.365 73.655 110.415 ;
        RECT 71.020 110.025 71.350 110.225 ;
        RECT 71.520 110.025 71.850 110.225 ;
        RECT 72.020 110.025 72.440 110.225 ;
        RECT 72.615 110.055 73.310 110.225 ;
        RECT 72.615 109.805 72.785 110.055 ;
        RECT 73.480 109.805 73.655 110.365 ;
        RECT 65.545 108.665 69.055 109.755 ;
        RECT 70.350 109.635 72.785 109.805 ;
        RECT 70.350 108.835 70.680 109.635 ;
        RECT 70.850 108.665 71.180 109.465 ;
        RECT 71.480 108.835 71.810 109.635 ;
        RECT 72.455 108.665 72.705 109.465 ;
        RECT 72.975 108.665 73.145 109.805 ;
        RECT 73.315 108.835 73.655 109.805 ;
        RECT 73.830 109.675 74.180 110.325 ;
        RECT 74.350 109.505 74.580 110.495 ;
        RECT 73.915 109.335 74.580 109.505 ;
        RECT 73.915 108.835 74.085 109.335 ;
        RECT 74.255 108.665 74.585 109.165 ;
        RECT 74.755 108.835 74.940 110.955 ;
        RECT 75.195 110.755 75.445 111.215 ;
        RECT 75.615 110.765 75.950 110.935 ;
        RECT 76.145 110.765 76.820 110.935 ;
        RECT 75.615 110.625 75.785 110.765 ;
        RECT 75.110 109.635 75.390 110.585 ;
        RECT 75.560 110.495 75.785 110.625 ;
        RECT 75.560 109.390 75.730 110.495 ;
        RECT 75.955 110.345 76.480 110.565 ;
        RECT 75.900 109.580 76.140 110.175 ;
        RECT 76.310 109.645 76.480 110.345 ;
        RECT 76.650 109.985 76.820 110.765 ;
        RECT 77.140 110.715 77.510 111.215 ;
        RECT 77.690 110.765 78.095 110.935 ;
        RECT 78.265 110.765 79.050 110.935 ;
        RECT 77.690 110.535 77.860 110.765 ;
        RECT 77.030 110.235 77.860 110.535 ;
        RECT 78.245 110.265 78.710 110.595 ;
        RECT 77.030 110.205 77.230 110.235 ;
        RECT 77.350 109.985 77.520 110.055 ;
        RECT 76.650 109.815 77.520 109.985 ;
        RECT 77.010 109.725 77.520 109.815 ;
        RECT 75.560 109.260 75.865 109.390 ;
        RECT 76.310 109.280 76.840 109.645 ;
        RECT 75.180 108.665 75.445 109.125 ;
        RECT 75.615 108.835 75.865 109.260 ;
        RECT 77.010 109.110 77.180 109.725 ;
        RECT 76.075 108.940 77.180 109.110 ;
        RECT 77.350 108.665 77.520 109.465 ;
        RECT 77.690 109.165 77.860 110.235 ;
        RECT 78.030 109.335 78.220 110.055 ;
        RECT 78.390 109.305 78.710 110.265 ;
        RECT 78.880 110.305 79.050 110.765 ;
        RECT 79.325 110.685 79.535 111.215 ;
        RECT 79.795 110.475 80.125 111.000 ;
        RECT 80.295 110.605 80.465 111.215 ;
        RECT 80.635 110.560 80.965 110.995 ;
        RECT 80.635 110.475 81.015 110.560 ;
        RECT 79.925 110.305 80.125 110.475 ;
        RECT 80.790 110.435 81.015 110.475 ;
        RECT 78.880 109.975 79.755 110.305 ;
        RECT 79.925 109.975 80.675 110.305 ;
        RECT 77.690 108.835 77.940 109.165 ;
        RECT 78.880 109.135 79.050 109.975 ;
        RECT 79.925 109.770 80.115 109.975 ;
        RECT 80.845 109.855 81.015 110.435 ;
        RECT 80.800 109.805 81.015 109.855 ;
        RECT 79.220 109.395 80.115 109.770 ;
        RECT 80.625 109.725 81.015 109.805 ;
        RECT 81.185 110.415 81.525 111.045 ;
        RECT 81.695 110.415 81.945 111.215 ;
        RECT 82.135 110.565 82.465 111.045 ;
        RECT 82.635 110.755 82.860 111.215 ;
        RECT 83.030 110.565 83.360 111.045 ;
        RECT 81.185 109.805 81.360 110.415 ;
        RECT 82.135 110.395 83.360 110.565 ;
        RECT 83.990 110.435 84.490 111.045 ;
        RECT 81.530 110.055 82.225 110.225 ;
        RECT 82.055 109.805 82.225 110.055 ;
        RECT 82.400 110.025 82.820 110.225 ;
        RECT 82.990 110.025 83.320 110.225 ;
        RECT 83.490 110.025 83.820 110.225 ;
        RECT 83.990 109.805 84.160 110.435 ;
        RECT 84.345 109.975 84.695 110.225 ;
        RECT 78.165 108.965 79.050 109.135 ;
        RECT 79.230 108.665 79.545 109.165 ;
        RECT 79.775 108.835 80.115 109.395 ;
        RECT 80.285 108.665 80.455 109.675 ;
        RECT 80.625 108.880 80.955 109.725 ;
        RECT 81.185 108.835 81.525 109.805 ;
        RECT 81.695 108.665 81.865 109.805 ;
        RECT 82.055 109.635 84.490 109.805 ;
        RECT 82.135 108.665 82.385 109.465 ;
        RECT 83.030 108.835 83.360 109.635 ;
        RECT 83.660 108.665 83.990 109.465 ;
        RECT 84.160 108.835 84.490 109.635 ;
        RECT 84.870 109.615 85.205 111.035 ;
        RECT 85.385 110.845 86.130 111.215 ;
        RECT 86.695 110.675 86.950 111.035 ;
        RECT 87.130 110.845 87.460 111.215 ;
        RECT 87.640 110.675 87.865 111.035 ;
        RECT 85.380 110.485 87.865 110.675 ;
        RECT 85.380 109.795 85.605 110.485 ;
        RECT 88.545 110.465 89.755 111.215 ;
        RECT 85.805 109.975 86.085 110.305 ;
        RECT 86.265 109.975 86.840 110.305 ;
        RECT 87.020 109.975 87.455 110.305 ;
        RECT 87.635 109.975 87.905 110.305 ;
        RECT 85.380 109.615 87.875 109.795 ;
        RECT 84.870 108.845 85.135 109.615 ;
        RECT 85.305 108.665 85.635 109.385 ;
        RECT 85.825 109.205 87.015 109.435 ;
        RECT 85.825 108.845 86.085 109.205 ;
        RECT 86.255 108.665 86.585 109.035 ;
        RECT 86.755 108.845 87.015 109.205 ;
        RECT 87.585 108.845 87.875 109.615 ;
        RECT 88.545 109.755 89.065 110.295 ;
        RECT 89.235 109.925 89.755 110.465 ;
        RECT 100.090 110.950 100.760 114.210 ;
        RECT 101.430 113.640 105.470 113.810 ;
        RECT 101.090 111.580 101.260 113.580 ;
        RECT 105.640 111.580 105.810 113.580 ;
        RECT 101.430 111.350 105.470 111.520 ;
        RECT 106.150 110.950 106.320 114.210 ;
        RECT 100.090 110.780 106.320 110.950 ;
        RECT 88.545 108.665 89.755 109.755 ;
        RECT 12.100 108.495 89.840 108.665 ;
        RECT 12.185 107.405 13.395 108.495 ;
        RECT 13.655 107.825 13.825 108.325 ;
        RECT 13.995 107.995 14.325 108.495 ;
        RECT 13.655 107.655 14.320 107.825 ;
        RECT 12.185 106.695 12.705 107.235 ;
        RECT 12.875 106.865 13.395 107.405 ;
        RECT 13.570 106.835 13.920 107.485 ;
        RECT 12.185 105.945 13.395 106.695 ;
        RECT 14.090 106.665 14.320 107.655 ;
        RECT 13.655 106.495 14.320 106.665 ;
        RECT 13.655 106.205 13.825 106.495 ;
        RECT 13.995 105.945 14.325 106.325 ;
        RECT 14.495 106.205 14.680 108.325 ;
        RECT 14.920 108.035 15.185 108.495 ;
        RECT 15.355 107.900 15.605 108.325 ;
        RECT 15.815 108.050 16.920 108.220 ;
        RECT 15.300 107.770 15.605 107.900 ;
        RECT 14.850 106.575 15.130 107.525 ;
        RECT 15.300 106.665 15.470 107.770 ;
        RECT 15.640 106.985 15.880 107.580 ;
        RECT 16.050 107.515 16.580 107.880 ;
        RECT 16.050 106.815 16.220 107.515 ;
        RECT 16.750 107.435 16.920 108.050 ;
        RECT 17.090 107.695 17.260 108.495 ;
        RECT 17.430 107.995 17.680 108.325 ;
        RECT 17.905 108.025 18.790 108.195 ;
        RECT 16.750 107.345 17.260 107.435 ;
        RECT 15.300 106.535 15.525 106.665 ;
        RECT 15.695 106.595 16.220 106.815 ;
        RECT 16.390 107.175 17.260 107.345 ;
        RECT 14.935 105.945 15.185 106.405 ;
        RECT 15.355 106.395 15.525 106.535 ;
        RECT 16.390 106.395 16.560 107.175 ;
        RECT 17.090 107.105 17.260 107.175 ;
        RECT 16.770 106.925 16.970 106.955 ;
        RECT 17.430 106.925 17.600 107.995 ;
        RECT 17.770 107.105 17.960 107.825 ;
        RECT 16.770 106.625 17.600 106.925 ;
        RECT 18.130 106.895 18.450 107.855 ;
        RECT 15.355 106.225 15.690 106.395 ;
        RECT 15.885 106.225 16.560 106.395 ;
        RECT 16.880 105.945 17.250 106.445 ;
        RECT 17.430 106.395 17.600 106.625 ;
        RECT 17.985 106.565 18.450 106.895 ;
        RECT 18.620 107.185 18.790 108.025 ;
        RECT 18.970 107.995 19.285 108.495 ;
        RECT 19.515 107.765 19.855 108.325 ;
        RECT 18.960 107.390 19.855 107.765 ;
        RECT 20.025 107.485 20.195 108.495 ;
        RECT 19.665 107.185 19.855 107.390 ;
        RECT 20.365 107.435 20.695 108.280 ;
        RECT 20.365 107.355 20.755 107.435 ;
        RECT 20.925 107.405 22.135 108.495 ;
        RECT 22.315 107.775 22.645 108.495 ;
        RECT 20.540 107.305 20.755 107.355 ;
        RECT 18.620 106.855 19.495 107.185 ;
        RECT 19.665 106.855 20.415 107.185 ;
        RECT 18.620 106.395 18.790 106.855 ;
        RECT 19.665 106.685 19.865 106.855 ;
        RECT 20.585 106.725 20.755 107.305 ;
        RECT 20.530 106.685 20.755 106.725 ;
        RECT 17.430 106.225 17.835 106.395 ;
        RECT 18.005 106.225 18.790 106.395 ;
        RECT 19.065 105.945 19.275 106.475 ;
        RECT 19.535 106.160 19.865 106.685 ;
        RECT 20.375 106.600 20.755 106.685 ;
        RECT 20.925 106.695 21.445 107.235 ;
        RECT 21.615 106.865 22.135 107.405 ;
        RECT 22.305 107.135 22.535 107.475 ;
        RECT 22.825 107.135 23.040 108.250 ;
        RECT 23.235 107.550 23.565 108.325 ;
        RECT 23.735 107.720 24.445 108.495 ;
        RECT 23.235 107.335 24.385 107.550 ;
        RECT 22.305 106.935 22.635 107.135 ;
        RECT 22.825 106.955 23.275 107.135 ;
        RECT 22.945 106.935 23.275 106.955 ;
        RECT 23.445 106.935 23.915 107.165 ;
        RECT 24.100 106.765 24.385 107.335 ;
        RECT 24.615 106.890 24.895 108.325 ;
        RECT 25.065 107.330 25.355 108.495 ;
        RECT 25.525 107.405 27.195 108.495 ;
        RECT 20.035 105.945 20.205 106.555 ;
        RECT 20.375 106.165 20.705 106.600 ;
        RECT 20.925 105.945 22.135 106.695 ;
        RECT 22.305 106.575 23.485 106.765 ;
        RECT 22.305 106.115 22.645 106.575 ;
        RECT 23.155 106.495 23.485 106.575 ;
        RECT 23.675 106.575 24.385 106.765 ;
        RECT 23.675 106.435 23.975 106.575 ;
        RECT 23.660 106.425 23.975 106.435 ;
        RECT 23.650 106.415 23.975 106.425 ;
        RECT 23.640 106.410 23.975 106.415 ;
        RECT 22.815 105.945 22.985 106.405 ;
        RECT 23.635 106.400 23.975 106.410 ;
        RECT 23.630 106.395 23.975 106.400 ;
        RECT 23.625 106.385 23.975 106.395 ;
        RECT 23.620 106.380 23.975 106.385 ;
        RECT 23.615 106.115 23.975 106.380 ;
        RECT 24.215 105.945 24.385 106.405 ;
        RECT 24.555 106.115 24.895 106.890 ;
        RECT 25.525 106.715 26.275 107.235 ;
        RECT 26.445 106.885 27.195 107.405 ;
        RECT 27.365 107.355 27.635 108.325 ;
        RECT 27.845 107.695 28.125 108.495 ;
        RECT 28.295 107.985 29.950 108.275 ;
        RECT 30.125 107.985 30.425 108.495 ;
        RECT 30.595 107.815 30.925 108.325 ;
        RECT 31.095 107.985 31.725 108.495 ;
        RECT 32.305 107.985 32.685 108.155 ;
        RECT 32.855 107.985 33.155 108.495 ;
        RECT 32.515 107.815 32.685 107.985 ;
        RECT 33.435 107.825 33.605 108.325 ;
        RECT 33.775 107.995 34.105 108.495 ;
        RECT 28.360 107.645 29.950 107.815 ;
        RECT 28.360 107.525 28.530 107.645 ;
        RECT 27.805 107.355 28.530 107.525 ;
        RECT 25.065 105.945 25.355 106.670 ;
        RECT 25.525 105.945 27.195 106.715 ;
        RECT 27.365 106.620 27.535 107.355 ;
        RECT 27.805 107.185 27.975 107.355 ;
        RECT 27.705 106.855 27.975 107.185 ;
        RECT 28.145 106.855 28.550 107.185 ;
        RECT 28.720 106.855 29.430 107.475 ;
        RECT 29.630 107.355 29.950 107.645 ;
        RECT 30.125 107.645 32.345 107.815 ;
        RECT 27.805 106.685 27.975 106.855 ;
        RECT 27.365 106.275 27.635 106.620 ;
        RECT 27.805 106.515 29.415 106.685 ;
        RECT 29.600 106.615 29.950 107.185 ;
        RECT 30.125 106.685 30.295 107.645 ;
        RECT 30.465 107.305 32.005 107.475 ;
        RECT 30.465 106.855 30.710 107.305 ;
        RECT 30.970 106.935 31.665 107.135 ;
        RECT 31.835 107.105 32.005 107.305 ;
        RECT 32.175 107.445 32.345 107.645 ;
        RECT 32.515 107.615 33.175 107.815 ;
        RECT 33.435 107.655 34.100 107.825 ;
        RECT 32.175 107.275 32.835 107.445 ;
        RECT 31.835 106.935 32.435 107.105 ;
        RECT 32.665 106.855 32.835 107.275 ;
        RECT 27.825 105.945 28.205 106.345 ;
        RECT 28.375 106.165 28.545 106.515 ;
        RECT 28.715 105.945 29.045 106.345 ;
        RECT 29.245 106.165 29.415 106.515 ;
        RECT 29.615 105.945 29.945 106.445 ;
        RECT 30.125 106.140 30.590 106.685 ;
        RECT 31.095 105.945 31.265 106.765 ;
        RECT 31.435 106.685 32.345 106.765 ;
        RECT 33.005 106.685 33.175 107.615 ;
        RECT 33.350 106.835 33.700 107.485 ;
        RECT 31.435 106.595 32.685 106.685 ;
        RECT 31.435 106.115 31.765 106.595 ;
        RECT 32.175 106.515 32.685 106.595 ;
        RECT 31.935 105.945 32.285 106.335 ;
        RECT 32.455 106.115 32.685 106.515 ;
        RECT 32.855 106.205 33.175 106.685 ;
        RECT 33.870 106.665 34.100 107.655 ;
        RECT 33.435 106.495 34.100 106.665 ;
        RECT 33.435 106.205 33.605 106.495 ;
        RECT 33.775 105.945 34.105 106.325 ;
        RECT 34.275 106.205 34.460 108.325 ;
        RECT 34.700 108.035 34.965 108.495 ;
        RECT 35.135 107.900 35.385 108.325 ;
        RECT 35.595 108.050 36.700 108.220 ;
        RECT 35.080 107.770 35.385 107.900 ;
        RECT 34.630 106.575 34.910 107.525 ;
        RECT 35.080 106.665 35.250 107.770 ;
        RECT 35.420 106.985 35.660 107.580 ;
        RECT 35.830 107.515 36.360 107.880 ;
        RECT 35.830 106.815 36.000 107.515 ;
        RECT 36.530 107.435 36.700 108.050 ;
        RECT 36.870 107.695 37.040 108.495 ;
        RECT 37.210 107.995 37.460 108.325 ;
        RECT 37.685 108.025 38.570 108.195 ;
        RECT 36.530 107.345 37.040 107.435 ;
        RECT 35.080 106.535 35.305 106.665 ;
        RECT 35.475 106.595 36.000 106.815 ;
        RECT 36.170 107.175 37.040 107.345 ;
        RECT 34.715 105.945 34.965 106.405 ;
        RECT 35.135 106.395 35.305 106.535 ;
        RECT 36.170 106.395 36.340 107.175 ;
        RECT 36.870 107.105 37.040 107.175 ;
        RECT 36.550 106.925 36.750 106.955 ;
        RECT 37.210 106.925 37.380 107.995 ;
        RECT 37.550 107.105 37.740 107.825 ;
        RECT 36.550 106.625 37.380 106.925 ;
        RECT 37.910 106.895 38.230 107.855 ;
        RECT 35.135 106.225 35.470 106.395 ;
        RECT 35.665 106.225 36.340 106.395 ;
        RECT 36.660 105.945 37.030 106.445 ;
        RECT 37.210 106.395 37.380 106.625 ;
        RECT 37.765 106.565 38.230 106.895 ;
        RECT 38.400 107.185 38.570 108.025 ;
        RECT 38.750 107.995 39.065 108.495 ;
        RECT 39.295 107.765 39.635 108.325 ;
        RECT 38.740 107.390 39.635 107.765 ;
        RECT 39.805 107.485 39.975 108.495 ;
        RECT 39.445 107.185 39.635 107.390 ;
        RECT 40.145 107.435 40.475 108.280 ;
        RECT 40.145 107.355 40.535 107.435 ;
        RECT 40.705 107.405 44.215 108.495 ;
        RECT 40.320 107.305 40.535 107.355 ;
        RECT 38.400 106.855 39.275 107.185 ;
        RECT 39.445 106.855 40.195 107.185 ;
        RECT 38.400 106.395 38.570 106.855 ;
        RECT 39.445 106.685 39.645 106.855 ;
        RECT 40.365 106.725 40.535 107.305 ;
        RECT 40.310 106.685 40.535 106.725 ;
        RECT 37.210 106.225 37.615 106.395 ;
        RECT 37.785 106.225 38.570 106.395 ;
        RECT 38.845 105.945 39.055 106.475 ;
        RECT 39.315 106.160 39.645 106.685 ;
        RECT 40.155 106.600 40.535 106.685 ;
        RECT 40.705 106.715 42.355 107.235 ;
        RECT 42.525 106.885 44.215 107.405 ;
        RECT 44.590 107.525 44.920 108.325 ;
        RECT 45.090 107.695 45.420 108.495 ;
        RECT 45.720 107.525 46.050 108.325 ;
        RECT 46.695 107.695 46.945 108.495 ;
        RECT 44.590 107.355 47.025 107.525 ;
        RECT 47.215 107.355 47.385 108.495 ;
        RECT 47.555 107.355 47.895 108.325 ;
        RECT 48.115 108.035 48.325 108.495 ;
        RECT 48.815 107.905 49.315 108.325 ;
        RECT 44.385 106.935 44.735 107.185 ;
        RECT 44.920 106.725 45.090 107.355 ;
        RECT 45.260 106.935 45.590 107.135 ;
        RECT 45.760 106.935 46.090 107.135 ;
        RECT 46.260 106.935 46.680 107.135 ;
        RECT 46.855 107.105 47.025 107.355 ;
        RECT 47.665 107.305 47.895 107.355 ;
        RECT 46.855 106.935 47.550 107.105 ;
        RECT 39.815 105.945 39.985 106.555 ;
        RECT 40.155 106.165 40.485 106.600 ;
        RECT 40.705 105.945 44.215 106.715 ;
        RECT 44.590 106.115 45.090 106.725 ;
        RECT 45.720 106.595 46.945 106.765 ;
        RECT 47.720 106.745 47.895 107.305 ;
        RECT 45.720 106.115 46.050 106.595 ;
        RECT 46.220 105.945 46.445 106.405 ;
        RECT 46.615 106.115 46.945 106.595 ;
        RECT 47.135 105.945 47.385 106.745 ;
        RECT 47.555 106.115 47.895 106.745 ;
        RECT 48.065 106.525 48.305 107.850 ;
        RECT 48.475 107.695 49.315 107.905 ;
        RECT 48.475 106.685 48.645 107.695 ;
        RECT 48.815 107.275 49.215 107.525 ;
        RECT 49.505 107.475 49.705 108.265 ;
        RECT 49.385 107.305 49.705 107.475 ;
        RECT 49.875 107.315 50.195 108.495 ;
        RECT 50.825 107.330 51.115 108.495 ;
        RECT 51.290 107.355 51.610 108.495 ;
        RECT 48.815 106.855 48.985 107.275 ;
        RECT 49.385 107.105 49.565 107.305 ;
        RECT 51.790 107.185 51.985 108.235 ;
        RECT 52.165 107.645 52.495 108.325 ;
        RECT 52.695 107.695 52.950 108.495 ;
        RECT 52.165 107.365 52.515 107.645 ;
        RECT 54.050 107.545 54.315 108.315 ;
        RECT 54.485 107.775 54.815 108.495 ;
        RECT 55.005 107.955 55.265 108.315 ;
        RECT 55.435 108.125 55.765 108.495 ;
        RECT 55.935 107.955 56.195 108.315 ;
        RECT 55.005 107.725 56.195 107.955 ;
        RECT 56.765 107.545 57.055 108.315 ;
        RECT 51.350 107.135 51.610 107.185 ;
        RECT 49.200 106.935 49.565 107.105 ;
        RECT 49.735 106.935 50.195 107.135 ;
        RECT 51.345 106.965 51.610 107.135 ;
        RECT 51.350 106.855 51.610 106.965 ;
        RECT 51.790 106.855 52.175 107.185 ;
        RECT 52.345 106.985 52.515 107.365 ;
        RECT 52.705 107.155 52.950 107.515 ;
        RECT 52.345 106.815 52.865 106.985 ;
        RECT 52.695 106.795 52.865 106.815 ;
        RECT 49.165 106.685 50.195 106.725 ;
        RECT 48.475 106.505 48.825 106.685 ;
        RECT 48.995 106.555 50.195 106.685 ;
        RECT 48.995 106.335 49.325 106.555 ;
        RECT 48.065 106.155 49.325 106.335 ;
        RECT 49.515 105.945 49.685 106.385 ;
        RECT 49.855 106.140 50.195 106.555 ;
        RECT 50.825 105.945 51.115 106.670 ;
        RECT 51.290 106.475 52.505 106.645 ;
        RECT 51.290 106.125 51.580 106.475 ;
        RECT 51.775 105.945 52.105 106.305 ;
        RECT 52.275 106.170 52.505 106.475 ;
        RECT 52.695 106.625 52.895 106.795 ;
        RECT 52.695 106.250 52.865 106.625 ;
        RECT 54.050 106.125 54.385 107.545 ;
        RECT 54.560 107.365 57.055 107.545 ;
        RECT 57.265 107.405 60.775 108.495 ;
        RECT 61.945 107.865 62.125 108.325 ;
        RECT 62.295 108.035 62.545 108.495 ;
        RECT 62.715 108.115 63.045 108.285 ;
        RECT 63.215 108.230 63.470 108.325 ;
        RECT 62.715 107.865 62.885 108.115 ;
        RECT 63.215 108.060 64.355 108.230 ;
        RECT 64.615 108.095 64.945 108.495 ;
        RECT 63.215 107.925 63.470 108.060 ;
        RECT 61.945 107.695 62.885 107.865 ;
        RECT 63.060 107.755 63.470 107.925 ;
        RECT 64.185 107.835 64.355 108.060 ;
        RECT 54.560 106.675 54.785 107.365 ;
        RECT 54.985 106.855 55.265 107.185 ;
        RECT 55.445 106.855 56.020 107.185 ;
        RECT 56.200 106.855 56.635 107.185 ;
        RECT 56.815 106.855 57.085 107.185 ;
        RECT 57.265 106.715 58.915 107.235 ;
        RECT 59.085 106.885 60.775 107.405 ;
        RECT 54.560 106.485 57.045 106.675 ;
        RECT 54.565 105.945 55.310 106.315 ;
        RECT 55.875 106.125 56.130 106.485 ;
        RECT 56.310 105.945 56.640 106.315 ;
        RECT 56.820 106.125 57.045 106.485 ;
        RECT 57.265 105.945 60.775 106.715 ;
        RECT 61.920 106.625 62.180 107.515 ;
        RECT 62.380 107.215 62.860 107.515 ;
        RECT 62.380 106.625 62.640 107.215 ;
        RECT 63.060 106.730 63.230 107.755 ;
        RECT 63.750 107.575 63.920 107.765 ;
        RECT 64.185 107.665 64.945 107.835 ;
        RECT 62.880 106.560 63.230 106.730 ;
        RECT 63.400 107.405 63.920 107.575 ;
        RECT 63.400 106.685 63.570 107.405 ;
        RECT 63.760 106.855 64.050 107.235 ;
        RECT 64.220 106.855 64.550 107.475 ;
        RECT 64.775 107.185 64.945 107.665 ;
        RECT 65.115 107.385 65.375 108.325 ;
        RECT 65.635 107.585 65.805 108.315 ;
        RECT 65.985 107.765 66.315 108.495 ;
        RECT 66.485 107.585 66.675 108.315 ;
        RECT 65.635 107.385 66.675 107.585 ;
        RECT 64.775 106.855 65.030 107.185 ;
        RECT 61.905 105.945 62.305 106.455 ;
        RECT 62.880 106.115 63.050 106.560 ;
        RECT 63.400 106.515 64.280 106.685 ;
        RECT 65.200 106.670 65.375 107.385 ;
        RECT 66.845 107.205 67.175 108.315 ;
        RECT 67.365 108.085 67.695 108.495 ;
        RECT 67.865 107.905 68.125 108.295 ;
        RECT 68.305 108.060 73.650 108.495 ;
        RECT 65.580 106.855 65.870 107.205 ;
        RECT 66.065 106.855 66.460 107.205 ;
        RECT 66.640 106.905 67.175 107.205 ;
        RECT 67.365 107.705 68.125 107.905 ;
        RECT 67.365 107.025 67.705 107.705 ;
        RECT 63.220 105.945 63.940 106.345 ;
        RECT 64.110 106.115 64.280 106.515 ;
        RECT 64.515 105.945 64.945 106.390 ;
        RECT 65.115 106.115 65.375 106.670 ;
        RECT 65.565 105.945 65.895 106.675 ;
        RECT 66.065 106.235 66.275 106.855 ;
        RECT 66.640 106.655 66.885 106.905 ;
        RECT 66.455 106.125 66.885 106.655 ;
        RECT 67.065 105.945 67.295 106.725 ;
        RECT 67.475 106.575 67.705 107.025 ;
        RECT 67.885 106.835 68.115 107.525 ;
        RECT 67.475 106.125 67.855 106.575 ;
        RECT 69.890 106.490 70.230 107.320 ;
        RECT 71.710 106.810 72.060 108.060 ;
        RECT 74.750 107.345 75.010 108.495 ;
        RECT 75.185 107.420 75.440 108.325 ;
        RECT 75.610 107.735 75.940 108.495 ;
        RECT 76.155 107.565 76.325 108.325 ;
        RECT 68.305 105.945 73.650 106.490 ;
        RECT 74.750 105.945 75.010 106.785 ;
        RECT 75.185 106.690 75.355 107.420 ;
        RECT 75.610 107.395 76.325 107.565 ;
        RECT 75.610 107.185 75.780 107.395 ;
        RECT 76.585 107.330 76.875 108.495 ;
        RECT 77.135 107.825 77.305 108.325 ;
        RECT 77.475 107.995 77.805 108.495 ;
        RECT 77.135 107.655 77.800 107.825 ;
        RECT 75.525 106.855 75.780 107.185 ;
        RECT 75.185 106.115 75.440 106.690 ;
        RECT 75.610 106.665 75.780 106.855 ;
        RECT 76.060 106.845 76.415 107.215 ;
        RECT 77.050 106.835 77.400 107.485 ;
        RECT 75.610 106.495 76.325 106.665 ;
        RECT 75.610 105.945 75.940 106.325 ;
        RECT 76.155 106.115 76.325 106.495 ;
        RECT 76.585 105.945 76.875 106.670 ;
        RECT 77.570 106.665 77.800 107.655 ;
        RECT 77.135 106.495 77.800 106.665 ;
        RECT 77.135 106.205 77.305 106.495 ;
        RECT 77.475 105.945 77.805 106.325 ;
        RECT 77.975 106.205 78.160 108.325 ;
        RECT 78.400 108.035 78.665 108.495 ;
        RECT 78.835 107.900 79.085 108.325 ;
        RECT 79.295 108.050 80.400 108.220 ;
        RECT 78.780 107.770 79.085 107.900 ;
        RECT 78.330 106.575 78.610 107.525 ;
        RECT 78.780 106.665 78.950 107.770 ;
        RECT 79.120 106.985 79.360 107.580 ;
        RECT 79.530 107.515 80.060 107.880 ;
        RECT 79.530 106.815 79.700 107.515 ;
        RECT 80.230 107.435 80.400 108.050 ;
        RECT 80.570 107.695 80.740 108.495 ;
        RECT 80.910 107.995 81.160 108.325 ;
        RECT 81.385 108.025 82.270 108.195 ;
        RECT 80.230 107.345 80.740 107.435 ;
        RECT 78.780 106.535 79.005 106.665 ;
        RECT 79.175 106.595 79.700 106.815 ;
        RECT 79.870 107.175 80.740 107.345 ;
        RECT 78.415 105.945 78.665 106.405 ;
        RECT 78.835 106.395 79.005 106.535 ;
        RECT 79.870 106.395 80.040 107.175 ;
        RECT 80.570 107.105 80.740 107.175 ;
        RECT 80.250 106.925 80.450 106.955 ;
        RECT 80.910 106.925 81.080 107.995 ;
        RECT 81.250 107.105 81.440 107.825 ;
        RECT 80.250 106.625 81.080 106.925 ;
        RECT 81.610 106.895 81.930 107.855 ;
        RECT 78.835 106.225 79.170 106.395 ;
        RECT 79.365 106.225 80.040 106.395 ;
        RECT 80.360 105.945 80.730 106.445 ;
        RECT 80.910 106.395 81.080 106.625 ;
        RECT 81.465 106.565 81.930 106.895 ;
        RECT 82.100 107.185 82.270 108.025 ;
        RECT 82.450 107.995 82.765 108.495 ;
        RECT 82.995 107.765 83.335 108.325 ;
        RECT 82.440 107.390 83.335 107.765 ;
        RECT 83.505 107.485 83.675 108.495 ;
        RECT 83.145 107.185 83.335 107.390 ;
        RECT 83.845 107.435 84.175 108.280 ;
        RECT 84.870 108.105 85.205 108.325 ;
        RECT 86.210 108.115 86.565 108.495 ;
        RECT 84.870 107.485 85.125 108.105 ;
        RECT 85.375 107.945 85.605 107.985 ;
        RECT 86.735 107.945 86.985 108.325 ;
        RECT 85.375 107.745 86.985 107.945 ;
        RECT 85.375 107.655 85.560 107.745 ;
        RECT 86.150 107.735 86.985 107.745 ;
        RECT 87.235 107.715 87.485 108.495 ;
        RECT 87.655 107.645 87.915 108.325 ;
        RECT 85.715 107.545 86.045 107.575 ;
        RECT 85.715 107.485 87.515 107.545 ;
        RECT 83.845 107.355 84.235 107.435 ;
        RECT 84.020 107.305 84.235 107.355 ;
        RECT 84.870 107.375 87.575 107.485 ;
        RECT 84.870 107.315 86.045 107.375 ;
        RECT 87.375 107.340 87.575 107.375 ;
        RECT 82.100 106.855 82.975 107.185 ;
        RECT 83.145 106.855 83.895 107.185 ;
        RECT 82.100 106.395 82.270 106.855 ;
        RECT 83.145 106.685 83.345 106.855 ;
        RECT 84.065 106.725 84.235 107.305 ;
        RECT 84.865 106.935 85.355 107.135 ;
        RECT 85.545 106.935 86.020 107.145 ;
        RECT 84.010 106.685 84.235 106.725 ;
        RECT 80.910 106.225 81.315 106.395 ;
        RECT 81.485 106.225 82.270 106.395 ;
        RECT 82.545 105.945 82.755 106.475 ;
        RECT 83.015 106.160 83.345 106.685 ;
        RECT 83.855 106.600 84.235 106.685 ;
        RECT 83.515 105.945 83.685 106.555 ;
        RECT 83.855 106.165 84.185 106.600 ;
        RECT 84.870 105.945 85.325 106.710 ;
        RECT 85.800 106.535 86.020 106.935 ;
        RECT 86.265 106.935 86.595 107.145 ;
        RECT 86.265 106.535 86.475 106.935 ;
        RECT 86.765 106.900 87.175 107.205 ;
        RECT 87.405 106.765 87.575 107.340 ;
        RECT 87.305 106.645 87.575 106.765 ;
        RECT 86.730 106.600 87.575 106.645 ;
        RECT 86.730 106.475 87.485 106.600 ;
        RECT 86.730 106.325 86.900 106.475 ;
        RECT 87.745 106.445 87.915 107.645 ;
        RECT 88.545 107.405 89.755 108.495 ;
        RECT 100.090 107.520 100.760 110.780 ;
        RECT 101.430 110.210 105.470 110.380 ;
        RECT 101.090 108.150 101.260 110.150 ;
        RECT 105.640 108.150 105.810 110.150 ;
        RECT 101.430 107.920 105.470 108.090 ;
        RECT 106.150 107.520 106.320 110.780 ;
        RECT 100.090 107.510 106.320 107.520 ;
        RECT 107.910 116.780 117.740 116.820 ;
        RECT 120.510 116.800 126.250 116.810 ;
        RECT 107.910 116.650 118.540 116.780 ;
        RECT 107.910 114.390 108.080 116.650 ;
        RECT 108.805 116.080 116.845 116.250 ;
        RECT 108.420 115.020 108.590 116.020 ;
        RECT 117.060 115.020 117.230 116.020 ;
        RECT 108.805 114.790 116.845 114.960 ;
        RECT 117.570 114.390 118.540 116.650 ;
        RECT 107.910 114.220 118.540 114.390 ;
        RECT 107.910 110.960 108.080 114.220 ;
        RECT 108.805 113.650 116.845 113.820 ;
        RECT 108.420 111.590 108.590 113.590 ;
        RECT 117.060 111.590 117.230 113.590 ;
        RECT 108.805 111.360 116.845 111.530 ;
        RECT 117.570 110.960 118.540 114.220 ;
        RECT 107.910 110.790 118.540 110.960 ;
        RECT 107.910 107.530 108.080 110.790 ;
        RECT 108.805 110.220 116.845 110.390 ;
        RECT 108.420 108.160 108.590 110.160 ;
        RECT 117.060 108.160 117.230 110.160 ;
        RECT 108.805 107.930 116.845 108.100 ;
        RECT 117.570 107.530 118.540 110.790 ;
        RECT 100.090 107.410 106.330 107.510 ;
        RECT 88.545 106.865 89.065 107.405 ;
        RECT 89.235 106.695 89.755 107.235 ;
        RECT 85.600 106.115 86.900 106.325 ;
        RECT 87.155 105.945 87.485 106.305 ;
        RECT 87.655 106.115 87.915 106.445 ;
        RECT 88.545 105.945 89.755 106.695 ;
        RECT 100.080 106.850 106.330 107.410 ;
        RECT 100.080 106.830 105.250 106.850 ;
        RECT 100.080 106.760 104.070 106.830 ;
        RECT 12.100 105.775 89.840 105.945 ;
        RECT 12.185 105.025 13.395 105.775 ;
        RECT 12.185 104.485 12.705 105.025 ;
        RECT 13.565 105.005 15.235 105.775 ;
        RECT 15.455 105.385 15.785 105.775 ;
        RECT 15.955 105.205 16.125 105.525 ;
        RECT 16.295 105.385 16.625 105.775 ;
        RECT 17.040 105.375 17.995 105.545 ;
        RECT 15.405 105.035 17.655 105.205 ;
        RECT 12.875 104.315 13.395 104.855 ;
        RECT 13.565 104.485 14.315 105.005 ;
        RECT 14.485 104.315 15.235 104.835 ;
        RECT 12.185 103.225 13.395 104.315 ;
        RECT 13.565 103.225 15.235 104.315 ;
        RECT 15.405 104.075 15.575 105.035 ;
        RECT 15.745 104.415 15.990 104.865 ;
        RECT 16.160 104.585 16.710 104.785 ;
        RECT 16.880 104.615 17.255 104.785 ;
        RECT 16.880 104.415 17.050 104.615 ;
        RECT 17.425 104.535 17.655 105.035 ;
        RECT 15.745 104.245 17.050 104.415 ;
        RECT 17.825 104.495 17.995 105.375 ;
        RECT 18.165 104.940 18.455 105.775 ;
        RECT 18.625 105.275 18.925 105.605 ;
        RECT 19.095 105.295 19.370 105.775 ;
        RECT 17.825 104.325 18.455 104.495 ;
        RECT 15.405 103.395 15.785 104.075 ;
        RECT 16.375 103.225 16.545 104.075 ;
        RECT 16.715 103.905 17.955 104.075 ;
        RECT 16.715 103.395 17.045 103.905 ;
        RECT 17.215 103.225 17.385 103.735 ;
        RECT 17.555 103.395 17.955 103.905 ;
        RECT 18.135 103.395 18.455 104.325 ;
        RECT 18.625 104.365 18.795 105.275 ;
        RECT 19.550 105.125 19.845 105.515 ;
        RECT 20.015 105.295 20.270 105.775 ;
        RECT 20.445 105.125 20.705 105.515 ;
        RECT 20.875 105.295 21.155 105.775 ;
        RECT 21.890 105.315 22.640 105.605 ;
        RECT 23.150 105.315 23.480 105.775 ;
        RECT 18.965 104.535 19.315 105.105 ;
        RECT 19.550 104.955 21.200 105.125 ;
        RECT 19.485 104.615 20.625 104.785 ;
        RECT 19.485 104.365 19.655 104.615 ;
        RECT 20.795 104.445 21.200 104.955 ;
        RECT 18.625 104.195 19.655 104.365 ;
        RECT 20.445 104.275 21.200 104.445 ;
        RECT 18.625 103.395 18.935 104.195 ;
        RECT 20.445 104.025 20.705 104.275 ;
        RECT 19.105 103.225 19.415 104.025 ;
        RECT 19.585 103.855 20.705 104.025 ;
        RECT 19.585 103.395 19.845 103.855 ;
        RECT 20.015 103.225 20.270 103.685 ;
        RECT 20.445 103.395 20.705 103.855 ;
        RECT 20.875 103.225 21.160 104.095 ;
        RECT 21.890 104.025 22.260 105.315 ;
        RECT 23.700 105.125 23.970 105.335 ;
        RECT 24.610 105.270 24.945 105.775 ;
        RECT 25.115 105.205 25.355 105.580 ;
        RECT 25.635 105.445 25.805 105.590 ;
        RECT 25.635 105.250 26.010 105.445 ;
        RECT 26.370 105.280 26.765 105.775 ;
        RECT 22.635 104.955 23.970 105.125 ;
        RECT 22.635 104.785 22.805 104.955 ;
        RECT 22.430 104.535 22.805 104.785 ;
        RECT 22.975 104.545 23.450 104.785 ;
        RECT 23.620 104.545 23.970 104.785 ;
        RECT 22.635 104.365 22.805 104.535 ;
        RECT 22.635 104.195 23.970 104.365 ;
        RECT 24.665 104.245 24.965 105.095 ;
        RECT 25.135 105.055 25.355 105.205 ;
        RECT 25.135 104.725 25.670 105.055 ;
        RECT 25.840 104.915 26.010 105.250 ;
        RECT 26.935 105.085 27.175 105.605 ;
        RECT 23.690 104.035 23.970 104.195 ;
        RECT 25.135 104.075 25.370 104.725 ;
        RECT 25.840 104.555 26.825 104.915 ;
        RECT 21.890 103.855 23.060 104.025 ;
        RECT 22.345 103.225 22.560 103.685 ;
        RECT 22.730 103.395 23.060 103.855 ;
        RECT 23.230 103.225 23.480 104.025 ;
        RECT 24.695 103.845 25.370 104.075 ;
        RECT 25.540 104.535 26.825 104.555 ;
        RECT 25.540 104.385 26.400 104.535 ;
        RECT 24.695 103.415 24.865 103.845 ;
        RECT 25.035 103.225 25.365 103.675 ;
        RECT 25.540 103.440 25.825 104.385 ;
        RECT 27.000 104.280 27.175 105.085 ;
        RECT 27.405 104.955 27.635 105.775 ;
        RECT 27.805 104.975 28.135 105.605 ;
        RECT 27.385 104.535 27.715 104.785 ;
        RECT 27.885 104.375 28.135 104.975 ;
        RECT 28.305 104.955 28.515 105.775 ;
        RECT 28.745 105.005 30.415 105.775 ;
        RECT 30.585 105.035 31.075 105.605 ;
        RECT 31.245 105.205 31.475 105.605 ;
        RECT 31.645 105.375 32.065 105.775 ;
        RECT 32.235 105.205 32.405 105.605 ;
        RECT 31.245 105.035 32.405 105.205 ;
        RECT 32.575 105.035 33.025 105.775 ;
        RECT 33.195 105.035 33.635 105.595 ;
        RECT 28.745 104.485 29.495 105.005 ;
        RECT 26.000 103.905 26.695 104.215 ;
        RECT 26.005 103.225 26.690 103.695 ;
        RECT 26.870 103.495 27.175 104.280 ;
        RECT 27.405 103.225 27.635 104.365 ;
        RECT 27.805 103.395 28.135 104.375 ;
        RECT 28.305 103.225 28.515 104.365 ;
        RECT 29.665 104.315 30.415 104.835 ;
        RECT 28.745 103.225 30.415 104.315 ;
        RECT 30.585 104.365 30.755 105.035 ;
        RECT 30.925 104.535 31.330 104.865 ;
        RECT 30.585 104.195 31.355 104.365 ;
        RECT 30.595 103.225 30.925 104.025 ;
        RECT 31.105 103.565 31.355 104.195 ;
        RECT 31.545 103.735 31.795 104.865 ;
        RECT 31.995 104.535 32.240 104.865 ;
        RECT 32.425 104.585 32.815 104.865 ;
        RECT 31.995 103.735 32.195 104.535 ;
        RECT 32.985 104.415 33.155 104.865 ;
        RECT 32.365 104.245 33.155 104.415 ;
        RECT 32.365 103.565 32.535 104.245 ;
        RECT 31.105 103.395 32.535 103.565 ;
        RECT 32.705 103.225 33.020 104.075 ;
        RECT 33.325 104.025 33.635 105.035 ;
        RECT 33.195 103.395 33.635 104.025 ;
        RECT 33.805 105.100 34.075 105.445 ;
        RECT 34.265 105.375 34.645 105.775 ;
        RECT 34.815 105.205 34.985 105.555 ;
        RECT 35.155 105.375 35.485 105.775 ;
        RECT 35.685 105.205 35.855 105.555 ;
        RECT 36.055 105.275 36.385 105.775 ;
        RECT 33.805 104.365 33.975 105.100 ;
        RECT 34.245 105.035 35.855 105.205 ;
        RECT 34.245 104.865 34.415 105.035 ;
        RECT 34.145 104.535 34.415 104.865 ;
        RECT 34.585 104.535 34.990 104.865 ;
        RECT 34.245 104.365 34.415 104.535 ;
        RECT 33.805 103.395 34.075 104.365 ;
        RECT 34.245 104.195 34.970 104.365 ;
        RECT 35.160 104.245 35.870 104.865 ;
        RECT 36.040 104.535 36.390 105.105 ;
        RECT 36.565 105.025 37.775 105.775 ;
        RECT 37.945 105.050 38.235 105.775 ;
        RECT 36.565 104.485 37.085 105.025 ;
        RECT 38.405 105.005 40.995 105.775 ;
        RECT 41.255 105.225 41.425 105.515 ;
        RECT 41.595 105.395 41.925 105.775 ;
        RECT 41.255 105.055 41.920 105.225 ;
        RECT 34.800 104.075 34.970 104.195 ;
        RECT 36.070 104.075 36.390 104.365 ;
        RECT 37.255 104.315 37.775 104.855 ;
        RECT 38.405 104.485 39.615 105.005 ;
        RECT 34.285 103.225 34.565 104.025 ;
        RECT 34.800 103.905 36.390 104.075 ;
        RECT 34.735 103.445 36.390 103.735 ;
        RECT 36.565 103.225 37.775 104.315 ;
        RECT 37.945 103.225 38.235 104.390 ;
        RECT 39.785 104.315 40.995 104.835 ;
        RECT 38.405 103.225 40.995 104.315 ;
        RECT 41.170 104.235 41.520 104.885 ;
        RECT 41.690 104.065 41.920 105.055 ;
        RECT 41.255 103.895 41.920 104.065 ;
        RECT 41.255 103.395 41.425 103.895 ;
        RECT 41.595 103.225 41.925 103.725 ;
        RECT 42.095 103.395 42.280 105.515 ;
        RECT 42.535 105.315 42.785 105.775 ;
        RECT 42.955 105.325 43.290 105.495 ;
        RECT 43.485 105.325 44.160 105.495 ;
        RECT 42.955 105.185 43.125 105.325 ;
        RECT 42.450 104.195 42.730 105.145 ;
        RECT 42.900 105.055 43.125 105.185 ;
        RECT 42.900 103.950 43.070 105.055 ;
        RECT 43.295 104.905 43.820 105.125 ;
        RECT 43.240 104.140 43.480 104.735 ;
        RECT 43.650 104.205 43.820 104.905 ;
        RECT 43.990 104.545 44.160 105.325 ;
        RECT 44.480 105.275 44.850 105.775 ;
        RECT 45.030 105.325 45.435 105.495 ;
        RECT 45.605 105.325 46.390 105.495 ;
        RECT 45.030 105.095 45.200 105.325 ;
        RECT 44.370 104.795 45.200 105.095 ;
        RECT 45.585 104.825 46.050 105.155 ;
        RECT 44.370 104.765 44.570 104.795 ;
        RECT 44.690 104.545 44.860 104.615 ;
        RECT 43.990 104.375 44.860 104.545 ;
        RECT 44.350 104.285 44.860 104.375 ;
        RECT 42.900 103.820 43.205 103.950 ;
        RECT 43.650 103.840 44.180 104.205 ;
        RECT 42.520 103.225 42.785 103.685 ;
        RECT 42.955 103.395 43.205 103.820 ;
        RECT 44.350 103.670 44.520 104.285 ;
        RECT 43.415 103.500 44.520 103.670 ;
        RECT 44.690 103.225 44.860 104.025 ;
        RECT 45.030 103.725 45.200 104.795 ;
        RECT 45.370 103.895 45.560 104.615 ;
        RECT 45.730 103.865 46.050 104.825 ;
        RECT 46.220 104.865 46.390 105.325 ;
        RECT 46.665 105.245 46.875 105.775 ;
        RECT 47.135 105.035 47.465 105.560 ;
        RECT 47.635 105.165 47.805 105.775 ;
        RECT 47.975 105.120 48.305 105.555 ;
        RECT 47.975 105.035 48.355 105.120 ;
        RECT 47.265 104.865 47.465 105.035 ;
        RECT 48.130 104.995 48.355 105.035 ;
        RECT 46.220 104.535 47.095 104.865 ;
        RECT 47.265 104.535 48.015 104.865 ;
        RECT 45.030 103.395 45.280 103.725 ;
        RECT 46.220 103.695 46.390 104.535 ;
        RECT 47.265 104.330 47.455 104.535 ;
        RECT 48.185 104.415 48.355 104.995 ;
        RECT 48.525 104.955 48.785 105.775 ;
        RECT 48.955 104.955 49.285 105.375 ;
        RECT 49.465 105.290 50.255 105.555 ;
        RECT 49.035 104.865 49.285 104.955 ;
        RECT 48.140 104.365 48.355 104.415 ;
        RECT 46.560 103.955 47.455 104.330 ;
        RECT 47.965 104.285 48.355 104.365 ;
        RECT 45.505 103.525 46.390 103.695 ;
        RECT 46.570 103.225 46.885 103.725 ;
        RECT 47.115 103.395 47.455 103.955 ;
        RECT 47.625 103.225 47.795 104.235 ;
        RECT 47.965 103.440 48.295 104.285 ;
        RECT 48.525 103.905 48.865 104.785 ;
        RECT 49.035 104.615 49.830 104.865 ;
        RECT 48.525 103.225 48.785 103.735 ;
        RECT 49.035 103.395 49.205 104.615 ;
        RECT 50.000 104.435 50.255 105.290 ;
        RECT 50.425 105.135 50.625 105.555 ;
        RECT 50.815 105.315 51.145 105.775 ;
        RECT 50.425 104.615 50.835 105.135 ;
        RECT 51.315 105.125 51.575 105.605 ;
        RECT 51.005 104.435 51.235 104.865 ;
        RECT 49.445 104.265 51.235 104.435 ;
        RECT 49.445 103.900 49.695 104.265 ;
        RECT 49.865 103.905 50.195 104.095 ;
        RECT 50.415 103.970 51.130 104.265 ;
        RECT 51.405 104.095 51.575 105.125 ;
        RECT 51.835 105.225 52.005 105.515 ;
        RECT 52.175 105.395 52.505 105.775 ;
        RECT 51.835 105.055 52.500 105.225 ;
        RECT 51.750 104.235 52.100 104.885 ;
        RECT 49.865 103.730 50.060 103.905 ;
        RECT 49.445 103.225 50.060 103.730 ;
        RECT 50.230 103.395 50.705 103.735 ;
        RECT 50.875 103.225 51.090 103.770 ;
        RECT 51.300 103.395 51.575 104.095 ;
        RECT 52.270 104.065 52.500 105.055 ;
        RECT 51.835 103.895 52.500 104.065 ;
        RECT 51.835 103.395 52.005 103.895 ;
        RECT 52.175 103.225 52.505 103.725 ;
        RECT 52.675 103.395 52.860 105.515 ;
        RECT 53.115 105.315 53.365 105.775 ;
        RECT 53.535 105.325 53.870 105.495 ;
        RECT 54.065 105.325 54.740 105.495 ;
        RECT 53.535 105.185 53.705 105.325 ;
        RECT 53.030 104.195 53.310 105.145 ;
        RECT 53.480 105.055 53.705 105.185 ;
        RECT 53.480 103.950 53.650 105.055 ;
        RECT 53.875 104.905 54.400 105.125 ;
        RECT 53.820 104.140 54.060 104.735 ;
        RECT 54.230 104.205 54.400 104.905 ;
        RECT 54.570 104.545 54.740 105.325 ;
        RECT 55.060 105.275 55.430 105.775 ;
        RECT 55.610 105.325 56.015 105.495 ;
        RECT 56.185 105.325 56.970 105.495 ;
        RECT 55.610 105.095 55.780 105.325 ;
        RECT 54.950 104.795 55.780 105.095 ;
        RECT 56.165 104.825 56.630 105.155 ;
        RECT 54.950 104.765 55.150 104.795 ;
        RECT 55.270 104.545 55.440 104.615 ;
        RECT 54.570 104.375 55.440 104.545 ;
        RECT 54.930 104.285 55.440 104.375 ;
        RECT 53.480 103.820 53.785 103.950 ;
        RECT 54.230 103.840 54.760 104.205 ;
        RECT 53.100 103.225 53.365 103.685 ;
        RECT 53.535 103.395 53.785 103.820 ;
        RECT 54.930 103.670 55.100 104.285 ;
        RECT 53.995 103.500 55.100 103.670 ;
        RECT 55.270 103.225 55.440 104.025 ;
        RECT 55.610 103.725 55.780 104.795 ;
        RECT 55.950 103.895 56.140 104.615 ;
        RECT 56.310 103.865 56.630 104.825 ;
        RECT 56.800 104.865 56.970 105.325 ;
        RECT 57.245 105.245 57.455 105.775 ;
        RECT 57.715 105.035 58.045 105.560 ;
        RECT 58.215 105.165 58.385 105.775 ;
        RECT 58.555 105.120 58.885 105.555 ;
        RECT 58.555 105.035 58.935 105.120 ;
        RECT 57.845 104.865 58.045 105.035 ;
        RECT 58.710 104.995 58.935 105.035 ;
        RECT 56.800 104.535 57.675 104.865 ;
        RECT 57.845 104.535 58.595 104.865 ;
        RECT 55.610 103.395 55.860 103.725 ;
        RECT 56.800 103.695 56.970 104.535 ;
        RECT 57.845 104.330 58.035 104.535 ;
        RECT 58.765 104.415 58.935 104.995 ;
        RECT 59.575 104.965 59.845 105.775 ;
        RECT 60.015 104.965 60.345 105.605 ;
        RECT 60.515 104.965 60.755 105.775 ;
        RECT 59.565 104.535 59.915 104.785 ;
        RECT 58.720 104.365 58.935 104.415 ;
        RECT 60.085 104.365 60.255 104.965 ;
        RECT 60.425 104.535 60.775 104.785 ;
        RECT 57.140 103.955 58.035 104.330 ;
        RECT 58.545 104.285 58.935 104.365 ;
        RECT 56.085 103.525 56.970 103.695 ;
        RECT 57.150 103.225 57.465 103.725 ;
        RECT 57.695 103.395 58.035 103.955 ;
        RECT 58.205 103.225 58.375 104.235 ;
        RECT 58.545 103.440 58.875 104.285 ;
        RECT 59.575 103.225 59.905 104.365 ;
        RECT 60.085 104.195 60.765 104.365 ;
        RECT 60.435 103.410 60.765 104.195 ;
        RECT 60.955 103.405 61.215 105.595 ;
        RECT 61.475 105.405 62.145 105.775 ;
        RECT 62.325 105.225 62.635 105.595 ;
        RECT 61.405 105.025 62.635 105.225 ;
        RECT 61.405 104.355 61.695 105.025 ;
        RECT 62.815 104.845 63.045 105.485 ;
        RECT 63.225 105.045 63.515 105.775 ;
        RECT 63.705 105.050 63.995 105.775 ;
        RECT 64.165 104.975 64.860 105.605 ;
        RECT 65.065 104.975 65.375 105.775 ;
        RECT 66.010 105.010 66.465 105.775 ;
        RECT 66.740 105.395 68.040 105.605 ;
        RECT 68.295 105.415 68.625 105.775 ;
        RECT 67.870 105.245 68.040 105.395 ;
        RECT 68.795 105.275 69.055 105.605 ;
        RECT 68.825 105.265 69.055 105.275 ;
        RECT 61.875 104.535 62.340 104.845 ;
        RECT 62.520 104.535 63.045 104.845 ;
        RECT 63.225 104.535 63.525 104.865 ;
        RECT 64.185 104.535 64.520 104.785 ;
        RECT 61.405 104.135 62.175 104.355 ;
        RECT 61.385 103.225 61.725 103.955 ;
        RECT 61.905 103.405 62.175 104.135 ;
        RECT 62.355 104.115 63.515 104.355 ;
        RECT 62.355 103.405 62.585 104.115 ;
        RECT 62.755 103.225 63.085 103.935 ;
        RECT 63.255 103.405 63.515 104.115 ;
        RECT 63.705 103.225 63.995 104.390 ;
        RECT 64.690 104.375 64.860 104.975 ;
        RECT 65.030 104.535 65.365 104.805 ;
        RECT 66.940 104.785 67.160 105.185 ;
        RECT 66.005 104.585 66.495 104.785 ;
        RECT 66.685 104.575 67.160 104.785 ;
        RECT 67.405 104.785 67.615 105.185 ;
        RECT 67.870 105.120 68.625 105.245 ;
        RECT 67.870 105.075 68.715 105.120 ;
        RECT 68.445 104.955 68.715 105.075 ;
        RECT 67.405 104.575 67.735 104.785 ;
        RECT 67.905 104.515 68.315 104.820 ;
        RECT 64.165 103.225 64.425 104.365 ;
        RECT 64.595 103.395 64.925 104.375 ;
        RECT 65.095 103.225 65.375 104.365 ;
        RECT 66.010 104.345 67.185 104.405 ;
        RECT 68.545 104.380 68.715 104.955 ;
        RECT 68.515 104.345 68.715 104.380 ;
        RECT 66.010 104.235 68.715 104.345 ;
        RECT 66.010 103.615 66.265 104.235 ;
        RECT 66.855 104.175 68.655 104.235 ;
        RECT 66.855 104.145 67.185 104.175 ;
        RECT 68.885 104.075 69.055 105.265 ;
        RECT 66.515 103.975 66.700 104.065 ;
        RECT 67.290 103.975 68.125 103.985 ;
        RECT 66.515 103.775 68.125 103.975 ;
        RECT 66.515 103.735 66.745 103.775 ;
        RECT 66.010 103.395 66.345 103.615 ;
        RECT 67.350 103.225 67.705 103.605 ;
        RECT 67.875 103.395 68.125 103.775 ;
        RECT 68.375 103.225 68.625 104.005 ;
        RECT 68.795 103.395 69.055 104.075 ;
        RECT 69.230 105.035 69.485 105.605 ;
        RECT 69.655 105.375 69.985 105.775 ;
        RECT 70.410 105.240 70.940 105.605 ;
        RECT 70.410 105.205 70.585 105.240 ;
        RECT 69.655 105.035 70.585 105.205 ;
        RECT 69.230 104.365 69.400 105.035 ;
        RECT 69.655 104.865 69.825 105.035 ;
        RECT 69.570 104.535 69.825 104.865 ;
        RECT 70.050 104.535 70.245 104.865 ;
        RECT 69.230 103.395 69.565 104.365 ;
        RECT 69.735 103.225 69.905 104.365 ;
        RECT 70.075 103.565 70.245 104.535 ;
        RECT 70.415 103.905 70.585 105.035 ;
        RECT 70.755 104.245 70.925 105.045 ;
        RECT 71.130 104.755 71.405 105.605 ;
        RECT 71.125 104.585 71.405 104.755 ;
        RECT 71.130 104.445 71.405 104.585 ;
        RECT 71.575 104.245 71.765 105.605 ;
        RECT 71.945 105.240 72.455 105.775 ;
        RECT 72.675 104.965 72.920 105.570 ;
        RECT 73.365 105.035 73.750 105.605 ;
        RECT 73.920 105.315 74.245 105.775 ;
        RECT 74.765 105.145 75.045 105.605 ;
        RECT 71.965 104.795 73.195 104.965 ;
        RECT 70.755 104.075 71.765 104.245 ;
        RECT 71.935 104.230 72.685 104.420 ;
        RECT 70.415 103.735 71.540 103.905 ;
        RECT 71.935 103.565 72.105 104.230 ;
        RECT 72.855 103.985 73.195 104.795 ;
        RECT 70.075 103.395 72.105 103.565 ;
        RECT 72.275 103.225 72.445 103.985 ;
        RECT 72.680 103.575 73.195 103.985 ;
        RECT 73.365 104.365 73.645 105.035 ;
        RECT 73.920 104.975 75.045 105.145 ;
        RECT 73.920 104.865 74.370 104.975 ;
        RECT 73.815 104.535 74.370 104.865 ;
        RECT 75.235 104.805 75.635 105.605 ;
        RECT 76.035 105.315 76.305 105.775 ;
        RECT 76.475 105.145 76.760 105.605 ;
        RECT 73.365 103.395 73.750 104.365 ;
        RECT 73.920 104.075 74.370 104.535 ;
        RECT 74.540 104.245 75.635 104.805 ;
        RECT 73.920 103.855 75.045 104.075 ;
        RECT 73.920 103.225 74.245 103.685 ;
        RECT 74.765 103.395 75.045 103.855 ;
        RECT 75.235 103.395 75.635 104.245 ;
        RECT 75.805 104.975 76.760 105.145 ;
        RECT 77.045 104.975 77.385 105.605 ;
        RECT 77.555 104.975 77.805 105.775 ;
        RECT 77.995 105.125 78.325 105.605 ;
        RECT 78.495 105.315 78.720 105.775 ;
        RECT 78.890 105.125 79.220 105.605 ;
        RECT 75.805 104.075 76.015 104.975 ;
        RECT 76.185 104.245 76.875 104.805 ;
        RECT 77.045 104.365 77.220 104.975 ;
        RECT 77.995 104.955 79.220 105.125 ;
        RECT 79.850 104.995 80.350 105.605 ;
        RECT 81.275 105.225 81.445 105.515 ;
        RECT 81.615 105.395 81.945 105.775 ;
        RECT 81.275 105.055 81.940 105.225 ;
        RECT 77.390 104.615 78.085 104.785 ;
        RECT 77.915 104.365 78.085 104.615 ;
        RECT 78.260 104.585 78.680 104.785 ;
        RECT 78.850 104.585 79.180 104.785 ;
        RECT 79.350 104.585 79.680 104.785 ;
        RECT 79.850 104.365 80.020 104.995 ;
        RECT 80.205 104.535 80.555 104.785 ;
        RECT 75.805 103.855 76.760 104.075 ;
        RECT 76.035 103.225 76.305 103.685 ;
        RECT 76.475 103.395 76.760 103.855 ;
        RECT 77.045 103.395 77.385 104.365 ;
        RECT 77.555 103.225 77.725 104.365 ;
        RECT 77.915 104.195 80.350 104.365 ;
        RECT 81.190 104.235 81.540 104.885 ;
        RECT 77.995 103.225 78.245 104.025 ;
        RECT 78.890 103.395 79.220 104.195 ;
        RECT 79.520 103.225 79.850 104.025 ;
        RECT 80.020 103.395 80.350 104.195 ;
        RECT 81.710 104.065 81.940 105.055 ;
        RECT 81.275 103.895 81.940 104.065 ;
        RECT 81.275 103.395 81.445 103.895 ;
        RECT 81.615 103.225 81.945 103.725 ;
        RECT 82.115 103.395 82.300 105.515 ;
        RECT 82.555 105.315 82.805 105.775 ;
        RECT 82.975 105.325 83.310 105.495 ;
        RECT 83.505 105.325 84.180 105.495 ;
        RECT 82.975 105.185 83.145 105.325 ;
        RECT 82.470 104.195 82.750 105.145 ;
        RECT 82.920 105.055 83.145 105.185 ;
        RECT 82.920 103.950 83.090 105.055 ;
        RECT 83.315 104.905 83.840 105.125 ;
        RECT 83.260 104.140 83.500 104.735 ;
        RECT 83.670 104.205 83.840 104.905 ;
        RECT 84.010 104.545 84.180 105.325 ;
        RECT 84.500 105.275 84.870 105.775 ;
        RECT 85.050 105.325 85.455 105.495 ;
        RECT 85.625 105.325 86.410 105.495 ;
        RECT 85.050 105.095 85.220 105.325 ;
        RECT 84.390 104.795 85.220 105.095 ;
        RECT 85.605 104.825 86.070 105.155 ;
        RECT 84.390 104.765 84.590 104.795 ;
        RECT 84.710 104.545 84.880 104.615 ;
        RECT 84.010 104.375 84.880 104.545 ;
        RECT 84.370 104.285 84.880 104.375 ;
        RECT 82.920 103.820 83.225 103.950 ;
        RECT 83.670 103.840 84.200 104.205 ;
        RECT 82.540 103.225 82.805 103.685 ;
        RECT 82.975 103.395 83.225 103.820 ;
        RECT 84.370 103.670 84.540 104.285 ;
        RECT 83.435 103.500 84.540 103.670 ;
        RECT 84.710 103.225 84.880 104.025 ;
        RECT 85.050 103.725 85.220 104.795 ;
        RECT 85.390 103.895 85.580 104.615 ;
        RECT 85.750 103.865 86.070 104.825 ;
        RECT 86.240 104.865 86.410 105.325 ;
        RECT 86.685 105.245 86.895 105.775 ;
        RECT 87.155 105.035 87.485 105.560 ;
        RECT 87.655 105.165 87.825 105.775 ;
        RECT 87.995 105.120 88.325 105.555 ;
        RECT 87.995 105.035 88.375 105.120 ;
        RECT 87.285 104.865 87.485 105.035 ;
        RECT 88.150 104.995 88.375 105.035 ;
        RECT 88.545 105.025 89.755 105.775 ;
        RECT 100.080 105.490 102.000 106.760 ;
        RECT 103.510 106.750 104.070 106.760 ;
        RECT 103.740 105.660 104.070 106.750 ;
        RECT 104.440 106.280 105.480 106.450 ;
        RECT 104.440 105.840 105.480 106.010 ;
        RECT 105.650 105.980 105.820 106.310 ;
        RECT 103.900 105.440 104.070 105.660 ;
        RECT 106.160 105.440 106.330 106.850 ;
        RECT 103.900 105.270 106.330 105.440 ;
        RECT 107.910 107.360 118.540 107.530 ;
        RECT 120.020 116.640 126.250 116.800 ;
        RECT 120.020 114.380 120.690 116.640 ;
        RECT 121.360 116.070 125.400 116.240 ;
        RECT 121.020 115.010 121.190 116.010 ;
        RECT 125.570 115.010 125.740 116.010 ;
        RECT 121.360 114.780 125.400 114.950 ;
        RECT 126.080 114.380 126.250 116.640 ;
        RECT 120.020 114.210 126.250 114.380 ;
        RECT 120.020 110.950 120.690 114.210 ;
        RECT 121.360 113.640 125.400 113.810 ;
        RECT 121.020 111.580 121.190 113.580 ;
        RECT 125.570 111.580 125.740 113.580 ;
        RECT 121.360 111.350 125.400 111.520 ;
        RECT 126.080 110.950 126.250 114.210 ;
        RECT 120.020 110.780 126.250 110.950 ;
        RECT 120.020 107.520 120.690 110.780 ;
        RECT 121.360 110.210 125.400 110.380 ;
        RECT 121.020 108.150 121.190 110.150 ;
        RECT 125.570 108.150 125.740 110.150 ;
        RECT 121.360 107.920 125.400 108.090 ;
        RECT 126.080 107.520 126.250 110.780 ;
        RECT 120.020 107.510 126.250 107.520 ;
        RECT 127.840 116.780 137.670 116.820 ;
        RECT 140.540 116.800 146.280 116.810 ;
        RECT 127.840 116.650 138.470 116.780 ;
        RECT 127.840 114.390 128.010 116.650 ;
        RECT 128.735 116.080 136.775 116.250 ;
        RECT 128.350 115.020 128.520 116.020 ;
        RECT 136.990 115.020 137.160 116.020 ;
        RECT 128.735 114.790 136.775 114.960 ;
        RECT 137.500 114.390 138.470 116.650 ;
        RECT 127.840 114.220 138.470 114.390 ;
        RECT 127.840 110.960 128.010 114.220 ;
        RECT 128.735 113.650 136.775 113.820 ;
        RECT 128.350 111.590 128.520 113.590 ;
        RECT 136.990 111.590 137.160 113.590 ;
        RECT 128.735 111.360 136.775 111.530 ;
        RECT 137.500 110.960 138.470 114.220 ;
        RECT 127.840 110.790 138.470 110.960 ;
        RECT 127.840 107.530 128.010 110.790 ;
        RECT 128.735 110.220 136.775 110.390 ;
        RECT 128.350 108.160 128.520 110.160 ;
        RECT 136.990 108.160 137.160 110.160 ;
        RECT 128.735 107.930 136.775 108.100 ;
        RECT 137.500 107.530 138.470 110.790 ;
        RECT 120.020 107.410 126.260 107.510 ;
        RECT 107.910 105.100 108.080 107.360 ;
        RECT 108.805 106.790 116.845 106.960 ;
        RECT 108.420 105.730 108.590 106.730 ;
        RECT 117.060 105.730 117.230 106.730 ;
        RECT 108.805 105.500 116.845 105.670 ;
        RECT 117.570 105.100 118.540 107.360 ;
        RECT 120.010 106.850 126.260 107.410 ;
        RECT 120.010 106.830 125.180 106.850 ;
        RECT 120.010 106.760 124.000 106.830 ;
        RECT 120.010 106.250 121.930 106.760 ;
        RECT 123.440 106.750 124.000 106.760 ;
        RECT 107.910 105.070 118.540 105.100 ;
        RECT 86.240 104.535 87.115 104.865 ;
        RECT 87.285 104.535 88.035 104.865 ;
        RECT 85.050 103.395 85.300 103.725 ;
        RECT 86.240 103.695 86.410 104.535 ;
        RECT 87.285 104.330 87.475 104.535 ;
        RECT 88.205 104.415 88.375 104.995 ;
        RECT 88.160 104.365 88.375 104.415 ;
        RECT 86.580 103.955 87.475 104.330 ;
        RECT 87.985 104.285 88.375 104.365 ;
        RECT 88.545 104.315 89.065 104.855 ;
        RECT 89.235 104.485 89.755 105.025 ;
        RECT 107.880 104.960 118.540 105.070 ;
        RECT 106.130 104.910 118.540 104.960 ;
        RECT 101.790 104.740 118.540 104.910 ;
        RECT 85.525 103.525 86.410 103.695 ;
        RECT 86.590 103.225 86.905 103.725 ;
        RECT 87.135 103.395 87.475 103.955 ;
        RECT 87.645 103.225 87.815 104.235 ;
        RECT 87.985 103.440 88.315 104.285 ;
        RECT 88.545 103.225 89.755 104.315 ;
        RECT 101.790 103.330 101.960 104.740 ;
        RECT 102.330 104.170 105.370 104.340 ;
        RECT 102.330 103.730 105.370 103.900 ;
        RECT 105.585 103.870 105.755 104.200 ;
        RECT 106.090 103.980 118.540 104.740 ;
        RECT 120.000 105.490 121.930 106.250 ;
        RECT 123.670 105.660 124.000 106.750 ;
        RECT 124.370 106.280 125.410 106.450 ;
        RECT 124.370 105.840 125.410 106.010 ;
        RECT 125.580 105.980 125.750 106.310 ;
        RECT 106.090 103.970 118.430 103.980 ;
        RECT 106.090 103.960 111.970 103.970 ;
        RECT 106.090 103.940 106.660 103.960 ;
        RECT 107.880 103.950 111.970 103.960 ;
        RECT 106.100 103.330 106.270 103.940 ;
        RECT 12.100 103.055 89.840 103.225 ;
        RECT 101.790 103.160 106.270 103.330 ;
        RECT 12.185 101.965 13.395 103.055 ;
        RECT 13.565 102.620 18.910 103.055 ;
        RECT 19.085 102.620 24.430 103.055 ;
        RECT 12.185 101.255 12.705 101.795 ;
        RECT 12.875 101.425 13.395 101.965 ;
        RECT 12.185 100.505 13.395 101.255 ;
        RECT 15.150 101.050 15.490 101.880 ;
        RECT 16.970 101.370 17.320 102.620 ;
        RECT 20.670 101.050 21.010 101.880 ;
        RECT 22.490 101.370 22.840 102.620 ;
        RECT 25.065 101.890 25.355 103.055 ;
        RECT 25.525 102.620 30.870 103.055 ;
        RECT 13.565 100.505 18.910 101.050 ;
        RECT 19.085 100.505 24.430 101.050 ;
        RECT 25.065 100.505 25.355 101.230 ;
        RECT 27.110 101.050 27.450 101.880 ;
        RECT 28.930 101.370 29.280 102.620 ;
        RECT 31.045 101.965 34.555 103.055 ;
        RECT 34.725 101.965 35.935 103.055 ;
        RECT 31.045 101.275 32.695 101.795 ;
        RECT 32.865 101.445 34.555 101.965 ;
        RECT 25.525 100.505 30.870 101.050 ;
        RECT 31.045 100.505 34.555 101.275 ;
        RECT 34.725 101.255 35.245 101.795 ;
        RECT 35.415 101.425 35.935 101.965 ;
        RECT 36.115 101.915 36.445 103.055 ;
        RECT 36.975 102.085 37.305 102.870 ;
        RECT 37.600 102.425 37.885 102.885 ;
        RECT 38.055 102.595 38.325 103.055 ;
        RECT 37.600 102.205 38.555 102.425 ;
        RECT 36.625 101.915 37.305 102.085 ;
        RECT 36.105 101.495 36.455 101.745 ;
        RECT 36.625 101.315 36.795 101.915 ;
        RECT 36.965 101.495 37.315 101.745 ;
        RECT 37.485 101.475 38.175 102.035 ;
        RECT 34.725 100.505 35.935 101.255 ;
        RECT 36.115 100.505 36.385 101.315 ;
        RECT 36.555 100.675 36.885 101.315 ;
        RECT 37.055 100.505 37.295 101.315 ;
        RECT 38.345 101.305 38.555 102.205 ;
        RECT 37.600 101.135 38.555 101.305 ;
        RECT 38.725 102.035 39.125 102.885 ;
        RECT 39.315 102.425 39.595 102.885 ;
        RECT 40.115 102.595 40.440 103.055 ;
        RECT 39.315 102.205 40.440 102.425 ;
        RECT 38.725 101.475 39.820 102.035 ;
        RECT 39.990 101.745 40.440 102.205 ;
        RECT 40.610 101.915 40.995 102.885 ;
        RECT 41.225 101.995 41.555 102.840 ;
        RECT 41.725 102.045 41.895 103.055 ;
        RECT 42.065 102.325 42.405 102.885 ;
        RECT 42.635 102.555 42.950 103.055 ;
        RECT 43.130 102.585 44.015 102.755 ;
        RECT 37.600 100.675 37.885 101.135 ;
        RECT 38.055 100.505 38.325 100.965 ;
        RECT 38.725 100.675 39.125 101.475 ;
        RECT 39.990 101.415 40.545 101.745 ;
        RECT 39.990 101.305 40.440 101.415 ;
        RECT 39.315 101.135 40.440 101.305 ;
        RECT 40.715 101.245 40.995 101.915 ;
        RECT 39.315 100.675 39.595 101.135 ;
        RECT 40.115 100.505 40.440 100.965 ;
        RECT 40.610 100.675 40.995 101.245 ;
        RECT 41.165 101.915 41.555 101.995 ;
        RECT 42.065 101.950 42.960 102.325 ;
        RECT 41.165 101.865 41.380 101.915 ;
        RECT 41.165 101.285 41.335 101.865 ;
        RECT 42.065 101.745 42.255 101.950 ;
        RECT 43.130 101.745 43.300 102.585 ;
        RECT 44.240 102.555 44.490 102.885 ;
        RECT 41.505 101.415 42.255 101.745 ;
        RECT 42.425 101.415 43.300 101.745 ;
        RECT 41.165 101.245 41.390 101.285 ;
        RECT 42.055 101.245 42.255 101.415 ;
        RECT 41.165 101.160 41.545 101.245 ;
        RECT 41.215 100.725 41.545 101.160 ;
        RECT 41.715 100.505 41.885 101.115 ;
        RECT 42.055 100.720 42.385 101.245 ;
        RECT 42.645 100.505 42.855 101.035 ;
        RECT 43.130 100.955 43.300 101.415 ;
        RECT 43.470 101.455 43.790 102.415 ;
        RECT 43.960 101.665 44.150 102.385 ;
        RECT 44.320 101.485 44.490 102.555 ;
        RECT 44.660 102.255 44.830 103.055 ;
        RECT 45.000 102.610 46.105 102.780 ;
        RECT 45.000 101.995 45.170 102.610 ;
        RECT 46.315 102.460 46.565 102.885 ;
        RECT 46.735 102.595 47.000 103.055 ;
        RECT 45.340 102.075 45.870 102.440 ;
        RECT 46.315 102.330 46.620 102.460 ;
        RECT 44.660 101.905 45.170 101.995 ;
        RECT 44.660 101.735 45.530 101.905 ;
        RECT 44.660 101.665 44.830 101.735 ;
        RECT 44.950 101.485 45.150 101.515 ;
        RECT 43.470 101.125 43.935 101.455 ;
        RECT 44.320 101.185 45.150 101.485 ;
        RECT 44.320 100.955 44.490 101.185 ;
        RECT 43.130 100.785 43.915 100.955 ;
        RECT 44.085 100.785 44.490 100.955 ;
        RECT 44.670 100.505 45.040 101.005 ;
        RECT 45.360 100.955 45.530 101.735 ;
        RECT 45.700 101.375 45.870 102.075 ;
        RECT 46.040 101.545 46.280 102.140 ;
        RECT 45.700 101.155 46.225 101.375 ;
        RECT 46.450 101.225 46.620 102.330 ;
        RECT 46.395 101.095 46.620 101.225 ;
        RECT 46.790 101.135 47.070 102.085 ;
        RECT 46.395 100.955 46.565 101.095 ;
        RECT 45.360 100.785 46.035 100.955 ;
        RECT 46.230 100.785 46.565 100.955 ;
        RECT 46.735 100.505 46.985 100.965 ;
        RECT 47.240 100.765 47.425 102.885 ;
        RECT 47.595 102.555 47.925 103.055 ;
        RECT 48.095 102.385 48.265 102.885 ;
        RECT 47.600 102.215 48.265 102.385 ;
        RECT 48.630 102.255 48.885 103.055 ;
        RECT 47.600 101.225 47.830 102.215 ;
        RECT 49.055 102.085 49.385 102.885 ;
        RECT 49.555 102.255 49.725 103.055 ;
        RECT 49.895 102.085 50.225 102.885 ;
        RECT 48.000 101.395 48.350 102.045 ;
        RECT 48.525 101.915 50.225 102.085 ;
        RECT 50.395 101.915 50.655 103.055 ;
        RECT 48.525 101.325 48.805 101.915 ;
        RECT 50.825 101.890 51.115 103.055 ;
        RECT 51.285 101.915 51.545 102.885 ;
        RECT 51.740 102.645 52.070 103.055 ;
        RECT 52.270 102.465 52.440 102.885 ;
        RECT 52.655 102.645 53.325 103.055 ;
        RECT 53.560 102.465 53.730 102.885 ;
        RECT 54.035 102.615 54.365 103.055 ;
        RECT 51.715 102.295 53.730 102.465 ;
        RECT 54.535 102.435 54.710 102.885 ;
        RECT 48.975 101.495 49.725 101.745 ;
        RECT 49.895 101.495 50.655 101.745 ;
        RECT 47.600 101.055 48.265 101.225 ;
        RECT 48.525 101.075 49.385 101.325 ;
        RECT 49.555 101.135 50.655 101.305 ;
        RECT 47.595 100.505 47.925 100.885 ;
        RECT 48.095 100.765 48.265 101.055 ;
        RECT 48.635 100.885 48.965 100.905 ;
        RECT 49.555 100.885 49.805 101.135 ;
        RECT 48.635 100.675 49.805 100.885 ;
        RECT 49.975 100.505 50.145 100.965 ;
        RECT 50.315 100.675 50.655 101.135 ;
        RECT 50.825 100.505 51.115 101.230 ;
        RECT 51.285 101.225 51.455 101.915 ;
        RECT 51.715 101.745 51.885 102.295 ;
        RECT 51.625 101.415 51.885 101.745 ;
        RECT 51.285 100.760 51.625 101.225 ;
        RECT 52.055 101.085 52.395 102.115 ;
        RECT 52.585 101.015 52.855 102.115 ;
        RECT 51.290 100.715 51.625 100.760 ;
        RECT 51.795 100.505 52.125 100.885 ;
        RECT 52.585 100.845 52.895 101.015 ;
        RECT 52.585 100.840 52.855 100.845 ;
        RECT 53.080 100.840 53.360 102.115 ;
        RECT 53.560 101.005 53.730 102.295 ;
        RECT 54.080 102.265 54.710 102.435 ;
        RECT 55.055 102.435 55.225 102.865 ;
        RECT 55.395 102.605 55.725 103.055 ;
        RECT 54.080 101.745 54.250 102.265 ;
        RECT 55.055 102.205 55.730 102.435 ;
        RECT 53.900 101.415 54.250 101.745 ;
        RECT 54.430 101.415 54.795 102.095 ;
        RECT 54.080 101.245 54.250 101.415 ;
        RECT 54.080 101.075 54.710 101.245 ;
        RECT 55.025 101.185 55.325 102.035 ;
        RECT 55.495 101.555 55.730 102.205 ;
        RECT 55.900 101.895 56.185 102.840 ;
        RECT 56.365 102.585 57.050 103.055 ;
        RECT 56.360 102.065 57.055 102.375 ;
        RECT 57.230 102.000 57.535 102.785 ;
        RECT 57.815 102.435 57.985 102.865 ;
        RECT 58.155 102.605 58.485 103.055 ;
        RECT 57.815 102.205 58.490 102.435 ;
        RECT 55.900 101.745 56.760 101.895 ;
        RECT 55.900 101.725 57.185 101.745 ;
        RECT 55.495 101.225 56.030 101.555 ;
        RECT 56.200 101.365 57.185 101.725 ;
        RECT 55.495 101.075 55.715 101.225 ;
        RECT 53.560 100.675 53.790 101.005 ;
        RECT 54.035 100.505 54.365 100.885 ;
        RECT 54.535 100.675 54.710 101.075 ;
        RECT 54.970 100.505 55.305 101.010 ;
        RECT 55.475 100.700 55.715 101.075 ;
        RECT 56.200 101.030 56.370 101.365 ;
        RECT 57.360 101.195 57.535 102.000 ;
        RECT 55.995 100.835 56.370 101.030 ;
        RECT 55.995 100.690 56.165 100.835 ;
        RECT 56.730 100.505 57.125 101.000 ;
        RECT 57.295 100.675 57.535 101.195 ;
        RECT 57.785 101.185 58.085 102.035 ;
        RECT 58.255 101.555 58.490 102.205 ;
        RECT 58.660 101.895 58.945 102.840 ;
        RECT 59.125 102.585 59.810 103.055 ;
        RECT 59.120 102.065 59.815 102.375 ;
        RECT 59.990 102.000 60.295 102.785 ;
        RECT 58.660 101.745 59.520 101.895 ;
        RECT 58.660 101.725 59.945 101.745 ;
        RECT 58.255 101.225 58.790 101.555 ;
        RECT 58.960 101.365 59.945 101.725 ;
        RECT 58.255 101.075 58.475 101.225 ;
        RECT 57.730 100.505 58.065 101.010 ;
        RECT 58.235 100.700 58.475 101.075 ;
        RECT 58.960 101.030 59.130 101.365 ;
        RECT 60.120 101.195 60.295 102.000 ;
        RECT 61.560 102.045 61.860 102.885 ;
        RECT 62.055 102.215 62.305 103.055 ;
        RECT 62.895 102.465 63.700 102.885 ;
        RECT 62.475 102.295 64.040 102.465 ;
        RECT 62.475 102.045 62.645 102.295 ;
        RECT 61.560 101.875 62.645 102.045 ;
        RECT 61.405 101.415 61.735 101.705 ;
        RECT 61.905 101.245 62.075 101.875 ;
        RECT 62.815 101.745 63.135 102.125 ;
        RECT 63.325 102.035 63.700 102.125 ;
        RECT 63.305 101.865 63.700 102.035 ;
        RECT 63.870 102.045 64.040 102.295 ;
        RECT 64.210 102.215 64.540 103.055 ;
        RECT 64.710 102.295 65.375 102.885 ;
        RECT 63.870 101.875 64.790 102.045 ;
        RECT 62.245 101.495 62.575 101.705 ;
        RECT 62.755 101.495 63.135 101.745 ;
        RECT 63.325 101.705 63.700 101.865 ;
        RECT 64.620 101.705 64.790 101.875 ;
        RECT 63.325 101.495 63.810 101.705 ;
        RECT 64.000 101.495 64.450 101.705 ;
        RECT 64.620 101.495 64.955 101.705 ;
        RECT 65.125 101.325 65.375 102.295 ;
        RECT 65.545 101.915 65.825 103.055 ;
        RECT 65.995 101.905 66.325 102.885 ;
        RECT 66.495 101.915 66.755 103.055 ;
        RECT 67.935 102.385 68.105 102.885 ;
        RECT 68.275 102.555 68.605 103.055 ;
        RECT 67.935 102.215 68.600 102.385 ;
        RECT 65.555 101.475 65.890 101.745 ;
        RECT 58.755 100.835 59.130 101.030 ;
        RECT 58.755 100.690 58.925 100.835 ;
        RECT 59.490 100.505 59.885 101.000 ;
        RECT 60.055 100.675 60.295 101.195 ;
        RECT 61.565 101.065 62.075 101.245 ;
        RECT 62.480 101.155 64.180 101.325 ;
        RECT 62.480 101.065 62.865 101.155 ;
        RECT 61.565 100.675 61.895 101.065 ;
        RECT 62.065 100.725 63.250 100.895 ;
        RECT 63.510 100.505 63.680 100.975 ;
        RECT 63.850 100.690 64.180 101.155 ;
        RECT 64.350 100.505 64.520 101.325 ;
        RECT 64.690 100.685 65.375 101.325 ;
        RECT 66.060 101.305 66.230 101.905 ;
        RECT 66.400 101.495 66.735 101.745 ;
        RECT 67.850 101.395 68.200 102.045 ;
        RECT 65.545 100.505 65.855 101.305 ;
        RECT 66.060 100.675 66.755 101.305 ;
        RECT 68.370 101.225 68.600 102.215 ;
        RECT 67.935 101.055 68.600 101.225 ;
        RECT 67.935 100.765 68.105 101.055 ;
        RECT 68.275 100.505 68.605 100.885 ;
        RECT 68.775 100.765 68.960 102.885 ;
        RECT 69.200 102.595 69.465 103.055 ;
        RECT 69.635 102.460 69.885 102.885 ;
        RECT 70.095 102.610 71.200 102.780 ;
        RECT 69.580 102.330 69.885 102.460 ;
        RECT 69.130 101.135 69.410 102.085 ;
        RECT 69.580 101.225 69.750 102.330 ;
        RECT 69.920 101.545 70.160 102.140 ;
        RECT 70.330 102.075 70.860 102.440 ;
        RECT 70.330 101.375 70.500 102.075 ;
        RECT 71.030 101.995 71.200 102.610 ;
        RECT 71.370 102.255 71.540 103.055 ;
        RECT 71.710 102.555 71.960 102.885 ;
        RECT 72.185 102.585 73.070 102.755 ;
        RECT 71.030 101.905 71.540 101.995 ;
        RECT 69.580 101.095 69.805 101.225 ;
        RECT 69.975 101.155 70.500 101.375 ;
        RECT 70.670 101.735 71.540 101.905 ;
        RECT 69.215 100.505 69.465 100.965 ;
        RECT 69.635 100.955 69.805 101.095 ;
        RECT 70.670 100.955 70.840 101.735 ;
        RECT 71.370 101.665 71.540 101.735 ;
        RECT 71.050 101.485 71.250 101.515 ;
        RECT 71.710 101.485 71.880 102.555 ;
        RECT 72.050 101.665 72.240 102.385 ;
        RECT 71.050 101.185 71.880 101.485 ;
        RECT 72.410 101.455 72.730 102.415 ;
        RECT 69.635 100.785 69.970 100.955 ;
        RECT 70.165 100.785 70.840 100.955 ;
        RECT 71.160 100.505 71.530 101.005 ;
        RECT 71.710 100.955 71.880 101.185 ;
        RECT 72.265 101.125 72.730 101.455 ;
        RECT 72.900 101.745 73.070 102.585 ;
        RECT 73.250 102.555 73.565 103.055 ;
        RECT 73.795 102.325 74.135 102.885 ;
        RECT 73.240 101.950 74.135 102.325 ;
        RECT 74.305 102.045 74.475 103.055 ;
        RECT 73.945 101.745 74.135 101.950 ;
        RECT 74.645 101.995 74.975 102.840 ;
        RECT 74.645 101.915 75.035 101.995 ;
        RECT 74.820 101.865 75.035 101.915 ;
        RECT 72.900 101.415 73.775 101.745 ;
        RECT 73.945 101.415 74.695 101.745 ;
        RECT 72.900 100.955 73.070 101.415 ;
        RECT 73.945 101.245 74.145 101.415 ;
        RECT 74.865 101.285 75.035 101.865 ;
        RECT 74.810 101.245 75.035 101.285 ;
        RECT 71.710 100.785 72.115 100.955 ;
        RECT 72.285 100.785 73.070 100.955 ;
        RECT 73.345 100.505 73.555 101.035 ;
        RECT 73.815 100.720 74.145 101.245 ;
        RECT 74.655 101.160 75.035 101.245 ;
        RECT 75.205 101.980 75.475 102.885 ;
        RECT 75.645 102.295 75.975 103.055 ;
        RECT 76.155 102.125 76.325 102.885 ;
        RECT 75.205 101.180 75.375 101.980 ;
        RECT 75.660 101.955 76.325 102.125 ;
        RECT 75.660 101.810 75.830 101.955 ;
        RECT 76.585 101.890 76.875 103.055 ;
        RECT 77.970 102.105 78.235 102.875 ;
        RECT 78.405 102.335 78.735 103.055 ;
        RECT 78.925 102.515 79.185 102.875 ;
        RECT 79.355 102.685 79.685 103.055 ;
        RECT 79.855 102.515 80.115 102.875 ;
        RECT 78.925 102.285 80.115 102.515 ;
        RECT 80.685 102.105 80.975 102.875 ;
        RECT 75.545 101.480 75.830 101.810 ;
        RECT 75.660 101.225 75.830 101.480 ;
        RECT 76.065 101.405 76.395 101.775 ;
        RECT 74.315 100.505 74.485 101.115 ;
        RECT 74.655 100.725 74.985 101.160 ;
        RECT 75.205 100.675 75.465 101.180 ;
        RECT 75.660 101.055 76.325 101.225 ;
        RECT 75.645 100.505 75.975 100.885 ;
        RECT 76.155 100.675 76.325 101.055 ;
        RECT 76.585 100.505 76.875 101.230 ;
        RECT 77.970 100.685 78.305 102.105 ;
        RECT 78.480 101.925 80.975 102.105 ;
        RECT 78.480 101.235 78.705 101.925 ;
        RECT 81.185 101.915 81.525 102.885 ;
        RECT 81.695 101.915 81.865 103.055 ;
        RECT 82.135 102.255 82.385 103.055 ;
        RECT 83.030 102.085 83.360 102.885 ;
        RECT 83.660 102.255 83.990 103.055 ;
        RECT 84.160 102.085 84.490 102.885 ;
        RECT 82.055 101.915 84.490 102.085 ;
        RECT 84.865 102.205 85.125 102.885 ;
        RECT 85.295 102.275 85.545 103.055 ;
        RECT 85.795 102.505 86.045 102.885 ;
        RECT 86.215 102.675 86.570 103.055 ;
        RECT 87.575 102.665 87.910 102.885 ;
        RECT 87.175 102.505 87.405 102.545 ;
        RECT 85.795 102.305 87.405 102.505 ;
        RECT 85.795 102.295 86.630 102.305 ;
        RECT 87.220 102.215 87.405 102.305 ;
        RECT 78.905 101.415 79.185 101.745 ;
        RECT 79.365 101.415 79.940 101.745 ;
        RECT 80.120 101.415 80.555 101.745 ;
        RECT 80.735 101.415 81.005 101.745 ;
        RECT 81.185 101.305 81.360 101.915 ;
        RECT 82.055 101.665 82.225 101.915 ;
        RECT 81.530 101.495 82.225 101.665 ;
        RECT 82.400 101.495 82.820 101.695 ;
        RECT 82.990 101.495 83.320 101.695 ;
        RECT 83.490 101.495 83.820 101.695 ;
        RECT 78.480 101.045 80.965 101.235 ;
        RECT 78.485 100.505 79.230 100.875 ;
        RECT 79.795 100.685 80.050 101.045 ;
        RECT 80.230 100.505 80.560 100.875 ;
        RECT 80.740 100.685 80.965 101.045 ;
        RECT 81.185 100.675 81.525 101.305 ;
        RECT 81.695 100.505 81.945 101.305 ;
        RECT 82.135 101.155 83.360 101.325 ;
        RECT 82.135 100.675 82.465 101.155 ;
        RECT 82.635 100.505 82.860 100.965 ;
        RECT 83.030 100.675 83.360 101.155 ;
        RECT 83.990 101.285 84.160 101.915 ;
        RECT 84.345 101.495 84.695 101.745 ;
        RECT 83.990 100.675 84.490 101.285 ;
        RECT 84.865 101.015 85.035 102.205 ;
        RECT 86.735 102.105 87.065 102.135 ;
        RECT 85.265 102.045 87.065 102.105 ;
        RECT 87.655 102.045 87.910 102.665 ;
        RECT 85.205 101.935 87.910 102.045 ;
        RECT 85.205 101.900 85.405 101.935 ;
        RECT 85.205 101.325 85.375 101.900 ;
        RECT 86.735 101.875 87.910 101.935 ;
        RECT 88.545 101.965 89.755 103.055 ;
        RECT 120.000 102.740 120.960 105.490 ;
        RECT 123.830 105.440 124.000 105.660 ;
        RECT 126.090 105.440 126.260 106.850 ;
        RECT 123.830 105.270 126.260 105.440 ;
        RECT 127.840 107.360 138.470 107.530 ;
        RECT 140.050 116.640 146.280 116.800 ;
        RECT 140.050 114.380 140.720 116.640 ;
        RECT 141.390 116.070 145.430 116.240 ;
        RECT 141.050 115.010 141.220 116.010 ;
        RECT 145.600 115.010 145.770 116.010 ;
        RECT 141.390 114.780 145.430 114.950 ;
        RECT 146.110 114.380 146.280 116.640 ;
        RECT 140.050 114.210 146.280 114.380 ;
        RECT 140.050 110.950 140.720 114.210 ;
        RECT 141.390 113.640 145.430 113.810 ;
        RECT 141.050 111.580 141.220 113.580 ;
        RECT 145.600 111.580 145.770 113.580 ;
        RECT 141.390 111.350 145.430 111.520 ;
        RECT 146.110 110.950 146.280 114.210 ;
        RECT 140.050 110.780 146.280 110.950 ;
        RECT 140.050 107.520 140.720 110.780 ;
        RECT 141.390 110.210 145.430 110.380 ;
        RECT 141.050 108.150 141.220 110.150 ;
        RECT 145.600 108.150 145.770 110.150 ;
        RECT 141.390 107.920 145.430 108.090 ;
        RECT 146.110 107.520 146.280 110.780 ;
        RECT 140.050 107.510 146.280 107.520 ;
        RECT 147.870 116.780 157.700 116.820 ;
        RECT 147.870 116.650 158.500 116.780 ;
        RECT 147.870 114.390 148.040 116.650 ;
        RECT 148.765 116.080 156.805 116.250 ;
        RECT 148.380 115.020 148.550 116.020 ;
        RECT 157.020 115.020 157.190 116.020 ;
        RECT 148.765 114.790 156.805 114.960 ;
        RECT 157.530 114.390 158.500 116.650 ;
        RECT 147.870 114.220 158.500 114.390 ;
        RECT 147.870 110.960 148.040 114.220 ;
        RECT 148.765 113.650 156.805 113.820 ;
        RECT 148.380 111.590 148.550 113.590 ;
        RECT 157.020 111.590 157.190 113.590 ;
        RECT 148.765 111.360 156.805 111.530 ;
        RECT 157.530 110.960 158.500 114.220 ;
        RECT 147.870 110.790 158.500 110.960 ;
        RECT 147.870 107.530 148.040 110.790 ;
        RECT 148.765 110.220 156.805 110.390 ;
        RECT 148.380 108.160 148.550 110.160 ;
        RECT 157.020 108.160 157.190 110.160 ;
        RECT 148.765 107.930 156.805 108.100 ;
        RECT 157.530 107.530 158.500 110.790 ;
        RECT 140.050 107.410 146.290 107.510 ;
        RECT 127.840 105.100 128.010 107.360 ;
        RECT 128.735 106.790 136.775 106.960 ;
        RECT 128.350 105.730 128.520 106.730 ;
        RECT 136.990 105.730 137.160 106.730 ;
        RECT 128.735 105.500 136.775 105.670 ;
        RECT 137.500 105.100 138.470 107.360 ;
        RECT 140.040 106.850 146.290 107.410 ;
        RECT 140.040 106.830 145.210 106.850 ;
        RECT 140.040 106.760 144.030 106.830 ;
        RECT 140.040 105.490 141.960 106.760 ;
        RECT 143.470 106.750 144.030 106.760 ;
        RECT 143.700 105.660 144.030 106.750 ;
        RECT 144.400 106.280 145.440 106.450 ;
        RECT 144.400 105.840 145.440 106.010 ;
        RECT 145.610 105.980 145.780 106.310 ;
        RECT 143.860 105.440 144.030 105.660 ;
        RECT 146.120 105.440 146.290 106.850 ;
        RECT 143.860 105.270 146.290 105.440 ;
        RECT 147.870 107.360 158.500 107.530 ;
        RECT 127.840 105.070 138.470 105.100 ;
        RECT 147.870 105.100 148.040 107.360 ;
        RECT 148.765 106.790 156.805 106.960 ;
        RECT 148.380 105.730 148.550 106.730 ;
        RECT 157.020 105.730 157.190 106.730 ;
        RECT 148.765 105.500 156.805 105.670 ;
        RECT 157.530 105.100 158.500 107.360 ;
        RECT 147.870 105.070 158.500 105.100 ;
        RECT 127.810 104.960 138.470 105.070 ;
        RECT 147.840 104.960 158.500 105.070 ;
        RECT 126.060 104.910 138.470 104.960 ;
        RECT 146.090 104.910 158.500 104.960 ;
        RECT 121.720 104.740 138.470 104.910 ;
        RECT 121.720 103.330 121.890 104.740 ;
        RECT 122.260 104.170 125.300 104.340 ;
        RECT 122.260 103.730 125.300 103.900 ;
        RECT 125.515 103.870 125.685 104.200 ;
        RECT 126.020 103.980 138.470 104.740 ;
        RECT 141.750 104.740 158.500 104.910 ;
        RECT 126.020 103.970 138.360 103.980 ;
        RECT 126.020 103.960 131.900 103.970 ;
        RECT 126.020 103.940 126.590 103.960 ;
        RECT 127.810 103.950 131.900 103.960 ;
        RECT 126.030 103.330 126.200 103.940 ;
        RECT 121.720 103.160 126.200 103.330 ;
        RECT 141.750 103.330 141.920 104.740 ;
        RECT 142.290 104.170 145.330 104.340 ;
        RECT 142.290 103.730 145.330 103.900 ;
        RECT 145.545 103.870 145.715 104.200 ;
        RECT 146.050 103.980 158.500 104.740 ;
        RECT 146.050 103.970 158.390 103.980 ;
        RECT 146.050 103.960 151.930 103.970 ;
        RECT 146.050 103.940 146.620 103.960 ;
        RECT 147.840 103.950 151.930 103.960 ;
        RECT 146.060 103.330 146.230 103.940 ;
        RECT 141.750 103.160 146.230 103.330 ;
        RECT 120.000 102.570 158.300 102.740 ;
        RECT 85.605 101.460 86.015 101.765 ;
        RECT 86.185 101.495 86.515 101.705 ;
        RECT 85.205 101.205 85.475 101.325 ;
        RECT 85.205 101.160 86.050 101.205 ;
        RECT 85.295 101.035 86.050 101.160 ;
        RECT 86.305 101.095 86.515 101.495 ;
        RECT 86.760 101.495 87.235 101.705 ;
        RECT 87.425 101.495 87.915 101.695 ;
        RECT 86.760 101.095 86.980 101.495 ;
        RECT 88.545 101.425 89.065 101.965 ;
        RECT 84.865 101.005 85.095 101.015 ;
        RECT 84.865 100.675 85.125 101.005 ;
        RECT 85.880 100.885 86.050 101.035 ;
        RECT 85.295 100.505 85.625 100.865 ;
        RECT 85.880 100.675 87.180 100.885 ;
        RECT 87.455 100.505 87.910 101.270 ;
        RECT 89.235 101.255 89.755 101.795 ;
        RECT 120.000 101.720 134.620 102.570 ;
        RECT 120.000 101.650 120.960 101.720 ;
        RECT 88.545 100.505 89.755 101.255 ;
        RECT 12.100 100.335 89.840 100.505 ;
        RECT 100.030 100.395 112.740 101.005 ;
        RECT 12.185 99.585 13.395 100.335 ;
        RECT 12.185 99.045 12.705 99.585 ;
        RECT 13.565 99.565 17.075 100.335 ;
        RECT 12.875 98.875 13.395 99.415 ;
        RECT 13.565 99.045 15.215 99.565 ;
        RECT 18.185 99.525 18.425 100.335 ;
        RECT 18.595 99.525 18.925 100.165 ;
        RECT 19.095 99.525 19.365 100.335 ;
        RECT 19.545 99.790 24.890 100.335 ;
        RECT 26.050 99.945 28.060 100.115 ;
        RECT 15.385 98.875 17.075 99.395 ;
        RECT 18.165 99.095 18.515 99.345 ;
        RECT 18.685 98.925 18.855 99.525 ;
        RECT 19.025 99.095 19.375 99.345 ;
        RECT 21.130 98.960 21.470 99.790 ;
        RECT 25.985 99.515 27.640 99.775 ;
        RECT 27.810 99.685 28.060 99.945 ;
        RECT 28.250 99.865 28.520 100.335 ;
        RECT 28.690 99.695 29.020 100.165 ;
        RECT 29.190 99.865 29.360 100.335 ;
        RECT 29.530 99.695 29.860 100.165 ;
        RECT 30.030 99.865 30.200 100.335 ;
        RECT 30.370 99.695 30.700 100.165 ;
        RECT 30.870 99.865 31.040 100.335 ;
        RECT 31.210 99.695 31.540 100.165 ;
        RECT 28.590 99.685 31.540 99.695 ;
        RECT 27.810 99.515 31.540 99.685 ;
        RECT 31.710 99.515 31.985 100.335 ;
        RECT 32.160 99.695 32.490 100.165 ;
        RECT 32.660 99.865 32.830 100.335 ;
        RECT 33.000 99.695 33.330 100.165 ;
        RECT 33.500 99.865 33.670 100.335 ;
        RECT 33.840 99.945 35.850 100.165 ;
        RECT 33.840 99.695 34.090 99.945 ;
        RECT 32.160 99.515 34.090 99.695 ;
        RECT 34.260 99.515 35.935 99.775 ;
        RECT 25.985 99.485 26.215 99.515 ;
        RECT 12.185 97.785 13.395 98.875 ;
        RECT 13.565 97.785 17.075 98.875 ;
        RECT 18.175 98.755 18.855 98.925 ;
        RECT 18.175 97.970 18.505 98.755 ;
        RECT 19.035 97.785 19.365 98.925 ;
        RECT 22.950 98.220 23.300 99.470 ;
        RECT 25.985 98.975 26.205 99.485 ;
        RECT 26.375 99.145 28.420 99.345 ;
        RECT 28.590 99.145 30.460 99.345 ;
        RECT 30.630 99.145 33.845 99.345 ;
        RECT 34.165 99.145 35.530 99.345 ;
        RECT 28.250 98.975 28.420 99.145 ;
        RECT 30.290 98.975 30.460 99.145 ;
        RECT 34.165 98.975 34.335 99.145 ;
        RECT 35.700 98.975 35.935 99.515 ;
        RECT 36.105 99.565 37.775 100.335 ;
        RECT 37.945 99.610 38.235 100.335 ;
        RECT 36.105 99.045 36.855 99.565 ;
        RECT 38.405 99.535 38.715 100.335 ;
        RECT 38.920 99.535 39.615 100.165 ;
        RECT 25.985 98.755 28.060 98.975 ;
        RECT 28.250 98.805 30.120 98.975 ;
        RECT 30.290 98.805 34.335 98.975 ;
        RECT 34.720 98.805 35.935 98.975 ;
        RECT 37.025 98.875 37.775 99.395 ;
        RECT 38.415 99.095 38.750 99.365 ;
        RECT 19.545 97.785 24.890 98.220 ;
        RECT 25.985 97.955 26.340 98.755 ;
        RECT 26.510 97.785 26.760 98.585 ;
        RECT 26.930 97.955 27.180 98.755 ;
        RECT 27.770 98.635 28.060 98.755 ;
        RECT 34.720 98.635 34.970 98.805 ;
        RECT 27.350 97.785 27.600 98.585 ;
        RECT 27.770 98.375 29.860 98.635 ;
        RECT 30.030 98.415 31.985 98.635 ;
        RECT 27.770 97.955 28.060 98.375 ;
        RECT 30.030 98.205 30.240 98.415 ;
        RECT 28.270 97.955 30.240 98.205 ;
        RECT 30.410 97.785 30.660 98.245 ;
        RECT 30.830 97.955 31.080 98.415 ;
        RECT 31.250 97.785 31.500 98.245 ;
        RECT 31.670 97.955 31.985 98.415 ;
        RECT 32.200 98.415 34.970 98.635 ;
        RECT 32.200 97.955 32.450 98.415 ;
        RECT 32.620 97.785 32.870 98.245 ;
        RECT 33.040 97.955 33.290 98.415 ;
        RECT 33.460 97.785 33.710 98.245 ;
        RECT 33.880 97.955 34.130 98.415 ;
        RECT 34.300 97.785 34.550 98.245 ;
        RECT 34.720 97.955 34.970 98.415 ;
        RECT 35.140 97.785 35.390 98.585 ;
        RECT 35.560 97.955 35.935 98.805 ;
        RECT 36.105 97.785 37.775 98.875 ;
        RECT 37.945 97.785 38.235 98.950 ;
        RECT 38.920 98.935 39.090 99.535 ;
        RECT 39.845 99.515 40.055 100.335 ;
        RECT 40.225 99.535 40.555 100.165 ;
        RECT 39.260 99.095 39.595 99.345 ;
        RECT 40.225 98.935 40.475 99.535 ;
        RECT 40.725 99.515 40.955 100.335 ;
        RECT 42.175 99.785 42.345 100.075 ;
        RECT 42.515 99.955 42.845 100.335 ;
        RECT 42.175 99.615 42.840 99.785 ;
        RECT 40.645 99.095 40.975 99.345 ;
        RECT 38.405 97.785 38.685 98.925 ;
        RECT 38.855 97.955 39.185 98.935 ;
        RECT 39.355 97.785 39.615 98.925 ;
        RECT 39.845 97.785 40.055 98.925 ;
        RECT 40.225 97.955 40.555 98.935 ;
        RECT 40.725 97.785 40.955 98.925 ;
        RECT 42.090 98.795 42.440 99.445 ;
        RECT 42.610 98.625 42.840 99.615 ;
        RECT 42.175 98.455 42.840 98.625 ;
        RECT 42.175 97.955 42.345 98.455 ;
        RECT 42.515 97.785 42.845 98.285 ;
        RECT 43.015 97.955 43.200 100.075 ;
        RECT 43.455 99.875 43.705 100.335 ;
        RECT 43.875 99.885 44.210 100.055 ;
        RECT 44.405 99.885 45.080 100.055 ;
        RECT 43.875 99.745 44.045 99.885 ;
        RECT 43.370 98.755 43.650 99.705 ;
        RECT 43.820 99.615 44.045 99.745 ;
        RECT 43.820 98.510 43.990 99.615 ;
        RECT 44.215 99.465 44.740 99.685 ;
        RECT 44.160 98.700 44.400 99.295 ;
        RECT 44.570 98.765 44.740 99.465 ;
        RECT 44.910 99.105 45.080 99.885 ;
        RECT 45.400 99.835 45.770 100.335 ;
        RECT 45.950 99.885 46.355 100.055 ;
        RECT 46.525 99.885 47.310 100.055 ;
        RECT 45.950 99.655 46.120 99.885 ;
        RECT 45.290 99.355 46.120 99.655 ;
        RECT 46.505 99.385 46.970 99.715 ;
        RECT 45.290 99.325 45.490 99.355 ;
        RECT 45.610 99.105 45.780 99.175 ;
        RECT 44.910 98.935 45.780 99.105 ;
        RECT 45.270 98.845 45.780 98.935 ;
        RECT 43.820 98.380 44.125 98.510 ;
        RECT 44.570 98.400 45.100 98.765 ;
        RECT 43.440 97.785 43.705 98.245 ;
        RECT 43.875 97.955 44.125 98.380 ;
        RECT 45.270 98.230 45.440 98.845 ;
        RECT 44.335 98.060 45.440 98.230 ;
        RECT 45.610 97.785 45.780 98.585 ;
        RECT 45.950 98.285 46.120 99.355 ;
        RECT 46.290 98.455 46.480 99.175 ;
        RECT 46.650 98.425 46.970 99.385 ;
        RECT 47.140 99.425 47.310 99.885 ;
        RECT 47.585 99.805 47.795 100.335 ;
        RECT 48.055 99.595 48.385 100.120 ;
        RECT 48.555 99.725 48.725 100.335 ;
        RECT 48.895 99.680 49.225 100.115 ;
        RECT 49.450 99.830 49.785 100.335 ;
        RECT 49.955 99.765 50.195 100.140 ;
        RECT 50.475 100.005 50.645 100.150 ;
        RECT 50.475 99.810 50.850 100.005 ;
        RECT 51.210 99.840 51.605 100.335 ;
        RECT 48.895 99.595 49.275 99.680 ;
        RECT 48.185 99.425 48.385 99.595 ;
        RECT 49.050 99.555 49.275 99.595 ;
        RECT 47.140 99.095 48.015 99.425 ;
        RECT 48.185 99.095 48.935 99.425 ;
        RECT 45.950 97.955 46.200 98.285 ;
        RECT 47.140 98.255 47.310 99.095 ;
        RECT 48.185 98.890 48.375 99.095 ;
        RECT 49.105 98.975 49.275 99.555 ;
        RECT 49.060 98.925 49.275 98.975 ;
        RECT 47.480 98.515 48.375 98.890 ;
        RECT 48.885 98.845 49.275 98.925 ;
        RECT 46.425 98.085 47.310 98.255 ;
        RECT 47.490 97.785 47.805 98.285 ;
        RECT 48.035 97.955 48.375 98.515 ;
        RECT 48.545 97.785 48.715 98.795 ;
        RECT 48.885 98.000 49.215 98.845 ;
        RECT 49.505 98.805 49.805 99.655 ;
        RECT 49.975 99.615 50.195 99.765 ;
        RECT 49.975 99.285 50.510 99.615 ;
        RECT 50.680 99.475 50.850 99.810 ;
        RECT 51.775 99.645 52.015 100.165 ;
        RECT 49.975 98.635 50.210 99.285 ;
        RECT 50.680 99.115 51.665 99.475 ;
        RECT 49.535 98.405 50.210 98.635 ;
        RECT 50.380 99.095 51.665 99.115 ;
        RECT 50.380 98.945 51.240 99.095 ;
        RECT 49.535 97.975 49.705 98.405 ;
        RECT 49.875 97.785 50.205 98.235 ;
        RECT 50.380 98.000 50.665 98.945 ;
        RECT 51.840 98.840 52.015 99.645 ;
        RECT 53.125 99.705 53.465 100.165 ;
        RECT 53.635 99.875 53.805 100.335 ;
        RECT 53.975 99.955 55.145 100.165 ;
        RECT 55.425 99.955 56.315 100.125 ;
        RECT 53.975 99.705 54.225 99.955 ;
        RECT 54.815 99.935 55.145 99.955 ;
        RECT 53.125 99.535 54.225 99.705 ;
        RECT 54.395 99.515 55.255 99.765 ;
        RECT 53.125 99.095 53.885 99.345 ;
        RECT 54.055 99.095 54.805 99.345 ;
        RECT 54.975 98.925 55.255 99.515 ;
        RECT 55.425 99.400 55.975 99.785 ;
        RECT 56.145 99.230 56.315 99.955 ;
        RECT 50.840 98.465 51.535 98.775 ;
        RECT 50.845 97.785 51.530 98.255 ;
        RECT 51.710 98.055 52.015 98.840 ;
        RECT 53.125 97.785 53.385 98.925 ;
        RECT 53.555 98.755 55.255 98.925 ;
        RECT 55.425 99.160 56.315 99.230 ;
        RECT 56.485 99.655 56.705 100.115 ;
        RECT 56.875 99.795 57.125 100.335 ;
        RECT 57.295 99.685 57.555 100.165 ;
        RECT 57.745 99.825 57.985 100.335 ;
        RECT 58.155 99.825 58.445 100.165 ;
        RECT 58.675 99.825 58.990 100.335 ;
        RECT 56.485 99.630 56.735 99.655 ;
        RECT 56.485 99.205 56.815 99.630 ;
        RECT 55.425 99.135 56.320 99.160 ;
        RECT 55.425 99.120 56.330 99.135 ;
        RECT 55.425 99.105 56.335 99.120 ;
        RECT 55.425 99.100 56.345 99.105 ;
        RECT 55.425 99.090 56.350 99.100 ;
        RECT 55.425 99.080 56.355 99.090 ;
        RECT 55.425 99.075 56.365 99.080 ;
        RECT 55.425 99.065 56.375 99.075 ;
        RECT 55.425 99.060 56.385 99.065 ;
        RECT 53.555 97.955 53.885 98.755 ;
        RECT 54.055 97.785 54.225 98.585 ;
        RECT 54.395 97.955 54.725 98.755 ;
        RECT 55.425 98.610 55.685 99.060 ;
        RECT 56.050 99.055 56.385 99.060 ;
        RECT 56.050 99.050 56.400 99.055 ;
        RECT 56.050 99.040 56.415 99.050 ;
        RECT 56.050 99.035 56.440 99.040 ;
        RECT 56.985 99.035 57.215 99.430 ;
        RECT 56.050 99.030 57.215 99.035 ;
        RECT 56.080 98.995 57.215 99.030 ;
        RECT 56.115 98.970 57.215 98.995 ;
        RECT 56.145 98.940 57.215 98.970 ;
        RECT 56.165 98.910 57.215 98.940 ;
        RECT 56.185 98.880 57.215 98.910 ;
        RECT 56.255 98.870 57.215 98.880 ;
        RECT 56.280 98.860 57.215 98.870 ;
        RECT 56.300 98.845 57.215 98.860 ;
        RECT 56.320 98.830 57.215 98.845 ;
        RECT 56.325 98.820 57.110 98.830 ;
        RECT 56.340 98.785 57.110 98.820 ;
        RECT 54.895 97.785 55.150 98.585 ;
        RECT 55.855 98.465 56.185 98.710 ;
        RECT 56.355 98.535 57.110 98.785 ;
        RECT 57.385 98.655 57.555 99.685 ;
        RECT 57.790 99.315 57.985 99.655 ;
        RECT 57.785 99.145 57.985 99.315 ;
        RECT 57.790 99.095 57.985 99.145 ;
        RECT 58.155 98.925 58.335 99.825 ;
        RECT 59.160 99.765 59.330 100.035 ;
        RECT 59.500 99.935 59.830 100.335 ;
        RECT 58.505 99.095 58.915 99.655 ;
        RECT 59.160 99.595 59.855 99.765 ;
        RECT 60.965 99.605 61.255 100.335 ;
        RECT 59.085 98.925 59.255 99.425 ;
        RECT 55.855 98.440 56.040 98.465 ;
        RECT 55.425 98.340 56.040 98.440 ;
        RECT 55.425 97.785 56.030 98.340 ;
        RECT 56.205 97.955 56.685 98.295 ;
        RECT 56.855 97.785 57.110 98.330 ;
        RECT 57.280 97.955 57.555 98.655 ;
        RECT 57.795 98.755 59.255 98.925 ;
        RECT 57.795 98.580 58.155 98.755 ;
        RECT 59.425 98.585 59.855 99.595 ;
        RECT 60.955 99.095 61.255 99.425 ;
        RECT 61.435 99.405 61.665 100.045 ;
        RECT 61.845 99.785 62.155 100.155 ;
        RECT 62.335 99.965 63.005 100.335 ;
        RECT 61.845 99.585 63.075 99.785 ;
        RECT 61.435 99.095 61.960 99.405 ;
        RECT 62.140 99.095 62.605 99.405 ;
        RECT 62.785 98.915 63.075 99.585 ;
        RECT 58.740 97.785 58.910 98.585 ;
        RECT 59.080 98.415 59.855 98.585 ;
        RECT 60.965 98.675 62.125 98.915 ;
        RECT 59.080 97.955 59.410 98.415 ;
        RECT 59.580 97.785 59.750 98.245 ;
        RECT 60.965 97.965 61.225 98.675 ;
        RECT 61.395 97.785 61.725 98.495 ;
        RECT 61.895 97.965 62.125 98.675 ;
        RECT 62.305 98.695 63.075 98.915 ;
        RECT 62.305 97.965 62.575 98.695 ;
        RECT 62.755 97.785 63.095 98.515 ;
        RECT 63.265 97.965 63.525 100.155 ;
        RECT 63.705 99.610 63.995 100.335 ;
        RECT 64.165 99.565 65.835 100.335 ;
        RECT 66.095 99.785 66.265 100.075 ;
        RECT 66.435 99.955 66.765 100.335 ;
        RECT 66.095 99.615 66.760 99.785 ;
        RECT 64.165 99.045 64.915 99.565 ;
        RECT 63.705 97.785 63.995 98.950 ;
        RECT 65.085 98.875 65.835 99.395 ;
        RECT 64.165 97.785 65.835 98.875 ;
        RECT 66.010 98.795 66.360 99.445 ;
        RECT 66.530 98.625 66.760 99.615 ;
        RECT 66.095 98.455 66.760 98.625 ;
        RECT 66.095 97.955 66.265 98.455 ;
        RECT 66.435 97.785 66.765 98.285 ;
        RECT 66.935 97.955 67.120 100.075 ;
        RECT 67.375 99.875 67.625 100.335 ;
        RECT 67.795 99.885 68.130 100.055 ;
        RECT 68.325 99.885 69.000 100.055 ;
        RECT 67.795 99.745 67.965 99.885 ;
        RECT 67.290 98.755 67.570 99.705 ;
        RECT 67.740 99.615 67.965 99.745 ;
        RECT 67.740 98.510 67.910 99.615 ;
        RECT 68.135 99.465 68.660 99.685 ;
        RECT 68.080 98.700 68.320 99.295 ;
        RECT 68.490 98.765 68.660 99.465 ;
        RECT 68.830 99.105 69.000 99.885 ;
        RECT 69.320 99.835 69.690 100.335 ;
        RECT 69.870 99.885 70.275 100.055 ;
        RECT 70.445 99.885 71.230 100.055 ;
        RECT 69.870 99.655 70.040 99.885 ;
        RECT 69.210 99.355 70.040 99.655 ;
        RECT 70.425 99.385 70.890 99.715 ;
        RECT 69.210 99.325 69.410 99.355 ;
        RECT 69.530 99.105 69.700 99.175 ;
        RECT 68.830 98.935 69.700 99.105 ;
        RECT 69.190 98.845 69.700 98.935 ;
        RECT 67.740 98.380 68.045 98.510 ;
        RECT 68.490 98.400 69.020 98.765 ;
        RECT 67.360 97.785 67.625 98.245 ;
        RECT 67.795 97.955 68.045 98.380 ;
        RECT 69.190 98.230 69.360 98.845 ;
        RECT 68.255 98.060 69.360 98.230 ;
        RECT 69.530 97.785 69.700 98.585 ;
        RECT 69.870 98.285 70.040 99.355 ;
        RECT 70.210 98.455 70.400 99.175 ;
        RECT 70.570 98.425 70.890 99.385 ;
        RECT 71.060 99.425 71.230 99.885 ;
        RECT 71.505 99.805 71.715 100.335 ;
        RECT 71.975 99.595 72.305 100.120 ;
        RECT 72.475 99.725 72.645 100.335 ;
        RECT 72.815 99.680 73.145 100.115 ;
        RECT 72.815 99.595 73.195 99.680 ;
        RECT 72.105 99.425 72.305 99.595 ;
        RECT 72.970 99.555 73.195 99.595 ;
        RECT 71.060 99.095 71.935 99.425 ;
        RECT 72.105 99.095 72.855 99.425 ;
        RECT 69.870 97.955 70.120 98.285 ;
        RECT 71.060 98.255 71.230 99.095 ;
        RECT 72.105 98.890 72.295 99.095 ;
        RECT 73.025 98.975 73.195 99.555 ;
        RECT 72.980 98.925 73.195 98.975 ;
        RECT 71.400 98.515 72.295 98.890 ;
        RECT 72.805 98.845 73.195 98.925 ;
        RECT 73.365 99.595 73.750 100.165 ;
        RECT 73.920 99.875 74.245 100.335 ;
        RECT 74.765 99.705 75.045 100.165 ;
        RECT 73.365 98.925 73.645 99.595 ;
        RECT 73.920 99.535 75.045 99.705 ;
        RECT 73.920 99.425 74.370 99.535 ;
        RECT 73.815 99.095 74.370 99.425 ;
        RECT 75.235 99.365 75.635 100.165 ;
        RECT 76.035 99.875 76.305 100.335 ;
        RECT 76.475 99.705 76.760 100.165 ;
        RECT 70.345 98.085 71.230 98.255 ;
        RECT 71.410 97.785 71.725 98.285 ;
        RECT 71.955 97.955 72.295 98.515 ;
        RECT 72.465 97.785 72.635 98.795 ;
        RECT 72.805 98.000 73.135 98.845 ;
        RECT 73.365 97.955 73.750 98.925 ;
        RECT 73.920 98.635 74.370 99.095 ;
        RECT 74.540 98.805 75.635 99.365 ;
        RECT 73.920 98.415 75.045 98.635 ;
        RECT 73.920 97.785 74.245 98.245 ;
        RECT 74.765 97.955 75.045 98.415 ;
        RECT 75.235 97.955 75.635 98.805 ;
        RECT 75.805 99.535 76.760 99.705 ;
        RECT 75.805 98.635 76.015 99.535 ;
        RECT 77.050 99.495 77.310 100.335 ;
        RECT 77.485 99.590 77.740 100.165 ;
        RECT 77.910 99.955 78.240 100.335 ;
        RECT 78.455 99.785 78.625 100.165 ;
        RECT 77.910 99.615 78.625 99.785 ;
        RECT 78.975 99.785 79.145 100.075 ;
        RECT 79.315 99.955 79.645 100.335 ;
        RECT 78.975 99.615 79.640 99.785 ;
        RECT 76.185 98.805 76.875 99.365 ;
        RECT 75.805 98.415 76.760 98.635 ;
        RECT 76.035 97.785 76.305 98.245 ;
        RECT 76.475 97.955 76.760 98.415 ;
        RECT 77.050 97.785 77.310 98.935 ;
        RECT 77.485 98.860 77.655 99.590 ;
        RECT 77.910 99.425 78.080 99.615 ;
        RECT 77.825 99.095 78.080 99.425 ;
        RECT 77.910 98.885 78.080 99.095 ;
        RECT 78.360 99.065 78.715 99.435 ;
        RECT 77.485 97.955 77.740 98.860 ;
        RECT 77.910 98.715 78.625 98.885 ;
        RECT 78.890 98.795 79.240 99.445 ;
        RECT 77.910 97.785 78.240 98.545 ;
        RECT 78.455 97.955 78.625 98.715 ;
        RECT 79.410 98.625 79.640 99.615 ;
        RECT 78.975 98.455 79.640 98.625 ;
        RECT 78.975 97.955 79.145 98.455 ;
        RECT 79.315 97.785 79.645 98.285 ;
        RECT 79.815 97.955 80.000 100.075 ;
        RECT 80.255 99.875 80.505 100.335 ;
        RECT 80.675 99.885 81.010 100.055 ;
        RECT 81.205 99.885 81.880 100.055 ;
        RECT 80.675 99.745 80.845 99.885 ;
        RECT 80.170 98.755 80.450 99.705 ;
        RECT 80.620 99.615 80.845 99.745 ;
        RECT 80.620 98.510 80.790 99.615 ;
        RECT 81.015 99.465 81.540 99.685 ;
        RECT 80.960 98.700 81.200 99.295 ;
        RECT 81.370 98.765 81.540 99.465 ;
        RECT 81.710 99.105 81.880 99.885 ;
        RECT 82.200 99.835 82.570 100.335 ;
        RECT 82.750 99.885 83.155 100.055 ;
        RECT 83.325 99.885 84.110 100.055 ;
        RECT 82.750 99.655 82.920 99.885 ;
        RECT 82.090 99.355 82.920 99.655 ;
        RECT 83.305 99.385 83.770 99.715 ;
        RECT 82.090 99.325 82.290 99.355 ;
        RECT 82.410 99.105 82.580 99.175 ;
        RECT 81.710 98.935 82.580 99.105 ;
        RECT 82.070 98.845 82.580 98.935 ;
        RECT 80.620 98.380 80.925 98.510 ;
        RECT 81.370 98.400 81.900 98.765 ;
        RECT 80.240 97.785 80.505 98.245 ;
        RECT 80.675 97.955 80.925 98.380 ;
        RECT 82.070 98.230 82.240 98.845 ;
        RECT 81.135 98.060 82.240 98.230 ;
        RECT 82.410 97.785 82.580 98.585 ;
        RECT 82.750 98.285 82.920 99.355 ;
        RECT 83.090 98.455 83.280 99.175 ;
        RECT 83.450 98.425 83.770 99.385 ;
        RECT 83.940 99.425 84.110 99.885 ;
        RECT 84.385 99.805 84.595 100.335 ;
        RECT 84.855 99.595 85.185 100.120 ;
        RECT 85.355 99.725 85.525 100.335 ;
        RECT 85.695 99.680 86.025 100.115 ;
        RECT 86.410 99.825 86.650 100.335 ;
        RECT 86.830 99.825 87.110 100.155 ;
        RECT 87.340 99.825 87.555 100.335 ;
        RECT 85.695 99.595 86.075 99.680 ;
        RECT 84.985 99.425 85.185 99.595 ;
        RECT 85.850 99.555 86.075 99.595 ;
        RECT 83.940 99.095 84.815 99.425 ;
        RECT 84.985 99.095 85.735 99.425 ;
        RECT 82.750 97.955 83.000 98.285 ;
        RECT 83.940 98.255 84.110 99.095 ;
        RECT 84.985 98.890 85.175 99.095 ;
        RECT 85.905 98.975 86.075 99.555 ;
        RECT 86.305 99.095 86.660 99.655 ;
        RECT 85.860 98.925 86.075 98.975 ;
        RECT 86.830 98.925 87.000 99.825 ;
        RECT 87.170 99.095 87.435 99.655 ;
        RECT 87.725 99.595 88.340 100.165 ;
        RECT 87.685 98.925 87.855 99.425 ;
        RECT 84.280 98.515 85.175 98.890 ;
        RECT 85.685 98.845 86.075 98.925 ;
        RECT 83.225 98.085 84.110 98.255 ;
        RECT 84.290 97.785 84.605 98.285 ;
        RECT 84.835 97.955 85.175 98.515 ;
        RECT 85.345 97.785 85.515 98.795 ;
        RECT 85.685 98.000 86.015 98.845 ;
        RECT 86.430 98.755 87.855 98.925 ;
        RECT 86.430 98.580 86.820 98.755 ;
        RECT 87.305 97.785 87.635 98.585 ;
        RECT 88.025 98.575 88.340 99.595 ;
        RECT 88.545 99.585 89.755 100.335 ;
        RECT 87.805 97.955 88.340 98.575 ;
        RECT 88.545 98.875 89.065 99.415 ;
        RECT 89.235 99.045 89.755 99.585 ;
        RECT 99.980 100.195 112.790 100.395 ;
        RECT 88.545 97.785 89.755 98.875 ;
        RECT 12.100 97.615 89.840 97.785 ;
        RECT 12.185 96.525 13.395 97.615 ;
        RECT 12.185 95.815 12.705 96.355 ;
        RECT 12.875 95.985 13.395 96.525 ;
        RECT 13.565 96.745 13.840 97.445 ;
        RECT 14.010 97.070 14.265 97.615 ;
        RECT 14.435 97.105 14.915 97.445 ;
        RECT 15.090 97.060 15.695 97.615 ;
        RECT 15.080 96.960 15.695 97.060 ;
        RECT 15.080 96.935 15.265 96.960 ;
        RECT 12.185 95.065 13.395 95.815 ;
        RECT 13.565 95.715 13.735 96.745 ;
        RECT 14.010 96.615 14.765 96.865 ;
        RECT 14.935 96.690 15.265 96.935 ;
        RECT 14.010 96.580 14.780 96.615 ;
        RECT 14.010 96.570 14.795 96.580 ;
        RECT 13.905 96.555 14.800 96.570 ;
        RECT 13.905 96.540 14.820 96.555 ;
        RECT 13.905 96.530 14.840 96.540 ;
        RECT 13.905 96.520 14.865 96.530 ;
        RECT 13.905 96.490 14.935 96.520 ;
        RECT 13.905 96.460 14.955 96.490 ;
        RECT 13.905 96.430 14.975 96.460 ;
        RECT 13.905 96.405 15.005 96.430 ;
        RECT 13.905 96.370 15.040 96.405 ;
        RECT 13.905 96.365 15.070 96.370 ;
        RECT 13.905 95.970 14.135 96.365 ;
        RECT 14.680 96.360 15.070 96.365 ;
        RECT 14.705 96.350 15.070 96.360 ;
        RECT 14.720 96.345 15.070 96.350 ;
        RECT 14.735 96.340 15.070 96.345 ;
        RECT 15.435 96.340 15.695 96.790 ;
        RECT 14.735 96.335 15.695 96.340 ;
        RECT 14.745 96.325 15.695 96.335 ;
        RECT 14.755 96.320 15.695 96.325 ;
        RECT 14.765 96.310 15.695 96.320 ;
        RECT 14.770 96.300 15.695 96.310 ;
        RECT 14.775 96.295 15.695 96.300 ;
        RECT 14.785 96.280 15.695 96.295 ;
        RECT 14.790 96.265 15.695 96.280 ;
        RECT 14.800 96.240 15.695 96.265 ;
        RECT 14.305 95.770 14.635 96.195 ;
        RECT 13.565 95.235 13.825 95.715 ;
        RECT 13.995 95.065 14.245 95.605 ;
        RECT 14.415 95.285 14.635 95.770 ;
        RECT 14.805 96.170 15.695 96.240 ;
        RECT 15.865 96.745 16.140 97.445 ;
        RECT 16.310 97.070 16.565 97.615 ;
        RECT 16.735 97.105 17.215 97.445 ;
        RECT 17.390 97.060 17.995 97.615 ;
        RECT 17.380 96.960 17.995 97.060 ;
        RECT 17.380 96.935 17.565 96.960 ;
        RECT 14.805 95.445 14.975 96.170 ;
        RECT 15.145 95.615 15.695 96.000 ;
        RECT 15.865 95.715 16.035 96.745 ;
        RECT 16.310 96.615 17.065 96.865 ;
        RECT 17.235 96.690 17.565 96.935 ;
        RECT 16.310 96.580 17.080 96.615 ;
        RECT 16.310 96.570 17.095 96.580 ;
        RECT 16.205 96.555 17.100 96.570 ;
        RECT 16.205 96.540 17.120 96.555 ;
        RECT 16.205 96.530 17.140 96.540 ;
        RECT 16.205 96.520 17.165 96.530 ;
        RECT 16.205 96.490 17.235 96.520 ;
        RECT 16.205 96.460 17.255 96.490 ;
        RECT 16.205 96.430 17.275 96.460 ;
        RECT 16.205 96.405 17.305 96.430 ;
        RECT 16.205 96.370 17.340 96.405 ;
        RECT 16.205 96.365 17.370 96.370 ;
        RECT 16.205 95.970 16.435 96.365 ;
        RECT 16.980 96.360 17.370 96.365 ;
        RECT 17.005 96.350 17.370 96.360 ;
        RECT 17.020 96.345 17.370 96.350 ;
        RECT 17.035 96.340 17.370 96.345 ;
        RECT 17.735 96.340 17.995 96.790 ;
        RECT 18.635 96.475 18.965 97.615 ;
        RECT 19.495 96.645 19.825 97.430 ;
        RECT 20.005 96.795 20.350 97.615 ;
        RECT 19.145 96.475 19.825 96.645 ;
        RECT 17.035 96.335 17.995 96.340 ;
        RECT 17.045 96.325 17.995 96.335 ;
        RECT 17.055 96.320 17.995 96.325 ;
        RECT 17.065 96.310 17.995 96.320 ;
        RECT 17.070 96.300 17.995 96.310 ;
        RECT 17.075 96.295 17.995 96.300 ;
        RECT 17.085 96.280 17.995 96.295 ;
        RECT 17.090 96.265 17.995 96.280 ;
        RECT 17.100 96.240 17.995 96.265 ;
        RECT 16.605 95.770 16.935 96.195 ;
        RECT 14.805 95.275 15.695 95.445 ;
        RECT 15.865 95.235 16.125 95.715 ;
        RECT 16.295 95.065 16.545 95.605 ;
        RECT 16.715 95.285 16.935 95.770 ;
        RECT 17.105 96.170 17.995 96.240 ;
        RECT 17.105 95.445 17.275 96.170 ;
        RECT 18.625 96.055 18.975 96.305 ;
        RECT 17.445 95.615 17.995 96.000 ;
        RECT 19.145 95.875 19.315 96.475 ;
        RECT 19.485 96.055 19.835 96.305 ;
        RECT 20.005 96.055 20.350 96.625 ;
        RECT 20.520 96.305 20.695 97.405 ;
        RECT 20.865 97.035 21.195 97.270 ;
        RECT 21.485 97.215 21.885 97.615 ;
        RECT 22.755 97.215 23.085 97.615 ;
        RECT 20.865 96.865 22.945 97.035 ;
        RECT 20.865 96.475 21.420 96.865 ;
        RECT 20.520 96.055 21.080 96.305 ;
        RECT 21.250 96.225 21.420 96.475 ;
        RECT 21.590 96.475 22.605 96.695 ;
        RECT 22.775 96.595 22.945 96.865 ;
        RECT 23.255 96.775 23.515 97.445 ;
        RECT 21.590 96.335 21.865 96.475 ;
        RECT 22.775 96.425 23.170 96.595 ;
        RECT 21.250 96.055 21.445 96.225 ;
        RECT 17.105 95.275 17.995 95.445 ;
        RECT 18.635 95.065 18.905 95.875 ;
        RECT 19.075 95.235 19.405 95.875 ;
        RECT 19.575 95.065 19.815 95.875 ;
        RECT 20.005 95.705 21.105 95.885 ;
        RECT 20.005 95.300 20.345 95.705 ;
        RECT 20.515 95.065 20.685 95.535 ;
        RECT 20.855 95.300 21.105 95.705 ;
        RECT 21.275 95.670 21.445 96.055 ;
        RECT 21.275 95.300 21.525 95.670 ;
        RECT 21.695 95.545 21.865 96.335 ;
        RECT 22.035 95.885 22.210 96.080 ;
        RECT 22.380 96.055 22.830 96.255 ;
        RECT 23.000 95.975 23.170 96.425 ;
        RECT 22.035 95.715 22.530 95.885 ;
        RECT 23.340 95.805 23.515 96.775 ;
        RECT 23.685 96.475 23.945 97.615 ;
        RECT 24.115 96.465 24.445 97.445 ;
        RECT 24.615 96.475 24.895 97.615 ;
        RECT 23.705 96.055 24.040 96.305 ;
        RECT 24.210 95.865 24.380 96.465 ;
        RECT 25.065 96.450 25.355 97.615 ;
        RECT 25.565 96.475 25.795 97.615 ;
        RECT 25.965 96.465 26.295 97.445 ;
        RECT 26.465 96.475 26.675 97.615 ;
        RECT 26.905 96.525 28.575 97.615 ;
        RECT 24.550 96.035 24.885 96.305 ;
        RECT 25.545 96.055 25.875 96.305 ;
        RECT 22.310 95.575 22.530 95.715 ;
        RECT 21.695 95.375 22.140 95.545 ;
        RECT 22.310 95.405 22.535 95.575 ;
        RECT 22.310 95.360 22.530 95.405 ;
        RECT 22.810 95.065 22.980 95.730 ;
        RECT 23.175 95.235 23.515 95.805 ;
        RECT 23.685 95.235 24.380 95.865 ;
        RECT 24.585 95.065 24.895 95.865 ;
        RECT 25.065 95.065 25.355 95.790 ;
        RECT 25.565 95.065 25.795 95.885 ;
        RECT 26.045 95.865 26.295 96.465 ;
        RECT 25.965 95.235 26.295 95.865 ;
        RECT 26.465 95.065 26.675 95.885 ;
        RECT 26.905 95.835 27.655 96.355 ;
        RECT 27.825 96.005 28.575 96.525 ;
        RECT 29.240 96.825 29.775 97.445 ;
        RECT 26.905 95.065 28.575 95.835 ;
        RECT 29.240 95.805 29.555 96.825 ;
        RECT 29.945 96.815 30.275 97.615 ;
        RECT 30.760 96.645 31.150 96.820 ;
        RECT 32.920 96.815 33.170 97.615 ;
        RECT 33.340 96.985 33.670 97.445 ;
        RECT 33.840 97.155 34.055 97.615 ;
        RECT 34.725 97.180 40.070 97.615 ;
        RECT 33.340 96.815 34.510 96.985 ;
        RECT 29.725 96.475 31.150 96.645 ;
        RECT 32.430 96.645 32.710 96.805 ;
        RECT 32.430 96.475 33.765 96.645 ;
        RECT 29.725 95.975 29.895 96.475 ;
        RECT 29.240 95.235 29.855 95.805 ;
        RECT 30.145 95.745 30.410 96.305 ;
        RECT 30.580 95.575 30.750 96.475 ;
        RECT 33.595 96.305 33.765 96.475 ;
        RECT 30.920 95.745 31.275 96.305 ;
        RECT 32.430 96.055 32.780 96.295 ;
        RECT 32.950 96.055 33.425 96.295 ;
        RECT 33.595 96.055 33.970 96.305 ;
        RECT 33.595 95.885 33.765 96.055 ;
        RECT 32.430 95.715 33.765 95.885 ;
        RECT 30.025 95.065 30.240 95.575 ;
        RECT 30.470 95.245 30.750 95.575 ;
        RECT 30.930 95.065 31.170 95.575 ;
        RECT 32.430 95.505 32.700 95.715 ;
        RECT 34.140 95.525 34.510 96.815 ;
        RECT 36.310 95.610 36.650 96.440 ;
        RECT 38.130 95.930 38.480 97.180 ;
        RECT 40.245 96.525 42.835 97.615 ;
        RECT 40.245 95.835 41.455 96.355 ;
        RECT 41.625 96.005 42.835 96.525 ;
        RECT 43.015 96.645 43.345 97.430 ;
        RECT 43.015 96.475 43.695 96.645 ;
        RECT 43.875 96.475 44.205 97.615 ;
        RECT 44.385 96.765 44.645 97.445 ;
        RECT 44.815 96.835 45.065 97.615 ;
        RECT 45.315 97.065 45.565 97.445 ;
        RECT 45.735 97.235 46.090 97.615 ;
        RECT 47.095 97.225 47.430 97.445 ;
        RECT 46.695 97.065 46.925 97.105 ;
        RECT 45.315 96.865 46.925 97.065 ;
        RECT 45.315 96.855 46.150 96.865 ;
        RECT 46.740 96.775 46.925 96.865 ;
        RECT 43.005 96.055 43.355 96.305 ;
        RECT 43.525 95.875 43.695 96.475 ;
        RECT 43.865 96.055 44.215 96.305 ;
        RECT 32.920 95.065 33.250 95.525 ;
        RECT 33.760 95.235 34.510 95.525 ;
        RECT 34.725 95.065 40.070 95.610 ;
        RECT 40.245 95.065 42.835 95.835 ;
        RECT 43.025 95.065 43.265 95.875 ;
        RECT 43.435 95.235 43.765 95.875 ;
        RECT 43.935 95.065 44.205 95.875 ;
        RECT 44.385 95.565 44.555 96.765 ;
        RECT 46.255 96.665 46.585 96.695 ;
        RECT 44.785 96.605 46.585 96.665 ;
        RECT 47.175 96.605 47.430 97.225 ;
        RECT 44.725 96.495 47.430 96.605 ;
        RECT 44.725 96.460 44.925 96.495 ;
        RECT 44.725 95.885 44.895 96.460 ;
        RECT 46.255 96.435 47.430 96.495 ;
        RECT 45.125 96.020 45.535 96.325 ;
        RECT 45.705 96.055 46.035 96.265 ;
        RECT 44.725 95.765 44.995 95.885 ;
        RECT 44.725 95.720 45.570 95.765 ;
        RECT 44.815 95.595 45.570 95.720 ;
        RECT 45.825 95.655 46.035 96.055 ;
        RECT 46.280 96.055 46.755 96.265 ;
        RECT 46.945 96.055 47.435 96.255 ;
        RECT 46.280 95.655 46.500 96.055 ;
        RECT 47.605 96.010 47.885 97.445 ;
        RECT 48.055 96.840 48.765 97.615 ;
        RECT 48.935 96.670 49.265 97.445 ;
        RECT 48.115 96.455 49.265 96.670 ;
        RECT 44.385 95.235 44.645 95.565 ;
        RECT 45.400 95.445 45.570 95.595 ;
        RECT 44.815 95.065 45.145 95.425 ;
        RECT 45.400 95.235 46.700 95.445 ;
        RECT 46.975 95.065 47.430 95.830 ;
        RECT 47.605 95.235 47.945 96.010 ;
        RECT 48.115 95.885 48.400 96.455 ;
        RECT 48.585 96.055 49.055 96.285 ;
        RECT 49.460 96.255 49.675 97.370 ;
        RECT 49.855 96.895 50.185 97.615 ;
        RECT 49.965 96.255 50.195 96.595 ;
        RECT 50.825 96.450 51.115 97.615 ;
        RECT 51.295 96.805 51.590 97.615 ;
        RECT 51.770 96.305 52.015 97.445 ;
        RECT 52.190 96.805 52.450 97.615 ;
        RECT 53.050 97.610 59.325 97.615 ;
        RECT 52.630 96.305 52.880 97.440 ;
        RECT 53.050 96.815 53.310 97.610 ;
        RECT 53.480 96.715 53.740 97.440 ;
        RECT 53.910 96.885 54.170 97.610 ;
        RECT 54.340 96.715 54.600 97.440 ;
        RECT 54.770 96.885 55.030 97.610 ;
        RECT 55.200 96.715 55.460 97.440 ;
        RECT 55.630 96.885 55.890 97.610 ;
        RECT 56.060 96.715 56.320 97.440 ;
        RECT 56.490 96.885 56.735 97.610 ;
        RECT 56.905 96.715 57.165 97.440 ;
        RECT 57.350 96.885 57.595 97.610 ;
        RECT 57.765 96.715 58.025 97.440 ;
        RECT 58.210 96.885 58.455 97.610 ;
        RECT 58.625 96.715 58.885 97.440 ;
        RECT 59.070 96.885 59.325 97.610 ;
        RECT 53.480 96.700 58.885 96.715 ;
        RECT 59.495 96.700 59.785 97.440 ;
        RECT 59.955 96.870 60.225 97.615 ;
        RECT 60.485 97.180 65.830 97.615 ;
        RECT 53.480 96.475 60.225 96.700 ;
        RECT 49.225 96.075 49.675 96.255 ;
        RECT 49.225 96.055 49.555 96.075 ;
        RECT 49.865 96.055 50.195 96.255 ;
        RECT 48.115 95.695 48.825 95.885 ;
        RECT 48.525 95.555 48.825 95.695 ;
        RECT 49.015 95.695 50.195 95.885 ;
        RECT 49.015 95.615 49.345 95.695 ;
        RECT 48.525 95.545 48.840 95.555 ;
        RECT 48.525 95.535 48.850 95.545 ;
        RECT 48.525 95.530 48.860 95.535 ;
        RECT 48.115 95.065 48.285 95.525 ;
        RECT 48.525 95.520 48.865 95.530 ;
        RECT 48.525 95.515 48.870 95.520 ;
        RECT 48.525 95.505 48.875 95.515 ;
        RECT 48.525 95.500 48.880 95.505 ;
        RECT 48.525 95.235 48.885 95.500 ;
        RECT 49.515 95.065 49.685 95.525 ;
        RECT 49.855 95.235 50.195 95.695 ;
        RECT 50.825 95.065 51.115 95.790 ;
        RECT 51.285 95.745 51.600 96.305 ;
        RECT 51.770 96.055 58.890 96.305 ;
        RECT 51.285 95.065 51.590 95.575 ;
        RECT 51.770 95.245 52.020 96.055 ;
        RECT 52.190 95.065 52.450 95.590 ;
        RECT 52.630 95.245 52.880 96.055 ;
        RECT 59.060 95.885 60.225 96.475 ;
        RECT 53.480 95.715 60.225 95.885 ;
        RECT 53.050 95.065 53.310 95.625 ;
        RECT 53.480 95.260 53.740 95.715 ;
        RECT 53.910 95.065 54.170 95.545 ;
        RECT 54.340 95.260 54.600 95.715 ;
        RECT 54.770 95.065 55.030 95.545 ;
        RECT 55.200 95.260 55.460 95.715 ;
        RECT 55.630 95.065 55.875 95.545 ;
        RECT 56.045 95.260 56.320 95.715 ;
        RECT 56.490 95.065 56.735 95.545 ;
        RECT 56.905 95.260 57.165 95.715 ;
        RECT 57.345 95.065 57.595 95.545 ;
        RECT 57.765 95.260 58.025 95.715 ;
        RECT 58.205 95.065 58.455 95.545 ;
        RECT 58.625 95.260 58.885 95.715 ;
        RECT 59.065 95.065 59.325 95.545 ;
        RECT 59.495 95.260 59.755 95.715 ;
        RECT 62.070 95.610 62.410 96.440 ;
        RECT 63.890 95.930 64.240 97.180 ;
        RECT 66.005 96.525 67.675 97.615 ;
        RECT 66.005 95.835 66.755 96.355 ;
        RECT 66.925 96.005 67.675 96.525 ;
        RECT 67.850 96.475 68.185 97.445 ;
        RECT 68.355 96.475 68.525 97.615 ;
        RECT 68.695 97.275 70.725 97.445 ;
        RECT 59.925 95.065 60.225 95.545 ;
        RECT 60.485 95.065 65.830 95.610 ;
        RECT 66.005 95.065 67.675 95.835 ;
        RECT 67.850 95.805 68.020 96.475 ;
        RECT 68.695 96.305 68.865 97.275 ;
        RECT 68.190 95.975 68.445 96.305 ;
        RECT 68.670 95.975 68.865 96.305 ;
        RECT 69.035 96.935 70.160 97.105 ;
        RECT 68.275 95.805 68.445 95.975 ;
        RECT 69.035 95.805 69.205 96.935 ;
        RECT 67.850 95.235 68.105 95.805 ;
        RECT 68.275 95.635 69.205 95.805 ;
        RECT 69.375 96.595 70.385 96.765 ;
        RECT 69.375 95.795 69.545 96.595 ;
        RECT 69.750 96.255 70.025 96.395 ;
        RECT 69.745 96.085 70.025 96.255 ;
        RECT 69.030 95.600 69.205 95.635 ;
        RECT 68.275 95.065 68.605 95.465 ;
        RECT 69.030 95.235 69.560 95.600 ;
        RECT 69.750 95.235 70.025 96.085 ;
        RECT 70.195 95.235 70.385 96.595 ;
        RECT 70.555 96.610 70.725 97.275 ;
        RECT 70.895 96.855 71.065 97.615 ;
        RECT 71.300 96.855 71.815 97.265 ;
        RECT 70.555 96.420 71.305 96.610 ;
        RECT 71.475 96.045 71.815 96.855 ;
        RECT 71.985 96.525 73.195 97.615 ;
        RECT 70.585 95.875 71.815 96.045 ;
        RECT 70.565 95.065 71.075 95.600 ;
        RECT 71.295 95.270 71.540 95.875 ;
        RECT 71.985 95.815 72.505 96.355 ;
        RECT 72.675 95.985 73.195 96.525 ;
        RECT 73.365 96.765 73.625 97.445 ;
        RECT 73.795 96.835 74.045 97.615 ;
        RECT 74.295 97.065 74.545 97.445 ;
        RECT 74.715 97.235 75.070 97.615 ;
        RECT 76.075 97.225 76.410 97.445 ;
        RECT 75.675 97.065 75.905 97.105 ;
        RECT 74.295 96.865 75.905 97.065 ;
        RECT 74.295 96.855 75.130 96.865 ;
        RECT 75.720 96.775 75.905 96.865 ;
        RECT 71.985 95.065 73.195 95.815 ;
        RECT 73.365 95.575 73.535 96.765 ;
        RECT 75.235 96.665 75.565 96.695 ;
        RECT 73.765 96.605 75.565 96.665 ;
        RECT 76.155 96.605 76.410 97.225 ;
        RECT 73.705 96.495 76.410 96.605 ;
        RECT 73.705 96.460 73.905 96.495 ;
        RECT 73.705 95.885 73.875 96.460 ;
        RECT 75.235 96.435 76.410 96.495 ;
        RECT 76.585 96.450 76.875 97.615 ;
        RECT 77.135 96.685 77.305 97.445 ;
        RECT 77.485 96.855 77.815 97.615 ;
        RECT 77.135 96.515 77.800 96.685 ;
        RECT 77.985 96.540 78.255 97.445 ;
        RECT 77.630 96.370 77.800 96.515 ;
        RECT 74.105 96.020 74.515 96.325 ;
        RECT 74.685 96.055 75.015 96.265 ;
        RECT 73.705 95.765 73.975 95.885 ;
        RECT 73.705 95.720 74.550 95.765 ;
        RECT 73.795 95.595 74.550 95.720 ;
        RECT 74.805 95.655 75.015 96.055 ;
        RECT 75.260 96.055 75.735 96.265 ;
        RECT 75.925 96.055 76.415 96.255 ;
        RECT 75.260 95.655 75.480 96.055 ;
        RECT 77.065 95.965 77.395 96.335 ;
        RECT 77.630 96.040 77.915 96.370 ;
        RECT 73.365 95.565 73.595 95.575 ;
        RECT 73.365 95.235 73.625 95.565 ;
        RECT 74.380 95.445 74.550 95.595 ;
        RECT 73.795 95.065 74.125 95.425 ;
        RECT 74.380 95.235 75.680 95.445 ;
        RECT 75.955 95.065 76.410 95.830 ;
        RECT 76.585 95.065 76.875 95.790 ;
        RECT 77.630 95.785 77.800 96.040 ;
        RECT 77.135 95.615 77.800 95.785 ;
        RECT 78.085 95.740 78.255 96.540 ;
        RECT 77.135 95.235 77.305 95.615 ;
        RECT 77.485 95.065 77.815 95.445 ;
        RECT 77.995 95.235 78.255 95.740 ;
        RECT 78.425 96.475 78.765 97.445 ;
        RECT 78.935 96.475 79.105 97.615 ;
        RECT 79.375 96.815 79.625 97.615 ;
        RECT 80.270 96.645 80.600 97.445 ;
        RECT 80.900 96.815 81.230 97.615 ;
        RECT 81.400 96.645 81.730 97.445 ;
        RECT 79.295 96.475 81.730 96.645 ;
        RECT 82.140 96.825 82.675 97.445 ;
        RECT 78.425 95.865 78.600 96.475 ;
        RECT 79.295 96.225 79.465 96.475 ;
        RECT 78.770 96.055 79.465 96.225 ;
        RECT 79.640 96.055 80.060 96.255 ;
        RECT 80.230 96.055 80.560 96.255 ;
        RECT 80.730 96.055 81.060 96.255 ;
        RECT 78.425 95.235 78.765 95.865 ;
        RECT 78.935 95.065 79.185 95.865 ;
        RECT 79.375 95.715 80.600 95.885 ;
        RECT 79.375 95.235 79.705 95.715 ;
        RECT 79.875 95.065 80.100 95.525 ;
        RECT 80.270 95.235 80.600 95.715 ;
        RECT 81.230 95.845 81.400 96.475 ;
        RECT 81.585 96.055 81.935 96.305 ;
        RECT 81.230 95.235 81.730 95.845 ;
        RECT 82.140 95.805 82.455 96.825 ;
        RECT 82.845 96.815 83.175 97.615 ;
        RECT 83.660 96.645 84.050 96.820 ;
        RECT 82.625 96.475 84.050 96.645 ;
        RECT 84.590 96.645 84.980 96.820 ;
        RECT 85.465 96.815 85.795 97.615 ;
        RECT 85.965 96.825 86.500 97.445 ;
        RECT 84.590 96.475 86.015 96.645 ;
        RECT 82.625 95.975 82.795 96.475 ;
        RECT 82.140 95.235 82.755 95.805 ;
        RECT 83.045 95.745 83.310 96.305 ;
        RECT 83.480 95.575 83.650 96.475 ;
        RECT 83.820 95.745 84.175 96.305 ;
        RECT 84.465 95.745 84.820 96.305 ;
        RECT 84.990 95.575 85.160 96.475 ;
        RECT 85.330 95.745 85.595 96.305 ;
        RECT 85.845 95.975 86.015 96.475 ;
        RECT 86.185 95.805 86.500 96.825 ;
        RECT 86.710 96.465 86.970 97.615 ;
        RECT 87.145 96.540 87.400 97.445 ;
        RECT 87.570 96.855 87.900 97.615 ;
        RECT 88.115 96.685 88.285 97.445 ;
        RECT 82.925 95.065 83.140 95.575 ;
        RECT 83.370 95.245 83.650 95.575 ;
        RECT 83.830 95.065 84.070 95.575 ;
        RECT 84.570 95.065 84.810 95.575 ;
        RECT 84.990 95.245 85.270 95.575 ;
        RECT 85.500 95.065 85.715 95.575 ;
        RECT 85.885 95.235 86.500 95.805 ;
        RECT 86.710 95.065 86.970 95.905 ;
        RECT 87.145 95.810 87.315 96.540 ;
        RECT 87.570 96.515 88.285 96.685 ;
        RECT 88.545 96.525 89.755 97.615 ;
        RECT 87.570 96.305 87.740 96.515 ;
        RECT 87.485 95.975 87.740 96.305 ;
        RECT 87.145 95.235 87.400 95.810 ;
        RECT 87.570 95.785 87.740 95.975 ;
        RECT 88.020 95.965 88.375 96.335 ;
        RECT 88.545 95.985 89.065 96.525 ;
        RECT 89.235 95.815 89.755 96.355 ;
        RECT 87.570 95.615 88.285 95.785 ;
        RECT 87.570 95.065 87.900 95.445 ;
        RECT 88.115 95.235 88.285 95.615 ;
        RECT 88.545 95.065 89.755 95.815 ;
        RECT 12.100 94.895 89.840 95.065 ;
        RECT 12.185 94.145 13.395 94.895 ;
        RECT 14.575 94.345 14.745 94.635 ;
        RECT 14.915 94.515 15.245 94.895 ;
        RECT 14.575 94.175 15.240 94.345 ;
        RECT 12.185 93.605 12.705 94.145 ;
        RECT 12.875 93.435 13.395 93.975 ;
        RECT 12.185 92.345 13.395 93.435 ;
        RECT 14.490 93.355 14.840 94.005 ;
        RECT 15.010 93.185 15.240 94.175 ;
        RECT 14.575 93.015 15.240 93.185 ;
        RECT 14.575 92.515 14.745 93.015 ;
        RECT 14.915 92.345 15.245 92.845 ;
        RECT 15.415 92.515 15.600 94.635 ;
        RECT 15.855 94.435 16.105 94.895 ;
        RECT 16.275 94.445 16.610 94.615 ;
        RECT 16.805 94.445 17.480 94.615 ;
        RECT 16.275 94.305 16.445 94.445 ;
        RECT 15.770 93.315 16.050 94.265 ;
        RECT 16.220 94.175 16.445 94.305 ;
        RECT 16.220 93.070 16.390 94.175 ;
        RECT 16.615 94.025 17.140 94.245 ;
        RECT 16.560 93.260 16.800 93.855 ;
        RECT 16.970 93.325 17.140 94.025 ;
        RECT 17.310 93.665 17.480 94.445 ;
        RECT 17.800 94.395 18.170 94.895 ;
        RECT 18.350 94.445 18.755 94.615 ;
        RECT 18.925 94.445 19.710 94.615 ;
        RECT 18.350 94.215 18.520 94.445 ;
        RECT 17.690 93.915 18.520 94.215 ;
        RECT 18.905 93.945 19.370 94.275 ;
        RECT 17.690 93.885 17.890 93.915 ;
        RECT 18.010 93.665 18.180 93.735 ;
        RECT 17.310 93.495 18.180 93.665 ;
        RECT 17.670 93.405 18.180 93.495 ;
        RECT 16.220 92.940 16.525 93.070 ;
        RECT 16.970 92.960 17.500 93.325 ;
        RECT 15.840 92.345 16.105 92.805 ;
        RECT 16.275 92.515 16.525 92.940 ;
        RECT 17.670 92.790 17.840 93.405 ;
        RECT 16.735 92.620 17.840 92.790 ;
        RECT 18.010 92.345 18.180 93.145 ;
        RECT 18.350 92.845 18.520 93.915 ;
        RECT 18.690 93.015 18.880 93.735 ;
        RECT 19.050 92.985 19.370 93.945 ;
        RECT 19.540 93.985 19.710 94.445 ;
        RECT 19.985 94.365 20.195 94.895 ;
        RECT 20.455 94.155 20.785 94.680 ;
        RECT 20.955 94.285 21.125 94.895 ;
        RECT 21.295 94.240 21.625 94.675 ;
        RECT 21.295 94.155 21.675 94.240 ;
        RECT 20.585 93.985 20.785 94.155 ;
        RECT 21.450 94.115 21.675 94.155 ;
        RECT 19.540 93.655 20.415 93.985 ;
        RECT 20.585 93.655 21.335 93.985 ;
        RECT 18.350 92.515 18.600 92.845 ;
        RECT 19.540 92.815 19.710 93.655 ;
        RECT 20.585 93.450 20.775 93.655 ;
        RECT 21.505 93.535 21.675 94.115 ;
        RECT 22.315 94.085 22.585 94.895 ;
        RECT 22.755 94.085 23.085 94.725 ;
        RECT 23.255 94.085 23.495 94.895 ;
        RECT 23.775 94.345 23.945 94.635 ;
        RECT 24.115 94.515 24.445 94.895 ;
        RECT 23.775 94.175 24.440 94.345 ;
        RECT 22.305 93.655 22.655 93.905 ;
        RECT 21.460 93.485 21.675 93.535 ;
        RECT 22.825 93.485 22.995 94.085 ;
        RECT 23.165 93.655 23.515 93.905 ;
        RECT 19.880 93.075 20.775 93.450 ;
        RECT 21.285 93.405 21.675 93.485 ;
        RECT 18.825 92.645 19.710 92.815 ;
        RECT 19.890 92.345 20.205 92.845 ;
        RECT 20.435 92.515 20.775 93.075 ;
        RECT 20.945 92.345 21.115 93.355 ;
        RECT 21.285 92.560 21.615 93.405 ;
        RECT 22.315 92.345 22.645 93.485 ;
        RECT 22.825 93.315 23.505 93.485 ;
        RECT 23.690 93.355 24.040 94.005 ;
        RECT 23.175 92.530 23.505 93.315 ;
        RECT 24.210 93.185 24.440 94.175 ;
        RECT 23.775 93.015 24.440 93.185 ;
        RECT 23.775 92.515 23.945 93.015 ;
        RECT 24.115 92.345 24.445 92.845 ;
        RECT 24.615 92.515 24.800 94.635 ;
        RECT 25.055 94.435 25.305 94.895 ;
        RECT 25.475 94.445 25.810 94.615 ;
        RECT 26.005 94.445 26.680 94.615 ;
        RECT 25.475 94.305 25.645 94.445 ;
        RECT 24.970 93.315 25.250 94.265 ;
        RECT 25.420 94.175 25.645 94.305 ;
        RECT 25.420 93.070 25.590 94.175 ;
        RECT 25.815 94.025 26.340 94.245 ;
        RECT 25.760 93.260 26.000 93.855 ;
        RECT 26.170 93.325 26.340 94.025 ;
        RECT 26.510 93.665 26.680 94.445 ;
        RECT 27.000 94.395 27.370 94.895 ;
        RECT 27.550 94.445 27.955 94.615 ;
        RECT 28.125 94.445 28.910 94.615 ;
        RECT 27.550 94.215 27.720 94.445 ;
        RECT 26.890 93.915 27.720 94.215 ;
        RECT 28.105 93.945 28.570 94.275 ;
        RECT 26.890 93.885 27.090 93.915 ;
        RECT 27.210 93.665 27.380 93.735 ;
        RECT 26.510 93.495 27.380 93.665 ;
        RECT 26.870 93.405 27.380 93.495 ;
        RECT 25.420 92.940 25.725 93.070 ;
        RECT 26.170 92.960 26.700 93.325 ;
        RECT 25.040 92.345 25.305 92.805 ;
        RECT 25.475 92.515 25.725 92.940 ;
        RECT 26.870 92.790 27.040 93.405 ;
        RECT 25.935 92.620 27.040 92.790 ;
        RECT 27.210 92.345 27.380 93.145 ;
        RECT 27.550 92.845 27.720 93.915 ;
        RECT 27.890 93.015 28.080 93.735 ;
        RECT 28.250 92.985 28.570 93.945 ;
        RECT 28.740 93.985 28.910 94.445 ;
        RECT 29.185 94.365 29.395 94.895 ;
        RECT 29.655 94.155 29.985 94.680 ;
        RECT 30.155 94.285 30.325 94.895 ;
        RECT 30.495 94.240 30.825 94.675 ;
        RECT 30.495 94.155 30.875 94.240 ;
        RECT 29.785 93.985 29.985 94.155 ;
        RECT 30.650 94.115 30.875 94.155 ;
        RECT 28.740 93.655 29.615 93.985 ;
        RECT 29.785 93.655 30.535 93.985 ;
        RECT 27.550 92.515 27.800 92.845 ;
        RECT 28.740 92.815 28.910 93.655 ;
        RECT 29.785 93.450 29.975 93.655 ;
        RECT 30.705 93.535 30.875 94.115 ;
        RECT 31.045 94.145 32.255 94.895 ;
        RECT 32.425 94.515 33.315 94.685 ;
        RECT 31.045 93.605 31.565 94.145 ;
        RECT 30.660 93.485 30.875 93.535 ;
        RECT 29.080 93.075 29.975 93.450 ;
        RECT 30.485 93.405 30.875 93.485 ;
        RECT 31.735 93.435 32.255 93.975 ;
        RECT 32.425 93.960 32.975 94.345 ;
        RECT 33.145 93.790 33.315 94.515 ;
        RECT 28.025 92.645 28.910 92.815 ;
        RECT 29.090 92.345 29.405 92.845 ;
        RECT 29.635 92.515 29.975 93.075 ;
        RECT 30.145 92.345 30.315 93.355 ;
        RECT 30.485 92.560 30.815 93.405 ;
        RECT 31.045 92.345 32.255 93.435 ;
        RECT 32.425 93.720 33.315 93.790 ;
        RECT 33.485 94.190 33.705 94.675 ;
        RECT 33.875 94.355 34.125 94.895 ;
        RECT 34.295 94.245 34.555 94.725 ;
        RECT 33.485 93.765 33.815 94.190 ;
        RECT 32.425 93.695 33.320 93.720 ;
        RECT 32.425 93.680 33.330 93.695 ;
        RECT 32.425 93.665 33.335 93.680 ;
        RECT 32.425 93.660 33.345 93.665 ;
        RECT 32.425 93.650 33.350 93.660 ;
        RECT 32.425 93.640 33.355 93.650 ;
        RECT 32.425 93.635 33.365 93.640 ;
        RECT 32.425 93.625 33.375 93.635 ;
        RECT 32.425 93.620 33.385 93.625 ;
        RECT 32.425 93.170 32.685 93.620 ;
        RECT 33.050 93.615 33.385 93.620 ;
        RECT 33.050 93.610 33.400 93.615 ;
        RECT 33.050 93.600 33.415 93.610 ;
        RECT 33.050 93.595 33.440 93.600 ;
        RECT 33.985 93.595 34.215 93.990 ;
        RECT 33.050 93.590 34.215 93.595 ;
        RECT 33.080 93.555 34.215 93.590 ;
        RECT 33.115 93.530 34.215 93.555 ;
        RECT 33.145 93.500 34.215 93.530 ;
        RECT 33.165 93.470 34.215 93.500 ;
        RECT 33.185 93.440 34.215 93.470 ;
        RECT 33.255 93.430 34.215 93.440 ;
        RECT 33.280 93.420 34.215 93.430 ;
        RECT 33.300 93.405 34.215 93.420 ;
        RECT 33.320 93.390 34.215 93.405 ;
        RECT 33.325 93.380 34.110 93.390 ;
        RECT 33.340 93.345 34.110 93.380 ;
        RECT 32.855 93.025 33.185 93.270 ;
        RECT 33.355 93.095 34.110 93.345 ;
        RECT 34.385 93.215 34.555 94.245 ;
        RECT 34.745 94.165 35.035 94.895 ;
        RECT 34.735 93.655 35.035 93.985 ;
        RECT 35.215 93.965 35.445 94.605 ;
        RECT 35.625 94.345 35.935 94.715 ;
        RECT 36.115 94.525 36.785 94.895 ;
        RECT 35.625 94.145 36.855 94.345 ;
        RECT 35.215 93.655 35.740 93.965 ;
        RECT 35.920 93.655 36.385 93.965 ;
        RECT 36.565 93.475 36.855 94.145 ;
        RECT 32.855 93.000 33.040 93.025 ;
        RECT 32.425 92.900 33.040 93.000 ;
        RECT 32.425 92.345 33.030 92.900 ;
        RECT 33.205 92.515 33.685 92.855 ;
        RECT 33.855 92.345 34.110 92.890 ;
        RECT 34.280 92.515 34.555 93.215 ;
        RECT 34.745 93.235 35.905 93.475 ;
        RECT 34.745 92.525 35.005 93.235 ;
        RECT 35.175 92.345 35.505 93.055 ;
        RECT 35.675 92.525 35.905 93.235 ;
        RECT 36.085 93.255 36.855 93.475 ;
        RECT 36.085 92.525 36.355 93.255 ;
        RECT 36.535 92.345 36.875 93.075 ;
        RECT 37.045 92.525 37.305 94.715 ;
        RECT 37.945 94.170 38.235 94.895 ;
        RECT 38.405 94.350 43.750 94.895 ;
        RECT 39.990 93.520 40.330 94.350 ;
        RECT 43.925 94.125 47.435 94.895 ;
        RECT 47.605 94.145 48.815 94.895 ;
        RECT 49.000 94.325 49.255 94.675 ;
        RECT 49.425 94.495 49.755 94.895 ;
        RECT 49.925 94.325 50.095 94.675 ;
        RECT 50.265 94.495 50.645 94.895 ;
        RECT 49.000 94.155 50.665 94.325 ;
        RECT 50.835 94.220 51.110 94.565 ;
        RECT 37.945 92.345 38.235 93.510 ;
        RECT 41.810 92.780 42.160 94.030 ;
        RECT 43.925 93.605 45.575 94.125 ;
        RECT 45.745 93.435 47.435 93.955 ;
        RECT 47.605 93.605 48.125 94.145 ;
        RECT 50.495 93.985 50.665 94.155 ;
        RECT 48.295 93.435 48.815 93.975 ;
        RECT 48.985 93.655 49.330 93.985 ;
        RECT 49.500 93.655 50.325 93.985 ;
        RECT 50.495 93.655 50.770 93.985 ;
        RECT 38.405 92.345 43.750 92.780 ;
        RECT 43.925 92.345 47.435 93.435 ;
        RECT 47.605 92.345 48.815 93.435 ;
        RECT 49.005 93.195 49.330 93.485 ;
        RECT 49.500 93.365 49.695 93.655 ;
        RECT 50.495 93.485 50.665 93.655 ;
        RECT 50.940 93.485 51.110 94.220 ;
        RECT 51.345 94.075 51.555 94.895 ;
        RECT 51.725 94.095 52.055 94.725 ;
        RECT 51.725 93.495 51.975 94.095 ;
        RECT 52.225 94.075 52.455 94.895 ;
        RECT 52.710 94.435 53.460 94.725 ;
        RECT 53.970 94.435 54.300 94.895 ;
        RECT 52.145 93.655 52.475 93.905 ;
        RECT 50.005 93.315 50.665 93.485 ;
        RECT 50.005 93.195 50.175 93.315 ;
        RECT 49.005 93.025 50.175 93.195 ;
        RECT 48.985 92.565 50.175 92.855 ;
        RECT 50.345 92.345 50.625 93.145 ;
        RECT 50.835 92.515 51.110 93.485 ;
        RECT 51.345 92.345 51.555 93.485 ;
        RECT 51.725 92.515 52.055 93.495 ;
        RECT 52.225 92.345 52.455 93.485 ;
        RECT 52.710 93.145 53.080 94.435 ;
        RECT 54.520 94.245 54.790 94.455 ;
        RECT 53.455 94.075 54.790 94.245 ;
        RECT 54.965 94.145 56.175 94.895 ;
        RECT 56.365 94.385 56.605 94.895 ;
        RECT 56.775 94.385 57.065 94.725 ;
        RECT 57.295 94.385 57.610 94.895 ;
        RECT 53.455 93.905 53.625 94.075 ;
        RECT 53.250 93.655 53.625 93.905 ;
        RECT 53.795 93.665 54.270 93.905 ;
        RECT 54.440 93.665 54.790 93.905 ;
        RECT 53.455 93.485 53.625 93.655 ;
        RECT 54.965 93.605 55.485 94.145 ;
        RECT 56.405 94.045 56.605 94.215 ;
        RECT 53.455 93.315 54.790 93.485 ;
        RECT 55.655 93.435 56.175 93.975 ;
        RECT 56.410 93.655 56.605 94.045 ;
        RECT 56.775 93.485 56.955 94.385 ;
        RECT 57.780 94.325 57.950 94.595 ;
        RECT 58.120 94.495 58.450 94.895 ;
        RECT 57.125 93.655 57.535 94.215 ;
        RECT 57.780 94.155 58.475 94.325 ;
        RECT 57.705 93.485 57.875 93.985 ;
        RECT 54.510 93.155 54.790 93.315 ;
        RECT 52.710 92.975 53.880 93.145 ;
        RECT 53.165 92.345 53.380 92.805 ;
        RECT 53.550 92.515 53.880 92.975 ;
        RECT 54.050 92.345 54.300 93.145 ;
        RECT 54.965 92.345 56.175 93.435 ;
        RECT 56.415 93.315 57.875 93.485 ;
        RECT 56.415 93.140 56.775 93.315 ;
        RECT 58.045 93.145 58.475 94.155 ;
        RECT 58.650 94.075 58.925 94.895 ;
        RECT 59.095 94.255 59.425 94.725 ;
        RECT 59.595 94.425 59.765 94.895 ;
        RECT 59.935 94.255 60.265 94.725 ;
        RECT 60.435 94.425 60.725 94.895 ;
        RECT 59.095 94.245 60.265 94.255 ;
        RECT 59.095 94.075 60.695 94.245 ;
        RECT 60.950 94.075 61.225 94.895 ;
        RECT 61.395 94.255 61.725 94.725 ;
        RECT 61.895 94.425 62.065 94.895 ;
        RECT 62.235 94.255 62.565 94.725 ;
        RECT 62.735 94.425 63.025 94.895 ;
        RECT 61.395 94.245 62.565 94.255 ;
        RECT 61.395 94.075 62.995 94.245 ;
        RECT 63.705 94.170 63.995 94.895 ;
        RECT 64.165 94.350 69.510 94.895 ;
        RECT 58.650 93.705 59.370 93.905 ;
        RECT 59.540 93.705 60.310 93.905 ;
        RECT 60.480 93.535 60.695 94.075 ;
        RECT 60.950 93.705 61.670 93.905 ;
        RECT 61.840 93.705 62.610 93.905 ;
        RECT 62.780 93.535 62.995 94.075 ;
        RECT 57.360 92.345 57.530 93.145 ;
        RECT 57.700 92.975 58.475 93.145 ;
        RECT 58.650 93.315 59.765 93.525 ;
        RECT 57.700 92.515 58.030 92.975 ;
        RECT 58.200 92.345 58.370 92.805 ;
        RECT 58.650 92.515 58.925 93.315 ;
        RECT 59.095 92.345 59.425 93.145 ;
        RECT 59.595 92.685 59.765 93.315 ;
        RECT 59.935 93.315 60.695 93.535 ;
        RECT 60.950 93.315 62.065 93.525 ;
        RECT 59.935 92.855 60.265 93.315 ;
        RECT 60.435 92.685 60.735 93.145 ;
        RECT 59.595 92.515 60.735 92.685 ;
        RECT 60.950 92.515 61.225 93.315 ;
        RECT 61.395 92.345 61.725 93.145 ;
        RECT 61.895 92.685 62.065 93.315 ;
        RECT 62.235 93.365 63.015 93.535 ;
        RECT 65.750 93.520 66.090 94.350 ;
        RECT 69.685 94.125 71.355 94.895 ;
        RECT 62.235 93.315 62.995 93.365 ;
        RECT 62.235 92.855 62.565 93.315 ;
        RECT 62.735 92.685 63.035 93.145 ;
        RECT 61.895 92.515 63.035 92.685 ;
        RECT 63.705 92.345 63.995 93.510 ;
        RECT 67.570 92.780 67.920 94.030 ;
        RECT 69.685 93.605 70.435 94.125 ;
        RECT 71.530 94.055 71.790 94.895 ;
        RECT 71.965 94.150 72.220 94.725 ;
        RECT 72.390 94.515 72.720 94.895 ;
        RECT 72.935 94.345 73.105 94.725 ;
        RECT 72.390 94.175 73.105 94.345 ;
        RECT 70.605 93.435 71.355 93.955 ;
        RECT 64.165 92.345 69.510 92.780 ;
        RECT 69.685 92.345 71.355 93.435 ;
        RECT 71.530 92.345 71.790 93.495 ;
        RECT 71.965 93.420 72.135 94.150 ;
        RECT 72.390 93.985 72.560 94.175 ;
        RECT 73.370 94.055 73.630 94.895 ;
        RECT 73.805 94.150 74.060 94.725 ;
        RECT 74.230 94.515 74.560 94.895 ;
        RECT 74.775 94.345 74.945 94.725 ;
        RECT 74.230 94.175 74.945 94.345 ;
        RECT 72.305 93.655 72.560 93.985 ;
        RECT 72.390 93.445 72.560 93.655 ;
        RECT 72.840 93.625 73.195 93.995 ;
        RECT 71.965 92.515 72.220 93.420 ;
        RECT 72.390 93.275 73.105 93.445 ;
        RECT 72.390 92.345 72.720 93.105 ;
        RECT 72.935 92.515 73.105 93.275 ;
        RECT 73.370 92.345 73.630 93.495 ;
        RECT 73.805 93.420 73.975 94.150 ;
        RECT 74.230 93.985 74.400 94.175 ;
        RECT 75.210 94.055 75.470 94.895 ;
        RECT 75.645 94.150 75.900 94.725 ;
        RECT 76.070 94.515 76.400 94.895 ;
        RECT 76.615 94.345 76.785 94.725 ;
        RECT 77.210 94.385 77.450 94.895 ;
        RECT 77.630 94.385 77.910 94.715 ;
        RECT 78.140 94.385 78.355 94.895 ;
        RECT 76.070 94.175 76.785 94.345 ;
        RECT 74.145 93.655 74.400 93.985 ;
        RECT 74.230 93.445 74.400 93.655 ;
        RECT 74.680 93.625 75.035 93.995 ;
        RECT 73.805 92.515 74.060 93.420 ;
        RECT 74.230 93.275 74.945 93.445 ;
        RECT 74.230 92.345 74.560 93.105 ;
        RECT 74.775 92.515 74.945 93.275 ;
        RECT 75.210 92.345 75.470 93.495 ;
        RECT 75.645 93.420 75.815 94.150 ;
        RECT 76.070 93.985 76.240 94.175 ;
        RECT 75.985 93.655 76.240 93.985 ;
        RECT 76.070 93.445 76.240 93.655 ;
        RECT 76.520 93.625 76.875 93.995 ;
        RECT 77.105 93.655 77.460 94.215 ;
        RECT 77.630 93.485 77.800 94.385 ;
        RECT 77.970 93.655 78.235 94.215 ;
        RECT 78.525 94.155 79.140 94.725 ;
        RECT 79.455 94.515 80.625 94.725 ;
        RECT 79.455 94.495 79.785 94.515 ;
        RECT 78.485 93.485 78.655 93.985 ;
        RECT 75.645 92.515 75.900 93.420 ;
        RECT 76.070 93.275 76.785 93.445 ;
        RECT 76.070 92.345 76.400 93.105 ;
        RECT 76.615 92.515 76.785 93.275 ;
        RECT 77.230 93.315 78.655 93.485 ;
        RECT 77.230 93.140 77.620 93.315 ;
        RECT 78.105 92.345 78.435 93.145 ;
        RECT 78.825 93.135 79.140 94.155 ;
        RECT 79.345 94.075 80.205 94.325 ;
        RECT 80.375 94.265 80.625 94.515 ;
        RECT 80.795 94.435 80.965 94.895 ;
        RECT 81.135 94.265 81.475 94.725 ;
        RECT 80.375 94.095 81.475 94.265 ;
        RECT 81.735 94.345 81.905 94.725 ;
        RECT 82.120 94.515 82.450 94.895 ;
        RECT 81.735 94.175 82.450 94.345 ;
        RECT 79.345 93.485 79.625 94.075 ;
        RECT 79.795 93.655 80.545 93.905 ;
        RECT 80.715 93.655 81.475 93.905 ;
        RECT 81.645 93.625 82.000 93.995 ;
        RECT 82.280 93.985 82.450 94.175 ;
        RECT 82.620 94.150 82.875 94.725 ;
        RECT 82.280 93.655 82.535 93.985 ;
        RECT 79.345 93.315 81.045 93.485 ;
        RECT 78.605 92.515 79.140 93.135 ;
        RECT 79.450 92.345 79.705 93.145 ;
        RECT 79.875 92.515 80.205 93.315 ;
        RECT 80.375 92.345 80.545 93.145 ;
        RECT 80.715 92.515 81.045 93.315 ;
        RECT 81.215 92.345 81.475 93.485 ;
        RECT 82.280 93.445 82.450 93.655 ;
        RECT 81.735 93.275 82.450 93.445 ;
        RECT 82.705 93.420 82.875 94.150 ;
        RECT 83.050 94.055 83.310 94.895 ;
        RECT 83.945 94.395 84.205 94.725 ;
        RECT 84.375 94.535 84.705 94.895 ;
        RECT 84.960 94.515 86.260 94.725 ;
        RECT 83.945 94.385 84.175 94.395 ;
        RECT 81.735 92.515 81.905 93.275 ;
        RECT 82.120 92.345 82.450 93.105 ;
        RECT 82.620 92.515 82.875 93.420 ;
        RECT 83.050 92.345 83.310 93.495 ;
        RECT 83.945 93.195 84.115 94.385 ;
        RECT 84.960 94.365 85.130 94.515 ;
        RECT 84.375 94.240 85.130 94.365 ;
        RECT 84.285 94.195 85.130 94.240 ;
        RECT 84.285 94.075 84.555 94.195 ;
        RECT 84.285 93.500 84.455 94.075 ;
        RECT 84.685 93.635 85.095 93.940 ;
        RECT 85.385 93.905 85.595 94.305 ;
        RECT 85.265 93.695 85.595 93.905 ;
        RECT 85.840 93.905 86.060 94.305 ;
        RECT 86.535 94.130 86.990 94.895 ;
        RECT 87.165 94.145 88.375 94.895 ;
        RECT 88.545 94.145 89.755 94.895 ;
        RECT 85.840 93.695 86.315 93.905 ;
        RECT 86.505 93.705 86.995 93.905 ;
        RECT 87.165 93.605 87.685 94.145 ;
        RECT 84.285 93.465 84.485 93.500 ;
        RECT 85.815 93.465 86.990 93.525 ;
        RECT 84.285 93.355 86.990 93.465 ;
        RECT 87.855 93.435 88.375 93.975 ;
        RECT 84.345 93.295 86.145 93.355 ;
        RECT 85.815 93.265 86.145 93.295 ;
        RECT 83.945 92.515 84.205 93.195 ;
        RECT 84.375 92.345 84.625 93.125 ;
        RECT 84.875 93.095 85.710 93.105 ;
        RECT 86.300 93.095 86.485 93.185 ;
        RECT 84.875 92.895 86.485 93.095 ;
        RECT 84.875 92.515 85.125 92.895 ;
        RECT 86.255 92.855 86.485 92.895 ;
        RECT 86.735 92.735 86.990 93.355 ;
        RECT 85.295 92.345 85.650 92.725 ;
        RECT 86.655 92.515 86.990 92.735 ;
        RECT 87.165 92.345 88.375 93.435 ;
        RECT 88.545 93.435 89.065 93.975 ;
        RECT 89.235 93.605 89.755 94.145 ;
        RECT 88.545 92.345 89.755 93.435 ;
        RECT 99.980 93.085 100.150 100.195 ;
        RECT 100.550 93.815 100.720 99.855 ;
        RECT 100.990 93.815 101.160 99.855 ;
        RECT 100.690 93.430 101.020 93.600 ;
        RECT 101.560 93.085 101.730 100.195 ;
        RECT 102.130 93.815 102.300 99.855 ;
        RECT 102.570 93.815 102.740 99.855 ;
        RECT 102.270 93.430 102.600 93.600 ;
        RECT 103.140 93.085 103.310 100.195 ;
        RECT 103.710 93.815 103.880 99.855 ;
        RECT 104.150 93.815 104.320 99.855 ;
        RECT 103.850 93.430 104.180 93.600 ;
        RECT 104.720 93.085 104.890 100.195 ;
        RECT 105.290 93.815 105.460 99.855 ;
        RECT 105.730 93.815 105.900 99.855 ;
        RECT 105.430 93.430 105.760 93.600 ;
        RECT 106.300 93.085 106.470 100.195 ;
        RECT 106.870 93.815 107.040 99.855 ;
        RECT 107.310 93.815 107.480 99.855 ;
        RECT 107.010 93.430 107.340 93.600 ;
        RECT 107.880 93.085 108.050 100.195 ;
        RECT 108.450 93.815 108.620 99.855 ;
        RECT 108.890 93.815 109.060 99.855 ;
        RECT 108.590 93.430 108.920 93.600 ;
        RECT 109.460 93.085 109.630 100.195 ;
        RECT 110.030 93.815 110.200 99.855 ;
        RECT 110.470 93.815 110.640 99.855 ;
        RECT 110.170 93.430 110.500 93.600 ;
        RECT 111.040 93.085 111.210 100.195 ;
        RECT 111.610 93.815 111.780 99.855 ;
        RECT 112.050 93.815 112.220 99.855 ;
        RECT 111.750 93.430 112.080 93.600 ;
        RECT 112.620 93.085 112.790 100.195 ;
        RECT 134.450 96.750 134.620 101.720 ;
        RECT 135.100 99.930 135.450 102.090 ;
        RECT 135.100 97.230 135.450 99.390 ;
        RECT 135.930 96.750 136.100 102.570 ;
        RECT 136.580 99.930 136.930 102.090 ;
        RECT 136.580 97.230 136.930 99.390 ;
        RECT 137.410 96.750 137.580 102.570 ;
        RECT 138.060 99.930 138.410 102.090 ;
        RECT 138.060 97.230 138.410 99.390 ;
        RECT 138.890 96.750 139.060 102.570 ;
        RECT 139.540 99.930 139.890 102.090 ;
        RECT 139.540 97.230 139.890 99.390 ;
        RECT 140.370 96.750 140.540 102.570 ;
        RECT 141.020 99.930 141.370 102.090 ;
        RECT 141.020 97.230 141.370 99.390 ;
        RECT 141.850 96.750 142.020 102.570 ;
        RECT 142.500 99.930 142.850 102.090 ;
        RECT 142.500 97.230 142.850 99.390 ;
        RECT 143.330 96.750 143.500 102.570 ;
        RECT 143.980 99.930 144.330 102.090 ;
        RECT 143.980 97.230 144.330 99.390 ;
        RECT 144.810 96.750 144.980 102.570 ;
        RECT 145.460 99.930 145.810 102.090 ;
        RECT 145.460 97.230 145.810 99.390 ;
        RECT 146.290 96.750 146.460 102.570 ;
        RECT 146.940 99.930 147.290 102.090 ;
        RECT 146.940 97.230 147.290 99.390 ;
        RECT 147.770 96.750 147.940 102.570 ;
        RECT 148.420 99.930 148.770 102.090 ;
        RECT 148.420 97.230 148.770 99.390 ;
        RECT 149.250 96.750 149.420 102.570 ;
        RECT 149.900 99.930 150.250 102.090 ;
        RECT 149.900 97.230 150.250 99.390 ;
        RECT 150.730 96.750 150.900 102.570 ;
        RECT 151.380 99.930 151.730 102.090 ;
        RECT 151.380 97.230 151.730 99.390 ;
        RECT 152.210 96.750 152.380 102.570 ;
        RECT 152.860 99.930 153.210 102.090 ;
        RECT 152.860 97.230 153.210 99.390 ;
        RECT 153.690 96.750 153.860 102.570 ;
        RECT 154.340 99.930 154.690 102.090 ;
        RECT 154.340 97.230 154.690 99.390 ;
        RECT 155.170 96.750 155.340 102.570 ;
        RECT 155.820 99.930 156.170 102.090 ;
        RECT 155.820 97.230 156.170 99.390 ;
        RECT 156.650 96.750 156.820 102.570 ;
        RECT 157.300 99.930 157.650 102.090 ;
        RECT 157.300 97.230 157.650 99.390 ;
        RECT 158.130 96.750 158.300 102.570 ;
        RECT 134.450 96.580 158.300 96.750 ;
        RECT 99.980 92.915 112.790 93.085 ;
        RECT 12.100 92.175 89.840 92.345 ;
        RECT 12.185 91.085 13.395 92.175 ;
        RECT 13.655 91.505 13.825 92.005 ;
        RECT 13.995 91.675 14.325 92.175 ;
        RECT 13.655 91.335 14.320 91.505 ;
        RECT 12.185 90.375 12.705 90.915 ;
        RECT 12.875 90.545 13.395 91.085 ;
        RECT 13.570 90.515 13.920 91.165 ;
        RECT 12.185 89.625 13.395 90.375 ;
        RECT 14.090 90.345 14.320 91.335 ;
        RECT 13.655 90.175 14.320 90.345 ;
        RECT 13.655 89.885 13.825 90.175 ;
        RECT 13.995 89.625 14.325 90.005 ;
        RECT 14.495 89.885 14.680 92.005 ;
        RECT 14.920 91.715 15.185 92.175 ;
        RECT 15.355 91.580 15.605 92.005 ;
        RECT 15.815 91.730 16.920 91.900 ;
        RECT 15.300 91.450 15.605 91.580 ;
        RECT 14.850 90.255 15.130 91.205 ;
        RECT 15.300 90.345 15.470 91.450 ;
        RECT 15.640 90.665 15.880 91.260 ;
        RECT 16.050 91.195 16.580 91.560 ;
        RECT 16.050 90.495 16.220 91.195 ;
        RECT 16.750 91.115 16.920 91.730 ;
        RECT 17.090 91.375 17.260 92.175 ;
        RECT 17.430 91.675 17.680 92.005 ;
        RECT 17.905 91.705 18.790 91.875 ;
        RECT 16.750 91.025 17.260 91.115 ;
        RECT 15.300 90.215 15.525 90.345 ;
        RECT 15.695 90.275 16.220 90.495 ;
        RECT 16.390 90.855 17.260 91.025 ;
        RECT 14.935 89.625 15.185 90.085 ;
        RECT 15.355 90.075 15.525 90.215 ;
        RECT 16.390 90.075 16.560 90.855 ;
        RECT 17.090 90.785 17.260 90.855 ;
        RECT 16.770 90.605 16.970 90.635 ;
        RECT 17.430 90.605 17.600 91.675 ;
        RECT 17.770 90.785 17.960 91.505 ;
        RECT 16.770 90.305 17.600 90.605 ;
        RECT 18.130 90.575 18.450 91.535 ;
        RECT 15.355 89.905 15.690 90.075 ;
        RECT 15.885 89.905 16.560 90.075 ;
        RECT 16.880 89.625 17.250 90.125 ;
        RECT 17.430 90.075 17.600 90.305 ;
        RECT 17.985 90.245 18.450 90.575 ;
        RECT 18.620 90.865 18.790 91.705 ;
        RECT 18.970 91.675 19.285 92.175 ;
        RECT 19.515 91.445 19.855 92.005 ;
        RECT 18.960 91.070 19.855 91.445 ;
        RECT 20.025 91.165 20.195 92.175 ;
        RECT 19.665 90.865 19.855 91.070 ;
        RECT 20.365 91.115 20.695 91.960 ;
        RECT 21.850 91.795 22.185 92.175 ;
        RECT 20.365 91.035 20.755 91.115 ;
        RECT 20.540 90.985 20.755 91.035 ;
        RECT 18.620 90.535 19.495 90.865 ;
        RECT 19.665 90.535 20.415 90.865 ;
        RECT 18.620 90.075 18.790 90.535 ;
        RECT 19.665 90.365 19.865 90.535 ;
        RECT 20.585 90.405 20.755 90.985 ;
        RECT 20.530 90.365 20.755 90.405 ;
        RECT 17.430 89.905 17.835 90.075 ;
        RECT 18.005 89.905 18.790 90.075 ;
        RECT 19.065 89.625 19.275 90.155 ;
        RECT 19.535 89.840 19.865 90.365 ;
        RECT 20.375 90.280 20.755 90.365 ;
        RECT 21.845 90.305 22.085 91.615 ;
        RECT 22.355 91.205 22.605 92.005 ;
        RECT 22.825 91.455 23.155 92.175 ;
        RECT 23.340 91.205 23.590 92.005 ;
        RECT 24.055 91.375 24.385 92.175 ;
        RECT 24.555 91.745 24.895 92.005 ;
        RECT 22.255 91.035 24.445 91.205 ;
        RECT 20.035 89.625 20.205 90.235 ;
        RECT 20.375 89.845 20.705 90.280 ;
        RECT 22.255 90.125 22.425 91.035 ;
        RECT 24.130 90.865 24.445 91.035 ;
        RECT 21.930 89.795 22.425 90.125 ;
        RECT 22.645 89.900 22.995 90.865 ;
        RECT 23.175 89.895 23.475 90.865 ;
        RECT 23.655 89.895 23.935 90.865 ;
        RECT 24.130 90.615 24.460 90.865 ;
        RECT 24.115 89.625 24.385 90.425 ;
        RECT 24.635 90.345 24.895 91.745 ;
        RECT 25.065 91.010 25.355 92.175 ;
        RECT 25.530 91.785 25.865 92.005 ;
        RECT 26.870 91.795 27.225 92.175 ;
        RECT 25.530 91.165 25.785 91.785 ;
        RECT 26.035 91.625 26.265 91.665 ;
        RECT 27.395 91.625 27.645 92.005 ;
        RECT 26.035 91.425 27.645 91.625 ;
        RECT 26.035 91.335 26.220 91.425 ;
        RECT 26.810 91.415 27.645 91.425 ;
        RECT 27.895 91.395 28.145 92.175 ;
        RECT 28.315 91.325 28.575 92.005 ;
        RECT 26.375 91.225 26.705 91.255 ;
        RECT 26.375 91.165 28.175 91.225 ;
        RECT 25.530 91.055 28.235 91.165 ;
        RECT 25.530 90.995 26.705 91.055 ;
        RECT 28.035 91.020 28.235 91.055 ;
        RECT 25.525 90.615 26.015 90.815 ;
        RECT 26.205 90.615 26.680 90.825 ;
        RECT 24.555 89.835 24.895 90.345 ;
        RECT 25.065 89.625 25.355 90.350 ;
        RECT 25.530 89.625 25.985 90.390 ;
        RECT 26.460 90.215 26.680 90.615 ;
        RECT 26.925 90.615 27.255 90.825 ;
        RECT 26.925 90.215 27.135 90.615 ;
        RECT 27.425 90.580 27.835 90.885 ;
        RECT 28.065 90.445 28.235 91.020 ;
        RECT 27.965 90.325 28.235 90.445 ;
        RECT 27.390 90.280 28.235 90.325 ;
        RECT 27.390 90.155 28.145 90.280 ;
        RECT 27.390 90.005 27.560 90.155 ;
        RECT 28.405 90.135 28.575 91.325 ;
        RECT 28.800 91.305 29.085 92.175 ;
        RECT 29.255 91.545 29.515 92.005 ;
        RECT 29.690 91.715 29.945 92.175 ;
        RECT 30.115 91.545 30.375 92.005 ;
        RECT 29.255 91.375 30.375 91.545 ;
        RECT 30.545 91.375 30.855 92.175 ;
        RECT 29.255 91.125 29.515 91.375 ;
        RECT 31.025 91.205 31.335 92.005 ;
        RECT 28.760 90.955 29.515 91.125 ;
        RECT 30.305 91.035 31.335 91.205 ;
        RECT 31.505 91.035 31.785 92.175 ;
        RECT 28.760 90.445 29.165 90.955 ;
        RECT 30.305 90.785 30.475 91.035 ;
        RECT 29.335 90.615 30.475 90.785 ;
        RECT 28.760 90.275 30.410 90.445 ;
        RECT 30.645 90.295 30.995 90.865 ;
        RECT 28.345 90.125 28.575 90.135 ;
        RECT 26.260 89.795 27.560 90.005 ;
        RECT 27.815 89.625 28.145 89.985 ;
        RECT 28.315 89.795 28.575 90.125 ;
        RECT 28.805 89.625 29.085 90.105 ;
        RECT 29.255 89.885 29.515 90.275 ;
        RECT 29.690 89.625 29.945 90.105 ;
        RECT 30.115 89.885 30.410 90.275 ;
        RECT 31.165 90.125 31.335 91.035 ;
        RECT 31.955 91.025 32.285 92.005 ;
        RECT 32.455 91.035 32.715 92.175 ;
        RECT 32.975 91.505 33.145 92.005 ;
        RECT 33.315 91.675 33.645 92.175 ;
        RECT 32.975 91.335 33.640 91.505 ;
        RECT 31.515 90.595 31.850 90.865 ;
        RECT 32.020 90.425 32.190 91.025 ;
        RECT 32.360 90.615 32.695 90.865 ;
        RECT 32.890 90.515 33.240 91.165 ;
        RECT 30.590 89.625 30.865 90.105 ;
        RECT 31.035 89.795 31.335 90.125 ;
        RECT 31.505 89.625 31.815 90.425 ;
        RECT 32.020 89.795 32.715 90.425 ;
        RECT 33.410 90.345 33.640 91.335 ;
        RECT 32.975 90.175 33.640 90.345 ;
        RECT 32.975 89.885 33.145 90.175 ;
        RECT 33.315 89.625 33.645 90.005 ;
        RECT 33.815 89.885 34.000 92.005 ;
        RECT 34.240 91.715 34.505 92.175 ;
        RECT 34.675 91.580 34.925 92.005 ;
        RECT 35.135 91.730 36.240 91.900 ;
        RECT 34.620 91.450 34.925 91.580 ;
        RECT 34.170 90.255 34.450 91.205 ;
        RECT 34.620 90.345 34.790 91.450 ;
        RECT 34.960 90.665 35.200 91.260 ;
        RECT 35.370 91.195 35.900 91.560 ;
        RECT 35.370 90.495 35.540 91.195 ;
        RECT 36.070 91.115 36.240 91.730 ;
        RECT 36.410 91.375 36.580 92.175 ;
        RECT 36.750 91.675 37.000 92.005 ;
        RECT 37.225 91.705 38.110 91.875 ;
        RECT 36.070 91.025 36.580 91.115 ;
        RECT 34.620 90.215 34.845 90.345 ;
        RECT 35.015 90.275 35.540 90.495 ;
        RECT 35.710 90.855 36.580 91.025 ;
        RECT 34.255 89.625 34.505 90.085 ;
        RECT 34.675 90.075 34.845 90.215 ;
        RECT 35.710 90.075 35.880 90.855 ;
        RECT 36.410 90.785 36.580 90.855 ;
        RECT 36.090 90.605 36.290 90.635 ;
        RECT 36.750 90.605 36.920 91.675 ;
        RECT 37.090 90.785 37.280 91.505 ;
        RECT 36.090 90.305 36.920 90.605 ;
        RECT 37.450 90.575 37.770 91.535 ;
        RECT 34.675 89.905 35.010 90.075 ;
        RECT 35.205 89.905 35.880 90.075 ;
        RECT 36.200 89.625 36.570 90.125 ;
        RECT 36.750 90.075 36.920 90.305 ;
        RECT 37.305 90.245 37.770 90.575 ;
        RECT 37.940 90.865 38.110 91.705 ;
        RECT 38.290 91.675 38.605 92.175 ;
        RECT 38.835 91.445 39.175 92.005 ;
        RECT 38.280 91.070 39.175 91.445 ;
        RECT 39.345 91.165 39.515 92.175 ;
        RECT 38.985 90.865 39.175 91.070 ;
        RECT 39.685 91.115 40.015 91.960 ;
        RECT 40.305 91.115 40.635 91.960 ;
        RECT 40.805 91.165 40.975 92.175 ;
        RECT 41.145 91.445 41.485 92.005 ;
        RECT 41.715 91.675 42.030 92.175 ;
        RECT 42.210 91.705 43.095 91.875 ;
        RECT 39.685 91.035 40.075 91.115 ;
        RECT 39.860 90.985 40.075 91.035 ;
        RECT 37.940 90.535 38.815 90.865 ;
        RECT 38.985 90.535 39.735 90.865 ;
        RECT 37.940 90.075 38.110 90.535 ;
        RECT 38.985 90.365 39.185 90.535 ;
        RECT 39.905 90.405 40.075 90.985 ;
        RECT 39.850 90.365 40.075 90.405 ;
        RECT 36.750 89.905 37.155 90.075 ;
        RECT 37.325 89.905 38.110 90.075 ;
        RECT 38.385 89.625 38.595 90.155 ;
        RECT 38.855 89.840 39.185 90.365 ;
        RECT 39.695 90.280 40.075 90.365 ;
        RECT 40.245 91.035 40.635 91.115 ;
        RECT 41.145 91.070 42.040 91.445 ;
        RECT 40.245 90.985 40.460 91.035 ;
        RECT 40.245 90.405 40.415 90.985 ;
        RECT 41.145 90.865 41.335 91.070 ;
        RECT 42.210 90.865 42.380 91.705 ;
        RECT 43.320 91.675 43.570 92.005 ;
        RECT 40.585 90.535 41.335 90.865 ;
        RECT 41.505 90.535 42.380 90.865 ;
        RECT 40.245 90.365 40.470 90.405 ;
        RECT 41.135 90.365 41.335 90.535 ;
        RECT 40.245 90.280 40.625 90.365 ;
        RECT 39.355 89.625 39.525 90.235 ;
        RECT 39.695 89.845 40.025 90.280 ;
        RECT 40.295 89.845 40.625 90.280 ;
        RECT 40.795 89.625 40.965 90.235 ;
        RECT 41.135 89.840 41.465 90.365 ;
        RECT 41.725 89.625 41.935 90.155 ;
        RECT 42.210 90.075 42.380 90.535 ;
        RECT 42.550 90.575 42.870 91.535 ;
        RECT 43.040 90.785 43.230 91.505 ;
        RECT 43.400 90.605 43.570 91.675 ;
        RECT 43.740 91.375 43.910 92.175 ;
        RECT 44.080 91.730 45.185 91.900 ;
        RECT 44.080 91.115 44.250 91.730 ;
        RECT 45.395 91.580 45.645 92.005 ;
        RECT 45.815 91.715 46.080 92.175 ;
        RECT 44.420 91.195 44.950 91.560 ;
        RECT 45.395 91.450 45.700 91.580 ;
        RECT 43.740 91.025 44.250 91.115 ;
        RECT 43.740 90.855 44.610 91.025 ;
        RECT 43.740 90.785 43.910 90.855 ;
        RECT 44.030 90.605 44.230 90.635 ;
        RECT 42.550 90.245 43.015 90.575 ;
        RECT 43.400 90.305 44.230 90.605 ;
        RECT 43.400 90.075 43.570 90.305 ;
        RECT 42.210 89.905 42.995 90.075 ;
        RECT 43.165 89.905 43.570 90.075 ;
        RECT 43.750 89.625 44.120 90.125 ;
        RECT 44.440 90.075 44.610 90.855 ;
        RECT 44.780 90.495 44.950 91.195 ;
        RECT 45.120 90.665 45.360 91.260 ;
        RECT 44.780 90.275 45.305 90.495 ;
        RECT 45.530 90.345 45.700 91.450 ;
        RECT 45.475 90.215 45.700 90.345 ;
        RECT 45.870 90.255 46.150 91.205 ;
        RECT 45.475 90.075 45.645 90.215 ;
        RECT 44.440 89.905 45.115 90.075 ;
        RECT 45.310 89.905 45.645 90.075 ;
        RECT 45.815 89.625 46.065 90.085 ;
        RECT 46.320 89.885 46.505 92.005 ;
        RECT 46.675 91.675 47.005 92.175 ;
        RECT 47.175 91.505 47.345 92.005 ;
        RECT 46.680 91.335 47.345 91.505 ;
        RECT 46.680 90.345 46.910 91.335 ;
        RECT 47.080 90.515 47.430 91.165 ;
        RECT 47.605 91.085 50.195 92.175 ;
        RECT 47.605 90.395 48.815 90.915 ;
        RECT 48.985 90.565 50.195 91.085 ;
        RECT 50.825 91.010 51.115 92.175 ;
        RECT 51.285 91.085 52.955 92.175 ;
        RECT 51.285 90.395 52.035 90.915 ;
        RECT 52.205 90.565 52.955 91.085 ;
        RECT 53.125 91.035 53.405 92.175 ;
        RECT 53.575 91.025 53.905 92.005 ;
        RECT 54.075 91.035 54.335 92.175 ;
        RECT 54.505 91.620 55.110 92.175 ;
        RECT 55.285 91.665 55.765 92.005 ;
        RECT 55.935 91.630 56.190 92.175 ;
        RECT 54.505 91.520 55.120 91.620 ;
        RECT 54.935 91.495 55.120 91.520 ;
        RECT 53.135 90.595 53.470 90.865 ;
        RECT 53.640 90.425 53.810 91.025 ;
        RECT 54.505 90.900 54.765 91.350 ;
        RECT 54.935 91.250 55.265 91.495 ;
        RECT 55.435 91.175 56.190 91.425 ;
        RECT 56.360 91.305 56.635 92.005 ;
        RECT 55.420 91.140 56.190 91.175 ;
        RECT 55.405 91.130 56.190 91.140 ;
        RECT 55.400 91.115 56.295 91.130 ;
        RECT 55.380 91.100 56.295 91.115 ;
        RECT 55.360 91.090 56.295 91.100 ;
        RECT 55.335 91.080 56.295 91.090 ;
        RECT 55.265 91.050 56.295 91.080 ;
        RECT 55.245 91.020 56.295 91.050 ;
        RECT 55.225 90.990 56.295 91.020 ;
        RECT 55.195 90.965 56.295 90.990 ;
        RECT 55.160 90.930 56.295 90.965 ;
        RECT 55.130 90.925 56.295 90.930 ;
        RECT 55.130 90.920 55.520 90.925 ;
        RECT 55.130 90.910 55.495 90.920 ;
        RECT 55.130 90.905 55.480 90.910 ;
        RECT 55.130 90.900 55.465 90.905 ;
        RECT 54.505 90.895 55.465 90.900 ;
        RECT 54.505 90.885 55.455 90.895 ;
        RECT 54.505 90.880 55.445 90.885 ;
        RECT 54.505 90.870 55.435 90.880 ;
        RECT 53.980 90.615 54.315 90.865 ;
        RECT 54.505 90.860 55.430 90.870 ;
        RECT 54.505 90.855 55.425 90.860 ;
        RECT 54.505 90.840 55.415 90.855 ;
        RECT 54.505 90.825 55.410 90.840 ;
        RECT 54.505 90.800 55.400 90.825 ;
        RECT 54.505 90.730 55.395 90.800 ;
        RECT 46.680 90.175 47.345 90.345 ;
        RECT 46.675 89.625 47.005 90.005 ;
        RECT 47.175 89.885 47.345 90.175 ;
        RECT 47.605 89.625 50.195 90.395 ;
        RECT 50.825 89.625 51.115 90.350 ;
        RECT 51.285 89.625 52.955 90.395 ;
        RECT 53.125 89.625 53.435 90.425 ;
        RECT 53.640 89.795 54.335 90.425 ;
        RECT 54.505 90.175 55.055 90.560 ;
        RECT 55.225 90.005 55.395 90.730 ;
        RECT 54.505 89.835 55.395 90.005 ;
        RECT 55.565 90.330 55.895 90.755 ;
        RECT 56.065 90.530 56.295 90.925 ;
        RECT 55.565 90.305 55.815 90.330 ;
        RECT 55.565 89.845 55.785 90.305 ;
        RECT 56.465 90.275 56.635 91.305 ;
        RECT 55.955 89.625 56.205 90.165 ;
        RECT 56.375 89.795 56.635 90.275 ;
        RECT 57.270 91.035 57.545 92.005 ;
        RECT 57.755 91.375 58.035 92.175 ;
        RECT 58.205 91.665 59.395 91.955 ;
        RECT 58.205 91.325 59.375 91.495 ;
        RECT 58.205 91.205 58.375 91.325 ;
        RECT 57.715 91.035 58.375 91.205 ;
        RECT 57.270 90.300 57.440 91.035 ;
        RECT 57.715 90.865 57.885 91.035 ;
        RECT 58.685 90.865 58.880 91.155 ;
        RECT 59.050 91.035 59.375 91.325 ;
        RECT 59.570 91.035 59.890 92.175 ;
        RECT 60.070 90.865 60.265 91.915 ;
        RECT 60.445 91.325 60.775 92.005 ;
        RECT 60.975 91.375 61.230 92.175 ;
        RECT 60.445 91.045 60.795 91.325 ;
        RECT 61.590 91.205 61.980 91.380 ;
        RECT 62.465 91.375 62.795 92.175 ;
        RECT 62.965 91.385 63.500 92.005 ;
        RECT 63.705 91.740 69.050 92.175 ;
        RECT 57.610 90.535 57.885 90.865 ;
        RECT 58.055 90.535 58.880 90.865 ;
        RECT 59.050 90.535 59.395 90.865 ;
        RECT 59.630 90.815 59.890 90.865 ;
        RECT 59.625 90.645 59.890 90.815 ;
        RECT 59.630 90.535 59.890 90.645 ;
        RECT 60.070 90.535 60.455 90.865 ;
        RECT 60.625 90.665 60.795 91.045 ;
        RECT 60.985 90.835 61.230 91.195 ;
        RECT 61.590 91.035 63.015 91.205 ;
        RECT 57.715 90.365 57.885 90.535 ;
        RECT 60.625 90.495 61.145 90.665 ;
        RECT 57.270 89.955 57.545 90.300 ;
        RECT 57.715 90.195 59.380 90.365 ;
        RECT 57.735 89.625 58.115 90.025 ;
        RECT 58.285 89.845 58.455 90.195 ;
        RECT 58.625 89.625 58.955 90.025 ;
        RECT 59.125 89.845 59.380 90.195 ;
        RECT 59.570 90.155 60.785 90.325 ;
        RECT 59.570 89.805 59.860 90.155 ;
        RECT 60.055 89.625 60.385 89.985 ;
        RECT 60.555 89.850 60.785 90.155 ;
        RECT 60.975 89.930 61.145 90.495 ;
        RECT 61.465 90.305 61.820 90.865 ;
        RECT 61.990 90.135 62.160 91.035 ;
        RECT 62.330 90.305 62.595 90.865 ;
        RECT 62.845 90.535 63.015 91.035 ;
        RECT 63.185 90.365 63.500 91.385 ;
        RECT 61.570 89.625 61.810 90.135 ;
        RECT 61.990 89.805 62.270 90.135 ;
        RECT 62.500 89.625 62.715 90.135 ;
        RECT 62.885 89.795 63.500 90.365 ;
        RECT 65.290 90.170 65.630 91.000 ;
        RECT 67.110 90.490 67.460 91.740 ;
        RECT 69.225 91.085 70.895 92.175 ;
        RECT 69.225 90.395 69.975 90.915 ;
        RECT 70.145 90.565 70.895 91.085 ;
        RECT 71.585 91.035 71.795 92.175 ;
        RECT 71.965 91.025 72.295 92.005 ;
        RECT 72.465 91.035 72.695 92.175 ;
        RECT 73.110 91.205 73.440 92.005 ;
        RECT 73.610 91.375 73.940 92.175 ;
        RECT 74.240 91.205 74.570 92.005 ;
        RECT 75.215 91.375 75.465 92.175 ;
        RECT 73.110 91.035 75.545 91.205 ;
        RECT 75.735 91.035 75.905 92.175 ;
        RECT 76.075 91.035 76.415 92.005 ;
        RECT 63.705 89.625 69.050 90.170 ;
        RECT 69.225 89.625 70.895 90.395 ;
        RECT 71.585 89.625 71.795 90.445 ;
        RECT 71.965 90.425 72.215 91.025 ;
        RECT 72.385 90.615 72.715 90.865 ;
        RECT 72.905 90.615 73.255 90.865 ;
        RECT 71.965 89.795 72.295 90.425 ;
        RECT 72.465 89.625 72.695 90.445 ;
        RECT 73.440 90.405 73.610 91.035 ;
        RECT 73.780 90.615 74.110 90.815 ;
        RECT 74.280 90.615 74.610 90.815 ;
        RECT 74.780 90.615 75.200 90.815 ;
        RECT 75.375 90.785 75.545 91.035 ;
        RECT 75.375 90.615 76.070 90.785 ;
        RECT 76.240 90.475 76.415 91.035 ;
        RECT 76.585 91.010 76.875 92.175 ;
        RECT 77.135 91.505 77.305 92.005 ;
        RECT 77.475 91.675 77.805 92.175 ;
        RECT 77.135 91.335 77.800 91.505 ;
        RECT 77.050 90.515 77.400 91.165 ;
        RECT 73.110 89.795 73.610 90.405 ;
        RECT 74.240 90.275 75.465 90.445 ;
        RECT 76.185 90.425 76.415 90.475 ;
        RECT 74.240 89.795 74.570 90.275 ;
        RECT 74.740 89.625 74.965 90.085 ;
        RECT 75.135 89.795 75.465 90.275 ;
        RECT 75.655 89.625 75.905 90.425 ;
        RECT 76.075 89.795 76.415 90.425 ;
        RECT 76.585 89.625 76.875 90.350 ;
        RECT 77.570 90.345 77.800 91.335 ;
        RECT 77.135 90.175 77.800 90.345 ;
        RECT 77.135 89.885 77.305 90.175 ;
        RECT 77.475 89.625 77.805 90.005 ;
        RECT 77.975 89.885 78.160 92.005 ;
        RECT 78.400 91.715 78.665 92.175 ;
        RECT 78.835 91.580 79.085 92.005 ;
        RECT 79.295 91.730 80.400 91.900 ;
        RECT 78.780 91.450 79.085 91.580 ;
        RECT 78.330 90.255 78.610 91.205 ;
        RECT 78.780 90.345 78.950 91.450 ;
        RECT 79.120 90.665 79.360 91.260 ;
        RECT 79.530 91.195 80.060 91.560 ;
        RECT 79.530 90.495 79.700 91.195 ;
        RECT 80.230 91.115 80.400 91.730 ;
        RECT 80.570 91.375 80.740 92.175 ;
        RECT 80.910 91.675 81.160 92.005 ;
        RECT 81.385 91.705 82.270 91.875 ;
        RECT 80.230 91.025 80.740 91.115 ;
        RECT 78.780 90.215 79.005 90.345 ;
        RECT 79.175 90.275 79.700 90.495 ;
        RECT 79.870 90.855 80.740 91.025 ;
        RECT 78.415 89.625 78.665 90.085 ;
        RECT 78.835 90.075 79.005 90.215 ;
        RECT 79.870 90.075 80.040 90.855 ;
        RECT 80.570 90.785 80.740 90.855 ;
        RECT 80.250 90.605 80.450 90.635 ;
        RECT 80.910 90.605 81.080 91.675 ;
        RECT 81.250 90.785 81.440 91.505 ;
        RECT 80.250 90.305 81.080 90.605 ;
        RECT 81.610 90.575 81.930 91.535 ;
        RECT 78.835 89.905 79.170 90.075 ;
        RECT 79.365 89.905 80.040 90.075 ;
        RECT 80.360 89.625 80.730 90.125 ;
        RECT 80.910 90.075 81.080 90.305 ;
        RECT 81.465 90.245 81.930 90.575 ;
        RECT 82.100 90.865 82.270 91.705 ;
        RECT 82.450 91.675 82.765 92.175 ;
        RECT 82.995 91.445 83.335 92.005 ;
        RECT 82.440 91.070 83.335 91.445 ;
        RECT 83.505 91.165 83.675 92.175 ;
        RECT 83.145 90.865 83.335 91.070 ;
        RECT 83.845 91.115 84.175 91.960 ;
        RECT 83.845 91.035 84.235 91.115 ;
        RECT 84.020 90.985 84.235 91.035 ;
        RECT 82.100 90.535 82.975 90.865 ;
        RECT 83.145 90.535 83.895 90.865 ;
        RECT 82.100 90.075 82.270 90.535 ;
        RECT 83.145 90.365 83.345 90.535 ;
        RECT 84.065 90.405 84.235 90.985 ;
        RECT 84.010 90.365 84.235 90.405 ;
        RECT 80.910 89.905 81.315 90.075 ;
        RECT 81.485 89.905 82.270 90.075 ;
        RECT 82.545 89.625 82.755 90.155 ;
        RECT 83.015 89.840 83.345 90.365 ;
        RECT 83.855 90.280 84.235 90.365 ;
        RECT 84.405 91.035 84.745 92.005 ;
        RECT 84.915 91.035 85.085 92.175 ;
        RECT 85.355 91.375 85.605 92.175 ;
        RECT 86.250 91.205 86.580 92.005 ;
        RECT 86.880 91.375 87.210 92.175 ;
        RECT 87.380 91.205 87.710 92.005 ;
        RECT 85.275 91.035 87.710 91.205 ;
        RECT 88.545 91.085 89.755 92.175 ;
        RECT 99.990 91.675 112.800 91.845 ;
        RECT 84.405 90.425 84.580 91.035 ;
        RECT 85.275 90.785 85.445 91.035 ;
        RECT 84.750 90.615 85.445 90.785 ;
        RECT 85.620 90.615 86.040 90.815 ;
        RECT 86.210 90.615 86.540 90.815 ;
        RECT 86.710 90.615 87.040 90.815 ;
        RECT 83.515 89.625 83.685 90.235 ;
        RECT 83.855 89.845 84.185 90.280 ;
        RECT 84.405 89.795 84.745 90.425 ;
        RECT 84.915 89.625 85.165 90.425 ;
        RECT 85.355 90.275 86.580 90.445 ;
        RECT 85.355 89.795 85.685 90.275 ;
        RECT 85.855 89.625 86.080 90.085 ;
        RECT 86.250 89.795 86.580 90.275 ;
        RECT 87.210 90.405 87.380 91.035 ;
        RECT 87.565 90.615 87.915 90.865 ;
        RECT 88.545 90.545 89.065 91.085 ;
        RECT 87.210 89.795 87.710 90.405 ;
        RECT 89.235 90.375 89.755 90.915 ;
        RECT 88.545 89.625 89.755 90.375 ;
        RECT 12.100 89.455 89.840 89.625 ;
        RECT 12.185 88.705 13.395 89.455 ;
        RECT 13.655 88.905 13.825 89.195 ;
        RECT 13.995 89.075 14.325 89.455 ;
        RECT 13.655 88.735 14.320 88.905 ;
        RECT 12.185 88.165 12.705 88.705 ;
        RECT 12.875 87.995 13.395 88.535 ;
        RECT 12.185 86.905 13.395 87.995 ;
        RECT 13.570 87.915 13.920 88.565 ;
        RECT 14.090 87.745 14.320 88.735 ;
        RECT 13.655 87.575 14.320 87.745 ;
        RECT 13.655 87.075 13.825 87.575 ;
        RECT 13.995 86.905 14.325 87.405 ;
        RECT 14.495 87.075 14.680 89.195 ;
        RECT 14.935 88.995 15.185 89.455 ;
        RECT 15.355 89.005 15.690 89.175 ;
        RECT 15.885 89.005 16.560 89.175 ;
        RECT 15.355 88.865 15.525 89.005 ;
        RECT 14.850 87.875 15.130 88.825 ;
        RECT 15.300 88.735 15.525 88.865 ;
        RECT 15.300 87.630 15.470 88.735 ;
        RECT 15.695 88.585 16.220 88.805 ;
        RECT 15.640 87.820 15.880 88.415 ;
        RECT 16.050 87.885 16.220 88.585 ;
        RECT 16.390 88.225 16.560 89.005 ;
        RECT 16.880 88.955 17.250 89.455 ;
        RECT 17.430 89.005 17.835 89.175 ;
        RECT 18.005 89.005 18.790 89.175 ;
        RECT 17.430 88.775 17.600 89.005 ;
        RECT 16.770 88.475 17.600 88.775 ;
        RECT 17.985 88.505 18.450 88.835 ;
        RECT 16.770 88.445 16.970 88.475 ;
        RECT 17.090 88.225 17.260 88.295 ;
        RECT 16.390 88.055 17.260 88.225 ;
        RECT 16.750 87.965 17.260 88.055 ;
        RECT 15.300 87.500 15.605 87.630 ;
        RECT 16.050 87.520 16.580 87.885 ;
        RECT 14.920 86.905 15.185 87.365 ;
        RECT 15.355 87.075 15.605 87.500 ;
        RECT 16.750 87.350 16.920 87.965 ;
        RECT 15.815 87.180 16.920 87.350 ;
        RECT 17.090 86.905 17.260 87.705 ;
        RECT 17.430 87.405 17.600 88.475 ;
        RECT 17.770 87.575 17.960 88.295 ;
        RECT 18.130 87.545 18.450 88.505 ;
        RECT 18.620 88.545 18.790 89.005 ;
        RECT 19.065 88.925 19.275 89.455 ;
        RECT 19.535 88.715 19.865 89.240 ;
        RECT 20.035 88.845 20.205 89.455 ;
        RECT 20.375 88.800 20.705 89.235 ;
        RECT 20.375 88.715 20.755 88.800 ;
        RECT 19.665 88.545 19.865 88.715 ;
        RECT 20.530 88.675 20.755 88.715 ;
        RECT 18.620 88.215 19.495 88.545 ;
        RECT 19.665 88.215 20.415 88.545 ;
        RECT 17.430 87.075 17.680 87.405 ;
        RECT 18.620 87.375 18.790 88.215 ;
        RECT 19.665 88.010 19.855 88.215 ;
        RECT 20.585 88.095 20.755 88.675 ;
        RECT 20.540 88.045 20.755 88.095 ;
        RECT 18.960 87.635 19.855 88.010 ;
        RECT 20.365 87.965 20.755 88.045 ;
        RECT 20.925 88.735 21.265 89.245 ;
        RECT 17.905 87.205 18.790 87.375 ;
        RECT 18.970 86.905 19.285 87.405 ;
        RECT 19.515 87.075 19.855 87.635 ;
        RECT 20.025 86.905 20.195 87.915 ;
        RECT 20.365 87.120 20.695 87.965 ;
        RECT 20.925 87.335 21.185 88.735 ;
        RECT 21.435 88.655 21.705 89.455 ;
        RECT 21.360 88.215 21.690 88.465 ;
        RECT 21.885 88.215 22.165 89.185 ;
        RECT 22.345 88.215 22.645 89.185 ;
        RECT 22.825 88.215 23.175 89.180 ;
        RECT 23.395 88.955 23.890 89.285 ;
        RECT 21.375 88.045 21.690 88.215 ;
        RECT 23.395 88.045 23.565 88.955 ;
        RECT 21.375 87.875 23.565 88.045 ;
        RECT 20.925 87.075 21.265 87.335 ;
        RECT 21.435 86.905 21.765 87.705 ;
        RECT 22.230 87.075 22.480 87.875 ;
        RECT 22.665 86.905 22.995 87.625 ;
        RECT 23.215 87.075 23.465 87.875 ;
        RECT 23.735 87.465 23.975 88.775 ;
        RECT 24.180 88.715 24.795 89.285 ;
        RECT 24.965 88.945 25.180 89.455 ;
        RECT 25.410 88.945 25.690 89.275 ;
        RECT 25.870 88.945 26.110 89.455 ;
        RECT 26.490 88.995 27.240 89.285 ;
        RECT 27.750 88.995 28.080 89.455 ;
        RECT 24.180 87.695 24.495 88.715 ;
        RECT 24.665 88.045 24.835 88.545 ;
        RECT 25.085 88.215 25.350 88.775 ;
        RECT 25.520 88.045 25.690 88.945 ;
        RECT 25.860 88.215 26.215 88.775 ;
        RECT 24.665 87.875 26.090 88.045 ;
        RECT 23.635 86.905 23.970 87.285 ;
        RECT 24.180 87.075 24.715 87.695 ;
        RECT 24.885 86.905 25.215 87.705 ;
        RECT 25.700 87.700 26.090 87.875 ;
        RECT 26.490 87.705 26.860 88.995 ;
        RECT 28.300 88.805 28.570 89.015 ;
        RECT 27.235 88.635 28.570 88.805 ;
        RECT 28.745 88.995 29.305 89.285 ;
        RECT 29.475 88.995 29.725 89.455 ;
        RECT 27.235 88.465 27.405 88.635 ;
        RECT 27.030 88.215 27.405 88.465 ;
        RECT 27.575 88.225 28.050 88.465 ;
        RECT 28.220 88.225 28.570 88.465 ;
        RECT 27.235 88.045 27.405 88.215 ;
        RECT 27.235 87.875 28.570 88.045 ;
        RECT 28.290 87.715 28.570 87.875 ;
        RECT 26.490 87.535 27.660 87.705 ;
        RECT 26.945 86.905 27.160 87.365 ;
        RECT 27.330 87.075 27.660 87.535 ;
        RECT 27.830 86.905 28.080 87.705 ;
        RECT 28.745 87.625 28.995 88.995 ;
        RECT 30.345 88.825 30.675 89.185 ;
        RECT 31.505 89.075 32.395 89.245 ;
        RECT 29.285 88.635 30.675 88.825 ;
        RECT 29.285 88.545 29.455 88.635 ;
        RECT 29.165 88.215 29.455 88.545 ;
        RECT 31.505 88.520 32.055 88.905 ;
        RECT 29.625 88.215 29.965 88.465 ;
        RECT 30.185 88.215 30.860 88.465 ;
        RECT 32.225 88.350 32.395 89.075 ;
        RECT 29.285 87.965 29.455 88.215 ;
        RECT 29.285 87.795 30.225 87.965 ;
        RECT 30.595 87.855 30.860 88.215 ;
        RECT 31.505 88.280 32.395 88.350 ;
        RECT 32.565 88.750 32.785 89.235 ;
        RECT 32.955 88.915 33.205 89.455 ;
        RECT 33.375 88.805 33.635 89.285 ;
        RECT 32.565 88.325 32.895 88.750 ;
        RECT 31.505 88.255 32.400 88.280 ;
        RECT 31.505 88.240 32.410 88.255 ;
        RECT 31.505 88.225 32.415 88.240 ;
        RECT 31.505 88.220 32.425 88.225 ;
        RECT 31.505 88.210 32.430 88.220 ;
        RECT 31.505 88.200 32.435 88.210 ;
        RECT 31.505 88.195 32.445 88.200 ;
        RECT 31.505 88.185 32.455 88.195 ;
        RECT 31.505 88.180 32.465 88.185 ;
        RECT 28.745 87.075 29.205 87.625 ;
        RECT 29.395 86.905 29.725 87.625 ;
        RECT 29.925 87.245 30.225 87.795 ;
        RECT 31.505 87.730 31.765 88.180 ;
        RECT 32.130 88.175 32.465 88.180 ;
        RECT 32.130 88.170 32.480 88.175 ;
        RECT 32.130 88.160 32.495 88.170 ;
        RECT 32.130 88.155 32.520 88.160 ;
        RECT 33.065 88.155 33.295 88.550 ;
        RECT 32.130 88.150 33.295 88.155 ;
        RECT 32.160 88.115 33.295 88.150 ;
        RECT 32.195 88.090 33.295 88.115 ;
        RECT 32.225 88.060 33.295 88.090 ;
        RECT 32.245 88.030 33.295 88.060 ;
        RECT 32.265 88.000 33.295 88.030 ;
        RECT 32.335 87.990 33.295 88.000 ;
        RECT 32.360 87.980 33.295 87.990 ;
        RECT 32.380 87.965 33.295 87.980 ;
        RECT 32.400 87.950 33.295 87.965 ;
        RECT 32.405 87.940 33.190 87.950 ;
        RECT 32.420 87.905 33.190 87.940 ;
        RECT 31.935 87.585 32.265 87.830 ;
        RECT 32.435 87.655 33.190 87.905 ;
        RECT 33.465 87.775 33.635 88.805 ;
        RECT 33.805 88.635 34.065 89.455 ;
        RECT 34.235 88.635 34.565 89.055 ;
        RECT 34.745 88.970 35.535 89.235 ;
        RECT 34.315 88.545 34.565 88.635 ;
        RECT 30.395 86.905 30.675 87.575 ;
        RECT 31.935 87.560 32.120 87.585 ;
        RECT 31.505 87.460 32.120 87.560 ;
        RECT 31.505 86.905 32.110 87.460 ;
        RECT 32.285 87.075 32.765 87.415 ;
        RECT 32.935 86.905 33.190 87.450 ;
        RECT 33.360 87.075 33.635 87.775 ;
        RECT 33.805 87.585 34.145 88.465 ;
        RECT 34.315 88.295 35.110 88.545 ;
        RECT 33.805 86.905 34.065 87.415 ;
        RECT 34.315 87.075 34.485 88.295 ;
        RECT 35.280 88.115 35.535 88.970 ;
        RECT 35.705 88.815 35.905 89.235 ;
        RECT 36.095 88.995 36.425 89.455 ;
        RECT 35.705 88.295 36.115 88.815 ;
        RECT 36.595 88.805 36.855 89.285 ;
        RECT 36.285 88.115 36.515 88.545 ;
        RECT 34.725 87.945 36.515 88.115 ;
        RECT 34.725 87.580 34.975 87.945 ;
        RECT 35.145 87.585 35.475 87.775 ;
        RECT 35.695 87.650 36.410 87.945 ;
        RECT 36.685 87.775 36.855 88.805 ;
        RECT 37.945 88.730 38.235 89.455 ;
        RECT 38.405 88.705 39.615 89.455 ;
        RECT 38.405 88.165 38.925 88.705 ;
        RECT 39.785 88.635 40.045 89.455 ;
        RECT 40.215 88.635 40.545 89.055 ;
        RECT 40.725 88.970 41.515 89.235 ;
        RECT 40.295 88.545 40.545 88.635 ;
        RECT 35.145 87.410 35.340 87.585 ;
        RECT 34.725 86.905 35.340 87.410 ;
        RECT 35.510 87.075 35.985 87.415 ;
        RECT 36.155 86.905 36.370 87.450 ;
        RECT 36.580 87.075 36.855 87.775 ;
        RECT 37.945 86.905 38.235 88.070 ;
        RECT 39.095 87.995 39.615 88.535 ;
        RECT 38.405 86.905 39.615 87.995 ;
        RECT 39.785 87.585 40.125 88.465 ;
        RECT 40.295 88.295 41.090 88.545 ;
        RECT 39.785 86.905 40.045 87.415 ;
        RECT 40.295 87.075 40.465 88.295 ;
        RECT 41.260 88.115 41.515 88.970 ;
        RECT 41.685 88.815 41.885 89.235 ;
        RECT 42.075 88.995 42.405 89.455 ;
        RECT 41.685 88.295 42.095 88.815 ;
        RECT 42.575 88.805 42.835 89.285 ;
        RECT 43.170 88.945 43.410 89.455 ;
        RECT 43.590 88.945 43.870 89.275 ;
        RECT 44.100 88.945 44.315 89.455 ;
        RECT 42.265 88.115 42.495 88.545 ;
        RECT 40.705 87.945 42.495 88.115 ;
        RECT 40.705 87.580 40.955 87.945 ;
        RECT 41.125 87.585 41.455 87.775 ;
        RECT 41.675 87.650 42.390 87.945 ;
        RECT 42.665 87.775 42.835 88.805 ;
        RECT 43.065 88.215 43.420 88.775 ;
        RECT 43.590 88.045 43.760 88.945 ;
        RECT 43.930 88.215 44.195 88.775 ;
        RECT 44.485 88.715 45.100 89.285 ;
        RECT 44.445 88.045 44.615 88.545 ;
        RECT 41.125 87.410 41.320 87.585 ;
        RECT 40.705 86.905 41.320 87.410 ;
        RECT 41.490 87.075 41.965 87.415 ;
        RECT 42.135 86.905 42.350 87.450 ;
        RECT 42.560 87.075 42.835 87.775 ;
        RECT 43.190 87.875 44.615 88.045 ;
        RECT 43.190 87.700 43.580 87.875 ;
        RECT 44.065 86.905 44.395 87.705 ;
        RECT 44.785 87.695 45.100 88.715 ;
        RECT 45.305 88.685 48.815 89.455 ;
        RECT 48.985 88.705 50.195 89.455 ;
        RECT 45.305 88.165 46.955 88.685 ;
        RECT 47.125 87.995 48.815 88.515 ;
        RECT 48.985 88.165 49.505 88.705 ;
        RECT 50.375 88.645 50.645 89.455 ;
        RECT 50.815 88.645 51.145 89.285 ;
        RECT 51.315 88.645 51.555 89.455 ;
        RECT 49.675 87.995 50.195 88.535 ;
        RECT 50.365 88.215 50.715 88.465 ;
        RECT 50.885 88.045 51.055 88.645 ;
        RECT 51.750 88.615 52.010 89.455 ;
        RECT 52.185 88.710 52.440 89.285 ;
        RECT 52.610 89.075 52.940 89.455 ;
        RECT 53.155 88.905 53.325 89.285 ;
        RECT 52.610 88.735 53.325 88.905 ;
        RECT 51.225 88.215 51.575 88.465 ;
        RECT 44.565 87.075 45.100 87.695 ;
        RECT 45.305 86.905 48.815 87.995 ;
        RECT 48.985 86.905 50.195 87.995 ;
        RECT 50.375 86.905 50.705 88.045 ;
        RECT 50.885 87.875 51.565 88.045 ;
        RECT 51.235 87.090 51.565 87.875 ;
        RECT 51.750 86.905 52.010 88.055 ;
        RECT 52.185 87.980 52.355 88.710 ;
        RECT 52.610 88.545 52.780 88.735 ;
        RECT 53.585 88.715 54.025 89.275 ;
        RECT 54.195 88.715 54.645 89.455 ;
        RECT 54.815 88.885 54.985 89.285 ;
        RECT 55.155 89.055 55.575 89.455 ;
        RECT 55.745 88.885 55.975 89.285 ;
        RECT 54.815 88.715 55.975 88.885 ;
        RECT 56.145 88.715 56.635 89.285 ;
        RECT 52.525 88.215 52.780 88.545 ;
        RECT 52.610 88.005 52.780 88.215 ;
        RECT 53.060 88.185 53.415 88.555 ;
        RECT 52.185 87.075 52.440 87.980 ;
        RECT 52.610 87.835 53.325 88.005 ;
        RECT 52.610 86.905 52.940 87.665 ;
        RECT 53.155 87.075 53.325 87.835 ;
        RECT 53.585 87.705 53.895 88.715 ;
        RECT 54.065 88.095 54.235 88.545 ;
        RECT 54.405 88.265 54.795 88.545 ;
        RECT 54.980 88.215 55.225 88.545 ;
        RECT 54.065 87.925 54.855 88.095 ;
        RECT 53.585 87.075 54.025 87.705 ;
        RECT 54.200 86.905 54.515 87.755 ;
        RECT 54.685 87.245 54.855 87.925 ;
        RECT 55.025 87.415 55.225 88.215 ;
        RECT 55.425 87.415 55.675 88.545 ;
        RECT 55.890 88.215 56.295 88.545 ;
        RECT 56.465 88.045 56.635 88.715 ;
        RECT 55.865 87.875 56.635 88.045 ;
        RECT 56.810 88.780 57.085 89.125 ;
        RECT 57.275 89.055 57.655 89.455 ;
        RECT 57.825 88.885 57.995 89.235 ;
        RECT 58.165 89.055 58.495 89.455 ;
        RECT 58.665 88.885 58.920 89.235 ;
        RECT 56.810 88.045 56.980 88.780 ;
        RECT 57.255 88.715 58.920 88.885 ;
        RECT 59.120 88.885 59.375 89.235 ;
        RECT 59.545 89.055 59.875 89.455 ;
        RECT 60.045 88.885 60.215 89.235 ;
        RECT 60.385 89.055 60.765 89.455 ;
        RECT 59.120 88.715 60.785 88.885 ;
        RECT 60.955 88.780 61.230 89.125 ;
        RECT 61.405 89.075 62.295 89.245 ;
        RECT 57.255 88.545 57.425 88.715 ;
        RECT 60.615 88.545 60.785 88.715 ;
        RECT 57.150 88.215 57.425 88.545 ;
        RECT 57.595 88.215 58.420 88.545 ;
        RECT 58.590 88.215 58.935 88.545 ;
        RECT 59.105 88.215 59.450 88.545 ;
        RECT 59.620 88.215 60.445 88.545 ;
        RECT 60.615 88.215 60.890 88.545 ;
        RECT 57.255 88.045 57.425 88.215 ;
        RECT 55.865 87.245 56.115 87.875 ;
        RECT 54.685 87.075 56.115 87.245 ;
        RECT 56.295 86.905 56.625 87.705 ;
        RECT 56.810 87.075 57.085 88.045 ;
        RECT 57.255 87.875 57.915 88.045 ;
        RECT 58.225 87.925 58.420 88.215 ;
        RECT 57.745 87.755 57.915 87.875 ;
        RECT 58.590 87.755 58.915 88.045 ;
        RECT 57.295 86.905 57.575 87.705 ;
        RECT 57.745 87.585 58.915 87.755 ;
        RECT 59.125 87.755 59.450 88.045 ;
        RECT 59.620 87.925 59.815 88.215 ;
        RECT 60.615 88.045 60.785 88.215 ;
        RECT 61.060 88.045 61.230 88.780 ;
        RECT 61.405 88.520 61.955 88.905 ;
        RECT 62.125 88.350 62.295 89.075 ;
        RECT 60.125 87.875 60.785 88.045 ;
        RECT 60.125 87.755 60.295 87.875 ;
        RECT 59.125 87.585 60.295 87.755 ;
        RECT 57.745 87.125 58.935 87.415 ;
        RECT 59.105 87.125 60.295 87.415 ;
        RECT 60.465 86.905 60.745 87.705 ;
        RECT 60.955 87.075 61.230 88.045 ;
        RECT 61.405 88.280 62.295 88.350 ;
        RECT 62.465 88.750 62.685 89.235 ;
        RECT 62.855 88.915 63.105 89.455 ;
        RECT 63.275 88.805 63.535 89.285 ;
        RECT 62.465 88.325 62.795 88.750 ;
        RECT 61.405 88.255 62.300 88.280 ;
        RECT 61.405 88.240 62.310 88.255 ;
        RECT 61.405 88.225 62.315 88.240 ;
        RECT 61.405 88.220 62.325 88.225 ;
        RECT 61.405 88.210 62.330 88.220 ;
        RECT 61.405 88.200 62.335 88.210 ;
        RECT 61.405 88.195 62.345 88.200 ;
        RECT 61.405 88.185 62.355 88.195 ;
        RECT 61.405 88.180 62.365 88.185 ;
        RECT 61.405 87.730 61.665 88.180 ;
        RECT 62.030 88.175 62.365 88.180 ;
        RECT 62.030 88.170 62.380 88.175 ;
        RECT 62.030 88.160 62.395 88.170 ;
        RECT 62.030 88.155 62.420 88.160 ;
        RECT 62.965 88.155 63.195 88.550 ;
        RECT 62.030 88.150 63.195 88.155 ;
        RECT 62.060 88.115 63.195 88.150 ;
        RECT 62.095 88.090 63.195 88.115 ;
        RECT 62.125 88.060 63.195 88.090 ;
        RECT 62.145 88.030 63.195 88.060 ;
        RECT 62.165 88.000 63.195 88.030 ;
        RECT 62.235 87.990 63.195 88.000 ;
        RECT 62.260 87.980 63.195 87.990 ;
        RECT 62.280 87.965 63.195 87.980 ;
        RECT 62.300 87.950 63.195 87.965 ;
        RECT 62.305 87.940 63.090 87.950 ;
        RECT 62.320 87.905 63.090 87.940 ;
        RECT 61.835 87.585 62.165 87.830 ;
        RECT 62.335 87.655 63.090 87.905 ;
        RECT 63.365 87.775 63.535 88.805 ;
        RECT 63.705 88.730 63.995 89.455 ;
        RECT 64.165 88.805 64.425 89.285 ;
        RECT 64.595 88.915 64.845 89.455 ;
        RECT 61.835 87.560 62.020 87.585 ;
        RECT 61.405 87.460 62.020 87.560 ;
        RECT 61.405 86.905 62.010 87.460 ;
        RECT 62.185 87.075 62.665 87.415 ;
        RECT 62.835 86.905 63.090 87.450 ;
        RECT 63.260 87.075 63.535 87.775 ;
        RECT 63.705 86.905 63.995 88.070 ;
        RECT 64.165 87.775 64.335 88.805 ;
        RECT 65.015 88.775 65.235 89.235 ;
        RECT 64.985 88.750 65.235 88.775 ;
        RECT 64.505 88.155 64.735 88.550 ;
        RECT 64.905 88.325 65.235 88.750 ;
        RECT 65.405 89.075 66.295 89.245 ;
        RECT 65.405 88.350 65.575 89.075 ;
        RECT 65.745 88.520 66.295 88.905 ;
        RECT 66.465 88.705 67.675 89.455 ;
        RECT 65.405 88.280 66.295 88.350 ;
        RECT 65.400 88.255 66.295 88.280 ;
        RECT 65.390 88.240 66.295 88.255 ;
        RECT 65.385 88.225 66.295 88.240 ;
        RECT 65.375 88.220 66.295 88.225 ;
        RECT 65.370 88.210 66.295 88.220 ;
        RECT 65.365 88.200 66.295 88.210 ;
        RECT 65.355 88.195 66.295 88.200 ;
        RECT 65.345 88.185 66.295 88.195 ;
        RECT 65.335 88.180 66.295 88.185 ;
        RECT 65.335 88.175 65.670 88.180 ;
        RECT 65.320 88.170 65.670 88.175 ;
        RECT 65.305 88.160 65.670 88.170 ;
        RECT 65.280 88.155 65.670 88.160 ;
        RECT 64.505 88.150 65.670 88.155 ;
        RECT 64.505 88.115 65.640 88.150 ;
        RECT 64.505 88.090 65.605 88.115 ;
        RECT 64.505 88.060 65.575 88.090 ;
        RECT 64.505 88.030 65.555 88.060 ;
        RECT 64.505 88.000 65.535 88.030 ;
        RECT 64.505 87.990 65.465 88.000 ;
        RECT 64.505 87.980 65.440 87.990 ;
        RECT 64.505 87.965 65.420 87.980 ;
        RECT 64.505 87.950 65.400 87.965 ;
        RECT 64.610 87.940 65.395 87.950 ;
        RECT 64.610 87.905 65.380 87.940 ;
        RECT 64.165 87.075 64.440 87.775 ;
        RECT 64.610 87.655 65.365 87.905 ;
        RECT 65.535 87.585 65.865 87.830 ;
        RECT 66.035 87.730 66.295 88.180 ;
        RECT 66.465 88.165 66.985 88.705 ;
        RECT 67.885 88.635 68.115 89.455 ;
        RECT 68.285 88.655 68.615 89.285 ;
        RECT 67.155 87.995 67.675 88.535 ;
        RECT 67.865 88.215 68.195 88.465 ;
        RECT 68.365 88.055 68.615 88.655 ;
        RECT 68.785 88.635 68.995 89.455 ;
        RECT 69.230 88.615 69.490 89.455 ;
        RECT 69.665 88.710 69.920 89.285 ;
        RECT 70.090 89.075 70.420 89.455 ;
        RECT 70.635 88.905 70.805 89.285 ;
        RECT 71.085 88.945 71.325 89.455 ;
        RECT 71.495 88.945 71.785 89.285 ;
        RECT 72.015 88.945 72.330 89.455 ;
        RECT 70.090 88.735 70.805 88.905 ;
        RECT 65.680 87.560 65.865 87.585 ;
        RECT 65.680 87.460 66.295 87.560 ;
        RECT 64.610 86.905 64.865 87.450 ;
        RECT 65.035 87.075 65.515 87.415 ;
        RECT 65.690 86.905 66.295 87.460 ;
        RECT 66.465 86.905 67.675 87.995 ;
        RECT 67.885 86.905 68.115 88.045 ;
        RECT 68.285 87.075 68.615 88.055 ;
        RECT 68.785 86.905 68.995 88.045 ;
        RECT 69.230 86.905 69.490 88.055 ;
        RECT 69.665 87.980 69.835 88.710 ;
        RECT 70.090 88.545 70.260 88.735 ;
        RECT 70.005 88.215 70.260 88.545 ;
        RECT 70.090 88.005 70.260 88.215 ;
        RECT 70.540 88.185 70.895 88.555 ;
        RECT 71.130 88.435 71.325 88.775 ;
        RECT 71.125 88.265 71.325 88.435 ;
        RECT 71.130 88.215 71.325 88.265 ;
        RECT 71.495 88.045 71.675 88.945 ;
        RECT 72.500 88.885 72.670 89.155 ;
        RECT 72.840 89.055 73.170 89.455 ;
        RECT 71.845 88.215 72.255 88.775 ;
        RECT 72.500 88.715 73.195 88.885 ;
        RECT 72.425 88.045 72.595 88.545 ;
        RECT 69.665 87.075 69.920 87.980 ;
        RECT 70.090 87.835 70.805 88.005 ;
        RECT 70.090 86.905 70.420 87.665 ;
        RECT 70.635 87.075 70.805 87.835 ;
        RECT 71.135 87.875 72.595 88.045 ;
        RECT 71.135 87.700 71.495 87.875 ;
        RECT 72.765 87.705 73.195 88.715 ;
        RECT 73.370 88.635 73.645 89.455 ;
        RECT 73.815 88.815 74.145 89.285 ;
        RECT 74.315 88.985 74.485 89.455 ;
        RECT 74.655 88.815 74.985 89.285 ;
        RECT 75.155 88.985 75.445 89.455 ;
        RECT 73.815 88.805 74.985 88.815 ;
        RECT 73.815 88.635 75.415 88.805 ;
        RECT 73.370 88.265 74.090 88.465 ;
        RECT 74.260 88.265 75.030 88.465 ;
        RECT 75.200 88.095 75.415 88.635 ;
        RECT 72.080 86.905 72.250 87.705 ;
        RECT 72.420 87.535 73.195 87.705 ;
        RECT 73.370 87.875 74.485 88.085 ;
        RECT 72.420 87.075 72.750 87.535 ;
        RECT 72.920 86.905 73.090 87.365 ;
        RECT 73.370 87.075 73.645 87.875 ;
        RECT 73.815 86.905 74.145 87.705 ;
        RECT 74.315 87.245 74.485 87.875 ;
        RECT 74.655 87.875 75.415 88.095 ;
        RECT 76.620 88.715 77.235 89.285 ;
        RECT 77.405 88.945 77.620 89.455 ;
        RECT 77.850 88.945 78.130 89.275 ;
        RECT 78.310 88.945 78.550 89.455 ;
        RECT 78.885 88.995 79.445 89.285 ;
        RECT 79.615 88.995 79.865 89.455 ;
        RECT 74.655 87.415 74.985 87.875 ;
        RECT 75.155 87.245 75.455 87.705 ;
        RECT 74.315 87.075 75.455 87.245 ;
        RECT 76.620 87.695 76.935 88.715 ;
        RECT 77.105 88.045 77.275 88.545 ;
        RECT 77.525 88.215 77.790 88.775 ;
        RECT 77.960 88.045 78.130 88.945 ;
        RECT 78.300 88.215 78.655 88.775 ;
        RECT 77.105 87.875 78.530 88.045 ;
        RECT 76.620 87.075 77.155 87.695 ;
        RECT 77.325 86.905 77.655 87.705 ;
        RECT 78.140 87.700 78.530 87.875 ;
        RECT 78.885 87.625 79.135 88.995 ;
        RECT 80.485 88.825 80.815 89.185 ;
        RECT 79.425 88.635 80.815 88.825 ;
        RECT 81.275 88.905 81.445 89.195 ;
        RECT 81.615 89.075 81.945 89.455 ;
        RECT 81.275 88.735 81.940 88.905 ;
        RECT 79.425 88.545 79.595 88.635 ;
        RECT 79.305 88.215 79.595 88.545 ;
        RECT 79.765 88.215 80.105 88.465 ;
        RECT 80.325 88.215 81.000 88.465 ;
        RECT 79.425 87.965 79.595 88.215 ;
        RECT 79.425 87.795 80.365 87.965 ;
        RECT 80.735 87.855 81.000 88.215 ;
        RECT 81.190 87.915 81.540 88.565 ;
        RECT 78.885 87.075 79.345 87.625 ;
        RECT 79.535 86.905 79.865 87.625 ;
        RECT 80.065 87.245 80.365 87.795 ;
        RECT 81.710 87.745 81.940 88.735 ;
        RECT 81.275 87.575 81.940 87.745 ;
        RECT 80.535 86.905 80.815 87.575 ;
        RECT 81.275 87.075 81.445 87.575 ;
        RECT 81.615 86.905 81.945 87.405 ;
        RECT 82.115 87.075 82.300 89.195 ;
        RECT 82.555 88.995 82.805 89.455 ;
        RECT 82.975 89.005 83.310 89.175 ;
        RECT 83.505 89.005 84.180 89.175 ;
        RECT 82.975 88.865 83.145 89.005 ;
        RECT 82.470 87.875 82.750 88.825 ;
        RECT 82.920 88.735 83.145 88.865 ;
        RECT 82.920 87.630 83.090 88.735 ;
        RECT 83.315 88.585 83.840 88.805 ;
        RECT 83.260 87.820 83.500 88.415 ;
        RECT 83.670 87.885 83.840 88.585 ;
        RECT 84.010 88.225 84.180 89.005 ;
        RECT 84.500 88.955 84.870 89.455 ;
        RECT 85.050 89.005 85.455 89.175 ;
        RECT 85.625 89.005 86.410 89.175 ;
        RECT 85.050 88.775 85.220 89.005 ;
        RECT 84.390 88.475 85.220 88.775 ;
        RECT 85.605 88.505 86.070 88.835 ;
        RECT 84.390 88.445 84.590 88.475 ;
        RECT 84.710 88.225 84.880 88.295 ;
        RECT 84.010 88.055 84.880 88.225 ;
        RECT 84.370 87.965 84.880 88.055 ;
        RECT 82.920 87.500 83.225 87.630 ;
        RECT 83.670 87.520 84.200 87.885 ;
        RECT 82.540 86.905 82.805 87.365 ;
        RECT 82.975 87.075 83.225 87.500 ;
        RECT 84.370 87.350 84.540 87.965 ;
        RECT 83.435 87.180 84.540 87.350 ;
        RECT 84.710 86.905 84.880 87.705 ;
        RECT 85.050 87.405 85.220 88.475 ;
        RECT 85.390 87.575 85.580 88.295 ;
        RECT 85.750 87.545 86.070 88.505 ;
        RECT 86.240 88.545 86.410 89.005 ;
        RECT 86.685 88.925 86.895 89.455 ;
        RECT 87.155 88.715 87.485 89.240 ;
        RECT 87.655 88.845 87.825 89.455 ;
        RECT 87.995 88.800 88.325 89.235 ;
        RECT 87.995 88.715 88.375 88.800 ;
        RECT 87.285 88.545 87.485 88.715 ;
        RECT 88.150 88.675 88.375 88.715 ;
        RECT 88.545 88.705 89.755 89.455 ;
        RECT 86.240 88.215 87.115 88.545 ;
        RECT 87.285 88.215 88.035 88.545 ;
        RECT 85.050 87.075 85.300 87.405 ;
        RECT 86.240 87.375 86.410 88.215 ;
        RECT 87.285 88.010 87.475 88.215 ;
        RECT 88.205 88.095 88.375 88.675 ;
        RECT 88.160 88.045 88.375 88.095 ;
        RECT 86.580 87.635 87.475 88.010 ;
        RECT 87.985 87.965 88.375 88.045 ;
        RECT 88.545 87.995 89.065 88.535 ;
        RECT 89.235 88.165 89.755 88.705 ;
        RECT 99.990 88.605 100.160 91.675 ;
        RECT 100.700 91.165 101.030 91.335 ;
        RECT 100.560 88.955 100.730 90.995 ;
        RECT 101.000 88.955 101.170 90.995 ;
        RECT 101.570 88.605 101.740 91.675 ;
        RECT 102.280 91.165 102.610 91.335 ;
        RECT 102.140 88.955 102.310 90.995 ;
        RECT 102.580 88.955 102.750 90.995 ;
        RECT 103.150 88.605 103.320 91.675 ;
        RECT 103.860 91.165 104.190 91.335 ;
        RECT 103.720 88.955 103.890 90.995 ;
        RECT 104.160 88.955 104.330 90.995 ;
        RECT 104.730 88.605 104.900 91.675 ;
        RECT 105.440 91.165 105.770 91.335 ;
        RECT 105.300 88.955 105.470 90.995 ;
        RECT 105.740 88.955 105.910 90.995 ;
        RECT 106.310 88.605 106.480 91.675 ;
        RECT 107.020 91.165 107.350 91.335 ;
        RECT 106.880 88.955 107.050 90.995 ;
        RECT 107.320 88.955 107.490 90.995 ;
        RECT 107.890 88.605 108.060 91.675 ;
        RECT 108.600 91.165 108.930 91.335 ;
        RECT 108.460 88.955 108.630 90.995 ;
        RECT 108.900 88.955 109.070 90.995 ;
        RECT 109.470 88.605 109.640 91.675 ;
        RECT 110.180 91.165 110.510 91.335 ;
        RECT 110.040 88.955 110.210 90.995 ;
        RECT 110.480 88.955 110.650 90.995 ;
        RECT 111.050 88.605 111.220 91.675 ;
        RECT 111.760 91.165 112.090 91.335 ;
        RECT 111.620 88.955 111.790 90.995 ;
        RECT 112.060 88.955 112.230 90.995 ;
        RECT 112.630 88.605 112.800 91.675 ;
        RECT 99.990 88.415 112.800 88.605 ;
        RECT 85.525 87.205 86.410 87.375 ;
        RECT 86.590 86.905 86.905 87.405 ;
        RECT 87.135 87.075 87.475 87.635 ;
        RECT 87.645 86.905 87.815 87.915 ;
        RECT 87.985 87.120 88.315 87.965 ;
        RECT 88.545 86.905 89.755 87.995 ;
        RECT 100.070 87.785 112.760 88.415 ;
        RECT 99.990 87.615 113.480 87.785 ;
        RECT 12.100 86.735 89.840 86.905 ;
        RECT 12.185 85.645 13.395 86.735 ;
        RECT 12.185 84.935 12.705 85.475 ;
        RECT 12.875 85.105 13.395 85.645 ;
        RECT 14.485 85.865 14.760 86.565 ;
        RECT 14.970 86.190 15.185 86.735 ;
        RECT 15.355 86.225 15.830 86.565 ;
        RECT 16.000 86.230 16.615 86.735 ;
        RECT 16.000 86.055 16.195 86.230 ;
        RECT 12.185 84.185 13.395 84.935 ;
        RECT 14.485 84.835 14.655 85.865 ;
        RECT 14.930 85.695 15.645 85.990 ;
        RECT 15.865 85.865 16.195 86.055 ;
        RECT 16.365 85.695 16.615 86.060 ;
        RECT 14.825 85.525 16.615 85.695 ;
        RECT 14.825 85.095 15.055 85.525 ;
        RECT 14.485 84.355 14.745 84.835 ;
        RECT 15.225 84.825 15.635 85.345 ;
        RECT 14.915 84.185 15.245 84.645 ;
        RECT 15.435 84.405 15.635 84.825 ;
        RECT 15.805 84.670 16.060 85.525 ;
        RECT 16.855 85.345 17.025 86.565 ;
        RECT 17.275 86.225 17.535 86.735 ;
        RECT 16.230 85.095 17.025 85.345 ;
        RECT 17.195 85.175 17.535 86.055 ;
        RECT 18.625 85.595 18.885 86.735 ;
        RECT 19.125 86.225 20.740 86.555 ;
        RECT 19.135 85.425 19.305 85.985 ;
        RECT 19.565 85.885 20.740 86.055 ;
        RECT 20.910 85.935 21.190 86.735 ;
        RECT 19.565 85.595 19.895 85.885 ;
        RECT 20.570 85.765 20.740 85.885 ;
        RECT 20.065 85.425 20.310 85.715 ;
        RECT 20.570 85.595 21.230 85.765 ;
        RECT 21.400 85.595 21.675 86.565 ;
        RECT 21.845 86.225 22.105 86.735 ;
        RECT 21.060 85.425 21.230 85.595 ;
        RECT 18.630 85.175 18.965 85.425 ;
        RECT 16.775 85.005 17.025 85.095 ;
        RECT 19.135 85.095 19.850 85.425 ;
        RECT 20.065 85.095 20.890 85.425 ;
        RECT 21.060 85.095 21.335 85.425 ;
        RECT 19.135 85.005 19.385 85.095 ;
        RECT 15.805 84.405 16.595 84.670 ;
        RECT 16.775 84.585 17.105 85.005 ;
        RECT 17.275 84.185 17.535 85.005 ;
        RECT 18.625 84.185 18.885 85.005 ;
        RECT 19.055 84.585 19.385 85.005 ;
        RECT 21.060 84.925 21.230 85.095 ;
        RECT 19.565 84.755 21.230 84.925 ;
        RECT 21.505 84.860 21.675 85.595 ;
        RECT 21.845 85.175 22.185 86.055 ;
        RECT 22.355 85.345 22.525 86.565 ;
        RECT 22.765 86.230 23.380 86.735 ;
        RECT 22.765 85.695 23.015 86.060 ;
        RECT 23.185 86.055 23.380 86.230 ;
        RECT 23.550 86.225 24.025 86.565 ;
        RECT 24.195 86.190 24.410 86.735 ;
        RECT 23.185 85.865 23.515 86.055 ;
        RECT 23.735 85.695 24.450 85.990 ;
        RECT 24.620 85.865 24.895 86.565 ;
        RECT 22.765 85.525 24.555 85.695 ;
        RECT 22.355 85.095 23.150 85.345 ;
        RECT 22.355 85.005 22.605 85.095 ;
        RECT 19.565 84.355 19.825 84.755 ;
        RECT 19.995 84.185 20.325 84.585 ;
        RECT 20.495 84.405 20.665 84.755 ;
        RECT 20.835 84.185 21.210 84.585 ;
        RECT 21.400 84.515 21.675 84.860 ;
        RECT 21.845 84.185 22.105 85.005 ;
        RECT 22.275 84.585 22.605 85.005 ;
        RECT 23.320 84.670 23.575 85.525 ;
        RECT 22.785 84.405 23.575 84.670 ;
        RECT 23.745 84.825 24.155 85.345 ;
        RECT 24.325 85.095 24.555 85.525 ;
        RECT 24.725 84.835 24.895 85.865 ;
        RECT 25.065 85.570 25.355 86.735 ;
        RECT 25.730 85.765 26.060 86.565 ;
        RECT 26.230 85.935 26.560 86.735 ;
        RECT 26.860 85.765 27.190 86.565 ;
        RECT 27.835 85.935 28.085 86.735 ;
        RECT 25.730 85.595 28.165 85.765 ;
        RECT 28.355 85.595 28.525 86.735 ;
        RECT 28.695 85.595 29.035 86.565 ;
        RECT 29.255 86.275 29.465 86.735 ;
        RECT 29.955 86.145 30.455 86.565 ;
        RECT 25.525 85.175 25.875 85.425 ;
        RECT 26.060 84.965 26.230 85.595 ;
        RECT 26.400 85.175 26.730 85.375 ;
        RECT 26.900 85.175 27.230 85.375 ;
        RECT 27.400 85.175 27.820 85.375 ;
        RECT 27.995 85.345 28.165 85.595 ;
        RECT 27.995 85.175 28.690 85.345 ;
        RECT 23.745 84.405 23.945 84.825 ;
        RECT 24.135 84.185 24.465 84.645 ;
        RECT 24.635 84.355 24.895 84.835 ;
        RECT 25.065 84.185 25.355 84.910 ;
        RECT 25.730 84.355 26.230 84.965 ;
        RECT 26.860 84.835 28.085 85.005 ;
        RECT 28.860 84.985 29.035 85.595 ;
        RECT 26.860 84.355 27.190 84.835 ;
        RECT 27.360 84.185 27.585 84.645 ;
        RECT 27.755 84.355 28.085 84.835 ;
        RECT 28.275 84.185 28.525 84.985 ;
        RECT 28.695 84.355 29.035 84.985 ;
        RECT 29.205 84.765 29.445 86.090 ;
        RECT 29.615 85.935 30.455 86.145 ;
        RECT 29.615 84.925 29.785 85.935 ;
        RECT 29.955 85.515 30.355 85.765 ;
        RECT 30.645 85.715 30.845 86.505 ;
        RECT 30.525 85.545 30.845 85.715 ;
        RECT 31.015 85.555 31.335 86.735 ;
        RECT 31.505 85.595 31.785 86.735 ;
        RECT 31.955 85.585 32.285 86.565 ;
        RECT 32.455 85.595 32.715 86.735 ;
        RECT 33.840 85.945 34.375 86.565 ;
        RECT 29.955 85.095 30.125 85.515 ;
        RECT 30.525 85.345 30.705 85.545 ;
        RECT 30.340 85.175 30.705 85.345 ;
        RECT 30.875 85.175 31.335 85.375 ;
        RECT 31.515 85.155 31.850 85.425 ;
        RECT 32.020 84.985 32.190 85.585 ;
        RECT 32.360 85.175 32.695 85.425 ;
        RECT 30.305 84.925 31.335 84.965 ;
        RECT 29.615 84.745 29.965 84.925 ;
        RECT 30.135 84.795 31.335 84.925 ;
        RECT 30.135 84.575 30.465 84.795 ;
        RECT 29.205 84.395 30.465 84.575 ;
        RECT 30.655 84.185 30.825 84.625 ;
        RECT 30.995 84.380 31.335 84.795 ;
        RECT 31.505 84.185 31.815 84.985 ;
        RECT 32.020 84.355 32.715 84.985 ;
        RECT 33.840 84.925 34.155 85.945 ;
        RECT 34.545 85.935 34.875 86.735 ;
        RECT 35.360 85.765 35.750 85.940 ;
        RECT 34.325 85.595 35.750 85.765 ;
        RECT 36.195 85.725 36.365 86.565 ;
        RECT 36.535 86.395 37.705 86.565 ;
        RECT 36.535 85.895 36.865 86.395 ;
        RECT 37.375 86.355 37.705 86.395 ;
        RECT 37.895 86.315 38.250 86.735 ;
        RECT 37.035 86.135 37.265 86.225 ;
        RECT 38.420 86.135 38.670 86.565 ;
        RECT 37.035 85.895 38.670 86.135 ;
        RECT 38.840 85.975 39.170 86.735 ;
        RECT 39.340 85.895 39.595 86.565 ;
        RECT 34.325 85.095 34.495 85.595 ;
        RECT 33.840 84.355 34.455 84.925 ;
        RECT 34.745 84.865 35.010 85.425 ;
        RECT 35.180 84.695 35.350 85.595 ;
        RECT 36.195 85.555 39.255 85.725 ;
        RECT 35.520 84.865 35.875 85.425 ;
        RECT 36.110 85.175 36.460 85.385 ;
        RECT 36.630 85.175 37.075 85.375 ;
        RECT 37.245 85.175 37.720 85.375 ;
        RECT 36.195 84.835 37.260 85.005 ;
        RECT 34.625 84.185 34.840 84.695 ;
        RECT 35.070 84.365 35.350 84.695 ;
        RECT 35.530 84.185 35.770 84.695 ;
        RECT 36.195 84.355 36.365 84.835 ;
        RECT 36.535 84.185 36.865 84.665 ;
        RECT 37.090 84.605 37.260 84.835 ;
        RECT 37.440 84.775 37.720 85.175 ;
        RECT 37.990 85.175 38.320 85.375 ;
        RECT 38.490 85.175 38.855 85.375 ;
        RECT 37.990 84.775 38.275 85.175 ;
        RECT 39.085 85.005 39.255 85.555 ;
        RECT 38.455 84.835 39.255 85.005 ;
        RECT 38.455 84.605 38.625 84.835 ;
        RECT 39.425 84.765 39.595 85.895 ;
        RECT 39.845 85.675 40.175 86.520 ;
        RECT 40.345 85.725 40.515 86.735 ;
        RECT 40.685 86.005 41.025 86.565 ;
        RECT 41.255 86.235 41.570 86.735 ;
        RECT 41.750 86.265 42.635 86.435 ;
        RECT 39.785 85.595 40.175 85.675 ;
        RECT 40.685 85.630 41.580 86.005 ;
        RECT 39.785 85.545 40.000 85.595 ;
        RECT 39.785 84.965 39.955 85.545 ;
        RECT 40.685 85.425 40.875 85.630 ;
        RECT 41.750 85.425 41.920 86.265 ;
        RECT 42.860 86.235 43.110 86.565 ;
        RECT 40.125 85.095 40.875 85.425 ;
        RECT 41.045 85.095 41.920 85.425 ;
        RECT 39.785 84.925 40.010 84.965 ;
        RECT 40.675 84.925 40.875 85.095 ;
        RECT 39.785 84.840 40.165 84.925 ;
        RECT 39.410 84.695 39.595 84.765 ;
        RECT 39.385 84.685 39.595 84.695 ;
        RECT 37.090 84.355 38.625 84.605 ;
        RECT 38.795 84.185 39.125 84.665 ;
        RECT 39.340 84.355 39.595 84.685 ;
        RECT 39.835 84.405 40.165 84.840 ;
        RECT 40.335 84.185 40.505 84.795 ;
        RECT 40.675 84.400 41.005 84.925 ;
        RECT 41.265 84.185 41.475 84.715 ;
        RECT 41.750 84.635 41.920 85.095 ;
        RECT 42.090 85.135 42.410 86.095 ;
        RECT 42.580 85.345 42.770 86.065 ;
        RECT 42.940 85.165 43.110 86.235 ;
        RECT 43.280 85.935 43.450 86.735 ;
        RECT 43.620 86.290 44.725 86.460 ;
        RECT 43.620 85.675 43.790 86.290 ;
        RECT 44.935 86.140 45.185 86.565 ;
        RECT 45.355 86.275 45.620 86.735 ;
        RECT 43.960 85.755 44.490 86.120 ;
        RECT 44.935 86.010 45.240 86.140 ;
        RECT 43.280 85.585 43.790 85.675 ;
        RECT 43.280 85.415 44.150 85.585 ;
        RECT 43.280 85.345 43.450 85.415 ;
        RECT 43.570 85.165 43.770 85.195 ;
        RECT 42.090 84.805 42.555 85.135 ;
        RECT 42.940 84.865 43.770 85.165 ;
        RECT 42.940 84.635 43.110 84.865 ;
        RECT 41.750 84.465 42.535 84.635 ;
        RECT 42.705 84.465 43.110 84.635 ;
        RECT 43.290 84.185 43.660 84.685 ;
        RECT 43.980 84.635 44.150 85.415 ;
        RECT 44.320 85.055 44.490 85.755 ;
        RECT 44.660 85.225 44.900 85.820 ;
        RECT 44.320 84.835 44.845 85.055 ;
        RECT 45.070 84.905 45.240 86.010 ;
        RECT 45.015 84.775 45.240 84.905 ;
        RECT 45.410 84.815 45.690 85.765 ;
        RECT 45.015 84.635 45.185 84.775 ;
        RECT 43.980 84.465 44.655 84.635 ;
        RECT 44.850 84.465 45.185 84.635 ;
        RECT 45.355 84.185 45.605 84.645 ;
        RECT 45.860 84.445 46.045 86.565 ;
        RECT 46.215 86.235 46.545 86.735 ;
        RECT 46.715 86.065 46.885 86.565 ;
        RECT 46.220 85.895 46.885 86.065 ;
        RECT 46.220 84.905 46.450 85.895 ;
        RECT 47.145 85.865 47.420 86.565 ;
        RECT 47.630 86.190 47.845 86.735 ;
        RECT 48.015 86.225 48.490 86.565 ;
        RECT 48.660 86.230 49.275 86.735 ;
        RECT 48.660 86.055 48.855 86.230 ;
        RECT 46.620 85.075 46.970 85.725 ;
        RECT 46.220 84.735 46.885 84.905 ;
        RECT 46.215 84.185 46.545 84.565 ;
        RECT 46.715 84.445 46.885 84.735 ;
        RECT 47.145 84.835 47.315 85.865 ;
        RECT 47.590 85.695 48.305 85.990 ;
        RECT 48.525 85.865 48.855 86.055 ;
        RECT 49.025 85.695 49.275 86.060 ;
        RECT 47.485 85.525 49.275 85.695 ;
        RECT 47.485 85.095 47.715 85.525 ;
        RECT 47.145 84.355 47.405 84.835 ;
        RECT 47.885 84.825 48.295 85.345 ;
        RECT 47.575 84.185 47.905 84.645 ;
        RECT 48.095 84.405 48.295 84.825 ;
        RECT 48.465 84.670 48.720 85.525 ;
        RECT 49.515 85.345 49.685 86.565 ;
        RECT 49.935 86.225 50.195 86.735 ;
        RECT 48.890 85.095 49.685 85.345 ;
        RECT 49.855 85.175 50.195 86.055 ;
        RECT 50.825 85.570 51.115 86.735 ;
        RECT 51.290 85.595 51.610 86.735 ;
        RECT 51.790 85.425 51.985 86.475 ;
        RECT 52.165 85.885 52.495 86.565 ;
        RECT 52.695 85.935 52.950 86.735 ;
        RECT 52.165 85.605 52.515 85.885 ;
        RECT 51.350 85.375 51.610 85.425 ;
        RECT 51.345 85.205 51.610 85.375 ;
        RECT 51.350 85.095 51.610 85.205 ;
        RECT 51.790 85.095 52.175 85.425 ;
        RECT 52.345 85.225 52.515 85.605 ;
        RECT 52.705 85.395 52.950 85.755 ;
        RECT 49.435 85.005 49.685 85.095 ;
        RECT 52.345 85.055 52.865 85.225 ;
        RECT 48.465 84.405 49.255 84.670 ;
        RECT 49.435 84.585 49.765 85.005 ;
        RECT 49.935 84.185 50.195 85.005 ;
        RECT 50.825 84.185 51.115 84.910 ;
        RECT 51.290 84.715 52.505 84.885 ;
        RECT 51.290 84.365 51.580 84.715 ;
        RECT 51.775 84.185 52.105 84.545 ;
        RECT 52.275 84.410 52.505 84.715 ;
        RECT 52.695 84.490 52.865 85.055 ;
        RECT 53.125 84.465 53.405 86.565 ;
        RECT 53.595 85.975 54.380 86.735 ;
        RECT 54.775 85.905 55.160 86.565 ;
        RECT 54.775 85.805 55.185 85.905 ;
        RECT 53.575 85.595 55.185 85.805 ;
        RECT 55.485 85.715 55.685 86.505 ;
        RECT 53.575 84.995 53.850 85.595 ;
        RECT 55.355 85.545 55.685 85.715 ;
        RECT 55.855 85.555 56.175 86.735 ;
        RECT 56.385 85.595 56.615 86.735 ;
        RECT 56.785 85.585 57.115 86.565 ;
        RECT 57.285 85.595 57.495 86.735 ;
        RECT 57.930 85.765 58.260 86.565 ;
        RECT 58.430 85.935 58.760 86.735 ;
        RECT 59.060 85.765 59.390 86.565 ;
        RECT 60.035 85.935 60.285 86.735 ;
        RECT 57.930 85.595 60.365 85.765 ;
        RECT 60.555 85.595 60.725 86.735 ;
        RECT 60.895 85.595 61.235 86.565 ;
        RECT 55.355 85.425 55.535 85.545 ;
        RECT 54.020 85.175 54.375 85.425 ;
        RECT 54.570 85.175 55.035 85.425 ;
        RECT 55.205 85.175 55.535 85.425 ;
        RECT 55.710 85.175 56.175 85.375 ;
        RECT 56.365 85.175 56.695 85.425 ;
        RECT 53.575 84.815 54.825 84.995 ;
        RECT 54.460 84.745 54.825 84.815 ;
        RECT 54.995 84.795 56.175 84.965 ;
        RECT 53.635 84.185 53.805 84.645 ;
        RECT 54.995 84.575 55.325 84.795 ;
        RECT 54.075 84.395 55.325 84.575 ;
        RECT 55.495 84.185 55.665 84.625 ;
        RECT 55.835 84.380 56.175 84.795 ;
        RECT 56.385 84.185 56.615 85.005 ;
        RECT 56.865 84.985 57.115 85.585 ;
        RECT 57.725 85.175 58.075 85.425 ;
        RECT 56.785 84.355 57.115 84.985 ;
        RECT 57.285 84.185 57.495 85.005 ;
        RECT 58.260 84.965 58.430 85.595 ;
        RECT 58.600 85.175 58.930 85.375 ;
        RECT 59.100 85.175 59.430 85.375 ;
        RECT 59.600 85.175 60.020 85.375 ;
        RECT 60.195 85.345 60.365 85.595 ;
        RECT 60.195 85.175 60.890 85.345 ;
        RECT 57.930 84.355 58.430 84.965 ;
        RECT 59.060 84.835 60.285 85.005 ;
        RECT 61.060 84.985 61.235 85.595 ;
        RECT 62.480 85.725 62.780 86.565 ;
        RECT 62.975 85.895 63.225 86.735 ;
        RECT 63.815 86.145 64.620 86.565 ;
        RECT 63.395 85.975 64.960 86.145 ;
        RECT 63.395 85.725 63.565 85.975 ;
        RECT 62.480 85.555 63.565 85.725 ;
        RECT 62.325 85.095 62.655 85.385 ;
        RECT 59.060 84.355 59.390 84.835 ;
        RECT 59.560 84.185 59.785 84.645 ;
        RECT 59.955 84.355 60.285 84.835 ;
        RECT 60.475 84.185 60.725 84.985 ;
        RECT 60.895 84.355 61.235 84.985 ;
        RECT 62.825 84.925 62.995 85.555 ;
        RECT 63.735 85.425 64.055 85.805 ;
        RECT 64.245 85.715 64.620 85.805 ;
        RECT 64.225 85.545 64.620 85.715 ;
        RECT 64.790 85.725 64.960 85.975 ;
        RECT 65.130 85.895 65.460 86.735 ;
        RECT 65.630 85.975 66.295 86.565 ;
        RECT 64.790 85.555 65.710 85.725 ;
        RECT 63.165 85.175 63.495 85.385 ;
        RECT 63.675 85.175 64.055 85.425 ;
        RECT 64.245 85.385 64.620 85.545 ;
        RECT 65.540 85.385 65.710 85.555 ;
        RECT 64.245 85.175 64.730 85.385 ;
        RECT 64.920 85.175 65.370 85.385 ;
        RECT 65.540 85.175 65.875 85.385 ;
        RECT 66.045 85.005 66.295 85.975 ;
        RECT 66.470 86.345 66.805 86.565 ;
        RECT 67.810 86.355 68.165 86.735 ;
        RECT 66.470 85.725 66.725 86.345 ;
        RECT 66.975 86.185 67.205 86.225 ;
        RECT 68.335 86.185 68.585 86.565 ;
        RECT 66.975 85.985 68.585 86.185 ;
        RECT 66.975 85.895 67.160 85.985 ;
        RECT 67.750 85.975 68.585 85.985 ;
        RECT 68.835 85.955 69.085 86.735 ;
        RECT 69.255 85.885 69.515 86.565 ;
        RECT 67.315 85.785 67.645 85.815 ;
        RECT 67.315 85.725 69.115 85.785 ;
        RECT 66.470 85.615 69.175 85.725 ;
        RECT 66.470 85.555 67.645 85.615 ;
        RECT 68.975 85.580 69.175 85.615 ;
        RECT 66.465 85.175 66.955 85.375 ;
        RECT 67.145 85.175 67.620 85.385 ;
        RECT 62.485 84.745 62.995 84.925 ;
        RECT 63.400 84.835 65.100 85.005 ;
        RECT 63.400 84.745 63.785 84.835 ;
        RECT 62.485 84.355 62.815 84.745 ;
        RECT 62.985 84.405 64.170 84.575 ;
        RECT 64.430 84.185 64.600 84.655 ;
        RECT 64.770 84.370 65.100 84.835 ;
        RECT 65.270 84.185 65.440 85.005 ;
        RECT 65.610 84.365 66.295 85.005 ;
        RECT 66.470 84.185 66.925 84.950 ;
        RECT 67.400 84.775 67.620 85.175 ;
        RECT 67.865 85.175 68.195 85.385 ;
        RECT 67.865 84.775 68.075 85.175 ;
        RECT 68.365 85.140 68.775 85.445 ;
        RECT 69.005 85.005 69.175 85.580 ;
        RECT 68.905 84.885 69.175 85.005 ;
        RECT 68.330 84.840 69.175 84.885 ;
        RECT 68.330 84.715 69.085 84.840 ;
        RECT 68.330 84.565 68.500 84.715 ;
        RECT 69.345 84.695 69.515 85.885 ;
        RECT 69.870 85.765 70.260 85.940 ;
        RECT 70.745 85.935 71.075 86.735 ;
        RECT 71.245 85.945 71.780 86.565 ;
        RECT 72.905 86.230 73.535 86.735 ;
        RECT 69.870 85.595 71.295 85.765 ;
        RECT 69.745 84.865 70.100 85.425 ;
        RECT 70.270 84.695 70.440 85.595 ;
        RECT 70.610 84.865 70.875 85.425 ;
        RECT 71.125 85.095 71.295 85.595 ;
        RECT 71.465 84.925 71.780 85.945 ;
        RECT 72.920 85.695 73.175 86.060 ;
        RECT 73.345 86.055 73.535 86.230 ;
        RECT 73.715 86.225 74.190 86.565 ;
        RECT 73.345 85.865 73.675 86.055 ;
        RECT 73.900 85.695 74.150 85.990 ;
        RECT 74.375 85.890 74.590 86.735 ;
        RECT 74.790 85.895 75.065 86.565 ;
        RECT 72.920 85.525 74.710 85.695 ;
        RECT 74.895 85.545 75.065 85.895 ;
        RECT 75.235 85.725 75.495 86.735 ;
        RECT 76.585 85.570 76.875 86.735 ;
        RECT 77.045 86.230 77.675 86.735 ;
        RECT 77.060 85.695 77.315 86.060 ;
        RECT 77.485 86.055 77.675 86.230 ;
        RECT 77.855 86.225 78.330 86.565 ;
        RECT 77.485 85.865 77.815 86.055 ;
        RECT 78.040 85.695 78.290 85.990 ;
        RECT 78.515 85.890 78.730 86.735 ;
        RECT 78.930 85.895 79.205 86.565 ;
        RECT 69.285 84.685 69.515 84.695 ;
        RECT 67.200 84.355 68.500 84.565 ;
        RECT 68.755 84.185 69.085 84.545 ;
        RECT 69.255 84.355 69.515 84.685 ;
        RECT 69.850 84.185 70.090 84.695 ;
        RECT 70.270 84.365 70.550 84.695 ;
        RECT 70.780 84.185 70.995 84.695 ;
        RECT 71.165 84.355 71.780 84.925 ;
        RECT 72.905 84.865 73.290 85.345 ;
        RECT 73.460 84.670 73.715 85.525 ;
        RECT 72.925 84.405 73.715 84.670 ;
        RECT 73.885 84.850 74.295 85.345 ;
        RECT 74.480 85.095 74.710 85.525 ;
        RECT 74.880 85.025 75.495 85.545 ;
        RECT 77.060 85.525 78.850 85.695 ;
        RECT 79.035 85.545 79.205 85.895 ;
        RECT 79.375 85.725 79.635 86.735 ;
        RECT 79.805 85.595 80.065 86.735 ;
        RECT 80.235 85.765 80.565 86.565 ;
        RECT 80.735 85.935 80.905 86.735 ;
        RECT 81.075 85.765 81.405 86.565 ;
        RECT 81.575 85.935 81.830 86.735 ;
        RECT 82.110 85.785 82.375 86.555 ;
        RECT 82.545 86.015 82.875 86.735 ;
        RECT 83.065 86.195 83.325 86.555 ;
        RECT 83.495 86.365 83.825 86.735 ;
        RECT 83.995 86.195 84.255 86.555 ;
        RECT 83.065 85.965 84.255 86.195 ;
        RECT 84.825 85.785 85.115 86.555 ;
        RECT 80.235 85.595 81.935 85.765 ;
        RECT 73.885 84.405 74.115 84.850 ;
        RECT 74.880 84.815 75.050 85.025 ;
        RECT 74.295 84.185 74.625 84.680 ;
        RECT 74.800 84.355 75.050 84.815 ;
        RECT 75.220 84.185 75.495 84.845 ;
        RECT 76.585 84.185 76.875 84.910 ;
        RECT 77.045 84.865 77.430 85.345 ;
        RECT 77.600 84.670 77.855 85.525 ;
        RECT 77.065 84.405 77.855 84.670 ;
        RECT 78.025 84.850 78.435 85.345 ;
        RECT 78.620 85.095 78.850 85.525 ;
        RECT 79.020 85.025 79.635 85.545 ;
        RECT 79.805 85.175 80.565 85.425 ;
        RECT 80.735 85.175 81.485 85.425 ;
        RECT 78.025 84.405 78.255 84.850 ;
        RECT 79.020 84.815 79.190 85.025 ;
        RECT 81.655 85.005 81.935 85.595 ;
        RECT 78.435 84.185 78.765 84.680 ;
        RECT 78.940 84.355 79.190 84.815 ;
        RECT 79.360 84.185 79.635 84.845 ;
        RECT 79.805 84.815 80.905 84.985 ;
        RECT 79.805 84.355 80.145 84.815 ;
        RECT 80.315 84.185 80.485 84.645 ;
        RECT 80.655 84.565 80.905 84.815 ;
        RECT 81.075 84.755 81.935 85.005 ;
        RECT 81.495 84.565 81.825 84.585 ;
        RECT 80.655 84.355 81.825 84.565 ;
        RECT 82.110 84.365 82.445 85.785 ;
        RECT 82.620 85.605 85.115 85.785 ;
        RECT 85.325 85.885 85.585 86.565 ;
        RECT 85.755 85.955 86.005 86.735 ;
        RECT 86.255 86.185 86.505 86.565 ;
        RECT 86.675 86.355 87.030 86.735 ;
        RECT 88.035 86.345 88.370 86.565 ;
        RECT 87.635 86.185 87.865 86.225 ;
        RECT 86.255 85.985 87.865 86.185 ;
        RECT 86.255 85.975 87.090 85.985 ;
        RECT 87.680 85.895 87.865 85.985 ;
        RECT 82.620 84.915 82.845 85.605 ;
        RECT 83.045 85.095 83.325 85.425 ;
        RECT 83.505 85.095 84.080 85.425 ;
        RECT 84.260 85.095 84.695 85.425 ;
        RECT 84.875 85.095 85.145 85.425 ;
        RECT 82.620 84.725 85.105 84.915 ;
        RECT 82.625 84.185 83.370 84.555 ;
        RECT 83.935 84.365 84.190 84.725 ;
        RECT 84.370 84.185 84.700 84.555 ;
        RECT 84.880 84.365 85.105 84.725 ;
        RECT 85.325 84.685 85.495 85.885 ;
        RECT 87.195 85.785 87.525 85.815 ;
        RECT 85.725 85.725 87.525 85.785 ;
        RECT 88.115 85.725 88.370 86.345 ;
        RECT 85.665 85.615 88.370 85.725 ;
        RECT 85.665 85.580 85.865 85.615 ;
        RECT 85.665 85.005 85.835 85.580 ;
        RECT 87.195 85.555 88.370 85.615 ;
        RECT 88.545 85.645 89.755 86.735 ;
        RECT 86.065 85.140 86.475 85.445 ;
        RECT 86.645 85.175 86.975 85.385 ;
        RECT 85.665 84.885 85.935 85.005 ;
        RECT 85.665 84.840 86.510 84.885 ;
        RECT 85.755 84.715 86.510 84.840 ;
        RECT 86.765 84.775 86.975 85.175 ;
        RECT 87.220 85.175 87.695 85.385 ;
        RECT 87.885 85.175 88.375 85.375 ;
        RECT 87.220 84.775 87.440 85.175 ;
        RECT 88.545 85.105 89.065 85.645 ;
        RECT 85.325 84.355 85.585 84.685 ;
        RECT 86.340 84.565 86.510 84.715 ;
        RECT 85.755 84.185 86.085 84.545 ;
        RECT 86.340 84.355 87.640 84.565 ;
        RECT 87.915 84.185 88.370 84.950 ;
        RECT 89.235 84.935 89.755 85.475 ;
        RECT 88.545 84.185 89.755 84.935 ;
        RECT 12.100 84.015 89.840 84.185 ;
        RECT 12.185 83.265 13.395 84.015 ;
        RECT 12.185 82.725 12.705 83.265 ;
        RECT 13.565 83.245 16.155 84.015 ;
        RECT 12.875 82.555 13.395 83.095 ;
        RECT 13.565 82.725 14.775 83.245 ;
        RECT 16.335 83.205 16.605 84.015 ;
        RECT 16.775 83.205 17.105 83.845 ;
        RECT 17.275 83.205 17.515 84.015 ;
        RECT 17.705 83.265 18.915 84.015 ;
        RECT 14.945 82.555 16.155 83.075 ;
        RECT 16.325 82.775 16.675 83.025 ;
        RECT 16.845 82.605 17.015 83.205 ;
        RECT 17.185 82.775 17.535 83.025 ;
        RECT 17.705 82.725 18.225 83.265 ;
        RECT 19.095 83.205 19.365 84.015 ;
        RECT 19.535 83.205 19.865 83.845 ;
        RECT 20.035 83.205 20.275 84.015 ;
        RECT 20.465 83.470 25.810 84.015 ;
        RECT 12.185 81.465 13.395 82.555 ;
        RECT 13.565 81.465 16.155 82.555 ;
        RECT 16.335 81.465 16.665 82.605 ;
        RECT 16.845 82.435 17.525 82.605 ;
        RECT 18.395 82.555 18.915 83.095 ;
        RECT 19.085 82.775 19.435 83.025 ;
        RECT 19.605 82.605 19.775 83.205 ;
        RECT 19.945 82.775 20.295 83.025 ;
        RECT 22.050 82.640 22.390 83.470 ;
        RECT 25.985 83.245 29.495 84.015 ;
        RECT 29.665 83.265 30.875 84.015 ;
        RECT 31.080 83.275 31.695 83.845 ;
        RECT 31.865 83.505 32.080 84.015 ;
        RECT 32.310 83.505 32.590 83.835 ;
        RECT 32.770 83.505 33.010 84.015 ;
        RECT 17.195 81.650 17.525 82.435 ;
        RECT 17.705 81.465 18.915 82.555 ;
        RECT 19.095 81.465 19.425 82.605 ;
        RECT 19.605 82.435 20.285 82.605 ;
        RECT 19.955 81.650 20.285 82.435 ;
        RECT 23.870 81.900 24.220 83.150 ;
        RECT 25.985 82.725 27.635 83.245 ;
        RECT 27.805 82.555 29.495 83.075 ;
        RECT 29.665 82.725 30.185 83.265 ;
        RECT 30.355 82.555 30.875 83.095 ;
        RECT 20.465 81.465 25.810 81.900 ;
        RECT 25.985 81.465 29.495 82.555 ;
        RECT 29.665 81.465 30.875 82.555 ;
        RECT 31.080 82.255 31.395 83.275 ;
        RECT 31.565 82.605 31.735 83.105 ;
        RECT 31.985 82.775 32.250 83.335 ;
        RECT 32.420 82.605 32.590 83.505 ;
        RECT 33.545 83.385 33.875 83.745 ;
        RECT 34.495 83.555 34.745 84.015 ;
        RECT 34.915 83.555 35.475 83.845 ;
        RECT 32.760 82.775 33.115 83.335 ;
        RECT 33.545 83.195 34.935 83.385 ;
        RECT 34.765 83.105 34.935 83.195 ;
        RECT 33.360 82.775 34.035 83.025 ;
        RECT 34.255 82.775 34.595 83.025 ;
        RECT 34.765 82.775 35.055 83.105 ;
        RECT 31.565 82.435 32.990 82.605 ;
        RECT 31.080 81.635 31.615 82.255 ;
        RECT 31.785 81.465 32.115 82.265 ;
        RECT 32.600 82.260 32.990 82.435 ;
        RECT 33.360 82.415 33.625 82.775 ;
        RECT 34.765 82.525 34.935 82.775 ;
        RECT 33.995 82.355 34.935 82.525 ;
        RECT 33.545 81.465 33.825 82.135 ;
        RECT 33.995 81.805 34.295 82.355 ;
        RECT 35.225 82.185 35.475 83.555 ;
        RECT 35.810 83.505 36.050 84.015 ;
        RECT 36.230 83.505 36.510 83.835 ;
        RECT 36.740 83.505 36.955 84.015 ;
        RECT 35.705 82.775 36.060 83.335 ;
        RECT 36.230 82.605 36.400 83.505 ;
        RECT 36.570 82.775 36.835 83.335 ;
        RECT 37.125 83.275 37.740 83.845 ;
        RECT 37.945 83.290 38.235 84.015 ;
        RECT 38.955 83.465 39.125 83.755 ;
        RECT 39.295 83.635 39.625 84.015 ;
        RECT 38.955 83.295 39.620 83.465 ;
        RECT 37.085 82.605 37.255 83.105 ;
        RECT 35.830 82.435 37.255 82.605 ;
        RECT 35.830 82.260 36.220 82.435 ;
        RECT 34.495 81.465 34.825 82.185 ;
        RECT 35.015 81.635 35.475 82.185 ;
        RECT 36.705 81.465 37.035 82.265 ;
        RECT 37.425 82.255 37.740 83.275 ;
        RECT 37.205 81.635 37.740 82.255 ;
        RECT 37.945 81.465 38.235 82.630 ;
        RECT 38.870 82.475 39.220 83.125 ;
        RECT 39.390 82.305 39.620 83.295 ;
        RECT 38.955 82.135 39.620 82.305 ;
        RECT 38.955 81.635 39.125 82.135 ;
        RECT 39.295 81.465 39.625 81.965 ;
        RECT 39.795 81.635 39.980 83.755 ;
        RECT 40.235 83.555 40.485 84.015 ;
        RECT 40.655 83.565 40.990 83.735 ;
        RECT 41.185 83.565 41.860 83.735 ;
        RECT 40.655 83.425 40.825 83.565 ;
        RECT 40.150 82.435 40.430 83.385 ;
        RECT 40.600 83.295 40.825 83.425 ;
        RECT 40.600 82.190 40.770 83.295 ;
        RECT 40.995 83.145 41.520 83.365 ;
        RECT 40.940 82.380 41.180 82.975 ;
        RECT 41.350 82.445 41.520 83.145 ;
        RECT 41.690 82.785 41.860 83.565 ;
        RECT 42.180 83.515 42.550 84.015 ;
        RECT 42.730 83.565 43.135 83.735 ;
        RECT 43.305 83.565 44.090 83.735 ;
        RECT 42.730 83.335 42.900 83.565 ;
        RECT 42.070 83.035 42.900 83.335 ;
        RECT 43.285 83.065 43.750 83.395 ;
        RECT 42.070 83.005 42.270 83.035 ;
        RECT 42.390 82.785 42.560 82.855 ;
        RECT 41.690 82.615 42.560 82.785 ;
        RECT 42.050 82.525 42.560 82.615 ;
        RECT 40.600 82.060 40.905 82.190 ;
        RECT 41.350 82.080 41.880 82.445 ;
        RECT 40.220 81.465 40.485 81.925 ;
        RECT 40.655 81.635 40.905 82.060 ;
        RECT 42.050 81.910 42.220 82.525 ;
        RECT 41.115 81.740 42.220 81.910 ;
        RECT 42.390 81.465 42.560 82.265 ;
        RECT 42.730 81.965 42.900 83.035 ;
        RECT 43.070 82.135 43.260 82.855 ;
        RECT 43.430 82.105 43.750 83.065 ;
        RECT 43.920 83.105 44.090 83.565 ;
        RECT 44.365 83.485 44.575 84.015 ;
        RECT 44.835 83.275 45.165 83.800 ;
        RECT 45.335 83.405 45.505 84.015 ;
        RECT 45.675 83.360 46.005 83.795 ;
        RECT 45.675 83.275 46.055 83.360 ;
        RECT 44.965 83.105 45.165 83.275 ;
        RECT 45.830 83.235 46.055 83.275 ;
        RECT 43.920 82.775 44.795 83.105 ;
        RECT 44.965 82.775 45.715 83.105 ;
        RECT 42.730 81.635 42.980 81.965 ;
        RECT 43.920 81.935 44.090 82.775 ;
        RECT 44.965 82.570 45.155 82.775 ;
        RECT 45.885 82.655 46.055 83.235 ;
        RECT 46.225 83.265 47.435 84.015 ;
        RECT 47.695 83.465 47.865 83.755 ;
        RECT 48.035 83.635 48.365 84.015 ;
        RECT 47.695 83.295 48.360 83.465 ;
        RECT 46.225 82.725 46.745 83.265 ;
        RECT 45.840 82.605 46.055 82.655 ;
        RECT 44.260 82.195 45.155 82.570 ;
        RECT 45.665 82.525 46.055 82.605 ;
        RECT 46.915 82.555 47.435 83.095 ;
        RECT 43.205 81.765 44.090 81.935 ;
        RECT 44.270 81.465 44.585 81.965 ;
        RECT 44.815 81.635 45.155 82.195 ;
        RECT 45.325 81.465 45.495 82.475 ;
        RECT 45.665 81.680 45.995 82.525 ;
        RECT 46.225 81.465 47.435 82.555 ;
        RECT 47.610 82.475 47.960 83.125 ;
        RECT 48.130 82.305 48.360 83.295 ;
        RECT 47.695 82.135 48.360 82.305 ;
        RECT 47.695 81.635 47.865 82.135 ;
        RECT 48.035 81.465 48.365 81.965 ;
        RECT 48.535 81.635 48.720 83.755 ;
        RECT 48.975 83.555 49.225 84.015 ;
        RECT 49.395 83.565 49.730 83.735 ;
        RECT 49.925 83.565 50.600 83.735 ;
        RECT 49.395 83.425 49.565 83.565 ;
        RECT 48.890 82.435 49.170 83.385 ;
        RECT 49.340 83.295 49.565 83.425 ;
        RECT 49.340 82.190 49.510 83.295 ;
        RECT 49.735 83.145 50.260 83.365 ;
        RECT 49.680 82.380 49.920 82.975 ;
        RECT 50.090 82.445 50.260 83.145 ;
        RECT 50.430 82.785 50.600 83.565 ;
        RECT 50.920 83.515 51.290 84.015 ;
        RECT 51.470 83.565 51.875 83.735 ;
        RECT 52.045 83.565 52.830 83.735 ;
        RECT 51.470 83.335 51.640 83.565 ;
        RECT 50.810 83.035 51.640 83.335 ;
        RECT 52.025 83.065 52.490 83.395 ;
        RECT 50.810 83.005 51.010 83.035 ;
        RECT 51.130 82.785 51.300 82.855 ;
        RECT 50.430 82.615 51.300 82.785 ;
        RECT 50.790 82.525 51.300 82.615 ;
        RECT 49.340 82.060 49.645 82.190 ;
        RECT 50.090 82.080 50.620 82.445 ;
        RECT 48.960 81.465 49.225 81.925 ;
        RECT 49.395 81.635 49.645 82.060 ;
        RECT 50.790 81.910 50.960 82.525 ;
        RECT 49.855 81.740 50.960 81.910 ;
        RECT 51.130 81.465 51.300 82.265 ;
        RECT 51.470 81.965 51.640 83.035 ;
        RECT 51.810 82.135 52.000 82.855 ;
        RECT 52.170 82.105 52.490 83.065 ;
        RECT 52.660 83.105 52.830 83.565 ;
        RECT 53.105 83.485 53.315 84.015 ;
        RECT 53.575 83.275 53.905 83.800 ;
        RECT 54.075 83.405 54.245 84.015 ;
        RECT 54.415 83.360 54.745 83.795 ;
        RECT 54.970 83.540 55.305 83.800 ;
        RECT 55.475 83.615 55.805 84.015 ;
        RECT 55.975 83.615 57.590 83.785 ;
        RECT 54.415 83.275 54.795 83.360 ;
        RECT 53.705 83.105 53.905 83.275 ;
        RECT 54.570 83.235 54.795 83.275 ;
        RECT 52.660 82.775 53.535 83.105 ;
        RECT 53.705 82.775 54.455 83.105 ;
        RECT 51.470 81.635 51.720 81.965 ;
        RECT 52.660 81.935 52.830 82.775 ;
        RECT 53.705 82.570 53.895 82.775 ;
        RECT 54.625 82.655 54.795 83.235 ;
        RECT 54.580 82.605 54.795 82.655 ;
        RECT 53.000 82.195 53.895 82.570 ;
        RECT 54.405 82.525 54.795 82.605 ;
        RECT 51.945 81.765 52.830 81.935 ;
        RECT 53.010 81.465 53.325 81.965 ;
        RECT 53.555 81.635 53.895 82.195 ;
        RECT 54.065 81.465 54.235 82.475 ;
        RECT 54.405 81.680 54.735 82.525 ;
        RECT 54.970 82.185 55.225 83.540 ;
        RECT 55.975 83.445 56.145 83.615 ;
        RECT 55.585 83.275 56.145 83.445 ;
        RECT 56.410 83.335 56.680 83.435 ;
        RECT 56.870 83.335 57.160 83.435 ;
        RECT 55.585 83.105 55.755 83.275 ;
        RECT 56.405 83.165 56.680 83.335 ;
        RECT 56.865 83.165 57.160 83.335 ;
        RECT 55.450 82.775 55.755 83.105 ;
        RECT 55.950 82.995 56.200 83.105 ;
        RECT 55.945 82.825 56.200 82.995 ;
        RECT 55.950 82.775 56.200 82.825 ;
        RECT 56.410 82.775 56.680 83.165 ;
        RECT 56.870 82.775 57.160 83.165 ;
        RECT 57.330 82.775 57.750 83.440 ;
        RECT 58.135 83.295 58.465 84.015 ;
        RECT 58.645 83.215 58.955 84.015 ;
        RECT 59.160 83.215 59.855 83.845 ;
        RECT 60.230 83.235 60.730 83.845 ;
        RECT 58.060 82.775 58.410 83.105 ;
        RECT 58.655 82.775 58.990 83.045 ;
        RECT 55.585 82.605 55.755 82.775 ;
        RECT 58.205 82.655 58.410 82.775 ;
        RECT 55.585 82.435 57.955 82.605 ;
        RECT 58.205 82.485 58.415 82.655 ;
        RECT 59.160 82.615 59.330 83.215 ;
        RECT 59.500 82.775 59.835 83.025 ;
        RECT 60.025 82.775 60.375 83.025 ;
        RECT 54.970 81.675 55.305 82.185 ;
        RECT 55.555 81.465 55.885 82.265 ;
        RECT 56.130 82.055 57.555 82.225 ;
        RECT 56.130 81.635 56.415 82.055 ;
        RECT 56.670 81.465 57.000 81.885 ;
        RECT 57.225 81.805 57.555 82.055 ;
        RECT 57.785 81.975 57.955 82.435 ;
        RECT 58.215 81.805 58.385 82.305 ;
        RECT 57.225 81.635 58.385 81.805 ;
        RECT 58.645 81.465 58.925 82.605 ;
        RECT 59.095 81.635 59.425 82.615 ;
        RECT 60.560 82.605 60.730 83.235 ;
        RECT 61.360 83.365 61.690 83.845 ;
        RECT 61.860 83.555 62.085 84.015 ;
        RECT 62.255 83.365 62.585 83.845 ;
        RECT 61.360 83.195 62.585 83.365 ;
        RECT 62.775 83.215 63.025 84.015 ;
        RECT 63.195 83.215 63.535 83.845 ;
        RECT 63.705 83.290 63.995 84.015 ;
        RECT 64.170 83.250 64.625 84.015 ;
        RECT 64.900 83.635 66.200 83.845 ;
        RECT 66.455 83.655 66.785 84.015 ;
        RECT 66.030 83.485 66.200 83.635 ;
        RECT 66.955 83.515 67.215 83.845 ;
        RECT 66.985 83.505 67.215 83.515 ;
        RECT 60.900 82.825 61.230 83.025 ;
        RECT 61.400 82.825 61.730 83.025 ;
        RECT 61.900 82.825 62.320 83.025 ;
        RECT 62.495 82.855 63.190 83.025 ;
        RECT 62.495 82.605 62.665 82.855 ;
        RECT 63.360 82.605 63.535 83.215 ;
        RECT 65.100 83.025 65.320 83.425 ;
        RECT 64.165 82.825 64.655 83.025 ;
        RECT 64.845 82.815 65.320 83.025 ;
        RECT 65.565 83.025 65.775 83.425 ;
        RECT 66.030 83.360 66.785 83.485 ;
        RECT 66.030 83.315 66.875 83.360 ;
        RECT 66.605 83.195 66.875 83.315 ;
        RECT 65.565 82.815 65.895 83.025 ;
        RECT 66.065 82.755 66.475 83.060 ;
        RECT 59.595 81.465 59.855 82.605 ;
        RECT 60.230 82.435 62.665 82.605 ;
        RECT 60.230 81.635 60.560 82.435 ;
        RECT 60.730 81.465 61.060 82.265 ;
        RECT 61.360 81.635 61.690 82.435 ;
        RECT 62.335 81.465 62.585 82.265 ;
        RECT 62.855 81.465 63.025 82.605 ;
        RECT 63.195 81.635 63.535 82.605 ;
        RECT 63.705 81.465 63.995 82.630 ;
        RECT 64.170 82.585 65.345 82.645 ;
        RECT 66.705 82.620 66.875 83.195 ;
        RECT 66.675 82.585 66.875 82.620 ;
        RECT 64.170 82.475 66.875 82.585 ;
        RECT 64.170 81.855 64.425 82.475 ;
        RECT 65.015 82.415 66.815 82.475 ;
        RECT 65.015 82.385 65.345 82.415 ;
        RECT 67.045 82.315 67.215 83.505 ;
        RECT 64.675 82.215 64.860 82.305 ;
        RECT 65.450 82.215 66.285 82.225 ;
        RECT 64.675 82.015 66.285 82.215 ;
        RECT 64.675 81.975 64.905 82.015 ;
        RECT 64.170 81.635 64.505 81.855 ;
        RECT 65.510 81.465 65.865 81.845 ;
        RECT 66.035 81.635 66.285 82.015 ;
        RECT 66.535 81.465 66.785 82.245 ;
        RECT 66.955 81.635 67.215 82.315 ;
        RECT 67.390 83.275 67.645 83.845 ;
        RECT 67.815 83.615 68.145 84.015 ;
        RECT 68.570 83.480 69.100 83.845 ;
        RECT 68.570 83.445 68.745 83.480 ;
        RECT 67.815 83.275 68.745 83.445 ;
        RECT 67.390 82.605 67.560 83.275 ;
        RECT 67.815 83.105 67.985 83.275 ;
        RECT 67.730 82.775 67.985 83.105 ;
        RECT 68.210 82.775 68.405 83.105 ;
        RECT 67.390 81.635 67.725 82.605 ;
        RECT 67.895 81.465 68.065 82.605 ;
        RECT 68.235 81.805 68.405 82.775 ;
        RECT 68.575 82.145 68.745 83.275 ;
        RECT 68.915 82.485 69.085 83.285 ;
        RECT 69.290 82.995 69.565 83.845 ;
        RECT 69.285 82.825 69.565 82.995 ;
        RECT 69.290 82.685 69.565 82.825 ;
        RECT 69.735 82.485 69.925 83.845 ;
        RECT 70.105 83.480 70.615 84.015 ;
        RECT 70.835 83.205 71.080 83.810 ;
        RECT 71.525 83.275 71.910 83.845 ;
        RECT 72.080 83.555 72.405 84.015 ;
        RECT 72.925 83.385 73.205 83.845 ;
        RECT 70.125 83.035 71.355 83.205 ;
        RECT 68.915 82.315 69.925 82.485 ;
        RECT 70.095 82.470 70.845 82.660 ;
        RECT 68.575 81.975 69.700 82.145 ;
        RECT 70.095 81.805 70.265 82.470 ;
        RECT 71.015 82.225 71.355 83.035 ;
        RECT 68.235 81.635 70.265 81.805 ;
        RECT 70.435 81.465 70.605 82.225 ;
        RECT 70.840 81.815 71.355 82.225 ;
        RECT 71.525 82.605 71.805 83.275 ;
        RECT 72.080 83.215 73.205 83.385 ;
        RECT 72.080 83.105 72.530 83.215 ;
        RECT 71.975 82.775 72.530 83.105 ;
        RECT 73.395 83.045 73.795 83.845 ;
        RECT 74.195 83.555 74.465 84.015 ;
        RECT 74.635 83.385 74.920 83.845 ;
        RECT 71.525 81.635 71.910 82.605 ;
        RECT 72.080 82.315 72.530 82.775 ;
        RECT 72.700 82.485 73.795 83.045 ;
        RECT 72.080 82.095 73.205 82.315 ;
        RECT 72.080 81.465 72.405 81.925 ;
        RECT 72.925 81.635 73.205 82.095 ;
        RECT 73.395 81.635 73.795 82.485 ;
        RECT 73.965 83.215 74.920 83.385 ;
        RECT 75.865 83.385 76.195 83.745 ;
        RECT 76.825 83.555 77.075 84.015 ;
        RECT 77.245 83.555 77.795 83.845 ;
        RECT 73.965 82.315 74.175 83.215 ;
        RECT 75.865 83.195 77.255 83.385 ;
        RECT 77.085 83.105 77.255 83.195 ;
        RECT 74.345 82.485 75.035 83.045 ;
        RECT 75.665 82.775 76.355 83.025 ;
        RECT 76.585 82.775 76.915 83.025 ;
        RECT 77.085 82.775 77.375 83.105 ;
        RECT 75.665 82.335 75.980 82.775 ;
        RECT 77.085 82.525 77.255 82.775 ;
        RECT 76.315 82.355 77.255 82.525 ;
        RECT 73.965 82.095 74.920 82.315 ;
        RECT 74.195 81.465 74.465 81.925 ;
        RECT 74.635 81.635 74.920 82.095 ;
        RECT 75.865 81.465 76.145 82.135 ;
        RECT 76.315 81.805 76.615 82.355 ;
        RECT 77.545 82.185 77.795 83.555 ;
        RECT 77.965 83.215 78.255 84.015 ;
        RECT 78.425 83.215 78.765 83.845 ;
        RECT 78.935 83.215 79.185 84.015 ;
        RECT 79.375 83.365 79.705 83.845 ;
        RECT 79.875 83.555 80.100 84.015 ;
        RECT 80.270 83.365 80.600 83.845 ;
        RECT 78.425 82.605 78.600 83.215 ;
        RECT 79.375 83.195 80.600 83.365 ;
        RECT 81.230 83.235 81.730 83.845 ;
        RECT 78.770 82.855 79.465 83.025 ;
        RECT 79.295 82.605 79.465 82.855 ;
        RECT 79.640 82.825 80.060 83.025 ;
        RECT 80.230 82.825 80.560 83.025 ;
        RECT 80.730 82.825 81.060 83.025 ;
        RECT 81.230 82.605 81.400 83.235 ;
        RECT 82.105 83.215 82.445 83.845 ;
        RECT 82.615 83.215 82.865 84.015 ;
        RECT 83.055 83.365 83.385 83.845 ;
        RECT 83.555 83.555 83.780 84.015 ;
        RECT 83.950 83.365 84.280 83.845 ;
        RECT 81.585 82.775 81.935 83.025 ;
        RECT 82.105 82.605 82.280 83.215 ;
        RECT 83.055 83.195 84.280 83.365 ;
        RECT 84.910 83.235 85.410 83.845 ;
        RECT 85.820 83.275 86.435 83.845 ;
        RECT 86.605 83.505 86.820 84.015 ;
        RECT 87.050 83.505 87.330 83.835 ;
        RECT 87.510 83.505 87.750 84.015 ;
        RECT 82.450 82.855 83.145 83.025 ;
        RECT 82.975 82.605 83.145 82.855 ;
        RECT 83.320 82.825 83.740 83.025 ;
        RECT 83.910 82.825 84.240 83.025 ;
        RECT 84.410 82.825 84.740 83.025 ;
        RECT 84.910 82.605 85.080 83.235 ;
        RECT 85.265 82.775 85.615 83.025 ;
        RECT 76.825 81.465 77.155 82.185 ;
        RECT 77.345 81.635 77.795 82.185 ;
        RECT 77.965 81.465 78.255 82.605 ;
        RECT 78.425 81.635 78.765 82.605 ;
        RECT 78.935 81.465 79.105 82.605 ;
        RECT 79.295 82.435 81.730 82.605 ;
        RECT 79.375 81.465 79.625 82.265 ;
        RECT 80.270 81.635 80.600 82.435 ;
        RECT 80.900 81.465 81.230 82.265 ;
        RECT 81.400 81.635 81.730 82.435 ;
        RECT 82.105 81.635 82.445 82.605 ;
        RECT 82.615 81.465 82.785 82.605 ;
        RECT 82.975 82.435 85.410 82.605 ;
        RECT 83.055 81.465 83.305 82.265 ;
        RECT 83.950 81.635 84.280 82.435 ;
        RECT 84.580 81.465 84.910 82.265 ;
        RECT 85.080 81.635 85.410 82.435 ;
        RECT 85.820 82.255 86.135 83.275 ;
        RECT 86.305 82.605 86.475 83.105 ;
        RECT 86.725 82.775 86.990 83.335 ;
        RECT 87.160 82.605 87.330 83.505 ;
        RECT 87.500 82.775 87.855 83.335 ;
        RECT 88.545 83.265 89.755 84.015 ;
        RECT 86.305 82.435 87.730 82.605 ;
        RECT 85.820 81.635 86.355 82.255 ;
        RECT 86.525 81.465 86.855 82.265 ;
        RECT 87.340 82.260 87.730 82.435 ;
        RECT 88.545 82.555 89.065 83.095 ;
        RECT 89.235 82.725 89.755 83.265 ;
        RECT 88.545 81.465 89.755 82.555 ;
        RECT 12.100 81.295 89.840 81.465 ;
        RECT 12.185 80.205 13.395 81.295 ;
        RECT 13.565 80.860 18.910 81.295 ;
        RECT 12.185 79.495 12.705 80.035 ;
        RECT 12.875 79.665 13.395 80.205 ;
        RECT 12.185 78.745 13.395 79.495 ;
        RECT 15.150 79.290 15.490 80.120 ;
        RECT 16.970 79.610 17.320 80.860 ;
        RECT 19.085 80.205 22.595 81.295 ;
        RECT 19.085 79.515 20.735 80.035 ;
        RECT 20.905 79.685 22.595 80.205 ;
        RECT 23.265 80.155 23.495 81.295 ;
        RECT 23.665 80.145 23.995 81.125 ;
        RECT 24.165 80.155 24.375 81.295 ;
        RECT 23.245 79.735 23.575 79.985 ;
        RECT 13.565 78.745 18.910 79.290 ;
        RECT 19.085 78.745 22.595 79.515 ;
        RECT 23.265 78.745 23.495 79.565 ;
        RECT 23.745 79.545 23.995 80.145 ;
        RECT 25.065 80.130 25.355 81.295 ;
        RECT 25.525 80.205 27.195 81.295 ;
        RECT 27.830 80.495 28.145 81.295 ;
        RECT 28.410 80.940 29.490 81.110 ;
        RECT 28.410 80.325 28.580 80.940 ;
        RECT 23.665 78.915 23.995 79.545 ;
        RECT 24.165 78.745 24.375 79.565 ;
        RECT 25.525 79.515 26.275 80.035 ;
        RECT 26.445 79.685 27.195 80.205 ;
        RECT 25.065 78.745 25.355 79.470 ;
        RECT 25.525 78.745 27.195 79.515 ;
        RECT 27.825 79.315 28.095 80.325 ;
        RECT 28.265 80.155 28.580 80.325 ;
        RECT 28.265 79.485 28.435 80.155 ;
        RECT 28.750 79.985 28.985 80.665 ;
        RECT 29.155 80.155 29.490 80.940 ;
        RECT 29.710 80.155 30.005 81.295 ;
        RECT 30.265 80.325 30.595 81.125 ;
        RECT 30.765 80.495 30.935 81.295 ;
        RECT 31.105 80.325 31.435 81.125 ;
        RECT 31.605 80.495 31.775 81.295 ;
        RECT 31.945 80.345 32.275 81.125 ;
        RECT 32.445 80.835 32.615 81.295 ;
        RECT 31.945 80.325 32.715 80.345 ;
        RECT 30.265 80.155 32.715 80.325 ;
        RECT 28.605 79.655 28.985 79.985 ;
        RECT 29.155 79.655 29.490 79.985 ;
        RECT 29.685 79.735 32.195 79.985 ;
        RECT 32.365 79.565 32.715 80.155 ;
        RECT 28.265 79.315 29.490 79.485 ;
        RECT 27.895 78.745 28.225 79.145 ;
        RECT 28.395 79.045 28.565 79.315 ;
        RECT 28.735 78.745 29.065 79.145 ;
        RECT 29.235 79.045 29.490 79.315 ;
        RECT 30.345 79.385 32.715 79.565 ;
        RECT 32.885 79.690 33.165 81.125 ;
        RECT 33.335 80.520 34.045 81.295 ;
        RECT 34.215 80.350 34.545 81.125 ;
        RECT 33.395 80.135 34.545 80.350 ;
        RECT 29.710 78.745 29.975 79.205 ;
        RECT 30.345 78.915 30.515 79.385 ;
        RECT 30.765 78.745 30.935 79.205 ;
        RECT 31.185 78.915 31.355 79.385 ;
        RECT 31.605 78.745 31.775 79.205 ;
        RECT 32.025 78.915 32.195 79.385 ;
        RECT 32.365 78.745 32.615 79.210 ;
        RECT 32.885 78.915 33.225 79.690 ;
        RECT 33.395 79.565 33.680 80.135 ;
        RECT 33.865 79.735 34.335 79.965 ;
        RECT 34.740 79.935 34.955 81.050 ;
        RECT 35.135 80.575 35.465 81.295 ;
        RECT 35.245 79.935 35.475 80.275 ;
        RECT 34.505 79.755 34.955 79.935 ;
        RECT 34.505 79.735 34.835 79.755 ;
        RECT 35.145 79.735 35.475 79.935 ;
        RECT 35.645 79.690 35.925 81.125 ;
        RECT 36.095 80.520 36.805 81.295 ;
        RECT 36.975 80.350 37.305 81.125 ;
        RECT 36.155 80.135 37.305 80.350 ;
        RECT 33.395 79.375 34.105 79.565 ;
        RECT 33.805 79.235 34.105 79.375 ;
        RECT 34.295 79.375 35.475 79.565 ;
        RECT 34.295 79.295 34.625 79.375 ;
        RECT 33.805 79.225 34.120 79.235 ;
        RECT 33.805 79.215 34.130 79.225 ;
        RECT 33.805 79.210 34.140 79.215 ;
        RECT 33.395 78.745 33.565 79.205 ;
        RECT 33.805 79.200 34.145 79.210 ;
        RECT 33.805 79.195 34.150 79.200 ;
        RECT 33.805 79.185 34.155 79.195 ;
        RECT 33.805 79.180 34.160 79.185 ;
        RECT 33.805 78.915 34.165 79.180 ;
        RECT 34.795 78.745 34.965 79.205 ;
        RECT 35.135 78.915 35.475 79.375 ;
        RECT 35.645 78.915 35.985 79.690 ;
        RECT 36.155 79.565 36.440 80.135 ;
        RECT 36.625 79.735 37.095 79.965 ;
        RECT 37.500 79.935 37.715 81.050 ;
        RECT 37.895 80.575 38.225 81.295 ;
        RECT 38.885 80.405 39.145 81.115 ;
        RECT 39.315 80.585 39.645 81.295 ;
        RECT 39.815 80.405 40.045 81.115 ;
        RECT 38.005 79.935 38.235 80.275 ;
        RECT 38.885 80.165 40.045 80.405 ;
        RECT 40.225 80.385 40.495 81.115 ;
        RECT 40.675 80.565 41.015 81.295 ;
        RECT 40.225 80.165 40.995 80.385 ;
        RECT 37.265 79.755 37.715 79.935 ;
        RECT 37.265 79.735 37.595 79.755 ;
        RECT 37.905 79.735 38.235 79.935 ;
        RECT 38.875 79.655 39.175 79.985 ;
        RECT 39.355 79.675 39.880 79.985 ;
        RECT 40.060 79.675 40.525 79.985 ;
        RECT 36.155 79.375 36.865 79.565 ;
        RECT 36.565 79.235 36.865 79.375 ;
        RECT 37.055 79.375 38.235 79.565 ;
        RECT 37.055 79.295 37.385 79.375 ;
        RECT 36.565 79.225 36.880 79.235 ;
        RECT 36.565 79.215 36.890 79.225 ;
        RECT 36.565 79.210 36.900 79.215 ;
        RECT 36.155 78.745 36.325 79.205 ;
        RECT 36.565 79.200 36.905 79.210 ;
        RECT 36.565 79.195 36.910 79.200 ;
        RECT 36.565 79.185 36.915 79.195 ;
        RECT 36.565 79.180 36.920 79.185 ;
        RECT 36.565 78.915 36.925 79.180 ;
        RECT 37.555 78.745 37.725 79.205 ;
        RECT 37.895 78.915 38.235 79.375 ;
        RECT 38.885 78.745 39.175 79.475 ;
        RECT 39.355 79.035 39.585 79.675 ;
        RECT 40.705 79.495 40.995 80.165 ;
        RECT 39.765 79.295 40.995 79.495 ;
        RECT 39.765 78.925 40.075 79.295 ;
        RECT 40.255 78.745 40.925 79.115 ;
        RECT 41.185 78.925 41.445 81.115 ;
        RECT 41.625 80.205 43.295 81.295 ;
        RECT 43.465 80.460 43.810 81.295 ;
        RECT 43.985 80.290 44.240 81.095 ;
        RECT 44.410 80.460 44.670 81.295 ;
        RECT 44.845 80.290 45.100 81.095 ;
        RECT 45.270 80.460 45.530 81.295 ;
        RECT 45.700 80.290 45.960 81.095 ;
        RECT 46.130 80.460 46.515 81.295 ;
        RECT 46.690 80.725 47.010 81.125 ;
        RECT 41.625 79.515 42.375 80.035 ;
        RECT 42.545 79.685 43.295 80.205 ;
        RECT 43.485 80.120 46.515 80.290 ;
        RECT 43.485 79.555 43.655 80.120 ;
        RECT 43.825 79.725 46.040 79.950 ;
        RECT 46.215 79.555 46.515 80.120 ;
        RECT 41.625 78.745 43.295 79.515 ;
        RECT 43.485 79.385 46.515 79.555 ;
        RECT 46.690 80.275 46.860 80.725 ;
        RECT 47.180 80.495 47.490 81.295 ;
        RECT 47.660 80.665 47.990 81.125 ;
        RECT 48.160 80.835 48.330 81.295 ;
        RECT 48.500 80.665 48.830 81.125 ;
        RECT 49.000 80.835 49.250 81.295 ;
        RECT 49.440 80.835 49.690 81.295 ;
        RECT 47.660 80.615 48.830 80.665 ;
        RECT 49.860 80.665 50.110 81.125 ;
        RECT 50.360 80.835 50.650 81.295 ;
        RECT 49.860 80.615 50.650 80.665 ;
        RECT 47.660 80.445 50.650 80.615 ;
        RECT 46.690 80.105 50.250 80.275 ;
        RECT 43.945 78.745 44.240 79.215 ;
        RECT 44.410 78.940 44.670 79.385 ;
        RECT 44.840 78.745 45.100 79.215 ;
        RECT 45.270 78.940 45.525 79.385 ;
        RECT 46.690 79.315 46.860 80.105 ;
        RECT 47.030 79.735 47.380 79.935 ;
        RECT 47.660 79.735 48.340 79.935 ;
        RECT 48.550 79.735 49.740 79.935 ;
        RECT 49.920 79.735 50.250 80.105 ;
        RECT 50.450 79.565 50.650 80.445 ;
        RECT 50.825 80.130 51.115 81.295 ;
        RECT 51.290 80.155 51.625 81.125 ;
        RECT 51.795 80.155 51.965 81.295 ;
        RECT 52.135 80.955 54.165 81.125 ;
        RECT 45.695 78.745 45.995 79.215 ;
        RECT 46.690 78.915 47.010 79.315 ;
        RECT 47.180 78.745 47.490 79.565 ;
        RECT 47.660 79.375 49.350 79.565 ;
        RECT 47.660 78.915 47.990 79.375 ;
        RECT 48.600 79.295 49.350 79.375 ;
        RECT 48.160 78.745 48.410 79.205 ;
        RECT 49.520 79.125 49.690 79.565 ;
        RECT 49.860 79.295 50.650 79.565 ;
        RECT 51.290 79.485 51.460 80.155 ;
        RECT 52.135 79.985 52.305 80.955 ;
        RECT 51.630 79.655 51.885 79.985 ;
        RECT 52.110 79.655 52.305 79.985 ;
        RECT 52.475 80.615 53.600 80.785 ;
        RECT 51.715 79.485 51.885 79.655 ;
        RECT 52.475 79.485 52.645 80.615 ;
        RECT 48.600 78.915 50.650 79.125 ;
        RECT 50.825 78.745 51.115 79.470 ;
        RECT 51.290 78.915 51.545 79.485 ;
        RECT 51.715 79.315 52.645 79.485 ;
        RECT 52.815 80.275 53.825 80.445 ;
        RECT 52.815 79.475 52.985 80.275 ;
        RECT 53.190 79.935 53.465 80.075 ;
        RECT 53.185 79.765 53.465 79.935 ;
        RECT 52.470 79.280 52.645 79.315 ;
        RECT 51.715 78.745 52.045 79.145 ;
        RECT 52.470 78.915 53.000 79.280 ;
        RECT 53.190 78.915 53.465 79.765 ;
        RECT 53.635 78.915 53.825 80.275 ;
        RECT 53.995 80.290 54.165 80.955 ;
        RECT 54.335 80.535 54.505 81.295 ;
        RECT 54.740 80.535 55.255 80.945 ;
        RECT 53.995 80.100 54.745 80.290 ;
        RECT 54.915 79.725 55.255 80.535 ;
        RECT 55.425 80.205 56.635 81.295 ;
        RECT 56.805 80.785 57.065 81.295 ;
        RECT 54.025 79.555 55.255 79.725 ;
        RECT 54.005 78.745 54.515 79.280 ;
        RECT 54.735 78.950 54.980 79.555 ;
        RECT 55.425 79.495 55.945 80.035 ;
        RECT 56.115 79.665 56.635 80.205 ;
        RECT 56.805 79.735 57.145 80.615 ;
        RECT 57.315 79.905 57.485 81.125 ;
        RECT 57.725 80.790 58.340 81.295 ;
        RECT 57.725 80.255 57.975 80.620 ;
        RECT 58.145 80.615 58.340 80.790 ;
        RECT 58.510 80.785 58.985 81.125 ;
        RECT 59.155 80.750 59.370 81.295 ;
        RECT 58.145 80.425 58.475 80.615 ;
        RECT 58.695 80.255 59.410 80.550 ;
        RECT 59.580 80.425 59.855 81.125 ;
        RECT 60.025 80.785 61.215 81.075 ;
        RECT 57.725 80.085 59.515 80.255 ;
        RECT 57.315 79.655 58.110 79.905 ;
        RECT 57.315 79.565 57.565 79.655 ;
        RECT 55.425 78.745 56.635 79.495 ;
        RECT 56.805 78.745 57.065 79.565 ;
        RECT 57.235 79.145 57.565 79.565 ;
        RECT 58.280 79.230 58.535 80.085 ;
        RECT 57.745 78.965 58.535 79.230 ;
        RECT 58.705 79.385 59.115 79.905 ;
        RECT 59.285 79.655 59.515 80.085 ;
        RECT 59.685 79.395 59.855 80.425 ;
        RECT 60.045 80.445 61.215 80.615 ;
        RECT 61.385 80.495 61.665 81.295 ;
        RECT 60.045 80.155 60.370 80.445 ;
        RECT 61.045 80.325 61.215 80.445 ;
        RECT 60.540 79.985 60.735 80.275 ;
        RECT 61.045 80.155 61.705 80.325 ;
        RECT 61.875 80.155 62.150 81.125 ;
        RECT 61.535 79.985 61.705 80.155 ;
        RECT 60.025 79.655 60.370 79.985 ;
        RECT 60.540 79.655 61.365 79.985 ;
        RECT 61.535 79.655 61.810 79.985 ;
        RECT 61.535 79.485 61.705 79.655 ;
        RECT 58.705 78.965 58.905 79.385 ;
        RECT 59.095 78.745 59.425 79.205 ;
        RECT 59.595 78.915 59.855 79.395 ;
        RECT 60.040 79.315 61.705 79.485 ;
        RECT 61.980 79.420 62.150 80.155 ;
        RECT 62.330 80.905 62.665 81.125 ;
        RECT 63.670 80.915 64.025 81.295 ;
        RECT 62.330 80.285 62.585 80.905 ;
        RECT 62.835 80.745 63.065 80.785 ;
        RECT 64.195 80.745 64.445 81.125 ;
        RECT 62.835 80.545 64.445 80.745 ;
        RECT 62.835 80.455 63.020 80.545 ;
        RECT 63.610 80.535 64.445 80.545 ;
        RECT 64.695 80.515 64.945 81.295 ;
        RECT 65.115 80.445 65.375 81.125 ;
        RECT 65.635 80.625 65.805 81.125 ;
        RECT 65.975 80.795 66.305 81.295 ;
        RECT 65.635 80.455 66.300 80.625 ;
        RECT 63.175 80.345 63.505 80.375 ;
        RECT 63.175 80.285 64.975 80.345 ;
        RECT 62.330 80.175 65.035 80.285 ;
        RECT 62.330 80.115 63.505 80.175 ;
        RECT 64.835 80.140 65.035 80.175 ;
        RECT 62.325 79.735 62.815 79.935 ;
        RECT 63.005 79.735 63.480 79.945 ;
        RECT 60.040 78.965 60.295 79.315 ;
        RECT 60.465 78.745 60.795 79.145 ;
        RECT 60.965 78.965 61.135 79.315 ;
        RECT 61.305 78.745 61.685 79.145 ;
        RECT 61.875 79.075 62.150 79.420 ;
        RECT 62.330 78.745 62.785 79.510 ;
        RECT 63.260 79.335 63.480 79.735 ;
        RECT 63.725 79.735 64.055 79.945 ;
        RECT 63.725 79.335 63.935 79.735 ;
        RECT 64.225 79.700 64.635 80.005 ;
        RECT 64.865 79.565 65.035 80.140 ;
        RECT 64.765 79.445 65.035 79.565 ;
        RECT 64.190 79.400 65.035 79.445 ;
        RECT 64.190 79.275 64.945 79.400 ;
        RECT 64.190 79.125 64.360 79.275 ;
        RECT 65.205 79.255 65.375 80.445 ;
        RECT 65.550 79.635 65.900 80.285 ;
        RECT 66.070 79.465 66.300 80.455 ;
        RECT 65.145 79.245 65.375 79.255 ;
        RECT 63.060 78.915 64.360 79.125 ;
        RECT 64.615 78.745 64.945 79.105 ;
        RECT 65.115 78.915 65.375 79.245 ;
        RECT 65.635 79.295 66.300 79.465 ;
        RECT 65.635 79.005 65.805 79.295 ;
        RECT 65.975 78.745 66.305 79.125 ;
        RECT 66.475 79.005 66.660 81.125 ;
        RECT 66.900 80.835 67.165 81.295 ;
        RECT 67.335 80.700 67.585 81.125 ;
        RECT 67.795 80.850 68.900 81.020 ;
        RECT 67.280 80.570 67.585 80.700 ;
        RECT 66.830 79.375 67.110 80.325 ;
        RECT 67.280 79.465 67.450 80.570 ;
        RECT 67.620 79.785 67.860 80.380 ;
        RECT 68.030 80.315 68.560 80.680 ;
        RECT 68.030 79.615 68.200 80.315 ;
        RECT 68.730 80.235 68.900 80.850 ;
        RECT 69.070 80.495 69.240 81.295 ;
        RECT 69.410 80.795 69.660 81.125 ;
        RECT 69.885 80.825 70.770 80.995 ;
        RECT 68.730 80.145 69.240 80.235 ;
        RECT 67.280 79.335 67.505 79.465 ;
        RECT 67.675 79.395 68.200 79.615 ;
        RECT 68.370 79.975 69.240 80.145 ;
        RECT 66.915 78.745 67.165 79.205 ;
        RECT 67.335 79.195 67.505 79.335 ;
        RECT 68.370 79.195 68.540 79.975 ;
        RECT 69.070 79.905 69.240 79.975 ;
        RECT 68.750 79.725 68.950 79.755 ;
        RECT 69.410 79.725 69.580 80.795 ;
        RECT 69.750 79.905 69.940 80.625 ;
        RECT 68.750 79.425 69.580 79.725 ;
        RECT 70.110 79.695 70.430 80.655 ;
        RECT 67.335 79.025 67.670 79.195 ;
        RECT 67.865 79.025 68.540 79.195 ;
        RECT 68.860 78.745 69.230 79.245 ;
        RECT 69.410 79.195 69.580 79.425 ;
        RECT 69.965 79.365 70.430 79.695 ;
        RECT 70.600 79.985 70.770 80.825 ;
        RECT 70.950 80.795 71.265 81.295 ;
        RECT 71.495 80.565 71.835 81.125 ;
        RECT 70.940 80.190 71.835 80.565 ;
        RECT 72.005 80.285 72.175 81.295 ;
        RECT 71.645 79.985 71.835 80.190 ;
        RECT 72.345 80.235 72.675 81.080 ;
        RECT 73.090 80.325 73.480 80.500 ;
        RECT 73.965 80.495 74.295 81.295 ;
        RECT 74.465 80.505 75.000 81.125 ;
        RECT 72.345 80.155 72.735 80.235 ;
        RECT 73.090 80.155 74.515 80.325 ;
        RECT 72.520 80.105 72.735 80.155 ;
        RECT 70.600 79.655 71.475 79.985 ;
        RECT 71.645 79.655 72.395 79.985 ;
        RECT 70.600 79.195 70.770 79.655 ;
        RECT 71.645 79.485 71.845 79.655 ;
        RECT 72.565 79.525 72.735 80.105 ;
        RECT 72.510 79.485 72.735 79.525 ;
        RECT 69.410 79.025 69.815 79.195 ;
        RECT 69.985 79.025 70.770 79.195 ;
        RECT 71.045 78.745 71.255 79.275 ;
        RECT 71.515 78.960 71.845 79.485 ;
        RECT 72.355 79.400 72.735 79.485 ;
        RECT 72.965 79.425 73.320 79.985 ;
        RECT 72.015 78.745 72.185 79.355 ;
        RECT 72.355 78.965 72.685 79.400 ;
        RECT 73.490 79.255 73.660 80.155 ;
        RECT 73.830 79.425 74.095 79.985 ;
        RECT 74.345 79.655 74.515 80.155 ;
        RECT 74.685 79.485 75.000 80.505 ;
        RECT 75.245 80.155 75.475 81.295 ;
        RECT 75.645 80.145 75.975 81.125 ;
        RECT 76.145 80.155 76.355 81.295 ;
        RECT 75.225 79.735 75.555 79.985 ;
        RECT 73.070 78.745 73.310 79.255 ;
        RECT 73.490 78.925 73.770 79.255 ;
        RECT 74.000 78.745 74.215 79.255 ;
        RECT 74.385 78.915 75.000 79.485 ;
        RECT 75.245 78.745 75.475 79.565 ;
        RECT 75.725 79.545 75.975 80.145 ;
        RECT 76.585 80.130 76.875 81.295 ;
        RECT 77.050 80.955 78.130 81.110 ;
        RECT 77.050 80.940 78.195 80.955 ;
        RECT 77.050 80.155 77.385 80.940 ;
        RECT 77.960 80.785 78.195 80.940 ;
        RECT 77.555 79.985 77.790 80.665 ;
        RECT 77.960 80.325 78.130 80.785 ;
        RECT 78.395 80.495 78.710 81.295 ;
        RECT 78.975 80.625 79.145 81.125 ;
        RECT 79.315 80.795 79.645 81.295 ;
        RECT 78.975 80.455 79.640 80.625 ;
        RECT 77.960 80.155 78.275 80.325 ;
        RECT 77.050 79.655 77.385 79.985 ;
        RECT 77.555 79.655 77.935 79.985 ;
        RECT 75.645 78.915 75.975 79.545 ;
        RECT 76.145 78.745 76.355 79.565 ;
        RECT 78.105 79.485 78.275 80.155 ;
        RECT 76.585 78.745 76.875 79.470 ;
        RECT 77.050 79.315 78.275 79.485 ;
        RECT 78.445 79.315 78.715 80.325 ;
        RECT 78.890 79.635 79.240 80.285 ;
        RECT 79.410 79.465 79.640 80.455 ;
        RECT 77.050 79.045 77.305 79.315 ;
        RECT 77.475 78.745 77.805 79.145 ;
        RECT 77.975 79.045 78.145 79.315 ;
        RECT 78.975 79.295 79.640 79.465 ;
        RECT 78.315 78.745 78.645 79.145 ;
        RECT 78.975 79.005 79.145 79.295 ;
        RECT 79.315 78.745 79.645 79.125 ;
        RECT 79.815 79.005 80.000 81.125 ;
        RECT 80.240 80.835 80.505 81.295 ;
        RECT 80.675 80.700 80.925 81.125 ;
        RECT 81.135 80.850 82.240 81.020 ;
        RECT 80.620 80.570 80.925 80.700 ;
        RECT 80.170 79.375 80.450 80.325 ;
        RECT 80.620 79.465 80.790 80.570 ;
        RECT 80.960 79.785 81.200 80.380 ;
        RECT 81.370 80.315 81.900 80.680 ;
        RECT 81.370 79.615 81.540 80.315 ;
        RECT 82.070 80.235 82.240 80.850 ;
        RECT 82.410 80.495 82.580 81.295 ;
        RECT 82.750 80.795 83.000 81.125 ;
        RECT 83.225 80.825 84.110 80.995 ;
        RECT 82.070 80.145 82.580 80.235 ;
        RECT 80.620 79.335 80.845 79.465 ;
        RECT 81.015 79.395 81.540 79.615 ;
        RECT 81.710 79.975 82.580 80.145 ;
        RECT 80.255 78.745 80.505 79.205 ;
        RECT 80.675 79.195 80.845 79.335 ;
        RECT 81.710 79.195 81.880 79.975 ;
        RECT 82.410 79.905 82.580 79.975 ;
        RECT 82.090 79.725 82.290 79.755 ;
        RECT 82.750 79.725 82.920 80.795 ;
        RECT 83.090 79.905 83.280 80.625 ;
        RECT 82.090 79.425 82.920 79.725 ;
        RECT 83.450 79.695 83.770 80.655 ;
        RECT 80.675 79.025 81.010 79.195 ;
        RECT 81.205 79.025 81.880 79.195 ;
        RECT 82.200 78.745 82.570 79.245 ;
        RECT 82.750 79.195 82.920 79.425 ;
        RECT 83.305 79.365 83.770 79.695 ;
        RECT 83.940 79.985 84.110 80.825 ;
        RECT 84.290 80.795 84.605 81.295 ;
        RECT 84.835 80.565 85.175 81.125 ;
        RECT 84.280 80.190 85.175 80.565 ;
        RECT 85.345 80.285 85.515 81.295 ;
        RECT 84.985 79.985 85.175 80.190 ;
        RECT 85.685 80.235 86.015 81.080 ;
        RECT 86.430 80.325 86.820 80.500 ;
        RECT 87.305 80.495 87.635 81.295 ;
        RECT 87.805 80.505 88.340 81.125 ;
        RECT 85.685 80.155 86.075 80.235 ;
        RECT 86.430 80.155 87.855 80.325 ;
        RECT 85.860 80.105 86.075 80.155 ;
        RECT 83.940 79.655 84.815 79.985 ;
        RECT 84.985 79.655 85.735 79.985 ;
        RECT 83.940 79.195 84.110 79.655 ;
        RECT 84.985 79.485 85.185 79.655 ;
        RECT 85.905 79.525 86.075 80.105 ;
        RECT 85.850 79.485 86.075 79.525 ;
        RECT 82.750 79.025 83.155 79.195 ;
        RECT 83.325 79.025 84.110 79.195 ;
        RECT 84.385 78.745 84.595 79.275 ;
        RECT 84.855 78.960 85.185 79.485 ;
        RECT 85.695 79.400 86.075 79.485 ;
        RECT 86.305 79.425 86.660 79.985 ;
        RECT 85.355 78.745 85.525 79.355 ;
        RECT 85.695 78.965 86.025 79.400 ;
        RECT 86.830 79.255 87.000 80.155 ;
        RECT 87.170 79.425 87.435 79.985 ;
        RECT 87.685 79.655 87.855 80.155 ;
        RECT 88.025 79.485 88.340 80.505 ;
        RECT 88.545 80.205 89.755 81.295 ;
        RECT 99.990 81.095 100.160 87.615 ;
        RECT 100.640 84.975 100.990 87.135 ;
        RECT 100.640 81.575 100.990 83.735 ;
        RECT 101.470 81.095 101.640 87.615 ;
        RECT 102.120 84.975 102.470 87.135 ;
        RECT 102.120 81.575 102.470 83.735 ;
        RECT 102.950 81.095 103.120 87.615 ;
        RECT 103.600 84.975 103.950 87.135 ;
        RECT 103.600 81.575 103.950 83.735 ;
        RECT 104.430 81.095 104.600 87.615 ;
        RECT 105.080 84.975 105.430 87.135 ;
        RECT 105.080 81.575 105.430 83.735 ;
        RECT 105.910 81.095 106.080 87.615 ;
        RECT 106.560 84.975 106.910 87.135 ;
        RECT 106.560 81.575 106.910 83.735 ;
        RECT 107.390 81.095 107.560 87.615 ;
        RECT 108.040 84.975 108.390 87.135 ;
        RECT 108.040 81.575 108.390 83.735 ;
        RECT 108.870 81.095 109.040 87.615 ;
        RECT 109.520 84.975 109.870 87.135 ;
        RECT 109.520 81.575 109.870 83.735 ;
        RECT 110.350 81.095 110.520 87.615 ;
        RECT 111.000 84.975 111.350 87.135 ;
        RECT 111.000 81.575 111.350 83.735 ;
        RECT 111.830 81.095 112.000 87.615 ;
        RECT 112.480 84.975 112.830 87.135 ;
        RECT 112.480 81.575 112.830 83.735 ;
        RECT 113.310 81.095 113.480 87.615 ;
        RECT 99.990 80.925 113.480 81.095 ;
        RECT 88.545 79.665 89.065 80.205 ;
        RECT 89.235 79.495 89.755 80.035 ;
        RECT 86.410 78.745 86.650 79.255 ;
        RECT 86.830 78.925 87.110 79.255 ;
        RECT 87.340 78.745 87.555 79.255 ;
        RECT 87.725 78.915 88.340 79.485 ;
        RECT 88.545 78.745 89.755 79.495 ;
        RECT 12.100 78.575 89.840 78.745 ;
        RECT 12.185 77.825 13.395 78.575 ;
        RECT 12.185 77.285 12.705 77.825 ;
        RECT 13.565 77.805 15.235 78.575 ;
        RECT 12.875 77.115 13.395 77.655 ;
        RECT 13.565 77.285 14.315 77.805 ;
        RECT 15.865 77.775 16.560 78.405 ;
        RECT 16.765 77.775 17.075 78.575 ;
        RECT 17.245 78.030 22.590 78.575 ;
        RECT 14.485 77.115 15.235 77.635 ;
        RECT 15.885 77.335 16.220 77.585 ;
        RECT 16.390 77.175 16.560 77.775 ;
        RECT 16.730 77.335 17.065 77.605 ;
        RECT 18.830 77.200 19.170 78.030 ;
        RECT 23.685 77.775 23.995 78.575 ;
        RECT 24.200 77.775 24.895 78.405 ;
        RECT 25.065 78.195 25.955 78.365 ;
        RECT 12.185 76.025 13.395 77.115 ;
        RECT 13.565 76.025 15.235 77.115 ;
        RECT 15.865 76.025 16.125 77.165 ;
        RECT 16.295 76.195 16.625 77.175 ;
        RECT 16.795 76.025 17.075 77.165 ;
        RECT 20.650 76.460 21.000 77.710 ;
        RECT 23.695 77.335 24.030 77.605 ;
        RECT 24.200 77.175 24.370 77.775 ;
        RECT 25.065 77.640 25.615 78.025 ;
        RECT 24.540 77.335 24.875 77.585 ;
        RECT 25.785 77.470 25.955 78.195 ;
        RECT 25.065 77.400 25.955 77.470 ;
        RECT 26.125 77.870 26.345 78.355 ;
        RECT 26.515 78.035 26.765 78.575 ;
        RECT 26.935 77.925 27.195 78.405 ;
        RECT 26.125 77.445 26.455 77.870 ;
        RECT 25.065 77.375 25.960 77.400 ;
        RECT 25.065 77.360 25.970 77.375 ;
        RECT 25.065 77.345 25.975 77.360 ;
        RECT 25.065 77.340 25.985 77.345 ;
        RECT 25.065 77.330 25.990 77.340 ;
        RECT 25.065 77.320 25.995 77.330 ;
        RECT 25.065 77.315 26.005 77.320 ;
        RECT 25.065 77.305 26.015 77.315 ;
        RECT 25.065 77.300 26.025 77.305 ;
        RECT 17.245 76.025 22.590 76.460 ;
        RECT 23.685 76.025 23.965 77.165 ;
        RECT 24.135 76.195 24.465 77.175 ;
        RECT 24.635 76.025 24.895 77.165 ;
        RECT 25.065 76.850 25.325 77.300 ;
        RECT 25.690 77.295 26.025 77.300 ;
        RECT 25.690 77.290 26.040 77.295 ;
        RECT 25.690 77.280 26.055 77.290 ;
        RECT 25.690 77.275 26.080 77.280 ;
        RECT 26.625 77.275 26.855 77.670 ;
        RECT 25.690 77.270 26.855 77.275 ;
        RECT 25.720 77.235 26.855 77.270 ;
        RECT 25.755 77.210 26.855 77.235 ;
        RECT 25.785 77.180 26.855 77.210 ;
        RECT 25.805 77.150 26.855 77.180 ;
        RECT 25.825 77.120 26.855 77.150 ;
        RECT 25.895 77.110 26.855 77.120 ;
        RECT 25.920 77.100 26.855 77.110 ;
        RECT 25.940 77.085 26.855 77.100 ;
        RECT 25.960 77.070 26.855 77.085 ;
        RECT 25.965 77.060 26.750 77.070 ;
        RECT 25.980 77.025 26.750 77.060 ;
        RECT 25.495 76.705 25.825 76.950 ;
        RECT 25.995 76.775 26.750 77.025 ;
        RECT 27.025 76.895 27.195 77.925 ;
        RECT 27.565 77.945 27.895 78.305 ;
        RECT 28.515 78.115 28.765 78.575 ;
        RECT 28.935 78.115 29.495 78.405 ;
        RECT 27.565 77.755 28.955 77.945 ;
        RECT 28.785 77.665 28.955 77.755 ;
        RECT 27.380 77.335 28.055 77.585 ;
        RECT 28.275 77.335 28.615 77.585 ;
        RECT 28.785 77.335 29.075 77.665 ;
        RECT 27.380 76.975 27.645 77.335 ;
        RECT 28.785 77.085 28.955 77.335 ;
        RECT 25.495 76.680 25.680 76.705 ;
        RECT 25.065 76.580 25.680 76.680 ;
        RECT 25.065 76.025 25.670 76.580 ;
        RECT 25.845 76.195 26.325 76.535 ;
        RECT 26.495 76.025 26.750 76.570 ;
        RECT 26.920 76.195 27.195 76.895 ;
        RECT 28.015 76.915 28.955 77.085 ;
        RECT 27.565 76.025 27.845 76.695 ;
        RECT 28.015 76.365 28.315 76.915 ;
        RECT 29.245 76.745 29.495 78.115 ;
        RECT 29.715 77.920 30.045 78.355 ;
        RECT 30.215 77.965 30.385 78.575 ;
        RECT 29.665 77.835 30.045 77.920 ;
        RECT 30.555 77.835 30.885 78.360 ;
        RECT 31.145 78.045 31.355 78.575 ;
        RECT 31.630 78.125 32.415 78.295 ;
        RECT 32.585 78.125 32.990 78.295 ;
        RECT 29.665 77.795 29.890 77.835 ;
        RECT 29.665 77.215 29.835 77.795 ;
        RECT 30.555 77.665 30.755 77.835 ;
        RECT 31.630 77.665 31.800 78.125 ;
        RECT 30.005 77.335 30.755 77.665 ;
        RECT 30.925 77.335 31.800 77.665 ;
        RECT 29.665 77.165 29.880 77.215 ;
        RECT 29.665 77.085 30.055 77.165 ;
        RECT 28.515 76.025 28.845 76.745 ;
        RECT 29.035 76.195 29.495 76.745 ;
        RECT 29.725 76.240 30.055 77.085 ;
        RECT 30.565 77.130 30.755 77.335 ;
        RECT 30.225 76.025 30.395 77.035 ;
        RECT 30.565 76.755 31.460 77.130 ;
        RECT 30.565 76.195 30.905 76.755 ;
        RECT 31.135 76.025 31.450 76.525 ;
        RECT 31.630 76.495 31.800 77.335 ;
        RECT 31.970 77.625 32.435 77.955 ;
        RECT 32.820 77.895 32.990 78.125 ;
        RECT 33.170 78.075 33.540 78.575 ;
        RECT 33.860 78.125 34.535 78.295 ;
        RECT 34.730 78.125 35.065 78.295 ;
        RECT 31.970 76.665 32.290 77.625 ;
        RECT 32.820 77.595 33.650 77.895 ;
        RECT 32.460 76.695 32.650 77.415 ;
        RECT 32.820 76.525 32.990 77.595 ;
        RECT 33.450 77.565 33.650 77.595 ;
        RECT 33.160 77.345 33.330 77.415 ;
        RECT 33.860 77.345 34.030 78.125 ;
        RECT 34.895 77.985 35.065 78.125 ;
        RECT 35.235 78.115 35.485 78.575 ;
        RECT 33.160 77.175 34.030 77.345 ;
        RECT 34.200 77.705 34.725 77.925 ;
        RECT 34.895 77.855 35.120 77.985 ;
        RECT 33.160 77.085 33.670 77.175 ;
        RECT 31.630 76.325 32.515 76.495 ;
        RECT 32.740 76.195 32.990 76.525 ;
        RECT 33.160 76.025 33.330 76.825 ;
        RECT 33.500 76.470 33.670 77.085 ;
        RECT 34.200 77.005 34.370 77.705 ;
        RECT 33.840 76.640 34.370 77.005 ;
        RECT 34.540 76.940 34.780 77.535 ;
        RECT 34.950 76.750 35.120 77.855 ;
        RECT 35.290 76.995 35.570 77.945 ;
        RECT 34.815 76.620 35.120 76.750 ;
        RECT 33.500 76.300 34.605 76.470 ;
        RECT 34.815 76.195 35.065 76.620 ;
        RECT 35.235 76.025 35.500 76.485 ;
        RECT 35.740 76.195 35.925 78.315 ;
        RECT 36.095 78.195 36.425 78.575 ;
        RECT 36.595 78.025 36.765 78.315 ;
        RECT 36.100 77.855 36.765 78.025 ;
        RECT 36.100 76.865 36.330 77.855 ;
        RECT 37.945 77.850 38.235 78.575 ;
        RECT 38.580 77.925 38.910 78.405 ;
        RECT 39.080 78.095 39.330 78.575 ;
        RECT 39.500 77.925 39.830 78.405 ;
        RECT 40.000 78.095 40.250 78.575 ;
        RECT 40.420 78.095 40.750 78.405 ;
        RECT 40.420 77.925 40.590 78.095 ;
        RECT 41.115 77.925 41.455 78.405 ;
        RECT 41.685 78.115 41.930 78.575 ;
        RECT 38.580 77.755 40.590 77.925 ;
        RECT 40.760 77.755 41.455 77.925 ;
        RECT 36.500 77.035 36.850 77.685 ;
        RECT 38.460 77.335 39.040 77.585 ;
        RECT 39.210 77.245 39.540 77.585 ;
        RECT 39.710 77.415 40.040 77.585 ;
        RECT 36.100 76.695 36.765 76.865 ;
        RECT 36.095 76.025 36.425 76.525 ;
        RECT 36.595 76.195 36.765 76.695 ;
        RECT 37.945 76.025 38.235 77.190 ;
        RECT 38.580 76.025 38.910 77.165 ;
        RECT 39.210 76.535 39.550 77.245 ;
        RECT 39.155 76.365 39.550 76.535 ;
        RECT 39.210 76.305 39.550 76.365 ;
        RECT 39.720 76.305 40.040 77.415 ;
        RECT 40.220 77.415 40.550 77.585 ;
        RECT 40.220 76.305 40.525 77.415 ;
        RECT 40.760 77.175 40.930 77.755 ;
        RECT 41.100 77.385 41.435 77.585 ;
        RECT 41.625 77.335 41.940 77.945 ;
        RECT 42.110 77.585 42.360 78.395 ;
        RECT 42.530 78.050 42.790 78.575 ;
        RECT 42.960 77.925 43.220 78.380 ;
        RECT 43.390 78.095 43.650 78.575 ;
        RECT 43.820 77.925 44.080 78.380 ;
        RECT 44.250 78.095 44.510 78.575 ;
        RECT 44.680 77.925 44.940 78.380 ;
        RECT 45.110 78.095 45.370 78.575 ;
        RECT 45.540 77.925 45.800 78.380 ;
        RECT 45.970 78.095 46.270 78.575 ;
        RECT 46.775 78.025 46.945 78.315 ;
        RECT 47.115 78.195 47.445 78.575 ;
        RECT 42.960 77.755 46.270 77.925 ;
        RECT 46.775 77.855 47.440 78.025 ;
        RECT 42.110 77.335 45.130 77.585 ;
        RECT 40.695 76.195 41.025 77.175 ;
        RECT 41.195 76.025 41.455 77.215 ;
        RECT 41.635 76.025 41.930 77.135 ;
        RECT 42.110 76.200 42.360 77.335 ;
        RECT 45.300 77.165 46.270 77.755 ;
        RECT 42.530 76.025 42.790 77.135 ;
        RECT 42.960 76.925 46.270 77.165 ;
        RECT 46.690 77.035 47.040 77.685 ;
        RECT 42.960 76.200 43.220 76.925 ;
        RECT 43.390 76.025 43.650 76.755 ;
        RECT 43.820 76.200 44.080 76.925 ;
        RECT 44.250 76.025 44.510 76.755 ;
        RECT 44.680 76.200 44.940 76.925 ;
        RECT 45.110 76.025 45.370 76.755 ;
        RECT 45.540 76.200 45.800 76.925 ;
        RECT 47.210 76.865 47.440 77.855 ;
        RECT 45.970 76.025 46.265 76.755 ;
        RECT 46.775 76.695 47.440 76.865 ;
        RECT 46.775 76.195 46.945 76.695 ;
        RECT 47.115 76.025 47.445 76.525 ;
        RECT 47.615 76.195 47.800 78.315 ;
        RECT 48.055 78.115 48.305 78.575 ;
        RECT 48.475 78.125 48.810 78.295 ;
        RECT 49.005 78.125 49.680 78.295 ;
        RECT 48.475 77.985 48.645 78.125 ;
        RECT 47.970 76.995 48.250 77.945 ;
        RECT 48.420 77.855 48.645 77.985 ;
        RECT 48.420 76.750 48.590 77.855 ;
        RECT 48.815 77.705 49.340 77.925 ;
        RECT 48.760 76.940 49.000 77.535 ;
        RECT 49.170 77.005 49.340 77.705 ;
        RECT 49.510 77.345 49.680 78.125 ;
        RECT 50.000 78.075 50.370 78.575 ;
        RECT 50.550 78.125 50.955 78.295 ;
        RECT 51.125 78.125 51.910 78.295 ;
        RECT 50.550 77.895 50.720 78.125 ;
        RECT 49.890 77.595 50.720 77.895 ;
        RECT 51.105 77.625 51.570 77.955 ;
        RECT 49.890 77.565 50.090 77.595 ;
        RECT 50.210 77.345 50.380 77.415 ;
        RECT 49.510 77.175 50.380 77.345 ;
        RECT 49.870 77.085 50.380 77.175 ;
        RECT 48.420 76.620 48.725 76.750 ;
        RECT 49.170 76.640 49.700 77.005 ;
        RECT 48.040 76.025 48.305 76.485 ;
        RECT 48.475 76.195 48.725 76.620 ;
        RECT 49.870 76.470 50.040 77.085 ;
        RECT 48.935 76.300 50.040 76.470 ;
        RECT 50.210 76.025 50.380 76.825 ;
        RECT 50.550 76.525 50.720 77.595 ;
        RECT 50.890 76.695 51.080 77.415 ;
        RECT 51.250 76.665 51.570 77.625 ;
        RECT 51.740 77.665 51.910 78.125 ;
        RECT 52.185 78.045 52.395 78.575 ;
        RECT 52.655 77.835 52.985 78.360 ;
        RECT 53.155 77.965 53.325 78.575 ;
        RECT 53.495 77.920 53.825 78.355 ;
        RECT 53.495 77.835 53.875 77.920 ;
        RECT 52.785 77.665 52.985 77.835 ;
        RECT 53.650 77.795 53.875 77.835 ;
        RECT 51.740 77.335 52.615 77.665 ;
        RECT 52.785 77.335 53.535 77.665 ;
        RECT 50.550 76.195 50.800 76.525 ;
        RECT 51.740 76.495 51.910 77.335 ;
        RECT 52.785 77.130 52.975 77.335 ;
        RECT 53.705 77.215 53.875 77.795 ;
        RECT 54.045 77.825 55.255 78.575 ;
        RECT 55.460 77.835 56.075 78.405 ;
        RECT 56.245 78.065 56.460 78.575 ;
        RECT 56.690 78.065 56.970 78.395 ;
        RECT 57.150 78.065 57.390 78.575 ;
        RECT 54.045 77.285 54.565 77.825 ;
        RECT 53.660 77.165 53.875 77.215 ;
        RECT 52.080 76.755 52.975 77.130 ;
        RECT 53.485 77.085 53.875 77.165 ;
        RECT 54.735 77.115 55.255 77.655 ;
        RECT 51.025 76.325 51.910 76.495 ;
        RECT 52.090 76.025 52.405 76.525 ;
        RECT 52.635 76.195 52.975 76.755 ;
        RECT 53.145 76.025 53.315 77.035 ;
        RECT 53.485 76.240 53.815 77.085 ;
        RECT 54.045 76.025 55.255 77.115 ;
        RECT 55.460 76.815 55.775 77.835 ;
        RECT 55.945 77.165 56.115 77.665 ;
        RECT 56.365 77.335 56.630 77.895 ;
        RECT 56.800 77.165 56.970 78.065 ;
        RECT 58.845 77.945 59.175 78.305 ;
        RECT 59.795 78.115 60.045 78.575 ;
        RECT 60.215 78.115 60.775 78.405 ;
        RECT 57.140 77.335 57.495 77.895 ;
        RECT 58.845 77.755 60.235 77.945 ;
        RECT 60.065 77.665 60.235 77.755 ;
        RECT 58.660 77.335 59.335 77.585 ;
        RECT 59.555 77.335 59.895 77.585 ;
        RECT 60.065 77.335 60.355 77.665 ;
        RECT 55.945 76.995 57.370 77.165 ;
        RECT 55.460 76.195 55.995 76.815 ;
        RECT 56.165 76.025 56.495 76.825 ;
        RECT 56.980 76.820 57.370 76.995 ;
        RECT 58.660 76.975 58.925 77.335 ;
        RECT 60.065 77.085 60.235 77.335 ;
        RECT 59.295 76.915 60.235 77.085 ;
        RECT 58.845 76.025 59.125 76.695 ;
        RECT 59.295 76.365 59.595 76.915 ;
        RECT 60.525 76.745 60.775 78.115 ;
        RECT 59.795 76.025 60.125 76.745 ;
        RECT 60.315 76.195 60.775 76.745 ;
        RECT 60.945 78.075 61.245 78.405 ;
        RECT 61.415 78.095 61.690 78.575 ;
        RECT 60.945 77.165 61.115 78.075 ;
        RECT 61.870 77.925 62.165 78.315 ;
        RECT 62.335 78.095 62.590 78.575 ;
        RECT 62.765 77.925 63.025 78.315 ;
        RECT 63.195 78.095 63.475 78.575 ;
        RECT 61.285 77.335 61.635 77.905 ;
        RECT 61.870 77.755 63.520 77.925 ;
        RECT 63.705 77.850 63.995 78.575 ;
        RECT 64.280 77.945 64.565 78.405 ;
        RECT 64.735 78.115 65.005 78.575 ;
        RECT 64.280 77.775 65.235 77.945 ;
        RECT 61.805 77.415 62.945 77.585 ;
        RECT 61.805 77.165 61.975 77.415 ;
        RECT 63.115 77.245 63.520 77.755 ;
        RECT 60.945 76.995 61.975 77.165 ;
        RECT 62.765 77.075 63.520 77.245 ;
        RECT 60.945 76.195 61.255 76.995 ;
        RECT 62.765 76.825 63.025 77.075 ;
        RECT 61.425 76.025 61.735 76.825 ;
        RECT 61.905 76.655 63.025 76.825 ;
        RECT 61.905 76.195 62.165 76.655 ;
        RECT 62.335 76.025 62.590 76.485 ;
        RECT 62.765 76.195 63.025 76.655 ;
        RECT 63.195 76.025 63.480 76.895 ;
        RECT 63.705 76.025 63.995 77.190 ;
        RECT 64.165 77.045 64.855 77.605 ;
        RECT 65.025 76.875 65.235 77.775 ;
        RECT 64.280 76.655 65.235 76.875 ;
        RECT 65.405 77.605 65.805 78.405 ;
        RECT 65.995 77.945 66.275 78.405 ;
        RECT 66.795 78.115 67.120 78.575 ;
        RECT 65.995 77.775 67.120 77.945 ;
        RECT 67.290 77.835 67.675 78.405 ;
        RECT 66.670 77.665 67.120 77.775 ;
        RECT 65.405 77.045 66.500 77.605 ;
        RECT 66.670 77.335 67.225 77.665 ;
        RECT 64.280 76.195 64.565 76.655 ;
        RECT 64.735 76.025 65.005 76.485 ;
        RECT 65.405 76.195 65.805 77.045 ;
        RECT 66.670 76.875 67.120 77.335 ;
        RECT 67.395 77.165 67.675 77.835 ;
        RECT 65.995 76.655 67.120 76.875 ;
        RECT 65.995 76.195 66.275 76.655 ;
        RECT 66.795 76.025 67.120 76.485 ;
        RECT 67.290 76.195 67.675 77.165 ;
        RECT 68.310 77.835 68.565 78.405 ;
        RECT 68.735 78.175 69.065 78.575 ;
        RECT 69.490 78.040 70.020 78.405 ;
        RECT 69.490 78.005 69.665 78.040 ;
        RECT 68.735 77.835 69.665 78.005 ;
        RECT 68.310 77.165 68.480 77.835 ;
        RECT 68.735 77.665 68.905 77.835 ;
        RECT 68.650 77.335 68.905 77.665 ;
        RECT 69.130 77.335 69.325 77.665 ;
        RECT 68.310 76.195 68.645 77.165 ;
        RECT 68.815 76.025 68.985 77.165 ;
        RECT 69.155 76.365 69.325 77.335 ;
        RECT 69.495 76.705 69.665 77.835 ;
        RECT 69.835 77.045 70.005 77.845 ;
        RECT 70.210 77.555 70.485 78.405 ;
        RECT 70.205 77.385 70.485 77.555 ;
        RECT 70.210 77.245 70.485 77.385 ;
        RECT 70.655 77.045 70.845 78.405 ;
        RECT 71.025 78.040 71.535 78.575 ;
        RECT 71.755 77.765 72.000 78.370 ;
        RECT 72.445 77.835 72.830 78.405 ;
        RECT 73.000 78.115 73.325 78.575 ;
        RECT 73.845 77.945 74.125 78.405 ;
        RECT 71.045 77.595 72.275 77.765 ;
        RECT 69.835 76.875 70.845 77.045 ;
        RECT 71.015 77.030 71.765 77.220 ;
        RECT 69.495 76.535 70.620 76.705 ;
        RECT 71.015 76.365 71.185 77.030 ;
        RECT 71.935 76.785 72.275 77.595 ;
        RECT 69.155 76.195 71.185 76.365 ;
        RECT 71.355 76.025 71.525 76.785 ;
        RECT 71.760 76.375 72.275 76.785 ;
        RECT 72.445 77.165 72.725 77.835 ;
        RECT 73.000 77.775 74.125 77.945 ;
        RECT 73.000 77.665 73.450 77.775 ;
        RECT 72.895 77.335 73.450 77.665 ;
        RECT 74.315 77.605 74.715 78.405 ;
        RECT 75.115 78.115 75.385 78.575 ;
        RECT 75.555 77.945 75.840 78.405 ;
        RECT 76.195 78.175 76.525 78.575 ;
        RECT 76.695 78.005 76.865 78.275 ;
        RECT 77.035 78.175 77.365 78.575 ;
        RECT 77.535 78.005 77.790 78.275 ;
        RECT 72.445 76.195 72.830 77.165 ;
        RECT 73.000 76.875 73.450 77.335 ;
        RECT 73.620 77.045 74.715 77.605 ;
        RECT 73.000 76.655 74.125 76.875 ;
        RECT 73.000 76.025 73.325 76.485 ;
        RECT 73.845 76.195 74.125 76.655 ;
        RECT 74.315 76.195 74.715 77.045 ;
        RECT 74.885 77.775 75.840 77.945 ;
        RECT 74.885 76.875 75.095 77.775 ;
        RECT 75.265 77.045 75.955 77.605 ;
        RECT 76.125 76.995 76.395 78.005 ;
        RECT 76.565 77.835 77.790 78.005 ;
        RECT 78.055 78.025 78.225 78.405 ;
        RECT 78.405 78.195 78.735 78.575 ;
        RECT 78.055 77.855 78.720 78.025 ;
        RECT 78.915 77.900 79.175 78.405 ;
        RECT 76.565 77.165 76.735 77.835 ;
        RECT 76.905 77.335 77.285 77.665 ;
        RECT 77.455 77.335 77.790 77.665 ;
        RECT 76.565 76.995 76.880 77.165 ;
        RECT 74.885 76.655 75.840 76.875 ;
        RECT 75.115 76.025 75.385 76.485 ;
        RECT 75.555 76.195 75.840 76.655 ;
        RECT 76.130 76.025 76.445 76.825 ;
        RECT 76.710 76.380 76.880 76.995 ;
        RECT 77.050 76.655 77.285 77.335 ;
        RECT 77.985 77.305 78.315 77.675 ;
        RECT 78.550 77.600 78.720 77.855 ;
        RECT 78.550 77.270 78.835 77.600 ;
        RECT 77.455 76.380 77.790 77.165 ;
        RECT 78.550 77.125 78.720 77.270 ;
        RECT 76.710 76.210 77.790 76.380 ;
        RECT 78.055 76.955 78.720 77.125 ;
        RECT 79.005 77.100 79.175 77.900 ;
        RECT 79.435 78.025 79.605 78.315 ;
        RECT 79.775 78.195 80.105 78.575 ;
        RECT 79.435 77.855 80.100 78.025 ;
        RECT 78.055 76.195 78.225 76.955 ;
        RECT 78.405 76.025 78.735 76.785 ;
        RECT 78.905 76.195 79.175 77.100 ;
        RECT 79.350 77.035 79.700 77.685 ;
        RECT 79.870 76.865 80.100 77.855 ;
        RECT 79.435 76.695 80.100 76.865 ;
        RECT 79.435 76.195 79.605 76.695 ;
        RECT 79.775 76.025 80.105 76.525 ;
        RECT 80.275 76.195 80.460 78.315 ;
        RECT 80.715 78.115 80.965 78.575 ;
        RECT 81.135 78.125 81.470 78.295 ;
        RECT 81.665 78.125 82.340 78.295 ;
        RECT 81.135 77.985 81.305 78.125 ;
        RECT 80.630 76.995 80.910 77.945 ;
        RECT 81.080 77.855 81.305 77.985 ;
        RECT 81.080 76.750 81.250 77.855 ;
        RECT 81.475 77.705 82.000 77.925 ;
        RECT 81.420 76.940 81.660 77.535 ;
        RECT 81.830 77.005 82.000 77.705 ;
        RECT 82.170 77.345 82.340 78.125 ;
        RECT 82.660 78.075 83.030 78.575 ;
        RECT 83.210 78.125 83.615 78.295 ;
        RECT 83.785 78.125 84.570 78.295 ;
        RECT 83.210 77.895 83.380 78.125 ;
        RECT 82.550 77.595 83.380 77.895 ;
        RECT 83.765 77.625 84.230 77.955 ;
        RECT 82.550 77.565 82.750 77.595 ;
        RECT 82.870 77.345 83.040 77.415 ;
        RECT 82.170 77.175 83.040 77.345 ;
        RECT 82.530 77.085 83.040 77.175 ;
        RECT 81.080 76.620 81.385 76.750 ;
        RECT 81.830 76.640 82.360 77.005 ;
        RECT 80.700 76.025 80.965 76.485 ;
        RECT 81.135 76.195 81.385 76.620 ;
        RECT 82.530 76.470 82.700 77.085 ;
        RECT 81.595 76.300 82.700 76.470 ;
        RECT 82.870 76.025 83.040 76.825 ;
        RECT 83.210 76.525 83.380 77.595 ;
        RECT 83.550 76.695 83.740 77.415 ;
        RECT 83.910 76.665 84.230 77.625 ;
        RECT 84.400 77.665 84.570 78.125 ;
        RECT 84.845 78.045 85.055 78.575 ;
        RECT 85.315 77.835 85.645 78.360 ;
        RECT 85.815 77.965 85.985 78.575 ;
        RECT 86.155 77.920 86.485 78.355 ;
        RECT 86.795 78.025 86.965 78.405 ;
        RECT 87.180 78.195 87.510 78.575 ;
        RECT 86.155 77.835 86.535 77.920 ;
        RECT 86.795 77.855 87.510 78.025 ;
        RECT 85.445 77.665 85.645 77.835 ;
        RECT 86.310 77.795 86.535 77.835 ;
        RECT 84.400 77.335 85.275 77.665 ;
        RECT 85.445 77.335 86.195 77.665 ;
        RECT 83.210 76.195 83.460 76.525 ;
        RECT 84.400 76.495 84.570 77.335 ;
        RECT 85.445 77.130 85.635 77.335 ;
        RECT 86.365 77.215 86.535 77.795 ;
        RECT 86.705 77.305 87.060 77.675 ;
        RECT 87.340 77.665 87.510 77.855 ;
        RECT 87.680 77.830 87.935 78.405 ;
        RECT 87.340 77.335 87.595 77.665 ;
        RECT 86.320 77.165 86.535 77.215 ;
        RECT 84.740 76.755 85.635 77.130 ;
        RECT 86.145 77.085 86.535 77.165 ;
        RECT 87.340 77.125 87.510 77.335 ;
        RECT 83.685 76.325 84.570 76.495 ;
        RECT 84.750 76.025 85.065 76.525 ;
        RECT 85.295 76.195 85.635 76.755 ;
        RECT 85.805 76.025 85.975 77.035 ;
        RECT 86.145 76.240 86.475 77.085 ;
        RECT 86.795 76.955 87.510 77.125 ;
        RECT 87.765 77.100 87.935 77.830 ;
        RECT 88.110 77.735 88.370 78.575 ;
        RECT 88.545 77.825 89.755 78.575 ;
        RECT 86.795 76.195 86.965 76.955 ;
        RECT 87.180 76.025 87.510 76.785 ;
        RECT 87.680 76.195 87.935 77.100 ;
        RECT 88.110 76.025 88.370 77.175 ;
        RECT 88.545 77.115 89.065 77.655 ;
        RECT 89.235 77.285 89.755 77.825 ;
        RECT 88.545 76.025 89.755 77.115 ;
        RECT 12.100 75.855 89.840 76.025 ;
        RECT 12.185 74.765 13.395 75.855 ;
        RECT 13.655 75.185 13.825 75.685 ;
        RECT 13.995 75.355 14.325 75.855 ;
        RECT 13.655 75.015 14.320 75.185 ;
        RECT 12.185 74.055 12.705 74.595 ;
        RECT 12.875 74.225 13.395 74.765 ;
        RECT 13.570 74.195 13.920 74.845 ;
        RECT 12.185 73.305 13.395 74.055 ;
        RECT 14.090 74.025 14.320 75.015 ;
        RECT 13.655 73.855 14.320 74.025 ;
        RECT 13.655 73.565 13.825 73.855 ;
        RECT 13.995 73.305 14.325 73.685 ;
        RECT 14.495 73.565 14.680 75.685 ;
        RECT 14.920 75.395 15.185 75.855 ;
        RECT 15.355 75.260 15.605 75.685 ;
        RECT 15.815 75.410 16.920 75.580 ;
        RECT 15.300 75.130 15.605 75.260 ;
        RECT 14.850 73.935 15.130 74.885 ;
        RECT 15.300 74.025 15.470 75.130 ;
        RECT 15.640 74.345 15.880 74.940 ;
        RECT 16.050 74.875 16.580 75.240 ;
        RECT 16.050 74.175 16.220 74.875 ;
        RECT 16.750 74.795 16.920 75.410 ;
        RECT 17.090 75.055 17.260 75.855 ;
        RECT 17.430 75.355 17.680 75.685 ;
        RECT 17.905 75.385 18.790 75.555 ;
        RECT 16.750 74.705 17.260 74.795 ;
        RECT 15.300 73.895 15.525 74.025 ;
        RECT 15.695 73.955 16.220 74.175 ;
        RECT 16.390 74.535 17.260 74.705 ;
        RECT 14.935 73.305 15.185 73.765 ;
        RECT 15.355 73.755 15.525 73.895 ;
        RECT 16.390 73.755 16.560 74.535 ;
        RECT 17.090 74.465 17.260 74.535 ;
        RECT 16.770 74.285 16.970 74.315 ;
        RECT 17.430 74.285 17.600 75.355 ;
        RECT 17.770 74.465 17.960 75.185 ;
        RECT 16.770 73.985 17.600 74.285 ;
        RECT 18.130 74.255 18.450 75.215 ;
        RECT 15.355 73.585 15.690 73.755 ;
        RECT 15.885 73.585 16.560 73.755 ;
        RECT 16.880 73.305 17.250 73.805 ;
        RECT 17.430 73.755 17.600 73.985 ;
        RECT 17.985 73.925 18.450 74.255 ;
        RECT 18.620 74.545 18.790 75.385 ;
        RECT 18.970 75.355 19.285 75.855 ;
        RECT 19.515 75.125 19.855 75.685 ;
        RECT 18.960 74.750 19.855 75.125 ;
        RECT 20.025 74.845 20.195 75.855 ;
        RECT 19.665 74.545 19.855 74.750 ;
        RECT 20.365 74.795 20.695 75.640 ;
        RECT 21.395 75.245 21.725 75.675 ;
        RECT 21.905 75.415 22.100 75.855 ;
        RECT 22.270 75.245 22.600 75.675 ;
        RECT 21.395 75.075 22.600 75.245 ;
        RECT 20.365 74.715 20.755 74.795 ;
        RECT 21.395 74.745 22.290 75.075 ;
        RECT 22.770 74.905 23.045 75.675 ;
        RECT 23.230 75.055 23.485 75.855 ;
        RECT 23.685 75.005 24.015 75.685 ;
        RECT 20.540 74.665 20.755 74.715 ;
        RECT 18.620 74.215 19.495 74.545 ;
        RECT 19.665 74.215 20.415 74.545 ;
        RECT 18.620 73.755 18.790 74.215 ;
        RECT 19.665 74.045 19.865 74.215 ;
        RECT 20.585 74.085 20.755 74.665 ;
        RECT 22.460 74.715 23.045 74.905 ;
        RECT 21.400 74.215 21.695 74.545 ;
        RECT 21.875 74.215 22.290 74.545 ;
        RECT 20.530 74.045 20.755 74.085 ;
        RECT 17.430 73.585 17.835 73.755 ;
        RECT 18.005 73.585 18.790 73.755 ;
        RECT 19.065 73.305 19.275 73.835 ;
        RECT 19.535 73.520 19.865 74.045 ;
        RECT 20.375 73.960 20.755 74.045 ;
        RECT 20.035 73.305 20.205 73.915 ;
        RECT 20.375 73.525 20.705 73.960 ;
        RECT 21.395 73.305 21.695 74.035 ;
        RECT 21.875 73.595 22.105 74.215 ;
        RECT 22.460 74.045 22.635 74.715 ;
        RECT 22.305 73.865 22.635 74.045 ;
        RECT 22.805 73.895 23.045 74.545 ;
        RECT 23.230 74.515 23.475 74.875 ;
        RECT 23.665 74.725 24.015 75.005 ;
        RECT 23.665 74.345 23.835 74.725 ;
        RECT 24.195 74.545 24.390 75.595 ;
        RECT 24.570 74.715 24.890 75.855 ;
        RECT 25.065 74.690 25.355 75.855 ;
        RECT 25.525 74.885 25.815 75.685 ;
        RECT 25.985 75.055 26.220 75.855 ;
        RECT 26.405 75.515 27.940 75.685 ;
        RECT 26.405 74.885 26.735 75.515 ;
        RECT 25.525 74.715 26.735 74.885 ;
        RECT 23.315 74.175 23.835 74.345 ;
        RECT 24.005 74.215 24.390 74.545 ;
        RECT 24.570 74.495 24.830 74.545 ;
        RECT 24.570 74.325 24.835 74.495 ;
        RECT 24.570 74.215 24.830 74.325 ;
        RECT 25.525 74.215 25.770 74.545 ;
        RECT 23.315 74.155 23.485 74.175 ;
        RECT 23.285 73.985 23.485 74.155 ;
        RECT 25.940 74.045 26.110 74.715 ;
        RECT 26.905 74.545 27.140 75.290 ;
        RECT 26.280 74.215 26.680 74.545 ;
        RECT 26.850 74.215 27.140 74.545 ;
        RECT 27.330 74.545 27.600 75.290 ;
        RECT 27.770 74.885 27.940 75.515 ;
        RECT 28.110 75.055 28.515 75.855 ;
        RECT 27.770 74.715 28.515 74.885 ;
        RECT 27.330 74.215 27.670 74.545 ;
        RECT 27.840 74.215 28.175 74.545 ;
        RECT 28.345 74.215 28.515 74.715 ;
        RECT 28.685 74.290 29.035 75.685 ;
        RECT 29.675 74.745 29.970 75.855 ;
        RECT 30.150 74.545 30.400 75.680 ;
        RECT 30.570 74.745 30.830 75.855 ;
        RECT 31.000 74.955 31.260 75.680 ;
        RECT 31.430 75.125 31.690 75.855 ;
        RECT 31.860 74.955 32.120 75.680 ;
        RECT 32.290 75.125 32.550 75.855 ;
        RECT 32.720 74.955 32.980 75.680 ;
        RECT 33.150 75.125 33.410 75.855 ;
        RECT 33.580 74.955 33.840 75.680 ;
        RECT 34.010 75.125 34.305 75.855 ;
        RECT 31.000 74.715 34.310 74.955 ;
        RECT 34.725 74.765 36.395 75.855 ;
        RECT 37.140 75.225 37.425 75.685 ;
        RECT 37.595 75.395 37.865 75.855 ;
        RECT 37.140 75.005 38.095 75.225 ;
        RECT 22.305 73.485 22.530 73.865 ;
        RECT 22.700 73.305 23.030 73.695 ;
        RECT 23.315 73.610 23.485 73.985 ;
        RECT 23.675 73.835 24.890 74.005 ;
        RECT 23.675 73.530 23.905 73.835 ;
        RECT 24.075 73.305 24.405 73.665 ;
        RECT 24.600 73.485 24.890 73.835 ;
        RECT 25.065 73.305 25.355 74.030 ;
        RECT 25.525 73.475 26.110 74.045 ;
        RECT 26.360 73.875 27.755 74.045 ;
        RECT 26.360 73.530 26.690 73.875 ;
        RECT 26.905 73.305 27.280 73.705 ;
        RECT 27.460 73.530 27.755 73.875 ;
        RECT 27.925 73.305 28.595 74.045 ;
        RECT 28.765 73.475 29.035 74.290 ;
        RECT 29.665 73.935 29.980 74.545 ;
        RECT 30.150 74.295 33.170 74.545 ;
        RECT 29.725 73.305 29.970 73.765 ;
        RECT 30.150 73.485 30.400 74.295 ;
        RECT 33.340 74.125 34.310 74.715 ;
        RECT 31.000 73.955 34.310 74.125 ;
        RECT 34.725 74.075 35.475 74.595 ;
        RECT 35.645 74.245 36.395 74.765 ;
        RECT 37.025 74.275 37.715 74.835 ;
        RECT 37.885 74.105 38.095 75.005 ;
        RECT 30.570 73.305 30.830 73.830 ;
        RECT 31.000 73.500 31.260 73.955 ;
        RECT 31.430 73.305 31.690 73.785 ;
        RECT 31.860 73.500 32.120 73.955 ;
        RECT 32.290 73.305 32.550 73.785 ;
        RECT 32.720 73.500 32.980 73.955 ;
        RECT 33.150 73.305 33.410 73.785 ;
        RECT 33.580 73.500 33.840 73.955 ;
        RECT 34.010 73.305 34.310 73.785 ;
        RECT 34.725 73.305 36.395 74.075 ;
        RECT 37.140 73.935 38.095 74.105 ;
        RECT 38.265 74.835 38.665 75.685 ;
        RECT 38.855 75.225 39.135 75.685 ;
        RECT 39.655 75.395 39.980 75.855 ;
        RECT 38.855 75.005 39.980 75.225 ;
        RECT 38.265 74.275 39.360 74.835 ;
        RECT 39.530 74.545 39.980 75.005 ;
        RECT 40.150 74.715 40.535 75.685 ;
        RECT 40.705 74.780 41.045 75.855 ;
        RECT 41.230 75.345 43.280 75.635 ;
        RECT 37.140 73.475 37.425 73.935 ;
        RECT 37.595 73.305 37.865 73.765 ;
        RECT 38.265 73.475 38.665 74.275 ;
        RECT 39.530 74.215 40.085 74.545 ;
        RECT 39.530 74.105 39.980 74.215 ;
        RECT 38.855 73.935 39.980 74.105 ;
        RECT 40.255 74.045 40.535 74.715 ;
        RECT 41.215 74.545 41.455 75.140 ;
        RECT 41.650 75.005 43.280 75.175 ;
        RECT 43.450 75.055 43.730 75.855 ;
        RECT 41.650 74.715 41.970 75.005 ;
        RECT 43.110 74.885 43.280 75.005 ;
        RECT 38.855 73.475 39.135 73.935 ;
        RECT 39.655 73.305 39.980 73.765 ;
        RECT 40.150 73.475 40.535 74.045 ;
        RECT 40.705 73.975 41.045 74.545 ;
        RECT 41.215 74.215 41.870 74.545 ;
        RECT 42.140 74.215 42.880 74.835 ;
        RECT 43.110 74.715 43.770 74.885 ;
        RECT 43.940 74.715 44.215 75.685 ;
        RECT 44.385 74.765 45.595 75.855 ;
        RECT 43.600 74.545 43.770 74.715 ;
        RECT 43.050 74.215 43.430 74.545 ;
        RECT 43.600 74.215 43.875 74.545 ;
        RECT 40.705 73.305 41.045 73.805 ;
        RECT 41.215 73.525 41.460 74.215 ;
        RECT 43.600 74.045 43.770 74.215 ;
        RECT 42.185 73.875 43.770 74.045 ;
        RECT 44.045 73.980 44.215 74.715 ;
        RECT 41.655 73.305 41.985 73.805 ;
        RECT 42.185 73.525 42.355 73.875 ;
        RECT 42.530 73.305 42.860 73.705 ;
        RECT 43.030 73.525 43.200 73.875 ;
        RECT 43.370 73.305 43.750 73.705 ;
        RECT 43.940 73.635 44.215 73.980 ;
        RECT 44.385 74.055 44.905 74.595 ;
        RECT 45.075 74.225 45.595 74.765 ;
        RECT 45.765 74.715 46.150 75.685 ;
        RECT 46.320 75.395 46.645 75.855 ;
        RECT 47.165 75.225 47.445 75.685 ;
        RECT 46.320 75.005 47.445 75.225 ;
        RECT 44.385 73.305 45.595 74.055 ;
        RECT 45.765 74.045 46.045 74.715 ;
        RECT 46.320 74.545 46.770 75.005 ;
        RECT 47.635 74.835 48.035 75.685 ;
        RECT 48.435 75.395 48.705 75.855 ;
        RECT 48.875 75.225 49.160 75.685 ;
        RECT 46.215 74.215 46.770 74.545 ;
        RECT 46.940 74.275 48.035 74.835 ;
        RECT 46.320 74.105 46.770 74.215 ;
        RECT 45.765 73.475 46.150 74.045 ;
        RECT 46.320 73.935 47.445 74.105 ;
        RECT 46.320 73.305 46.645 73.765 ;
        RECT 47.165 73.475 47.445 73.935 ;
        RECT 47.635 73.475 48.035 74.275 ;
        RECT 48.205 75.005 49.160 75.225 ;
        RECT 48.205 74.105 48.415 75.005 ;
        RECT 48.585 74.275 49.275 74.835 ;
        RECT 49.445 74.765 50.655 75.855 ;
        RECT 48.205 73.935 49.160 74.105 ;
        RECT 48.435 73.305 48.705 73.765 ;
        RECT 48.875 73.475 49.160 73.935 ;
        RECT 49.445 74.055 49.965 74.595 ;
        RECT 50.135 74.225 50.655 74.765 ;
        RECT 50.825 74.690 51.115 75.855 ;
        RECT 51.285 74.765 54.795 75.855 ;
        RECT 51.285 74.075 52.935 74.595 ;
        RECT 53.105 74.245 54.795 74.765 ;
        RECT 55.975 74.925 56.145 75.685 ;
        RECT 56.360 75.095 56.690 75.855 ;
        RECT 55.975 74.755 56.690 74.925 ;
        RECT 56.860 74.780 57.115 75.685 ;
        RECT 55.885 74.205 56.240 74.575 ;
        RECT 56.520 74.545 56.690 74.755 ;
        RECT 56.520 74.215 56.775 74.545 ;
        RECT 49.445 73.305 50.655 74.055 ;
        RECT 50.825 73.305 51.115 74.030 ;
        RECT 51.285 73.305 54.795 74.075 ;
        RECT 56.520 74.025 56.690 74.215 ;
        RECT 56.945 74.050 57.115 74.780 ;
        RECT 57.290 74.705 57.550 75.855 ;
        RECT 57.735 74.885 58.065 75.685 ;
        RECT 58.235 75.055 58.465 75.855 ;
        RECT 58.635 74.885 58.965 75.685 ;
        RECT 57.735 74.715 58.965 74.885 ;
        RECT 59.135 74.715 59.390 75.855 ;
        RECT 59.680 75.225 59.965 75.685 ;
        RECT 60.135 75.395 60.405 75.855 ;
        RECT 59.680 75.005 60.635 75.225 ;
        RECT 57.725 74.215 58.035 74.545 ;
        RECT 55.975 73.855 56.690 74.025 ;
        RECT 55.975 73.475 56.145 73.855 ;
        RECT 56.360 73.305 56.690 73.685 ;
        RECT 56.860 73.475 57.115 74.050 ;
        RECT 57.290 73.305 57.550 74.145 ;
        RECT 57.735 73.815 58.065 74.045 ;
        RECT 58.240 73.985 58.615 74.545 ;
        RECT 58.785 73.815 58.965 74.715 ;
        RECT 59.150 73.965 59.370 74.545 ;
        RECT 59.565 74.275 60.255 74.835 ;
        RECT 60.425 74.105 60.635 75.005 ;
        RECT 57.735 73.475 58.965 73.815 ;
        RECT 59.680 73.935 60.635 74.105 ;
        RECT 60.805 74.835 61.205 75.685 ;
        RECT 61.395 75.225 61.675 75.685 ;
        RECT 62.195 75.395 62.520 75.855 ;
        RECT 61.395 75.005 62.520 75.225 ;
        RECT 60.805 74.275 61.900 74.835 ;
        RECT 62.070 74.545 62.520 75.005 ;
        RECT 62.690 74.715 63.075 75.685 ;
        RECT 59.135 73.305 59.390 73.795 ;
        RECT 59.680 73.475 59.965 73.935 ;
        RECT 60.135 73.305 60.405 73.765 ;
        RECT 60.805 73.475 61.205 74.275 ;
        RECT 62.070 74.215 62.625 74.545 ;
        RECT 62.070 74.105 62.520 74.215 ;
        RECT 61.395 73.935 62.520 74.105 ;
        RECT 62.795 74.045 63.075 74.715 ;
        RECT 63.250 75.465 63.585 75.685 ;
        RECT 64.590 75.475 64.945 75.855 ;
        RECT 63.250 74.845 63.505 75.465 ;
        RECT 63.755 75.305 63.985 75.345 ;
        RECT 65.115 75.305 65.365 75.685 ;
        RECT 63.755 75.105 65.365 75.305 ;
        RECT 63.755 75.015 63.940 75.105 ;
        RECT 64.530 75.095 65.365 75.105 ;
        RECT 65.615 75.075 65.865 75.855 ;
        RECT 66.035 75.005 66.295 75.685 ;
        RECT 66.555 75.185 66.725 75.685 ;
        RECT 66.895 75.355 67.225 75.855 ;
        RECT 66.555 75.015 67.220 75.185 ;
        RECT 64.095 74.905 64.425 74.935 ;
        RECT 64.095 74.845 65.895 74.905 ;
        RECT 63.250 74.735 65.955 74.845 ;
        RECT 63.250 74.675 64.425 74.735 ;
        RECT 65.755 74.700 65.955 74.735 ;
        RECT 63.245 74.295 63.735 74.495 ;
        RECT 63.925 74.295 64.400 74.505 ;
        RECT 61.395 73.475 61.675 73.935 ;
        RECT 62.195 73.305 62.520 73.765 ;
        RECT 62.690 73.475 63.075 74.045 ;
        RECT 63.250 73.305 63.705 74.070 ;
        RECT 64.180 73.895 64.400 74.295 ;
        RECT 64.645 74.295 64.975 74.505 ;
        RECT 64.645 73.895 64.855 74.295 ;
        RECT 65.145 74.260 65.555 74.565 ;
        RECT 65.785 74.125 65.955 74.700 ;
        RECT 65.685 74.005 65.955 74.125 ;
        RECT 65.110 73.960 65.955 74.005 ;
        RECT 65.110 73.835 65.865 73.960 ;
        RECT 65.110 73.685 65.280 73.835 ;
        RECT 66.125 73.815 66.295 75.005 ;
        RECT 66.470 74.195 66.820 74.845 ;
        RECT 66.990 74.025 67.220 75.015 ;
        RECT 66.065 73.805 66.295 73.815 ;
        RECT 63.980 73.475 65.280 73.685 ;
        RECT 65.535 73.305 65.865 73.665 ;
        RECT 66.035 73.475 66.295 73.805 ;
        RECT 66.555 73.855 67.220 74.025 ;
        RECT 66.555 73.565 66.725 73.855 ;
        RECT 66.895 73.305 67.225 73.685 ;
        RECT 67.395 73.565 67.580 75.685 ;
        RECT 67.820 75.395 68.085 75.855 ;
        RECT 68.255 75.260 68.505 75.685 ;
        RECT 68.715 75.410 69.820 75.580 ;
        RECT 68.200 75.130 68.505 75.260 ;
        RECT 67.750 73.935 68.030 74.885 ;
        RECT 68.200 74.025 68.370 75.130 ;
        RECT 68.540 74.345 68.780 74.940 ;
        RECT 68.950 74.875 69.480 75.240 ;
        RECT 68.950 74.175 69.120 74.875 ;
        RECT 69.650 74.795 69.820 75.410 ;
        RECT 69.990 75.055 70.160 75.855 ;
        RECT 70.330 75.355 70.580 75.685 ;
        RECT 70.805 75.385 71.690 75.555 ;
        RECT 69.650 74.705 70.160 74.795 ;
        RECT 68.200 73.895 68.425 74.025 ;
        RECT 68.595 73.955 69.120 74.175 ;
        RECT 69.290 74.535 70.160 74.705 ;
        RECT 67.835 73.305 68.085 73.765 ;
        RECT 68.255 73.755 68.425 73.895 ;
        RECT 69.290 73.755 69.460 74.535 ;
        RECT 69.990 74.465 70.160 74.535 ;
        RECT 69.670 74.285 69.870 74.315 ;
        RECT 70.330 74.285 70.500 75.355 ;
        RECT 70.670 74.465 70.860 75.185 ;
        RECT 69.670 73.985 70.500 74.285 ;
        RECT 71.030 74.255 71.350 75.215 ;
        RECT 68.255 73.585 68.590 73.755 ;
        RECT 68.785 73.585 69.460 73.755 ;
        RECT 69.780 73.305 70.150 73.805 ;
        RECT 70.330 73.755 70.500 73.985 ;
        RECT 70.885 73.925 71.350 74.255 ;
        RECT 71.520 74.545 71.690 75.385 ;
        RECT 71.870 75.355 72.185 75.855 ;
        RECT 72.415 75.125 72.755 75.685 ;
        RECT 71.860 74.750 72.755 75.125 ;
        RECT 72.925 74.845 73.095 75.855 ;
        RECT 72.565 74.545 72.755 74.750 ;
        RECT 73.265 74.795 73.595 75.640 ;
        RECT 73.265 74.715 73.655 74.795 ;
        RECT 73.440 74.665 73.655 74.715 ;
        RECT 74.750 74.705 75.010 75.855 ;
        RECT 75.185 74.780 75.440 75.685 ;
        RECT 75.610 75.095 75.940 75.855 ;
        RECT 76.155 74.925 76.325 75.685 ;
        RECT 71.520 74.215 72.395 74.545 ;
        RECT 72.565 74.215 73.315 74.545 ;
        RECT 71.520 73.755 71.690 74.215 ;
        RECT 72.565 74.045 72.765 74.215 ;
        RECT 73.485 74.085 73.655 74.665 ;
        RECT 73.430 74.045 73.655 74.085 ;
        RECT 70.330 73.585 70.735 73.755 ;
        RECT 70.905 73.585 71.690 73.755 ;
        RECT 71.965 73.305 72.175 73.835 ;
        RECT 72.435 73.520 72.765 74.045 ;
        RECT 73.275 73.960 73.655 74.045 ;
        RECT 72.935 73.305 73.105 73.915 ;
        RECT 73.275 73.525 73.605 73.960 ;
        RECT 74.750 73.305 75.010 74.145 ;
        RECT 75.185 74.050 75.355 74.780 ;
        RECT 75.610 74.755 76.325 74.925 ;
        RECT 75.610 74.545 75.780 74.755 ;
        RECT 76.585 74.690 76.875 75.855 ;
        RECT 77.045 74.715 77.430 75.685 ;
        RECT 77.600 75.395 77.925 75.855 ;
        RECT 78.445 75.225 78.725 75.685 ;
        RECT 77.600 75.005 78.725 75.225 ;
        RECT 75.525 74.215 75.780 74.545 ;
        RECT 75.185 73.475 75.440 74.050 ;
        RECT 75.610 74.025 75.780 74.215 ;
        RECT 76.060 74.205 76.415 74.575 ;
        RECT 77.045 74.045 77.325 74.715 ;
        RECT 77.600 74.545 78.050 75.005 ;
        RECT 78.915 74.835 79.315 75.685 ;
        RECT 79.715 75.395 79.985 75.855 ;
        RECT 80.155 75.225 80.440 75.685 ;
        RECT 80.730 75.430 81.065 75.855 ;
        RECT 81.235 75.250 81.420 75.655 ;
        RECT 77.495 74.215 78.050 74.545 ;
        RECT 78.220 74.275 79.315 74.835 ;
        RECT 77.600 74.105 78.050 74.215 ;
        RECT 75.610 73.855 76.325 74.025 ;
        RECT 75.610 73.305 75.940 73.685 ;
        RECT 76.155 73.475 76.325 73.855 ;
        RECT 76.585 73.305 76.875 74.030 ;
        RECT 77.045 73.475 77.430 74.045 ;
        RECT 77.600 73.935 78.725 74.105 ;
        RECT 77.600 73.305 77.925 73.765 ;
        RECT 78.445 73.475 78.725 73.935 ;
        RECT 78.915 73.475 79.315 74.275 ;
        RECT 79.485 75.005 80.440 75.225 ;
        RECT 80.755 75.075 81.420 75.250 ;
        RECT 81.625 75.075 81.955 75.855 ;
        RECT 79.485 74.105 79.695 75.005 ;
        RECT 79.865 74.275 80.555 74.835 ;
        RECT 79.485 73.935 80.440 74.105 ;
        RECT 79.715 73.305 79.985 73.765 ;
        RECT 80.155 73.475 80.440 73.935 ;
        RECT 80.755 74.045 81.095 75.075 ;
        RECT 82.125 74.885 82.395 75.655 ;
        RECT 81.265 74.715 82.395 74.885 ;
        RECT 82.655 74.925 82.825 75.685 ;
        RECT 83.040 75.095 83.370 75.855 ;
        RECT 82.655 74.755 83.370 74.925 ;
        RECT 83.540 74.780 83.795 75.685 ;
        RECT 81.265 74.215 81.515 74.715 ;
        RECT 80.755 73.875 81.440 74.045 ;
        RECT 81.695 73.965 82.055 74.545 ;
        RECT 80.730 73.305 81.065 73.705 ;
        RECT 81.235 73.475 81.440 73.875 ;
        RECT 82.225 73.805 82.395 74.715 ;
        RECT 82.565 74.205 82.920 74.575 ;
        RECT 83.200 74.545 83.370 74.755 ;
        RECT 83.200 74.215 83.455 74.545 ;
        RECT 83.200 74.025 83.370 74.215 ;
        RECT 83.625 74.050 83.795 74.780 ;
        RECT 83.970 74.705 84.230 75.855 ;
        RECT 84.405 75.005 84.665 75.685 ;
        RECT 84.835 75.075 85.085 75.855 ;
        RECT 85.335 75.305 85.585 75.685 ;
        RECT 85.755 75.475 86.110 75.855 ;
        RECT 87.115 75.465 87.450 75.685 ;
        RECT 86.715 75.305 86.945 75.345 ;
        RECT 85.335 75.105 86.945 75.305 ;
        RECT 85.335 75.095 86.170 75.105 ;
        RECT 86.760 75.015 86.945 75.105 ;
        RECT 81.650 73.305 81.925 73.785 ;
        RECT 82.135 73.475 82.395 73.805 ;
        RECT 82.655 73.855 83.370 74.025 ;
        RECT 82.655 73.475 82.825 73.855 ;
        RECT 83.040 73.305 83.370 73.685 ;
        RECT 83.540 73.475 83.795 74.050 ;
        RECT 83.970 73.305 84.230 74.145 ;
        RECT 84.405 73.805 84.575 75.005 ;
        RECT 86.275 74.905 86.605 74.935 ;
        RECT 84.805 74.845 86.605 74.905 ;
        RECT 87.195 74.845 87.450 75.465 ;
        RECT 84.745 74.735 87.450 74.845 ;
        RECT 84.745 74.700 84.945 74.735 ;
        RECT 84.745 74.125 84.915 74.700 ;
        RECT 86.275 74.675 87.450 74.735 ;
        RECT 88.545 74.765 89.755 75.855 ;
        RECT 99.990 75.105 100.160 80.925 ;
        RECT 100.640 78.285 100.990 80.445 ;
        RECT 100.640 75.585 100.990 77.745 ;
        RECT 101.470 75.105 101.640 80.925 ;
        RECT 102.120 78.285 102.470 80.445 ;
        RECT 102.120 75.585 102.470 77.745 ;
        RECT 102.950 75.105 103.120 80.925 ;
        RECT 103.600 78.285 103.950 80.445 ;
        RECT 103.600 75.585 103.950 77.745 ;
        RECT 104.430 75.105 104.600 80.925 ;
        RECT 105.080 78.285 105.430 80.445 ;
        RECT 105.080 75.585 105.430 77.745 ;
        RECT 105.910 75.105 106.080 80.925 ;
        RECT 106.560 78.285 106.910 80.445 ;
        RECT 106.560 75.585 106.910 77.745 ;
        RECT 107.390 75.105 107.560 80.925 ;
        RECT 108.040 78.285 108.390 80.445 ;
        RECT 108.040 75.585 108.390 77.745 ;
        RECT 108.870 75.105 109.040 80.925 ;
        RECT 109.520 78.285 109.870 80.445 ;
        RECT 109.520 75.585 109.870 77.745 ;
        RECT 110.350 75.105 110.520 80.925 ;
        RECT 99.990 74.935 110.520 75.105 ;
        RECT 85.145 74.260 85.555 74.565 ;
        RECT 85.725 74.295 86.055 74.505 ;
        RECT 84.745 74.005 85.015 74.125 ;
        RECT 84.745 73.960 85.590 74.005 ;
        RECT 84.835 73.835 85.590 73.960 ;
        RECT 85.845 73.895 86.055 74.295 ;
        RECT 86.300 74.295 86.775 74.505 ;
        RECT 86.965 74.295 87.455 74.495 ;
        RECT 86.300 73.895 86.520 74.295 ;
        RECT 88.545 74.225 89.065 74.765 ;
        RECT 84.405 73.475 84.665 73.805 ;
        RECT 85.420 73.685 85.590 73.835 ;
        RECT 84.835 73.305 85.165 73.665 ;
        RECT 85.420 73.475 86.720 73.685 ;
        RECT 86.995 73.305 87.450 74.070 ;
        RECT 89.235 74.055 89.755 74.595 ;
        RECT 88.545 73.305 89.755 74.055 ;
        RECT 12.100 73.135 89.840 73.305 ;
        RECT 12.185 72.385 13.395 73.135 ;
        RECT 14.485 72.415 14.825 72.925 ;
        RECT 12.185 71.845 12.705 72.385 ;
        RECT 12.875 71.675 13.395 72.215 ;
        RECT 12.185 70.585 13.395 71.675 ;
        RECT 14.485 71.015 14.745 72.415 ;
        RECT 14.995 72.335 15.265 73.135 ;
        RECT 14.920 71.895 15.250 72.145 ;
        RECT 15.445 71.895 15.725 72.865 ;
        RECT 15.905 71.895 16.205 72.865 ;
        RECT 16.385 71.895 16.735 72.860 ;
        RECT 16.955 72.635 17.450 72.965 ;
        RECT 14.935 71.725 15.250 71.895 ;
        RECT 16.955 71.725 17.125 72.635 ;
        RECT 14.935 71.555 17.125 71.725 ;
        RECT 14.485 70.755 14.825 71.015 ;
        RECT 14.995 70.585 15.325 71.385 ;
        RECT 15.790 70.755 16.040 71.555 ;
        RECT 16.225 70.585 16.555 71.305 ;
        RECT 16.775 70.755 17.025 71.555 ;
        RECT 17.295 71.145 17.535 72.455 ;
        RECT 17.740 72.395 18.355 72.965 ;
        RECT 18.525 72.625 18.740 73.135 ;
        RECT 18.970 72.625 19.250 72.955 ;
        RECT 19.430 72.625 19.670 73.135 ;
        RECT 17.740 71.375 18.055 72.395 ;
        RECT 18.225 71.725 18.395 72.225 ;
        RECT 18.645 71.895 18.910 72.455 ;
        RECT 19.080 71.725 19.250 72.625 ;
        RECT 19.420 71.895 19.775 72.455 ;
        RECT 20.015 72.405 20.315 73.135 ;
        RECT 20.495 72.225 20.725 72.845 ;
        RECT 20.925 72.575 21.150 72.955 ;
        RECT 21.320 72.745 21.650 73.135 ;
        RECT 20.925 72.395 21.255 72.575 ;
        RECT 20.020 71.895 20.315 72.225 ;
        RECT 20.495 71.895 20.910 72.225 ;
        RECT 21.080 71.725 21.255 72.395 ;
        RECT 21.425 71.895 21.665 72.545 ;
        RECT 22.045 72.505 22.375 72.865 ;
        RECT 22.995 72.675 23.245 73.135 ;
        RECT 23.415 72.675 23.975 72.965 ;
        RECT 22.045 72.315 23.435 72.505 ;
        RECT 23.265 72.225 23.435 72.315 ;
        RECT 21.860 71.895 22.535 72.145 ;
        RECT 22.755 71.895 23.095 72.145 ;
        RECT 23.265 71.895 23.555 72.225 ;
        RECT 18.225 71.555 19.650 71.725 ;
        RECT 17.195 70.585 17.530 70.965 ;
        RECT 17.740 70.755 18.275 71.375 ;
        RECT 18.445 70.585 18.775 71.385 ;
        RECT 19.260 71.380 19.650 71.555 ;
        RECT 20.015 71.365 20.910 71.695 ;
        RECT 21.080 71.535 21.665 71.725 ;
        RECT 21.860 71.535 22.125 71.895 ;
        RECT 23.265 71.645 23.435 71.895 ;
        RECT 20.015 71.195 21.220 71.365 ;
        RECT 20.015 70.765 20.345 71.195 ;
        RECT 20.525 70.585 20.720 71.025 ;
        RECT 20.890 70.765 21.220 71.195 ;
        RECT 21.390 70.765 21.665 71.535 ;
        RECT 22.495 71.475 23.435 71.645 ;
        RECT 22.045 70.585 22.325 71.255 ;
        RECT 22.495 70.925 22.795 71.475 ;
        RECT 23.725 71.305 23.975 72.675 ;
        RECT 22.995 70.585 23.325 71.305 ;
        RECT 23.515 70.755 23.975 71.305 ;
        RECT 24.145 72.550 24.455 72.965 ;
        RECT 24.650 72.755 24.980 73.135 ;
        RECT 25.150 72.795 26.555 72.965 ;
        RECT 25.150 72.565 25.320 72.795 ;
        RECT 24.145 71.435 24.315 72.550 ;
        RECT 24.625 72.395 25.320 72.565 ;
        RECT 26.385 72.565 26.555 72.795 ;
        RECT 26.825 72.735 27.155 73.135 ;
        RECT 27.395 72.565 27.565 72.965 ;
        RECT 24.625 72.225 24.795 72.395 ;
        RECT 24.485 71.895 24.795 72.225 ;
        RECT 24.965 71.895 25.300 72.225 ;
        RECT 25.570 71.895 25.765 72.470 ;
        RECT 26.025 72.225 26.215 72.455 ;
        RECT 26.385 72.395 27.565 72.565 ;
        RECT 28.745 72.315 29.005 73.135 ;
        RECT 29.175 72.315 29.505 72.735 ;
        RECT 29.685 72.650 30.475 72.915 ;
        RECT 29.255 72.225 29.505 72.315 ;
        RECT 26.025 71.895 26.370 72.225 ;
        RECT 26.680 71.895 27.155 72.225 ;
        RECT 27.410 71.895 27.595 72.225 ;
        RECT 24.625 71.725 24.795 71.895 ;
        RECT 24.625 71.555 27.565 71.725 ;
        RECT 24.145 70.795 24.485 71.435 ;
        RECT 25.075 71.215 26.635 71.385 ;
        RECT 24.655 70.585 24.900 71.045 ;
        RECT 25.075 70.755 25.325 71.215 ;
        RECT 25.515 70.585 26.185 70.965 ;
        RECT 26.385 70.755 26.635 71.215 ;
        RECT 27.395 70.755 27.565 71.555 ;
        RECT 28.745 71.265 29.085 72.145 ;
        RECT 29.255 71.975 30.050 72.225 ;
        RECT 28.745 70.585 29.005 71.095 ;
        RECT 29.255 70.755 29.425 71.975 ;
        RECT 30.220 71.795 30.475 72.650 ;
        RECT 30.645 72.495 30.845 72.915 ;
        RECT 31.035 72.675 31.365 73.135 ;
        RECT 30.645 71.975 31.055 72.495 ;
        RECT 31.535 72.485 31.795 72.965 ;
        RECT 31.225 71.795 31.455 72.225 ;
        RECT 29.665 71.625 31.455 71.795 ;
        RECT 29.665 71.260 29.915 71.625 ;
        RECT 30.085 71.265 30.415 71.455 ;
        RECT 30.635 71.330 31.350 71.625 ;
        RECT 31.625 71.455 31.795 72.485 ;
        RECT 32.125 72.575 32.455 72.965 ;
        RECT 32.625 72.745 33.810 72.915 ;
        RECT 34.070 72.665 34.240 73.135 ;
        RECT 32.125 72.395 32.635 72.575 ;
        RECT 31.965 71.935 32.295 72.225 ;
        RECT 32.465 71.765 32.635 72.395 ;
        RECT 33.040 72.485 33.425 72.575 ;
        RECT 34.410 72.485 34.740 72.950 ;
        RECT 33.040 72.315 34.740 72.485 ;
        RECT 34.910 72.315 35.080 73.135 ;
        RECT 35.250 72.315 35.935 72.955 ;
        RECT 36.565 72.335 36.875 73.135 ;
        RECT 37.080 72.335 37.775 72.965 ;
        RECT 37.945 72.410 38.235 73.135 ;
        RECT 32.805 71.935 33.135 72.145 ;
        RECT 33.315 71.895 33.695 72.145 ;
        RECT 30.085 71.090 30.280 71.265 ;
        RECT 29.665 70.585 30.280 71.090 ;
        RECT 30.450 70.755 30.925 71.095 ;
        RECT 31.095 70.585 31.310 71.130 ;
        RECT 31.520 70.755 31.795 71.455 ;
        RECT 32.120 71.595 33.205 71.765 ;
        RECT 32.120 70.755 32.420 71.595 ;
        RECT 32.615 70.585 32.865 71.425 ;
        RECT 33.035 71.345 33.205 71.595 ;
        RECT 33.375 71.515 33.695 71.895 ;
        RECT 33.885 71.935 34.370 72.145 ;
        RECT 34.560 71.935 35.010 72.145 ;
        RECT 35.180 71.935 35.515 72.145 ;
        RECT 33.885 71.775 34.260 71.935 ;
        RECT 33.865 71.605 34.260 71.775 ;
        RECT 35.180 71.765 35.350 71.935 ;
        RECT 33.885 71.515 34.260 71.605 ;
        RECT 34.430 71.595 35.350 71.765 ;
        RECT 34.430 71.345 34.600 71.595 ;
        RECT 33.035 71.175 34.600 71.345 ;
        RECT 33.455 70.755 34.260 71.175 ;
        RECT 34.770 70.585 35.100 71.425 ;
        RECT 35.685 71.345 35.935 72.315 ;
        RECT 36.575 71.895 36.910 72.165 ;
        RECT 37.080 71.775 37.250 72.335 ;
        RECT 38.465 72.315 38.675 73.135 ;
        RECT 38.845 72.335 39.175 72.965 ;
        RECT 37.420 71.895 37.755 72.145 ;
        RECT 37.080 71.735 37.255 71.775 ;
        RECT 35.270 70.755 35.935 71.345 ;
        RECT 36.565 70.585 36.845 71.725 ;
        RECT 37.015 70.755 37.345 71.735 ;
        RECT 37.515 70.585 37.775 71.725 ;
        RECT 37.945 70.585 38.235 71.750 ;
        RECT 38.845 71.735 39.095 72.335 ;
        RECT 39.345 72.315 39.575 73.135 ;
        RECT 39.835 72.480 40.165 72.915 ;
        RECT 40.335 72.525 40.505 73.135 ;
        RECT 39.785 72.395 40.165 72.480 ;
        RECT 40.675 72.395 41.005 72.920 ;
        RECT 41.265 72.605 41.475 73.135 ;
        RECT 41.750 72.685 42.535 72.855 ;
        RECT 42.705 72.685 43.110 72.855 ;
        RECT 39.785 72.355 40.010 72.395 ;
        RECT 39.265 71.895 39.595 72.145 ;
        RECT 39.785 71.775 39.955 72.355 ;
        RECT 40.675 72.225 40.875 72.395 ;
        RECT 41.750 72.225 41.920 72.685 ;
        RECT 40.125 71.895 40.875 72.225 ;
        RECT 41.045 71.895 41.920 72.225 ;
        RECT 38.465 70.585 38.675 71.725 ;
        RECT 38.845 70.755 39.175 71.735 ;
        RECT 39.785 71.725 40.000 71.775 ;
        RECT 39.345 70.585 39.575 71.725 ;
        RECT 39.785 71.645 40.175 71.725 ;
        RECT 39.845 70.800 40.175 71.645 ;
        RECT 40.685 71.690 40.875 71.895 ;
        RECT 40.345 70.585 40.515 71.595 ;
        RECT 40.685 71.315 41.580 71.690 ;
        RECT 40.685 70.755 41.025 71.315 ;
        RECT 41.255 70.585 41.570 71.085 ;
        RECT 41.750 71.055 41.920 71.895 ;
        RECT 42.090 72.185 42.555 72.515 ;
        RECT 42.940 72.455 43.110 72.685 ;
        RECT 43.290 72.635 43.660 73.135 ;
        RECT 43.980 72.685 44.655 72.855 ;
        RECT 44.850 72.685 45.185 72.855 ;
        RECT 42.090 71.225 42.410 72.185 ;
        RECT 42.940 72.155 43.770 72.455 ;
        RECT 42.580 71.255 42.770 71.975 ;
        RECT 42.940 71.085 43.110 72.155 ;
        RECT 43.570 72.125 43.770 72.155 ;
        RECT 43.280 71.905 43.450 71.975 ;
        RECT 43.980 71.905 44.150 72.685 ;
        RECT 45.015 72.545 45.185 72.685 ;
        RECT 45.355 72.675 45.605 73.135 ;
        RECT 43.280 71.735 44.150 71.905 ;
        RECT 44.320 72.265 44.845 72.485 ;
        RECT 45.015 72.415 45.240 72.545 ;
        RECT 43.280 71.645 43.790 71.735 ;
        RECT 41.750 70.885 42.635 71.055 ;
        RECT 42.860 70.755 43.110 71.085 ;
        RECT 43.280 70.585 43.450 71.385 ;
        RECT 43.620 71.030 43.790 71.645 ;
        RECT 44.320 71.565 44.490 72.265 ;
        RECT 43.960 71.200 44.490 71.565 ;
        RECT 44.660 71.500 44.900 72.095 ;
        RECT 45.070 71.310 45.240 72.415 ;
        RECT 45.410 71.555 45.690 72.505 ;
        RECT 44.935 71.180 45.240 71.310 ;
        RECT 43.620 70.860 44.725 71.030 ;
        RECT 44.935 70.755 45.185 71.180 ;
        RECT 45.355 70.585 45.620 71.045 ;
        RECT 45.860 70.755 46.045 72.875 ;
        RECT 46.215 72.755 46.545 73.135 ;
        RECT 46.715 72.585 46.885 72.875 ;
        RECT 46.220 72.415 46.885 72.585 ;
        RECT 46.220 71.425 46.450 72.415 ;
        RECT 47.165 72.405 47.495 73.135 ;
        RECT 46.620 71.595 46.970 72.245 ;
        RECT 47.665 72.225 47.875 72.845 ;
        RECT 48.055 72.425 48.485 72.955 ;
        RECT 47.180 71.875 47.470 72.225 ;
        RECT 47.665 71.875 48.060 72.225 ;
        RECT 48.240 72.175 48.485 72.425 ;
        RECT 48.665 72.355 48.895 73.135 ;
        RECT 49.075 72.505 49.455 72.955 ;
        RECT 48.240 71.875 48.775 72.175 ;
        RECT 49.075 72.055 49.305 72.505 ;
        RECT 49.910 72.395 50.165 72.965 ;
        RECT 50.335 72.735 50.665 73.135 ;
        RECT 51.090 72.600 51.620 72.965 ;
        RECT 51.090 72.565 51.265 72.600 ;
        RECT 50.335 72.395 51.265 72.565 ;
        RECT 47.235 71.495 48.275 71.695 ;
        RECT 46.220 71.255 46.885 71.425 ;
        RECT 46.215 70.585 46.545 71.085 ;
        RECT 46.715 70.755 46.885 71.255 ;
        RECT 47.235 70.765 47.405 71.495 ;
        RECT 47.585 70.585 47.915 71.315 ;
        RECT 48.085 70.765 48.275 71.495 ;
        RECT 48.445 70.765 48.775 71.875 ;
        RECT 48.965 71.375 49.305 72.055 ;
        RECT 49.485 71.555 49.715 72.245 ;
        RECT 49.910 71.725 50.080 72.395 ;
        RECT 50.335 72.225 50.505 72.395 ;
        RECT 50.250 71.895 50.505 72.225 ;
        RECT 50.730 71.895 50.925 72.225 ;
        RECT 48.965 71.175 49.725 71.375 ;
        RECT 48.965 70.585 49.295 70.995 ;
        RECT 49.465 70.785 49.725 71.175 ;
        RECT 49.910 70.755 50.245 71.725 ;
        RECT 50.415 70.585 50.585 71.725 ;
        RECT 50.755 70.925 50.925 71.895 ;
        RECT 51.095 71.265 51.265 72.395 ;
        RECT 51.435 71.605 51.605 72.405 ;
        RECT 51.810 72.115 52.085 72.965 ;
        RECT 51.805 71.945 52.085 72.115 ;
        RECT 51.810 71.805 52.085 71.945 ;
        RECT 52.255 71.605 52.445 72.965 ;
        RECT 52.625 72.600 53.135 73.135 ;
        RECT 53.355 72.325 53.600 72.930 ;
        RECT 54.045 72.395 54.430 72.965 ;
        RECT 54.600 72.675 54.925 73.135 ;
        RECT 55.445 72.505 55.725 72.965 ;
        RECT 52.645 72.155 53.875 72.325 ;
        RECT 51.435 71.435 52.445 71.605 ;
        RECT 52.615 71.590 53.365 71.780 ;
        RECT 51.095 71.095 52.220 71.265 ;
        RECT 52.615 70.925 52.785 71.590 ;
        RECT 53.535 71.345 53.875 72.155 ;
        RECT 50.755 70.755 52.785 70.925 ;
        RECT 52.955 70.585 53.125 71.345 ;
        RECT 53.360 70.935 53.875 71.345 ;
        RECT 54.045 71.725 54.325 72.395 ;
        RECT 54.600 72.335 55.725 72.505 ;
        RECT 54.600 72.225 55.050 72.335 ;
        RECT 54.495 71.895 55.050 72.225 ;
        RECT 55.915 72.165 56.315 72.965 ;
        RECT 56.715 72.675 56.985 73.135 ;
        RECT 57.155 72.505 57.440 72.965 ;
        RECT 54.045 70.755 54.430 71.725 ;
        RECT 54.600 71.435 55.050 71.895 ;
        RECT 55.220 71.605 56.315 72.165 ;
        RECT 54.600 71.215 55.725 71.435 ;
        RECT 54.600 70.585 54.925 71.045 ;
        RECT 55.445 70.755 55.725 71.215 ;
        RECT 55.915 70.755 56.315 71.605 ;
        RECT 56.485 72.335 57.440 72.505 ;
        RECT 58.650 72.395 58.905 72.965 ;
        RECT 59.075 72.735 59.405 73.135 ;
        RECT 59.830 72.600 60.360 72.965 ;
        RECT 59.830 72.565 60.005 72.600 ;
        RECT 59.075 72.395 60.005 72.565 ;
        RECT 60.550 72.455 60.825 72.965 ;
        RECT 56.485 71.435 56.695 72.335 ;
        RECT 56.865 71.605 57.555 72.165 ;
        RECT 58.650 71.725 58.820 72.395 ;
        RECT 59.075 72.225 59.245 72.395 ;
        RECT 58.990 71.895 59.245 72.225 ;
        RECT 59.470 71.895 59.665 72.225 ;
        RECT 56.485 71.215 57.440 71.435 ;
        RECT 56.715 70.585 56.985 71.045 ;
        RECT 57.155 70.755 57.440 71.215 ;
        RECT 58.650 70.755 58.985 71.725 ;
        RECT 59.155 70.585 59.325 71.725 ;
        RECT 59.495 70.925 59.665 71.895 ;
        RECT 59.835 71.265 60.005 72.395 ;
        RECT 60.175 71.605 60.345 72.405 ;
        RECT 60.545 72.285 60.825 72.455 ;
        RECT 60.550 71.805 60.825 72.285 ;
        RECT 60.995 71.605 61.185 72.965 ;
        RECT 61.365 72.600 61.875 73.135 ;
        RECT 62.095 72.325 62.340 72.930 ;
        RECT 63.705 72.410 63.995 73.135 ;
        RECT 64.170 72.395 64.425 72.965 ;
        RECT 64.595 72.735 64.925 73.135 ;
        RECT 65.350 72.600 65.880 72.965 ;
        RECT 66.070 72.795 66.345 72.965 ;
        RECT 66.065 72.625 66.345 72.795 ;
        RECT 65.350 72.565 65.525 72.600 ;
        RECT 64.595 72.395 65.525 72.565 ;
        RECT 61.385 72.155 62.615 72.325 ;
        RECT 60.175 71.435 61.185 71.605 ;
        RECT 61.355 71.590 62.105 71.780 ;
        RECT 59.835 71.095 60.960 71.265 ;
        RECT 61.355 70.925 61.525 71.590 ;
        RECT 62.275 71.345 62.615 72.155 ;
        RECT 59.495 70.755 61.525 70.925 ;
        RECT 61.695 70.585 61.865 71.345 ;
        RECT 62.100 70.935 62.615 71.345 ;
        RECT 63.705 70.585 63.995 71.750 ;
        RECT 64.170 71.725 64.340 72.395 ;
        RECT 64.595 72.225 64.765 72.395 ;
        RECT 64.510 71.895 64.765 72.225 ;
        RECT 64.990 71.895 65.185 72.225 ;
        RECT 64.170 70.755 64.505 71.725 ;
        RECT 64.675 70.585 64.845 71.725 ;
        RECT 65.015 70.925 65.185 71.895 ;
        RECT 65.355 71.265 65.525 72.395 ;
        RECT 65.695 71.605 65.865 72.405 ;
        RECT 66.070 71.805 66.345 72.625 ;
        RECT 66.515 71.605 66.705 72.965 ;
        RECT 66.885 72.600 67.395 73.135 ;
        RECT 67.615 72.325 67.860 72.930 ;
        RECT 68.770 72.395 69.025 72.965 ;
        RECT 69.195 72.735 69.525 73.135 ;
        RECT 69.950 72.600 70.480 72.965 ;
        RECT 70.670 72.795 70.945 72.965 ;
        RECT 70.665 72.625 70.945 72.795 ;
        RECT 69.950 72.565 70.125 72.600 ;
        RECT 69.195 72.395 70.125 72.565 ;
        RECT 66.905 72.155 68.135 72.325 ;
        RECT 65.695 71.435 66.705 71.605 ;
        RECT 66.875 71.590 67.625 71.780 ;
        RECT 65.355 71.095 66.480 71.265 ;
        RECT 66.875 70.925 67.045 71.590 ;
        RECT 67.795 71.345 68.135 72.155 ;
        RECT 65.015 70.755 67.045 70.925 ;
        RECT 67.215 70.585 67.385 71.345 ;
        RECT 67.620 70.935 68.135 71.345 ;
        RECT 68.770 71.725 68.940 72.395 ;
        RECT 69.195 72.225 69.365 72.395 ;
        RECT 69.110 71.895 69.365 72.225 ;
        RECT 69.590 71.895 69.785 72.225 ;
        RECT 68.770 70.755 69.105 71.725 ;
        RECT 69.275 70.585 69.445 71.725 ;
        RECT 69.615 70.925 69.785 71.895 ;
        RECT 69.955 71.265 70.125 72.395 ;
        RECT 70.295 71.605 70.465 72.405 ;
        RECT 70.670 71.805 70.945 72.625 ;
        RECT 71.115 71.605 71.305 72.965 ;
        RECT 71.485 72.600 71.995 73.135 ;
        RECT 72.215 72.325 72.460 72.930 ;
        RECT 72.910 72.395 73.165 72.965 ;
        RECT 73.335 72.735 73.665 73.135 ;
        RECT 74.090 72.600 74.620 72.965 ;
        RECT 74.810 72.795 75.085 72.965 ;
        RECT 74.805 72.625 75.085 72.795 ;
        RECT 74.090 72.565 74.265 72.600 ;
        RECT 73.335 72.395 74.265 72.565 ;
        RECT 71.505 72.155 72.735 72.325 ;
        RECT 70.295 71.435 71.305 71.605 ;
        RECT 71.475 71.590 72.225 71.780 ;
        RECT 69.955 71.095 71.080 71.265 ;
        RECT 71.475 70.925 71.645 71.590 ;
        RECT 72.395 71.345 72.735 72.155 ;
        RECT 69.615 70.755 71.645 70.925 ;
        RECT 71.815 70.585 71.985 71.345 ;
        RECT 72.220 70.935 72.735 71.345 ;
        RECT 72.910 71.725 73.080 72.395 ;
        RECT 73.335 72.225 73.505 72.395 ;
        RECT 73.250 71.895 73.505 72.225 ;
        RECT 73.730 71.895 73.925 72.225 ;
        RECT 72.910 70.755 73.245 71.725 ;
        RECT 73.415 70.585 73.585 71.725 ;
        RECT 73.755 70.925 73.925 71.895 ;
        RECT 74.095 71.265 74.265 72.395 ;
        RECT 74.435 71.605 74.605 72.405 ;
        RECT 74.810 71.805 75.085 72.625 ;
        RECT 75.255 71.605 75.445 72.965 ;
        RECT 75.625 72.600 76.135 73.135 ;
        RECT 76.355 72.325 76.600 72.930 ;
        RECT 77.045 72.395 77.430 72.965 ;
        RECT 77.600 72.675 77.925 73.135 ;
        RECT 78.445 72.505 78.725 72.965 ;
        RECT 75.645 72.155 76.875 72.325 ;
        RECT 74.435 71.435 75.445 71.605 ;
        RECT 75.615 71.590 76.365 71.780 ;
        RECT 74.095 71.095 75.220 71.265 ;
        RECT 75.615 70.925 75.785 71.590 ;
        RECT 76.535 71.345 76.875 72.155 ;
        RECT 73.755 70.755 75.785 70.925 ;
        RECT 75.955 70.585 76.125 71.345 ;
        RECT 76.360 70.935 76.875 71.345 ;
        RECT 77.045 71.725 77.325 72.395 ;
        RECT 77.600 72.335 78.725 72.505 ;
        RECT 77.600 72.225 78.050 72.335 ;
        RECT 77.495 71.895 78.050 72.225 ;
        RECT 78.915 72.165 79.315 72.965 ;
        RECT 79.715 72.675 79.985 73.135 ;
        RECT 80.155 72.505 80.440 72.965 ;
        RECT 80.835 72.755 82.005 72.965 ;
        RECT 80.835 72.735 81.165 72.755 ;
        RECT 77.045 70.755 77.430 71.725 ;
        RECT 77.600 71.435 78.050 71.895 ;
        RECT 78.220 71.605 79.315 72.165 ;
        RECT 77.600 71.215 78.725 71.435 ;
        RECT 77.600 70.585 77.925 71.045 ;
        RECT 78.445 70.755 78.725 71.215 ;
        RECT 78.915 70.755 79.315 71.605 ;
        RECT 79.485 72.335 80.440 72.505 ;
        RECT 79.485 71.435 79.695 72.335 ;
        RECT 80.725 72.315 81.585 72.565 ;
        RECT 81.755 72.505 82.005 72.755 ;
        RECT 82.175 72.675 82.345 73.135 ;
        RECT 82.515 72.505 82.855 72.965 ;
        RECT 81.755 72.335 82.855 72.505 ;
        RECT 83.115 72.585 83.285 72.965 ;
        RECT 83.465 72.755 83.795 73.135 ;
        RECT 83.115 72.415 83.780 72.585 ;
        RECT 83.975 72.460 84.235 72.965 ;
        RECT 79.865 71.605 80.555 72.165 ;
        RECT 80.725 71.725 81.005 72.315 ;
        RECT 81.175 71.895 81.925 72.145 ;
        RECT 82.095 71.895 82.855 72.145 ;
        RECT 83.045 71.865 83.375 72.235 ;
        RECT 83.610 72.160 83.780 72.415 ;
        RECT 83.610 71.830 83.895 72.160 ;
        RECT 80.725 71.555 82.425 71.725 ;
        RECT 79.485 71.215 80.440 71.435 ;
        RECT 79.715 70.585 79.985 71.045 ;
        RECT 80.155 70.755 80.440 71.215 ;
        RECT 80.830 70.585 81.085 71.385 ;
        RECT 81.255 70.755 81.585 71.555 ;
        RECT 81.755 70.585 81.925 71.385 ;
        RECT 82.095 70.755 82.425 71.555 ;
        RECT 82.595 70.585 82.855 71.725 ;
        RECT 83.610 71.685 83.780 71.830 ;
        RECT 83.115 71.515 83.780 71.685 ;
        RECT 84.065 71.660 84.235 72.460 ;
        RECT 84.410 72.370 84.865 73.135 ;
        RECT 85.140 72.755 86.440 72.965 ;
        RECT 86.695 72.775 87.025 73.135 ;
        RECT 86.270 72.605 86.440 72.755 ;
        RECT 87.195 72.635 87.455 72.965 ;
        RECT 85.340 72.145 85.560 72.545 ;
        RECT 84.405 71.945 84.895 72.145 ;
        RECT 85.085 71.935 85.560 72.145 ;
        RECT 85.805 72.145 86.015 72.545 ;
        RECT 86.270 72.480 87.025 72.605 ;
        RECT 86.270 72.435 87.115 72.480 ;
        RECT 86.845 72.315 87.115 72.435 ;
        RECT 85.805 71.935 86.135 72.145 ;
        RECT 86.305 71.875 86.715 72.180 ;
        RECT 83.115 70.755 83.285 71.515 ;
        RECT 83.465 70.585 83.795 71.345 ;
        RECT 83.965 70.755 84.235 71.660 ;
        RECT 84.410 71.705 85.585 71.765 ;
        RECT 86.945 71.740 87.115 72.315 ;
        RECT 86.915 71.705 87.115 71.740 ;
        RECT 84.410 71.595 87.115 71.705 ;
        RECT 84.410 70.975 84.665 71.595 ;
        RECT 85.255 71.535 87.055 71.595 ;
        RECT 85.255 71.505 85.585 71.535 ;
        RECT 87.285 71.435 87.455 72.635 ;
        RECT 88.545 72.385 89.755 73.135 ;
        RECT 84.915 71.335 85.100 71.425 ;
        RECT 85.690 71.335 86.525 71.345 ;
        RECT 84.915 71.135 86.525 71.335 ;
        RECT 84.915 71.095 85.145 71.135 ;
        RECT 84.410 70.755 84.745 70.975 ;
        RECT 85.750 70.585 86.105 70.965 ;
        RECT 86.275 70.755 86.525 71.135 ;
        RECT 86.775 70.585 87.025 71.365 ;
        RECT 87.195 70.755 87.455 71.435 ;
        RECT 88.545 71.675 89.065 72.215 ;
        RECT 89.235 71.845 89.755 72.385 ;
        RECT 88.545 70.585 89.755 71.675 ;
        RECT 12.100 70.415 89.840 70.585 ;
        RECT 12.185 69.325 13.395 70.415 ;
        RECT 12.185 68.615 12.705 69.155 ;
        RECT 12.875 68.785 13.395 69.325 ;
        RECT 14.035 69.465 14.310 70.235 ;
        RECT 14.480 69.805 14.810 70.235 ;
        RECT 14.980 69.975 15.175 70.415 ;
        RECT 15.355 69.805 15.685 70.235 ;
        RECT 14.480 69.635 15.685 69.805 ;
        RECT 15.865 69.860 16.470 70.415 ;
        RECT 16.645 69.905 17.125 70.245 ;
        RECT 17.295 69.870 17.550 70.415 ;
        RECT 15.865 69.760 16.480 69.860 ;
        RECT 14.035 69.275 14.620 69.465 ;
        RECT 14.790 69.305 15.685 69.635 ;
        RECT 16.295 69.735 16.480 69.760 ;
        RECT 12.185 67.865 13.395 68.615 ;
        RECT 14.035 68.455 14.275 69.105 ;
        RECT 14.445 68.605 14.620 69.275 ;
        RECT 15.865 69.140 16.125 69.590 ;
        RECT 16.295 69.490 16.625 69.735 ;
        RECT 16.795 69.415 17.550 69.665 ;
        RECT 17.720 69.545 17.995 70.245 ;
        RECT 16.780 69.380 17.550 69.415 ;
        RECT 16.765 69.370 17.550 69.380 ;
        RECT 16.760 69.355 17.655 69.370 ;
        RECT 16.740 69.340 17.655 69.355 ;
        RECT 16.720 69.330 17.655 69.340 ;
        RECT 16.695 69.320 17.655 69.330 ;
        RECT 16.625 69.290 17.655 69.320 ;
        RECT 16.605 69.260 17.655 69.290 ;
        RECT 16.585 69.230 17.655 69.260 ;
        RECT 16.555 69.205 17.655 69.230 ;
        RECT 16.520 69.170 17.655 69.205 ;
        RECT 16.490 69.165 17.655 69.170 ;
        RECT 16.490 69.160 16.880 69.165 ;
        RECT 16.490 69.150 16.855 69.160 ;
        RECT 16.490 69.145 16.840 69.150 ;
        RECT 16.490 69.140 16.825 69.145 ;
        RECT 15.865 69.135 16.825 69.140 ;
        RECT 15.865 69.125 16.815 69.135 ;
        RECT 15.865 69.120 16.805 69.125 ;
        RECT 15.865 69.110 16.795 69.120 ;
        RECT 14.790 68.775 15.205 69.105 ;
        RECT 15.385 68.775 15.680 69.105 ;
        RECT 15.865 69.100 16.790 69.110 ;
        RECT 15.865 69.095 16.785 69.100 ;
        RECT 15.865 69.080 16.775 69.095 ;
        RECT 15.865 69.065 16.770 69.080 ;
        RECT 15.865 69.040 16.760 69.065 ;
        RECT 15.865 68.970 16.755 69.040 ;
        RECT 14.445 68.425 14.775 68.605 ;
        RECT 14.050 67.865 14.380 68.255 ;
        RECT 14.550 68.045 14.775 68.425 ;
        RECT 14.975 68.155 15.205 68.775 ;
        RECT 15.385 67.865 15.685 68.595 ;
        RECT 15.865 68.415 16.415 68.800 ;
        RECT 16.585 68.245 16.755 68.970 ;
        RECT 15.865 68.075 16.755 68.245 ;
        RECT 16.925 68.570 17.255 68.995 ;
        RECT 17.425 68.770 17.655 69.165 ;
        RECT 16.925 68.085 17.145 68.570 ;
        RECT 17.825 68.515 17.995 69.545 ;
        RECT 17.315 67.865 17.565 68.405 ;
        RECT 17.735 68.035 17.995 68.515 ;
        RECT 18.165 69.985 18.505 70.245 ;
        RECT 18.165 68.585 18.425 69.985 ;
        RECT 18.675 69.615 19.005 70.415 ;
        RECT 19.470 69.445 19.720 70.245 ;
        RECT 19.905 69.695 20.235 70.415 ;
        RECT 20.455 69.445 20.705 70.245 ;
        RECT 20.875 70.035 21.210 70.415 ;
        RECT 18.615 69.275 20.805 69.445 ;
        RECT 18.615 69.105 18.930 69.275 ;
        RECT 18.600 68.855 18.930 69.105 ;
        RECT 18.165 68.075 18.505 68.585 ;
        RECT 18.675 67.865 18.945 68.665 ;
        RECT 19.125 68.135 19.405 69.105 ;
        RECT 19.585 68.135 19.885 69.105 ;
        RECT 20.065 68.140 20.415 69.105 ;
        RECT 20.635 68.365 20.805 69.275 ;
        RECT 20.975 68.545 21.215 69.855 ;
        RECT 22.305 68.810 22.585 70.245 ;
        RECT 22.755 69.640 23.465 70.415 ;
        RECT 23.635 69.470 23.965 70.245 ;
        RECT 22.815 69.255 23.965 69.470 ;
        RECT 20.635 68.035 21.130 68.365 ;
        RECT 22.305 68.035 22.645 68.810 ;
        RECT 22.815 68.685 23.100 69.255 ;
        RECT 23.285 68.855 23.755 69.085 ;
        RECT 24.160 69.055 24.375 70.170 ;
        RECT 24.555 69.695 24.885 70.415 ;
        RECT 24.665 69.055 24.895 69.395 ;
        RECT 25.065 69.250 25.355 70.415 ;
        RECT 25.525 69.325 27.195 70.415 ;
        RECT 27.370 70.035 27.705 70.415 ;
        RECT 23.925 68.875 24.375 69.055 ;
        RECT 23.925 68.855 24.255 68.875 ;
        RECT 24.565 68.855 24.895 69.055 ;
        RECT 22.815 68.495 23.525 68.685 ;
        RECT 23.225 68.355 23.525 68.495 ;
        RECT 23.715 68.495 24.895 68.685 ;
        RECT 25.525 68.635 26.275 69.155 ;
        RECT 26.445 68.805 27.195 69.325 ;
        RECT 23.715 68.415 24.045 68.495 ;
        RECT 23.225 68.345 23.540 68.355 ;
        RECT 23.225 68.335 23.550 68.345 ;
        RECT 23.225 68.330 23.560 68.335 ;
        RECT 22.815 67.865 22.985 68.325 ;
        RECT 23.225 68.320 23.565 68.330 ;
        RECT 23.225 68.315 23.570 68.320 ;
        RECT 23.225 68.305 23.575 68.315 ;
        RECT 23.225 68.300 23.580 68.305 ;
        RECT 23.225 68.035 23.585 68.300 ;
        RECT 24.215 67.865 24.385 68.325 ;
        RECT 24.555 68.035 24.895 68.495 ;
        RECT 25.065 67.865 25.355 68.590 ;
        RECT 25.525 67.865 27.195 68.635 ;
        RECT 27.365 68.545 27.605 69.855 ;
        RECT 27.875 69.445 28.125 70.245 ;
        RECT 28.345 69.695 28.675 70.415 ;
        RECT 28.860 69.445 29.110 70.245 ;
        RECT 29.575 69.615 29.905 70.415 ;
        RECT 30.075 69.985 30.415 70.245 ;
        RECT 27.775 69.275 29.965 69.445 ;
        RECT 27.775 68.365 27.945 69.275 ;
        RECT 29.650 69.105 29.965 69.275 ;
        RECT 27.450 68.035 27.945 68.365 ;
        RECT 28.165 68.140 28.515 69.105 ;
        RECT 28.695 68.135 28.995 69.105 ;
        RECT 29.175 68.135 29.455 69.105 ;
        RECT 29.650 68.855 29.980 69.105 ;
        RECT 29.635 67.865 29.905 68.665 ;
        RECT 30.155 68.585 30.415 69.985 ;
        RECT 30.675 69.745 30.845 70.245 ;
        RECT 31.015 69.915 31.345 70.415 ;
        RECT 30.675 69.575 31.340 69.745 ;
        RECT 30.590 68.755 30.940 69.405 ;
        RECT 31.110 68.585 31.340 69.575 ;
        RECT 30.075 68.075 30.415 68.585 ;
        RECT 30.675 68.415 31.340 68.585 ;
        RECT 30.675 68.125 30.845 68.415 ;
        RECT 31.015 67.865 31.345 68.245 ;
        RECT 31.515 68.125 31.700 70.245 ;
        RECT 31.940 69.955 32.205 70.415 ;
        RECT 32.375 69.820 32.625 70.245 ;
        RECT 32.835 69.970 33.940 70.140 ;
        RECT 32.320 69.690 32.625 69.820 ;
        RECT 31.870 68.495 32.150 69.445 ;
        RECT 32.320 68.585 32.490 69.690 ;
        RECT 32.660 68.905 32.900 69.500 ;
        RECT 33.070 69.435 33.600 69.800 ;
        RECT 33.070 68.735 33.240 69.435 ;
        RECT 33.770 69.355 33.940 69.970 ;
        RECT 34.110 69.615 34.280 70.415 ;
        RECT 34.450 69.915 34.700 70.245 ;
        RECT 34.925 69.945 35.810 70.115 ;
        RECT 33.770 69.265 34.280 69.355 ;
        RECT 32.320 68.455 32.545 68.585 ;
        RECT 32.715 68.515 33.240 68.735 ;
        RECT 33.410 69.095 34.280 69.265 ;
        RECT 31.955 67.865 32.205 68.325 ;
        RECT 32.375 68.315 32.545 68.455 ;
        RECT 33.410 68.315 33.580 69.095 ;
        RECT 34.110 69.025 34.280 69.095 ;
        RECT 33.790 68.845 33.990 68.875 ;
        RECT 34.450 68.845 34.620 69.915 ;
        RECT 34.790 69.025 34.980 69.745 ;
        RECT 33.790 68.545 34.620 68.845 ;
        RECT 35.150 68.815 35.470 69.775 ;
        RECT 32.375 68.145 32.710 68.315 ;
        RECT 32.905 68.145 33.580 68.315 ;
        RECT 33.900 67.865 34.270 68.365 ;
        RECT 34.450 68.315 34.620 68.545 ;
        RECT 35.005 68.485 35.470 68.815 ;
        RECT 35.640 69.105 35.810 69.945 ;
        RECT 35.990 69.915 36.305 70.415 ;
        RECT 36.535 69.685 36.875 70.245 ;
        RECT 35.980 69.310 36.875 69.685 ;
        RECT 37.045 69.405 37.215 70.415 ;
        RECT 36.685 69.105 36.875 69.310 ;
        RECT 37.385 69.355 37.715 70.200 ;
        RECT 37.385 69.275 37.775 69.355 ;
        RECT 37.560 69.225 37.775 69.275 ;
        RECT 35.640 68.775 36.515 69.105 ;
        RECT 36.685 68.775 37.435 69.105 ;
        RECT 35.640 68.315 35.810 68.775 ;
        RECT 36.685 68.605 36.885 68.775 ;
        RECT 37.605 68.645 37.775 69.225 ;
        RECT 37.550 68.605 37.775 68.645 ;
        RECT 34.450 68.145 34.855 68.315 ;
        RECT 35.025 68.145 35.810 68.315 ;
        RECT 36.085 67.865 36.295 68.395 ;
        RECT 36.555 68.080 36.885 68.605 ;
        RECT 37.395 68.520 37.775 68.605 ;
        RECT 37.055 67.865 37.225 68.475 ;
        RECT 37.395 68.085 37.725 68.520 ;
        RECT 37.955 68.045 38.215 70.235 ;
        RECT 38.385 69.685 38.725 70.415 ;
        RECT 38.905 69.505 39.175 70.235 ;
        RECT 38.405 69.285 39.175 69.505 ;
        RECT 39.355 69.525 39.585 70.235 ;
        RECT 39.755 69.705 40.085 70.415 ;
        RECT 40.255 69.525 40.515 70.235 ;
        RECT 40.795 69.745 40.965 70.245 ;
        RECT 41.135 69.915 41.465 70.415 ;
        RECT 40.795 69.575 41.460 69.745 ;
        RECT 39.355 69.285 40.515 69.525 ;
        RECT 38.405 68.615 38.695 69.285 ;
        RECT 38.875 68.795 39.340 69.105 ;
        RECT 39.520 68.795 40.045 69.105 ;
        RECT 38.405 68.415 39.635 68.615 ;
        RECT 38.475 67.865 39.145 68.235 ;
        RECT 39.325 68.045 39.635 68.415 ;
        RECT 39.815 68.155 40.045 68.795 ;
        RECT 40.225 68.775 40.525 69.105 ;
        RECT 40.710 68.755 41.060 69.405 ;
        RECT 40.225 67.865 40.515 68.595 ;
        RECT 41.230 68.585 41.460 69.575 ;
        RECT 40.795 68.415 41.460 68.585 ;
        RECT 40.795 68.125 40.965 68.415 ;
        RECT 41.135 67.865 41.465 68.245 ;
        RECT 41.635 68.125 41.820 70.245 ;
        RECT 42.060 69.955 42.325 70.415 ;
        RECT 42.495 69.820 42.745 70.245 ;
        RECT 42.955 69.970 44.060 70.140 ;
        RECT 42.440 69.690 42.745 69.820 ;
        RECT 41.990 68.495 42.270 69.445 ;
        RECT 42.440 68.585 42.610 69.690 ;
        RECT 42.780 68.905 43.020 69.500 ;
        RECT 43.190 69.435 43.720 69.800 ;
        RECT 43.190 68.735 43.360 69.435 ;
        RECT 43.890 69.355 44.060 69.970 ;
        RECT 44.230 69.615 44.400 70.415 ;
        RECT 44.570 69.915 44.820 70.245 ;
        RECT 45.045 69.945 45.930 70.115 ;
        RECT 43.890 69.265 44.400 69.355 ;
        RECT 42.440 68.455 42.665 68.585 ;
        RECT 42.835 68.515 43.360 68.735 ;
        RECT 43.530 69.095 44.400 69.265 ;
        RECT 42.075 67.865 42.325 68.325 ;
        RECT 42.495 68.315 42.665 68.455 ;
        RECT 43.530 68.315 43.700 69.095 ;
        RECT 44.230 69.025 44.400 69.095 ;
        RECT 43.910 68.845 44.110 68.875 ;
        RECT 44.570 68.845 44.740 69.915 ;
        RECT 44.910 69.025 45.100 69.745 ;
        RECT 43.910 68.545 44.740 68.845 ;
        RECT 45.270 68.815 45.590 69.775 ;
        RECT 42.495 68.145 42.830 68.315 ;
        RECT 43.025 68.145 43.700 68.315 ;
        RECT 44.020 67.865 44.390 68.365 ;
        RECT 44.570 68.315 44.740 68.545 ;
        RECT 45.125 68.485 45.590 68.815 ;
        RECT 45.760 69.105 45.930 69.945 ;
        RECT 46.110 69.915 46.425 70.415 ;
        RECT 46.655 69.685 46.995 70.245 ;
        RECT 46.100 69.310 46.995 69.685 ;
        RECT 47.165 69.405 47.335 70.415 ;
        RECT 46.805 69.105 46.995 69.310 ;
        RECT 47.505 69.355 47.835 70.200 ;
        RECT 48.250 69.445 48.640 69.620 ;
        RECT 49.125 69.615 49.455 70.415 ;
        RECT 49.625 69.625 50.160 70.245 ;
        RECT 47.505 69.275 47.895 69.355 ;
        RECT 48.250 69.275 49.675 69.445 ;
        RECT 47.680 69.225 47.895 69.275 ;
        RECT 45.760 68.775 46.635 69.105 ;
        RECT 46.805 68.775 47.555 69.105 ;
        RECT 45.760 68.315 45.930 68.775 ;
        RECT 46.805 68.605 47.005 68.775 ;
        RECT 47.725 68.645 47.895 69.225 ;
        RECT 47.670 68.605 47.895 68.645 ;
        RECT 44.570 68.145 44.975 68.315 ;
        RECT 45.145 68.145 45.930 68.315 ;
        RECT 46.205 67.865 46.415 68.395 ;
        RECT 46.675 68.080 47.005 68.605 ;
        RECT 47.515 68.520 47.895 68.605 ;
        RECT 48.125 68.545 48.480 69.105 ;
        RECT 47.175 67.865 47.345 68.475 ;
        RECT 47.515 68.085 47.845 68.520 ;
        RECT 48.650 68.375 48.820 69.275 ;
        RECT 48.990 68.545 49.255 69.105 ;
        RECT 49.505 68.775 49.675 69.275 ;
        RECT 49.845 68.605 50.160 69.625 ;
        RECT 50.825 69.250 51.115 70.415 ;
        RECT 51.345 69.275 51.555 70.415 ;
        RECT 51.725 69.265 52.055 70.245 ;
        RECT 52.225 69.275 52.455 70.415 ;
        RECT 52.670 69.275 53.005 70.245 ;
        RECT 53.175 69.275 53.345 70.415 ;
        RECT 53.515 70.075 55.545 70.245 ;
        RECT 48.230 67.865 48.470 68.375 ;
        RECT 48.650 68.045 48.930 68.375 ;
        RECT 49.160 67.865 49.375 68.375 ;
        RECT 49.545 68.035 50.160 68.605 ;
        RECT 50.825 67.865 51.115 68.590 ;
        RECT 51.345 67.865 51.555 68.685 ;
        RECT 51.725 68.665 51.975 69.265 ;
        RECT 52.145 68.855 52.475 69.105 ;
        RECT 51.725 68.035 52.055 68.665 ;
        RECT 52.225 67.865 52.455 68.685 ;
        RECT 52.670 68.605 52.840 69.275 ;
        RECT 53.515 69.105 53.685 70.075 ;
        RECT 53.010 68.775 53.265 69.105 ;
        RECT 53.490 68.775 53.685 69.105 ;
        RECT 53.855 69.735 54.980 69.905 ;
        RECT 53.095 68.605 53.265 68.775 ;
        RECT 53.855 68.605 54.025 69.735 ;
        RECT 52.670 68.035 52.925 68.605 ;
        RECT 53.095 68.435 54.025 68.605 ;
        RECT 54.195 69.395 55.205 69.565 ;
        RECT 54.195 68.595 54.365 69.395 ;
        RECT 54.570 69.055 54.845 69.195 ;
        RECT 54.565 68.885 54.845 69.055 ;
        RECT 53.850 68.400 54.025 68.435 ;
        RECT 53.095 67.865 53.425 68.265 ;
        RECT 53.850 68.035 54.380 68.400 ;
        RECT 54.570 68.035 54.845 68.885 ;
        RECT 55.015 68.035 55.205 69.395 ;
        RECT 55.375 69.410 55.545 70.075 ;
        RECT 55.715 69.655 55.885 70.415 ;
        RECT 56.120 69.655 56.635 70.065 ;
        RECT 55.375 69.220 56.125 69.410 ;
        RECT 56.295 68.845 56.635 69.655 ;
        RECT 56.865 69.355 57.195 70.200 ;
        RECT 57.365 69.405 57.535 70.415 ;
        RECT 57.705 69.685 58.045 70.245 ;
        RECT 58.275 69.915 58.590 70.415 ;
        RECT 58.770 69.945 59.655 70.115 ;
        RECT 55.405 68.675 56.635 68.845 ;
        RECT 56.805 69.275 57.195 69.355 ;
        RECT 57.705 69.310 58.600 69.685 ;
        RECT 56.805 69.225 57.020 69.275 ;
        RECT 55.385 67.865 55.895 68.400 ;
        RECT 56.115 68.070 56.360 68.675 ;
        RECT 56.805 68.645 56.975 69.225 ;
        RECT 57.705 69.105 57.895 69.310 ;
        RECT 58.770 69.105 58.940 69.945 ;
        RECT 59.880 69.915 60.130 70.245 ;
        RECT 57.145 68.775 57.895 69.105 ;
        RECT 58.065 68.775 58.940 69.105 ;
        RECT 56.805 68.605 57.030 68.645 ;
        RECT 57.695 68.605 57.895 68.775 ;
        RECT 56.805 68.520 57.185 68.605 ;
        RECT 56.855 68.085 57.185 68.520 ;
        RECT 57.355 67.865 57.525 68.475 ;
        RECT 57.695 68.080 58.025 68.605 ;
        RECT 58.285 67.865 58.495 68.395 ;
        RECT 58.770 68.315 58.940 68.775 ;
        RECT 59.110 68.815 59.430 69.775 ;
        RECT 59.600 69.025 59.790 69.745 ;
        RECT 59.960 68.845 60.130 69.915 ;
        RECT 60.300 69.615 60.470 70.415 ;
        RECT 60.640 69.970 61.745 70.140 ;
        RECT 60.640 69.355 60.810 69.970 ;
        RECT 61.955 69.820 62.205 70.245 ;
        RECT 62.375 69.955 62.640 70.415 ;
        RECT 60.980 69.435 61.510 69.800 ;
        RECT 61.955 69.690 62.260 69.820 ;
        RECT 60.300 69.265 60.810 69.355 ;
        RECT 60.300 69.095 61.170 69.265 ;
        RECT 60.300 69.025 60.470 69.095 ;
        RECT 60.590 68.845 60.790 68.875 ;
        RECT 59.110 68.485 59.575 68.815 ;
        RECT 59.960 68.545 60.790 68.845 ;
        RECT 59.960 68.315 60.130 68.545 ;
        RECT 58.770 68.145 59.555 68.315 ;
        RECT 59.725 68.145 60.130 68.315 ;
        RECT 60.310 67.865 60.680 68.365 ;
        RECT 61.000 68.315 61.170 69.095 ;
        RECT 61.340 68.735 61.510 69.435 ;
        RECT 61.680 68.905 61.920 69.500 ;
        RECT 61.340 68.515 61.865 68.735 ;
        RECT 62.090 68.585 62.260 69.690 ;
        RECT 62.035 68.455 62.260 68.585 ;
        RECT 62.430 68.495 62.710 69.445 ;
        RECT 62.035 68.315 62.205 68.455 ;
        RECT 61.000 68.145 61.675 68.315 ;
        RECT 61.870 68.145 62.205 68.315 ;
        RECT 62.375 67.865 62.625 68.325 ;
        RECT 62.880 68.125 63.065 70.245 ;
        RECT 63.235 69.915 63.565 70.415 ;
        RECT 63.735 69.745 63.905 70.245 ;
        RECT 63.240 69.575 63.905 69.745 ;
        RECT 63.240 68.585 63.470 69.575 ;
        RECT 63.640 68.755 63.990 69.405 ;
        RECT 64.630 69.265 64.890 70.415 ;
        RECT 65.065 69.340 65.320 70.245 ;
        RECT 65.490 69.655 65.820 70.415 ;
        RECT 66.035 69.485 66.205 70.245 ;
        RECT 66.555 69.745 66.725 70.245 ;
        RECT 66.895 69.915 67.225 70.415 ;
        RECT 66.555 69.575 67.220 69.745 ;
        RECT 63.240 68.415 63.905 68.585 ;
        RECT 63.235 67.865 63.565 68.245 ;
        RECT 63.735 68.125 63.905 68.415 ;
        RECT 64.630 67.865 64.890 68.705 ;
        RECT 65.065 68.610 65.235 69.340 ;
        RECT 65.490 69.315 66.205 69.485 ;
        RECT 65.490 69.105 65.660 69.315 ;
        RECT 65.405 68.775 65.660 69.105 ;
        RECT 65.065 68.035 65.320 68.610 ;
        RECT 65.490 68.585 65.660 68.775 ;
        RECT 65.940 68.765 66.295 69.135 ;
        RECT 66.470 68.755 66.820 69.405 ;
        RECT 66.990 68.585 67.220 69.575 ;
        RECT 65.490 68.415 66.205 68.585 ;
        RECT 65.490 67.865 65.820 68.245 ;
        RECT 66.035 68.035 66.205 68.415 ;
        RECT 66.555 68.415 67.220 68.585 ;
        RECT 66.555 68.125 66.725 68.415 ;
        RECT 66.895 67.865 67.225 68.245 ;
        RECT 67.395 68.125 67.580 70.245 ;
        RECT 67.820 69.955 68.085 70.415 ;
        RECT 68.255 69.820 68.505 70.245 ;
        RECT 68.715 69.970 69.820 70.140 ;
        RECT 68.200 69.690 68.505 69.820 ;
        RECT 67.750 68.495 68.030 69.445 ;
        RECT 68.200 68.585 68.370 69.690 ;
        RECT 68.540 68.905 68.780 69.500 ;
        RECT 68.950 69.435 69.480 69.800 ;
        RECT 68.950 68.735 69.120 69.435 ;
        RECT 69.650 69.355 69.820 69.970 ;
        RECT 69.990 69.615 70.160 70.415 ;
        RECT 70.330 69.915 70.580 70.245 ;
        RECT 70.805 69.945 71.690 70.115 ;
        RECT 69.650 69.265 70.160 69.355 ;
        RECT 68.200 68.455 68.425 68.585 ;
        RECT 68.595 68.515 69.120 68.735 ;
        RECT 69.290 69.095 70.160 69.265 ;
        RECT 67.835 67.865 68.085 68.325 ;
        RECT 68.255 68.315 68.425 68.455 ;
        RECT 69.290 68.315 69.460 69.095 ;
        RECT 69.990 69.025 70.160 69.095 ;
        RECT 69.670 68.845 69.870 68.875 ;
        RECT 70.330 68.845 70.500 69.915 ;
        RECT 70.670 69.025 70.860 69.745 ;
        RECT 69.670 68.545 70.500 68.845 ;
        RECT 71.030 68.815 71.350 69.775 ;
        RECT 68.255 68.145 68.590 68.315 ;
        RECT 68.785 68.145 69.460 68.315 ;
        RECT 69.780 67.865 70.150 68.365 ;
        RECT 70.330 68.315 70.500 68.545 ;
        RECT 70.885 68.485 71.350 68.815 ;
        RECT 71.520 69.105 71.690 69.945 ;
        RECT 71.870 69.915 72.185 70.415 ;
        RECT 72.415 69.685 72.755 70.245 ;
        RECT 71.860 69.310 72.755 69.685 ;
        RECT 72.925 69.405 73.095 70.415 ;
        RECT 72.565 69.105 72.755 69.310 ;
        RECT 73.265 69.355 73.595 70.200 ;
        RECT 73.265 69.275 73.655 69.355 ;
        RECT 73.835 69.275 74.165 70.415 ;
        RECT 73.440 69.225 73.655 69.275 ;
        RECT 71.520 68.775 72.395 69.105 ;
        RECT 72.565 68.775 73.315 69.105 ;
        RECT 71.520 68.315 71.690 68.775 ;
        RECT 72.565 68.605 72.765 68.775 ;
        RECT 73.485 68.645 73.655 69.225 ;
        RECT 73.430 68.605 73.655 68.645 ;
        RECT 70.330 68.145 70.735 68.315 ;
        RECT 70.905 68.145 71.690 68.315 ;
        RECT 71.965 67.865 72.175 68.395 ;
        RECT 72.435 68.080 72.765 68.605 ;
        RECT 73.275 68.520 73.655 68.605 ;
        RECT 73.825 68.525 74.165 69.105 ;
        RECT 74.335 69.075 74.695 70.245 ;
        RECT 74.895 69.245 75.225 70.415 ;
        RECT 75.425 69.075 75.755 70.245 ;
        RECT 75.955 69.245 76.285 70.415 ;
        RECT 76.585 69.250 76.875 70.415 ;
        RECT 77.055 69.305 77.350 70.415 ;
        RECT 77.530 69.105 77.780 70.240 ;
        RECT 77.950 69.305 78.210 70.415 ;
        RECT 78.380 69.515 78.640 70.240 ;
        RECT 78.810 69.685 79.070 70.415 ;
        RECT 79.240 69.515 79.500 70.240 ;
        RECT 79.670 69.685 79.930 70.415 ;
        RECT 80.100 69.515 80.360 70.240 ;
        RECT 80.530 69.685 80.790 70.415 ;
        RECT 80.960 69.515 81.220 70.240 ;
        RECT 81.390 69.685 81.685 70.415 ;
        RECT 78.380 69.275 81.690 69.515 ;
        RECT 74.335 68.795 75.755 69.075 ;
        RECT 72.935 67.865 73.105 68.475 ;
        RECT 73.275 68.085 73.605 68.520 ;
        RECT 74.335 68.460 74.695 68.795 ;
        RECT 73.835 67.865 74.165 68.355 ;
        RECT 74.335 68.035 74.955 68.460 ;
        RECT 75.415 67.865 75.745 68.555 ;
        RECT 76.585 67.865 76.875 68.590 ;
        RECT 77.045 68.495 77.360 69.105 ;
        RECT 77.530 68.855 80.550 69.105 ;
        RECT 77.105 67.865 77.350 68.325 ;
        RECT 77.530 68.045 77.780 68.855 ;
        RECT 80.720 68.685 81.690 69.275 ;
        RECT 78.380 68.515 81.690 68.685 ;
        RECT 82.105 69.275 82.445 70.245 ;
        RECT 82.615 69.275 82.785 70.415 ;
        RECT 83.055 69.615 83.305 70.415 ;
        RECT 83.950 69.445 84.280 70.245 ;
        RECT 84.580 69.615 84.910 70.415 ;
        RECT 85.080 69.445 85.410 70.245 ;
        RECT 82.975 69.275 85.410 69.445 ;
        RECT 85.970 69.445 86.360 69.620 ;
        RECT 86.845 69.615 87.175 70.415 ;
        RECT 87.345 69.625 87.880 70.245 ;
        RECT 85.970 69.275 87.395 69.445 ;
        RECT 82.105 68.665 82.280 69.275 ;
        RECT 82.975 69.025 83.145 69.275 ;
        RECT 82.450 68.855 83.145 69.025 ;
        RECT 83.320 68.855 83.740 69.055 ;
        RECT 83.910 68.855 84.240 69.055 ;
        RECT 84.410 68.855 84.740 69.055 ;
        RECT 77.950 67.865 78.210 68.390 ;
        RECT 78.380 68.060 78.640 68.515 ;
        RECT 78.810 67.865 79.070 68.345 ;
        RECT 79.240 68.060 79.500 68.515 ;
        RECT 79.670 67.865 79.930 68.345 ;
        RECT 80.100 68.060 80.360 68.515 ;
        RECT 80.530 67.865 80.790 68.345 ;
        RECT 80.960 68.060 81.220 68.515 ;
        RECT 81.390 67.865 81.690 68.345 ;
        RECT 82.105 68.035 82.445 68.665 ;
        RECT 82.615 67.865 82.865 68.665 ;
        RECT 83.055 68.515 84.280 68.685 ;
        RECT 83.055 68.035 83.385 68.515 ;
        RECT 83.555 67.865 83.780 68.325 ;
        RECT 83.950 68.035 84.280 68.515 ;
        RECT 84.910 68.645 85.080 69.275 ;
        RECT 85.265 68.855 85.615 69.105 ;
        RECT 84.910 68.035 85.410 68.645 ;
        RECT 85.845 68.545 86.200 69.105 ;
        RECT 86.370 68.375 86.540 69.275 ;
        RECT 86.710 68.545 86.975 69.105 ;
        RECT 87.225 68.775 87.395 69.275 ;
        RECT 87.565 68.605 87.880 69.625 ;
        RECT 88.545 69.325 89.755 70.415 ;
        RECT 88.545 68.785 89.065 69.325 ;
        RECT 89.235 68.615 89.755 69.155 ;
        RECT 85.950 67.865 86.190 68.375 ;
        RECT 86.370 68.045 86.650 68.375 ;
        RECT 86.880 67.865 87.095 68.375 ;
        RECT 87.265 68.035 87.880 68.605 ;
        RECT 88.545 67.865 89.755 68.615 ;
        RECT 12.100 67.695 89.840 67.865 ;
        RECT 12.185 66.945 13.395 67.695 ;
        RECT 13.615 67.040 13.945 67.475 ;
        RECT 14.115 67.085 14.285 67.695 ;
        RECT 13.565 66.955 13.945 67.040 ;
        RECT 14.455 66.955 14.785 67.480 ;
        RECT 15.045 67.165 15.255 67.695 ;
        RECT 15.530 67.245 16.315 67.415 ;
        RECT 16.485 67.245 16.890 67.415 ;
        RECT 12.185 66.405 12.705 66.945 ;
        RECT 13.565 66.915 13.790 66.955 ;
        RECT 12.875 66.235 13.395 66.775 ;
        RECT 12.185 65.145 13.395 66.235 ;
        RECT 13.565 66.335 13.735 66.915 ;
        RECT 14.455 66.785 14.655 66.955 ;
        RECT 15.530 66.785 15.700 67.245 ;
        RECT 13.905 66.455 14.655 66.785 ;
        RECT 14.825 66.455 15.700 66.785 ;
        RECT 13.565 66.285 13.780 66.335 ;
        RECT 13.565 66.205 13.955 66.285 ;
        RECT 13.625 65.360 13.955 66.205 ;
        RECT 14.465 66.250 14.655 66.455 ;
        RECT 14.125 65.145 14.295 66.155 ;
        RECT 14.465 65.875 15.360 66.250 ;
        RECT 14.465 65.315 14.805 65.875 ;
        RECT 15.035 65.145 15.350 65.645 ;
        RECT 15.530 65.615 15.700 66.455 ;
        RECT 15.870 66.745 16.335 67.075 ;
        RECT 16.720 67.015 16.890 67.245 ;
        RECT 17.070 67.195 17.440 67.695 ;
        RECT 17.760 67.245 18.435 67.415 ;
        RECT 18.630 67.245 18.965 67.415 ;
        RECT 15.870 65.785 16.190 66.745 ;
        RECT 16.720 66.715 17.550 67.015 ;
        RECT 16.360 65.815 16.550 66.535 ;
        RECT 16.720 65.645 16.890 66.715 ;
        RECT 17.350 66.685 17.550 66.715 ;
        RECT 17.060 66.465 17.230 66.535 ;
        RECT 17.760 66.465 17.930 67.245 ;
        RECT 18.795 67.105 18.965 67.245 ;
        RECT 19.135 67.235 19.385 67.695 ;
        RECT 17.060 66.295 17.930 66.465 ;
        RECT 18.100 66.825 18.625 67.045 ;
        RECT 18.795 66.975 19.020 67.105 ;
        RECT 17.060 66.205 17.570 66.295 ;
        RECT 15.530 65.445 16.415 65.615 ;
        RECT 16.640 65.315 16.890 65.645 ;
        RECT 17.060 65.145 17.230 65.945 ;
        RECT 17.400 65.590 17.570 66.205 ;
        RECT 18.100 66.125 18.270 66.825 ;
        RECT 17.740 65.760 18.270 66.125 ;
        RECT 18.440 66.060 18.680 66.655 ;
        RECT 18.850 65.870 19.020 66.975 ;
        RECT 19.190 66.115 19.470 67.065 ;
        RECT 18.715 65.740 19.020 65.870 ;
        RECT 17.400 65.420 18.505 65.590 ;
        RECT 18.715 65.315 18.965 65.740 ;
        RECT 19.135 65.145 19.400 65.605 ;
        RECT 19.640 65.315 19.825 67.435 ;
        RECT 19.995 67.315 20.325 67.695 ;
        RECT 20.495 67.145 20.665 67.435 ;
        RECT 20.000 66.975 20.665 67.145 ;
        RECT 20.925 67.045 21.185 67.525 ;
        RECT 21.355 67.155 21.605 67.695 ;
        RECT 20.000 65.985 20.230 66.975 ;
        RECT 20.400 66.155 20.750 66.805 ;
        RECT 20.925 66.015 21.095 67.045 ;
        RECT 21.775 66.990 21.995 67.475 ;
        RECT 21.265 66.395 21.495 66.790 ;
        RECT 21.665 66.565 21.995 66.990 ;
        RECT 22.165 67.315 23.055 67.485 ;
        RECT 22.165 66.590 22.335 67.315 ;
        RECT 23.225 67.195 23.485 67.525 ;
        RECT 23.695 67.215 23.970 67.695 ;
        RECT 22.505 66.760 23.055 67.145 ;
        RECT 22.165 66.520 23.055 66.590 ;
        RECT 22.160 66.495 23.055 66.520 ;
        RECT 22.150 66.480 23.055 66.495 ;
        RECT 22.145 66.465 23.055 66.480 ;
        RECT 22.135 66.460 23.055 66.465 ;
        RECT 22.130 66.450 23.055 66.460 ;
        RECT 22.125 66.440 23.055 66.450 ;
        RECT 22.115 66.435 23.055 66.440 ;
        RECT 22.105 66.425 23.055 66.435 ;
        RECT 22.095 66.420 23.055 66.425 ;
        RECT 22.095 66.415 22.430 66.420 ;
        RECT 22.080 66.410 22.430 66.415 ;
        RECT 22.065 66.400 22.430 66.410 ;
        RECT 22.040 66.395 22.430 66.400 ;
        RECT 21.265 66.390 22.430 66.395 ;
        RECT 21.265 66.355 22.400 66.390 ;
        RECT 21.265 66.330 22.365 66.355 ;
        RECT 21.265 66.300 22.335 66.330 ;
        RECT 21.265 66.270 22.315 66.300 ;
        RECT 21.265 66.240 22.295 66.270 ;
        RECT 21.265 66.230 22.225 66.240 ;
        RECT 21.265 66.220 22.200 66.230 ;
        RECT 21.265 66.205 22.180 66.220 ;
        RECT 21.265 66.190 22.160 66.205 ;
        RECT 21.370 66.180 22.155 66.190 ;
        RECT 21.370 66.145 22.140 66.180 ;
        RECT 20.000 65.815 20.665 65.985 ;
        RECT 19.995 65.145 20.325 65.645 ;
        RECT 20.495 65.315 20.665 65.815 ;
        RECT 20.925 65.315 21.200 66.015 ;
        RECT 21.370 65.895 22.125 66.145 ;
        RECT 22.295 65.825 22.625 66.070 ;
        RECT 22.795 65.970 23.055 66.420 ;
        RECT 23.225 66.285 23.395 67.195 ;
        RECT 24.180 67.125 24.385 67.525 ;
        RECT 24.555 67.295 24.890 67.695 ;
        RECT 23.565 66.455 23.925 67.035 ;
        RECT 24.180 66.955 24.865 67.125 ;
        RECT 24.105 66.285 24.355 66.785 ;
        RECT 23.225 66.115 24.355 66.285 ;
        RECT 22.440 65.800 22.625 65.825 ;
        RECT 22.440 65.700 23.055 65.800 ;
        RECT 21.370 65.145 21.625 65.690 ;
        RECT 21.795 65.315 22.275 65.655 ;
        RECT 22.450 65.145 23.055 65.700 ;
        RECT 23.225 65.345 23.495 66.115 ;
        RECT 24.525 65.925 24.865 66.955 ;
        RECT 25.525 67.085 25.865 67.500 ;
        RECT 26.035 67.255 26.205 67.695 ;
        RECT 26.375 67.305 27.625 67.485 ;
        RECT 26.375 67.085 26.705 67.305 ;
        RECT 27.895 67.235 28.065 67.695 ;
        RECT 25.525 66.915 26.705 67.085 ;
        RECT 26.875 67.065 27.240 67.135 ;
        RECT 26.875 66.885 28.125 67.065 ;
        RECT 25.525 66.505 25.990 66.705 ;
        RECT 26.165 66.455 26.495 66.705 ;
        RECT 26.665 66.675 27.130 66.705 ;
        RECT 26.665 66.505 27.135 66.675 ;
        RECT 26.665 66.455 27.130 66.505 ;
        RECT 27.325 66.455 27.680 66.705 ;
        RECT 26.165 66.335 26.345 66.455 ;
        RECT 23.665 65.145 23.995 65.925 ;
        RECT 24.200 65.750 24.865 65.925 ;
        RECT 24.200 65.345 24.385 65.750 ;
        RECT 24.555 65.145 24.890 65.570 ;
        RECT 25.525 65.145 25.845 66.325 ;
        RECT 26.015 66.165 26.345 66.335 ;
        RECT 27.850 66.285 28.125 66.885 ;
        RECT 26.015 65.375 26.215 66.165 ;
        RECT 26.515 66.075 28.125 66.285 ;
        RECT 26.515 65.975 26.925 66.075 ;
        RECT 26.540 65.315 26.925 65.975 ;
        RECT 27.320 65.145 28.105 65.905 ;
        RECT 28.295 65.315 28.575 67.415 ;
        RECT 28.765 66.885 29.005 67.695 ;
        RECT 29.175 66.885 29.505 67.525 ;
        RECT 29.675 66.885 29.945 67.695 ;
        RECT 30.125 66.945 31.335 67.695 ;
        RECT 31.505 67.045 31.765 67.525 ;
        RECT 31.935 67.235 32.265 67.695 ;
        RECT 32.455 67.055 32.655 67.475 ;
        RECT 28.745 66.455 29.095 66.705 ;
        RECT 29.265 66.285 29.435 66.885 ;
        RECT 29.605 66.455 29.955 66.705 ;
        RECT 30.125 66.405 30.645 66.945 ;
        RECT 28.755 66.115 29.435 66.285 ;
        RECT 28.755 65.330 29.085 66.115 ;
        RECT 29.615 65.145 29.945 66.285 ;
        RECT 30.815 66.235 31.335 66.775 ;
        RECT 30.125 65.145 31.335 66.235 ;
        RECT 31.505 66.015 31.675 67.045 ;
        RECT 31.845 66.355 32.075 66.785 ;
        RECT 32.245 66.535 32.655 67.055 ;
        RECT 32.825 67.210 33.615 67.475 ;
        RECT 32.825 66.355 33.080 67.210 ;
        RECT 33.795 66.875 34.125 67.295 ;
        RECT 34.295 66.875 34.555 67.695 ;
        RECT 33.795 66.785 34.045 66.875 ;
        RECT 33.250 66.535 34.045 66.785 ;
        RECT 31.845 66.185 33.635 66.355 ;
        RECT 31.505 65.315 31.780 66.015 ;
        RECT 31.950 65.890 32.665 66.185 ;
        RECT 32.885 65.825 33.215 66.015 ;
        RECT 31.990 65.145 32.205 65.690 ;
        RECT 32.375 65.315 32.850 65.655 ;
        RECT 33.020 65.650 33.215 65.825 ;
        RECT 33.385 65.820 33.635 66.185 ;
        RECT 33.020 65.145 33.635 65.650 ;
        RECT 33.875 65.315 34.045 66.535 ;
        RECT 34.215 65.825 34.555 66.705 ;
        RECT 34.295 65.145 34.555 65.655 ;
        RECT 34.735 65.325 34.995 67.515 ;
        RECT 35.255 67.325 35.925 67.695 ;
        RECT 36.105 67.145 36.415 67.515 ;
        RECT 35.185 66.945 36.415 67.145 ;
        RECT 35.185 66.275 35.475 66.945 ;
        RECT 36.595 66.765 36.825 67.405 ;
        RECT 37.005 66.965 37.295 67.695 ;
        RECT 37.945 66.970 38.235 67.695 ;
        RECT 38.405 66.945 39.615 67.695 ;
        RECT 39.875 67.145 40.045 67.525 ;
        RECT 40.225 67.315 40.555 67.695 ;
        RECT 39.875 66.975 40.540 67.145 ;
        RECT 40.735 67.020 40.995 67.525 ;
        RECT 41.165 67.315 42.055 67.485 ;
        RECT 35.655 66.455 36.120 66.765 ;
        RECT 36.300 66.455 36.825 66.765 ;
        RECT 37.005 66.455 37.305 66.785 ;
        RECT 38.405 66.405 38.925 66.945 ;
        RECT 35.185 66.055 35.955 66.275 ;
        RECT 35.165 65.145 35.505 65.875 ;
        RECT 35.685 65.325 35.955 66.055 ;
        RECT 36.135 66.035 37.295 66.275 ;
        RECT 36.135 65.325 36.365 66.035 ;
        RECT 36.535 65.145 36.865 65.855 ;
        RECT 37.035 65.325 37.295 66.035 ;
        RECT 37.945 65.145 38.235 66.310 ;
        RECT 39.095 66.235 39.615 66.775 ;
        RECT 39.805 66.425 40.135 66.795 ;
        RECT 40.370 66.720 40.540 66.975 ;
        RECT 40.370 66.390 40.655 66.720 ;
        RECT 40.370 66.245 40.540 66.390 ;
        RECT 38.405 65.145 39.615 66.235 ;
        RECT 39.875 66.075 40.540 66.245 ;
        RECT 40.825 66.220 40.995 67.020 ;
        RECT 41.165 66.760 41.715 67.145 ;
        RECT 41.885 66.590 42.055 67.315 ;
        RECT 39.875 65.315 40.045 66.075 ;
        RECT 40.225 65.145 40.555 65.905 ;
        RECT 40.725 65.315 40.995 66.220 ;
        RECT 41.165 66.520 42.055 66.590 ;
        RECT 42.225 66.990 42.445 67.475 ;
        RECT 42.615 67.155 42.865 67.695 ;
        RECT 43.035 67.045 43.295 67.525 ;
        RECT 42.225 66.565 42.555 66.990 ;
        RECT 41.165 66.495 42.060 66.520 ;
        RECT 41.165 66.480 42.070 66.495 ;
        RECT 41.165 66.465 42.075 66.480 ;
        RECT 41.165 66.460 42.085 66.465 ;
        RECT 41.165 66.450 42.090 66.460 ;
        RECT 41.165 66.440 42.095 66.450 ;
        RECT 41.165 66.435 42.105 66.440 ;
        RECT 41.165 66.425 42.115 66.435 ;
        RECT 41.165 66.420 42.125 66.425 ;
        RECT 41.165 65.970 41.425 66.420 ;
        RECT 41.790 66.415 42.125 66.420 ;
        RECT 41.790 66.410 42.140 66.415 ;
        RECT 41.790 66.400 42.155 66.410 ;
        RECT 41.790 66.395 42.180 66.400 ;
        RECT 42.725 66.395 42.955 66.790 ;
        RECT 41.790 66.390 42.955 66.395 ;
        RECT 41.820 66.355 42.955 66.390 ;
        RECT 41.855 66.330 42.955 66.355 ;
        RECT 41.885 66.300 42.955 66.330 ;
        RECT 41.905 66.270 42.955 66.300 ;
        RECT 41.925 66.240 42.955 66.270 ;
        RECT 41.995 66.230 42.955 66.240 ;
        RECT 42.020 66.220 42.955 66.230 ;
        RECT 42.040 66.205 42.955 66.220 ;
        RECT 42.060 66.190 42.955 66.205 ;
        RECT 42.065 66.180 42.850 66.190 ;
        RECT 42.080 66.145 42.850 66.180 ;
        RECT 41.595 65.825 41.925 66.070 ;
        RECT 42.095 65.895 42.850 66.145 ;
        RECT 43.125 66.015 43.295 67.045 ;
        RECT 43.465 66.925 45.135 67.695 ;
        RECT 45.855 67.145 46.025 67.435 ;
        RECT 46.195 67.315 46.525 67.695 ;
        RECT 45.855 66.975 46.520 67.145 ;
        RECT 43.465 66.405 44.215 66.925 ;
        RECT 44.385 66.235 45.135 66.755 ;
        RECT 41.595 65.800 41.780 65.825 ;
        RECT 41.165 65.700 41.780 65.800 ;
        RECT 41.165 65.145 41.770 65.700 ;
        RECT 41.945 65.315 42.425 65.655 ;
        RECT 42.595 65.145 42.850 65.690 ;
        RECT 43.020 65.315 43.295 66.015 ;
        RECT 43.465 65.145 45.135 66.235 ;
        RECT 45.770 66.155 46.120 66.805 ;
        RECT 46.290 65.985 46.520 66.975 ;
        RECT 45.855 65.815 46.520 65.985 ;
        RECT 45.855 65.315 46.025 65.815 ;
        RECT 46.195 65.145 46.525 65.645 ;
        RECT 46.695 65.315 46.880 67.435 ;
        RECT 47.135 67.235 47.385 67.695 ;
        RECT 47.555 67.245 47.890 67.415 ;
        RECT 48.085 67.245 48.760 67.415 ;
        RECT 47.555 67.105 47.725 67.245 ;
        RECT 47.050 66.115 47.330 67.065 ;
        RECT 47.500 66.975 47.725 67.105 ;
        RECT 47.500 65.870 47.670 66.975 ;
        RECT 47.895 66.825 48.420 67.045 ;
        RECT 47.840 66.060 48.080 66.655 ;
        RECT 48.250 66.125 48.420 66.825 ;
        RECT 48.590 66.465 48.760 67.245 ;
        RECT 49.080 67.195 49.450 67.695 ;
        RECT 49.630 67.245 50.035 67.415 ;
        RECT 50.205 67.245 50.990 67.415 ;
        RECT 49.630 67.015 49.800 67.245 ;
        RECT 48.970 66.715 49.800 67.015 ;
        RECT 50.185 66.745 50.650 67.075 ;
        RECT 48.970 66.685 49.170 66.715 ;
        RECT 49.290 66.465 49.460 66.535 ;
        RECT 48.590 66.295 49.460 66.465 ;
        RECT 48.950 66.205 49.460 66.295 ;
        RECT 47.500 65.740 47.805 65.870 ;
        RECT 48.250 65.760 48.780 66.125 ;
        RECT 47.120 65.145 47.385 65.605 ;
        RECT 47.555 65.315 47.805 65.740 ;
        RECT 48.950 65.590 49.120 66.205 ;
        RECT 48.015 65.420 49.120 65.590 ;
        RECT 49.290 65.145 49.460 65.945 ;
        RECT 49.630 65.645 49.800 66.715 ;
        RECT 49.970 65.815 50.160 66.535 ;
        RECT 50.330 65.785 50.650 66.745 ;
        RECT 50.820 66.785 50.990 67.245 ;
        RECT 51.265 67.165 51.475 67.695 ;
        RECT 51.735 66.955 52.065 67.480 ;
        RECT 52.235 67.085 52.405 67.695 ;
        RECT 52.575 67.040 52.905 67.475 ;
        RECT 53.145 67.185 53.385 67.695 ;
        RECT 52.575 66.955 52.955 67.040 ;
        RECT 51.865 66.785 52.065 66.955 ;
        RECT 52.730 66.915 52.955 66.955 ;
        RECT 50.820 66.455 51.695 66.785 ;
        RECT 51.865 66.455 52.615 66.785 ;
        RECT 49.630 65.315 49.880 65.645 ;
        RECT 50.820 65.615 50.990 66.455 ;
        RECT 51.865 66.250 52.055 66.455 ;
        RECT 52.785 66.335 52.955 66.915 ;
        RECT 53.130 66.455 53.385 67.015 ;
        RECT 53.555 66.955 53.885 67.490 ;
        RECT 54.100 66.955 54.270 67.695 ;
        RECT 54.480 67.045 54.810 67.515 ;
        RECT 54.980 67.215 55.150 67.695 ;
        RECT 55.320 67.045 55.650 67.515 ;
        RECT 55.820 67.215 55.990 67.695 ;
        RECT 52.740 66.285 52.955 66.335 ;
        RECT 53.555 66.285 53.735 66.955 ;
        RECT 54.480 66.875 56.175 67.045 ;
        RECT 56.395 67.040 56.725 67.475 ;
        RECT 56.895 67.085 57.065 67.695 ;
        RECT 53.905 66.455 54.280 66.785 ;
        RECT 54.450 66.535 55.660 66.705 ;
        RECT 54.450 66.285 54.655 66.535 ;
        RECT 55.830 66.285 56.175 66.875 ;
        RECT 51.160 65.875 52.055 66.250 ;
        RECT 52.565 66.205 52.955 66.285 ;
        RECT 50.105 65.445 50.990 65.615 ;
        RECT 51.170 65.145 51.485 65.645 ;
        RECT 51.715 65.315 52.055 65.875 ;
        RECT 52.225 65.145 52.395 66.155 ;
        RECT 52.565 65.360 52.895 66.205 ;
        RECT 53.195 66.115 54.655 66.285 ;
        RECT 55.320 66.115 56.175 66.285 ;
        RECT 56.345 66.955 56.725 67.040 ;
        RECT 57.235 66.955 57.565 67.480 ;
        RECT 57.825 67.165 58.035 67.695 ;
        RECT 58.310 67.245 59.095 67.415 ;
        RECT 59.265 67.245 59.670 67.415 ;
        RECT 56.345 66.915 56.570 66.955 ;
        RECT 56.345 66.335 56.515 66.915 ;
        RECT 57.235 66.785 57.435 66.955 ;
        RECT 58.310 66.785 58.480 67.245 ;
        RECT 56.685 66.455 57.435 66.785 ;
        RECT 57.605 66.455 58.480 66.785 ;
        RECT 56.345 66.285 56.560 66.335 ;
        RECT 56.345 66.205 56.735 66.285 ;
        RECT 53.195 65.315 53.555 66.115 ;
        RECT 55.320 65.945 55.650 66.115 ;
        RECT 54.100 65.145 54.270 65.945 ;
        RECT 54.480 65.775 55.650 65.945 ;
        RECT 54.480 65.315 54.810 65.775 ;
        RECT 54.980 65.145 55.150 65.605 ;
        RECT 55.320 65.315 55.650 65.775 ;
        RECT 55.820 65.145 55.990 65.945 ;
        RECT 56.405 65.360 56.735 66.205 ;
        RECT 57.245 66.250 57.435 66.455 ;
        RECT 56.905 65.145 57.075 66.155 ;
        RECT 57.245 65.875 58.140 66.250 ;
        RECT 57.245 65.315 57.585 65.875 ;
        RECT 57.815 65.145 58.130 65.645 ;
        RECT 58.310 65.615 58.480 66.455 ;
        RECT 58.650 66.745 59.115 67.075 ;
        RECT 59.500 67.015 59.670 67.245 ;
        RECT 59.850 67.195 60.220 67.695 ;
        RECT 60.540 67.245 61.215 67.415 ;
        RECT 61.410 67.245 61.745 67.415 ;
        RECT 58.650 65.785 58.970 66.745 ;
        RECT 59.500 66.715 60.330 67.015 ;
        RECT 59.140 65.815 59.330 66.535 ;
        RECT 59.500 65.645 59.670 66.715 ;
        RECT 60.130 66.685 60.330 66.715 ;
        RECT 59.840 66.465 60.010 66.535 ;
        RECT 60.540 66.465 60.710 67.245 ;
        RECT 61.575 67.105 61.745 67.245 ;
        RECT 61.915 67.235 62.165 67.695 ;
        RECT 59.840 66.295 60.710 66.465 ;
        RECT 60.880 66.825 61.405 67.045 ;
        RECT 61.575 66.975 61.800 67.105 ;
        RECT 59.840 66.205 60.350 66.295 ;
        RECT 58.310 65.445 59.195 65.615 ;
        RECT 59.420 65.315 59.670 65.645 ;
        RECT 59.840 65.145 60.010 65.945 ;
        RECT 60.180 65.590 60.350 66.205 ;
        RECT 60.880 66.125 61.050 66.825 ;
        RECT 60.520 65.760 61.050 66.125 ;
        RECT 61.220 66.060 61.460 66.655 ;
        RECT 61.630 65.870 61.800 66.975 ;
        RECT 61.970 66.115 62.250 67.065 ;
        RECT 61.495 65.740 61.800 65.870 ;
        RECT 60.180 65.420 61.285 65.590 ;
        RECT 61.495 65.315 61.745 65.740 ;
        RECT 61.915 65.145 62.180 65.605 ;
        RECT 62.420 65.315 62.605 67.435 ;
        RECT 62.775 67.315 63.105 67.695 ;
        RECT 63.275 67.145 63.445 67.435 ;
        RECT 62.780 66.975 63.445 67.145 ;
        RECT 62.780 65.985 63.010 66.975 ;
        RECT 63.705 66.970 63.995 67.695 ;
        RECT 64.165 66.925 66.755 67.695 ;
        RECT 67.015 67.145 67.185 67.435 ;
        RECT 67.355 67.315 67.685 67.695 ;
        RECT 67.015 66.975 67.680 67.145 ;
        RECT 63.180 66.155 63.530 66.805 ;
        RECT 64.165 66.405 65.375 66.925 ;
        RECT 62.780 65.815 63.445 65.985 ;
        RECT 62.775 65.145 63.105 65.645 ;
        RECT 63.275 65.315 63.445 65.815 ;
        RECT 63.705 65.145 63.995 66.310 ;
        RECT 65.545 66.235 66.755 66.755 ;
        RECT 64.165 65.145 66.755 66.235 ;
        RECT 66.930 66.155 67.280 66.805 ;
        RECT 67.450 65.985 67.680 66.975 ;
        RECT 67.015 65.815 67.680 65.985 ;
        RECT 67.015 65.315 67.185 65.815 ;
        RECT 67.355 65.145 67.685 65.645 ;
        RECT 67.855 65.315 68.040 67.435 ;
        RECT 68.295 67.235 68.545 67.695 ;
        RECT 68.715 67.245 69.050 67.415 ;
        RECT 69.245 67.245 69.920 67.415 ;
        RECT 68.715 67.105 68.885 67.245 ;
        RECT 68.210 66.115 68.490 67.065 ;
        RECT 68.660 66.975 68.885 67.105 ;
        RECT 68.660 65.870 68.830 66.975 ;
        RECT 69.055 66.825 69.580 67.045 ;
        RECT 69.000 66.060 69.240 66.655 ;
        RECT 69.410 66.125 69.580 66.825 ;
        RECT 69.750 66.465 69.920 67.245 ;
        RECT 70.240 67.195 70.610 67.695 ;
        RECT 70.790 67.245 71.195 67.415 ;
        RECT 71.365 67.245 72.150 67.415 ;
        RECT 70.790 67.015 70.960 67.245 ;
        RECT 70.130 66.715 70.960 67.015 ;
        RECT 71.345 66.745 71.810 67.075 ;
        RECT 70.130 66.685 70.330 66.715 ;
        RECT 70.450 66.465 70.620 66.535 ;
        RECT 69.750 66.295 70.620 66.465 ;
        RECT 70.110 66.205 70.620 66.295 ;
        RECT 68.660 65.740 68.965 65.870 ;
        RECT 69.410 65.760 69.940 66.125 ;
        RECT 68.280 65.145 68.545 65.605 ;
        RECT 68.715 65.315 68.965 65.740 ;
        RECT 70.110 65.590 70.280 66.205 ;
        RECT 69.175 65.420 70.280 65.590 ;
        RECT 70.450 65.145 70.620 65.945 ;
        RECT 70.790 65.645 70.960 66.715 ;
        RECT 71.130 65.815 71.320 66.535 ;
        RECT 71.490 65.785 71.810 66.745 ;
        RECT 71.980 66.785 72.150 67.245 ;
        RECT 72.425 67.165 72.635 67.695 ;
        RECT 72.895 66.955 73.225 67.480 ;
        RECT 73.395 67.085 73.565 67.695 ;
        RECT 73.735 67.040 74.065 67.475 ;
        RECT 73.735 66.955 74.115 67.040 ;
        RECT 73.025 66.785 73.225 66.955 ;
        RECT 73.890 66.915 74.115 66.955 ;
        RECT 71.980 66.455 72.855 66.785 ;
        RECT 73.025 66.455 73.775 66.785 ;
        RECT 70.790 65.315 71.040 65.645 ;
        RECT 71.980 65.615 72.150 66.455 ;
        RECT 73.025 66.250 73.215 66.455 ;
        RECT 73.945 66.335 74.115 66.915 ;
        RECT 74.290 66.855 74.550 67.695 ;
        RECT 74.725 66.950 74.980 67.525 ;
        RECT 75.150 67.315 75.480 67.695 ;
        RECT 75.695 67.145 75.865 67.525 ;
        RECT 75.150 66.975 75.865 67.145 ;
        RECT 76.325 67.065 76.655 67.425 ;
        RECT 77.275 67.235 77.525 67.695 ;
        RECT 77.695 67.235 78.255 67.525 ;
        RECT 73.900 66.285 74.115 66.335 ;
        RECT 72.320 65.875 73.215 66.250 ;
        RECT 73.725 66.205 74.115 66.285 ;
        RECT 71.265 65.445 72.150 65.615 ;
        RECT 72.330 65.145 72.645 65.645 ;
        RECT 72.875 65.315 73.215 65.875 ;
        RECT 73.385 65.145 73.555 66.155 ;
        RECT 73.725 65.360 74.055 66.205 ;
        RECT 74.290 65.145 74.550 66.295 ;
        RECT 74.725 66.220 74.895 66.950 ;
        RECT 75.150 66.785 75.320 66.975 ;
        RECT 76.325 66.875 77.715 67.065 ;
        RECT 75.065 66.455 75.320 66.785 ;
        RECT 75.150 66.245 75.320 66.455 ;
        RECT 75.600 66.425 75.955 66.795 ;
        RECT 77.545 66.785 77.715 66.875 ;
        RECT 76.140 66.455 76.815 66.705 ;
        RECT 77.035 66.455 77.375 66.705 ;
        RECT 77.545 66.455 77.835 66.785 ;
        RECT 74.725 65.315 74.980 66.220 ;
        RECT 75.150 66.075 75.865 66.245 ;
        RECT 76.140 66.095 76.405 66.455 ;
        RECT 77.545 66.205 77.715 66.455 ;
        RECT 75.150 65.145 75.480 65.905 ;
        RECT 75.695 65.315 75.865 66.075 ;
        RECT 76.775 66.035 77.715 66.205 ;
        RECT 76.325 65.145 76.605 65.815 ;
        RECT 76.775 65.485 77.075 66.035 ;
        RECT 78.005 65.865 78.255 67.235 ;
        RECT 78.590 67.185 78.830 67.695 ;
        RECT 79.010 67.185 79.290 67.515 ;
        RECT 79.520 67.185 79.735 67.695 ;
        RECT 78.485 66.455 78.840 67.015 ;
        RECT 79.010 66.285 79.180 67.185 ;
        RECT 79.350 66.455 79.615 67.015 ;
        RECT 79.905 66.955 80.520 67.525 ;
        RECT 81.275 67.145 81.445 67.435 ;
        RECT 81.615 67.315 81.945 67.695 ;
        RECT 81.275 66.975 81.940 67.145 ;
        RECT 79.865 66.285 80.035 66.785 ;
        RECT 78.610 66.115 80.035 66.285 ;
        RECT 78.610 65.940 79.000 66.115 ;
        RECT 77.275 65.145 77.605 65.865 ;
        RECT 77.795 65.315 78.255 65.865 ;
        RECT 79.485 65.145 79.815 65.945 ;
        RECT 80.205 65.935 80.520 66.955 ;
        RECT 81.190 66.155 81.540 66.805 ;
        RECT 81.710 65.985 81.940 66.975 ;
        RECT 79.985 65.315 80.520 65.935 ;
        RECT 81.275 65.815 81.940 65.985 ;
        RECT 81.275 65.315 81.445 65.815 ;
        RECT 81.615 65.145 81.945 65.645 ;
        RECT 82.115 65.315 82.300 67.435 ;
        RECT 82.555 67.235 82.805 67.695 ;
        RECT 82.975 67.245 83.310 67.415 ;
        RECT 83.505 67.245 84.180 67.415 ;
        RECT 82.975 67.105 83.145 67.245 ;
        RECT 82.470 66.115 82.750 67.065 ;
        RECT 82.920 66.975 83.145 67.105 ;
        RECT 82.920 65.870 83.090 66.975 ;
        RECT 83.315 66.825 83.840 67.045 ;
        RECT 83.260 66.060 83.500 66.655 ;
        RECT 83.670 66.125 83.840 66.825 ;
        RECT 84.010 66.465 84.180 67.245 ;
        RECT 84.500 67.195 84.870 67.695 ;
        RECT 85.050 67.245 85.455 67.415 ;
        RECT 85.625 67.245 86.410 67.415 ;
        RECT 85.050 67.015 85.220 67.245 ;
        RECT 84.390 66.715 85.220 67.015 ;
        RECT 85.605 66.745 86.070 67.075 ;
        RECT 84.390 66.685 84.590 66.715 ;
        RECT 84.710 66.465 84.880 66.535 ;
        RECT 84.010 66.295 84.880 66.465 ;
        RECT 84.370 66.205 84.880 66.295 ;
        RECT 82.920 65.740 83.225 65.870 ;
        RECT 83.670 65.760 84.200 66.125 ;
        RECT 82.540 65.145 82.805 65.605 ;
        RECT 82.975 65.315 83.225 65.740 ;
        RECT 84.370 65.590 84.540 66.205 ;
        RECT 83.435 65.420 84.540 65.590 ;
        RECT 84.710 65.145 84.880 65.945 ;
        RECT 85.050 65.645 85.220 66.715 ;
        RECT 85.390 65.815 85.580 66.535 ;
        RECT 85.750 65.785 86.070 66.745 ;
        RECT 86.240 66.785 86.410 67.245 ;
        RECT 86.685 67.165 86.895 67.695 ;
        RECT 87.155 66.955 87.485 67.480 ;
        RECT 87.655 67.085 87.825 67.695 ;
        RECT 87.995 67.040 88.325 67.475 ;
        RECT 87.995 66.955 88.375 67.040 ;
        RECT 87.285 66.785 87.485 66.955 ;
        RECT 88.150 66.915 88.375 66.955 ;
        RECT 88.545 66.945 89.755 67.695 ;
        RECT 86.240 66.455 87.115 66.785 ;
        RECT 87.285 66.455 88.035 66.785 ;
        RECT 85.050 65.315 85.300 65.645 ;
        RECT 86.240 65.615 86.410 66.455 ;
        RECT 87.285 66.250 87.475 66.455 ;
        RECT 88.205 66.335 88.375 66.915 ;
        RECT 88.160 66.285 88.375 66.335 ;
        RECT 86.580 65.875 87.475 66.250 ;
        RECT 87.985 66.205 88.375 66.285 ;
        RECT 88.545 66.235 89.065 66.775 ;
        RECT 89.235 66.405 89.755 66.945 ;
        RECT 85.525 65.445 86.410 65.615 ;
        RECT 86.590 65.145 86.905 65.645 ;
        RECT 87.135 65.315 87.475 65.875 ;
        RECT 87.645 65.145 87.815 66.155 ;
        RECT 87.985 65.360 88.315 66.205 ;
        RECT 88.545 65.145 89.755 66.235 ;
        RECT 12.100 64.975 89.840 65.145 ;
        RECT 12.185 63.885 13.395 64.975 ;
        RECT 13.655 64.305 13.825 64.805 ;
        RECT 13.995 64.475 14.325 64.975 ;
        RECT 13.655 64.135 14.320 64.305 ;
        RECT 12.185 63.175 12.705 63.715 ;
        RECT 12.875 63.345 13.395 63.885 ;
        RECT 13.570 63.315 13.920 63.965 ;
        RECT 12.185 62.425 13.395 63.175 ;
        RECT 14.090 63.145 14.320 64.135 ;
        RECT 13.655 62.975 14.320 63.145 ;
        RECT 13.655 62.685 13.825 62.975 ;
        RECT 13.995 62.425 14.325 62.805 ;
        RECT 14.495 62.685 14.680 64.805 ;
        RECT 14.920 64.515 15.185 64.975 ;
        RECT 15.355 64.380 15.605 64.805 ;
        RECT 15.815 64.530 16.920 64.700 ;
        RECT 15.300 64.250 15.605 64.380 ;
        RECT 14.850 63.055 15.130 64.005 ;
        RECT 15.300 63.145 15.470 64.250 ;
        RECT 15.640 63.465 15.880 64.060 ;
        RECT 16.050 63.995 16.580 64.360 ;
        RECT 16.050 63.295 16.220 63.995 ;
        RECT 16.750 63.915 16.920 64.530 ;
        RECT 17.090 64.175 17.260 64.975 ;
        RECT 17.430 64.475 17.680 64.805 ;
        RECT 17.905 64.505 18.790 64.675 ;
        RECT 16.750 63.825 17.260 63.915 ;
        RECT 15.300 63.015 15.525 63.145 ;
        RECT 15.695 63.075 16.220 63.295 ;
        RECT 16.390 63.655 17.260 63.825 ;
        RECT 14.935 62.425 15.185 62.885 ;
        RECT 15.355 62.875 15.525 63.015 ;
        RECT 16.390 62.875 16.560 63.655 ;
        RECT 17.090 63.585 17.260 63.655 ;
        RECT 16.770 63.405 16.970 63.435 ;
        RECT 17.430 63.405 17.600 64.475 ;
        RECT 17.770 63.585 17.960 64.305 ;
        RECT 16.770 63.105 17.600 63.405 ;
        RECT 18.130 63.375 18.450 64.335 ;
        RECT 15.355 62.705 15.690 62.875 ;
        RECT 15.885 62.705 16.560 62.875 ;
        RECT 16.880 62.425 17.250 62.925 ;
        RECT 17.430 62.875 17.600 63.105 ;
        RECT 17.985 63.045 18.450 63.375 ;
        RECT 18.620 63.665 18.790 64.505 ;
        RECT 18.970 64.475 19.285 64.975 ;
        RECT 19.515 64.245 19.855 64.805 ;
        RECT 18.960 63.870 19.855 64.245 ;
        RECT 20.025 63.965 20.195 64.975 ;
        RECT 19.665 63.665 19.855 63.870 ;
        RECT 20.365 63.915 20.695 64.760 ;
        RECT 20.935 64.005 21.265 64.790 ;
        RECT 20.365 63.835 20.755 63.915 ;
        RECT 20.935 63.835 21.615 64.005 ;
        RECT 21.795 63.835 22.125 64.975 ;
        RECT 22.305 63.885 24.895 64.975 ;
        RECT 20.540 63.785 20.755 63.835 ;
        RECT 18.620 63.335 19.495 63.665 ;
        RECT 19.665 63.335 20.415 63.665 ;
        RECT 18.620 62.875 18.790 63.335 ;
        RECT 19.665 63.165 19.865 63.335 ;
        RECT 20.585 63.205 20.755 63.785 ;
        RECT 20.925 63.415 21.275 63.665 ;
        RECT 21.445 63.235 21.615 63.835 ;
        RECT 21.785 63.415 22.135 63.665 ;
        RECT 20.530 63.165 20.755 63.205 ;
        RECT 17.430 62.705 17.835 62.875 ;
        RECT 18.005 62.705 18.790 62.875 ;
        RECT 19.065 62.425 19.275 62.955 ;
        RECT 19.535 62.640 19.865 63.165 ;
        RECT 20.375 63.080 20.755 63.165 ;
        RECT 20.035 62.425 20.205 63.035 ;
        RECT 20.375 62.645 20.705 63.080 ;
        RECT 20.945 62.425 21.185 63.235 ;
        RECT 21.355 62.595 21.685 63.235 ;
        RECT 21.855 62.425 22.125 63.235 ;
        RECT 22.305 63.195 23.515 63.715 ;
        RECT 23.685 63.365 24.895 63.885 ;
        RECT 25.065 63.810 25.355 64.975 ;
        RECT 25.525 63.885 28.115 64.975 ;
        RECT 25.525 63.195 26.735 63.715 ;
        RECT 26.905 63.365 28.115 63.885 ;
        RECT 28.285 63.835 28.545 64.975 ;
        RECT 28.715 63.825 29.045 64.805 ;
        RECT 29.215 63.835 29.495 64.975 ;
        RECT 29.665 63.835 29.945 64.975 ;
        RECT 30.115 63.825 30.445 64.805 ;
        RECT 30.615 63.835 30.875 64.975 ;
        RECT 31.045 63.885 32.715 64.975 ;
        RECT 28.305 63.415 28.640 63.665 ;
        RECT 28.810 63.225 28.980 63.825 ;
        RECT 30.180 63.785 30.355 63.825 ;
        RECT 29.150 63.395 29.485 63.665 ;
        RECT 29.675 63.395 30.010 63.665 ;
        RECT 30.180 63.225 30.350 63.785 ;
        RECT 30.520 63.415 30.855 63.665 ;
        RECT 22.305 62.425 24.895 63.195 ;
        RECT 25.065 62.425 25.355 63.150 ;
        RECT 25.525 62.425 28.115 63.195 ;
        RECT 28.285 62.595 28.980 63.225 ;
        RECT 29.185 62.425 29.495 63.225 ;
        RECT 29.665 62.425 29.975 63.225 ;
        RECT 30.180 62.595 30.875 63.225 ;
        RECT 31.045 63.195 31.795 63.715 ;
        RECT 31.965 63.365 32.715 63.885 ;
        RECT 32.885 64.105 33.160 64.805 ;
        RECT 33.330 64.430 33.585 64.975 ;
        RECT 33.755 64.465 34.235 64.805 ;
        RECT 34.410 64.420 35.015 64.975 ;
        RECT 35.185 64.540 40.530 64.975 ;
        RECT 40.705 64.540 46.050 64.975 ;
        RECT 34.400 64.320 35.015 64.420 ;
        RECT 34.400 64.295 34.585 64.320 ;
        RECT 31.045 62.425 32.715 63.195 ;
        RECT 32.885 63.075 33.055 64.105 ;
        RECT 33.330 63.975 34.085 64.225 ;
        RECT 34.255 64.050 34.585 64.295 ;
        RECT 33.330 63.940 34.100 63.975 ;
        RECT 33.330 63.930 34.115 63.940 ;
        RECT 33.225 63.915 34.120 63.930 ;
        RECT 33.225 63.900 34.140 63.915 ;
        RECT 33.225 63.890 34.160 63.900 ;
        RECT 33.225 63.880 34.185 63.890 ;
        RECT 33.225 63.850 34.255 63.880 ;
        RECT 33.225 63.820 34.275 63.850 ;
        RECT 33.225 63.790 34.295 63.820 ;
        RECT 33.225 63.765 34.325 63.790 ;
        RECT 33.225 63.730 34.360 63.765 ;
        RECT 33.225 63.725 34.390 63.730 ;
        RECT 33.225 63.330 33.455 63.725 ;
        RECT 34.000 63.720 34.390 63.725 ;
        RECT 34.025 63.710 34.390 63.720 ;
        RECT 34.040 63.705 34.390 63.710 ;
        RECT 34.055 63.700 34.390 63.705 ;
        RECT 34.755 63.700 35.015 64.150 ;
        RECT 34.055 63.695 35.015 63.700 ;
        RECT 34.065 63.685 35.015 63.695 ;
        RECT 34.075 63.680 35.015 63.685 ;
        RECT 34.085 63.670 35.015 63.680 ;
        RECT 34.090 63.660 35.015 63.670 ;
        RECT 34.095 63.655 35.015 63.660 ;
        RECT 34.105 63.640 35.015 63.655 ;
        RECT 34.110 63.625 35.015 63.640 ;
        RECT 34.120 63.600 35.015 63.625 ;
        RECT 33.625 63.130 33.955 63.555 ;
        RECT 32.885 62.595 33.145 63.075 ;
        RECT 33.315 62.425 33.565 62.965 ;
        RECT 33.735 62.645 33.955 63.130 ;
        RECT 34.125 63.530 35.015 63.600 ;
        RECT 34.125 62.805 34.295 63.530 ;
        RECT 34.465 62.975 35.015 63.360 ;
        RECT 36.770 62.970 37.110 63.800 ;
        RECT 38.590 63.290 38.940 64.540 ;
        RECT 42.290 62.970 42.630 63.800 ;
        RECT 44.110 63.290 44.460 64.540 ;
        RECT 46.225 63.885 47.895 64.975 ;
        RECT 48.525 64.420 49.130 64.975 ;
        RECT 49.305 64.465 49.785 64.805 ;
        RECT 49.955 64.430 50.210 64.975 ;
        RECT 48.525 64.320 49.140 64.420 ;
        RECT 48.955 64.295 49.140 64.320 ;
        RECT 46.225 63.195 46.975 63.715 ;
        RECT 47.145 63.365 47.895 63.885 ;
        RECT 48.525 63.700 48.785 64.150 ;
        RECT 48.955 64.050 49.285 64.295 ;
        RECT 49.455 63.975 50.210 64.225 ;
        RECT 50.380 64.105 50.655 64.805 ;
        RECT 49.440 63.940 50.210 63.975 ;
        RECT 49.425 63.930 50.210 63.940 ;
        RECT 49.420 63.915 50.315 63.930 ;
        RECT 49.400 63.900 50.315 63.915 ;
        RECT 49.380 63.890 50.315 63.900 ;
        RECT 49.355 63.880 50.315 63.890 ;
        RECT 49.285 63.850 50.315 63.880 ;
        RECT 49.265 63.820 50.315 63.850 ;
        RECT 49.245 63.790 50.315 63.820 ;
        RECT 49.215 63.765 50.315 63.790 ;
        RECT 49.180 63.730 50.315 63.765 ;
        RECT 49.150 63.725 50.315 63.730 ;
        RECT 49.150 63.720 49.540 63.725 ;
        RECT 49.150 63.710 49.515 63.720 ;
        RECT 49.150 63.705 49.500 63.710 ;
        RECT 49.150 63.700 49.485 63.705 ;
        RECT 48.525 63.695 49.485 63.700 ;
        RECT 48.525 63.685 49.475 63.695 ;
        RECT 48.525 63.680 49.465 63.685 ;
        RECT 48.525 63.670 49.455 63.680 ;
        RECT 48.525 63.660 49.450 63.670 ;
        RECT 48.525 63.655 49.445 63.660 ;
        RECT 48.525 63.640 49.435 63.655 ;
        RECT 48.525 63.625 49.430 63.640 ;
        RECT 48.525 63.600 49.420 63.625 ;
        RECT 48.525 63.530 49.415 63.600 ;
        RECT 34.125 62.635 35.015 62.805 ;
        RECT 35.185 62.425 40.530 62.970 ;
        RECT 40.705 62.425 46.050 62.970 ;
        RECT 46.225 62.425 47.895 63.195 ;
        RECT 48.525 62.975 49.075 63.360 ;
        RECT 49.245 62.805 49.415 63.530 ;
        RECT 48.525 62.635 49.415 62.805 ;
        RECT 49.585 63.130 49.915 63.555 ;
        RECT 50.085 63.330 50.315 63.725 ;
        RECT 49.585 62.645 49.805 63.130 ;
        RECT 50.485 63.075 50.655 64.105 ;
        RECT 50.825 63.810 51.115 64.975 ;
        RECT 51.285 64.465 52.485 64.705 ;
        RECT 52.665 64.550 52.995 64.975 ;
        RECT 53.510 64.550 53.870 64.975 ;
        RECT 54.075 64.380 54.335 64.560 ;
        RECT 52.700 64.295 54.335 64.380 ;
        RECT 54.505 64.420 55.110 64.975 ;
        RECT 55.285 64.465 55.765 64.805 ;
        RECT 55.935 64.430 56.190 64.975 ;
        RECT 54.505 64.320 55.120 64.420 ;
        RECT 51.285 63.835 51.590 64.265 ;
        RECT 51.760 64.210 54.335 64.295 ;
        RECT 51.760 64.125 52.870 64.210 ;
        RECT 53.655 64.150 54.335 64.210 ;
        RECT 54.935 64.295 55.120 64.320 ;
        RECT 51.285 63.165 51.455 63.835 ;
        RECT 51.760 63.665 51.930 64.125 ;
        RECT 51.630 63.335 51.930 63.665 ;
        RECT 52.190 63.415 52.725 63.955 ;
        RECT 53.090 63.835 53.485 64.040 ;
        RECT 52.975 63.275 53.145 63.665 ;
        RECT 52.825 63.245 53.145 63.275 ;
        RECT 52.260 63.165 53.145 63.245 ;
        RECT 49.975 62.425 50.225 62.965 ;
        RECT 50.395 62.595 50.655 63.075 ;
        RECT 50.825 62.425 51.115 63.150 ;
        RECT 51.285 63.105 53.145 63.165 ;
        RECT 51.285 63.075 52.995 63.105 ;
        RECT 51.285 62.995 52.430 63.075 ;
        RECT 51.285 62.945 51.590 62.995 ;
        RECT 51.335 62.645 51.590 62.945 ;
        RECT 51.760 62.425 52.090 62.825 ;
        RECT 52.260 62.645 52.430 62.995 ;
        RECT 53.315 62.935 53.485 63.835 ;
        RECT 53.655 63.245 53.825 64.150 ;
        RECT 53.995 63.415 54.335 63.980 ;
        RECT 54.505 63.700 54.765 64.150 ;
        RECT 54.935 64.050 55.265 64.295 ;
        RECT 55.435 63.975 56.190 64.225 ;
        RECT 56.360 64.105 56.635 64.805 ;
        RECT 56.805 64.540 62.150 64.975 ;
        RECT 55.420 63.940 56.190 63.975 ;
        RECT 55.405 63.930 56.190 63.940 ;
        RECT 55.400 63.915 56.295 63.930 ;
        RECT 55.380 63.900 56.295 63.915 ;
        RECT 55.360 63.890 56.295 63.900 ;
        RECT 55.335 63.880 56.295 63.890 ;
        RECT 55.265 63.850 56.295 63.880 ;
        RECT 55.245 63.820 56.295 63.850 ;
        RECT 55.225 63.790 56.295 63.820 ;
        RECT 55.195 63.765 56.295 63.790 ;
        RECT 55.160 63.730 56.295 63.765 ;
        RECT 55.130 63.725 56.295 63.730 ;
        RECT 55.130 63.720 55.520 63.725 ;
        RECT 55.130 63.710 55.495 63.720 ;
        RECT 55.130 63.705 55.480 63.710 ;
        RECT 55.130 63.700 55.465 63.705 ;
        RECT 54.505 63.695 55.465 63.700 ;
        RECT 54.505 63.685 55.455 63.695 ;
        RECT 54.505 63.680 55.445 63.685 ;
        RECT 54.505 63.670 55.435 63.680 ;
        RECT 54.505 63.660 55.430 63.670 ;
        RECT 54.505 63.655 55.425 63.660 ;
        RECT 54.505 63.640 55.415 63.655 ;
        RECT 54.505 63.625 55.410 63.640 ;
        RECT 54.505 63.600 55.400 63.625 ;
        RECT 54.505 63.530 55.395 63.600 ;
        RECT 53.655 63.075 54.335 63.245 ;
        RECT 52.730 62.425 52.900 62.905 ;
        RECT 53.135 62.605 53.485 62.935 ;
        RECT 53.655 62.425 53.825 62.905 ;
        RECT 54.075 62.630 54.335 63.075 ;
        RECT 54.505 62.975 55.055 63.360 ;
        RECT 55.225 62.805 55.395 63.530 ;
        RECT 54.505 62.635 55.395 62.805 ;
        RECT 55.565 63.130 55.895 63.555 ;
        RECT 56.065 63.330 56.295 63.725 ;
        RECT 55.565 62.645 55.785 63.130 ;
        RECT 56.465 63.075 56.635 64.105 ;
        RECT 55.955 62.425 56.205 62.965 ;
        RECT 56.375 62.595 56.635 63.075 ;
        RECT 58.390 62.970 58.730 63.800 ;
        RECT 60.210 63.290 60.560 64.540 ;
        RECT 62.325 63.885 64.915 64.975 ;
        RECT 62.325 63.195 63.535 63.715 ;
        RECT 63.705 63.365 64.915 63.885 ;
        RECT 65.095 63.865 65.390 64.975 ;
        RECT 65.570 63.665 65.820 64.800 ;
        RECT 65.990 63.865 66.250 64.975 ;
        RECT 66.420 64.075 66.680 64.800 ;
        RECT 66.850 64.245 67.110 64.975 ;
        RECT 67.280 64.075 67.540 64.800 ;
        RECT 67.710 64.245 67.970 64.975 ;
        RECT 68.140 64.075 68.400 64.800 ;
        RECT 68.570 64.245 68.830 64.975 ;
        RECT 69.000 64.075 69.260 64.800 ;
        RECT 69.430 64.245 69.725 64.975 ;
        RECT 66.420 63.835 69.730 64.075 ;
        RECT 70.145 63.885 71.815 64.975 ;
        RECT 72.090 64.175 72.345 64.975 ;
        RECT 72.515 64.005 72.845 64.805 ;
        RECT 73.015 64.175 73.185 64.975 ;
        RECT 73.355 64.005 73.685 64.805 ;
        RECT 56.805 62.425 62.150 62.970 ;
        RECT 62.325 62.425 64.915 63.195 ;
        RECT 65.085 63.055 65.400 63.665 ;
        RECT 65.570 63.415 68.590 63.665 ;
        RECT 65.145 62.425 65.390 62.885 ;
        RECT 65.570 62.605 65.820 63.415 ;
        RECT 68.760 63.245 69.730 63.835 ;
        RECT 66.420 63.075 69.730 63.245 ;
        RECT 70.145 63.195 70.895 63.715 ;
        RECT 71.065 63.365 71.815 63.885 ;
        RECT 71.985 63.835 73.685 64.005 ;
        RECT 73.855 63.835 74.115 64.975 ;
        RECT 74.285 64.255 74.745 64.805 ;
        RECT 74.935 64.255 75.265 64.975 ;
        RECT 71.985 63.245 72.265 63.835 ;
        RECT 72.435 63.415 73.185 63.665 ;
        RECT 73.355 63.415 74.115 63.665 ;
        RECT 65.990 62.425 66.250 62.950 ;
        RECT 66.420 62.620 66.680 63.075 ;
        RECT 66.850 62.425 67.110 62.905 ;
        RECT 67.280 62.620 67.540 63.075 ;
        RECT 67.710 62.425 67.970 62.905 ;
        RECT 68.140 62.620 68.400 63.075 ;
        RECT 68.570 62.425 68.830 62.905 ;
        RECT 69.000 62.620 69.260 63.075 ;
        RECT 69.430 62.425 69.730 62.905 ;
        RECT 70.145 62.425 71.815 63.195 ;
        RECT 71.985 62.995 72.845 63.245 ;
        RECT 73.015 63.055 74.115 63.225 ;
        RECT 72.095 62.805 72.425 62.825 ;
        RECT 73.015 62.805 73.265 63.055 ;
        RECT 72.095 62.595 73.265 62.805 ;
        RECT 73.435 62.425 73.605 62.885 ;
        RECT 73.775 62.595 74.115 63.055 ;
        RECT 74.285 62.885 74.535 64.255 ;
        RECT 75.465 64.085 75.765 64.635 ;
        RECT 75.935 64.305 76.215 64.975 ;
        RECT 74.825 63.915 75.765 64.085 ;
        RECT 74.825 63.665 74.995 63.915 ;
        RECT 76.135 63.665 76.400 64.025 ;
        RECT 76.585 63.810 76.875 64.975 ;
        RECT 77.710 64.005 78.040 64.805 ;
        RECT 78.210 64.175 78.540 64.975 ;
        RECT 78.840 64.005 79.170 64.805 ;
        RECT 79.815 64.175 80.065 64.975 ;
        RECT 77.710 63.835 80.145 64.005 ;
        RECT 80.335 63.835 80.505 64.975 ;
        RECT 80.675 63.835 81.015 64.805 ;
        RECT 81.275 64.305 81.445 64.805 ;
        RECT 81.615 64.475 81.945 64.975 ;
        RECT 81.275 64.135 81.940 64.305 ;
        RECT 74.705 63.335 74.995 63.665 ;
        RECT 75.165 63.415 75.505 63.665 ;
        RECT 75.725 63.415 76.400 63.665 ;
        RECT 77.505 63.415 77.855 63.665 ;
        RECT 74.825 63.245 74.995 63.335 ;
        RECT 74.825 63.055 76.215 63.245 ;
        RECT 78.040 63.205 78.210 63.835 ;
        RECT 78.380 63.415 78.710 63.615 ;
        RECT 78.880 63.415 79.210 63.615 ;
        RECT 79.380 63.415 79.800 63.615 ;
        RECT 79.975 63.585 80.145 63.835 ;
        RECT 79.975 63.415 80.670 63.585 ;
        RECT 74.285 62.595 74.845 62.885 ;
        RECT 75.015 62.425 75.265 62.885 ;
        RECT 75.885 62.695 76.215 63.055 ;
        RECT 76.585 62.425 76.875 63.150 ;
        RECT 77.710 62.595 78.210 63.205 ;
        RECT 78.840 63.075 80.065 63.245 ;
        RECT 80.840 63.225 81.015 63.835 ;
        RECT 81.190 63.315 81.540 63.965 ;
        RECT 78.840 62.595 79.170 63.075 ;
        RECT 79.340 62.425 79.565 62.885 ;
        RECT 79.735 62.595 80.065 63.075 ;
        RECT 80.255 62.425 80.505 63.225 ;
        RECT 80.675 62.595 81.015 63.225 ;
        RECT 81.710 63.145 81.940 64.135 ;
        RECT 81.275 62.975 81.940 63.145 ;
        RECT 81.275 62.685 81.445 62.975 ;
        RECT 81.615 62.425 81.945 62.805 ;
        RECT 82.115 62.685 82.300 64.805 ;
        RECT 82.540 64.515 82.805 64.975 ;
        RECT 82.975 64.380 83.225 64.805 ;
        RECT 83.435 64.530 84.540 64.700 ;
        RECT 82.920 64.250 83.225 64.380 ;
        RECT 82.470 63.055 82.750 64.005 ;
        RECT 82.920 63.145 83.090 64.250 ;
        RECT 83.260 63.465 83.500 64.060 ;
        RECT 83.670 63.995 84.200 64.360 ;
        RECT 83.670 63.295 83.840 63.995 ;
        RECT 84.370 63.915 84.540 64.530 ;
        RECT 84.710 64.175 84.880 64.975 ;
        RECT 85.050 64.475 85.300 64.805 ;
        RECT 85.525 64.505 86.410 64.675 ;
        RECT 84.370 63.825 84.880 63.915 ;
        RECT 82.920 63.015 83.145 63.145 ;
        RECT 83.315 63.075 83.840 63.295 ;
        RECT 84.010 63.655 84.880 63.825 ;
        RECT 82.555 62.425 82.805 62.885 ;
        RECT 82.975 62.875 83.145 63.015 ;
        RECT 84.010 62.875 84.180 63.655 ;
        RECT 84.710 63.585 84.880 63.655 ;
        RECT 84.390 63.405 84.590 63.435 ;
        RECT 85.050 63.405 85.220 64.475 ;
        RECT 85.390 63.585 85.580 64.305 ;
        RECT 84.390 63.105 85.220 63.405 ;
        RECT 85.750 63.375 86.070 64.335 ;
        RECT 82.975 62.705 83.310 62.875 ;
        RECT 83.505 62.705 84.180 62.875 ;
        RECT 84.500 62.425 84.870 62.925 ;
        RECT 85.050 62.875 85.220 63.105 ;
        RECT 85.605 63.045 86.070 63.375 ;
        RECT 86.240 63.665 86.410 64.505 ;
        RECT 86.590 64.475 86.905 64.975 ;
        RECT 87.135 64.245 87.475 64.805 ;
        RECT 86.580 63.870 87.475 64.245 ;
        RECT 87.645 63.965 87.815 64.975 ;
        RECT 87.285 63.665 87.475 63.870 ;
        RECT 87.985 63.915 88.315 64.760 ;
        RECT 87.985 63.835 88.375 63.915 ;
        RECT 88.160 63.785 88.375 63.835 ;
        RECT 86.240 63.335 87.115 63.665 ;
        RECT 87.285 63.335 88.035 63.665 ;
        RECT 86.240 62.875 86.410 63.335 ;
        RECT 87.285 63.165 87.485 63.335 ;
        RECT 88.205 63.205 88.375 63.785 ;
        RECT 88.545 63.885 89.755 64.975 ;
        RECT 88.545 63.345 89.065 63.885 ;
        RECT 88.150 63.165 88.375 63.205 ;
        RECT 89.235 63.175 89.755 63.715 ;
        RECT 85.050 62.705 85.455 62.875 ;
        RECT 85.625 62.705 86.410 62.875 ;
        RECT 86.685 62.425 86.895 62.955 ;
        RECT 87.155 62.640 87.485 63.165 ;
        RECT 87.995 63.080 88.375 63.165 ;
        RECT 87.655 62.425 87.825 63.035 ;
        RECT 87.995 62.645 88.325 63.080 ;
        RECT 88.545 62.425 89.755 63.175 ;
        RECT 12.100 62.255 89.840 62.425 ;
        RECT 12.185 61.505 13.395 62.255 ;
        RECT 13.565 61.505 14.775 62.255 ;
        RECT 14.945 61.605 15.205 62.085 ;
        RECT 15.375 61.715 15.625 62.255 ;
        RECT 12.185 60.965 12.705 61.505 ;
        RECT 12.875 60.795 13.395 61.335 ;
        RECT 13.565 60.965 14.085 61.505 ;
        RECT 14.255 60.795 14.775 61.335 ;
        RECT 12.185 59.705 13.395 60.795 ;
        RECT 13.565 59.705 14.775 60.795 ;
        RECT 14.945 60.575 15.115 61.605 ;
        RECT 15.795 61.550 16.015 62.035 ;
        RECT 15.285 60.955 15.515 61.350 ;
        RECT 15.685 61.125 16.015 61.550 ;
        RECT 16.185 61.875 17.075 62.045 ;
        RECT 16.185 61.150 16.355 61.875 ;
        RECT 17.245 61.755 17.505 62.085 ;
        RECT 17.715 61.775 17.990 62.255 ;
        RECT 16.525 61.320 17.075 61.705 ;
        RECT 16.185 61.080 17.075 61.150 ;
        RECT 16.180 61.055 17.075 61.080 ;
        RECT 16.170 61.040 17.075 61.055 ;
        RECT 16.165 61.025 17.075 61.040 ;
        RECT 16.155 61.020 17.075 61.025 ;
        RECT 16.150 61.010 17.075 61.020 ;
        RECT 16.145 61.000 17.075 61.010 ;
        RECT 16.135 60.995 17.075 61.000 ;
        RECT 16.125 60.985 17.075 60.995 ;
        RECT 16.115 60.980 17.075 60.985 ;
        RECT 16.115 60.975 16.450 60.980 ;
        RECT 16.100 60.970 16.450 60.975 ;
        RECT 16.085 60.960 16.450 60.970 ;
        RECT 16.060 60.955 16.450 60.960 ;
        RECT 15.285 60.950 16.450 60.955 ;
        RECT 15.285 60.915 16.420 60.950 ;
        RECT 15.285 60.890 16.385 60.915 ;
        RECT 15.285 60.860 16.355 60.890 ;
        RECT 15.285 60.830 16.335 60.860 ;
        RECT 15.285 60.800 16.315 60.830 ;
        RECT 15.285 60.790 16.245 60.800 ;
        RECT 15.285 60.780 16.220 60.790 ;
        RECT 15.285 60.765 16.200 60.780 ;
        RECT 15.285 60.750 16.180 60.765 ;
        RECT 15.390 60.740 16.175 60.750 ;
        RECT 15.390 60.705 16.160 60.740 ;
        RECT 14.945 59.875 15.220 60.575 ;
        RECT 15.390 60.455 16.145 60.705 ;
        RECT 16.315 60.385 16.645 60.630 ;
        RECT 16.815 60.530 17.075 60.980 ;
        RECT 17.245 60.845 17.415 61.755 ;
        RECT 18.200 61.685 18.405 62.085 ;
        RECT 18.575 61.855 18.910 62.255 ;
        RECT 17.585 61.015 17.945 61.595 ;
        RECT 18.200 61.515 18.885 61.685 ;
        RECT 18.125 60.845 18.375 61.345 ;
        RECT 17.245 60.675 18.375 60.845 ;
        RECT 16.460 60.360 16.645 60.385 ;
        RECT 16.460 60.260 17.075 60.360 ;
        RECT 15.390 59.705 15.645 60.250 ;
        RECT 15.815 59.875 16.295 60.215 ;
        RECT 16.470 59.705 17.075 60.260 ;
        RECT 17.245 59.905 17.515 60.675 ;
        RECT 18.545 60.485 18.885 61.515 ;
        RECT 19.095 61.445 19.365 62.255 ;
        RECT 19.535 61.445 19.865 62.085 ;
        RECT 20.035 61.445 20.275 62.255 ;
        RECT 20.465 61.710 25.810 62.255 ;
        RECT 19.085 61.015 19.435 61.265 ;
        RECT 19.605 60.845 19.775 61.445 ;
        RECT 19.945 61.015 20.295 61.265 ;
        RECT 22.050 60.880 22.390 61.710 ;
        RECT 26.455 61.615 26.785 62.085 ;
        RECT 26.955 61.785 27.125 62.255 ;
        RECT 27.295 61.615 27.625 62.085 ;
        RECT 27.795 61.785 27.965 62.255 ;
        RECT 28.135 61.865 30.145 62.085 ;
        RECT 30.335 61.865 32.345 62.085 ;
        RECT 28.135 61.615 28.385 61.865 ;
        RECT 26.455 61.435 28.385 61.615 ;
        RECT 28.555 61.455 31.925 61.695 ;
        RECT 32.095 61.615 32.345 61.865 ;
        RECT 32.515 61.785 32.685 62.255 ;
        RECT 32.855 61.615 33.185 62.085 ;
        RECT 33.355 61.785 33.525 62.255 ;
        RECT 33.695 61.615 34.025 62.085 ;
        RECT 34.430 61.745 34.670 62.255 ;
        RECT 34.850 61.745 35.130 62.075 ;
        RECT 35.360 61.745 35.575 62.255 ;
        RECT 17.685 59.705 18.015 60.485 ;
        RECT 18.220 60.310 18.885 60.485 ;
        RECT 18.220 59.905 18.405 60.310 ;
        RECT 18.575 59.705 18.910 60.130 ;
        RECT 19.095 59.705 19.425 60.845 ;
        RECT 19.605 60.675 20.285 60.845 ;
        RECT 19.955 59.890 20.285 60.675 ;
        RECT 23.870 60.140 24.220 61.390 ;
        RECT 26.450 61.065 28.255 61.265 ;
        RECT 28.555 60.895 28.805 61.455 ;
        RECT 32.095 61.435 34.025 61.615 ;
        RECT 28.975 61.065 30.400 61.265 ;
        RECT 30.635 61.055 32.045 61.265 ;
        RECT 32.270 61.055 34.095 61.265 ;
        RECT 34.325 61.015 34.680 61.575 ;
        RECT 20.465 59.705 25.810 60.140 ;
        RECT 26.450 60.045 26.785 60.885 ;
        RECT 26.955 60.715 29.685 60.895 ;
        RECT 26.955 60.215 27.165 60.715 ;
        RECT 27.335 60.045 27.585 60.545 ;
        RECT 27.755 60.215 28.005 60.715 ;
        RECT 28.175 60.045 28.425 60.545 ;
        RECT 28.595 60.215 28.845 60.715 ;
        RECT 29.015 60.045 29.265 60.545 ;
        RECT 29.435 60.215 29.685 60.715 ;
        RECT 29.855 60.715 33.985 60.885 ;
        RECT 34.850 60.845 35.020 61.745 ;
        RECT 35.190 61.015 35.455 61.575 ;
        RECT 35.745 61.515 36.360 62.085 ;
        RECT 35.705 60.845 35.875 61.345 ;
        RECT 29.855 60.045 30.625 60.715 ;
        RECT 26.450 59.875 30.625 60.045 ;
        RECT 30.795 59.705 31.045 60.545 ;
        RECT 31.215 59.875 31.465 60.715 ;
        RECT 31.635 59.705 31.885 60.545 ;
        RECT 32.055 59.875 32.305 60.715 ;
        RECT 32.475 59.705 32.725 60.545 ;
        RECT 32.895 59.875 33.145 60.715 ;
        RECT 33.315 59.705 33.565 60.545 ;
        RECT 33.735 59.875 33.985 60.715 ;
        RECT 34.450 60.675 35.875 60.845 ;
        RECT 34.450 60.500 34.840 60.675 ;
        RECT 35.325 59.705 35.655 60.505 ;
        RECT 36.045 60.495 36.360 61.515 ;
        RECT 36.565 61.505 37.775 62.255 ;
        RECT 37.945 61.530 38.235 62.255 ;
        RECT 36.565 60.965 37.085 61.505 ;
        RECT 38.405 61.485 41.915 62.255 ;
        RECT 42.085 61.505 43.295 62.255 ;
        RECT 43.475 61.525 43.775 62.255 ;
        RECT 37.255 60.795 37.775 61.335 ;
        RECT 38.405 60.965 40.055 61.485 ;
        RECT 35.825 59.875 36.360 60.495 ;
        RECT 36.565 59.705 37.775 60.795 ;
        RECT 37.945 59.705 38.235 60.870 ;
        RECT 40.225 60.795 41.915 61.315 ;
        RECT 42.085 60.965 42.605 61.505 ;
        RECT 43.955 61.345 44.185 61.965 ;
        RECT 44.385 61.695 44.610 62.075 ;
        RECT 44.780 61.865 45.110 62.255 ;
        RECT 44.385 61.515 44.715 61.695 ;
        RECT 42.775 60.795 43.295 61.335 ;
        RECT 43.480 61.015 43.775 61.345 ;
        RECT 43.955 61.015 44.370 61.345 ;
        RECT 44.540 60.845 44.715 61.515 ;
        RECT 44.885 61.015 45.125 61.665 ;
        RECT 45.305 61.485 47.895 62.255 ;
        RECT 45.305 60.965 46.515 61.485 ;
        RECT 48.075 61.445 48.345 62.255 ;
        RECT 48.515 61.445 48.845 62.085 ;
        RECT 49.015 61.445 49.255 62.255 ;
        RECT 49.445 61.485 51.115 62.255 ;
        RECT 51.320 61.515 51.935 62.085 ;
        RECT 52.105 61.745 52.320 62.255 ;
        RECT 52.550 61.745 52.830 62.075 ;
        RECT 53.010 61.745 53.250 62.255 ;
        RECT 38.405 59.705 41.915 60.795 ;
        RECT 42.085 59.705 43.295 60.795 ;
        RECT 43.475 60.485 44.370 60.815 ;
        RECT 44.540 60.655 45.125 60.845 ;
        RECT 46.685 60.795 47.895 61.315 ;
        RECT 48.065 61.015 48.415 61.265 ;
        RECT 48.585 60.845 48.755 61.445 ;
        RECT 48.925 61.015 49.275 61.265 ;
        RECT 49.445 60.965 50.195 61.485 ;
        RECT 43.475 60.315 44.680 60.485 ;
        RECT 43.475 59.885 43.805 60.315 ;
        RECT 43.985 59.705 44.180 60.145 ;
        RECT 44.350 59.885 44.680 60.315 ;
        RECT 44.850 59.885 45.125 60.655 ;
        RECT 45.305 59.705 47.895 60.795 ;
        RECT 48.075 59.705 48.405 60.845 ;
        RECT 48.585 60.675 49.265 60.845 ;
        RECT 50.365 60.795 51.115 61.315 ;
        RECT 48.935 59.890 49.265 60.675 ;
        RECT 49.445 59.705 51.115 60.795 ;
        RECT 51.320 60.495 51.635 61.515 ;
        RECT 51.805 60.845 51.975 61.345 ;
        RECT 52.225 61.015 52.490 61.575 ;
        RECT 52.660 60.845 52.830 61.745 ;
        RECT 53.000 61.015 53.355 61.575 ;
        RECT 53.675 61.385 53.845 61.950 ;
        RECT 54.035 61.725 54.265 62.030 ;
        RECT 54.435 61.895 54.765 62.255 ;
        RECT 54.960 61.725 55.250 62.075 ;
        RECT 54.035 61.555 55.250 61.725 ;
        RECT 55.425 61.710 60.770 62.255 ;
        RECT 53.675 61.215 54.195 61.385 ;
        RECT 51.805 60.675 53.230 60.845 ;
        RECT 53.590 60.685 53.835 61.045 ;
        RECT 54.025 60.835 54.195 61.215 ;
        RECT 54.365 61.015 54.750 61.345 ;
        RECT 54.930 61.235 55.190 61.345 ;
        RECT 54.930 61.065 55.195 61.235 ;
        RECT 54.930 61.015 55.190 61.065 ;
        RECT 51.320 59.875 51.855 60.495 ;
        RECT 52.025 59.705 52.355 60.505 ;
        RECT 52.840 60.500 53.230 60.675 ;
        RECT 54.025 60.555 54.375 60.835 ;
        RECT 53.590 59.705 53.845 60.505 ;
        RECT 54.045 59.875 54.375 60.555 ;
        RECT 54.555 59.965 54.750 61.015 ;
        RECT 57.010 60.880 57.350 61.710 ;
        RECT 60.945 61.485 63.535 62.255 ;
        RECT 63.705 61.530 63.995 62.255 ;
        RECT 65.130 61.795 65.395 62.255 ;
        RECT 65.765 61.615 65.935 62.085 ;
        RECT 66.185 61.795 66.355 62.255 ;
        RECT 66.605 61.615 66.775 62.085 ;
        RECT 67.025 61.795 67.195 62.255 ;
        RECT 67.445 61.615 67.615 62.085 ;
        RECT 67.785 61.790 68.035 62.255 ;
        RECT 54.930 59.705 55.250 60.845 ;
        RECT 58.830 60.140 59.180 61.390 ;
        RECT 60.945 60.965 62.155 61.485 ;
        RECT 65.765 61.435 68.135 61.615 ;
        RECT 62.325 60.795 63.535 61.315 ;
        RECT 65.105 61.015 67.615 61.265 ;
        RECT 55.425 59.705 60.770 60.140 ;
        RECT 60.945 59.705 63.535 60.795 ;
        RECT 63.705 59.705 63.995 60.870 ;
        RECT 67.785 60.845 68.135 61.435 ;
        RECT 68.305 61.485 71.815 62.255 ;
        RECT 68.305 60.965 69.955 61.485 ;
        RECT 72.450 61.415 72.710 62.255 ;
        RECT 72.885 61.510 73.140 62.085 ;
        RECT 73.310 61.875 73.640 62.255 ;
        RECT 73.855 61.705 74.025 62.085 ;
        RECT 73.310 61.535 74.025 61.705 ;
        RECT 65.130 59.705 65.425 60.845 ;
        RECT 65.685 60.675 68.135 60.845 ;
        RECT 70.125 60.795 71.815 61.315 ;
        RECT 65.685 59.875 66.015 60.675 ;
        RECT 66.185 59.705 66.355 60.505 ;
        RECT 66.525 59.875 66.855 60.675 ;
        RECT 67.365 60.655 68.135 60.675 ;
        RECT 67.025 59.705 67.195 60.505 ;
        RECT 67.365 59.875 67.695 60.655 ;
        RECT 67.865 59.705 68.035 60.165 ;
        RECT 68.305 59.705 71.815 60.795 ;
        RECT 72.450 59.705 72.710 60.855 ;
        RECT 72.885 60.780 73.055 61.510 ;
        RECT 73.310 61.345 73.480 61.535 ;
        RECT 74.290 61.415 74.550 62.255 ;
        RECT 74.725 61.510 74.980 62.085 ;
        RECT 75.150 61.875 75.480 62.255 ;
        RECT 75.695 61.705 75.865 62.085 ;
        RECT 75.150 61.535 75.865 61.705 ;
        RECT 76.125 61.580 76.385 62.085 ;
        RECT 76.565 61.875 76.895 62.255 ;
        RECT 77.075 61.705 77.245 62.085 ;
        RECT 73.225 61.015 73.480 61.345 ;
        RECT 73.310 60.805 73.480 61.015 ;
        RECT 73.760 60.985 74.115 61.355 ;
        RECT 72.885 59.875 73.140 60.780 ;
        RECT 73.310 60.635 74.025 60.805 ;
        RECT 73.310 59.705 73.640 60.465 ;
        RECT 73.855 59.875 74.025 60.635 ;
        RECT 74.290 59.705 74.550 60.855 ;
        RECT 74.725 60.780 74.895 61.510 ;
        RECT 75.150 61.345 75.320 61.535 ;
        RECT 75.065 61.015 75.320 61.345 ;
        RECT 75.150 60.805 75.320 61.015 ;
        RECT 75.600 60.985 75.955 61.355 ;
        RECT 74.725 59.875 74.980 60.780 ;
        RECT 75.150 60.635 75.865 60.805 ;
        RECT 75.150 59.705 75.480 60.465 ;
        RECT 75.695 59.875 75.865 60.635 ;
        RECT 76.125 60.780 76.305 61.580 ;
        RECT 76.580 61.535 77.245 61.705 ;
        RECT 76.580 61.280 76.750 61.535 ;
        RECT 77.710 61.475 78.210 62.085 ;
        RECT 76.475 60.950 76.750 61.280 ;
        RECT 76.975 60.985 77.315 61.355 ;
        RECT 77.505 61.015 77.855 61.265 ;
        RECT 76.580 60.805 76.750 60.950 ;
        RECT 78.040 60.845 78.210 61.475 ;
        RECT 78.840 61.605 79.170 62.085 ;
        RECT 79.340 61.795 79.565 62.255 ;
        RECT 79.735 61.605 80.065 62.085 ;
        RECT 78.840 61.435 80.065 61.605 ;
        RECT 80.255 61.455 80.505 62.255 ;
        RECT 80.675 61.455 81.015 62.085 ;
        RECT 81.275 61.705 81.445 61.995 ;
        RECT 81.615 61.875 81.945 62.255 ;
        RECT 81.275 61.535 81.940 61.705 ;
        RECT 80.785 61.405 81.015 61.455 ;
        RECT 78.380 61.065 78.710 61.265 ;
        RECT 78.880 61.065 79.210 61.265 ;
        RECT 79.380 61.065 79.800 61.265 ;
        RECT 79.975 61.095 80.670 61.265 ;
        RECT 79.975 60.845 80.145 61.095 ;
        RECT 80.840 60.845 81.015 61.405 ;
        RECT 76.125 59.875 76.395 60.780 ;
        RECT 76.580 60.635 77.255 60.805 ;
        RECT 76.565 59.705 76.895 60.465 ;
        RECT 77.075 59.875 77.255 60.635 ;
        RECT 77.710 60.675 80.145 60.845 ;
        RECT 77.710 59.875 78.040 60.675 ;
        RECT 78.210 59.705 78.540 60.505 ;
        RECT 78.840 59.875 79.170 60.675 ;
        RECT 79.815 59.705 80.065 60.505 ;
        RECT 80.335 59.705 80.505 60.845 ;
        RECT 80.675 59.875 81.015 60.845 ;
        RECT 81.190 60.715 81.540 61.365 ;
        RECT 81.710 60.545 81.940 61.535 ;
        RECT 81.275 60.375 81.940 60.545 ;
        RECT 81.275 59.875 81.445 60.375 ;
        RECT 81.615 59.705 81.945 60.205 ;
        RECT 82.115 59.875 82.300 61.995 ;
        RECT 82.555 61.795 82.805 62.255 ;
        RECT 82.975 61.805 83.310 61.975 ;
        RECT 83.505 61.805 84.180 61.975 ;
        RECT 82.975 61.665 83.145 61.805 ;
        RECT 82.470 60.675 82.750 61.625 ;
        RECT 82.920 61.535 83.145 61.665 ;
        RECT 82.920 60.430 83.090 61.535 ;
        RECT 83.315 61.385 83.840 61.605 ;
        RECT 83.260 60.620 83.500 61.215 ;
        RECT 83.670 60.685 83.840 61.385 ;
        RECT 84.010 61.025 84.180 61.805 ;
        RECT 84.500 61.755 84.870 62.255 ;
        RECT 85.050 61.805 85.455 61.975 ;
        RECT 85.625 61.805 86.410 61.975 ;
        RECT 85.050 61.575 85.220 61.805 ;
        RECT 84.390 61.275 85.220 61.575 ;
        RECT 85.605 61.305 86.070 61.635 ;
        RECT 84.390 61.245 84.590 61.275 ;
        RECT 84.710 61.025 84.880 61.095 ;
        RECT 84.010 60.855 84.880 61.025 ;
        RECT 84.370 60.765 84.880 60.855 ;
        RECT 82.920 60.300 83.225 60.430 ;
        RECT 83.670 60.320 84.200 60.685 ;
        RECT 82.540 59.705 82.805 60.165 ;
        RECT 82.975 59.875 83.225 60.300 ;
        RECT 84.370 60.150 84.540 60.765 ;
        RECT 83.435 59.980 84.540 60.150 ;
        RECT 84.710 59.705 84.880 60.505 ;
        RECT 85.050 60.205 85.220 61.275 ;
        RECT 85.390 60.375 85.580 61.095 ;
        RECT 85.750 60.345 86.070 61.305 ;
        RECT 86.240 61.345 86.410 61.805 ;
        RECT 86.685 61.725 86.895 62.255 ;
        RECT 87.155 61.515 87.485 62.040 ;
        RECT 87.655 61.645 87.825 62.255 ;
        RECT 87.995 61.600 88.325 62.035 ;
        RECT 87.995 61.515 88.375 61.600 ;
        RECT 87.285 61.345 87.485 61.515 ;
        RECT 88.150 61.475 88.375 61.515 ;
        RECT 88.545 61.505 89.755 62.255 ;
        RECT 86.240 61.015 87.115 61.345 ;
        RECT 87.285 61.015 88.035 61.345 ;
        RECT 85.050 59.875 85.300 60.205 ;
        RECT 86.240 60.175 86.410 61.015 ;
        RECT 87.285 60.810 87.475 61.015 ;
        RECT 88.205 60.895 88.375 61.475 ;
        RECT 88.160 60.845 88.375 60.895 ;
        RECT 86.580 60.435 87.475 60.810 ;
        RECT 87.985 60.765 88.375 60.845 ;
        RECT 88.545 60.795 89.065 61.335 ;
        RECT 89.235 60.965 89.755 61.505 ;
        RECT 85.525 60.005 86.410 60.175 ;
        RECT 86.590 59.705 86.905 60.205 ;
        RECT 87.135 59.875 87.475 60.435 ;
        RECT 87.645 59.705 87.815 60.715 ;
        RECT 87.985 59.920 88.315 60.765 ;
        RECT 88.545 59.705 89.755 60.795 ;
        RECT 12.100 59.535 89.840 59.705 ;
        RECT 12.185 58.445 13.395 59.535 ;
        RECT 13.565 59.100 18.910 59.535 ;
        RECT 12.185 57.735 12.705 58.275 ;
        RECT 12.875 57.905 13.395 58.445 ;
        RECT 12.185 56.985 13.395 57.735 ;
        RECT 15.150 57.530 15.490 58.360 ;
        RECT 16.970 57.850 17.320 59.100 ;
        RECT 19.085 58.445 21.675 59.535 ;
        RECT 19.085 57.755 20.295 58.275 ;
        RECT 20.465 57.925 21.675 58.445 ;
        RECT 13.565 56.985 18.910 57.530 ;
        RECT 19.085 56.985 21.675 57.755 ;
        RECT 22.315 57.165 22.575 59.355 ;
        RECT 22.745 58.805 23.085 59.535 ;
        RECT 23.265 58.625 23.535 59.355 ;
        RECT 22.765 58.405 23.535 58.625 ;
        RECT 23.715 58.645 23.945 59.355 ;
        RECT 24.115 58.825 24.445 59.535 ;
        RECT 24.615 58.645 24.875 59.355 ;
        RECT 23.715 58.405 24.875 58.645 ;
        RECT 22.765 57.735 23.055 58.405 ;
        RECT 25.065 58.370 25.355 59.535 ;
        RECT 25.985 58.565 26.255 59.335 ;
        RECT 26.425 58.755 26.755 59.535 ;
        RECT 26.960 58.930 27.145 59.335 ;
        RECT 27.315 59.110 27.650 59.535 ;
        RECT 26.960 58.755 27.625 58.930 ;
        RECT 28.075 58.805 28.370 59.535 ;
        RECT 25.985 58.395 27.115 58.565 ;
        RECT 23.235 57.915 23.700 58.225 ;
        RECT 23.880 57.915 24.405 58.225 ;
        RECT 22.765 57.535 23.995 57.735 ;
        RECT 22.835 56.985 23.505 57.355 ;
        RECT 23.685 57.165 23.995 57.535 ;
        RECT 24.175 57.275 24.405 57.915 ;
        RECT 24.585 57.895 24.885 58.225 ;
        RECT 24.585 56.985 24.875 57.715 ;
        RECT 25.065 56.985 25.355 57.710 ;
        RECT 25.985 57.485 26.155 58.395 ;
        RECT 26.325 57.645 26.685 58.225 ;
        RECT 26.865 57.895 27.115 58.395 ;
        RECT 27.285 57.725 27.625 58.755 ;
        RECT 28.540 58.635 28.800 59.360 ;
        RECT 28.970 58.805 29.230 59.535 ;
        RECT 29.400 58.635 29.660 59.360 ;
        RECT 29.830 58.805 30.090 59.535 ;
        RECT 30.260 58.635 30.520 59.360 ;
        RECT 30.690 58.805 30.950 59.535 ;
        RECT 31.120 58.635 31.380 59.360 ;
        RECT 26.940 57.555 27.625 57.725 ;
        RECT 28.070 58.395 31.380 58.635 ;
        RECT 31.550 58.425 31.810 59.535 ;
        RECT 28.070 57.805 29.040 58.395 ;
        RECT 31.980 58.225 32.230 59.360 ;
        RECT 32.410 58.425 32.705 59.535 ;
        RECT 32.945 58.475 33.275 59.320 ;
        RECT 33.445 58.525 33.615 59.535 ;
        RECT 33.785 58.805 34.125 59.365 ;
        RECT 34.355 59.035 34.670 59.535 ;
        RECT 34.850 59.065 35.735 59.235 ;
        RECT 32.885 58.395 33.275 58.475 ;
        RECT 33.785 58.430 34.680 58.805 ;
        RECT 32.885 58.345 33.100 58.395 ;
        RECT 29.210 57.975 32.230 58.225 ;
        RECT 28.070 57.635 31.380 57.805 ;
        RECT 25.985 57.155 26.245 57.485 ;
        RECT 26.455 56.985 26.730 57.465 ;
        RECT 26.940 57.155 27.145 57.555 ;
        RECT 27.315 56.985 27.650 57.385 ;
        RECT 28.070 56.985 28.370 57.465 ;
        RECT 28.540 57.180 28.800 57.635 ;
        RECT 28.970 56.985 29.230 57.465 ;
        RECT 29.400 57.180 29.660 57.635 ;
        RECT 29.830 56.985 30.090 57.465 ;
        RECT 30.260 57.180 30.520 57.635 ;
        RECT 30.690 56.985 30.950 57.465 ;
        RECT 31.120 57.180 31.380 57.635 ;
        RECT 31.550 56.985 31.810 57.510 ;
        RECT 31.980 57.165 32.230 57.975 ;
        RECT 32.400 57.615 32.715 58.225 ;
        RECT 32.885 57.765 33.055 58.345 ;
        RECT 33.785 58.225 33.975 58.430 ;
        RECT 34.850 58.225 35.020 59.065 ;
        RECT 35.960 59.035 36.210 59.365 ;
        RECT 33.225 57.895 33.975 58.225 ;
        RECT 34.145 57.895 35.020 58.225 ;
        RECT 32.885 57.725 33.110 57.765 ;
        RECT 33.775 57.725 33.975 57.895 ;
        RECT 32.885 57.640 33.265 57.725 ;
        RECT 32.410 56.985 32.655 57.445 ;
        RECT 32.935 57.205 33.265 57.640 ;
        RECT 33.435 56.985 33.605 57.595 ;
        RECT 33.775 57.200 34.105 57.725 ;
        RECT 34.365 56.985 34.575 57.515 ;
        RECT 34.850 57.435 35.020 57.895 ;
        RECT 35.190 57.935 35.510 58.895 ;
        RECT 35.680 58.145 35.870 58.865 ;
        RECT 36.040 57.965 36.210 59.035 ;
        RECT 36.380 58.735 36.550 59.535 ;
        RECT 36.720 59.090 37.825 59.260 ;
        RECT 36.720 58.475 36.890 59.090 ;
        RECT 38.035 58.940 38.285 59.365 ;
        RECT 38.455 59.075 38.720 59.535 ;
        RECT 37.060 58.555 37.590 58.920 ;
        RECT 38.035 58.810 38.340 58.940 ;
        RECT 36.380 58.385 36.890 58.475 ;
        RECT 36.380 58.215 37.250 58.385 ;
        RECT 36.380 58.145 36.550 58.215 ;
        RECT 36.670 57.965 36.870 57.995 ;
        RECT 35.190 57.605 35.655 57.935 ;
        RECT 36.040 57.665 36.870 57.965 ;
        RECT 36.040 57.435 36.210 57.665 ;
        RECT 34.850 57.265 35.635 57.435 ;
        RECT 35.805 57.265 36.210 57.435 ;
        RECT 36.390 56.985 36.760 57.485 ;
        RECT 37.080 57.435 37.250 58.215 ;
        RECT 37.420 57.855 37.590 58.555 ;
        RECT 37.760 58.025 38.000 58.620 ;
        RECT 37.420 57.635 37.945 57.855 ;
        RECT 38.170 57.705 38.340 58.810 ;
        RECT 38.115 57.575 38.340 57.705 ;
        RECT 38.510 57.615 38.790 58.565 ;
        RECT 38.115 57.435 38.285 57.575 ;
        RECT 37.080 57.265 37.755 57.435 ;
        RECT 37.950 57.265 38.285 57.435 ;
        RECT 38.455 56.985 38.705 57.445 ;
        RECT 38.960 57.245 39.145 59.365 ;
        RECT 39.315 59.035 39.645 59.535 ;
        RECT 39.815 58.865 39.985 59.365 ;
        RECT 40.245 59.025 40.505 59.535 ;
        RECT 39.320 58.695 39.985 58.865 ;
        RECT 39.320 57.705 39.550 58.695 ;
        RECT 39.720 57.875 40.070 58.525 ;
        RECT 40.245 57.975 40.585 58.855 ;
        RECT 40.755 58.145 40.925 59.365 ;
        RECT 41.165 59.030 41.780 59.535 ;
        RECT 41.165 58.495 41.415 58.860 ;
        RECT 41.585 58.855 41.780 59.030 ;
        RECT 41.950 59.025 42.425 59.365 ;
        RECT 42.595 58.990 42.810 59.535 ;
        RECT 41.585 58.665 41.915 58.855 ;
        RECT 42.135 58.495 42.850 58.790 ;
        RECT 43.020 58.665 43.295 59.365 ;
        RECT 43.580 58.905 43.865 59.365 ;
        RECT 44.035 59.075 44.305 59.535 ;
        RECT 43.580 58.685 44.535 58.905 ;
        RECT 41.165 58.325 42.955 58.495 ;
        RECT 40.755 57.895 41.550 58.145 ;
        RECT 40.755 57.805 41.005 57.895 ;
        RECT 39.320 57.535 39.985 57.705 ;
        RECT 39.315 56.985 39.645 57.365 ;
        RECT 39.815 57.245 39.985 57.535 ;
        RECT 40.245 56.985 40.505 57.805 ;
        RECT 40.675 57.385 41.005 57.805 ;
        RECT 41.720 57.470 41.975 58.325 ;
        RECT 41.185 57.205 41.975 57.470 ;
        RECT 42.145 57.625 42.555 58.145 ;
        RECT 42.725 57.895 42.955 58.325 ;
        RECT 43.125 57.635 43.295 58.665 ;
        RECT 43.465 57.955 44.155 58.515 ;
        RECT 44.325 57.785 44.535 58.685 ;
        RECT 42.145 57.205 42.345 57.625 ;
        RECT 42.535 56.985 42.865 57.445 ;
        RECT 43.035 57.155 43.295 57.635 ;
        RECT 43.580 57.615 44.535 57.785 ;
        RECT 44.705 58.515 45.105 59.365 ;
        RECT 45.295 58.905 45.575 59.365 ;
        RECT 46.095 59.075 46.420 59.535 ;
        RECT 45.295 58.685 46.420 58.905 ;
        RECT 44.705 57.955 45.800 58.515 ;
        RECT 45.970 58.225 46.420 58.685 ;
        RECT 46.590 58.395 46.975 59.365 ;
        RECT 47.155 58.585 47.430 59.355 ;
        RECT 47.600 58.925 47.930 59.355 ;
        RECT 48.100 59.095 48.295 59.535 ;
        RECT 48.475 58.925 48.805 59.355 ;
        RECT 47.600 58.755 48.805 58.925 ;
        RECT 47.155 58.395 47.740 58.585 ;
        RECT 47.910 58.425 48.805 58.755 ;
        RECT 49.455 58.395 49.785 59.535 ;
        RECT 50.315 58.565 50.645 59.350 ;
        RECT 49.965 58.395 50.645 58.565 ;
        RECT 43.580 57.155 43.865 57.615 ;
        RECT 44.035 56.985 44.305 57.445 ;
        RECT 44.705 57.155 45.105 57.955 ;
        RECT 45.970 57.895 46.525 58.225 ;
        RECT 45.970 57.785 46.420 57.895 ;
        RECT 45.295 57.615 46.420 57.785 ;
        RECT 46.695 57.725 46.975 58.395 ;
        RECT 45.295 57.155 45.575 57.615 ;
        RECT 46.095 56.985 46.420 57.445 ;
        RECT 46.590 57.155 46.975 57.725 ;
        RECT 47.155 57.575 47.395 58.225 ;
        RECT 47.565 57.725 47.740 58.395 ;
        RECT 47.910 57.895 48.325 58.225 ;
        RECT 48.505 57.895 48.800 58.225 ;
        RECT 49.445 57.975 49.795 58.225 ;
        RECT 47.565 57.545 47.895 57.725 ;
        RECT 47.170 56.985 47.500 57.375 ;
        RECT 47.670 57.165 47.895 57.545 ;
        RECT 48.095 57.275 48.325 57.895 ;
        RECT 49.965 57.795 50.135 58.395 ;
        RECT 50.825 58.370 51.115 59.535 ;
        RECT 51.285 58.395 51.670 59.365 ;
        RECT 51.840 59.075 52.165 59.535 ;
        RECT 52.685 58.905 52.965 59.365 ;
        RECT 51.840 58.685 52.965 58.905 ;
        RECT 50.305 57.975 50.655 58.225 ;
        RECT 48.505 56.985 48.805 57.715 ;
        RECT 49.455 56.985 49.725 57.795 ;
        RECT 49.895 57.155 50.225 57.795 ;
        RECT 50.395 56.985 50.635 57.795 ;
        RECT 51.285 57.725 51.565 58.395 ;
        RECT 51.840 58.225 52.290 58.685 ;
        RECT 53.155 58.515 53.555 59.365 ;
        RECT 53.955 59.075 54.225 59.535 ;
        RECT 54.395 58.905 54.680 59.365 ;
        RECT 51.735 57.895 52.290 58.225 ;
        RECT 52.460 57.955 53.555 58.515 ;
        RECT 51.840 57.785 52.290 57.895 ;
        RECT 50.825 56.985 51.115 57.710 ;
        RECT 51.285 57.155 51.670 57.725 ;
        RECT 51.840 57.615 52.965 57.785 ;
        RECT 51.840 56.985 52.165 57.445 ;
        RECT 52.685 57.155 52.965 57.615 ;
        RECT 53.155 57.155 53.555 57.955 ;
        RECT 53.725 58.685 54.680 58.905 ;
        RECT 53.725 57.785 53.935 58.685 ;
        RECT 54.105 57.955 54.795 58.515 ;
        RECT 55.885 58.395 56.270 59.365 ;
        RECT 56.440 59.075 56.765 59.535 ;
        RECT 57.285 58.905 57.565 59.365 ;
        RECT 56.440 58.685 57.565 58.905 ;
        RECT 53.725 57.615 54.680 57.785 ;
        RECT 53.955 56.985 54.225 57.445 ;
        RECT 54.395 57.155 54.680 57.615 ;
        RECT 55.885 57.725 56.165 58.395 ;
        RECT 56.440 58.225 56.890 58.685 ;
        RECT 57.755 58.515 58.155 59.365 ;
        RECT 58.555 59.075 58.825 59.535 ;
        RECT 58.995 58.905 59.280 59.365 ;
        RECT 56.335 57.895 56.890 58.225 ;
        RECT 57.060 57.955 58.155 58.515 ;
        RECT 56.440 57.785 56.890 57.895 ;
        RECT 55.885 57.155 56.270 57.725 ;
        RECT 56.440 57.615 57.565 57.785 ;
        RECT 56.440 56.985 56.765 57.445 ;
        RECT 57.285 57.155 57.565 57.615 ;
        RECT 57.755 57.155 58.155 57.955 ;
        RECT 58.325 58.685 59.280 58.905 ;
        RECT 58.325 57.785 58.535 58.685 ;
        RECT 58.705 57.955 59.395 58.515 ;
        RECT 59.565 58.445 62.155 59.535 ;
        RECT 62.415 58.865 62.585 59.365 ;
        RECT 62.755 59.035 63.085 59.535 ;
        RECT 62.415 58.695 63.080 58.865 ;
        RECT 58.325 57.615 59.280 57.785 ;
        RECT 58.555 56.985 58.825 57.445 ;
        RECT 58.995 57.155 59.280 57.615 ;
        RECT 59.565 57.755 60.775 58.275 ;
        RECT 60.945 57.925 62.155 58.445 ;
        RECT 62.330 57.875 62.680 58.525 ;
        RECT 59.565 56.985 62.155 57.755 ;
        RECT 62.850 57.705 63.080 58.695 ;
        RECT 62.415 57.535 63.080 57.705 ;
        RECT 62.415 57.245 62.585 57.535 ;
        RECT 62.755 56.985 63.085 57.365 ;
        RECT 63.255 57.245 63.440 59.365 ;
        RECT 63.680 59.075 63.945 59.535 ;
        RECT 64.115 58.940 64.365 59.365 ;
        RECT 64.575 59.090 65.680 59.260 ;
        RECT 64.060 58.810 64.365 58.940 ;
        RECT 63.610 57.615 63.890 58.565 ;
        RECT 64.060 57.705 64.230 58.810 ;
        RECT 64.400 58.025 64.640 58.620 ;
        RECT 64.810 58.555 65.340 58.920 ;
        RECT 64.810 57.855 64.980 58.555 ;
        RECT 65.510 58.475 65.680 59.090 ;
        RECT 65.850 58.735 66.020 59.535 ;
        RECT 66.190 59.035 66.440 59.365 ;
        RECT 66.665 59.065 67.550 59.235 ;
        RECT 65.510 58.385 66.020 58.475 ;
        RECT 64.060 57.575 64.285 57.705 ;
        RECT 64.455 57.635 64.980 57.855 ;
        RECT 65.150 58.215 66.020 58.385 ;
        RECT 63.695 56.985 63.945 57.445 ;
        RECT 64.115 57.435 64.285 57.575 ;
        RECT 65.150 57.435 65.320 58.215 ;
        RECT 65.850 58.145 66.020 58.215 ;
        RECT 65.530 57.965 65.730 57.995 ;
        RECT 66.190 57.965 66.360 59.035 ;
        RECT 66.530 58.145 66.720 58.865 ;
        RECT 65.530 57.665 66.360 57.965 ;
        RECT 66.890 57.935 67.210 58.895 ;
        RECT 64.115 57.265 64.450 57.435 ;
        RECT 64.645 57.265 65.320 57.435 ;
        RECT 65.640 56.985 66.010 57.485 ;
        RECT 66.190 57.435 66.360 57.665 ;
        RECT 66.745 57.605 67.210 57.935 ;
        RECT 67.380 58.225 67.550 59.065 ;
        RECT 67.730 59.035 68.045 59.535 ;
        RECT 68.275 58.805 68.615 59.365 ;
        RECT 67.720 58.430 68.615 58.805 ;
        RECT 68.785 58.525 68.955 59.535 ;
        RECT 68.425 58.225 68.615 58.430 ;
        RECT 69.125 58.475 69.455 59.320 ;
        RECT 69.125 58.395 69.515 58.475 ;
        RECT 69.685 58.445 70.895 59.535 ;
        RECT 69.300 58.345 69.515 58.395 ;
        RECT 67.380 57.895 68.255 58.225 ;
        RECT 68.425 57.895 69.175 58.225 ;
        RECT 67.380 57.435 67.550 57.895 ;
        RECT 68.425 57.725 68.625 57.895 ;
        RECT 69.345 57.765 69.515 58.345 ;
        RECT 69.290 57.725 69.515 57.765 ;
        RECT 66.190 57.265 66.595 57.435 ;
        RECT 66.765 57.265 67.550 57.435 ;
        RECT 67.825 56.985 68.035 57.515 ;
        RECT 68.295 57.200 68.625 57.725 ;
        RECT 69.135 57.640 69.515 57.725 ;
        RECT 69.685 57.735 70.205 58.275 ;
        RECT 70.375 57.905 70.895 58.445 ;
        RECT 71.070 58.385 71.330 59.535 ;
        RECT 71.505 58.460 71.760 59.365 ;
        RECT 71.930 58.775 72.260 59.535 ;
        RECT 72.475 58.605 72.645 59.365 ;
        RECT 68.795 56.985 68.965 57.595 ;
        RECT 69.135 57.205 69.465 57.640 ;
        RECT 69.685 56.985 70.895 57.735 ;
        RECT 71.070 56.985 71.330 57.825 ;
        RECT 71.505 57.730 71.675 58.460 ;
        RECT 71.930 58.435 72.645 58.605 ;
        RECT 71.930 58.225 72.100 58.435 ;
        RECT 72.905 58.395 73.245 59.365 ;
        RECT 73.415 58.395 73.585 59.535 ;
        RECT 73.855 58.735 74.105 59.535 ;
        RECT 74.750 58.565 75.080 59.365 ;
        RECT 75.380 58.735 75.710 59.535 ;
        RECT 75.880 58.565 76.210 59.365 ;
        RECT 73.775 58.395 76.210 58.565 ;
        RECT 71.845 57.895 72.100 58.225 ;
        RECT 71.505 57.155 71.760 57.730 ;
        RECT 71.930 57.705 72.100 57.895 ;
        RECT 72.380 57.885 72.735 58.255 ;
        RECT 72.905 57.785 73.080 58.395 ;
        RECT 73.775 58.145 73.945 58.395 ;
        RECT 73.250 57.975 73.945 58.145 ;
        RECT 74.120 57.975 74.540 58.175 ;
        RECT 74.710 57.975 75.040 58.175 ;
        RECT 75.210 57.975 75.540 58.175 ;
        RECT 71.930 57.535 72.645 57.705 ;
        RECT 71.930 56.985 72.260 57.365 ;
        RECT 72.475 57.155 72.645 57.535 ;
        RECT 72.905 57.155 73.245 57.785 ;
        RECT 73.415 56.985 73.665 57.785 ;
        RECT 73.855 57.635 75.080 57.805 ;
        RECT 73.855 57.155 74.185 57.635 ;
        RECT 74.355 56.985 74.580 57.445 ;
        RECT 74.750 57.155 75.080 57.635 ;
        RECT 75.710 57.765 75.880 58.395 ;
        RECT 76.585 58.370 76.875 59.535 ;
        RECT 77.135 58.865 77.305 59.365 ;
        RECT 77.475 59.035 77.805 59.535 ;
        RECT 77.135 58.695 77.800 58.865 ;
        RECT 76.065 57.975 76.415 58.225 ;
        RECT 77.050 57.875 77.400 58.525 ;
        RECT 75.710 57.155 76.210 57.765 ;
        RECT 76.585 56.985 76.875 57.710 ;
        RECT 77.570 57.705 77.800 58.695 ;
        RECT 77.135 57.535 77.800 57.705 ;
        RECT 77.135 57.245 77.305 57.535 ;
        RECT 77.475 56.985 77.805 57.365 ;
        RECT 77.975 57.245 78.160 59.365 ;
        RECT 78.400 59.075 78.665 59.535 ;
        RECT 78.835 58.940 79.085 59.365 ;
        RECT 79.295 59.090 80.400 59.260 ;
        RECT 78.780 58.810 79.085 58.940 ;
        RECT 78.330 57.615 78.610 58.565 ;
        RECT 78.780 57.705 78.950 58.810 ;
        RECT 79.120 58.025 79.360 58.620 ;
        RECT 79.530 58.555 80.060 58.920 ;
        RECT 79.530 57.855 79.700 58.555 ;
        RECT 80.230 58.475 80.400 59.090 ;
        RECT 80.570 58.735 80.740 59.535 ;
        RECT 80.910 59.035 81.160 59.365 ;
        RECT 81.385 59.065 82.270 59.235 ;
        RECT 80.230 58.385 80.740 58.475 ;
        RECT 78.780 57.575 79.005 57.705 ;
        RECT 79.175 57.635 79.700 57.855 ;
        RECT 79.870 58.215 80.740 58.385 ;
        RECT 78.415 56.985 78.665 57.445 ;
        RECT 78.835 57.435 79.005 57.575 ;
        RECT 79.870 57.435 80.040 58.215 ;
        RECT 80.570 58.145 80.740 58.215 ;
        RECT 80.250 57.965 80.450 57.995 ;
        RECT 80.910 57.965 81.080 59.035 ;
        RECT 81.250 58.145 81.440 58.865 ;
        RECT 80.250 57.665 81.080 57.965 ;
        RECT 81.610 57.935 81.930 58.895 ;
        RECT 78.835 57.265 79.170 57.435 ;
        RECT 79.365 57.265 80.040 57.435 ;
        RECT 80.360 56.985 80.730 57.485 ;
        RECT 80.910 57.435 81.080 57.665 ;
        RECT 81.465 57.605 81.930 57.935 ;
        RECT 82.100 58.225 82.270 59.065 ;
        RECT 82.450 59.035 82.765 59.535 ;
        RECT 82.995 58.805 83.335 59.365 ;
        RECT 82.440 58.430 83.335 58.805 ;
        RECT 83.505 58.525 83.675 59.535 ;
        RECT 83.145 58.225 83.335 58.430 ;
        RECT 83.845 58.475 84.175 59.320 ;
        RECT 84.440 58.745 84.975 59.365 ;
        RECT 83.845 58.395 84.235 58.475 ;
        RECT 84.020 58.345 84.235 58.395 ;
        RECT 82.100 57.895 82.975 58.225 ;
        RECT 83.145 57.895 83.895 58.225 ;
        RECT 82.100 57.435 82.270 57.895 ;
        RECT 83.145 57.725 83.345 57.895 ;
        RECT 84.065 57.765 84.235 58.345 ;
        RECT 84.010 57.725 84.235 57.765 ;
        RECT 80.910 57.265 81.315 57.435 ;
        RECT 81.485 57.265 82.270 57.435 ;
        RECT 82.545 56.985 82.755 57.515 ;
        RECT 83.015 57.200 83.345 57.725 ;
        RECT 83.855 57.640 84.235 57.725 ;
        RECT 84.440 57.725 84.755 58.745 ;
        RECT 85.145 58.735 85.475 59.535 ;
        RECT 85.960 58.565 86.350 58.740 ;
        RECT 84.925 58.395 86.350 58.565 ;
        RECT 86.795 58.605 86.965 59.365 ;
        RECT 87.180 58.775 87.510 59.535 ;
        RECT 86.795 58.435 87.510 58.605 ;
        RECT 87.680 58.460 87.935 59.365 ;
        RECT 84.925 57.895 85.095 58.395 ;
        RECT 83.515 56.985 83.685 57.595 ;
        RECT 83.855 57.205 84.185 57.640 ;
        RECT 84.440 57.155 85.055 57.725 ;
        RECT 85.345 57.665 85.610 58.225 ;
        RECT 85.780 57.495 85.950 58.395 ;
        RECT 86.120 57.665 86.475 58.225 ;
        RECT 86.705 57.885 87.060 58.255 ;
        RECT 87.340 58.225 87.510 58.435 ;
        RECT 87.340 57.895 87.595 58.225 ;
        RECT 87.340 57.705 87.510 57.895 ;
        RECT 87.765 57.730 87.935 58.460 ;
        RECT 88.110 58.385 88.370 59.535 ;
        RECT 88.545 58.445 89.755 59.535 ;
        RECT 88.545 57.905 89.065 58.445 ;
        RECT 86.795 57.535 87.510 57.705 ;
        RECT 85.225 56.985 85.440 57.495 ;
        RECT 85.670 57.165 85.950 57.495 ;
        RECT 86.130 56.985 86.370 57.495 ;
        RECT 86.795 57.155 86.965 57.535 ;
        RECT 87.180 56.985 87.510 57.365 ;
        RECT 87.680 57.155 87.935 57.730 ;
        RECT 88.110 56.985 88.370 57.825 ;
        RECT 89.235 57.735 89.755 58.275 ;
        RECT 88.545 56.985 89.755 57.735 ;
        RECT 12.100 56.815 89.840 56.985 ;
        RECT 12.185 56.065 13.395 56.815 ;
        RECT 13.565 56.270 18.910 56.815 ;
        RECT 12.185 55.525 12.705 56.065 ;
        RECT 12.875 55.355 13.395 55.895 ;
        RECT 15.150 55.440 15.490 56.270 ;
        RECT 19.085 56.065 20.295 56.815 ;
        RECT 20.470 56.285 20.760 56.635 ;
        RECT 20.955 56.455 21.285 56.815 ;
        RECT 21.455 56.285 21.685 56.590 ;
        RECT 20.470 56.115 21.685 56.285 ;
        RECT 21.875 56.475 22.045 56.510 ;
        RECT 21.875 56.305 22.075 56.475 ;
        RECT 12.185 54.265 13.395 55.355 ;
        RECT 16.970 54.700 17.320 55.950 ;
        RECT 19.085 55.525 19.605 56.065 ;
        RECT 21.875 55.945 22.045 56.305 ;
        RECT 19.775 55.355 20.295 55.895 ;
        RECT 20.530 55.795 20.790 55.905 ;
        RECT 20.525 55.625 20.790 55.795 ;
        RECT 20.530 55.575 20.790 55.625 ;
        RECT 20.970 55.575 21.355 55.905 ;
        RECT 21.525 55.775 22.045 55.945 ;
        RECT 22.305 56.075 22.770 56.620 ;
        RECT 13.565 54.265 18.910 54.700 ;
        RECT 19.085 54.265 20.295 55.355 ;
        RECT 20.470 54.265 20.790 55.405 ;
        RECT 20.970 54.525 21.165 55.575 ;
        RECT 21.525 55.395 21.695 55.775 ;
        RECT 21.345 55.115 21.695 55.395 ;
        RECT 21.885 55.245 22.130 55.605 ;
        RECT 22.305 55.115 22.475 56.075 ;
        RECT 23.275 55.995 23.445 56.815 ;
        RECT 23.615 56.165 23.945 56.645 ;
        RECT 24.115 56.425 24.465 56.815 ;
        RECT 24.635 56.245 24.865 56.645 ;
        RECT 24.355 56.165 24.865 56.245 ;
        RECT 23.615 56.075 24.865 56.165 ;
        RECT 25.035 56.075 25.355 56.555 ;
        RECT 25.610 56.245 25.785 56.645 ;
        RECT 25.955 56.435 26.285 56.815 ;
        RECT 26.530 56.315 26.760 56.645 ;
        RECT 25.610 56.075 26.240 56.245 ;
        RECT 23.615 55.995 24.525 56.075 ;
        RECT 22.645 55.455 22.890 55.905 ;
        RECT 23.150 55.625 23.845 55.825 ;
        RECT 24.015 55.655 24.615 55.825 ;
        RECT 24.015 55.455 24.185 55.655 ;
        RECT 24.845 55.485 25.015 55.905 ;
        RECT 22.645 55.285 24.185 55.455 ;
        RECT 24.355 55.315 25.015 55.485 ;
        RECT 24.355 55.115 24.525 55.315 ;
        RECT 25.185 55.145 25.355 56.075 ;
        RECT 26.070 55.905 26.240 56.075 ;
        RECT 25.525 55.225 25.890 55.905 ;
        RECT 26.070 55.575 26.420 55.905 ;
        RECT 21.345 54.435 21.675 55.115 ;
        RECT 21.875 54.265 22.130 55.065 ;
        RECT 22.305 54.945 24.525 55.115 ;
        RECT 24.695 54.945 25.355 55.145 ;
        RECT 26.070 55.055 26.240 55.575 ;
        RECT 22.305 54.265 22.605 54.775 ;
        RECT 22.775 54.435 23.105 54.945 ;
        RECT 24.695 54.775 24.865 54.945 ;
        RECT 25.610 54.885 26.240 55.055 ;
        RECT 26.590 55.025 26.760 56.315 ;
        RECT 26.960 55.205 27.240 56.480 ;
        RECT 27.465 56.475 27.735 56.480 ;
        RECT 27.425 56.305 27.735 56.475 ;
        RECT 28.195 56.435 28.525 56.815 ;
        RECT 28.695 56.560 29.030 56.605 ;
        RECT 27.465 55.205 27.735 56.305 ;
        RECT 27.925 55.205 28.265 56.235 ;
        RECT 28.695 56.095 29.035 56.560 ;
        RECT 30.175 56.355 30.480 56.815 ;
        RECT 30.650 56.185 30.980 56.645 ;
        RECT 31.150 56.355 31.320 56.815 ;
        RECT 31.490 56.185 31.820 56.645 ;
        RECT 31.990 56.355 32.160 56.815 ;
        RECT 32.330 56.185 32.660 56.645 ;
        RECT 32.830 56.355 33.000 56.815 ;
        RECT 33.170 56.185 33.500 56.645 ;
        RECT 33.670 56.355 33.925 56.815 ;
        RECT 28.435 55.575 28.695 55.905 ;
        RECT 28.435 55.025 28.605 55.575 ;
        RECT 28.865 55.405 29.035 56.095 ;
        RECT 23.275 54.265 23.905 54.775 ;
        RECT 24.485 54.605 24.865 54.775 ;
        RECT 25.035 54.265 25.335 54.775 ;
        RECT 25.610 54.435 25.785 54.885 ;
        RECT 26.590 54.855 28.605 55.025 ;
        RECT 25.955 54.265 26.285 54.705 ;
        RECT 26.590 54.435 26.760 54.855 ;
        RECT 26.995 54.265 27.665 54.675 ;
        RECT 27.880 54.435 28.050 54.855 ;
        RECT 28.250 54.265 28.580 54.675 ;
        RECT 28.775 54.435 29.035 55.405 ;
        RECT 30.125 55.995 34.095 56.185 ;
        RECT 30.125 55.405 30.445 55.995 ;
        RECT 30.645 55.575 33.500 55.825 ;
        RECT 33.750 55.405 34.095 55.995 ;
        RECT 30.125 55.235 34.095 55.405 ;
        RECT 34.285 56.125 34.525 56.645 ;
        RECT 34.695 56.320 35.090 56.815 ;
        RECT 35.655 56.485 35.825 56.630 ;
        RECT 35.450 56.290 35.825 56.485 ;
        RECT 34.285 55.455 34.460 56.125 ;
        RECT 35.450 55.955 35.620 56.290 ;
        RECT 36.105 56.245 36.345 56.620 ;
        RECT 36.515 56.310 36.850 56.815 ;
        RECT 36.105 56.095 36.325 56.245 ;
        RECT 34.635 55.595 35.620 55.955 ;
        RECT 35.790 55.765 36.325 56.095 ;
        RECT 34.635 55.575 35.920 55.595 ;
        RECT 34.285 55.320 34.495 55.455 ;
        RECT 35.060 55.425 35.920 55.575 ;
        RECT 30.180 54.265 30.480 55.065 ;
        RECT 30.650 54.435 30.980 55.235 ;
        RECT 31.150 54.265 31.320 55.065 ;
        RECT 31.490 54.435 31.820 55.235 ;
        RECT 31.990 54.265 32.160 55.065 ;
        RECT 32.330 54.435 32.660 55.235 ;
        RECT 32.830 54.265 33.000 55.065 ;
        RECT 33.170 54.435 33.500 55.235 ;
        RECT 33.670 54.265 33.925 55.065 ;
        RECT 34.285 54.535 34.590 55.320 ;
        RECT 34.765 54.945 35.460 55.255 ;
        RECT 34.770 54.265 35.455 54.735 ;
        RECT 35.635 54.480 35.920 55.425 ;
        RECT 36.090 55.115 36.325 55.765 ;
        RECT 36.495 55.285 36.795 56.135 ;
        RECT 37.945 56.090 38.235 56.815 ;
        RECT 38.405 56.165 38.665 56.645 ;
        RECT 38.835 56.275 39.085 56.815 ;
        RECT 36.090 54.885 36.765 55.115 ;
        RECT 36.095 54.265 36.425 54.715 ;
        RECT 36.595 54.455 36.765 54.885 ;
        RECT 37.945 54.265 38.235 55.430 ;
        RECT 38.405 55.135 38.575 56.165 ;
        RECT 39.255 56.135 39.475 56.595 ;
        RECT 39.225 56.110 39.475 56.135 ;
        RECT 38.745 55.515 38.975 55.910 ;
        RECT 39.145 55.685 39.475 56.110 ;
        RECT 39.645 56.435 40.535 56.605 ;
        RECT 39.645 55.710 39.815 56.435 ;
        RECT 39.985 55.880 40.535 56.265 ;
        RECT 41.215 56.160 41.545 56.595 ;
        RECT 41.715 56.205 41.885 56.815 ;
        RECT 41.165 56.075 41.545 56.160 ;
        RECT 42.055 56.075 42.385 56.600 ;
        RECT 42.645 56.285 42.855 56.815 ;
        RECT 43.130 56.365 43.915 56.535 ;
        RECT 44.085 56.365 44.490 56.535 ;
        RECT 41.165 56.035 41.390 56.075 ;
        RECT 39.645 55.640 40.535 55.710 ;
        RECT 39.640 55.615 40.535 55.640 ;
        RECT 39.630 55.600 40.535 55.615 ;
        RECT 39.625 55.585 40.535 55.600 ;
        RECT 39.615 55.580 40.535 55.585 ;
        RECT 39.610 55.570 40.535 55.580 ;
        RECT 39.605 55.560 40.535 55.570 ;
        RECT 39.595 55.555 40.535 55.560 ;
        RECT 39.585 55.545 40.535 55.555 ;
        RECT 39.575 55.540 40.535 55.545 ;
        RECT 39.575 55.535 39.910 55.540 ;
        RECT 39.560 55.530 39.910 55.535 ;
        RECT 39.545 55.520 39.910 55.530 ;
        RECT 39.520 55.515 39.910 55.520 ;
        RECT 38.745 55.510 39.910 55.515 ;
        RECT 38.745 55.475 39.880 55.510 ;
        RECT 38.745 55.450 39.845 55.475 ;
        RECT 38.745 55.420 39.815 55.450 ;
        RECT 38.745 55.390 39.795 55.420 ;
        RECT 38.745 55.360 39.775 55.390 ;
        RECT 38.745 55.350 39.705 55.360 ;
        RECT 38.745 55.340 39.680 55.350 ;
        RECT 38.745 55.325 39.660 55.340 ;
        RECT 38.745 55.310 39.640 55.325 ;
        RECT 38.850 55.300 39.635 55.310 ;
        RECT 38.850 55.265 39.620 55.300 ;
        RECT 38.405 54.435 38.680 55.135 ;
        RECT 38.850 55.015 39.605 55.265 ;
        RECT 39.775 54.945 40.105 55.190 ;
        RECT 40.275 55.090 40.535 55.540 ;
        RECT 41.165 55.455 41.335 56.035 ;
        RECT 42.055 55.905 42.255 56.075 ;
        RECT 43.130 55.905 43.300 56.365 ;
        RECT 41.505 55.575 42.255 55.905 ;
        RECT 42.425 55.575 43.300 55.905 ;
        RECT 41.165 55.405 41.380 55.455 ;
        RECT 41.165 55.325 41.555 55.405 ;
        RECT 39.920 54.920 40.105 54.945 ;
        RECT 39.920 54.820 40.535 54.920 ;
        RECT 38.850 54.265 39.105 54.810 ;
        RECT 39.275 54.435 39.755 54.775 ;
        RECT 39.930 54.265 40.535 54.820 ;
        RECT 41.225 54.480 41.555 55.325 ;
        RECT 42.065 55.370 42.255 55.575 ;
        RECT 41.725 54.265 41.895 55.275 ;
        RECT 42.065 54.995 42.960 55.370 ;
        RECT 42.065 54.435 42.405 54.995 ;
        RECT 42.635 54.265 42.950 54.765 ;
        RECT 43.130 54.735 43.300 55.575 ;
        RECT 43.470 55.865 43.935 56.195 ;
        RECT 44.320 56.135 44.490 56.365 ;
        RECT 44.670 56.315 45.040 56.815 ;
        RECT 45.360 56.365 46.035 56.535 ;
        RECT 46.230 56.365 46.565 56.535 ;
        RECT 43.470 54.905 43.790 55.865 ;
        RECT 44.320 55.835 45.150 56.135 ;
        RECT 43.960 54.935 44.150 55.655 ;
        RECT 44.320 54.765 44.490 55.835 ;
        RECT 44.950 55.805 45.150 55.835 ;
        RECT 44.660 55.585 44.830 55.655 ;
        RECT 45.360 55.585 45.530 56.365 ;
        RECT 46.395 56.225 46.565 56.365 ;
        RECT 46.735 56.355 46.985 56.815 ;
        RECT 44.660 55.415 45.530 55.585 ;
        RECT 45.700 55.945 46.225 56.165 ;
        RECT 46.395 56.095 46.620 56.225 ;
        RECT 44.660 55.325 45.170 55.415 ;
        RECT 43.130 54.565 44.015 54.735 ;
        RECT 44.240 54.435 44.490 54.765 ;
        RECT 44.660 54.265 44.830 55.065 ;
        RECT 45.000 54.710 45.170 55.325 ;
        RECT 45.700 55.245 45.870 55.945 ;
        RECT 45.340 54.880 45.870 55.245 ;
        RECT 46.040 55.180 46.280 55.775 ;
        RECT 46.450 54.990 46.620 56.095 ;
        RECT 46.790 55.235 47.070 56.185 ;
        RECT 46.315 54.860 46.620 54.990 ;
        RECT 45.000 54.540 46.105 54.710 ;
        RECT 46.315 54.435 46.565 54.860 ;
        RECT 46.735 54.265 47.000 54.725 ;
        RECT 47.240 54.435 47.425 56.555 ;
        RECT 47.595 56.435 47.925 56.815 ;
        RECT 48.095 56.265 48.265 56.555 ;
        RECT 47.600 56.095 48.265 56.265 ;
        RECT 48.640 56.185 48.925 56.645 ;
        RECT 49.095 56.355 49.365 56.815 ;
        RECT 47.600 55.105 47.830 56.095 ;
        RECT 48.640 56.015 49.595 56.185 ;
        RECT 48.000 55.275 48.350 55.925 ;
        RECT 48.525 55.285 49.215 55.845 ;
        RECT 49.385 55.115 49.595 56.015 ;
        RECT 47.600 54.935 48.265 55.105 ;
        RECT 47.595 54.265 47.925 54.765 ;
        RECT 48.095 54.435 48.265 54.935 ;
        RECT 48.640 54.895 49.595 55.115 ;
        RECT 49.765 55.845 50.165 56.645 ;
        RECT 50.355 56.185 50.635 56.645 ;
        RECT 51.155 56.355 51.480 56.815 ;
        RECT 50.355 56.015 51.480 56.185 ;
        RECT 51.650 56.075 52.035 56.645 ;
        RECT 51.030 55.905 51.480 56.015 ;
        RECT 49.765 55.285 50.860 55.845 ;
        RECT 51.030 55.575 51.585 55.905 ;
        RECT 48.640 54.435 48.925 54.895 ;
        RECT 49.095 54.265 49.365 54.725 ;
        RECT 49.765 54.435 50.165 55.285 ;
        RECT 51.030 55.115 51.480 55.575 ;
        RECT 51.755 55.405 52.035 56.075 ;
        RECT 50.355 54.895 51.480 55.115 ;
        RECT 50.355 54.435 50.635 54.895 ;
        RECT 51.155 54.265 51.480 54.725 ;
        RECT 51.650 54.435 52.035 55.405 ;
        RECT 52.205 55.870 52.545 56.645 ;
        RECT 52.715 56.355 52.885 56.815 ;
        RECT 53.125 56.380 53.485 56.645 ;
        RECT 53.125 56.375 53.480 56.380 ;
        RECT 53.125 56.365 53.475 56.375 ;
        RECT 53.125 56.360 53.470 56.365 ;
        RECT 53.125 56.350 53.465 56.360 ;
        RECT 54.115 56.355 54.285 56.815 ;
        RECT 53.125 56.345 53.460 56.350 ;
        RECT 53.125 56.335 53.450 56.345 ;
        RECT 53.125 56.325 53.440 56.335 ;
        RECT 53.125 56.185 53.425 56.325 ;
        RECT 52.715 55.995 53.425 56.185 ;
        RECT 53.615 56.185 53.945 56.265 ;
        RECT 54.455 56.185 54.795 56.645 ;
        RECT 53.615 55.995 54.795 56.185 ;
        RECT 55.515 56.265 55.685 56.555 ;
        RECT 55.855 56.435 56.185 56.815 ;
        RECT 55.515 56.095 56.180 56.265 ;
        RECT 52.205 54.435 52.485 55.870 ;
        RECT 52.715 55.425 53.000 55.995 ;
        RECT 53.185 55.595 53.655 55.825 ;
        RECT 53.825 55.805 54.155 55.825 ;
        RECT 53.825 55.625 54.275 55.805 ;
        RECT 54.465 55.625 54.795 55.825 ;
        RECT 52.715 55.210 53.865 55.425 ;
        RECT 52.655 54.265 53.365 55.040 ;
        RECT 53.535 54.435 53.865 55.210 ;
        RECT 54.060 54.510 54.275 55.625 ;
        RECT 54.565 55.285 54.795 55.625 ;
        RECT 55.430 55.275 55.780 55.925 ;
        RECT 55.950 55.105 56.180 56.095 ;
        RECT 54.455 54.265 54.785 54.985 ;
        RECT 55.515 54.935 56.180 55.105 ;
        RECT 55.515 54.435 55.685 54.935 ;
        RECT 55.855 54.265 56.185 54.765 ;
        RECT 56.355 54.435 56.540 56.555 ;
        RECT 56.795 56.355 57.045 56.815 ;
        RECT 57.215 56.365 57.550 56.535 ;
        RECT 57.745 56.365 58.420 56.535 ;
        RECT 57.215 56.225 57.385 56.365 ;
        RECT 56.710 55.235 56.990 56.185 ;
        RECT 57.160 56.095 57.385 56.225 ;
        RECT 57.160 54.990 57.330 56.095 ;
        RECT 57.555 55.945 58.080 56.165 ;
        RECT 57.500 55.180 57.740 55.775 ;
        RECT 57.910 55.245 58.080 55.945 ;
        RECT 58.250 55.585 58.420 56.365 ;
        RECT 58.740 56.315 59.110 56.815 ;
        RECT 59.290 56.365 59.695 56.535 ;
        RECT 59.865 56.365 60.650 56.535 ;
        RECT 59.290 56.135 59.460 56.365 ;
        RECT 58.630 55.835 59.460 56.135 ;
        RECT 59.845 55.865 60.310 56.195 ;
        RECT 58.630 55.805 58.830 55.835 ;
        RECT 58.950 55.585 59.120 55.655 ;
        RECT 58.250 55.415 59.120 55.585 ;
        RECT 58.610 55.325 59.120 55.415 ;
        RECT 57.160 54.860 57.465 54.990 ;
        RECT 57.910 54.880 58.440 55.245 ;
        RECT 56.780 54.265 57.045 54.725 ;
        RECT 57.215 54.435 57.465 54.860 ;
        RECT 58.610 54.710 58.780 55.325 ;
        RECT 57.675 54.540 58.780 54.710 ;
        RECT 58.950 54.265 59.120 55.065 ;
        RECT 59.290 54.765 59.460 55.835 ;
        RECT 59.630 54.935 59.820 55.655 ;
        RECT 59.990 54.905 60.310 55.865 ;
        RECT 60.480 55.905 60.650 56.365 ;
        RECT 60.925 56.285 61.135 56.815 ;
        RECT 61.395 56.075 61.725 56.600 ;
        RECT 61.895 56.205 62.065 56.815 ;
        RECT 62.235 56.160 62.565 56.595 ;
        RECT 62.735 56.300 62.905 56.815 ;
        RECT 62.235 56.075 62.615 56.160 ;
        RECT 63.705 56.090 63.995 56.815 ;
        RECT 64.255 56.265 64.425 56.555 ;
        RECT 64.595 56.435 64.925 56.815 ;
        RECT 64.255 56.095 64.920 56.265 ;
        RECT 61.525 55.905 61.725 56.075 ;
        RECT 62.390 56.035 62.615 56.075 ;
        RECT 60.480 55.575 61.355 55.905 ;
        RECT 61.525 55.575 62.275 55.905 ;
        RECT 59.290 54.435 59.540 54.765 ;
        RECT 60.480 54.735 60.650 55.575 ;
        RECT 61.525 55.370 61.715 55.575 ;
        RECT 62.445 55.455 62.615 56.035 ;
        RECT 62.400 55.405 62.615 55.455 ;
        RECT 60.820 54.995 61.715 55.370 ;
        RECT 62.225 55.325 62.615 55.405 ;
        RECT 59.765 54.565 60.650 54.735 ;
        RECT 60.830 54.265 61.145 54.765 ;
        RECT 61.375 54.435 61.715 54.995 ;
        RECT 61.885 54.265 62.055 55.275 ;
        RECT 62.225 54.480 62.555 55.325 ;
        RECT 62.725 54.265 62.895 55.180 ;
        RECT 63.705 54.265 63.995 55.430 ;
        RECT 64.170 55.275 64.520 55.925 ;
        RECT 64.690 55.105 64.920 56.095 ;
        RECT 64.255 54.935 64.920 55.105 ;
        RECT 64.255 54.435 64.425 54.935 ;
        RECT 64.595 54.265 64.925 54.765 ;
        RECT 65.095 54.435 65.280 56.555 ;
        RECT 65.535 56.355 65.785 56.815 ;
        RECT 65.955 56.365 66.290 56.535 ;
        RECT 66.485 56.365 67.160 56.535 ;
        RECT 65.955 56.225 66.125 56.365 ;
        RECT 65.450 55.235 65.730 56.185 ;
        RECT 65.900 56.095 66.125 56.225 ;
        RECT 65.900 54.990 66.070 56.095 ;
        RECT 66.295 55.945 66.820 56.165 ;
        RECT 66.240 55.180 66.480 55.775 ;
        RECT 66.650 55.245 66.820 55.945 ;
        RECT 66.990 55.585 67.160 56.365 ;
        RECT 67.480 56.315 67.850 56.815 ;
        RECT 68.030 56.365 68.435 56.535 ;
        RECT 68.605 56.365 69.390 56.535 ;
        RECT 68.030 56.135 68.200 56.365 ;
        RECT 67.370 55.835 68.200 56.135 ;
        RECT 68.585 55.865 69.050 56.195 ;
        RECT 67.370 55.805 67.570 55.835 ;
        RECT 67.690 55.585 67.860 55.655 ;
        RECT 66.990 55.415 67.860 55.585 ;
        RECT 67.350 55.325 67.860 55.415 ;
        RECT 65.900 54.860 66.205 54.990 ;
        RECT 66.650 54.880 67.180 55.245 ;
        RECT 65.520 54.265 65.785 54.725 ;
        RECT 65.955 54.435 66.205 54.860 ;
        RECT 67.350 54.710 67.520 55.325 ;
        RECT 66.415 54.540 67.520 54.710 ;
        RECT 67.690 54.265 67.860 55.065 ;
        RECT 68.030 54.765 68.200 55.835 ;
        RECT 68.370 54.935 68.560 55.655 ;
        RECT 68.730 54.905 69.050 55.865 ;
        RECT 69.220 55.905 69.390 56.365 ;
        RECT 69.665 56.285 69.875 56.815 ;
        RECT 70.135 56.075 70.465 56.600 ;
        RECT 70.635 56.205 70.805 56.815 ;
        RECT 70.975 56.160 71.305 56.595 ;
        RECT 71.475 56.300 71.645 56.815 ;
        RECT 72.075 56.265 72.245 56.555 ;
        RECT 72.415 56.435 72.745 56.815 ;
        RECT 70.975 56.075 71.355 56.160 ;
        RECT 72.075 56.095 72.740 56.265 ;
        RECT 70.265 55.905 70.465 56.075 ;
        RECT 71.130 56.035 71.355 56.075 ;
        RECT 69.220 55.575 70.095 55.905 ;
        RECT 70.265 55.575 71.015 55.905 ;
        RECT 68.030 54.435 68.280 54.765 ;
        RECT 69.220 54.735 69.390 55.575 ;
        RECT 70.265 55.370 70.455 55.575 ;
        RECT 71.185 55.455 71.355 56.035 ;
        RECT 71.140 55.405 71.355 55.455 ;
        RECT 69.560 54.995 70.455 55.370 ;
        RECT 70.965 55.325 71.355 55.405 ;
        RECT 68.505 54.565 69.390 54.735 ;
        RECT 69.570 54.265 69.885 54.765 ;
        RECT 70.115 54.435 70.455 54.995 ;
        RECT 70.625 54.265 70.795 55.275 ;
        RECT 70.965 54.480 71.295 55.325 ;
        RECT 71.990 55.275 72.340 55.925 ;
        RECT 71.465 54.265 71.635 55.180 ;
        RECT 72.510 55.105 72.740 56.095 ;
        RECT 72.075 54.935 72.740 55.105 ;
        RECT 72.075 54.435 72.245 54.935 ;
        RECT 72.415 54.265 72.745 54.765 ;
        RECT 72.915 54.435 73.100 56.555 ;
        RECT 73.355 56.355 73.605 56.815 ;
        RECT 73.775 56.365 74.110 56.535 ;
        RECT 74.305 56.365 74.980 56.535 ;
        RECT 73.775 56.225 73.945 56.365 ;
        RECT 73.270 55.235 73.550 56.185 ;
        RECT 73.720 56.095 73.945 56.225 ;
        RECT 73.720 54.990 73.890 56.095 ;
        RECT 74.115 55.945 74.640 56.165 ;
        RECT 74.060 55.180 74.300 55.775 ;
        RECT 74.470 55.245 74.640 55.945 ;
        RECT 74.810 55.585 74.980 56.365 ;
        RECT 75.300 56.315 75.670 56.815 ;
        RECT 75.850 56.365 76.255 56.535 ;
        RECT 76.425 56.365 77.210 56.535 ;
        RECT 75.850 56.135 76.020 56.365 ;
        RECT 75.190 55.835 76.020 56.135 ;
        RECT 76.405 55.865 76.870 56.195 ;
        RECT 75.190 55.805 75.390 55.835 ;
        RECT 75.510 55.585 75.680 55.655 ;
        RECT 74.810 55.415 75.680 55.585 ;
        RECT 75.170 55.325 75.680 55.415 ;
        RECT 73.720 54.860 74.025 54.990 ;
        RECT 74.470 54.880 75.000 55.245 ;
        RECT 73.340 54.265 73.605 54.725 ;
        RECT 73.775 54.435 74.025 54.860 ;
        RECT 75.170 54.710 75.340 55.325 ;
        RECT 74.235 54.540 75.340 54.710 ;
        RECT 75.510 54.265 75.680 55.065 ;
        RECT 75.850 54.765 76.020 55.835 ;
        RECT 76.190 54.935 76.380 55.655 ;
        RECT 76.550 54.905 76.870 55.865 ;
        RECT 77.040 55.905 77.210 56.365 ;
        RECT 77.485 56.285 77.695 56.815 ;
        RECT 77.955 56.075 78.285 56.600 ;
        RECT 78.455 56.205 78.625 56.815 ;
        RECT 78.795 56.160 79.125 56.595 ;
        RECT 79.345 56.315 79.605 56.645 ;
        RECT 79.775 56.455 80.105 56.815 ;
        RECT 80.360 56.435 81.660 56.645 ;
        RECT 78.795 56.075 79.175 56.160 ;
        RECT 78.085 55.905 78.285 56.075 ;
        RECT 78.950 56.035 79.175 56.075 ;
        RECT 77.040 55.575 77.915 55.905 ;
        RECT 78.085 55.575 78.835 55.905 ;
        RECT 75.850 54.435 76.100 54.765 ;
        RECT 77.040 54.735 77.210 55.575 ;
        RECT 78.085 55.370 78.275 55.575 ;
        RECT 79.005 55.455 79.175 56.035 ;
        RECT 78.960 55.405 79.175 55.455 ;
        RECT 77.380 54.995 78.275 55.370 ;
        RECT 78.785 55.325 79.175 55.405 ;
        RECT 76.325 54.565 77.210 54.735 ;
        RECT 77.390 54.265 77.705 54.765 ;
        RECT 77.935 54.435 78.275 54.995 ;
        RECT 78.445 54.265 78.615 55.275 ;
        RECT 78.785 54.480 79.115 55.325 ;
        RECT 79.345 55.115 79.515 56.315 ;
        RECT 80.360 56.285 80.530 56.435 ;
        RECT 79.775 56.160 80.530 56.285 ;
        RECT 79.685 56.115 80.530 56.160 ;
        RECT 79.685 55.995 79.955 56.115 ;
        RECT 79.685 55.420 79.855 55.995 ;
        RECT 80.085 55.555 80.495 55.860 ;
        RECT 80.785 55.825 80.995 56.225 ;
        RECT 80.665 55.615 80.995 55.825 ;
        RECT 81.240 55.825 81.460 56.225 ;
        RECT 81.935 56.050 82.390 56.815 ;
        RECT 83.650 56.305 83.890 56.815 ;
        RECT 84.070 56.305 84.350 56.635 ;
        RECT 84.580 56.305 84.795 56.815 ;
        RECT 81.240 55.615 81.715 55.825 ;
        RECT 81.905 55.625 82.395 55.825 ;
        RECT 83.545 55.575 83.900 56.135 ;
        RECT 79.685 55.385 79.885 55.420 ;
        RECT 81.215 55.385 82.390 55.445 ;
        RECT 84.070 55.405 84.240 56.305 ;
        RECT 84.410 55.575 84.675 56.135 ;
        RECT 84.965 56.075 85.580 56.645 ;
        RECT 85.950 56.305 86.190 56.815 ;
        RECT 86.370 56.305 86.650 56.635 ;
        RECT 86.880 56.305 87.095 56.815 ;
        RECT 84.925 55.405 85.095 55.905 ;
        RECT 79.685 55.275 82.390 55.385 ;
        RECT 79.745 55.215 81.545 55.275 ;
        RECT 81.215 55.185 81.545 55.215 ;
        RECT 79.345 54.435 79.605 55.115 ;
        RECT 79.775 54.265 80.025 55.045 ;
        RECT 80.275 55.015 81.110 55.025 ;
        RECT 81.700 55.015 81.885 55.105 ;
        RECT 80.275 54.815 81.885 55.015 ;
        RECT 80.275 54.435 80.525 54.815 ;
        RECT 81.655 54.775 81.885 54.815 ;
        RECT 82.135 54.655 82.390 55.275 ;
        RECT 83.670 55.235 85.095 55.405 ;
        RECT 83.670 55.060 84.060 55.235 ;
        RECT 80.695 54.265 81.050 54.645 ;
        RECT 82.055 54.435 82.390 54.655 ;
        RECT 84.545 54.265 84.875 55.065 ;
        RECT 85.265 55.055 85.580 56.075 ;
        RECT 85.845 55.575 86.200 56.135 ;
        RECT 86.370 55.405 86.540 56.305 ;
        RECT 86.710 55.575 86.975 56.135 ;
        RECT 87.265 56.075 87.880 56.645 ;
        RECT 87.225 55.405 87.395 55.905 ;
        RECT 85.970 55.235 87.395 55.405 ;
        RECT 85.970 55.060 86.360 55.235 ;
        RECT 85.045 54.435 85.580 55.055 ;
        RECT 86.845 54.265 87.175 55.065 ;
        RECT 87.565 55.055 87.880 56.075 ;
        RECT 88.545 56.065 89.755 56.815 ;
        RECT 87.345 54.435 87.880 55.055 ;
        RECT 88.545 55.355 89.065 55.895 ;
        RECT 89.235 55.525 89.755 56.065 ;
        RECT 88.545 54.265 89.755 55.355 ;
        RECT 12.100 54.095 89.840 54.265 ;
        RECT 12.185 53.005 13.395 54.095 ;
        RECT 13.565 53.005 15.235 54.095 ;
        RECT 12.185 52.295 12.705 52.835 ;
        RECT 12.875 52.465 13.395 53.005 ;
        RECT 13.565 52.315 14.315 52.835 ;
        RECT 14.485 52.485 15.235 53.005 ;
        RECT 15.405 53.225 15.680 53.925 ;
        RECT 15.850 53.550 16.105 54.095 ;
        RECT 16.275 53.585 16.755 53.925 ;
        RECT 16.930 53.540 17.535 54.095 ;
        RECT 16.920 53.440 17.535 53.540 ;
        RECT 17.715 53.485 18.045 53.915 ;
        RECT 18.225 53.655 18.420 54.095 ;
        RECT 18.590 53.485 18.920 53.915 ;
        RECT 16.920 53.415 17.105 53.440 ;
        RECT 12.185 51.545 13.395 52.295 ;
        RECT 13.565 51.545 15.235 52.315 ;
        RECT 15.405 52.195 15.575 53.225 ;
        RECT 15.850 53.095 16.605 53.345 ;
        RECT 16.775 53.170 17.105 53.415 ;
        RECT 17.715 53.315 18.920 53.485 ;
        RECT 15.850 53.060 16.620 53.095 ;
        RECT 15.850 53.050 16.635 53.060 ;
        RECT 15.745 53.035 16.640 53.050 ;
        RECT 15.745 53.020 16.660 53.035 ;
        RECT 15.745 53.010 16.680 53.020 ;
        RECT 15.745 53.000 16.705 53.010 ;
        RECT 15.745 52.970 16.775 53.000 ;
        RECT 15.745 52.940 16.795 52.970 ;
        RECT 15.745 52.910 16.815 52.940 ;
        RECT 15.745 52.885 16.845 52.910 ;
        RECT 15.745 52.850 16.880 52.885 ;
        RECT 15.745 52.845 16.910 52.850 ;
        RECT 15.745 52.450 15.975 52.845 ;
        RECT 16.520 52.840 16.910 52.845 ;
        RECT 16.545 52.830 16.910 52.840 ;
        RECT 16.560 52.825 16.910 52.830 ;
        RECT 16.575 52.820 16.910 52.825 ;
        RECT 17.275 52.820 17.535 53.270 ;
        RECT 17.715 52.985 18.610 53.315 ;
        RECT 19.090 53.145 19.365 53.915 ;
        RECT 16.575 52.815 17.535 52.820 ;
        RECT 16.585 52.805 17.535 52.815 ;
        RECT 16.595 52.800 17.535 52.805 ;
        RECT 16.605 52.790 17.535 52.800 ;
        RECT 16.610 52.780 17.535 52.790 ;
        RECT 18.780 52.955 19.365 53.145 ;
        RECT 19.545 53.005 22.135 54.095 ;
        RECT 16.615 52.775 17.535 52.780 ;
        RECT 16.625 52.760 17.535 52.775 ;
        RECT 16.630 52.745 17.535 52.760 ;
        RECT 16.640 52.720 17.535 52.745 ;
        RECT 16.145 52.250 16.475 52.675 ;
        RECT 16.225 52.225 16.475 52.250 ;
        RECT 15.405 51.715 15.665 52.195 ;
        RECT 15.835 51.545 16.085 52.085 ;
        RECT 16.255 51.765 16.475 52.225 ;
        RECT 16.645 52.650 17.535 52.720 ;
        RECT 16.645 51.925 16.815 52.650 ;
        RECT 16.985 52.095 17.535 52.480 ;
        RECT 17.720 52.455 18.015 52.785 ;
        RECT 18.195 52.455 18.610 52.785 ;
        RECT 16.645 51.755 17.535 51.925 ;
        RECT 17.715 51.545 18.015 52.275 ;
        RECT 18.195 51.835 18.425 52.455 ;
        RECT 18.780 52.285 18.955 52.955 ;
        RECT 18.625 52.105 18.955 52.285 ;
        RECT 19.125 52.135 19.365 52.785 ;
        RECT 19.545 52.315 20.755 52.835 ;
        RECT 20.925 52.485 22.135 53.005 ;
        RECT 22.950 53.125 23.340 53.300 ;
        RECT 23.825 53.295 24.155 54.095 ;
        RECT 24.325 53.305 24.860 53.925 ;
        RECT 22.950 52.955 24.375 53.125 ;
        RECT 18.625 51.725 18.850 52.105 ;
        RECT 19.020 51.545 19.350 51.935 ;
        RECT 19.545 51.545 22.135 52.315 ;
        RECT 22.825 52.225 23.180 52.785 ;
        RECT 23.350 52.055 23.520 52.955 ;
        RECT 23.690 52.225 23.955 52.785 ;
        RECT 24.205 52.455 24.375 52.955 ;
        RECT 24.545 52.285 24.860 53.305 ;
        RECT 25.065 52.930 25.355 54.095 ;
        RECT 25.530 53.585 27.185 53.875 ;
        RECT 25.530 53.245 27.120 53.415 ;
        RECT 27.355 53.295 27.635 54.095 ;
        RECT 25.530 52.955 25.850 53.245 ;
        RECT 26.950 53.125 27.120 53.245 ;
        RECT 22.930 51.545 23.170 52.055 ;
        RECT 23.350 51.725 23.630 52.055 ;
        RECT 23.860 51.545 24.075 52.055 ;
        RECT 24.245 51.715 24.860 52.285 ;
        RECT 25.065 51.545 25.355 52.270 ;
        RECT 25.530 52.215 25.880 52.785 ;
        RECT 26.050 52.455 26.760 53.075 ;
        RECT 26.950 52.955 27.675 53.125 ;
        RECT 27.845 52.955 28.115 53.925 ;
        RECT 27.505 52.785 27.675 52.955 ;
        RECT 26.930 52.455 27.335 52.785 ;
        RECT 27.505 52.455 27.775 52.785 ;
        RECT 27.505 52.285 27.675 52.455 ;
        RECT 26.065 52.115 27.675 52.285 ;
        RECT 27.945 52.220 28.115 52.955 ;
        RECT 25.535 51.545 25.865 52.045 ;
        RECT 26.065 51.765 26.235 52.115 ;
        RECT 26.435 51.545 26.765 51.945 ;
        RECT 26.935 51.765 27.105 52.115 ;
        RECT 27.275 51.545 27.655 51.945 ;
        RECT 27.845 51.875 28.115 52.220 ;
        RECT 29.205 51.825 29.485 53.925 ;
        RECT 29.675 53.335 30.460 54.095 ;
        RECT 30.855 53.265 31.240 53.925 ;
        RECT 30.855 53.165 31.265 53.265 ;
        RECT 29.655 52.955 31.265 53.165 ;
        RECT 31.565 53.075 31.765 53.865 ;
        RECT 29.655 52.355 29.930 52.955 ;
        RECT 31.435 52.905 31.765 53.075 ;
        RECT 31.935 52.915 32.255 54.095 ;
        RECT 32.885 53.260 33.230 54.095 ;
        RECT 33.405 53.090 33.660 53.895 ;
        RECT 33.830 53.260 34.090 54.095 ;
        RECT 34.265 53.090 34.520 53.895 ;
        RECT 34.690 53.260 34.950 54.095 ;
        RECT 35.120 53.090 35.380 53.895 ;
        RECT 35.550 53.260 35.935 54.095 ;
        RECT 36.355 53.365 36.650 54.095 ;
        RECT 36.820 53.195 37.080 53.920 ;
        RECT 37.250 53.365 37.510 54.095 ;
        RECT 37.680 53.195 37.940 53.920 ;
        RECT 38.110 53.365 38.370 54.095 ;
        RECT 38.540 53.195 38.800 53.920 ;
        RECT 38.970 53.365 39.230 54.095 ;
        RECT 39.400 53.195 39.660 53.920 ;
        RECT 32.905 52.920 35.935 53.090 ;
        RECT 31.435 52.785 31.615 52.905 ;
        RECT 30.100 52.535 30.455 52.785 ;
        RECT 30.650 52.735 31.115 52.785 ;
        RECT 30.645 52.565 31.115 52.735 ;
        RECT 30.650 52.535 31.115 52.565 ;
        RECT 31.285 52.535 31.615 52.785 ;
        RECT 31.790 52.535 32.255 52.735 ;
        RECT 32.905 52.355 33.075 52.920 ;
        RECT 33.245 52.525 35.460 52.750 ;
        RECT 35.635 52.355 35.935 52.920 ;
        RECT 29.655 52.175 30.905 52.355 ;
        RECT 30.540 52.105 30.905 52.175 ;
        RECT 31.075 52.155 32.255 52.325 ;
        RECT 32.905 52.185 35.935 52.355 ;
        RECT 36.350 52.955 39.660 53.195 ;
        RECT 39.830 52.985 40.090 54.095 ;
        RECT 36.350 52.365 37.320 52.955 ;
        RECT 40.260 52.785 40.510 53.920 ;
        RECT 40.690 52.985 40.985 54.095 ;
        RECT 41.255 53.425 41.425 53.925 ;
        RECT 41.595 53.595 41.925 54.095 ;
        RECT 41.255 53.255 41.920 53.425 ;
        RECT 37.490 52.535 40.510 52.785 ;
        RECT 36.350 52.195 39.660 52.365 ;
        RECT 29.715 51.545 29.885 52.005 ;
        RECT 31.075 51.935 31.405 52.155 ;
        RECT 30.155 51.755 31.405 51.935 ;
        RECT 31.575 51.545 31.745 51.985 ;
        RECT 31.915 51.740 32.255 52.155 ;
        RECT 33.365 51.545 33.660 52.015 ;
        RECT 33.830 51.740 34.090 52.185 ;
        RECT 34.260 51.545 34.520 52.015 ;
        RECT 34.690 51.740 34.945 52.185 ;
        RECT 35.115 51.545 35.415 52.015 ;
        RECT 36.350 51.545 36.650 52.025 ;
        RECT 36.820 51.740 37.080 52.195 ;
        RECT 37.250 51.545 37.510 52.025 ;
        RECT 37.680 51.740 37.940 52.195 ;
        RECT 38.110 51.545 38.370 52.025 ;
        RECT 38.540 51.740 38.800 52.195 ;
        RECT 38.970 51.545 39.230 52.025 ;
        RECT 39.400 51.740 39.660 52.195 ;
        RECT 39.830 51.545 40.090 52.070 ;
        RECT 40.260 51.725 40.510 52.535 ;
        RECT 40.680 52.175 40.995 52.785 ;
        RECT 41.170 52.435 41.520 53.085 ;
        RECT 41.690 52.265 41.920 53.255 ;
        RECT 41.255 52.095 41.920 52.265 ;
        RECT 40.690 51.545 40.935 52.005 ;
        RECT 41.255 51.805 41.425 52.095 ;
        RECT 41.595 51.545 41.925 51.925 ;
        RECT 42.095 51.805 42.280 53.925 ;
        RECT 42.520 53.635 42.785 54.095 ;
        RECT 42.955 53.500 43.205 53.925 ;
        RECT 43.415 53.650 44.520 53.820 ;
        RECT 42.900 53.370 43.205 53.500 ;
        RECT 42.450 52.175 42.730 53.125 ;
        RECT 42.900 52.265 43.070 53.370 ;
        RECT 43.240 52.585 43.480 53.180 ;
        RECT 43.650 53.115 44.180 53.480 ;
        RECT 43.650 52.415 43.820 53.115 ;
        RECT 44.350 53.035 44.520 53.650 ;
        RECT 44.690 53.295 44.860 54.095 ;
        RECT 45.030 53.595 45.280 53.925 ;
        RECT 45.505 53.625 46.390 53.795 ;
        RECT 44.350 52.945 44.860 53.035 ;
        RECT 42.900 52.135 43.125 52.265 ;
        RECT 43.295 52.195 43.820 52.415 ;
        RECT 43.990 52.775 44.860 52.945 ;
        RECT 42.535 51.545 42.785 52.005 ;
        RECT 42.955 51.995 43.125 52.135 ;
        RECT 43.990 51.995 44.160 52.775 ;
        RECT 44.690 52.705 44.860 52.775 ;
        RECT 44.370 52.525 44.570 52.555 ;
        RECT 45.030 52.525 45.200 53.595 ;
        RECT 45.370 52.705 45.560 53.425 ;
        RECT 44.370 52.225 45.200 52.525 ;
        RECT 45.730 52.495 46.050 53.455 ;
        RECT 42.955 51.825 43.290 51.995 ;
        RECT 43.485 51.825 44.160 51.995 ;
        RECT 44.480 51.545 44.850 52.045 ;
        RECT 45.030 51.995 45.200 52.225 ;
        RECT 45.585 52.165 46.050 52.495 ;
        RECT 46.220 52.785 46.390 53.625 ;
        RECT 46.570 53.595 46.885 54.095 ;
        RECT 47.115 53.365 47.455 53.925 ;
        RECT 46.560 52.990 47.455 53.365 ;
        RECT 47.625 53.085 47.795 54.095 ;
        RECT 47.265 52.785 47.455 52.990 ;
        RECT 47.965 53.035 48.295 53.880 ;
        RECT 48.525 53.540 49.130 54.095 ;
        RECT 49.305 53.585 49.785 53.925 ;
        RECT 49.955 53.550 50.210 54.095 ;
        RECT 48.525 53.440 49.140 53.540 ;
        RECT 48.955 53.415 49.140 53.440 ;
        RECT 47.965 52.955 48.355 53.035 ;
        RECT 48.140 52.905 48.355 52.955 ;
        RECT 46.220 52.455 47.095 52.785 ;
        RECT 47.265 52.455 48.015 52.785 ;
        RECT 46.220 51.995 46.390 52.455 ;
        RECT 47.265 52.285 47.465 52.455 ;
        RECT 48.185 52.325 48.355 52.905 ;
        RECT 48.525 52.820 48.785 53.270 ;
        RECT 48.955 53.170 49.285 53.415 ;
        RECT 49.455 53.095 50.210 53.345 ;
        RECT 50.380 53.225 50.655 53.925 ;
        RECT 49.440 53.060 50.210 53.095 ;
        RECT 49.425 53.050 50.210 53.060 ;
        RECT 49.420 53.035 50.315 53.050 ;
        RECT 49.400 53.020 50.315 53.035 ;
        RECT 49.380 53.010 50.315 53.020 ;
        RECT 49.355 53.000 50.315 53.010 ;
        RECT 49.285 52.970 50.315 53.000 ;
        RECT 49.265 52.940 50.315 52.970 ;
        RECT 49.245 52.910 50.315 52.940 ;
        RECT 49.215 52.885 50.315 52.910 ;
        RECT 49.180 52.850 50.315 52.885 ;
        RECT 49.150 52.845 50.315 52.850 ;
        RECT 49.150 52.840 49.540 52.845 ;
        RECT 49.150 52.830 49.515 52.840 ;
        RECT 49.150 52.825 49.500 52.830 ;
        RECT 49.150 52.820 49.485 52.825 ;
        RECT 48.525 52.815 49.485 52.820 ;
        RECT 48.525 52.805 49.475 52.815 ;
        RECT 48.525 52.800 49.465 52.805 ;
        RECT 48.525 52.790 49.455 52.800 ;
        RECT 48.525 52.780 49.450 52.790 ;
        RECT 48.525 52.775 49.445 52.780 ;
        RECT 48.525 52.760 49.435 52.775 ;
        RECT 48.525 52.745 49.430 52.760 ;
        RECT 48.525 52.720 49.420 52.745 ;
        RECT 48.525 52.650 49.415 52.720 ;
        RECT 48.130 52.285 48.355 52.325 ;
        RECT 45.030 51.825 45.435 51.995 ;
        RECT 45.605 51.825 46.390 51.995 ;
        RECT 46.665 51.545 46.875 52.075 ;
        RECT 47.135 51.760 47.465 52.285 ;
        RECT 47.975 52.200 48.355 52.285 ;
        RECT 47.635 51.545 47.805 52.155 ;
        RECT 47.975 51.765 48.305 52.200 ;
        RECT 48.525 52.095 49.075 52.480 ;
        RECT 49.245 51.925 49.415 52.650 ;
        RECT 48.525 51.755 49.415 51.925 ;
        RECT 49.585 52.250 49.915 52.675 ;
        RECT 50.085 52.450 50.315 52.845 ;
        RECT 49.585 51.765 49.805 52.250 ;
        RECT 50.485 52.195 50.655 53.225 ;
        RECT 50.825 52.930 51.115 54.095 ;
        RECT 51.375 53.425 51.545 53.925 ;
        RECT 51.715 53.595 52.045 54.095 ;
        RECT 51.375 53.255 52.040 53.425 ;
        RECT 51.290 52.435 51.640 53.085 ;
        RECT 49.975 51.545 50.225 52.085 ;
        RECT 50.395 51.715 50.655 52.195 ;
        RECT 50.825 51.545 51.115 52.270 ;
        RECT 51.810 52.265 52.040 53.255 ;
        RECT 51.375 52.095 52.040 52.265 ;
        RECT 51.375 51.805 51.545 52.095 ;
        RECT 51.715 51.545 52.045 51.925 ;
        RECT 52.215 51.805 52.400 53.925 ;
        RECT 52.640 53.635 52.905 54.095 ;
        RECT 53.075 53.500 53.325 53.925 ;
        RECT 53.535 53.650 54.640 53.820 ;
        RECT 53.020 53.370 53.325 53.500 ;
        RECT 52.570 52.175 52.850 53.125 ;
        RECT 53.020 52.265 53.190 53.370 ;
        RECT 53.360 52.585 53.600 53.180 ;
        RECT 53.770 53.115 54.300 53.480 ;
        RECT 53.770 52.415 53.940 53.115 ;
        RECT 54.470 53.035 54.640 53.650 ;
        RECT 54.810 53.295 54.980 54.095 ;
        RECT 55.150 53.595 55.400 53.925 ;
        RECT 55.625 53.625 56.510 53.795 ;
        RECT 54.470 52.945 54.980 53.035 ;
        RECT 53.020 52.135 53.245 52.265 ;
        RECT 53.415 52.195 53.940 52.415 ;
        RECT 54.110 52.775 54.980 52.945 ;
        RECT 52.655 51.545 52.905 52.005 ;
        RECT 53.075 51.995 53.245 52.135 ;
        RECT 54.110 51.995 54.280 52.775 ;
        RECT 54.810 52.705 54.980 52.775 ;
        RECT 54.490 52.525 54.690 52.555 ;
        RECT 55.150 52.525 55.320 53.595 ;
        RECT 55.490 52.705 55.680 53.425 ;
        RECT 54.490 52.225 55.320 52.525 ;
        RECT 55.850 52.495 56.170 53.455 ;
        RECT 53.075 51.825 53.410 51.995 ;
        RECT 53.605 51.825 54.280 51.995 ;
        RECT 54.600 51.545 54.970 52.045 ;
        RECT 55.150 51.995 55.320 52.225 ;
        RECT 55.705 52.165 56.170 52.495 ;
        RECT 56.340 52.785 56.510 53.625 ;
        RECT 56.690 53.595 57.005 54.095 ;
        RECT 57.235 53.365 57.575 53.925 ;
        RECT 56.680 52.990 57.575 53.365 ;
        RECT 57.745 53.085 57.915 54.095 ;
        RECT 57.385 52.785 57.575 52.990 ;
        RECT 58.085 53.035 58.415 53.880 ;
        RECT 58.895 53.365 59.190 54.095 ;
        RECT 59.360 53.195 59.620 53.920 ;
        RECT 59.790 53.365 60.050 54.095 ;
        RECT 60.220 53.195 60.480 53.920 ;
        RECT 60.650 53.365 60.910 54.095 ;
        RECT 61.080 53.195 61.340 53.920 ;
        RECT 61.510 53.365 61.770 54.095 ;
        RECT 61.940 53.195 62.200 53.920 ;
        RECT 58.085 52.955 58.475 53.035 ;
        RECT 58.260 52.905 58.475 52.955 ;
        RECT 56.340 52.455 57.215 52.785 ;
        RECT 57.385 52.455 58.135 52.785 ;
        RECT 56.340 51.995 56.510 52.455 ;
        RECT 57.385 52.285 57.585 52.455 ;
        RECT 58.305 52.325 58.475 52.905 ;
        RECT 58.250 52.285 58.475 52.325 ;
        RECT 55.150 51.825 55.555 51.995 ;
        RECT 55.725 51.825 56.510 51.995 ;
        RECT 56.785 51.545 56.995 52.075 ;
        RECT 57.255 51.760 57.585 52.285 ;
        RECT 58.095 52.200 58.475 52.285 ;
        RECT 58.890 52.955 62.200 53.195 ;
        RECT 62.370 52.985 62.630 54.095 ;
        RECT 58.890 52.365 59.860 52.955 ;
        RECT 62.800 52.785 63.050 53.920 ;
        RECT 63.230 52.985 63.525 54.095 ;
        RECT 63.710 52.955 64.045 53.925 ;
        RECT 64.215 52.955 64.385 54.095 ;
        RECT 64.555 53.755 66.585 53.925 ;
        RECT 60.030 52.535 63.050 52.785 ;
        RECT 57.755 51.545 57.925 52.155 ;
        RECT 58.095 51.765 58.425 52.200 ;
        RECT 58.890 52.195 62.200 52.365 ;
        RECT 58.890 51.545 59.190 52.025 ;
        RECT 59.360 51.740 59.620 52.195 ;
        RECT 59.790 51.545 60.050 52.025 ;
        RECT 60.220 51.740 60.480 52.195 ;
        RECT 60.650 51.545 60.910 52.025 ;
        RECT 61.080 51.740 61.340 52.195 ;
        RECT 61.510 51.545 61.770 52.025 ;
        RECT 61.940 51.740 62.200 52.195 ;
        RECT 62.370 51.545 62.630 52.070 ;
        RECT 62.800 51.725 63.050 52.535 ;
        RECT 63.220 52.175 63.535 52.785 ;
        RECT 63.710 52.285 63.880 52.955 ;
        RECT 64.555 52.785 64.725 53.755 ;
        RECT 64.050 52.455 64.305 52.785 ;
        RECT 64.530 52.455 64.725 52.785 ;
        RECT 64.895 53.415 66.020 53.585 ;
        RECT 64.135 52.285 64.305 52.455 ;
        RECT 64.895 52.285 65.065 53.415 ;
        RECT 63.230 51.545 63.475 52.005 ;
        RECT 63.710 51.715 63.965 52.285 ;
        RECT 64.135 52.115 65.065 52.285 ;
        RECT 65.235 53.075 66.245 53.245 ;
        RECT 65.235 52.275 65.405 53.075 ;
        RECT 65.610 52.395 65.885 52.875 ;
        RECT 65.605 52.225 65.885 52.395 ;
        RECT 64.890 52.080 65.065 52.115 ;
        RECT 64.135 51.545 64.465 51.945 ;
        RECT 64.890 51.715 65.420 52.080 ;
        RECT 65.610 51.715 65.885 52.225 ;
        RECT 66.055 51.715 66.245 53.075 ;
        RECT 66.415 53.090 66.585 53.755 ;
        RECT 66.755 53.335 66.925 54.095 ;
        RECT 67.160 53.335 67.675 53.745 ;
        RECT 69.015 53.365 69.310 54.095 ;
        RECT 66.415 52.900 67.165 53.090 ;
        RECT 67.335 52.525 67.675 53.335 ;
        RECT 69.480 53.195 69.740 53.920 ;
        RECT 69.910 53.365 70.170 54.095 ;
        RECT 70.340 53.195 70.600 53.920 ;
        RECT 70.770 53.365 71.030 54.095 ;
        RECT 71.200 53.195 71.460 53.920 ;
        RECT 71.630 53.365 71.890 54.095 ;
        RECT 72.060 53.195 72.320 53.920 ;
        RECT 66.445 52.355 67.675 52.525 ;
        RECT 69.010 52.955 72.320 53.195 ;
        RECT 72.490 52.985 72.750 54.095 ;
        RECT 69.010 52.365 69.980 52.955 ;
        RECT 72.920 52.785 73.170 53.920 ;
        RECT 73.350 52.985 73.645 54.095 ;
        RECT 73.825 53.585 75.015 53.875 ;
        RECT 73.845 53.245 75.015 53.415 ;
        RECT 75.185 53.295 75.465 54.095 ;
        RECT 73.845 52.955 74.170 53.245 ;
        RECT 74.845 53.125 75.015 53.245 ;
        RECT 74.340 52.785 74.535 53.075 ;
        RECT 74.845 52.955 75.505 53.125 ;
        RECT 75.675 52.955 75.950 53.925 ;
        RECT 75.335 52.785 75.505 52.955 ;
        RECT 70.150 52.535 73.170 52.785 ;
        RECT 66.425 51.545 66.935 52.080 ;
        RECT 67.155 51.750 67.400 52.355 ;
        RECT 69.010 52.195 72.320 52.365 ;
        RECT 69.010 51.545 69.310 52.025 ;
        RECT 69.480 51.740 69.740 52.195 ;
        RECT 69.910 51.545 70.170 52.025 ;
        RECT 70.340 51.740 70.600 52.195 ;
        RECT 70.770 51.545 71.030 52.025 ;
        RECT 71.200 51.740 71.460 52.195 ;
        RECT 71.630 51.545 71.890 52.025 ;
        RECT 72.060 51.740 72.320 52.195 ;
        RECT 72.490 51.545 72.750 52.070 ;
        RECT 72.920 51.725 73.170 52.535 ;
        RECT 73.340 52.175 73.655 52.785 ;
        RECT 73.825 52.455 74.170 52.785 ;
        RECT 74.340 52.455 75.165 52.785 ;
        RECT 75.335 52.455 75.610 52.785 ;
        RECT 75.335 52.285 75.505 52.455 ;
        RECT 73.840 52.115 75.505 52.285 ;
        RECT 75.780 52.220 75.950 52.955 ;
        RECT 76.585 52.930 76.875 54.095 ;
        RECT 77.080 53.305 77.615 53.925 ;
        RECT 77.080 52.285 77.395 53.305 ;
        RECT 77.785 53.295 78.115 54.095 ;
        RECT 78.600 53.125 78.990 53.300 ;
        RECT 77.565 52.955 78.990 53.125 ;
        RECT 79.345 53.005 80.555 54.095 ;
        RECT 77.565 52.455 77.735 52.955 ;
        RECT 73.350 51.545 73.595 52.005 ;
        RECT 73.840 51.765 74.095 52.115 ;
        RECT 74.265 51.545 74.595 51.945 ;
        RECT 74.765 51.765 74.935 52.115 ;
        RECT 75.105 51.545 75.485 51.945 ;
        RECT 75.675 51.875 75.950 52.220 ;
        RECT 76.585 51.545 76.875 52.270 ;
        RECT 77.080 51.715 77.695 52.285 ;
        RECT 77.985 52.225 78.250 52.785 ;
        RECT 78.420 52.055 78.590 52.955 ;
        RECT 78.760 52.225 79.115 52.785 ;
        RECT 79.345 52.295 79.865 52.835 ;
        RECT 80.035 52.465 80.555 53.005 ;
        RECT 80.725 52.955 81.065 53.925 ;
        RECT 81.235 52.955 81.405 54.095 ;
        RECT 81.675 53.295 81.925 54.095 ;
        RECT 82.570 53.125 82.900 53.925 ;
        RECT 83.200 53.295 83.530 54.095 ;
        RECT 83.700 53.125 84.030 53.925 ;
        RECT 81.595 52.955 84.030 53.125 ;
        RECT 84.440 53.305 84.975 53.925 ;
        RECT 80.725 52.345 80.900 52.955 ;
        RECT 81.595 52.705 81.765 52.955 ;
        RECT 81.070 52.535 81.765 52.705 ;
        RECT 81.940 52.535 82.360 52.735 ;
        RECT 82.530 52.535 82.860 52.735 ;
        RECT 83.030 52.535 83.360 52.735 ;
        RECT 77.865 51.545 78.080 52.055 ;
        RECT 78.310 51.725 78.590 52.055 ;
        RECT 78.770 51.545 79.010 52.055 ;
        RECT 79.345 51.545 80.555 52.295 ;
        RECT 80.725 51.715 81.065 52.345 ;
        RECT 81.235 51.545 81.485 52.345 ;
        RECT 81.675 52.195 82.900 52.365 ;
        RECT 81.675 51.715 82.005 52.195 ;
        RECT 82.175 51.545 82.400 52.005 ;
        RECT 82.570 51.715 82.900 52.195 ;
        RECT 83.530 52.325 83.700 52.955 ;
        RECT 83.885 52.535 84.235 52.785 ;
        RECT 83.530 51.715 84.030 52.325 ;
        RECT 84.440 52.285 84.755 53.305 ;
        RECT 85.145 53.295 85.475 54.095 ;
        RECT 85.960 53.125 86.350 53.300 ;
        RECT 84.925 52.955 86.350 53.125 ;
        RECT 86.795 53.165 86.965 53.925 ;
        RECT 87.180 53.335 87.510 54.095 ;
        RECT 86.795 52.995 87.510 53.165 ;
        RECT 87.680 53.020 87.935 53.925 ;
        RECT 84.925 52.455 85.095 52.955 ;
        RECT 84.440 51.715 85.055 52.285 ;
        RECT 85.345 52.225 85.610 52.785 ;
        RECT 85.780 52.055 85.950 52.955 ;
        RECT 86.120 52.225 86.475 52.785 ;
        RECT 86.705 52.445 87.060 52.815 ;
        RECT 87.340 52.785 87.510 52.995 ;
        RECT 87.340 52.455 87.595 52.785 ;
        RECT 87.340 52.265 87.510 52.455 ;
        RECT 87.765 52.290 87.935 53.020 ;
        RECT 88.110 52.945 88.370 54.095 ;
        RECT 88.545 53.005 89.755 54.095 ;
        RECT 88.545 52.465 89.065 53.005 ;
        RECT 86.795 52.095 87.510 52.265 ;
        RECT 85.225 51.545 85.440 52.055 ;
        RECT 85.670 51.725 85.950 52.055 ;
        RECT 86.130 51.545 86.370 52.055 ;
        RECT 86.795 51.715 86.965 52.095 ;
        RECT 87.180 51.545 87.510 51.925 ;
        RECT 87.680 51.715 87.935 52.290 ;
        RECT 88.110 51.545 88.370 52.385 ;
        RECT 89.235 52.295 89.755 52.835 ;
        RECT 88.545 51.545 89.755 52.295 ;
        RECT 12.100 51.375 89.840 51.545 ;
        RECT 12.185 50.625 13.395 51.375 ;
        RECT 13.615 50.720 13.945 51.155 ;
        RECT 14.115 50.765 14.285 51.375 ;
        RECT 13.565 50.635 13.945 50.720 ;
        RECT 14.455 50.635 14.785 51.160 ;
        RECT 15.045 50.845 15.255 51.375 ;
        RECT 15.530 50.925 16.315 51.095 ;
        RECT 16.485 50.925 16.890 51.095 ;
        RECT 12.185 50.085 12.705 50.625 ;
        RECT 13.565 50.595 13.790 50.635 ;
        RECT 12.875 49.915 13.395 50.455 ;
        RECT 12.185 48.825 13.395 49.915 ;
        RECT 13.565 50.015 13.735 50.595 ;
        RECT 14.455 50.465 14.655 50.635 ;
        RECT 15.530 50.465 15.700 50.925 ;
        RECT 13.905 50.135 14.655 50.465 ;
        RECT 14.825 50.135 15.700 50.465 ;
        RECT 13.565 49.965 13.780 50.015 ;
        RECT 13.565 49.885 13.955 49.965 ;
        RECT 13.625 49.040 13.955 49.885 ;
        RECT 14.465 49.930 14.655 50.135 ;
        RECT 14.125 48.825 14.295 49.835 ;
        RECT 14.465 49.555 15.360 49.930 ;
        RECT 14.465 48.995 14.805 49.555 ;
        RECT 15.035 48.825 15.350 49.325 ;
        RECT 15.530 49.295 15.700 50.135 ;
        RECT 15.870 50.425 16.335 50.755 ;
        RECT 16.720 50.695 16.890 50.925 ;
        RECT 17.070 50.875 17.440 51.375 ;
        RECT 17.760 50.925 18.435 51.095 ;
        RECT 18.630 50.925 18.965 51.095 ;
        RECT 15.870 49.465 16.190 50.425 ;
        RECT 16.720 50.395 17.550 50.695 ;
        RECT 16.360 49.495 16.550 50.215 ;
        RECT 16.720 49.325 16.890 50.395 ;
        RECT 17.350 50.365 17.550 50.395 ;
        RECT 17.060 50.145 17.230 50.215 ;
        RECT 17.760 50.145 17.930 50.925 ;
        RECT 18.795 50.785 18.965 50.925 ;
        RECT 19.135 50.915 19.385 51.375 ;
        RECT 17.060 49.975 17.930 50.145 ;
        RECT 18.100 50.505 18.625 50.725 ;
        RECT 18.795 50.655 19.020 50.785 ;
        RECT 17.060 49.885 17.570 49.975 ;
        RECT 15.530 49.125 16.415 49.295 ;
        RECT 16.640 48.995 16.890 49.325 ;
        RECT 17.060 48.825 17.230 49.625 ;
        RECT 17.400 49.270 17.570 49.885 ;
        RECT 18.100 49.805 18.270 50.505 ;
        RECT 17.740 49.440 18.270 49.805 ;
        RECT 18.440 49.740 18.680 50.335 ;
        RECT 18.850 49.550 19.020 50.655 ;
        RECT 19.190 49.795 19.470 50.745 ;
        RECT 18.715 49.420 19.020 49.550 ;
        RECT 17.400 49.100 18.505 49.270 ;
        RECT 18.715 48.995 18.965 49.420 ;
        RECT 19.135 48.825 19.400 49.285 ;
        RECT 19.640 48.995 19.825 51.115 ;
        RECT 19.995 50.995 20.325 51.375 ;
        RECT 20.495 50.825 20.665 51.115 ;
        RECT 20.925 50.995 21.815 51.165 ;
        RECT 20.000 50.655 20.665 50.825 ;
        RECT 20.000 49.665 20.230 50.655 ;
        RECT 20.400 49.835 20.750 50.485 ;
        RECT 20.925 50.440 21.475 50.825 ;
        RECT 21.645 50.270 21.815 50.995 ;
        RECT 20.925 50.200 21.815 50.270 ;
        RECT 21.985 50.670 22.205 51.155 ;
        RECT 22.375 50.835 22.625 51.375 ;
        RECT 22.795 50.725 23.055 51.205 ;
        RECT 21.985 50.245 22.315 50.670 ;
        RECT 20.925 50.175 21.820 50.200 ;
        RECT 20.925 50.160 21.830 50.175 ;
        RECT 20.925 50.145 21.835 50.160 ;
        RECT 20.925 50.140 21.845 50.145 ;
        RECT 20.925 50.130 21.850 50.140 ;
        RECT 20.925 50.120 21.855 50.130 ;
        RECT 20.925 50.115 21.865 50.120 ;
        RECT 20.925 50.105 21.875 50.115 ;
        RECT 20.925 50.100 21.885 50.105 ;
        RECT 20.000 49.495 20.665 49.665 ;
        RECT 20.925 49.650 21.185 50.100 ;
        RECT 21.550 50.095 21.885 50.100 ;
        RECT 21.550 50.090 21.900 50.095 ;
        RECT 21.550 50.080 21.915 50.090 ;
        RECT 21.550 50.075 21.940 50.080 ;
        RECT 22.485 50.075 22.715 50.470 ;
        RECT 21.550 50.070 22.715 50.075 ;
        RECT 21.580 50.035 22.715 50.070 ;
        RECT 21.615 50.010 22.715 50.035 ;
        RECT 21.645 49.980 22.715 50.010 ;
        RECT 21.665 49.950 22.715 49.980 ;
        RECT 21.685 49.920 22.715 49.950 ;
        RECT 21.755 49.910 22.715 49.920 ;
        RECT 21.780 49.900 22.715 49.910 ;
        RECT 21.800 49.885 22.715 49.900 ;
        RECT 21.820 49.870 22.715 49.885 ;
        RECT 21.825 49.860 22.610 49.870 ;
        RECT 21.840 49.825 22.610 49.860 ;
        RECT 19.995 48.825 20.325 49.325 ;
        RECT 20.495 48.995 20.665 49.495 ;
        RECT 21.355 49.505 21.685 49.750 ;
        RECT 21.855 49.575 22.610 49.825 ;
        RECT 22.885 49.695 23.055 50.725 ;
        RECT 23.245 50.565 23.485 51.375 ;
        RECT 23.655 50.565 23.985 51.205 ;
        RECT 24.155 50.565 24.425 51.375 ;
        RECT 24.605 50.605 28.115 51.375 ;
        RECT 28.320 50.635 28.935 51.205 ;
        RECT 29.105 50.865 29.320 51.375 ;
        RECT 29.550 50.865 29.830 51.195 ;
        RECT 30.010 50.865 30.250 51.375 ;
        RECT 30.585 50.995 31.475 51.165 ;
        RECT 23.225 50.135 23.575 50.385 ;
        RECT 23.745 49.965 23.915 50.565 ;
        RECT 24.085 50.135 24.435 50.385 ;
        RECT 24.605 50.085 26.255 50.605 ;
        RECT 21.355 49.480 21.540 49.505 ;
        RECT 20.925 49.380 21.540 49.480 ;
        RECT 20.925 48.825 21.530 49.380 ;
        RECT 21.705 48.995 22.185 49.335 ;
        RECT 22.355 48.825 22.610 49.370 ;
        RECT 22.780 48.995 23.055 49.695 ;
        RECT 23.235 49.795 23.915 49.965 ;
        RECT 23.235 49.010 23.565 49.795 ;
        RECT 24.095 48.825 24.425 49.965 ;
        RECT 26.425 49.915 28.115 50.435 ;
        RECT 24.605 48.825 28.115 49.915 ;
        RECT 28.320 49.615 28.635 50.635 ;
        RECT 28.805 49.965 28.975 50.465 ;
        RECT 29.225 50.135 29.490 50.695 ;
        RECT 29.660 49.965 29.830 50.865 ;
        RECT 30.000 50.135 30.355 50.695 ;
        RECT 30.585 50.440 31.135 50.825 ;
        RECT 31.305 50.270 31.475 50.995 ;
        RECT 30.585 50.200 31.475 50.270 ;
        RECT 31.645 50.670 31.865 51.155 ;
        RECT 32.035 50.835 32.285 51.375 ;
        RECT 32.455 50.725 32.715 51.205 ;
        RECT 31.645 50.245 31.975 50.670 ;
        RECT 30.585 50.175 31.480 50.200 ;
        RECT 30.585 50.160 31.490 50.175 ;
        RECT 30.585 50.145 31.495 50.160 ;
        RECT 30.585 50.140 31.505 50.145 ;
        RECT 30.585 50.130 31.510 50.140 ;
        RECT 30.585 50.120 31.515 50.130 ;
        RECT 30.585 50.115 31.525 50.120 ;
        RECT 30.585 50.105 31.535 50.115 ;
        RECT 30.585 50.100 31.545 50.105 ;
        RECT 28.805 49.795 30.230 49.965 ;
        RECT 28.320 48.995 28.855 49.615 ;
        RECT 29.025 48.825 29.355 49.625 ;
        RECT 29.840 49.620 30.230 49.795 ;
        RECT 30.585 49.650 30.845 50.100 ;
        RECT 31.210 50.095 31.545 50.100 ;
        RECT 31.210 50.090 31.560 50.095 ;
        RECT 31.210 50.080 31.575 50.090 ;
        RECT 31.210 50.075 31.600 50.080 ;
        RECT 32.145 50.075 32.375 50.470 ;
        RECT 31.210 50.070 32.375 50.075 ;
        RECT 31.240 50.035 32.375 50.070 ;
        RECT 31.275 50.010 32.375 50.035 ;
        RECT 31.305 49.980 32.375 50.010 ;
        RECT 31.325 49.950 32.375 49.980 ;
        RECT 31.345 49.920 32.375 49.950 ;
        RECT 31.415 49.910 32.375 49.920 ;
        RECT 31.440 49.900 32.375 49.910 ;
        RECT 31.460 49.885 32.375 49.900 ;
        RECT 31.480 49.870 32.375 49.885 ;
        RECT 31.485 49.860 32.270 49.870 ;
        RECT 31.500 49.825 32.270 49.860 ;
        RECT 31.015 49.505 31.345 49.750 ;
        RECT 31.515 49.575 32.270 49.825 ;
        RECT 32.545 49.695 32.715 50.725 ;
        RECT 31.015 49.480 31.200 49.505 ;
        RECT 30.585 49.380 31.200 49.480 ;
        RECT 30.585 48.825 31.190 49.380 ;
        RECT 31.365 48.995 31.845 49.335 ;
        RECT 32.015 48.825 32.270 49.370 ;
        RECT 32.440 48.995 32.715 49.695 ;
        RECT 32.885 50.635 33.325 51.195 ;
        RECT 33.495 50.635 33.945 51.375 ;
        RECT 34.115 50.805 34.285 51.205 ;
        RECT 34.455 50.975 34.875 51.375 ;
        RECT 35.045 50.805 35.275 51.205 ;
        RECT 34.115 50.635 35.275 50.805 ;
        RECT 35.445 50.635 35.935 51.205 ;
        RECT 32.885 49.625 33.195 50.635 ;
        RECT 33.365 50.015 33.535 50.465 ;
        RECT 33.705 50.185 34.095 50.465 ;
        RECT 34.280 50.135 34.525 50.465 ;
        RECT 33.365 49.845 34.155 50.015 ;
        RECT 32.885 48.995 33.325 49.625 ;
        RECT 33.500 48.825 33.815 49.675 ;
        RECT 33.985 49.165 34.155 49.845 ;
        RECT 34.325 49.335 34.525 50.135 ;
        RECT 34.725 49.335 34.975 50.465 ;
        RECT 35.190 50.135 35.595 50.465 ;
        RECT 35.765 49.965 35.935 50.635 ;
        RECT 36.105 50.605 37.775 51.375 ;
        RECT 37.945 50.650 38.235 51.375 ;
        RECT 38.405 50.915 38.965 51.205 ;
        RECT 39.135 50.915 39.385 51.375 ;
        RECT 36.105 50.085 36.855 50.605 ;
        RECT 35.165 49.795 35.935 49.965 ;
        RECT 37.025 49.915 37.775 50.435 ;
        RECT 35.165 49.165 35.415 49.795 ;
        RECT 33.985 48.995 35.415 49.165 ;
        RECT 35.595 48.825 35.925 49.625 ;
        RECT 36.105 48.825 37.775 49.915 ;
        RECT 37.945 48.825 38.235 49.990 ;
        RECT 38.405 49.545 38.655 50.915 ;
        RECT 40.005 50.745 40.335 51.105 ;
        RECT 38.945 50.555 40.335 50.745 ;
        RECT 41.255 50.825 41.425 51.115 ;
        RECT 41.595 50.995 41.925 51.375 ;
        RECT 41.255 50.655 41.920 50.825 ;
        RECT 38.945 50.465 39.115 50.555 ;
        RECT 38.825 50.135 39.115 50.465 ;
        RECT 39.285 50.135 39.625 50.385 ;
        RECT 39.845 50.135 40.520 50.385 ;
        RECT 38.945 49.885 39.115 50.135 ;
        RECT 38.945 49.715 39.885 49.885 ;
        RECT 40.255 49.775 40.520 50.135 ;
        RECT 41.170 49.835 41.520 50.485 ;
        RECT 38.405 48.995 38.865 49.545 ;
        RECT 39.055 48.825 39.385 49.545 ;
        RECT 39.585 49.165 39.885 49.715 ;
        RECT 41.690 49.665 41.920 50.655 ;
        RECT 41.255 49.495 41.920 49.665 ;
        RECT 40.055 48.825 40.335 49.495 ;
        RECT 41.255 48.995 41.425 49.495 ;
        RECT 41.595 48.825 41.925 49.325 ;
        RECT 42.095 48.995 42.280 51.115 ;
        RECT 42.535 50.915 42.785 51.375 ;
        RECT 42.955 50.925 43.290 51.095 ;
        RECT 43.485 50.925 44.160 51.095 ;
        RECT 42.955 50.785 43.125 50.925 ;
        RECT 42.450 49.795 42.730 50.745 ;
        RECT 42.900 50.655 43.125 50.785 ;
        RECT 42.900 49.550 43.070 50.655 ;
        RECT 43.295 50.505 43.820 50.725 ;
        RECT 43.240 49.740 43.480 50.335 ;
        RECT 43.650 49.805 43.820 50.505 ;
        RECT 43.990 50.145 44.160 50.925 ;
        RECT 44.480 50.875 44.850 51.375 ;
        RECT 45.030 50.925 45.435 51.095 ;
        RECT 45.605 50.925 46.390 51.095 ;
        RECT 45.030 50.695 45.200 50.925 ;
        RECT 44.370 50.395 45.200 50.695 ;
        RECT 45.585 50.425 46.050 50.755 ;
        RECT 44.370 50.365 44.570 50.395 ;
        RECT 44.690 50.145 44.860 50.215 ;
        RECT 43.990 49.975 44.860 50.145 ;
        RECT 44.350 49.885 44.860 49.975 ;
        RECT 42.900 49.420 43.205 49.550 ;
        RECT 43.650 49.440 44.180 49.805 ;
        RECT 42.520 48.825 42.785 49.285 ;
        RECT 42.955 48.995 43.205 49.420 ;
        RECT 44.350 49.270 44.520 49.885 ;
        RECT 43.415 49.100 44.520 49.270 ;
        RECT 44.690 48.825 44.860 49.625 ;
        RECT 45.030 49.325 45.200 50.395 ;
        RECT 45.370 49.495 45.560 50.215 ;
        RECT 45.730 49.465 46.050 50.425 ;
        RECT 46.220 50.465 46.390 50.925 ;
        RECT 46.665 50.845 46.875 51.375 ;
        RECT 47.135 50.635 47.465 51.160 ;
        RECT 47.635 50.765 47.805 51.375 ;
        RECT 47.975 50.720 48.305 51.155 ;
        RECT 48.615 50.825 48.785 51.115 ;
        RECT 48.955 50.995 49.285 51.375 ;
        RECT 47.975 50.635 48.355 50.720 ;
        RECT 48.615 50.655 49.280 50.825 ;
        RECT 47.265 50.465 47.465 50.635 ;
        RECT 48.130 50.595 48.355 50.635 ;
        RECT 46.220 50.135 47.095 50.465 ;
        RECT 47.265 50.135 48.015 50.465 ;
        RECT 45.030 48.995 45.280 49.325 ;
        RECT 46.220 49.295 46.390 50.135 ;
        RECT 47.265 49.930 47.455 50.135 ;
        RECT 48.185 50.015 48.355 50.595 ;
        RECT 48.140 49.965 48.355 50.015 ;
        RECT 46.560 49.555 47.455 49.930 ;
        RECT 47.965 49.885 48.355 49.965 ;
        RECT 45.505 49.125 46.390 49.295 ;
        RECT 46.570 48.825 46.885 49.325 ;
        RECT 47.115 48.995 47.455 49.555 ;
        RECT 47.625 48.825 47.795 49.835 ;
        RECT 47.965 49.040 48.295 49.885 ;
        RECT 48.530 49.835 48.880 50.485 ;
        RECT 49.050 49.665 49.280 50.655 ;
        RECT 48.615 49.495 49.280 49.665 ;
        RECT 48.615 48.995 48.785 49.495 ;
        RECT 48.955 48.825 49.285 49.325 ;
        RECT 49.455 48.995 49.640 51.115 ;
        RECT 49.895 50.915 50.145 51.375 ;
        RECT 50.315 50.925 50.650 51.095 ;
        RECT 50.845 50.925 51.520 51.095 ;
        RECT 50.315 50.785 50.485 50.925 ;
        RECT 49.810 49.795 50.090 50.745 ;
        RECT 50.260 50.655 50.485 50.785 ;
        RECT 50.260 49.550 50.430 50.655 ;
        RECT 50.655 50.505 51.180 50.725 ;
        RECT 50.600 49.740 50.840 50.335 ;
        RECT 51.010 49.805 51.180 50.505 ;
        RECT 51.350 50.145 51.520 50.925 ;
        RECT 51.840 50.875 52.210 51.375 ;
        RECT 52.390 50.925 52.795 51.095 ;
        RECT 52.965 50.925 53.750 51.095 ;
        RECT 52.390 50.695 52.560 50.925 ;
        RECT 51.730 50.395 52.560 50.695 ;
        RECT 52.945 50.425 53.410 50.755 ;
        RECT 51.730 50.365 51.930 50.395 ;
        RECT 52.050 50.145 52.220 50.215 ;
        RECT 51.350 49.975 52.220 50.145 ;
        RECT 51.710 49.885 52.220 49.975 ;
        RECT 50.260 49.420 50.565 49.550 ;
        RECT 51.010 49.440 51.540 49.805 ;
        RECT 49.880 48.825 50.145 49.285 ;
        RECT 50.315 48.995 50.565 49.420 ;
        RECT 51.710 49.270 51.880 49.885 ;
        RECT 50.775 49.100 51.880 49.270 ;
        RECT 52.050 48.825 52.220 49.625 ;
        RECT 52.390 49.325 52.560 50.395 ;
        RECT 52.730 49.495 52.920 50.215 ;
        RECT 53.090 49.465 53.410 50.425 ;
        RECT 53.580 50.465 53.750 50.925 ;
        RECT 54.025 50.845 54.235 51.375 ;
        RECT 54.495 50.635 54.825 51.160 ;
        RECT 54.995 50.765 55.165 51.375 ;
        RECT 55.335 50.720 55.665 51.155 ;
        RECT 55.895 50.885 56.225 51.375 ;
        RECT 56.395 50.780 57.015 51.205 ;
        RECT 55.335 50.635 55.715 50.720 ;
        RECT 54.625 50.465 54.825 50.635 ;
        RECT 55.490 50.595 55.715 50.635 ;
        RECT 53.580 50.135 54.455 50.465 ;
        RECT 54.625 50.135 55.375 50.465 ;
        RECT 52.390 48.995 52.640 49.325 ;
        RECT 53.580 49.295 53.750 50.135 ;
        RECT 54.625 49.930 54.815 50.135 ;
        RECT 55.545 50.015 55.715 50.595 ;
        RECT 55.885 50.135 56.225 50.715 ;
        RECT 56.395 50.445 56.755 50.780 ;
        RECT 57.475 50.685 57.805 51.375 ;
        RECT 58.650 50.635 58.905 51.205 ;
        RECT 59.075 50.975 59.405 51.375 ;
        RECT 59.830 50.840 60.360 51.205 ;
        RECT 60.550 51.035 60.825 51.205 ;
        RECT 60.545 50.865 60.825 51.035 ;
        RECT 59.830 50.805 60.005 50.840 ;
        RECT 59.075 50.635 60.005 50.805 ;
        RECT 56.395 50.165 57.815 50.445 ;
        RECT 55.500 49.965 55.715 50.015 ;
        RECT 53.920 49.555 54.815 49.930 ;
        RECT 55.325 49.885 55.715 49.965 ;
        RECT 52.865 49.125 53.750 49.295 ;
        RECT 53.930 48.825 54.245 49.325 ;
        RECT 54.475 48.995 54.815 49.555 ;
        RECT 54.985 48.825 55.155 49.835 ;
        RECT 55.325 49.040 55.655 49.885 ;
        RECT 55.895 48.825 56.225 49.965 ;
        RECT 56.395 48.995 56.755 50.165 ;
        RECT 56.955 48.825 57.285 49.995 ;
        RECT 57.485 48.995 57.815 50.165 ;
        RECT 58.015 48.825 58.345 49.995 ;
        RECT 58.650 49.965 58.820 50.635 ;
        RECT 59.075 50.465 59.245 50.635 ;
        RECT 58.990 50.135 59.245 50.465 ;
        RECT 59.470 50.135 59.665 50.465 ;
        RECT 58.650 48.995 58.985 49.965 ;
        RECT 59.155 48.825 59.325 49.965 ;
        RECT 59.495 49.165 59.665 50.135 ;
        RECT 59.835 49.505 60.005 50.635 ;
        RECT 60.175 49.845 60.345 50.645 ;
        RECT 60.550 50.045 60.825 50.865 ;
        RECT 60.995 49.845 61.185 51.205 ;
        RECT 61.365 50.840 61.875 51.375 ;
        RECT 62.095 50.565 62.340 51.170 ;
        RECT 63.705 50.650 63.995 51.375 ;
        RECT 65.090 50.635 65.345 51.205 ;
        RECT 65.515 50.975 65.845 51.375 ;
        RECT 66.270 50.840 66.800 51.205 ;
        RECT 66.270 50.805 66.445 50.840 ;
        RECT 65.515 50.635 66.445 50.805 ;
        RECT 61.385 50.395 62.615 50.565 ;
        RECT 60.175 49.675 61.185 49.845 ;
        RECT 61.355 49.830 62.105 50.020 ;
        RECT 59.835 49.335 60.960 49.505 ;
        RECT 61.355 49.165 61.525 49.830 ;
        RECT 62.275 49.585 62.615 50.395 ;
        RECT 59.495 48.995 61.525 49.165 ;
        RECT 61.695 48.825 61.865 49.585 ;
        RECT 62.100 49.175 62.615 49.585 ;
        RECT 63.705 48.825 63.995 49.990 ;
        RECT 65.090 49.965 65.260 50.635 ;
        RECT 65.515 50.465 65.685 50.635 ;
        RECT 65.430 50.135 65.685 50.465 ;
        RECT 65.910 50.135 66.105 50.465 ;
        RECT 65.090 48.995 65.425 49.965 ;
        RECT 65.595 48.825 65.765 49.965 ;
        RECT 65.935 49.165 66.105 50.135 ;
        RECT 66.275 49.505 66.445 50.635 ;
        RECT 66.615 49.845 66.785 50.645 ;
        RECT 66.990 50.355 67.265 51.205 ;
        RECT 66.985 50.185 67.265 50.355 ;
        RECT 66.990 50.045 67.265 50.185 ;
        RECT 67.435 49.845 67.625 51.205 ;
        RECT 67.805 50.840 68.315 51.375 ;
        RECT 68.535 50.565 68.780 51.170 ;
        RECT 69.230 50.635 69.485 51.205 ;
        RECT 69.655 50.975 69.985 51.375 ;
        RECT 70.410 50.840 70.940 51.205 ;
        RECT 70.410 50.805 70.585 50.840 ;
        RECT 69.655 50.635 70.585 50.805 ;
        RECT 67.825 50.395 69.055 50.565 ;
        RECT 66.615 49.675 67.625 49.845 ;
        RECT 67.795 49.830 68.545 50.020 ;
        RECT 66.275 49.335 67.400 49.505 ;
        RECT 67.795 49.165 67.965 49.830 ;
        RECT 68.715 49.585 69.055 50.395 ;
        RECT 65.935 48.995 67.965 49.165 ;
        RECT 68.135 48.825 68.305 49.585 ;
        RECT 68.540 49.175 69.055 49.585 ;
        RECT 69.230 49.965 69.400 50.635 ;
        RECT 69.655 50.465 69.825 50.635 ;
        RECT 69.570 50.135 69.825 50.465 ;
        RECT 70.050 50.135 70.245 50.465 ;
        RECT 69.230 48.995 69.565 49.965 ;
        RECT 69.735 48.825 69.905 49.965 ;
        RECT 70.075 49.165 70.245 50.135 ;
        RECT 70.415 49.505 70.585 50.635 ;
        RECT 70.755 49.845 70.925 50.645 ;
        RECT 71.130 50.355 71.405 51.205 ;
        RECT 71.125 50.185 71.405 50.355 ;
        RECT 71.130 50.045 71.405 50.185 ;
        RECT 71.575 49.845 71.765 51.205 ;
        RECT 71.945 50.840 72.455 51.375 ;
        RECT 72.675 50.565 72.920 51.170 ;
        RECT 73.365 50.575 73.705 51.205 ;
        RECT 73.875 50.575 74.125 51.375 ;
        RECT 74.315 50.725 74.645 51.205 ;
        RECT 74.815 50.915 75.040 51.375 ;
        RECT 75.210 50.725 75.540 51.205 ;
        RECT 71.965 50.395 73.195 50.565 ;
        RECT 70.755 49.675 71.765 49.845 ;
        RECT 71.935 49.830 72.685 50.020 ;
        RECT 70.415 49.335 71.540 49.505 ;
        RECT 71.935 49.165 72.105 49.830 ;
        RECT 72.855 49.585 73.195 50.395 ;
        RECT 70.075 48.995 72.105 49.165 ;
        RECT 72.275 48.825 72.445 49.585 ;
        RECT 72.680 49.175 73.195 49.585 ;
        RECT 73.365 49.965 73.540 50.575 ;
        RECT 74.315 50.555 75.540 50.725 ;
        RECT 76.170 50.595 76.670 51.205 ;
        RECT 77.710 50.595 78.210 51.205 ;
        RECT 73.710 50.215 74.405 50.385 ;
        RECT 74.235 49.965 74.405 50.215 ;
        RECT 74.580 50.185 75.000 50.385 ;
        RECT 75.170 50.185 75.500 50.385 ;
        RECT 75.670 50.185 76.000 50.385 ;
        RECT 76.170 49.965 76.340 50.595 ;
        RECT 76.525 50.135 76.875 50.385 ;
        RECT 77.505 50.135 77.855 50.385 ;
        RECT 78.040 49.965 78.210 50.595 ;
        RECT 78.840 50.725 79.170 51.205 ;
        RECT 79.340 50.915 79.565 51.375 ;
        RECT 79.735 50.725 80.065 51.205 ;
        RECT 78.840 50.555 80.065 50.725 ;
        RECT 80.255 50.575 80.505 51.375 ;
        RECT 80.675 50.575 81.015 51.205 ;
        RECT 81.275 50.825 81.445 51.115 ;
        RECT 81.615 50.995 81.945 51.375 ;
        RECT 81.275 50.655 81.940 50.825 ;
        RECT 78.380 50.185 78.710 50.385 ;
        RECT 78.880 50.185 79.210 50.385 ;
        RECT 79.380 50.185 79.800 50.385 ;
        RECT 79.975 50.215 80.670 50.385 ;
        RECT 79.975 49.965 80.145 50.215 ;
        RECT 80.840 49.965 81.015 50.575 ;
        RECT 73.365 48.995 73.705 49.965 ;
        RECT 73.875 48.825 74.045 49.965 ;
        RECT 74.235 49.795 76.670 49.965 ;
        RECT 74.315 48.825 74.565 49.625 ;
        RECT 75.210 48.995 75.540 49.795 ;
        RECT 75.840 48.825 76.170 49.625 ;
        RECT 76.340 48.995 76.670 49.795 ;
        RECT 77.710 49.795 80.145 49.965 ;
        RECT 77.710 48.995 78.040 49.795 ;
        RECT 78.210 48.825 78.540 49.625 ;
        RECT 78.840 48.995 79.170 49.795 ;
        RECT 79.815 48.825 80.065 49.625 ;
        RECT 80.335 48.825 80.505 49.965 ;
        RECT 80.675 48.995 81.015 49.965 ;
        RECT 81.190 49.835 81.540 50.485 ;
        RECT 81.710 49.665 81.940 50.655 ;
        RECT 81.275 49.495 81.940 49.665 ;
        RECT 81.275 48.995 81.445 49.495 ;
        RECT 81.615 48.825 81.945 49.325 ;
        RECT 82.115 48.995 82.300 51.115 ;
        RECT 82.555 50.915 82.805 51.375 ;
        RECT 82.975 50.925 83.310 51.095 ;
        RECT 83.505 50.925 84.180 51.095 ;
        RECT 82.975 50.785 83.145 50.925 ;
        RECT 82.470 49.795 82.750 50.745 ;
        RECT 82.920 50.655 83.145 50.785 ;
        RECT 82.920 49.550 83.090 50.655 ;
        RECT 83.315 50.505 83.840 50.725 ;
        RECT 83.260 49.740 83.500 50.335 ;
        RECT 83.670 49.805 83.840 50.505 ;
        RECT 84.010 50.145 84.180 50.925 ;
        RECT 84.500 50.875 84.870 51.375 ;
        RECT 85.050 50.925 85.455 51.095 ;
        RECT 85.625 50.925 86.410 51.095 ;
        RECT 85.050 50.695 85.220 50.925 ;
        RECT 84.390 50.395 85.220 50.695 ;
        RECT 85.605 50.425 86.070 50.755 ;
        RECT 84.390 50.365 84.590 50.395 ;
        RECT 84.710 50.145 84.880 50.215 ;
        RECT 84.010 49.975 84.880 50.145 ;
        RECT 84.370 49.885 84.880 49.975 ;
        RECT 82.920 49.420 83.225 49.550 ;
        RECT 83.670 49.440 84.200 49.805 ;
        RECT 82.540 48.825 82.805 49.285 ;
        RECT 82.975 48.995 83.225 49.420 ;
        RECT 84.370 49.270 84.540 49.885 ;
        RECT 83.435 49.100 84.540 49.270 ;
        RECT 84.710 48.825 84.880 49.625 ;
        RECT 85.050 49.325 85.220 50.395 ;
        RECT 85.390 49.495 85.580 50.215 ;
        RECT 85.750 49.465 86.070 50.425 ;
        RECT 86.240 50.465 86.410 50.925 ;
        RECT 86.685 50.845 86.895 51.375 ;
        RECT 87.155 50.635 87.485 51.160 ;
        RECT 87.655 50.765 87.825 51.375 ;
        RECT 87.995 50.720 88.325 51.155 ;
        RECT 87.995 50.635 88.375 50.720 ;
        RECT 87.285 50.465 87.485 50.635 ;
        RECT 88.150 50.595 88.375 50.635 ;
        RECT 88.545 50.625 89.755 51.375 ;
        RECT 86.240 50.135 87.115 50.465 ;
        RECT 87.285 50.135 88.035 50.465 ;
        RECT 85.050 48.995 85.300 49.325 ;
        RECT 86.240 49.295 86.410 50.135 ;
        RECT 87.285 49.930 87.475 50.135 ;
        RECT 88.205 50.015 88.375 50.595 ;
        RECT 88.160 49.965 88.375 50.015 ;
        RECT 86.580 49.555 87.475 49.930 ;
        RECT 87.985 49.885 88.375 49.965 ;
        RECT 88.545 49.915 89.065 50.455 ;
        RECT 89.235 50.085 89.755 50.625 ;
        RECT 85.525 49.125 86.410 49.295 ;
        RECT 86.590 48.825 86.905 49.325 ;
        RECT 87.135 48.995 87.475 49.555 ;
        RECT 87.645 48.825 87.815 49.835 ;
        RECT 87.985 49.040 88.315 49.885 ;
        RECT 88.545 48.825 89.755 49.915 ;
        RECT 12.100 48.655 89.840 48.825 ;
        RECT 12.185 47.565 13.395 48.655 ;
        RECT 14.575 47.985 14.745 48.485 ;
        RECT 14.915 48.155 15.245 48.655 ;
        RECT 14.575 47.815 15.240 47.985 ;
        RECT 12.185 46.855 12.705 47.395 ;
        RECT 12.875 47.025 13.395 47.565 ;
        RECT 14.490 46.995 14.840 47.645 ;
        RECT 12.185 46.105 13.395 46.855 ;
        RECT 15.010 46.825 15.240 47.815 ;
        RECT 14.575 46.655 15.240 46.825 ;
        RECT 14.575 46.365 14.745 46.655 ;
        RECT 14.915 46.105 15.245 46.485 ;
        RECT 15.415 46.365 15.600 48.485 ;
        RECT 15.840 48.195 16.105 48.655 ;
        RECT 16.275 48.060 16.525 48.485 ;
        RECT 16.735 48.210 17.840 48.380 ;
        RECT 16.220 47.930 16.525 48.060 ;
        RECT 15.770 46.735 16.050 47.685 ;
        RECT 16.220 46.825 16.390 47.930 ;
        RECT 16.560 47.145 16.800 47.740 ;
        RECT 16.970 47.675 17.500 48.040 ;
        RECT 16.970 46.975 17.140 47.675 ;
        RECT 17.670 47.595 17.840 48.210 ;
        RECT 18.010 47.855 18.180 48.655 ;
        RECT 18.350 48.155 18.600 48.485 ;
        RECT 18.825 48.185 19.710 48.355 ;
        RECT 17.670 47.505 18.180 47.595 ;
        RECT 16.220 46.695 16.445 46.825 ;
        RECT 16.615 46.755 17.140 46.975 ;
        RECT 17.310 47.335 18.180 47.505 ;
        RECT 15.855 46.105 16.105 46.565 ;
        RECT 16.275 46.555 16.445 46.695 ;
        RECT 17.310 46.555 17.480 47.335 ;
        RECT 18.010 47.265 18.180 47.335 ;
        RECT 17.690 47.085 17.890 47.115 ;
        RECT 18.350 47.085 18.520 48.155 ;
        RECT 18.690 47.265 18.880 47.985 ;
        RECT 17.690 46.785 18.520 47.085 ;
        RECT 19.050 47.055 19.370 48.015 ;
        RECT 16.275 46.385 16.610 46.555 ;
        RECT 16.805 46.385 17.480 46.555 ;
        RECT 17.800 46.105 18.170 46.605 ;
        RECT 18.350 46.555 18.520 46.785 ;
        RECT 18.905 46.725 19.370 47.055 ;
        RECT 19.540 47.345 19.710 48.185 ;
        RECT 19.890 48.155 20.205 48.655 ;
        RECT 20.435 47.925 20.775 48.485 ;
        RECT 19.880 47.550 20.775 47.925 ;
        RECT 20.945 47.645 21.115 48.655 ;
        RECT 20.585 47.345 20.775 47.550 ;
        RECT 21.285 47.595 21.615 48.440 ;
        RECT 21.845 48.225 22.185 48.485 ;
        RECT 21.285 47.515 21.675 47.595 ;
        RECT 21.460 47.465 21.675 47.515 ;
        RECT 19.540 47.015 20.415 47.345 ;
        RECT 20.585 47.015 21.335 47.345 ;
        RECT 19.540 46.555 19.710 47.015 ;
        RECT 20.585 46.845 20.785 47.015 ;
        RECT 21.505 46.885 21.675 47.465 ;
        RECT 21.450 46.845 21.675 46.885 ;
        RECT 18.350 46.385 18.755 46.555 ;
        RECT 18.925 46.385 19.710 46.555 ;
        RECT 19.985 46.105 20.195 46.635 ;
        RECT 20.455 46.320 20.785 46.845 ;
        RECT 21.295 46.760 21.675 46.845 ;
        RECT 21.845 46.825 22.105 48.225 ;
        RECT 22.355 47.855 22.685 48.655 ;
        RECT 23.150 47.685 23.400 48.485 ;
        RECT 23.585 47.935 23.915 48.655 ;
        RECT 24.135 47.685 24.385 48.485 ;
        RECT 24.555 48.275 24.890 48.655 ;
        RECT 22.295 47.515 24.485 47.685 ;
        RECT 22.295 47.345 22.610 47.515 ;
        RECT 22.280 47.095 22.610 47.345 ;
        RECT 20.955 46.105 21.125 46.715 ;
        RECT 21.295 46.325 21.625 46.760 ;
        RECT 21.845 46.315 22.185 46.825 ;
        RECT 22.355 46.105 22.625 46.905 ;
        RECT 22.805 46.375 23.085 47.345 ;
        RECT 23.265 46.375 23.565 47.345 ;
        RECT 23.745 46.380 24.095 47.345 ;
        RECT 24.315 46.605 24.485 47.515 ;
        RECT 24.655 46.785 24.895 48.095 ;
        RECT 25.065 47.490 25.355 48.655 ;
        RECT 25.535 48.045 25.865 48.475 ;
        RECT 26.045 48.215 26.240 48.655 ;
        RECT 26.410 48.045 26.740 48.475 ;
        RECT 25.535 47.875 26.740 48.045 ;
        RECT 25.535 47.545 26.430 47.875 ;
        RECT 26.910 47.705 27.185 48.475 ;
        RECT 26.600 47.515 27.185 47.705 ;
        RECT 27.375 47.685 27.705 48.470 ;
        RECT 27.375 47.515 28.055 47.685 ;
        RECT 28.235 47.515 28.565 48.655 ;
        RECT 28.745 47.565 32.255 48.655 ;
        RECT 25.540 47.015 25.835 47.345 ;
        RECT 26.015 47.015 26.430 47.345 ;
        RECT 24.315 46.275 24.810 46.605 ;
        RECT 25.065 46.105 25.355 46.830 ;
        RECT 25.535 46.105 25.835 46.835 ;
        RECT 26.015 46.395 26.245 47.015 ;
        RECT 26.600 46.845 26.775 47.515 ;
        RECT 26.445 46.665 26.775 46.845 ;
        RECT 26.945 46.695 27.185 47.345 ;
        RECT 27.365 47.095 27.715 47.345 ;
        RECT 27.885 46.915 28.055 47.515 ;
        RECT 28.225 47.095 28.575 47.345 ;
        RECT 26.445 46.285 26.670 46.665 ;
        RECT 26.840 46.105 27.170 46.495 ;
        RECT 27.385 46.105 27.625 46.915 ;
        RECT 27.795 46.275 28.125 46.915 ;
        RECT 28.295 46.105 28.565 46.915 ;
        RECT 28.745 46.875 30.395 47.395 ;
        RECT 30.565 47.045 32.255 47.565 ;
        RECT 32.425 47.785 32.700 48.485 ;
        RECT 32.910 48.110 33.125 48.655 ;
        RECT 33.295 48.145 33.770 48.485 ;
        RECT 33.940 48.150 34.555 48.655 ;
        RECT 33.940 47.975 34.135 48.150 ;
        RECT 28.745 46.105 32.255 46.875 ;
        RECT 32.425 46.755 32.595 47.785 ;
        RECT 32.870 47.615 33.585 47.910 ;
        RECT 33.805 47.785 34.135 47.975 ;
        RECT 34.305 47.615 34.555 47.980 ;
        RECT 32.765 47.445 34.555 47.615 ;
        RECT 32.765 47.015 32.995 47.445 ;
        RECT 32.425 46.275 32.685 46.755 ;
        RECT 33.165 46.745 33.575 47.265 ;
        RECT 32.855 46.105 33.185 46.565 ;
        RECT 33.375 46.325 33.575 46.745 ;
        RECT 33.745 46.590 34.000 47.445 ;
        RECT 34.795 47.265 34.965 48.485 ;
        RECT 35.215 48.145 35.475 48.655 ;
        RECT 35.645 48.225 35.985 48.485 ;
        RECT 34.170 47.015 34.965 47.265 ;
        RECT 35.135 47.095 35.475 47.975 ;
        RECT 34.715 46.925 34.965 47.015 ;
        RECT 33.745 46.325 34.535 46.590 ;
        RECT 34.715 46.505 35.045 46.925 ;
        RECT 35.215 46.105 35.475 46.925 ;
        RECT 35.645 46.825 35.905 48.225 ;
        RECT 36.155 47.855 36.485 48.655 ;
        RECT 36.950 47.685 37.200 48.485 ;
        RECT 37.385 47.935 37.715 48.655 ;
        RECT 37.935 47.685 38.185 48.485 ;
        RECT 38.355 48.275 38.690 48.655 ;
        RECT 36.095 47.515 38.285 47.685 ;
        RECT 36.095 47.345 36.410 47.515 ;
        RECT 36.080 47.095 36.410 47.345 ;
        RECT 35.645 46.315 35.985 46.825 ;
        RECT 36.155 46.105 36.425 46.905 ;
        RECT 36.605 46.375 36.885 47.345 ;
        RECT 37.065 46.375 37.365 47.345 ;
        RECT 37.545 46.380 37.895 47.345 ;
        RECT 38.115 46.605 38.285 47.515 ;
        RECT 38.455 46.785 38.695 48.095 ;
        RECT 38.875 47.595 39.205 48.445 ;
        RECT 38.875 46.830 39.065 47.595 ;
        RECT 39.375 47.515 39.625 48.655 ;
        RECT 39.815 48.015 40.065 48.435 ;
        RECT 40.295 48.185 40.625 48.655 ;
        RECT 40.855 48.015 41.105 48.435 ;
        RECT 39.815 47.845 41.105 48.015 ;
        RECT 41.285 48.015 41.615 48.445 ;
        RECT 41.285 47.845 41.740 48.015 ;
        RECT 39.805 47.345 40.020 47.675 ;
        RECT 39.235 47.015 39.545 47.345 ;
        RECT 39.715 47.015 40.020 47.345 ;
        RECT 40.195 47.015 40.480 47.675 ;
        RECT 40.675 47.015 40.940 47.675 ;
        RECT 41.155 47.015 41.400 47.675 ;
        RECT 39.375 46.845 39.545 47.015 ;
        RECT 41.570 46.845 41.740 47.845 ;
        RECT 38.115 46.275 38.610 46.605 ;
        RECT 38.875 46.320 39.205 46.830 ;
        RECT 39.375 46.675 41.740 46.845 ;
        RECT 42.120 47.865 42.655 48.485 ;
        RECT 42.120 46.845 42.435 47.865 ;
        RECT 42.825 47.855 43.155 48.655 ;
        RECT 43.640 47.685 44.030 47.860 ;
        RECT 42.605 47.515 44.030 47.685 ;
        RECT 44.385 47.565 45.595 48.655 ;
        RECT 42.605 47.015 42.775 47.515 ;
        RECT 39.375 46.105 39.705 46.505 ;
        RECT 40.755 46.335 41.085 46.675 ;
        RECT 41.255 46.105 41.585 46.505 ;
        RECT 42.120 46.275 42.735 46.845 ;
        RECT 43.025 46.785 43.290 47.345 ;
        RECT 43.460 46.615 43.630 47.515 ;
        RECT 43.800 46.785 44.155 47.345 ;
        RECT 44.385 46.855 44.905 47.395 ;
        RECT 45.075 47.025 45.595 47.565 ;
        RECT 45.765 47.515 46.045 48.655 ;
        RECT 46.215 47.505 46.545 48.485 ;
        RECT 46.715 47.515 46.975 48.655 ;
        RECT 47.145 47.515 47.530 48.485 ;
        RECT 47.700 48.195 48.025 48.655 ;
        RECT 48.545 48.025 48.825 48.485 ;
        RECT 47.700 47.805 48.825 48.025 ;
        RECT 45.775 47.075 46.110 47.345 ;
        RECT 46.280 46.905 46.450 47.505 ;
        RECT 46.620 47.095 46.955 47.345 ;
        RECT 42.905 46.105 43.120 46.615 ;
        RECT 43.350 46.285 43.630 46.615 ;
        RECT 43.810 46.105 44.050 46.615 ;
        RECT 44.385 46.105 45.595 46.855 ;
        RECT 45.765 46.105 46.075 46.905 ;
        RECT 46.280 46.275 46.975 46.905 ;
        RECT 47.145 46.845 47.425 47.515 ;
        RECT 47.700 47.345 48.150 47.805 ;
        RECT 49.015 47.635 49.415 48.485 ;
        RECT 49.815 48.195 50.085 48.655 ;
        RECT 50.255 48.025 50.540 48.485 ;
        RECT 47.595 47.015 48.150 47.345 ;
        RECT 48.320 47.075 49.415 47.635 ;
        RECT 47.700 46.905 48.150 47.015 ;
        RECT 47.145 46.275 47.530 46.845 ;
        RECT 47.700 46.735 48.825 46.905 ;
        RECT 47.700 46.105 48.025 46.565 ;
        RECT 48.545 46.275 48.825 46.735 ;
        RECT 49.015 46.275 49.415 47.075 ;
        RECT 49.585 47.805 50.540 48.025 ;
        RECT 49.585 46.905 49.795 47.805 ;
        RECT 49.965 47.075 50.655 47.635 ;
        RECT 50.825 47.490 51.115 48.655 ;
        RECT 51.290 47.515 51.565 48.485 ;
        RECT 51.775 47.855 52.055 48.655 ;
        RECT 52.225 48.145 53.415 48.435 ;
        RECT 52.225 47.805 53.395 47.975 ;
        RECT 52.225 47.685 52.395 47.805 ;
        RECT 51.735 47.515 52.395 47.685 ;
        RECT 49.585 46.735 50.540 46.905 ;
        RECT 49.815 46.105 50.085 46.565 ;
        RECT 50.255 46.275 50.540 46.735 ;
        RECT 50.825 46.105 51.115 46.830 ;
        RECT 51.290 46.780 51.460 47.515 ;
        RECT 51.735 47.345 51.905 47.515 ;
        RECT 52.705 47.345 52.900 47.635 ;
        RECT 53.070 47.515 53.395 47.805 ;
        RECT 54.105 47.595 54.435 48.440 ;
        RECT 54.605 47.645 54.775 48.655 ;
        RECT 54.945 47.925 55.285 48.485 ;
        RECT 55.515 48.155 55.830 48.655 ;
        RECT 56.010 48.185 56.895 48.355 ;
        RECT 54.045 47.515 54.435 47.595 ;
        RECT 54.945 47.550 55.840 47.925 ;
        RECT 54.045 47.465 54.260 47.515 ;
        RECT 51.630 47.015 51.905 47.345 ;
        RECT 52.075 47.015 52.900 47.345 ;
        RECT 53.070 47.015 53.415 47.345 ;
        RECT 51.735 46.845 51.905 47.015 ;
        RECT 54.045 46.885 54.215 47.465 ;
        RECT 54.945 47.345 55.135 47.550 ;
        RECT 56.010 47.345 56.180 48.185 ;
        RECT 57.120 48.155 57.370 48.485 ;
        RECT 54.385 47.015 55.135 47.345 ;
        RECT 55.305 47.015 56.180 47.345 ;
        RECT 54.045 46.845 54.270 46.885 ;
        RECT 54.935 46.845 55.135 47.015 ;
        RECT 51.290 46.435 51.565 46.780 ;
        RECT 51.735 46.675 53.400 46.845 ;
        RECT 54.045 46.760 54.425 46.845 ;
        RECT 51.755 46.105 52.135 46.505 ;
        RECT 52.305 46.325 52.475 46.675 ;
        RECT 52.645 46.105 52.975 46.505 ;
        RECT 53.145 46.325 53.400 46.675 ;
        RECT 54.095 46.325 54.425 46.760 ;
        RECT 54.595 46.105 54.765 46.715 ;
        RECT 54.935 46.320 55.265 46.845 ;
        RECT 55.525 46.105 55.735 46.635 ;
        RECT 56.010 46.555 56.180 47.015 ;
        RECT 56.350 47.055 56.670 48.015 ;
        RECT 56.840 47.265 57.030 47.985 ;
        RECT 57.200 47.085 57.370 48.155 ;
        RECT 57.540 47.855 57.710 48.655 ;
        RECT 57.880 48.210 58.985 48.380 ;
        RECT 57.880 47.595 58.050 48.210 ;
        RECT 59.195 48.060 59.445 48.485 ;
        RECT 59.615 48.195 59.880 48.655 ;
        RECT 58.220 47.675 58.750 48.040 ;
        RECT 59.195 47.930 59.500 48.060 ;
        RECT 57.540 47.505 58.050 47.595 ;
        RECT 57.540 47.335 58.410 47.505 ;
        RECT 57.540 47.265 57.710 47.335 ;
        RECT 57.830 47.085 58.030 47.115 ;
        RECT 56.350 46.725 56.815 47.055 ;
        RECT 57.200 46.785 58.030 47.085 ;
        RECT 57.200 46.555 57.370 46.785 ;
        RECT 56.010 46.385 56.795 46.555 ;
        RECT 56.965 46.385 57.370 46.555 ;
        RECT 57.550 46.105 57.920 46.605 ;
        RECT 58.240 46.555 58.410 47.335 ;
        RECT 58.580 46.975 58.750 47.675 ;
        RECT 58.920 47.145 59.160 47.740 ;
        RECT 58.580 46.755 59.105 46.975 ;
        RECT 59.330 46.825 59.500 47.930 ;
        RECT 59.275 46.695 59.500 46.825 ;
        RECT 59.670 46.735 59.950 47.685 ;
        RECT 59.275 46.555 59.445 46.695 ;
        RECT 58.240 46.385 58.915 46.555 ;
        RECT 59.110 46.385 59.445 46.555 ;
        RECT 59.615 46.105 59.865 46.565 ;
        RECT 60.120 46.365 60.305 48.485 ;
        RECT 60.475 48.155 60.805 48.655 ;
        RECT 60.975 47.985 61.145 48.485 ;
        RECT 61.405 48.145 62.600 48.435 ;
        RECT 60.480 47.815 61.145 47.985 ;
        RECT 60.480 46.825 60.710 47.815 ;
        RECT 61.425 47.805 62.590 47.975 ;
        RECT 62.770 47.855 63.050 48.655 ;
        RECT 60.880 46.995 61.230 47.645 ;
        RECT 61.425 47.515 61.755 47.805 ;
        RECT 62.420 47.685 62.590 47.805 ;
        RECT 61.925 47.345 62.150 47.635 ;
        RECT 62.420 47.515 63.090 47.685 ;
        RECT 63.260 47.515 63.535 48.485 ;
        RECT 62.920 47.345 63.090 47.515 ;
        RECT 61.405 47.015 61.755 47.345 ;
        RECT 61.925 47.015 62.750 47.345 ;
        RECT 62.920 47.015 63.195 47.345 ;
        RECT 62.920 46.845 63.090 47.015 ;
        RECT 60.480 46.655 61.145 46.825 ;
        RECT 60.475 46.105 60.805 46.485 ;
        RECT 60.975 46.365 61.145 46.655 ;
        RECT 61.425 46.675 63.090 46.845 ;
        RECT 63.365 46.780 63.535 47.515 ;
        RECT 63.705 47.450 63.995 48.655 ;
        RECT 64.255 47.985 64.425 48.485 ;
        RECT 64.595 48.155 64.925 48.655 ;
        RECT 64.255 47.815 64.920 47.985 ;
        RECT 64.170 46.995 64.520 47.645 ;
        RECT 61.425 46.325 61.680 46.675 ;
        RECT 61.850 46.105 62.180 46.505 ;
        RECT 62.350 46.325 62.520 46.675 ;
        RECT 62.690 46.105 63.070 46.505 ;
        RECT 63.260 46.435 63.535 46.780 ;
        RECT 63.705 46.105 63.995 46.935 ;
        RECT 64.690 46.825 64.920 47.815 ;
        RECT 64.255 46.655 64.920 46.825 ;
        RECT 64.255 46.365 64.425 46.655 ;
        RECT 64.595 46.105 64.925 46.485 ;
        RECT 65.095 46.365 65.280 48.485 ;
        RECT 65.520 48.195 65.785 48.655 ;
        RECT 65.955 48.060 66.205 48.485 ;
        RECT 66.415 48.210 67.520 48.380 ;
        RECT 65.900 47.930 66.205 48.060 ;
        RECT 65.450 46.735 65.730 47.685 ;
        RECT 65.900 46.825 66.070 47.930 ;
        RECT 66.240 47.145 66.480 47.740 ;
        RECT 66.650 47.675 67.180 48.040 ;
        RECT 66.650 46.975 66.820 47.675 ;
        RECT 67.350 47.595 67.520 48.210 ;
        RECT 67.690 47.855 67.860 48.655 ;
        RECT 68.030 48.155 68.280 48.485 ;
        RECT 68.505 48.185 69.390 48.355 ;
        RECT 67.350 47.505 67.860 47.595 ;
        RECT 65.900 46.695 66.125 46.825 ;
        RECT 66.295 46.755 66.820 46.975 ;
        RECT 66.990 47.335 67.860 47.505 ;
        RECT 65.535 46.105 65.785 46.565 ;
        RECT 65.955 46.555 66.125 46.695 ;
        RECT 66.990 46.555 67.160 47.335 ;
        RECT 67.690 47.265 67.860 47.335 ;
        RECT 67.370 47.085 67.570 47.115 ;
        RECT 68.030 47.085 68.200 48.155 ;
        RECT 68.370 47.265 68.560 47.985 ;
        RECT 67.370 46.785 68.200 47.085 ;
        RECT 68.730 47.055 69.050 48.015 ;
        RECT 65.955 46.385 66.290 46.555 ;
        RECT 66.485 46.385 67.160 46.555 ;
        RECT 67.480 46.105 67.850 46.605 ;
        RECT 68.030 46.555 68.200 46.785 ;
        RECT 68.585 46.725 69.050 47.055 ;
        RECT 69.220 47.345 69.390 48.185 ;
        RECT 69.570 48.155 69.885 48.655 ;
        RECT 70.115 47.925 70.455 48.485 ;
        RECT 69.560 47.550 70.455 47.925 ;
        RECT 70.625 47.645 70.795 48.655 ;
        RECT 70.265 47.345 70.455 47.550 ;
        RECT 70.965 47.595 71.295 48.440 ;
        RECT 71.465 47.740 71.635 48.655 ;
        RECT 70.965 47.515 71.355 47.595 ;
        RECT 71.140 47.465 71.355 47.515 ;
        RECT 69.220 47.015 70.095 47.345 ;
        RECT 70.265 47.015 71.015 47.345 ;
        RECT 69.220 46.555 69.390 47.015 ;
        RECT 70.265 46.845 70.465 47.015 ;
        RECT 71.185 46.885 71.355 47.465 ;
        RECT 71.130 46.845 71.355 46.885 ;
        RECT 68.030 46.385 68.435 46.555 ;
        RECT 68.605 46.385 69.390 46.555 ;
        RECT 69.665 46.105 69.875 46.635 ;
        RECT 70.135 46.320 70.465 46.845 ;
        RECT 70.975 46.760 71.355 46.845 ;
        RECT 71.985 47.515 72.260 48.485 ;
        RECT 72.470 47.855 72.750 48.655 ;
        RECT 72.920 48.145 74.535 48.475 ;
        RECT 72.920 47.805 74.095 47.975 ;
        RECT 72.920 47.685 73.090 47.805 ;
        RECT 72.430 47.515 73.090 47.685 ;
        RECT 71.985 46.780 72.155 47.515 ;
        RECT 72.430 47.345 72.600 47.515 ;
        RECT 73.350 47.345 73.595 47.635 ;
        RECT 73.765 47.515 74.095 47.805 ;
        RECT 74.355 47.345 74.525 47.905 ;
        RECT 74.775 47.515 75.035 48.655 ;
        RECT 75.205 47.565 76.415 48.655 ;
        RECT 72.325 47.015 72.600 47.345 ;
        RECT 72.770 47.015 73.595 47.345 ;
        RECT 73.810 47.015 74.525 47.345 ;
        RECT 74.695 47.095 75.030 47.345 ;
        RECT 72.430 46.845 72.600 47.015 ;
        RECT 74.275 46.925 74.525 47.015 ;
        RECT 70.635 46.105 70.805 46.715 ;
        RECT 70.975 46.325 71.305 46.760 ;
        RECT 71.475 46.105 71.645 46.620 ;
        RECT 71.985 46.435 72.260 46.780 ;
        RECT 72.430 46.675 74.095 46.845 ;
        RECT 72.450 46.105 72.825 46.505 ;
        RECT 72.995 46.325 73.165 46.675 ;
        RECT 73.335 46.105 73.665 46.505 ;
        RECT 73.835 46.275 74.095 46.675 ;
        RECT 74.275 46.505 74.605 46.925 ;
        RECT 74.775 46.105 75.035 46.925 ;
        RECT 75.205 46.855 75.725 47.395 ;
        RECT 75.895 47.025 76.415 47.565 ;
        RECT 76.585 47.490 76.875 48.655 ;
        RECT 77.250 47.685 77.580 48.485 ;
        RECT 77.750 47.855 78.080 48.655 ;
        RECT 78.380 47.685 78.710 48.485 ;
        RECT 79.355 47.855 79.605 48.655 ;
        RECT 77.250 47.515 79.685 47.685 ;
        RECT 79.875 47.515 80.045 48.655 ;
        RECT 80.215 47.515 80.555 48.485 ;
        RECT 81.275 47.985 81.445 48.485 ;
        RECT 81.615 48.155 81.945 48.655 ;
        RECT 81.275 47.815 81.940 47.985 ;
        RECT 77.045 47.095 77.395 47.345 ;
        RECT 77.580 46.885 77.750 47.515 ;
        RECT 77.920 47.095 78.250 47.295 ;
        RECT 78.420 47.095 78.750 47.295 ;
        RECT 78.920 47.095 79.340 47.295 ;
        RECT 79.515 47.265 79.685 47.515 ;
        RECT 79.515 47.095 80.210 47.265 ;
        RECT 75.205 46.105 76.415 46.855 ;
        RECT 76.585 46.105 76.875 46.830 ;
        RECT 77.250 46.275 77.750 46.885 ;
        RECT 78.380 46.755 79.605 46.925 ;
        RECT 80.380 46.905 80.555 47.515 ;
        RECT 81.190 46.995 81.540 47.645 ;
        RECT 78.380 46.275 78.710 46.755 ;
        RECT 78.880 46.105 79.105 46.565 ;
        RECT 79.275 46.275 79.605 46.755 ;
        RECT 79.795 46.105 80.045 46.905 ;
        RECT 80.215 46.275 80.555 46.905 ;
        RECT 81.710 46.825 81.940 47.815 ;
        RECT 81.275 46.655 81.940 46.825 ;
        RECT 81.275 46.365 81.445 46.655 ;
        RECT 81.615 46.105 81.945 46.485 ;
        RECT 82.115 46.365 82.300 48.485 ;
        RECT 82.540 48.195 82.805 48.655 ;
        RECT 82.975 48.060 83.225 48.485 ;
        RECT 83.435 48.210 84.540 48.380 ;
        RECT 82.920 47.930 83.225 48.060 ;
        RECT 82.470 46.735 82.750 47.685 ;
        RECT 82.920 46.825 83.090 47.930 ;
        RECT 83.260 47.145 83.500 47.740 ;
        RECT 83.670 47.675 84.200 48.040 ;
        RECT 83.670 46.975 83.840 47.675 ;
        RECT 84.370 47.595 84.540 48.210 ;
        RECT 84.710 47.855 84.880 48.655 ;
        RECT 85.050 48.155 85.300 48.485 ;
        RECT 85.525 48.185 86.410 48.355 ;
        RECT 84.370 47.505 84.880 47.595 ;
        RECT 82.920 46.695 83.145 46.825 ;
        RECT 83.315 46.755 83.840 46.975 ;
        RECT 84.010 47.335 84.880 47.505 ;
        RECT 82.555 46.105 82.805 46.565 ;
        RECT 82.975 46.555 83.145 46.695 ;
        RECT 84.010 46.555 84.180 47.335 ;
        RECT 84.710 47.265 84.880 47.335 ;
        RECT 84.390 47.085 84.590 47.115 ;
        RECT 85.050 47.085 85.220 48.155 ;
        RECT 85.390 47.265 85.580 47.985 ;
        RECT 84.390 46.785 85.220 47.085 ;
        RECT 85.750 47.055 86.070 48.015 ;
        RECT 82.975 46.385 83.310 46.555 ;
        RECT 83.505 46.385 84.180 46.555 ;
        RECT 84.500 46.105 84.870 46.605 ;
        RECT 85.050 46.555 85.220 46.785 ;
        RECT 85.605 46.725 86.070 47.055 ;
        RECT 86.240 47.345 86.410 48.185 ;
        RECT 86.590 48.155 86.905 48.655 ;
        RECT 87.135 47.925 87.475 48.485 ;
        RECT 86.580 47.550 87.475 47.925 ;
        RECT 87.645 47.645 87.815 48.655 ;
        RECT 87.285 47.345 87.475 47.550 ;
        RECT 87.985 47.595 88.315 48.440 ;
        RECT 87.985 47.515 88.375 47.595 ;
        RECT 88.160 47.465 88.375 47.515 ;
        RECT 86.240 47.015 87.115 47.345 ;
        RECT 87.285 47.015 88.035 47.345 ;
        RECT 86.240 46.555 86.410 47.015 ;
        RECT 87.285 46.845 87.485 47.015 ;
        RECT 88.205 46.885 88.375 47.465 ;
        RECT 88.545 47.565 89.755 48.655 ;
        RECT 88.545 47.025 89.065 47.565 ;
        RECT 88.150 46.845 88.375 46.885 ;
        RECT 89.235 46.855 89.755 47.395 ;
        RECT 85.050 46.385 85.455 46.555 ;
        RECT 85.625 46.385 86.410 46.555 ;
        RECT 86.685 46.105 86.895 46.635 ;
        RECT 87.155 46.320 87.485 46.845 ;
        RECT 87.995 46.760 88.375 46.845 ;
        RECT 87.655 46.105 87.825 46.715 ;
        RECT 87.995 46.325 88.325 46.760 ;
        RECT 88.545 46.105 89.755 46.855 ;
        RECT 12.100 45.935 89.840 46.105 ;
        RECT 12.185 45.185 13.395 45.935 ;
        RECT 12.185 44.645 12.705 45.185 ;
        RECT 13.575 45.125 13.845 45.935 ;
        RECT 14.015 45.125 14.345 45.765 ;
        RECT 14.515 45.125 14.755 45.935 ;
        RECT 15.035 45.385 15.205 45.675 ;
        RECT 15.375 45.555 15.705 45.935 ;
        RECT 15.035 45.215 15.700 45.385 ;
        RECT 12.875 44.475 13.395 45.015 ;
        RECT 13.565 44.695 13.915 44.945 ;
        RECT 14.085 44.525 14.255 45.125 ;
        RECT 14.425 44.695 14.775 44.945 ;
        RECT 12.185 43.385 13.395 44.475 ;
        RECT 13.575 43.385 13.905 44.525 ;
        RECT 14.085 44.355 14.765 44.525 ;
        RECT 14.950 44.395 15.300 45.045 ;
        RECT 14.435 43.570 14.765 44.355 ;
        RECT 15.470 44.225 15.700 45.215 ;
        RECT 15.035 44.055 15.700 44.225 ;
        RECT 15.035 43.555 15.205 44.055 ;
        RECT 15.375 43.385 15.705 43.885 ;
        RECT 15.875 43.555 16.060 45.675 ;
        RECT 16.315 45.475 16.565 45.935 ;
        RECT 16.735 45.485 17.070 45.655 ;
        RECT 17.265 45.485 17.940 45.655 ;
        RECT 16.735 45.345 16.905 45.485 ;
        RECT 16.230 44.355 16.510 45.305 ;
        RECT 16.680 45.215 16.905 45.345 ;
        RECT 16.680 44.110 16.850 45.215 ;
        RECT 17.075 45.065 17.600 45.285 ;
        RECT 17.020 44.300 17.260 44.895 ;
        RECT 17.430 44.365 17.600 45.065 ;
        RECT 17.770 44.705 17.940 45.485 ;
        RECT 18.260 45.435 18.630 45.935 ;
        RECT 18.810 45.485 19.215 45.655 ;
        RECT 19.385 45.485 20.170 45.655 ;
        RECT 18.810 45.255 18.980 45.485 ;
        RECT 18.150 44.955 18.980 45.255 ;
        RECT 19.365 44.985 19.830 45.315 ;
        RECT 18.150 44.925 18.350 44.955 ;
        RECT 18.470 44.705 18.640 44.775 ;
        RECT 17.770 44.535 18.640 44.705 ;
        RECT 18.130 44.445 18.640 44.535 ;
        RECT 16.680 43.980 16.985 44.110 ;
        RECT 17.430 44.000 17.960 44.365 ;
        RECT 16.300 43.385 16.565 43.845 ;
        RECT 16.735 43.555 16.985 43.980 ;
        RECT 18.130 43.830 18.300 44.445 ;
        RECT 17.195 43.660 18.300 43.830 ;
        RECT 18.470 43.385 18.640 44.185 ;
        RECT 18.810 43.885 18.980 44.955 ;
        RECT 19.150 44.055 19.340 44.775 ;
        RECT 19.510 44.025 19.830 44.985 ;
        RECT 20.000 45.025 20.170 45.485 ;
        RECT 20.445 45.405 20.655 45.935 ;
        RECT 20.915 45.195 21.245 45.720 ;
        RECT 21.415 45.325 21.585 45.935 ;
        RECT 21.755 45.280 22.085 45.715 ;
        RECT 22.305 45.285 22.565 45.765 ;
        RECT 22.735 45.395 22.985 45.935 ;
        RECT 21.755 45.195 22.135 45.280 ;
        RECT 21.045 45.025 21.245 45.195 ;
        RECT 21.910 45.155 22.135 45.195 ;
        RECT 20.000 44.695 20.875 45.025 ;
        RECT 21.045 44.695 21.795 45.025 ;
        RECT 18.810 43.555 19.060 43.885 ;
        RECT 20.000 43.855 20.170 44.695 ;
        RECT 21.045 44.490 21.235 44.695 ;
        RECT 21.965 44.575 22.135 45.155 ;
        RECT 21.920 44.525 22.135 44.575 ;
        RECT 20.340 44.115 21.235 44.490 ;
        RECT 21.745 44.445 22.135 44.525 ;
        RECT 19.285 43.685 20.170 43.855 ;
        RECT 20.350 43.385 20.665 43.885 ;
        RECT 20.895 43.555 21.235 44.115 ;
        RECT 21.405 43.385 21.575 44.395 ;
        RECT 21.745 43.600 22.075 44.445 ;
        RECT 22.305 44.255 22.475 45.285 ;
        RECT 23.155 45.230 23.375 45.715 ;
        RECT 22.645 44.635 22.875 45.030 ;
        RECT 23.045 44.805 23.375 45.230 ;
        RECT 23.545 45.555 24.435 45.725 ;
        RECT 23.545 44.830 23.715 45.555 ;
        RECT 23.885 45.000 24.435 45.385 ;
        RECT 25.270 45.155 25.770 45.765 ;
        RECT 23.545 44.760 24.435 44.830 ;
        RECT 23.540 44.735 24.435 44.760 ;
        RECT 23.530 44.720 24.435 44.735 ;
        RECT 23.525 44.705 24.435 44.720 ;
        RECT 23.515 44.700 24.435 44.705 ;
        RECT 23.510 44.690 24.435 44.700 ;
        RECT 25.065 44.695 25.415 44.945 ;
        RECT 23.505 44.680 24.435 44.690 ;
        RECT 23.495 44.675 24.435 44.680 ;
        RECT 23.485 44.665 24.435 44.675 ;
        RECT 23.475 44.660 24.435 44.665 ;
        RECT 23.475 44.655 23.810 44.660 ;
        RECT 23.460 44.650 23.810 44.655 ;
        RECT 23.445 44.640 23.810 44.650 ;
        RECT 23.420 44.635 23.810 44.640 ;
        RECT 22.645 44.630 23.810 44.635 ;
        RECT 22.645 44.595 23.780 44.630 ;
        RECT 22.645 44.570 23.745 44.595 ;
        RECT 22.645 44.540 23.715 44.570 ;
        RECT 22.645 44.510 23.695 44.540 ;
        RECT 22.645 44.480 23.675 44.510 ;
        RECT 22.645 44.470 23.605 44.480 ;
        RECT 22.645 44.460 23.580 44.470 ;
        RECT 22.645 44.445 23.560 44.460 ;
        RECT 22.645 44.430 23.540 44.445 ;
        RECT 22.750 44.420 23.535 44.430 ;
        RECT 22.750 44.385 23.520 44.420 ;
        RECT 22.305 43.555 22.580 44.255 ;
        RECT 22.750 44.135 23.505 44.385 ;
        RECT 23.675 44.065 24.005 44.310 ;
        RECT 24.175 44.210 24.435 44.660 ;
        RECT 25.600 44.525 25.770 45.155 ;
        RECT 26.400 45.285 26.730 45.765 ;
        RECT 26.900 45.475 27.125 45.935 ;
        RECT 27.295 45.285 27.625 45.765 ;
        RECT 26.400 45.115 27.625 45.285 ;
        RECT 27.815 45.135 28.065 45.935 ;
        RECT 28.235 45.135 28.575 45.765 ;
        RECT 28.750 45.445 29.005 45.935 ;
        RECT 29.175 45.425 30.405 45.765 ;
        RECT 25.940 44.745 26.270 44.945 ;
        RECT 26.440 44.745 26.770 44.945 ;
        RECT 26.940 44.745 27.360 44.945 ;
        RECT 27.535 44.775 28.230 44.945 ;
        RECT 27.535 44.525 27.705 44.775 ;
        RECT 28.400 44.525 28.575 45.135 ;
        RECT 28.770 44.695 28.990 45.275 ;
        RECT 29.175 44.525 29.355 45.425 ;
        RECT 29.525 44.695 29.900 45.255 ;
        RECT 30.075 45.195 30.405 45.425 ;
        RECT 30.675 45.385 30.845 45.675 ;
        RECT 31.015 45.555 31.345 45.935 ;
        RECT 30.675 45.215 31.340 45.385 ;
        RECT 30.105 44.695 30.415 45.025 ;
        RECT 25.270 44.355 27.705 44.525 ;
        RECT 23.820 44.040 24.005 44.065 ;
        RECT 23.820 43.940 24.435 44.040 ;
        RECT 22.750 43.385 23.005 43.930 ;
        RECT 23.175 43.555 23.655 43.895 ;
        RECT 23.830 43.385 24.435 43.940 ;
        RECT 25.270 43.555 25.600 44.355 ;
        RECT 25.770 43.385 26.100 44.185 ;
        RECT 26.400 43.555 26.730 44.355 ;
        RECT 27.375 43.385 27.625 44.185 ;
        RECT 27.895 43.385 28.065 44.525 ;
        RECT 28.235 43.555 28.575 44.525 ;
        RECT 28.750 43.385 29.005 44.525 ;
        RECT 29.175 44.355 30.405 44.525 ;
        RECT 30.590 44.395 30.940 45.045 ;
        RECT 29.175 43.555 29.505 44.355 ;
        RECT 29.675 43.385 29.905 44.185 ;
        RECT 30.075 43.555 30.405 44.355 ;
        RECT 31.110 44.225 31.340 45.215 ;
        RECT 30.675 44.055 31.340 44.225 ;
        RECT 30.675 43.555 30.845 44.055 ;
        RECT 31.015 43.385 31.345 43.885 ;
        RECT 31.515 43.555 31.700 45.675 ;
        RECT 31.955 45.475 32.205 45.935 ;
        RECT 32.375 45.485 32.710 45.655 ;
        RECT 32.905 45.485 33.580 45.655 ;
        RECT 32.375 45.345 32.545 45.485 ;
        RECT 31.870 44.355 32.150 45.305 ;
        RECT 32.320 45.215 32.545 45.345 ;
        RECT 32.320 44.110 32.490 45.215 ;
        RECT 32.715 45.065 33.240 45.285 ;
        RECT 32.660 44.300 32.900 44.895 ;
        RECT 33.070 44.365 33.240 45.065 ;
        RECT 33.410 44.705 33.580 45.485 ;
        RECT 33.900 45.435 34.270 45.935 ;
        RECT 34.450 45.485 34.855 45.655 ;
        RECT 35.025 45.485 35.810 45.655 ;
        RECT 34.450 45.255 34.620 45.485 ;
        RECT 33.790 44.955 34.620 45.255 ;
        RECT 35.005 44.985 35.470 45.315 ;
        RECT 33.790 44.925 33.990 44.955 ;
        RECT 34.110 44.705 34.280 44.775 ;
        RECT 33.410 44.535 34.280 44.705 ;
        RECT 33.770 44.445 34.280 44.535 ;
        RECT 32.320 43.980 32.625 44.110 ;
        RECT 33.070 44.000 33.600 44.365 ;
        RECT 31.940 43.385 32.205 43.845 ;
        RECT 32.375 43.555 32.625 43.980 ;
        RECT 33.770 43.830 33.940 44.445 ;
        RECT 32.835 43.660 33.940 43.830 ;
        RECT 34.110 43.385 34.280 44.185 ;
        RECT 34.450 43.885 34.620 44.955 ;
        RECT 34.790 44.055 34.980 44.775 ;
        RECT 35.150 44.025 35.470 44.985 ;
        RECT 35.640 45.025 35.810 45.485 ;
        RECT 36.085 45.405 36.295 45.935 ;
        RECT 36.555 45.195 36.885 45.720 ;
        RECT 37.055 45.325 37.225 45.935 ;
        RECT 37.395 45.280 37.725 45.715 ;
        RECT 37.395 45.195 37.775 45.280 ;
        RECT 37.945 45.210 38.235 45.935 ;
        RECT 38.495 45.385 38.665 45.675 ;
        RECT 38.835 45.555 39.165 45.935 ;
        RECT 38.495 45.215 39.160 45.385 ;
        RECT 36.685 45.025 36.885 45.195 ;
        RECT 37.550 45.155 37.775 45.195 ;
        RECT 35.640 44.695 36.515 45.025 ;
        RECT 36.685 44.695 37.435 45.025 ;
        RECT 34.450 43.555 34.700 43.885 ;
        RECT 35.640 43.855 35.810 44.695 ;
        RECT 36.685 44.490 36.875 44.695 ;
        RECT 37.605 44.575 37.775 45.155 ;
        RECT 37.560 44.525 37.775 44.575 ;
        RECT 35.980 44.115 36.875 44.490 ;
        RECT 37.385 44.445 37.775 44.525 ;
        RECT 34.925 43.685 35.810 43.855 ;
        RECT 35.990 43.385 36.305 43.885 ;
        RECT 36.535 43.555 36.875 44.115 ;
        RECT 37.045 43.385 37.215 44.395 ;
        RECT 37.385 43.600 37.715 44.445 ;
        RECT 37.945 43.385 38.235 44.550 ;
        RECT 38.410 44.395 38.760 45.045 ;
        RECT 38.930 44.225 39.160 45.215 ;
        RECT 38.495 44.055 39.160 44.225 ;
        RECT 38.495 43.555 38.665 44.055 ;
        RECT 38.835 43.385 39.165 43.885 ;
        RECT 39.335 43.555 39.520 45.675 ;
        RECT 39.775 45.475 40.025 45.935 ;
        RECT 40.195 45.485 40.530 45.655 ;
        RECT 40.725 45.485 41.400 45.655 ;
        RECT 40.195 45.345 40.365 45.485 ;
        RECT 39.690 44.355 39.970 45.305 ;
        RECT 40.140 45.215 40.365 45.345 ;
        RECT 40.140 44.110 40.310 45.215 ;
        RECT 40.535 45.065 41.060 45.285 ;
        RECT 40.480 44.300 40.720 44.895 ;
        RECT 40.890 44.365 41.060 45.065 ;
        RECT 41.230 44.705 41.400 45.485 ;
        RECT 41.720 45.435 42.090 45.935 ;
        RECT 42.270 45.485 42.675 45.655 ;
        RECT 42.845 45.485 43.630 45.655 ;
        RECT 42.270 45.255 42.440 45.485 ;
        RECT 41.610 44.955 42.440 45.255 ;
        RECT 42.825 44.985 43.290 45.315 ;
        RECT 41.610 44.925 41.810 44.955 ;
        RECT 41.930 44.705 42.100 44.775 ;
        RECT 41.230 44.535 42.100 44.705 ;
        RECT 41.590 44.445 42.100 44.535 ;
        RECT 40.140 43.980 40.445 44.110 ;
        RECT 40.890 44.000 41.420 44.365 ;
        RECT 39.760 43.385 40.025 43.845 ;
        RECT 40.195 43.555 40.445 43.980 ;
        RECT 41.590 43.830 41.760 44.445 ;
        RECT 40.655 43.660 41.760 43.830 ;
        RECT 41.930 43.385 42.100 44.185 ;
        RECT 42.270 43.885 42.440 44.955 ;
        RECT 42.610 44.055 42.800 44.775 ;
        RECT 42.970 44.025 43.290 44.985 ;
        RECT 43.460 45.025 43.630 45.485 ;
        RECT 43.905 45.405 44.115 45.935 ;
        RECT 44.375 45.195 44.705 45.720 ;
        RECT 44.875 45.325 45.045 45.935 ;
        RECT 45.215 45.280 45.545 45.715 ;
        RECT 45.770 45.405 46.060 45.755 ;
        RECT 46.255 45.575 46.585 45.935 ;
        RECT 46.755 45.405 46.985 45.710 ;
        RECT 45.215 45.195 45.595 45.280 ;
        RECT 45.770 45.235 46.985 45.405 ;
        RECT 47.175 45.595 47.345 45.630 ;
        RECT 47.175 45.425 47.375 45.595 ;
        RECT 44.505 45.025 44.705 45.195 ;
        RECT 45.370 45.155 45.595 45.195 ;
        RECT 43.460 44.695 44.335 45.025 ;
        RECT 44.505 44.695 45.255 45.025 ;
        RECT 42.270 43.555 42.520 43.885 ;
        RECT 43.460 43.855 43.630 44.695 ;
        RECT 44.505 44.490 44.695 44.695 ;
        RECT 45.425 44.575 45.595 45.155 ;
        RECT 47.175 45.065 47.345 45.425 ;
        RECT 45.830 44.915 46.090 45.025 ;
        RECT 45.825 44.745 46.090 44.915 ;
        RECT 45.830 44.695 46.090 44.745 ;
        RECT 46.270 44.695 46.655 45.025 ;
        RECT 46.825 44.895 47.345 45.065 ;
        RECT 47.605 45.195 48.070 45.740 ;
        RECT 45.380 44.525 45.595 44.575 ;
        RECT 43.800 44.115 44.695 44.490 ;
        RECT 45.205 44.445 45.595 44.525 ;
        RECT 42.745 43.685 43.630 43.855 ;
        RECT 43.810 43.385 44.125 43.885 ;
        RECT 44.355 43.555 44.695 44.115 ;
        RECT 44.865 43.385 45.035 44.395 ;
        RECT 45.205 43.600 45.535 44.445 ;
        RECT 45.770 43.385 46.090 44.525 ;
        RECT 46.270 43.645 46.465 44.695 ;
        RECT 46.825 44.515 46.995 44.895 ;
        RECT 46.645 44.235 46.995 44.515 ;
        RECT 47.185 44.365 47.430 44.725 ;
        RECT 47.605 44.235 47.775 45.195 ;
        RECT 48.575 45.115 48.745 45.935 ;
        RECT 48.915 45.285 49.245 45.765 ;
        RECT 49.415 45.545 49.765 45.935 ;
        RECT 49.935 45.365 50.165 45.765 ;
        RECT 49.655 45.285 50.165 45.365 ;
        RECT 48.915 45.195 50.165 45.285 ;
        RECT 50.335 45.195 50.655 45.675 ;
        RECT 51.835 45.385 52.005 45.675 ;
        RECT 52.175 45.555 52.505 45.935 ;
        RECT 51.835 45.215 52.500 45.385 ;
        RECT 48.915 45.115 49.825 45.195 ;
        RECT 47.945 44.575 48.190 45.025 ;
        RECT 48.450 44.745 49.145 44.945 ;
        RECT 49.315 44.775 49.915 44.945 ;
        RECT 49.315 44.575 49.485 44.775 ;
        RECT 50.145 44.605 50.315 45.025 ;
        RECT 47.945 44.405 49.485 44.575 ;
        RECT 49.655 44.435 50.315 44.605 ;
        RECT 49.655 44.235 49.825 44.435 ;
        RECT 50.485 44.265 50.655 45.195 ;
        RECT 51.750 44.395 52.100 45.045 ;
        RECT 46.645 43.555 46.975 44.235 ;
        RECT 47.175 43.385 47.430 44.185 ;
        RECT 47.605 44.065 49.825 44.235 ;
        RECT 49.995 44.065 50.655 44.265 ;
        RECT 52.270 44.225 52.500 45.215 ;
        RECT 47.605 43.385 47.905 43.895 ;
        RECT 48.075 43.555 48.405 44.065 ;
        RECT 49.995 43.895 50.165 44.065 ;
        RECT 51.835 44.055 52.500 44.225 ;
        RECT 48.575 43.385 49.205 43.895 ;
        RECT 49.785 43.725 50.165 43.895 ;
        RECT 50.335 43.385 50.635 43.895 ;
        RECT 51.835 43.555 52.005 44.055 ;
        RECT 52.175 43.385 52.505 43.885 ;
        RECT 52.675 43.555 52.860 45.675 ;
        RECT 53.115 45.475 53.365 45.935 ;
        RECT 53.535 45.485 53.870 45.655 ;
        RECT 54.065 45.485 54.740 45.655 ;
        RECT 53.535 45.345 53.705 45.485 ;
        RECT 53.030 44.355 53.310 45.305 ;
        RECT 53.480 45.215 53.705 45.345 ;
        RECT 53.480 44.110 53.650 45.215 ;
        RECT 53.875 45.065 54.400 45.285 ;
        RECT 53.820 44.300 54.060 44.895 ;
        RECT 54.230 44.365 54.400 45.065 ;
        RECT 54.570 44.705 54.740 45.485 ;
        RECT 55.060 45.435 55.430 45.935 ;
        RECT 55.610 45.485 56.015 45.655 ;
        RECT 56.185 45.485 56.970 45.655 ;
        RECT 55.610 45.255 55.780 45.485 ;
        RECT 54.950 44.955 55.780 45.255 ;
        RECT 56.165 44.985 56.630 45.315 ;
        RECT 54.950 44.925 55.150 44.955 ;
        RECT 55.270 44.705 55.440 44.775 ;
        RECT 54.570 44.535 55.440 44.705 ;
        RECT 54.930 44.445 55.440 44.535 ;
        RECT 53.480 43.980 53.785 44.110 ;
        RECT 54.230 44.000 54.760 44.365 ;
        RECT 53.100 43.385 53.365 43.845 ;
        RECT 53.535 43.555 53.785 43.980 ;
        RECT 54.930 43.830 55.100 44.445 ;
        RECT 53.995 43.660 55.100 43.830 ;
        RECT 55.270 43.385 55.440 44.185 ;
        RECT 55.610 43.885 55.780 44.955 ;
        RECT 55.950 44.055 56.140 44.775 ;
        RECT 56.310 44.025 56.630 44.985 ;
        RECT 56.800 45.025 56.970 45.485 ;
        RECT 57.245 45.405 57.455 45.935 ;
        RECT 57.715 45.195 58.045 45.720 ;
        RECT 58.215 45.325 58.385 45.935 ;
        RECT 58.555 45.280 58.885 45.715 ;
        RECT 58.555 45.195 58.935 45.280 ;
        RECT 57.845 45.025 58.045 45.195 ;
        RECT 58.710 45.155 58.935 45.195 ;
        RECT 56.800 44.695 57.675 45.025 ;
        RECT 57.845 44.695 58.595 45.025 ;
        RECT 55.610 43.555 55.860 43.885 ;
        RECT 56.800 43.855 56.970 44.695 ;
        RECT 57.845 44.490 58.035 44.695 ;
        RECT 58.765 44.575 58.935 45.155 ;
        RECT 58.720 44.525 58.935 44.575 ;
        RECT 57.140 44.115 58.035 44.490 ;
        RECT 58.545 44.445 58.935 44.525 ;
        RECT 59.105 45.195 59.490 45.765 ;
        RECT 59.660 45.475 59.985 45.935 ;
        RECT 60.505 45.305 60.785 45.765 ;
        RECT 59.105 44.525 59.385 45.195 ;
        RECT 59.660 45.135 60.785 45.305 ;
        RECT 59.660 45.025 60.110 45.135 ;
        RECT 59.555 44.695 60.110 45.025 ;
        RECT 60.975 44.965 61.375 45.765 ;
        RECT 61.775 45.475 62.045 45.935 ;
        RECT 62.215 45.305 62.500 45.765 ;
        RECT 56.085 43.685 56.970 43.855 ;
        RECT 57.150 43.385 57.465 43.885 ;
        RECT 57.695 43.555 58.035 44.115 ;
        RECT 58.205 43.385 58.375 44.395 ;
        RECT 58.545 43.600 58.875 44.445 ;
        RECT 59.105 43.555 59.490 44.525 ;
        RECT 59.660 44.235 60.110 44.695 ;
        RECT 60.280 44.405 61.375 44.965 ;
        RECT 59.660 44.015 60.785 44.235 ;
        RECT 59.660 43.385 59.985 43.845 ;
        RECT 60.505 43.555 60.785 44.015 ;
        RECT 60.975 43.555 61.375 44.405 ;
        RECT 61.545 45.135 62.500 45.305 ;
        RECT 63.705 45.210 63.995 45.935 ;
        RECT 64.255 45.385 64.425 45.675 ;
        RECT 64.595 45.555 64.925 45.935 ;
        RECT 64.255 45.215 64.920 45.385 ;
        RECT 61.545 44.235 61.755 45.135 ;
        RECT 61.925 44.405 62.615 44.965 ;
        RECT 61.545 44.015 62.500 44.235 ;
        RECT 61.775 43.385 62.045 43.845 ;
        RECT 62.215 43.555 62.500 44.015 ;
        RECT 63.705 43.385 63.995 44.550 ;
        RECT 64.170 44.395 64.520 45.045 ;
        RECT 64.690 44.225 64.920 45.215 ;
        RECT 64.255 44.055 64.920 44.225 ;
        RECT 64.255 43.555 64.425 44.055 ;
        RECT 64.595 43.385 64.925 43.885 ;
        RECT 65.095 43.555 65.280 45.675 ;
        RECT 65.535 45.475 65.785 45.935 ;
        RECT 65.955 45.485 66.290 45.655 ;
        RECT 66.485 45.485 67.160 45.655 ;
        RECT 65.955 45.345 66.125 45.485 ;
        RECT 65.450 44.355 65.730 45.305 ;
        RECT 65.900 45.215 66.125 45.345 ;
        RECT 65.900 44.110 66.070 45.215 ;
        RECT 66.295 45.065 66.820 45.285 ;
        RECT 66.240 44.300 66.480 44.895 ;
        RECT 66.650 44.365 66.820 45.065 ;
        RECT 66.990 44.705 67.160 45.485 ;
        RECT 67.480 45.435 67.850 45.935 ;
        RECT 68.030 45.485 68.435 45.655 ;
        RECT 68.605 45.485 69.390 45.655 ;
        RECT 68.030 45.255 68.200 45.485 ;
        RECT 67.370 44.955 68.200 45.255 ;
        RECT 68.585 44.985 69.050 45.315 ;
        RECT 67.370 44.925 67.570 44.955 ;
        RECT 67.690 44.705 67.860 44.775 ;
        RECT 66.990 44.535 67.860 44.705 ;
        RECT 67.350 44.445 67.860 44.535 ;
        RECT 65.900 43.980 66.205 44.110 ;
        RECT 66.650 44.000 67.180 44.365 ;
        RECT 65.520 43.385 65.785 43.845 ;
        RECT 65.955 43.555 66.205 43.980 ;
        RECT 67.350 43.830 67.520 44.445 ;
        RECT 66.415 43.660 67.520 43.830 ;
        RECT 67.690 43.385 67.860 44.185 ;
        RECT 68.030 43.885 68.200 44.955 ;
        RECT 68.370 44.055 68.560 44.775 ;
        RECT 68.730 44.025 69.050 44.985 ;
        RECT 69.220 45.025 69.390 45.485 ;
        RECT 69.665 45.405 69.875 45.935 ;
        RECT 70.135 45.195 70.465 45.720 ;
        RECT 70.635 45.325 70.805 45.935 ;
        RECT 70.975 45.280 71.305 45.715 ;
        RECT 71.475 45.420 71.645 45.935 ;
        RECT 72.075 45.385 72.245 45.675 ;
        RECT 72.415 45.555 72.745 45.935 ;
        RECT 70.975 45.195 71.355 45.280 ;
        RECT 72.075 45.215 72.740 45.385 ;
        RECT 70.265 45.025 70.465 45.195 ;
        RECT 71.130 45.155 71.355 45.195 ;
        RECT 69.220 44.695 70.095 45.025 ;
        RECT 70.265 44.695 71.015 45.025 ;
        RECT 68.030 43.555 68.280 43.885 ;
        RECT 69.220 43.855 69.390 44.695 ;
        RECT 70.265 44.490 70.455 44.695 ;
        RECT 71.185 44.575 71.355 45.155 ;
        RECT 71.140 44.525 71.355 44.575 ;
        RECT 69.560 44.115 70.455 44.490 ;
        RECT 70.965 44.445 71.355 44.525 ;
        RECT 68.505 43.685 69.390 43.855 ;
        RECT 69.570 43.385 69.885 43.885 ;
        RECT 70.115 43.555 70.455 44.115 ;
        RECT 70.625 43.385 70.795 44.395 ;
        RECT 70.965 43.600 71.295 44.445 ;
        RECT 71.990 44.395 72.340 45.045 ;
        RECT 71.465 43.385 71.635 44.300 ;
        RECT 72.510 44.225 72.740 45.215 ;
        RECT 72.075 44.055 72.740 44.225 ;
        RECT 72.075 43.555 72.245 44.055 ;
        RECT 72.415 43.385 72.745 43.885 ;
        RECT 72.915 43.555 73.100 45.675 ;
        RECT 73.355 45.475 73.605 45.935 ;
        RECT 73.775 45.485 74.110 45.655 ;
        RECT 74.305 45.485 74.980 45.655 ;
        RECT 73.775 45.345 73.945 45.485 ;
        RECT 73.270 44.355 73.550 45.305 ;
        RECT 73.720 45.215 73.945 45.345 ;
        RECT 73.720 44.110 73.890 45.215 ;
        RECT 74.115 45.065 74.640 45.285 ;
        RECT 74.060 44.300 74.300 44.895 ;
        RECT 74.470 44.365 74.640 45.065 ;
        RECT 74.810 44.705 74.980 45.485 ;
        RECT 75.300 45.435 75.670 45.935 ;
        RECT 75.850 45.485 76.255 45.655 ;
        RECT 76.425 45.485 77.210 45.655 ;
        RECT 75.850 45.255 76.020 45.485 ;
        RECT 75.190 44.955 76.020 45.255 ;
        RECT 76.405 44.985 76.870 45.315 ;
        RECT 75.190 44.925 75.390 44.955 ;
        RECT 75.510 44.705 75.680 44.775 ;
        RECT 74.810 44.535 75.680 44.705 ;
        RECT 75.170 44.445 75.680 44.535 ;
        RECT 73.720 43.980 74.025 44.110 ;
        RECT 74.470 44.000 75.000 44.365 ;
        RECT 73.340 43.385 73.605 43.845 ;
        RECT 73.775 43.555 74.025 43.980 ;
        RECT 75.170 43.830 75.340 44.445 ;
        RECT 74.235 43.660 75.340 43.830 ;
        RECT 75.510 43.385 75.680 44.185 ;
        RECT 75.850 43.885 76.020 44.955 ;
        RECT 76.190 44.055 76.380 44.775 ;
        RECT 76.550 44.025 76.870 44.985 ;
        RECT 77.040 45.025 77.210 45.485 ;
        RECT 77.485 45.405 77.695 45.935 ;
        RECT 77.955 45.195 78.285 45.720 ;
        RECT 78.455 45.325 78.625 45.935 ;
        RECT 78.795 45.280 79.125 45.715 ;
        RECT 79.395 45.280 79.725 45.715 ;
        RECT 79.895 45.325 80.065 45.935 ;
        RECT 78.795 45.195 79.175 45.280 ;
        RECT 78.085 45.025 78.285 45.195 ;
        RECT 78.950 45.155 79.175 45.195 ;
        RECT 77.040 44.695 77.915 45.025 ;
        RECT 78.085 44.695 78.835 45.025 ;
        RECT 75.850 43.555 76.100 43.885 ;
        RECT 77.040 43.855 77.210 44.695 ;
        RECT 78.085 44.490 78.275 44.695 ;
        RECT 79.005 44.575 79.175 45.155 ;
        RECT 78.960 44.525 79.175 44.575 ;
        RECT 77.380 44.115 78.275 44.490 ;
        RECT 78.785 44.445 79.175 44.525 ;
        RECT 79.345 45.195 79.725 45.280 ;
        RECT 80.235 45.195 80.565 45.720 ;
        RECT 80.825 45.405 81.035 45.935 ;
        RECT 81.310 45.485 82.095 45.655 ;
        RECT 82.265 45.485 82.670 45.655 ;
        RECT 79.345 45.155 79.570 45.195 ;
        RECT 79.345 44.575 79.515 45.155 ;
        RECT 80.235 45.025 80.435 45.195 ;
        RECT 81.310 45.025 81.480 45.485 ;
        RECT 79.685 44.695 80.435 45.025 ;
        RECT 80.605 44.695 81.480 45.025 ;
        RECT 79.345 44.525 79.560 44.575 ;
        RECT 79.345 44.445 79.735 44.525 ;
        RECT 76.325 43.685 77.210 43.855 ;
        RECT 77.390 43.385 77.705 43.885 ;
        RECT 77.935 43.555 78.275 44.115 ;
        RECT 78.445 43.385 78.615 44.395 ;
        RECT 78.785 43.600 79.115 44.445 ;
        RECT 79.405 43.600 79.735 44.445 ;
        RECT 80.245 44.490 80.435 44.695 ;
        RECT 79.905 43.385 80.075 44.395 ;
        RECT 80.245 44.115 81.140 44.490 ;
        RECT 80.245 43.555 80.585 44.115 ;
        RECT 80.815 43.385 81.130 43.885 ;
        RECT 81.310 43.855 81.480 44.695 ;
        RECT 81.650 44.985 82.115 45.315 ;
        RECT 82.500 45.255 82.670 45.485 ;
        RECT 82.850 45.435 83.220 45.935 ;
        RECT 83.540 45.485 84.215 45.655 ;
        RECT 84.410 45.485 84.745 45.655 ;
        RECT 81.650 44.025 81.970 44.985 ;
        RECT 82.500 44.955 83.330 45.255 ;
        RECT 82.140 44.055 82.330 44.775 ;
        RECT 82.500 43.885 82.670 44.955 ;
        RECT 83.130 44.925 83.330 44.955 ;
        RECT 82.840 44.705 83.010 44.775 ;
        RECT 83.540 44.705 83.710 45.485 ;
        RECT 84.575 45.345 84.745 45.485 ;
        RECT 84.915 45.475 85.165 45.935 ;
        RECT 82.840 44.535 83.710 44.705 ;
        RECT 83.880 45.065 84.405 45.285 ;
        RECT 84.575 45.215 84.800 45.345 ;
        RECT 82.840 44.445 83.350 44.535 ;
        RECT 81.310 43.685 82.195 43.855 ;
        RECT 82.420 43.555 82.670 43.885 ;
        RECT 82.840 43.385 83.010 44.185 ;
        RECT 83.180 43.830 83.350 44.445 ;
        RECT 83.880 44.365 84.050 45.065 ;
        RECT 83.520 44.000 84.050 44.365 ;
        RECT 84.220 44.300 84.460 44.895 ;
        RECT 84.630 44.110 84.800 45.215 ;
        RECT 84.970 44.355 85.250 45.305 ;
        RECT 84.495 43.980 84.800 44.110 ;
        RECT 83.180 43.660 84.285 43.830 ;
        RECT 84.495 43.555 84.745 43.980 ;
        RECT 84.915 43.385 85.180 43.845 ;
        RECT 85.420 43.555 85.605 45.675 ;
        RECT 85.775 45.555 86.105 45.935 ;
        RECT 86.275 45.385 86.445 45.675 ;
        RECT 85.780 45.215 86.445 45.385 ;
        RECT 86.795 45.385 86.965 45.765 ;
        RECT 87.180 45.555 87.510 45.935 ;
        RECT 86.795 45.215 87.510 45.385 ;
        RECT 85.780 44.225 86.010 45.215 ;
        RECT 86.180 44.395 86.530 45.045 ;
        RECT 86.705 44.665 87.060 45.035 ;
        RECT 87.340 45.025 87.510 45.215 ;
        RECT 87.680 45.190 87.935 45.765 ;
        RECT 87.340 44.695 87.595 45.025 ;
        RECT 87.340 44.485 87.510 44.695 ;
        RECT 86.795 44.315 87.510 44.485 ;
        RECT 87.765 44.460 87.935 45.190 ;
        RECT 88.110 45.095 88.370 45.935 ;
        RECT 88.545 45.185 89.755 45.935 ;
        RECT 85.780 44.055 86.445 44.225 ;
        RECT 85.775 43.385 86.105 43.885 ;
        RECT 86.275 43.555 86.445 44.055 ;
        RECT 86.795 43.555 86.965 44.315 ;
        RECT 87.180 43.385 87.510 44.145 ;
        RECT 87.680 43.555 87.935 44.460 ;
        RECT 88.110 43.385 88.370 44.535 ;
        RECT 88.545 44.475 89.065 45.015 ;
        RECT 89.235 44.645 89.755 45.185 ;
        RECT 88.545 43.385 89.755 44.475 ;
        RECT 12.100 43.215 89.840 43.385 ;
        RECT 12.185 42.125 13.395 43.215 ;
        RECT 12.185 41.415 12.705 41.955 ;
        RECT 12.875 41.585 13.395 42.125 ;
        RECT 14.025 42.365 14.405 43.045 ;
        RECT 14.995 42.365 15.165 43.215 ;
        RECT 15.335 42.535 15.665 43.045 ;
        RECT 15.835 42.705 16.005 43.215 ;
        RECT 16.175 42.535 16.575 43.045 ;
        RECT 15.335 42.365 16.575 42.535 ;
        RECT 12.185 40.665 13.395 41.415 ;
        RECT 14.025 41.405 14.195 42.365 ;
        RECT 14.365 42.025 15.670 42.195 ;
        RECT 16.755 42.115 17.075 43.045 ;
        RECT 17.245 42.660 17.850 43.215 ;
        RECT 18.025 42.705 18.505 43.045 ;
        RECT 18.675 42.670 18.930 43.215 ;
        RECT 17.245 42.560 17.860 42.660 ;
        RECT 17.675 42.535 17.860 42.560 ;
        RECT 14.365 41.575 14.610 42.025 ;
        RECT 14.780 41.655 15.330 41.855 ;
        RECT 15.500 41.825 15.670 42.025 ;
        RECT 16.445 41.945 17.075 42.115 ;
        RECT 15.500 41.655 15.875 41.825 ;
        RECT 16.045 41.405 16.275 41.905 ;
        RECT 14.025 41.235 16.275 41.405 ;
        RECT 14.075 40.665 14.405 41.055 ;
        RECT 14.575 40.915 14.745 41.235 ;
        RECT 16.445 41.065 16.615 41.945 ;
        RECT 17.245 41.940 17.505 42.390 ;
        RECT 17.675 42.290 18.005 42.535 ;
        RECT 18.175 42.215 18.930 42.465 ;
        RECT 19.100 42.345 19.375 43.045 ;
        RECT 20.465 42.660 21.070 43.215 ;
        RECT 21.245 42.705 21.725 43.045 ;
        RECT 21.895 42.670 22.150 43.215 ;
        RECT 20.465 42.560 21.080 42.660 ;
        RECT 20.895 42.535 21.080 42.560 ;
        RECT 18.160 42.180 18.930 42.215 ;
        RECT 18.145 42.170 18.930 42.180 ;
        RECT 18.140 42.155 19.035 42.170 ;
        RECT 18.120 42.140 19.035 42.155 ;
        RECT 18.100 42.130 19.035 42.140 ;
        RECT 18.075 42.120 19.035 42.130 ;
        RECT 18.005 42.090 19.035 42.120 ;
        RECT 17.985 42.060 19.035 42.090 ;
        RECT 17.965 42.030 19.035 42.060 ;
        RECT 17.935 42.005 19.035 42.030 ;
        RECT 17.900 41.970 19.035 42.005 ;
        RECT 17.870 41.965 19.035 41.970 ;
        RECT 17.870 41.960 18.260 41.965 ;
        RECT 17.870 41.950 18.235 41.960 ;
        RECT 17.870 41.945 18.220 41.950 ;
        RECT 17.870 41.940 18.205 41.945 ;
        RECT 17.245 41.935 18.205 41.940 ;
        RECT 17.245 41.925 18.195 41.935 ;
        RECT 17.245 41.920 18.185 41.925 ;
        RECT 17.245 41.910 18.175 41.920 ;
        RECT 17.245 41.900 18.170 41.910 ;
        RECT 17.245 41.895 18.165 41.900 ;
        RECT 17.245 41.880 18.155 41.895 ;
        RECT 17.245 41.865 18.150 41.880 ;
        RECT 17.245 41.840 18.140 41.865 ;
        RECT 17.245 41.770 18.135 41.840 ;
        RECT 14.915 40.665 15.245 41.055 ;
        RECT 15.660 40.895 16.615 41.065 ;
        RECT 16.785 40.665 17.075 41.500 ;
        RECT 17.245 41.215 17.795 41.600 ;
        RECT 17.965 41.045 18.135 41.770 ;
        RECT 17.245 40.875 18.135 41.045 ;
        RECT 18.305 41.370 18.635 41.795 ;
        RECT 18.805 41.570 19.035 41.965 ;
        RECT 18.305 40.885 18.525 41.370 ;
        RECT 19.205 41.315 19.375 42.345 ;
        RECT 20.465 41.940 20.725 42.390 ;
        RECT 20.895 42.290 21.225 42.535 ;
        RECT 21.395 42.215 22.150 42.465 ;
        RECT 22.320 42.345 22.595 43.045 ;
        RECT 22.765 42.660 23.370 43.215 ;
        RECT 23.545 42.705 24.025 43.045 ;
        RECT 24.195 42.670 24.450 43.215 ;
        RECT 22.765 42.560 23.380 42.660 ;
        RECT 23.195 42.535 23.380 42.560 ;
        RECT 21.380 42.180 22.150 42.215 ;
        RECT 21.365 42.170 22.150 42.180 ;
        RECT 21.360 42.155 22.255 42.170 ;
        RECT 21.340 42.140 22.255 42.155 ;
        RECT 21.320 42.130 22.255 42.140 ;
        RECT 21.295 42.120 22.255 42.130 ;
        RECT 21.225 42.090 22.255 42.120 ;
        RECT 21.205 42.060 22.255 42.090 ;
        RECT 21.185 42.030 22.255 42.060 ;
        RECT 21.155 42.005 22.255 42.030 ;
        RECT 21.120 41.970 22.255 42.005 ;
        RECT 21.090 41.965 22.255 41.970 ;
        RECT 21.090 41.960 21.480 41.965 ;
        RECT 21.090 41.950 21.455 41.960 ;
        RECT 21.090 41.945 21.440 41.950 ;
        RECT 21.090 41.940 21.425 41.945 ;
        RECT 20.465 41.935 21.425 41.940 ;
        RECT 20.465 41.925 21.415 41.935 ;
        RECT 20.465 41.920 21.405 41.925 ;
        RECT 20.465 41.910 21.395 41.920 ;
        RECT 20.465 41.900 21.390 41.910 ;
        RECT 20.465 41.895 21.385 41.900 ;
        RECT 20.465 41.880 21.375 41.895 ;
        RECT 20.465 41.865 21.370 41.880 ;
        RECT 20.465 41.840 21.360 41.865 ;
        RECT 20.465 41.770 21.355 41.840 ;
        RECT 18.695 40.665 18.945 41.205 ;
        RECT 19.115 40.835 19.375 41.315 ;
        RECT 20.465 41.215 21.015 41.600 ;
        RECT 21.185 41.045 21.355 41.770 ;
        RECT 20.465 40.875 21.355 41.045 ;
        RECT 21.525 41.370 21.855 41.795 ;
        RECT 22.025 41.570 22.255 41.965 ;
        RECT 21.525 40.885 21.745 41.370 ;
        RECT 22.425 41.315 22.595 42.345 ;
        RECT 22.765 41.940 23.025 42.390 ;
        RECT 23.195 42.290 23.525 42.535 ;
        RECT 23.695 42.215 24.450 42.465 ;
        RECT 24.620 42.345 24.895 43.045 ;
        RECT 23.680 42.180 24.450 42.215 ;
        RECT 23.665 42.170 24.450 42.180 ;
        RECT 23.660 42.155 24.555 42.170 ;
        RECT 23.640 42.140 24.555 42.155 ;
        RECT 23.620 42.130 24.555 42.140 ;
        RECT 23.595 42.120 24.555 42.130 ;
        RECT 23.525 42.090 24.555 42.120 ;
        RECT 23.505 42.060 24.555 42.090 ;
        RECT 23.485 42.030 24.555 42.060 ;
        RECT 23.455 42.005 24.555 42.030 ;
        RECT 23.420 41.970 24.555 42.005 ;
        RECT 23.390 41.965 24.555 41.970 ;
        RECT 23.390 41.960 23.780 41.965 ;
        RECT 23.390 41.950 23.755 41.960 ;
        RECT 23.390 41.945 23.740 41.950 ;
        RECT 23.390 41.940 23.725 41.945 ;
        RECT 22.765 41.935 23.725 41.940 ;
        RECT 22.765 41.925 23.715 41.935 ;
        RECT 22.765 41.920 23.705 41.925 ;
        RECT 22.765 41.910 23.695 41.920 ;
        RECT 22.765 41.900 23.690 41.910 ;
        RECT 22.765 41.895 23.685 41.900 ;
        RECT 22.765 41.880 23.675 41.895 ;
        RECT 22.765 41.865 23.670 41.880 ;
        RECT 22.765 41.840 23.660 41.865 ;
        RECT 22.765 41.770 23.655 41.840 ;
        RECT 21.915 40.665 22.165 41.205 ;
        RECT 22.335 40.835 22.595 41.315 ;
        RECT 22.765 41.215 23.315 41.600 ;
        RECT 23.485 41.045 23.655 41.770 ;
        RECT 22.765 40.875 23.655 41.045 ;
        RECT 23.825 41.370 24.155 41.795 ;
        RECT 24.325 41.570 24.555 41.965 ;
        RECT 23.825 40.885 24.045 41.370 ;
        RECT 24.725 41.315 24.895 42.345 ;
        RECT 25.065 42.050 25.355 43.215 ;
        RECT 25.615 42.545 25.785 43.045 ;
        RECT 25.955 42.715 26.285 43.215 ;
        RECT 25.615 42.375 26.280 42.545 ;
        RECT 25.530 41.555 25.880 42.205 ;
        RECT 24.215 40.665 24.465 41.205 ;
        RECT 24.635 40.835 24.895 41.315 ;
        RECT 25.065 40.665 25.355 41.390 ;
        RECT 26.050 41.385 26.280 42.375 ;
        RECT 25.615 41.215 26.280 41.385 ;
        RECT 25.615 40.925 25.785 41.215 ;
        RECT 25.955 40.665 26.285 41.045 ;
        RECT 26.455 40.925 26.640 43.045 ;
        RECT 26.880 42.755 27.145 43.215 ;
        RECT 27.315 42.620 27.565 43.045 ;
        RECT 27.775 42.770 28.880 42.940 ;
        RECT 27.260 42.490 27.565 42.620 ;
        RECT 26.810 41.295 27.090 42.245 ;
        RECT 27.260 41.385 27.430 42.490 ;
        RECT 27.600 41.705 27.840 42.300 ;
        RECT 28.010 42.235 28.540 42.600 ;
        RECT 28.010 41.535 28.180 42.235 ;
        RECT 28.710 42.155 28.880 42.770 ;
        RECT 29.050 42.415 29.220 43.215 ;
        RECT 29.390 42.715 29.640 43.045 ;
        RECT 29.865 42.745 30.750 42.915 ;
        RECT 28.710 42.065 29.220 42.155 ;
        RECT 27.260 41.255 27.485 41.385 ;
        RECT 27.655 41.315 28.180 41.535 ;
        RECT 28.350 41.895 29.220 42.065 ;
        RECT 26.895 40.665 27.145 41.125 ;
        RECT 27.315 41.115 27.485 41.255 ;
        RECT 28.350 41.115 28.520 41.895 ;
        RECT 29.050 41.825 29.220 41.895 ;
        RECT 28.730 41.645 28.930 41.675 ;
        RECT 29.390 41.645 29.560 42.715 ;
        RECT 29.730 41.825 29.920 42.545 ;
        RECT 28.730 41.345 29.560 41.645 ;
        RECT 30.090 41.615 30.410 42.575 ;
        RECT 27.315 40.945 27.650 41.115 ;
        RECT 27.845 40.945 28.520 41.115 ;
        RECT 28.840 40.665 29.210 41.165 ;
        RECT 29.390 41.115 29.560 41.345 ;
        RECT 29.945 41.285 30.410 41.615 ;
        RECT 30.580 41.905 30.750 42.745 ;
        RECT 30.930 42.715 31.245 43.215 ;
        RECT 31.475 42.485 31.815 43.045 ;
        RECT 30.920 42.110 31.815 42.485 ;
        RECT 31.985 42.205 32.155 43.215 ;
        RECT 31.625 41.905 31.815 42.110 ;
        RECT 32.325 42.155 32.655 43.000 ;
        RECT 32.895 42.245 33.225 43.030 ;
        RECT 32.325 42.075 32.715 42.155 ;
        RECT 32.895 42.075 33.575 42.245 ;
        RECT 33.755 42.075 34.085 43.215 ;
        RECT 34.355 42.545 34.525 43.045 ;
        RECT 34.695 42.715 35.025 43.215 ;
        RECT 34.355 42.375 35.020 42.545 ;
        RECT 32.500 42.025 32.715 42.075 ;
        RECT 30.580 41.575 31.455 41.905 ;
        RECT 31.625 41.575 32.375 41.905 ;
        RECT 30.580 41.115 30.750 41.575 ;
        RECT 31.625 41.405 31.825 41.575 ;
        RECT 32.545 41.445 32.715 42.025 ;
        RECT 32.885 41.655 33.235 41.905 ;
        RECT 33.405 41.475 33.575 42.075 ;
        RECT 33.745 41.655 34.095 41.905 ;
        RECT 34.270 41.555 34.620 42.205 ;
        RECT 32.490 41.405 32.715 41.445 ;
        RECT 29.390 40.945 29.795 41.115 ;
        RECT 29.965 40.945 30.750 41.115 ;
        RECT 31.025 40.665 31.235 41.195 ;
        RECT 31.495 40.880 31.825 41.405 ;
        RECT 32.335 41.320 32.715 41.405 ;
        RECT 31.995 40.665 32.165 41.275 ;
        RECT 32.335 40.885 32.665 41.320 ;
        RECT 32.905 40.665 33.145 41.475 ;
        RECT 33.315 40.835 33.645 41.475 ;
        RECT 33.815 40.665 34.085 41.475 ;
        RECT 34.790 41.385 35.020 42.375 ;
        RECT 34.355 41.215 35.020 41.385 ;
        RECT 34.355 40.925 34.525 41.215 ;
        RECT 34.695 40.665 35.025 41.045 ;
        RECT 35.195 40.925 35.380 43.045 ;
        RECT 35.620 42.755 35.885 43.215 ;
        RECT 36.055 42.620 36.305 43.045 ;
        RECT 36.515 42.770 37.620 42.940 ;
        RECT 36.000 42.490 36.305 42.620 ;
        RECT 35.550 41.295 35.830 42.245 ;
        RECT 36.000 41.385 36.170 42.490 ;
        RECT 36.340 41.705 36.580 42.300 ;
        RECT 36.750 42.235 37.280 42.600 ;
        RECT 36.750 41.535 36.920 42.235 ;
        RECT 37.450 42.155 37.620 42.770 ;
        RECT 37.790 42.415 37.960 43.215 ;
        RECT 38.130 42.715 38.380 43.045 ;
        RECT 38.605 42.745 39.490 42.915 ;
        RECT 37.450 42.065 37.960 42.155 ;
        RECT 36.000 41.255 36.225 41.385 ;
        RECT 36.395 41.315 36.920 41.535 ;
        RECT 37.090 41.895 37.960 42.065 ;
        RECT 35.635 40.665 35.885 41.125 ;
        RECT 36.055 41.115 36.225 41.255 ;
        RECT 37.090 41.115 37.260 41.895 ;
        RECT 37.790 41.825 37.960 41.895 ;
        RECT 37.470 41.645 37.670 41.675 ;
        RECT 38.130 41.645 38.300 42.715 ;
        RECT 38.470 41.825 38.660 42.545 ;
        RECT 37.470 41.345 38.300 41.645 ;
        RECT 38.830 41.615 39.150 42.575 ;
        RECT 36.055 40.945 36.390 41.115 ;
        RECT 36.585 40.945 37.260 41.115 ;
        RECT 37.580 40.665 37.950 41.165 ;
        RECT 38.130 41.115 38.300 41.345 ;
        RECT 38.685 41.285 39.150 41.615 ;
        RECT 39.320 41.905 39.490 42.745 ;
        RECT 39.670 42.715 39.985 43.215 ;
        RECT 40.215 42.485 40.555 43.045 ;
        RECT 39.660 42.110 40.555 42.485 ;
        RECT 40.725 42.205 40.895 43.215 ;
        RECT 40.365 41.905 40.555 42.110 ;
        RECT 41.065 42.155 41.395 43.000 ;
        RECT 41.625 42.345 41.900 43.045 ;
        RECT 42.070 42.670 42.325 43.215 ;
        RECT 42.495 42.705 42.975 43.045 ;
        RECT 43.150 42.660 43.755 43.215 ;
        RECT 43.140 42.560 43.755 42.660 ;
        RECT 43.140 42.535 43.325 42.560 ;
        RECT 41.065 42.075 41.455 42.155 ;
        RECT 41.240 42.025 41.455 42.075 ;
        RECT 39.320 41.575 40.195 41.905 ;
        RECT 40.365 41.575 41.115 41.905 ;
        RECT 39.320 41.115 39.490 41.575 ;
        RECT 40.365 41.405 40.565 41.575 ;
        RECT 41.285 41.445 41.455 42.025 ;
        RECT 41.230 41.405 41.455 41.445 ;
        RECT 38.130 40.945 38.535 41.115 ;
        RECT 38.705 40.945 39.490 41.115 ;
        RECT 39.765 40.665 39.975 41.195 ;
        RECT 40.235 40.880 40.565 41.405 ;
        RECT 41.075 41.320 41.455 41.405 ;
        RECT 40.735 40.665 40.905 41.275 ;
        RECT 41.075 40.885 41.405 41.320 ;
        RECT 41.625 41.315 41.795 42.345 ;
        RECT 42.070 42.215 42.825 42.465 ;
        RECT 42.995 42.290 43.325 42.535 ;
        RECT 42.070 42.180 42.840 42.215 ;
        RECT 42.070 42.170 42.855 42.180 ;
        RECT 41.965 42.155 42.860 42.170 ;
        RECT 41.965 42.140 42.880 42.155 ;
        RECT 41.965 42.130 42.900 42.140 ;
        RECT 41.965 42.120 42.925 42.130 ;
        RECT 41.965 42.090 42.995 42.120 ;
        RECT 41.965 42.060 43.015 42.090 ;
        RECT 41.965 42.030 43.035 42.060 ;
        RECT 41.965 42.005 43.065 42.030 ;
        RECT 41.965 41.970 43.100 42.005 ;
        RECT 41.965 41.965 43.130 41.970 ;
        RECT 41.965 41.570 42.195 41.965 ;
        RECT 42.740 41.960 43.130 41.965 ;
        RECT 42.765 41.950 43.130 41.960 ;
        RECT 42.780 41.945 43.130 41.950 ;
        RECT 42.795 41.940 43.130 41.945 ;
        RECT 43.495 41.940 43.755 42.390 ;
        RECT 43.925 42.125 45.595 43.215 ;
        RECT 42.795 41.935 43.755 41.940 ;
        RECT 42.805 41.925 43.755 41.935 ;
        RECT 42.815 41.920 43.755 41.925 ;
        RECT 42.825 41.910 43.755 41.920 ;
        RECT 42.830 41.900 43.755 41.910 ;
        RECT 42.835 41.895 43.755 41.900 ;
        RECT 42.845 41.880 43.755 41.895 ;
        RECT 42.850 41.865 43.755 41.880 ;
        RECT 42.860 41.840 43.755 41.865 ;
        RECT 42.365 41.370 42.695 41.795 ;
        RECT 42.445 41.345 42.695 41.370 ;
        RECT 41.625 40.835 41.885 41.315 ;
        RECT 42.055 40.665 42.305 41.205 ;
        RECT 42.475 40.885 42.695 41.345 ;
        RECT 42.865 41.770 43.755 41.840 ;
        RECT 42.865 41.045 43.035 41.770 ;
        RECT 43.205 41.215 43.755 41.600 ;
        RECT 43.925 41.435 44.675 41.955 ;
        RECT 44.845 41.605 45.595 42.125 ;
        RECT 45.765 42.075 46.025 43.215 ;
        RECT 46.195 42.065 46.525 43.045 ;
        RECT 46.695 42.075 46.975 43.215 ;
        RECT 47.145 42.125 50.655 43.215 ;
        RECT 45.785 41.655 46.120 41.905 ;
        RECT 46.290 41.515 46.460 42.065 ;
        RECT 46.630 41.635 46.965 41.905 ;
        RECT 46.285 41.465 46.460 41.515 ;
        RECT 42.865 40.875 43.755 41.045 ;
        RECT 43.925 40.665 45.595 41.435 ;
        RECT 45.765 40.835 46.460 41.465 ;
        RECT 46.665 40.665 46.975 41.465 ;
        RECT 47.145 41.435 48.795 41.955 ;
        RECT 48.965 41.605 50.655 42.125 ;
        RECT 50.825 42.050 51.115 43.215 ;
        RECT 51.285 42.125 52.495 43.215 ;
        RECT 47.145 40.665 50.655 41.435 ;
        RECT 51.285 41.415 51.805 41.955 ;
        RECT 51.975 41.585 52.495 42.125 ;
        RECT 52.665 42.075 53.050 43.045 ;
        RECT 53.220 42.755 53.545 43.215 ;
        RECT 54.065 42.585 54.345 43.045 ;
        RECT 53.220 42.365 54.345 42.585 ;
        RECT 50.825 40.665 51.115 41.390 ;
        RECT 51.285 40.665 52.495 41.415 ;
        RECT 52.665 41.405 52.945 42.075 ;
        RECT 53.220 41.905 53.670 42.365 ;
        RECT 54.535 42.195 54.935 43.045 ;
        RECT 55.335 42.755 55.605 43.215 ;
        RECT 55.775 42.585 56.060 43.045 ;
        RECT 53.115 41.575 53.670 41.905 ;
        RECT 53.840 41.635 54.935 42.195 ;
        RECT 53.220 41.465 53.670 41.575 ;
        RECT 52.665 40.835 53.050 41.405 ;
        RECT 53.220 41.295 54.345 41.465 ;
        RECT 53.220 40.665 53.545 41.125 ;
        RECT 54.065 40.835 54.345 41.295 ;
        RECT 54.535 40.835 54.935 41.635 ;
        RECT 55.105 42.365 56.060 42.585 ;
        RECT 55.105 41.465 55.315 42.365 ;
        RECT 55.485 41.635 56.175 42.195 ;
        RECT 56.345 42.075 56.730 43.045 ;
        RECT 56.900 42.755 57.225 43.215 ;
        RECT 57.745 42.585 58.025 43.045 ;
        RECT 56.900 42.365 58.025 42.585 ;
        RECT 55.105 41.295 56.060 41.465 ;
        RECT 55.335 40.665 55.605 41.125 ;
        RECT 55.775 40.835 56.060 41.295 ;
        RECT 56.345 41.405 56.625 42.075 ;
        RECT 56.900 41.905 57.350 42.365 ;
        RECT 58.215 42.195 58.615 43.045 ;
        RECT 59.015 42.755 59.285 43.215 ;
        RECT 59.455 42.585 59.740 43.045 ;
        RECT 56.795 41.575 57.350 41.905 ;
        RECT 57.520 41.635 58.615 42.195 ;
        RECT 56.900 41.465 57.350 41.575 ;
        RECT 56.345 40.835 56.730 41.405 ;
        RECT 56.900 41.295 58.025 41.465 ;
        RECT 56.900 40.665 57.225 41.125 ;
        RECT 57.745 40.835 58.025 41.295 ;
        RECT 58.215 40.835 58.615 41.635 ;
        RECT 58.785 42.365 59.740 42.585 ;
        RECT 60.110 42.595 60.285 43.045 ;
        RECT 60.455 42.775 60.785 43.215 ;
        RECT 61.090 42.625 61.260 43.045 ;
        RECT 61.495 42.805 62.165 43.215 ;
        RECT 62.380 42.625 62.550 43.045 ;
        RECT 62.750 42.805 63.080 43.215 ;
        RECT 60.110 42.425 60.740 42.595 ;
        RECT 58.785 41.465 58.995 42.365 ;
        RECT 59.165 41.635 59.855 42.195 ;
        RECT 60.025 41.575 60.390 42.255 ;
        RECT 60.570 41.905 60.740 42.425 ;
        RECT 61.090 42.455 63.105 42.625 ;
        RECT 60.570 41.575 60.920 41.905 ;
        RECT 58.785 41.295 59.740 41.465 ;
        RECT 60.570 41.405 60.740 41.575 ;
        RECT 59.015 40.665 59.285 41.125 ;
        RECT 59.455 40.835 59.740 41.295 ;
        RECT 60.110 41.235 60.740 41.405 ;
        RECT 60.110 40.835 60.285 41.235 ;
        RECT 61.090 41.165 61.260 42.455 ;
        RECT 60.455 40.665 60.785 41.045 ;
        RECT 61.030 40.835 61.260 41.165 ;
        RECT 61.460 41.000 61.740 42.275 ;
        RECT 61.965 41.515 62.235 42.275 ;
        RECT 61.925 41.345 62.235 41.515 ;
        RECT 61.965 41.000 62.235 41.345 ;
        RECT 62.425 41.245 62.765 42.275 ;
        RECT 62.935 41.905 63.105 42.455 ;
        RECT 63.275 42.075 63.535 43.045 ;
        RECT 62.935 41.575 63.195 41.905 ;
        RECT 63.365 41.385 63.535 42.075 ;
        RECT 62.695 40.665 63.025 41.045 ;
        RECT 63.195 40.920 63.535 41.385 ;
        RECT 64.170 42.075 64.505 43.045 ;
        RECT 64.675 42.075 64.845 43.215 ;
        RECT 65.015 42.875 67.045 43.045 ;
        RECT 64.170 41.405 64.340 42.075 ;
        RECT 65.015 41.905 65.185 42.875 ;
        RECT 64.510 41.575 64.765 41.905 ;
        RECT 64.990 41.575 65.185 41.905 ;
        RECT 65.355 42.535 66.480 42.705 ;
        RECT 64.595 41.405 64.765 41.575 ;
        RECT 65.355 41.405 65.525 42.535 ;
        RECT 63.195 40.875 63.530 40.920 ;
        RECT 64.170 40.835 64.425 41.405 ;
        RECT 64.595 41.235 65.525 41.405 ;
        RECT 65.695 42.195 66.705 42.365 ;
        RECT 65.695 41.395 65.865 42.195 ;
        RECT 65.350 41.200 65.525 41.235 ;
        RECT 64.595 40.665 64.925 41.065 ;
        RECT 65.350 40.835 65.880 41.200 ;
        RECT 66.070 41.175 66.345 41.995 ;
        RECT 66.065 41.005 66.345 41.175 ;
        RECT 66.070 40.835 66.345 41.005 ;
        RECT 66.515 40.835 66.705 42.195 ;
        RECT 66.875 42.210 67.045 42.875 ;
        RECT 67.215 42.455 67.385 43.215 ;
        RECT 67.620 42.455 68.135 42.865 ;
        RECT 66.875 42.020 67.625 42.210 ;
        RECT 67.795 41.645 68.135 42.455 ;
        RECT 68.305 42.125 69.515 43.215 ;
        RECT 66.905 41.475 68.135 41.645 ;
        RECT 66.885 40.665 67.395 41.200 ;
        RECT 67.615 40.870 67.860 41.475 ;
        RECT 68.305 41.415 68.825 41.955 ;
        RECT 68.995 41.585 69.515 42.125 ;
        RECT 69.690 42.065 69.950 43.215 ;
        RECT 70.125 42.140 70.380 43.045 ;
        RECT 70.550 42.455 70.880 43.215 ;
        RECT 71.095 42.285 71.265 43.045 ;
        RECT 68.305 40.665 69.515 41.415 ;
        RECT 69.690 40.665 69.950 41.505 ;
        RECT 70.125 41.410 70.295 42.140 ;
        RECT 70.550 42.115 71.265 42.285 ;
        RECT 70.550 41.905 70.720 42.115 ;
        RECT 71.525 42.075 71.865 43.045 ;
        RECT 72.035 42.075 72.205 43.215 ;
        RECT 72.475 42.415 72.725 43.215 ;
        RECT 73.370 42.245 73.700 43.045 ;
        RECT 74.000 42.415 74.330 43.215 ;
        RECT 74.500 42.245 74.830 43.045 ;
        RECT 72.395 42.075 74.830 42.245 ;
        RECT 75.205 42.125 76.415 43.215 ;
        RECT 70.465 41.575 70.720 41.905 ;
        RECT 70.125 40.835 70.380 41.410 ;
        RECT 70.550 41.385 70.720 41.575 ;
        RECT 71.000 41.565 71.355 41.935 ;
        RECT 71.525 41.465 71.700 42.075 ;
        RECT 72.395 41.825 72.565 42.075 ;
        RECT 71.870 41.655 72.565 41.825 ;
        RECT 72.740 41.655 73.160 41.855 ;
        RECT 73.330 41.655 73.660 41.855 ;
        RECT 73.830 41.655 74.160 41.855 ;
        RECT 70.550 41.215 71.265 41.385 ;
        RECT 70.550 40.665 70.880 41.045 ;
        RECT 71.095 40.835 71.265 41.215 ;
        RECT 71.525 40.835 71.865 41.465 ;
        RECT 72.035 40.665 72.285 41.465 ;
        RECT 72.475 41.315 73.700 41.485 ;
        RECT 72.475 40.835 72.805 41.315 ;
        RECT 72.975 40.665 73.200 41.125 ;
        RECT 73.370 40.835 73.700 41.315 ;
        RECT 74.330 41.445 74.500 42.075 ;
        RECT 74.685 41.655 75.035 41.905 ;
        RECT 74.330 40.835 74.830 41.445 ;
        RECT 75.205 41.415 75.725 41.955 ;
        RECT 75.895 41.585 76.415 42.125 ;
        RECT 76.585 42.050 76.875 43.215 ;
        RECT 77.050 42.825 77.385 43.045 ;
        RECT 78.390 42.835 78.745 43.215 ;
        RECT 77.050 42.205 77.305 42.825 ;
        RECT 77.555 42.665 77.785 42.705 ;
        RECT 78.915 42.665 79.165 43.045 ;
        RECT 77.555 42.465 79.165 42.665 ;
        RECT 77.555 42.375 77.740 42.465 ;
        RECT 78.330 42.455 79.165 42.465 ;
        RECT 79.415 42.435 79.665 43.215 ;
        RECT 79.835 42.365 80.095 43.045 ;
        RECT 81.275 42.545 81.445 43.045 ;
        RECT 81.615 42.715 81.945 43.215 ;
        RECT 81.275 42.375 81.940 42.545 ;
        RECT 77.895 42.265 78.225 42.295 ;
        RECT 77.895 42.205 79.695 42.265 ;
        RECT 77.050 42.095 79.755 42.205 ;
        RECT 77.050 42.035 78.225 42.095 ;
        RECT 79.555 42.060 79.755 42.095 ;
        RECT 77.045 41.655 77.535 41.855 ;
        RECT 77.725 41.655 78.200 41.865 ;
        RECT 75.205 40.665 76.415 41.415 ;
        RECT 76.585 40.665 76.875 41.390 ;
        RECT 77.050 40.665 77.505 41.430 ;
        RECT 77.980 41.255 78.200 41.655 ;
        RECT 78.445 41.655 78.775 41.865 ;
        RECT 78.445 41.255 78.655 41.655 ;
        RECT 78.945 41.620 79.355 41.925 ;
        RECT 79.585 41.485 79.755 42.060 ;
        RECT 79.485 41.365 79.755 41.485 ;
        RECT 78.910 41.320 79.755 41.365 ;
        RECT 78.910 41.195 79.665 41.320 ;
        RECT 78.910 41.045 79.080 41.195 ;
        RECT 79.925 41.165 80.095 42.365 ;
        RECT 81.190 41.555 81.540 42.205 ;
        RECT 81.710 41.385 81.940 42.375 ;
        RECT 77.780 40.835 79.080 41.045 ;
        RECT 79.335 40.665 79.665 41.025 ;
        RECT 79.835 40.835 80.095 41.165 ;
        RECT 81.275 41.215 81.940 41.385 ;
        RECT 81.275 40.925 81.445 41.215 ;
        RECT 81.615 40.665 81.945 41.045 ;
        RECT 82.115 40.925 82.300 43.045 ;
        RECT 82.540 42.755 82.805 43.215 ;
        RECT 82.975 42.620 83.225 43.045 ;
        RECT 83.435 42.770 84.540 42.940 ;
        RECT 82.920 42.490 83.225 42.620 ;
        RECT 82.470 41.295 82.750 42.245 ;
        RECT 82.920 41.385 83.090 42.490 ;
        RECT 83.260 41.705 83.500 42.300 ;
        RECT 83.670 42.235 84.200 42.600 ;
        RECT 83.670 41.535 83.840 42.235 ;
        RECT 84.370 42.155 84.540 42.770 ;
        RECT 84.710 42.415 84.880 43.215 ;
        RECT 85.050 42.715 85.300 43.045 ;
        RECT 85.525 42.745 86.410 42.915 ;
        RECT 84.370 42.065 84.880 42.155 ;
        RECT 82.920 41.255 83.145 41.385 ;
        RECT 83.315 41.315 83.840 41.535 ;
        RECT 84.010 41.895 84.880 42.065 ;
        RECT 82.555 40.665 82.805 41.125 ;
        RECT 82.975 41.115 83.145 41.255 ;
        RECT 84.010 41.115 84.180 41.895 ;
        RECT 84.710 41.825 84.880 41.895 ;
        RECT 84.390 41.645 84.590 41.675 ;
        RECT 85.050 41.645 85.220 42.715 ;
        RECT 85.390 41.825 85.580 42.545 ;
        RECT 84.390 41.345 85.220 41.645 ;
        RECT 85.750 41.615 86.070 42.575 ;
        RECT 82.975 40.945 83.310 41.115 ;
        RECT 83.505 40.945 84.180 41.115 ;
        RECT 84.500 40.665 84.870 41.165 ;
        RECT 85.050 41.115 85.220 41.345 ;
        RECT 85.605 41.285 86.070 41.615 ;
        RECT 86.240 41.905 86.410 42.745 ;
        RECT 86.590 42.715 86.905 43.215 ;
        RECT 87.135 42.485 87.475 43.045 ;
        RECT 86.580 42.110 87.475 42.485 ;
        RECT 87.645 42.205 87.815 43.215 ;
        RECT 87.285 41.905 87.475 42.110 ;
        RECT 87.985 42.155 88.315 43.000 ;
        RECT 87.985 42.075 88.375 42.155 ;
        RECT 88.160 42.025 88.375 42.075 ;
        RECT 86.240 41.575 87.115 41.905 ;
        RECT 87.285 41.575 88.035 41.905 ;
        RECT 86.240 41.115 86.410 41.575 ;
        RECT 87.285 41.405 87.485 41.575 ;
        RECT 88.205 41.445 88.375 42.025 ;
        RECT 88.545 42.125 89.755 43.215 ;
        RECT 88.545 41.585 89.065 42.125 ;
        RECT 88.150 41.405 88.375 41.445 ;
        RECT 89.235 41.415 89.755 41.955 ;
        RECT 85.050 40.945 85.455 41.115 ;
        RECT 85.625 40.945 86.410 41.115 ;
        RECT 86.685 40.665 86.895 41.195 ;
        RECT 87.155 40.880 87.485 41.405 ;
        RECT 87.995 41.320 88.375 41.405 ;
        RECT 87.655 40.665 87.825 41.275 ;
        RECT 87.995 40.885 88.325 41.320 ;
        RECT 88.545 40.665 89.755 41.415 ;
        RECT 12.100 40.495 89.840 40.665 ;
        RECT 12.185 39.745 13.395 40.495 ;
        RECT 13.565 39.950 18.910 40.495 ;
        RECT 19.595 40.105 19.925 40.495 ;
        RECT 12.185 39.205 12.705 39.745 ;
        RECT 12.875 39.035 13.395 39.575 ;
        RECT 15.150 39.120 15.490 39.950 ;
        RECT 20.095 39.925 20.265 40.245 ;
        RECT 20.435 40.105 20.765 40.495 ;
        RECT 21.180 40.095 22.135 40.265 ;
        RECT 19.545 39.755 21.795 39.925 ;
        RECT 12.185 37.945 13.395 39.035 ;
        RECT 16.970 38.380 17.320 39.630 ;
        RECT 19.545 38.795 19.715 39.755 ;
        RECT 19.885 39.135 20.130 39.585 ;
        RECT 20.300 39.305 20.850 39.505 ;
        RECT 21.020 39.335 21.395 39.505 ;
        RECT 21.020 39.135 21.190 39.335 ;
        RECT 21.565 39.255 21.795 39.755 ;
        RECT 19.885 38.965 21.190 39.135 ;
        RECT 21.965 39.215 22.135 40.095 ;
        RECT 22.305 39.660 22.595 40.495 ;
        RECT 22.855 39.945 23.025 40.235 ;
        RECT 23.195 40.115 23.525 40.495 ;
        RECT 22.855 39.775 23.520 39.945 ;
        RECT 21.965 39.045 22.595 39.215 ;
        RECT 13.565 37.945 18.910 38.380 ;
        RECT 19.545 38.115 19.925 38.795 ;
        RECT 20.515 37.945 20.685 38.795 ;
        RECT 20.855 38.625 22.095 38.795 ;
        RECT 20.855 38.115 21.185 38.625 ;
        RECT 21.355 37.945 21.525 38.455 ;
        RECT 21.695 38.115 22.095 38.625 ;
        RECT 22.275 38.115 22.595 39.045 ;
        RECT 22.770 38.955 23.120 39.605 ;
        RECT 23.290 38.785 23.520 39.775 ;
        RECT 22.855 38.615 23.520 38.785 ;
        RECT 22.855 38.115 23.025 38.615 ;
        RECT 23.195 37.945 23.525 38.445 ;
        RECT 23.695 38.115 23.880 40.235 ;
        RECT 24.135 40.035 24.385 40.495 ;
        RECT 24.555 40.045 24.890 40.215 ;
        RECT 25.085 40.045 25.760 40.215 ;
        RECT 24.555 39.905 24.725 40.045 ;
        RECT 24.050 38.915 24.330 39.865 ;
        RECT 24.500 39.775 24.725 39.905 ;
        RECT 24.500 38.670 24.670 39.775 ;
        RECT 24.895 39.625 25.420 39.845 ;
        RECT 24.840 38.860 25.080 39.455 ;
        RECT 25.250 38.925 25.420 39.625 ;
        RECT 25.590 39.265 25.760 40.045 ;
        RECT 26.080 39.995 26.450 40.495 ;
        RECT 26.630 40.045 27.035 40.215 ;
        RECT 27.205 40.045 27.990 40.215 ;
        RECT 26.630 39.815 26.800 40.045 ;
        RECT 25.970 39.515 26.800 39.815 ;
        RECT 27.185 39.545 27.650 39.875 ;
        RECT 25.970 39.485 26.170 39.515 ;
        RECT 26.290 39.265 26.460 39.335 ;
        RECT 25.590 39.095 26.460 39.265 ;
        RECT 25.950 39.005 26.460 39.095 ;
        RECT 24.500 38.540 24.805 38.670 ;
        RECT 25.250 38.560 25.780 38.925 ;
        RECT 24.120 37.945 24.385 38.405 ;
        RECT 24.555 38.115 24.805 38.540 ;
        RECT 25.950 38.390 26.120 39.005 ;
        RECT 25.015 38.220 26.120 38.390 ;
        RECT 26.290 37.945 26.460 38.745 ;
        RECT 26.630 38.445 26.800 39.515 ;
        RECT 26.970 38.615 27.160 39.335 ;
        RECT 27.330 38.585 27.650 39.545 ;
        RECT 27.820 39.585 27.990 40.045 ;
        RECT 28.265 39.965 28.475 40.495 ;
        RECT 28.735 39.755 29.065 40.280 ;
        RECT 29.235 39.885 29.405 40.495 ;
        RECT 29.575 39.840 29.905 40.275 ;
        RECT 30.125 39.845 30.385 40.325 ;
        RECT 30.555 39.955 30.805 40.495 ;
        RECT 29.575 39.755 29.955 39.840 ;
        RECT 28.865 39.585 29.065 39.755 ;
        RECT 29.730 39.715 29.955 39.755 ;
        RECT 27.820 39.255 28.695 39.585 ;
        RECT 28.865 39.255 29.615 39.585 ;
        RECT 26.630 38.115 26.880 38.445 ;
        RECT 27.820 38.415 27.990 39.255 ;
        RECT 28.865 39.050 29.055 39.255 ;
        RECT 29.785 39.135 29.955 39.715 ;
        RECT 29.740 39.085 29.955 39.135 ;
        RECT 28.160 38.675 29.055 39.050 ;
        RECT 29.565 39.005 29.955 39.085 ;
        RECT 27.105 38.245 27.990 38.415 ;
        RECT 28.170 37.945 28.485 38.445 ;
        RECT 28.715 38.115 29.055 38.675 ;
        RECT 29.225 37.945 29.395 38.955 ;
        RECT 29.565 38.160 29.895 39.005 ;
        RECT 30.125 38.815 30.295 39.845 ;
        RECT 30.975 39.815 31.195 40.275 ;
        RECT 30.945 39.790 31.195 39.815 ;
        RECT 30.465 39.195 30.695 39.590 ;
        RECT 30.865 39.365 31.195 39.790 ;
        RECT 31.365 40.115 32.255 40.285 ;
        RECT 31.365 39.390 31.535 40.115 ;
        RECT 31.705 39.560 32.255 39.945 ;
        RECT 32.425 39.745 33.635 40.495 ;
        RECT 33.825 39.805 34.065 40.325 ;
        RECT 34.235 40.000 34.630 40.495 ;
        RECT 35.195 40.165 35.365 40.310 ;
        RECT 34.990 39.970 35.365 40.165 ;
        RECT 31.365 39.320 32.255 39.390 ;
        RECT 31.360 39.295 32.255 39.320 ;
        RECT 31.350 39.280 32.255 39.295 ;
        RECT 31.345 39.265 32.255 39.280 ;
        RECT 31.335 39.260 32.255 39.265 ;
        RECT 31.330 39.250 32.255 39.260 ;
        RECT 31.325 39.240 32.255 39.250 ;
        RECT 31.315 39.235 32.255 39.240 ;
        RECT 31.305 39.225 32.255 39.235 ;
        RECT 31.295 39.220 32.255 39.225 ;
        RECT 31.295 39.215 31.630 39.220 ;
        RECT 31.280 39.210 31.630 39.215 ;
        RECT 31.265 39.200 31.630 39.210 ;
        RECT 31.240 39.195 31.630 39.200 ;
        RECT 30.465 39.190 31.630 39.195 ;
        RECT 30.465 39.155 31.600 39.190 ;
        RECT 30.465 39.130 31.565 39.155 ;
        RECT 30.465 39.100 31.535 39.130 ;
        RECT 30.465 39.070 31.515 39.100 ;
        RECT 30.465 39.040 31.495 39.070 ;
        RECT 30.465 39.030 31.425 39.040 ;
        RECT 30.465 39.020 31.400 39.030 ;
        RECT 30.465 39.005 31.380 39.020 ;
        RECT 30.465 38.990 31.360 39.005 ;
        RECT 30.570 38.980 31.355 38.990 ;
        RECT 30.570 38.945 31.340 38.980 ;
        RECT 30.125 38.115 30.400 38.815 ;
        RECT 30.570 38.695 31.325 38.945 ;
        RECT 31.495 38.625 31.825 38.870 ;
        RECT 31.995 38.770 32.255 39.220 ;
        RECT 32.425 39.205 32.945 39.745 ;
        RECT 33.115 39.035 33.635 39.575 ;
        RECT 31.640 38.600 31.825 38.625 ;
        RECT 31.640 38.500 32.255 38.600 ;
        RECT 30.570 37.945 30.825 38.490 ;
        RECT 30.995 38.115 31.475 38.455 ;
        RECT 31.650 37.945 32.255 38.500 ;
        RECT 32.425 37.945 33.635 39.035 ;
        RECT 33.825 39.000 34.000 39.805 ;
        RECT 34.990 39.635 35.160 39.970 ;
        RECT 35.645 39.925 35.885 40.300 ;
        RECT 36.055 39.990 36.390 40.495 ;
        RECT 35.645 39.775 35.865 39.925 ;
        RECT 34.175 39.275 35.160 39.635 ;
        RECT 35.330 39.445 35.865 39.775 ;
        RECT 34.175 39.255 35.460 39.275 ;
        RECT 34.600 39.105 35.460 39.255 ;
        RECT 33.825 38.215 34.130 39.000 ;
        RECT 34.305 38.625 35.000 38.935 ;
        RECT 34.310 37.945 34.995 38.415 ;
        RECT 35.175 38.160 35.460 39.105 ;
        RECT 35.630 38.795 35.865 39.445 ;
        RECT 36.035 38.965 36.335 39.815 ;
        RECT 36.565 39.745 37.775 40.495 ;
        RECT 37.945 39.770 38.235 40.495 ;
        RECT 36.565 39.205 37.085 39.745 ;
        RECT 37.255 39.035 37.775 39.575 ;
        RECT 35.630 38.565 36.305 38.795 ;
        RECT 35.635 37.945 35.965 38.395 ;
        RECT 36.135 38.135 36.305 38.565 ;
        RECT 36.565 37.945 37.775 39.035 ;
        RECT 37.945 37.945 38.235 39.110 ;
        RECT 38.415 38.125 38.675 40.315 ;
        RECT 38.935 40.125 39.605 40.495 ;
        RECT 39.785 39.945 40.095 40.315 ;
        RECT 38.865 39.745 40.095 39.945 ;
        RECT 38.865 39.075 39.155 39.745 ;
        RECT 40.275 39.565 40.505 40.205 ;
        RECT 40.685 39.765 40.975 40.495 ;
        RECT 41.165 39.950 46.510 40.495 ;
        RECT 46.685 39.950 52.030 40.495 ;
        RECT 39.335 39.255 39.800 39.565 ;
        RECT 39.980 39.255 40.505 39.565 ;
        RECT 40.685 39.255 40.985 39.585 ;
        RECT 42.750 39.120 43.090 39.950 ;
        RECT 38.865 38.855 39.635 39.075 ;
        RECT 38.845 37.945 39.185 38.675 ;
        RECT 39.365 38.125 39.635 38.855 ;
        RECT 39.815 38.835 40.975 39.075 ;
        RECT 39.815 38.125 40.045 38.835 ;
        RECT 40.215 37.945 40.545 38.655 ;
        RECT 40.715 38.125 40.975 38.835 ;
        RECT 44.570 38.380 44.920 39.630 ;
        RECT 48.270 39.120 48.610 39.950 ;
        RECT 52.205 39.725 53.875 40.495 ;
        RECT 50.090 38.380 50.440 39.630 ;
        RECT 52.205 39.205 52.955 39.725 ;
        RECT 54.045 39.695 54.740 40.325 ;
        RECT 54.945 39.695 55.255 40.495 ;
        RECT 55.430 39.965 55.720 40.315 ;
        RECT 55.915 40.135 56.245 40.495 ;
        RECT 56.415 39.965 56.645 40.270 ;
        RECT 55.430 39.795 56.645 39.965 ;
        RECT 53.125 39.035 53.875 39.555 ;
        RECT 54.065 39.255 54.400 39.505 ;
        RECT 54.570 39.095 54.740 39.695 ;
        RECT 56.835 39.625 57.005 40.190 ;
        RECT 54.910 39.255 55.245 39.525 ;
        RECT 55.490 39.475 55.750 39.585 ;
        RECT 55.485 39.305 55.750 39.475 ;
        RECT 55.490 39.255 55.750 39.305 ;
        RECT 55.930 39.255 56.315 39.585 ;
        RECT 56.485 39.455 57.005 39.625 ;
        RECT 58.185 39.845 58.445 40.325 ;
        RECT 58.615 39.955 58.865 40.495 ;
        RECT 41.165 37.945 46.510 38.380 ;
        RECT 46.685 37.945 52.030 38.380 ;
        RECT 52.205 37.945 53.875 39.035 ;
        RECT 54.045 37.945 54.305 39.085 ;
        RECT 54.475 38.115 54.805 39.095 ;
        RECT 54.975 37.945 55.255 39.085 ;
        RECT 55.430 37.945 55.750 39.085 ;
        RECT 55.930 38.205 56.125 39.255 ;
        RECT 56.485 39.075 56.655 39.455 ;
        RECT 56.305 38.795 56.655 39.075 ;
        RECT 56.845 38.925 57.090 39.285 ;
        RECT 58.185 38.815 58.355 39.845 ;
        RECT 59.035 39.790 59.255 40.275 ;
        RECT 58.525 39.195 58.755 39.590 ;
        RECT 58.925 39.365 59.255 39.790 ;
        RECT 59.425 40.115 60.315 40.285 ;
        RECT 59.425 39.390 59.595 40.115 ;
        RECT 59.765 39.560 60.315 39.945 ;
        RECT 60.485 39.675 60.745 40.495 ;
        RECT 60.915 39.675 61.245 40.095 ;
        RECT 61.425 40.010 62.215 40.275 ;
        RECT 60.995 39.585 61.245 39.675 ;
        RECT 59.425 39.320 60.315 39.390 ;
        RECT 59.420 39.295 60.315 39.320 ;
        RECT 59.410 39.280 60.315 39.295 ;
        RECT 59.405 39.265 60.315 39.280 ;
        RECT 59.395 39.260 60.315 39.265 ;
        RECT 59.390 39.250 60.315 39.260 ;
        RECT 59.385 39.240 60.315 39.250 ;
        RECT 59.375 39.235 60.315 39.240 ;
        RECT 59.365 39.225 60.315 39.235 ;
        RECT 59.355 39.220 60.315 39.225 ;
        RECT 59.355 39.215 59.690 39.220 ;
        RECT 59.340 39.210 59.690 39.215 ;
        RECT 59.325 39.200 59.690 39.210 ;
        RECT 59.300 39.195 59.690 39.200 ;
        RECT 58.525 39.190 59.690 39.195 ;
        RECT 58.525 39.155 59.660 39.190 ;
        RECT 58.525 39.130 59.625 39.155 ;
        RECT 58.525 39.100 59.595 39.130 ;
        RECT 58.525 39.070 59.575 39.100 ;
        RECT 58.525 39.040 59.555 39.070 ;
        RECT 58.525 39.030 59.485 39.040 ;
        RECT 58.525 39.020 59.460 39.030 ;
        RECT 58.525 39.005 59.440 39.020 ;
        RECT 58.525 38.990 59.420 39.005 ;
        RECT 58.630 38.980 59.415 38.990 ;
        RECT 58.630 38.945 59.400 38.980 ;
        RECT 56.305 38.115 56.635 38.795 ;
        RECT 56.835 37.945 57.090 38.745 ;
        RECT 58.185 38.115 58.460 38.815 ;
        RECT 58.630 38.695 59.385 38.945 ;
        RECT 59.555 38.625 59.885 38.870 ;
        RECT 60.055 38.770 60.315 39.220 ;
        RECT 60.485 38.625 60.825 39.505 ;
        RECT 60.995 39.335 61.790 39.585 ;
        RECT 59.700 38.600 59.885 38.625 ;
        RECT 59.700 38.500 60.315 38.600 ;
        RECT 58.630 37.945 58.885 38.490 ;
        RECT 59.055 38.115 59.535 38.455 ;
        RECT 59.710 37.945 60.315 38.500 ;
        RECT 60.485 37.945 60.745 38.455 ;
        RECT 60.995 38.115 61.165 39.335 ;
        RECT 61.960 39.155 62.215 40.010 ;
        RECT 62.385 39.855 62.585 40.275 ;
        RECT 62.775 40.035 63.105 40.495 ;
        RECT 62.385 39.335 62.795 39.855 ;
        RECT 63.275 39.845 63.535 40.325 ;
        RECT 62.965 39.155 63.195 39.585 ;
        RECT 61.405 38.985 63.195 39.155 ;
        RECT 61.405 38.620 61.655 38.985 ;
        RECT 61.825 38.625 62.155 38.815 ;
        RECT 62.375 38.690 63.090 38.985 ;
        RECT 63.365 38.815 63.535 39.845 ;
        RECT 63.705 39.770 63.995 40.495 ;
        RECT 64.165 39.675 64.425 40.495 ;
        RECT 64.595 39.675 64.925 40.095 ;
        RECT 65.105 39.925 65.365 40.325 ;
        RECT 65.535 40.095 65.865 40.495 ;
        RECT 66.035 39.925 66.205 40.275 ;
        RECT 66.375 40.095 66.750 40.495 ;
        RECT 65.105 39.755 66.770 39.925 ;
        RECT 66.940 39.820 67.215 40.165 ;
        RECT 64.675 39.585 64.925 39.675 ;
        RECT 66.600 39.585 66.770 39.755 ;
        RECT 64.170 39.255 64.505 39.505 ;
        RECT 64.675 39.255 65.390 39.585 ;
        RECT 65.605 39.255 66.430 39.585 ;
        RECT 66.600 39.255 66.875 39.585 ;
        RECT 61.825 38.450 62.020 38.625 ;
        RECT 61.405 37.945 62.020 38.450 ;
        RECT 62.190 38.115 62.665 38.455 ;
        RECT 62.835 37.945 63.050 38.490 ;
        RECT 63.260 38.115 63.535 38.815 ;
        RECT 63.705 37.945 63.995 39.110 ;
        RECT 64.165 37.945 64.425 39.085 ;
        RECT 64.675 38.695 64.845 39.255 ;
        RECT 65.105 38.795 65.435 39.085 ;
        RECT 65.605 38.965 65.850 39.255 ;
        RECT 66.600 39.085 66.770 39.255 ;
        RECT 67.045 39.085 67.215 39.820 ;
        RECT 68.310 39.655 68.570 40.495 ;
        RECT 68.745 39.750 69.000 40.325 ;
        RECT 69.170 40.115 69.500 40.495 ;
        RECT 69.715 39.945 69.885 40.325 ;
        RECT 69.170 39.775 69.885 39.945 ;
        RECT 66.110 38.915 66.770 39.085 ;
        RECT 66.110 38.795 66.280 38.915 ;
        RECT 65.105 38.625 66.280 38.795 ;
        RECT 64.665 38.125 66.280 38.455 ;
        RECT 66.450 37.945 66.730 38.745 ;
        RECT 66.940 38.115 67.215 39.085 ;
        RECT 68.310 37.945 68.570 39.095 ;
        RECT 68.745 39.020 68.915 39.750 ;
        RECT 69.170 39.585 69.340 39.775 ;
        RECT 70.150 39.655 70.410 40.495 ;
        RECT 70.585 39.750 70.840 40.325 ;
        RECT 71.010 40.115 71.340 40.495 ;
        RECT 71.555 39.945 71.725 40.325 ;
        RECT 71.010 39.775 71.725 39.945 ;
        RECT 69.085 39.255 69.340 39.585 ;
        RECT 69.170 39.045 69.340 39.255 ;
        RECT 69.620 39.225 69.975 39.595 ;
        RECT 68.745 38.115 69.000 39.020 ;
        RECT 69.170 38.875 69.885 39.045 ;
        RECT 69.170 37.945 69.500 38.705 ;
        RECT 69.715 38.115 69.885 38.875 ;
        RECT 70.150 37.945 70.410 39.095 ;
        RECT 70.585 39.020 70.755 39.750 ;
        RECT 71.010 39.585 71.180 39.775 ;
        RECT 72.020 39.755 72.635 40.325 ;
        RECT 72.805 39.985 73.020 40.495 ;
        RECT 73.250 39.985 73.530 40.315 ;
        RECT 73.710 39.985 73.950 40.495 ;
        RECT 70.925 39.255 71.180 39.585 ;
        RECT 71.010 39.045 71.180 39.255 ;
        RECT 71.460 39.225 71.815 39.595 ;
        RECT 70.585 38.115 70.840 39.020 ;
        RECT 71.010 38.875 71.725 39.045 ;
        RECT 71.010 37.945 71.340 38.705 ;
        RECT 71.555 38.115 71.725 38.875 ;
        RECT 72.020 38.735 72.335 39.755 ;
        RECT 72.505 39.085 72.675 39.585 ;
        RECT 72.925 39.255 73.190 39.815 ;
        RECT 73.360 39.085 73.530 39.985 ;
        RECT 73.700 39.255 74.055 39.815 ;
        RECT 74.320 39.755 74.935 40.325 ;
        RECT 75.105 39.985 75.320 40.495 ;
        RECT 75.550 39.985 75.830 40.315 ;
        RECT 76.010 39.985 76.250 40.495 ;
        RECT 72.505 38.915 73.930 39.085 ;
        RECT 72.020 38.115 72.555 38.735 ;
        RECT 72.725 37.945 73.055 38.745 ;
        RECT 73.540 38.740 73.930 38.915 ;
        RECT 74.320 38.735 74.635 39.755 ;
        RECT 74.805 39.085 74.975 39.585 ;
        RECT 75.225 39.255 75.490 39.815 ;
        RECT 75.660 39.085 75.830 39.985 ;
        RECT 76.000 39.255 76.355 39.815 ;
        RECT 77.080 39.755 77.695 40.325 ;
        RECT 77.865 39.985 78.080 40.495 ;
        RECT 78.310 39.985 78.590 40.315 ;
        RECT 78.770 39.985 79.010 40.495 ;
        RECT 74.805 38.915 76.230 39.085 ;
        RECT 74.320 38.115 74.855 38.735 ;
        RECT 75.025 37.945 75.355 38.745 ;
        RECT 75.840 38.740 76.230 38.915 ;
        RECT 77.080 38.735 77.395 39.755 ;
        RECT 77.565 39.085 77.735 39.585 ;
        RECT 77.985 39.255 78.250 39.815 ;
        RECT 78.420 39.085 78.590 39.985 ;
        RECT 79.435 39.945 79.605 40.325 ;
        RECT 79.820 40.115 80.150 40.495 ;
        RECT 78.760 39.255 79.115 39.815 ;
        RECT 79.435 39.775 80.150 39.945 ;
        RECT 79.345 39.225 79.700 39.595 ;
        RECT 79.980 39.585 80.150 39.775 ;
        RECT 80.320 39.750 80.575 40.325 ;
        RECT 79.980 39.255 80.235 39.585 ;
        RECT 77.565 38.915 78.990 39.085 ;
        RECT 79.980 39.045 80.150 39.255 ;
        RECT 77.080 38.115 77.615 38.735 ;
        RECT 77.785 37.945 78.115 38.745 ;
        RECT 78.600 38.740 78.990 38.915 ;
        RECT 79.435 38.875 80.150 39.045 ;
        RECT 80.405 39.020 80.575 39.750 ;
        RECT 80.750 39.655 81.010 40.495 ;
        RECT 81.390 39.715 81.890 40.325 ;
        RECT 81.185 39.255 81.535 39.505 ;
        RECT 79.435 38.115 79.605 38.875 ;
        RECT 79.820 37.945 80.150 38.705 ;
        RECT 80.320 38.115 80.575 39.020 ;
        RECT 80.750 37.945 81.010 39.095 ;
        RECT 81.720 39.085 81.890 39.715 ;
        RECT 82.520 39.845 82.850 40.325 ;
        RECT 83.020 40.035 83.245 40.495 ;
        RECT 83.415 39.845 83.745 40.325 ;
        RECT 82.520 39.675 83.745 39.845 ;
        RECT 83.935 39.695 84.185 40.495 ;
        RECT 84.355 39.695 84.695 40.325 ;
        RECT 82.060 39.305 82.390 39.505 ;
        RECT 82.560 39.305 82.890 39.505 ;
        RECT 83.060 39.475 83.480 39.505 ;
        RECT 83.060 39.305 83.485 39.475 ;
        RECT 83.655 39.335 84.350 39.505 ;
        RECT 83.655 39.085 83.825 39.335 ;
        RECT 84.520 39.085 84.695 39.695 ;
        RECT 81.390 38.915 83.825 39.085 ;
        RECT 81.390 38.115 81.720 38.915 ;
        RECT 81.890 37.945 82.220 38.745 ;
        RECT 82.520 38.115 82.850 38.915 ;
        RECT 83.495 37.945 83.745 38.745 ;
        RECT 84.015 37.945 84.185 39.085 ;
        RECT 84.355 38.115 84.695 39.085 ;
        RECT 84.865 39.995 85.125 40.325 ;
        RECT 85.295 40.135 85.625 40.495 ;
        RECT 85.880 40.115 87.180 40.325 ;
        RECT 84.865 39.985 85.095 39.995 ;
        RECT 84.865 38.795 85.035 39.985 ;
        RECT 85.880 39.965 86.050 40.115 ;
        RECT 85.295 39.840 86.050 39.965 ;
        RECT 85.205 39.795 86.050 39.840 ;
        RECT 85.205 39.675 85.475 39.795 ;
        RECT 85.205 39.100 85.375 39.675 ;
        RECT 85.605 39.235 86.015 39.540 ;
        RECT 86.305 39.505 86.515 39.905 ;
        RECT 86.185 39.295 86.515 39.505 ;
        RECT 86.760 39.505 86.980 39.905 ;
        RECT 87.455 39.730 87.910 40.495 ;
        RECT 88.545 39.745 89.755 40.495 ;
        RECT 86.760 39.295 87.235 39.505 ;
        RECT 87.425 39.305 87.915 39.505 ;
        RECT 85.205 39.065 85.405 39.100 ;
        RECT 86.735 39.065 87.910 39.125 ;
        RECT 85.205 38.955 87.910 39.065 ;
        RECT 85.265 38.895 87.065 38.955 ;
        RECT 86.735 38.865 87.065 38.895 ;
        RECT 84.865 38.115 85.125 38.795 ;
        RECT 85.295 37.945 85.545 38.725 ;
        RECT 85.795 38.695 86.630 38.705 ;
        RECT 87.220 38.695 87.405 38.785 ;
        RECT 85.795 38.495 87.405 38.695 ;
        RECT 85.795 38.115 86.045 38.495 ;
        RECT 87.175 38.455 87.405 38.495 ;
        RECT 87.655 38.335 87.910 38.955 ;
        RECT 86.215 37.945 86.570 38.325 ;
        RECT 87.575 38.115 87.910 38.335 ;
        RECT 88.545 39.035 89.065 39.575 ;
        RECT 89.235 39.205 89.755 39.745 ;
        RECT 88.545 37.945 89.755 39.035 ;
        RECT 12.100 37.775 89.840 37.945 ;
        RECT 12.185 36.685 13.395 37.775 ;
        RECT 13.565 37.340 18.910 37.775 ;
        RECT 19.085 37.340 24.430 37.775 ;
        RECT 12.185 35.975 12.705 36.515 ;
        RECT 12.875 36.145 13.395 36.685 ;
        RECT 12.185 35.225 13.395 35.975 ;
        RECT 15.150 35.770 15.490 36.600 ;
        RECT 16.970 36.090 17.320 37.340 ;
        RECT 20.670 35.770 21.010 36.600 ;
        RECT 22.490 36.090 22.840 37.340 ;
        RECT 25.065 36.610 25.355 37.775 ;
        RECT 25.585 36.715 25.915 37.560 ;
        RECT 26.085 36.765 26.255 37.775 ;
        RECT 26.425 37.045 26.765 37.605 ;
        RECT 26.995 37.275 27.310 37.775 ;
        RECT 27.490 37.305 28.375 37.475 ;
        RECT 25.525 36.635 25.915 36.715 ;
        RECT 26.425 36.670 27.320 37.045 ;
        RECT 25.525 36.585 25.740 36.635 ;
        RECT 25.525 36.005 25.695 36.585 ;
        RECT 26.425 36.465 26.615 36.670 ;
        RECT 27.490 36.465 27.660 37.305 ;
        RECT 28.600 37.275 28.850 37.605 ;
        RECT 25.865 36.135 26.615 36.465 ;
        RECT 26.785 36.135 27.660 36.465 ;
        RECT 25.525 35.965 25.750 36.005 ;
        RECT 26.415 35.965 26.615 36.135 ;
        RECT 13.565 35.225 18.910 35.770 ;
        RECT 19.085 35.225 24.430 35.770 ;
        RECT 25.065 35.225 25.355 35.950 ;
        RECT 25.525 35.880 25.905 35.965 ;
        RECT 25.575 35.445 25.905 35.880 ;
        RECT 26.075 35.225 26.245 35.835 ;
        RECT 26.415 35.440 26.745 35.965 ;
        RECT 27.005 35.225 27.215 35.755 ;
        RECT 27.490 35.675 27.660 36.135 ;
        RECT 27.830 36.175 28.150 37.135 ;
        RECT 28.320 36.385 28.510 37.105 ;
        RECT 28.680 36.205 28.850 37.275 ;
        RECT 29.020 36.975 29.190 37.775 ;
        RECT 29.360 37.330 30.465 37.500 ;
        RECT 29.360 36.715 29.530 37.330 ;
        RECT 30.675 37.180 30.925 37.605 ;
        RECT 31.095 37.315 31.360 37.775 ;
        RECT 29.700 36.795 30.230 37.160 ;
        RECT 30.675 37.050 30.980 37.180 ;
        RECT 29.020 36.625 29.530 36.715 ;
        RECT 29.020 36.455 29.890 36.625 ;
        RECT 29.020 36.385 29.190 36.455 ;
        RECT 29.310 36.205 29.510 36.235 ;
        RECT 27.830 35.845 28.295 36.175 ;
        RECT 28.680 35.905 29.510 36.205 ;
        RECT 28.680 35.675 28.850 35.905 ;
        RECT 27.490 35.505 28.275 35.675 ;
        RECT 28.445 35.505 28.850 35.675 ;
        RECT 29.030 35.225 29.400 35.725 ;
        RECT 29.720 35.675 29.890 36.455 ;
        RECT 30.060 36.095 30.230 36.795 ;
        RECT 30.400 36.265 30.640 36.860 ;
        RECT 30.060 35.875 30.585 36.095 ;
        RECT 30.810 35.945 30.980 37.050 ;
        RECT 30.755 35.815 30.980 35.945 ;
        RECT 31.150 35.855 31.430 36.805 ;
        RECT 30.755 35.675 30.925 35.815 ;
        RECT 29.720 35.505 30.395 35.675 ;
        RECT 30.590 35.505 30.925 35.675 ;
        RECT 31.095 35.225 31.345 35.685 ;
        RECT 31.600 35.485 31.785 37.605 ;
        RECT 31.955 37.275 32.285 37.775 ;
        RECT 32.455 37.105 32.625 37.605 ;
        RECT 31.960 36.935 32.625 37.105 ;
        RECT 32.975 37.105 33.145 37.605 ;
        RECT 33.315 37.275 33.645 37.775 ;
        RECT 32.975 36.935 33.640 37.105 ;
        RECT 31.960 35.945 32.190 36.935 ;
        RECT 32.360 36.115 32.710 36.765 ;
        RECT 32.890 36.115 33.240 36.765 ;
        RECT 33.410 35.945 33.640 36.935 ;
        RECT 31.960 35.775 32.625 35.945 ;
        RECT 31.955 35.225 32.285 35.605 ;
        RECT 32.455 35.485 32.625 35.775 ;
        RECT 32.975 35.775 33.640 35.945 ;
        RECT 32.975 35.485 33.145 35.775 ;
        RECT 33.315 35.225 33.645 35.605 ;
        RECT 33.815 35.485 34.000 37.605 ;
        RECT 34.240 37.315 34.505 37.775 ;
        RECT 34.675 37.180 34.925 37.605 ;
        RECT 35.135 37.330 36.240 37.500 ;
        RECT 34.620 37.050 34.925 37.180 ;
        RECT 34.170 35.855 34.450 36.805 ;
        RECT 34.620 35.945 34.790 37.050 ;
        RECT 34.960 36.265 35.200 36.860 ;
        RECT 35.370 36.795 35.900 37.160 ;
        RECT 35.370 36.095 35.540 36.795 ;
        RECT 36.070 36.715 36.240 37.330 ;
        RECT 36.410 36.975 36.580 37.775 ;
        RECT 36.750 37.275 37.000 37.605 ;
        RECT 37.225 37.305 38.110 37.475 ;
        RECT 36.070 36.625 36.580 36.715 ;
        RECT 34.620 35.815 34.845 35.945 ;
        RECT 35.015 35.875 35.540 36.095 ;
        RECT 35.710 36.455 36.580 36.625 ;
        RECT 34.255 35.225 34.505 35.685 ;
        RECT 34.675 35.675 34.845 35.815 ;
        RECT 35.710 35.675 35.880 36.455 ;
        RECT 36.410 36.385 36.580 36.455 ;
        RECT 36.090 36.205 36.290 36.235 ;
        RECT 36.750 36.205 36.920 37.275 ;
        RECT 37.090 36.385 37.280 37.105 ;
        RECT 36.090 35.905 36.920 36.205 ;
        RECT 37.450 36.175 37.770 37.135 ;
        RECT 34.675 35.505 35.010 35.675 ;
        RECT 35.205 35.505 35.880 35.675 ;
        RECT 36.200 35.225 36.570 35.725 ;
        RECT 36.750 35.675 36.920 35.905 ;
        RECT 37.305 35.845 37.770 36.175 ;
        RECT 37.940 36.465 38.110 37.305 ;
        RECT 38.290 37.275 38.605 37.775 ;
        RECT 38.835 37.045 39.175 37.605 ;
        RECT 38.280 36.670 39.175 37.045 ;
        RECT 39.345 36.765 39.515 37.775 ;
        RECT 38.985 36.465 39.175 36.670 ;
        RECT 39.685 36.715 40.015 37.560 ;
        RECT 40.245 37.340 45.590 37.775 ;
        RECT 39.685 36.635 40.075 36.715 ;
        RECT 39.860 36.585 40.075 36.635 ;
        RECT 37.940 36.135 38.815 36.465 ;
        RECT 38.985 36.135 39.735 36.465 ;
        RECT 37.940 35.675 38.110 36.135 ;
        RECT 38.985 35.965 39.185 36.135 ;
        RECT 39.905 36.005 40.075 36.585 ;
        RECT 39.850 35.965 40.075 36.005 ;
        RECT 36.750 35.505 37.155 35.675 ;
        RECT 37.325 35.505 38.110 35.675 ;
        RECT 38.385 35.225 38.595 35.755 ;
        RECT 38.855 35.440 39.185 35.965 ;
        RECT 39.695 35.880 40.075 35.965 ;
        RECT 39.355 35.225 39.525 35.835 ;
        RECT 39.695 35.445 40.025 35.880 ;
        RECT 41.830 35.770 42.170 36.600 ;
        RECT 43.650 36.090 44.000 37.340 ;
        RECT 45.765 36.685 49.275 37.775 ;
        RECT 49.445 36.685 50.655 37.775 ;
        RECT 45.765 35.995 47.415 36.515 ;
        RECT 47.585 36.165 49.275 36.685 ;
        RECT 40.245 35.225 45.590 35.770 ;
        RECT 45.765 35.225 49.275 35.995 ;
        RECT 49.445 35.975 49.965 36.515 ;
        RECT 50.135 36.145 50.655 36.685 ;
        RECT 50.825 36.610 51.115 37.775 ;
        RECT 51.285 37.340 56.630 37.775 ;
        RECT 49.445 35.225 50.655 35.975 ;
        RECT 50.825 35.225 51.115 35.950 ;
        RECT 52.870 35.770 53.210 36.600 ;
        RECT 54.690 36.090 55.040 37.340 ;
        RECT 56.805 36.685 58.475 37.775 ;
        RECT 56.805 35.995 57.555 36.515 ;
        RECT 57.725 36.165 58.475 36.685 ;
        RECT 59.105 36.635 59.385 37.775 ;
        RECT 59.555 36.625 59.885 37.605 ;
        RECT 60.055 36.635 60.315 37.775 ;
        RECT 60.495 36.805 60.825 37.590 ;
        RECT 60.495 36.635 61.175 36.805 ;
        RECT 61.355 36.635 61.685 37.775 ;
        RECT 61.865 36.685 63.075 37.775 ;
        RECT 59.115 36.195 59.450 36.465 ;
        RECT 59.620 36.025 59.790 36.625 ;
        RECT 59.960 36.215 60.295 36.465 ;
        RECT 60.485 36.215 60.835 36.465 ;
        RECT 61.005 36.035 61.175 36.635 ;
        RECT 61.345 36.215 61.695 36.465 ;
        RECT 51.285 35.225 56.630 35.770 ;
        RECT 56.805 35.225 58.475 35.995 ;
        RECT 59.105 35.225 59.415 36.025 ;
        RECT 59.620 35.395 60.315 36.025 ;
        RECT 60.505 35.225 60.745 36.035 ;
        RECT 60.915 35.395 61.245 36.035 ;
        RECT 61.415 35.225 61.685 36.035 ;
        RECT 61.865 35.975 62.385 36.515 ;
        RECT 62.555 36.145 63.075 36.685 ;
        RECT 63.285 36.635 63.515 37.775 ;
        RECT 63.685 36.625 64.015 37.605 ;
        RECT 64.185 36.635 64.395 37.775 ;
        RECT 64.625 36.685 65.835 37.775 ;
        RECT 63.265 36.215 63.595 36.465 ;
        RECT 61.865 35.225 63.075 35.975 ;
        RECT 63.285 35.225 63.515 36.045 ;
        RECT 63.765 36.025 64.015 36.625 ;
        RECT 63.685 35.395 64.015 36.025 ;
        RECT 64.185 35.225 64.395 36.045 ;
        RECT 64.625 35.975 65.145 36.515 ;
        RECT 65.315 36.145 65.835 36.685 ;
        RECT 66.010 36.625 66.270 37.775 ;
        RECT 66.445 36.700 66.700 37.605 ;
        RECT 66.870 37.015 67.200 37.775 ;
        RECT 67.415 36.845 67.585 37.605 ;
        RECT 64.625 35.225 65.835 35.975 ;
        RECT 66.010 35.225 66.270 36.065 ;
        RECT 66.445 35.970 66.615 36.700 ;
        RECT 66.870 36.675 67.585 36.845 ;
        RECT 66.870 36.465 67.040 36.675 ;
        RECT 67.850 36.625 68.110 37.775 ;
        RECT 68.285 36.700 68.540 37.605 ;
        RECT 68.710 37.015 69.040 37.775 ;
        RECT 69.255 36.845 69.425 37.605 ;
        RECT 66.785 36.135 67.040 36.465 ;
        RECT 66.445 35.395 66.700 35.970 ;
        RECT 66.870 35.945 67.040 36.135 ;
        RECT 67.320 36.125 67.675 36.495 ;
        RECT 66.870 35.775 67.585 35.945 ;
        RECT 66.870 35.225 67.200 35.605 ;
        RECT 67.415 35.395 67.585 35.775 ;
        RECT 67.850 35.225 68.110 36.065 ;
        RECT 68.285 35.970 68.455 36.700 ;
        RECT 68.710 36.675 69.425 36.845 ;
        RECT 69.720 36.985 70.255 37.605 ;
        RECT 68.710 36.465 68.880 36.675 ;
        RECT 68.625 36.135 68.880 36.465 ;
        RECT 68.285 35.395 68.540 35.970 ;
        RECT 68.710 35.945 68.880 36.135 ;
        RECT 69.160 36.125 69.515 36.495 ;
        RECT 69.720 35.965 70.035 36.985 ;
        RECT 70.425 36.975 70.755 37.775 ;
        RECT 71.240 36.805 71.630 36.980 ;
        RECT 70.205 36.635 71.630 36.805 ;
        RECT 72.170 36.805 72.560 36.980 ;
        RECT 73.045 36.975 73.375 37.775 ;
        RECT 73.545 36.985 74.080 37.605 ;
        RECT 72.170 36.635 73.595 36.805 ;
        RECT 70.205 36.135 70.375 36.635 ;
        RECT 68.710 35.775 69.425 35.945 ;
        RECT 68.710 35.225 69.040 35.605 ;
        RECT 69.255 35.395 69.425 35.775 ;
        RECT 69.720 35.395 70.335 35.965 ;
        RECT 70.625 35.905 70.890 36.465 ;
        RECT 71.060 35.735 71.230 36.635 ;
        RECT 71.400 35.905 71.755 36.465 ;
        RECT 72.045 35.905 72.400 36.465 ;
        RECT 72.570 35.735 72.740 36.635 ;
        RECT 72.910 35.905 73.175 36.465 ;
        RECT 73.425 36.135 73.595 36.635 ;
        RECT 73.765 35.965 74.080 36.985 ;
        RECT 74.470 36.805 74.860 36.980 ;
        RECT 75.345 36.975 75.675 37.775 ;
        RECT 75.845 36.985 76.380 37.605 ;
        RECT 74.470 36.635 75.895 36.805 ;
        RECT 70.505 35.225 70.720 35.735 ;
        RECT 70.950 35.405 71.230 35.735 ;
        RECT 71.410 35.225 71.650 35.735 ;
        RECT 72.150 35.225 72.390 35.735 ;
        RECT 72.570 35.405 72.850 35.735 ;
        RECT 73.080 35.225 73.295 35.735 ;
        RECT 73.465 35.395 74.080 35.965 ;
        RECT 74.345 35.905 74.700 36.465 ;
        RECT 74.870 35.735 75.040 36.635 ;
        RECT 75.210 35.905 75.475 36.465 ;
        RECT 75.725 36.135 75.895 36.635 ;
        RECT 76.065 35.965 76.380 36.985 ;
        RECT 76.585 36.610 76.875 37.775 ;
        RECT 77.050 37.385 77.385 37.605 ;
        RECT 78.390 37.395 78.745 37.775 ;
        RECT 77.050 36.765 77.305 37.385 ;
        RECT 77.555 37.225 77.785 37.265 ;
        RECT 78.915 37.225 79.165 37.605 ;
        RECT 77.555 37.025 79.165 37.225 ;
        RECT 77.555 36.935 77.740 37.025 ;
        RECT 78.330 37.015 79.165 37.025 ;
        RECT 79.415 36.995 79.665 37.775 ;
        RECT 79.835 36.925 80.095 37.605 ;
        RECT 77.895 36.825 78.225 36.855 ;
        RECT 77.895 36.765 79.695 36.825 ;
        RECT 77.050 36.655 79.755 36.765 ;
        RECT 77.050 36.595 78.225 36.655 ;
        RECT 79.555 36.620 79.755 36.655 ;
        RECT 77.045 36.215 77.535 36.415 ;
        RECT 77.725 36.215 78.200 36.425 ;
        RECT 74.450 35.225 74.690 35.735 ;
        RECT 74.870 35.405 75.150 35.735 ;
        RECT 75.380 35.225 75.595 35.735 ;
        RECT 75.765 35.395 76.380 35.965 ;
        RECT 76.585 35.225 76.875 35.950 ;
        RECT 77.050 35.225 77.505 35.990 ;
        RECT 77.980 35.815 78.200 36.215 ;
        RECT 78.445 36.215 78.775 36.425 ;
        RECT 78.445 35.815 78.655 36.215 ;
        RECT 78.945 36.180 79.355 36.485 ;
        RECT 79.585 36.045 79.755 36.620 ;
        RECT 79.485 35.925 79.755 36.045 ;
        RECT 78.910 35.880 79.755 35.925 ;
        RECT 78.910 35.755 79.665 35.880 ;
        RECT 78.910 35.605 79.080 35.755 ;
        RECT 79.925 35.735 80.095 36.925 ;
        RECT 79.865 35.725 80.095 35.735 ;
        RECT 77.780 35.395 79.080 35.605 ;
        RECT 79.335 35.225 79.665 35.585 ;
        RECT 79.835 35.395 80.095 35.725 ;
        RECT 80.265 36.925 80.525 37.605 ;
        RECT 80.695 36.995 80.945 37.775 ;
        RECT 81.195 37.225 81.445 37.605 ;
        RECT 81.615 37.395 81.970 37.775 ;
        RECT 82.975 37.385 83.310 37.605 ;
        RECT 82.575 37.225 82.805 37.265 ;
        RECT 81.195 37.025 82.805 37.225 ;
        RECT 81.195 37.015 82.030 37.025 ;
        RECT 82.620 36.935 82.805 37.025 ;
        RECT 80.265 35.725 80.435 36.925 ;
        RECT 82.135 36.825 82.465 36.855 ;
        RECT 80.665 36.765 82.465 36.825 ;
        RECT 83.055 36.765 83.310 37.385 ;
        RECT 80.605 36.655 83.310 36.765 ;
        RECT 80.605 36.620 80.805 36.655 ;
        RECT 80.605 36.045 80.775 36.620 ;
        RECT 82.135 36.595 83.310 36.655 ;
        RECT 83.945 36.635 84.285 37.605 ;
        RECT 84.455 36.635 84.625 37.775 ;
        RECT 84.895 36.975 85.145 37.775 ;
        RECT 85.790 36.805 86.120 37.605 ;
        RECT 86.420 36.975 86.750 37.775 ;
        RECT 86.920 36.805 87.250 37.605 ;
        RECT 84.815 36.635 87.250 36.805 ;
        RECT 88.545 36.685 89.755 37.775 ;
        RECT 81.005 36.180 81.415 36.485 ;
        RECT 81.585 36.215 81.915 36.425 ;
        RECT 80.605 35.925 80.875 36.045 ;
        RECT 80.605 35.880 81.450 35.925 ;
        RECT 80.695 35.755 81.450 35.880 ;
        RECT 81.705 35.815 81.915 36.215 ;
        RECT 82.160 36.215 82.635 36.425 ;
        RECT 82.825 36.215 83.315 36.415 ;
        RECT 82.160 35.815 82.380 36.215 ;
        RECT 83.945 36.025 84.120 36.635 ;
        RECT 84.815 36.385 84.985 36.635 ;
        RECT 84.290 36.215 84.985 36.385 ;
        RECT 85.160 36.215 85.580 36.415 ;
        RECT 85.750 36.215 86.080 36.415 ;
        RECT 86.250 36.215 86.580 36.415 ;
        RECT 80.265 35.395 80.525 35.725 ;
        RECT 81.280 35.605 81.450 35.755 ;
        RECT 80.695 35.225 81.025 35.585 ;
        RECT 81.280 35.395 82.580 35.605 ;
        RECT 82.855 35.225 83.310 35.990 ;
        RECT 83.945 35.395 84.285 36.025 ;
        RECT 84.455 35.225 84.705 36.025 ;
        RECT 84.895 35.875 86.120 36.045 ;
        RECT 84.895 35.395 85.225 35.875 ;
        RECT 85.395 35.225 85.620 35.685 ;
        RECT 85.790 35.395 86.120 35.875 ;
        RECT 86.750 36.005 86.920 36.635 ;
        RECT 87.105 36.215 87.455 36.465 ;
        RECT 88.545 36.145 89.065 36.685 ;
        RECT 86.750 35.395 87.250 36.005 ;
        RECT 89.235 35.975 89.755 36.515 ;
        RECT 88.545 35.225 89.755 35.975 ;
        RECT 12.100 35.055 89.840 35.225 ;
        RECT 12.185 34.305 13.395 35.055 ;
        RECT 13.565 34.510 18.910 35.055 ;
        RECT 19.085 34.510 24.430 35.055 ;
        RECT 24.605 34.510 29.950 35.055 ;
        RECT 30.125 34.510 35.470 35.055 ;
        RECT 12.185 33.765 12.705 34.305 ;
        RECT 12.875 33.595 13.395 34.135 ;
        RECT 15.150 33.680 15.490 34.510 ;
        RECT 12.185 32.505 13.395 33.595 ;
        RECT 16.970 32.940 17.320 34.190 ;
        RECT 20.670 33.680 21.010 34.510 ;
        RECT 22.490 32.940 22.840 34.190 ;
        RECT 26.190 33.680 26.530 34.510 ;
        RECT 28.010 32.940 28.360 34.190 ;
        RECT 31.710 33.680 32.050 34.510 ;
        RECT 35.645 34.285 37.315 35.055 ;
        RECT 37.945 34.330 38.235 35.055 ;
        RECT 38.405 34.510 43.750 35.055 ;
        RECT 43.925 34.510 49.270 35.055 ;
        RECT 49.445 34.510 54.790 35.055 ;
        RECT 33.530 32.940 33.880 34.190 ;
        RECT 35.645 33.765 36.395 34.285 ;
        RECT 36.565 33.595 37.315 34.115 ;
        RECT 39.990 33.680 40.330 34.510 ;
        RECT 13.565 32.505 18.910 32.940 ;
        RECT 19.085 32.505 24.430 32.940 ;
        RECT 24.605 32.505 29.950 32.940 ;
        RECT 30.125 32.505 35.470 32.940 ;
        RECT 35.645 32.505 37.315 33.595 ;
        RECT 37.945 32.505 38.235 33.670 ;
        RECT 41.810 32.940 42.160 34.190 ;
        RECT 45.510 33.680 45.850 34.510 ;
        RECT 47.330 32.940 47.680 34.190 ;
        RECT 51.030 33.680 51.370 34.510 ;
        RECT 54.965 34.305 56.175 35.055 ;
        RECT 52.850 32.940 53.200 34.190 ;
        RECT 54.965 33.765 55.485 34.305 ;
        RECT 56.345 34.255 57.040 34.885 ;
        RECT 57.245 34.255 57.555 35.055 ;
        RECT 57.760 34.315 58.375 34.885 ;
        RECT 58.545 34.545 58.760 35.055 ;
        RECT 58.990 34.545 59.270 34.875 ;
        RECT 59.450 34.545 59.690 35.055 ;
        RECT 55.655 33.595 56.175 34.135 ;
        RECT 56.365 33.815 56.700 34.065 ;
        RECT 56.870 33.655 57.040 34.255 ;
        RECT 57.210 33.815 57.545 34.085 ;
        RECT 38.405 32.505 43.750 32.940 ;
        RECT 43.925 32.505 49.270 32.940 ;
        RECT 49.445 32.505 54.790 32.940 ;
        RECT 54.965 32.505 56.175 33.595 ;
        RECT 56.345 32.505 56.605 33.645 ;
        RECT 56.775 32.675 57.105 33.655 ;
        RECT 57.275 32.505 57.555 33.645 ;
        RECT 57.760 33.295 58.075 34.315 ;
        RECT 58.245 33.645 58.415 34.145 ;
        RECT 58.665 33.815 58.930 34.375 ;
        RECT 59.100 33.645 59.270 34.545 ;
        RECT 59.440 33.815 59.795 34.375 ;
        RECT 60.485 34.235 60.745 35.055 ;
        RECT 60.915 34.235 61.245 34.655 ;
        RECT 61.425 34.485 61.685 34.885 ;
        RECT 61.855 34.655 62.185 35.055 ;
        RECT 62.355 34.485 62.525 34.835 ;
        RECT 62.695 34.655 63.070 35.055 ;
        RECT 61.425 34.315 63.090 34.485 ;
        RECT 63.260 34.380 63.535 34.725 ;
        RECT 60.995 34.145 61.245 34.235 ;
        RECT 62.920 34.145 63.090 34.315 ;
        RECT 60.490 33.815 60.825 34.065 ;
        RECT 60.995 33.815 61.710 34.145 ;
        RECT 61.925 33.815 62.750 34.145 ;
        RECT 62.920 33.815 63.195 34.145 ;
        RECT 58.245 33.475 59.670 33.645 ;
        RECT 57.760 32.675 58.295 33.295 ;
        RECT 58.465 32.505 58.795 33.305 ;
        RECT 59.280 33.300 59.670 33.475 ;
        RECT 60.485 32.505 60.745 33.645 ;
        RECT 60.995 33.255 61.165 33.815 ;
        RECT 61.425 33.355 61.755 33.645 ;
        RECT 61.925 33.525 62.170 33.815 ;
        RECT 62.920 33.645 63.090 33.815 ;
        RECT 63.365 33.645 63.535 34.380 ;
        RECT 63.705 34.330 63.995 35.055 ;
        RECT 64.630 34.315 64.885 34.885 ;
        RECT 65.055 34.655 65.385 35.055 ;
        RECT 65.810 34.520 66.340 34.885 ;
        RECT 66.530 34.715 66.805 34.885 ;
        RECT 66.525 34.545 66.805 34.715 ;
        RECT 65.810 34.485 65.985 34.520 ;
        RECT 65.055 34.315 65.985 34.485 ;
        RECT 62.430 33.475 63.090 33.645 ;
        RECT 62.430 33.355 62.600 33.475 ;
        RECT 61.425 33.185 62.600 33.355 ;
        RECT 60.985 32.685 62.600 33.015 ;
        RECT 62.770 32.505 63.050 33.305 ;
        RECT 63.260 32.675 63.535 33.645 ;
        RECT 63.705 32.505 63.995 33.670 ;
        RECT 64.630 33.645 64.800 34.315 ;
        RECT 65.055 34.145 65.225 34.315 ;
        RECT 64.970 33.815 65.225 34.145 ;
        RECT 65.450 33.815 65.645 34.145 ;
        RECT 64.630 32.675 64.965 33.645 ;
        RECT 65.135 32.505 65.305 33.645 ;
        RECT 65.475 32.845 65.645 33.815 ;
        RECT 65.815 33.185 65.985 34.315 ;
        RECT 66.155 33.525 66.325 34.325 ;
        RECT 66.530 33.725 66.805 34.545 ;
        RECT 66.975 33.525 67.165 34.885 ;
        RECT 67.345 34.520 67.855 35.055 ;
        RECT 68.075 34.245 68.320 34.850 ;
        RECT 68.770 34.315 69.025 34.885 ;
        RECT 69.195 34.655 69.525 35.055 ;
        RECT 69.950 34.520 70.480 34.885 ;
        RECT 70.670 34.715 70.945 34.885 ;
        RECT 70.665 34.545 70.945 34.715 ;
        RECT 69.950 34.485 70.125 34.520 ;
        RECT 69.195 34.315 70.125 34.485 ;
        RECT 67.365 34.075 68.595 34.245 ;
        RECT 66.155 33.355 67.165 33.525 ;
        RECT 67.335 33.510 68.085 33.700 ;
        RECT 65.815 33.015 66.940 33.185 ;
        RECT 67.335 32.845 67.505 33.510 ;
        RECT 68.255 33.265 68.595 34.075 ;
        RECT 65.475 32.675 67.505 32.845 ;
        RECT 67.675 32.505 67.845 33.265 ;
        RECT 68.080 32.855 68.595 33.265 ;
        RECT 68.770 33.645 68.940 34.315 ;
        RECT 69.195 34.145 69.365 34.315 ;
        RECT 69.110 33.815 69.365 34.145 ;
        RECT 69.590 33.815 69.785 34.145 ;
        RECT 68.770 32.675 69.105 33.645 ;
        RECT 69.275 32.505 69.445 33.645 ;
        RECT 69.615 32.845 69.785 33.815 ;
        RECT 69.955 33.185 70.125 34.315 ;
        RECT 70.295 33.525 70.465 34.325 ;
        RECT 70.670 33.725 70.945 34.545 ;
        RECT 71.115 33.525 71.305 34.885 ;
        RECT 71.485 34.520 71.995 35.055 ;
        RECT 72.215 34.245 72.460 34.850 ;
        RECT 72.905 34.255 73.245 34.885 ;
        RECT 73.415 34.255 73.665 35.055 ;
        RECT 73.855 34.405 74.185 34.885 ;
        RECT 74.355 34.595 74.580 35.055 ;
        RECT 74.750 34.405 75.080 34.885 ;
        RECT 71.505 34.075 72.735 34.245 ;
        RECT 70.295 33.355 71.305 33.525 ;
        RECT 71.475 33.510 72.225 33.700 ;
        RECT 69.955 33.015 71.080 33.185 ;
        RECT 71.475 32.845 71.645 33.510 ;
        RECT 72.395 33.265 72.735 34.075 ;
        RECT 69.615 32.675 71.645 32.845 ;
        RECT 71.815 32.505 71.985 33.265 ;
        RECT 72.220 32.855 72.735 33.265 ;
        RECT 72.905 33.645 73.080 34.255 ;
        RECT 73.855 34.235 75.080 34.405 ;
        RECT 75.710 34.275 76.210 34.885 ;
        RECT 76.585 34.315 76.970 34.885 ;
        RECT 77.140 34.595 77.465 35.055 ;
        RECT 77.985 34.425 78.265 34.885 ;
        RECT 73.250 33.895 73.945 34.065 ;
        RECT 73.775 33.645 73.945 33.895 ;
        RECT 74.120 33.865 74.540 34.065 ;
        RECT 74.710 33.865 75.040 34.065 ;
        RECT 75.210 33.865 75.540 34.065 ;
        RECT 75.710 33.645 75.880 34.275 ;
        RECT 76.065 33.815 76.415 34.065 ;
        RECT 76.585 33.645 76.865 34.315 ;
        RECT 77.140 34.255 78.265 34.425 ;
        RECT 77.140 34.145 77.590 34.255 ;
        RECT 77.035 33.815 77.590 34.145 ;
        RECT 78.455 34.085 78.855 34.885 ;
        RECT 79.255 34.595 79.525 35.055 ;
        RECT 79.695 34.425 79.980 34.885 ;
        RECT 72.905 32.675 73.245 33.645 ;
        RECT 73.415 32.505 73.585 33.645 ;
        RECT 73.775 33.475 76.210 33.645 ;
        RECT 73.855 32.505 74.105 33.305 ;
        RECT 74.750 32.675 75.080 33.475 ;
        RECT 75.380 32.505 75.710 33.305 ;
        RECT 75.880 32.675 76.210 33.475 ;
        RECT 76.585 32.675 76.970 33.645 ;
        RECT 77.140 33.355 77.590 33.815 ;
        RECT 77.760 33.525 78.855 34.085 ;
        RECT 77.140 33.135 78.265 33.355 ;
        RECT 77.140 32.505 77.465 32.965 ;
        RECT 77.985 32.675 78.265 33.135 ;
        RECT 78.455 32.675 78.855 33.525 ;
        RECT 79.025 34.255 79.980 34.425 ;
        RECT 80.265 34.255 80.605 34.885 ;
        RECT 80.775 34.255 81.025 35.055 ;
        RECT 81.215 34.405 81.545 34.885 ;
        RECT 81.715 34.595 81.940 35.055 ;
        RECT 82.110 34.405 82.440 34.885 ;
        RECT 79.025 33.355 79.235 34.255 ;
        RECT 79.405 33.525 80.095 34.085 ;
        RECT 80.265 33.645 80.440 34.255 ;
        RECT 81.215 34.235 82.440 34.405 ;
        RECT 83.070 34.275 83.570 34.885 ;
        RECT 80.610 33.895 81.305 34.065 ;
        RECT 81.135 33.645 81.305 33.895 ;
        RECT 81.480 33.865 81.900 34.065 ;
        RECT 82.070 33.865 82.400 34.065 ;
        RECT 82.570 33.865 82.900 34.065 ;
        RECT 83.070 33.645 83.240 34.275 ;
        RECT 83.945 34.255 84.285 34.885 ;
        RECT 84.455 34.255 84.705 35.055 ;
        RECT 84.895 34.405 85.225 34.885 ;
        RECT 85.395 34.595 85.620 35.055 ;
        RECT 85.790 34.405 86.120 34.885 ;
        RECT 83.425 33.815 83.775 34.065 ;
        RECT 83.945 33.645 84.120 34.255 ;
        RECT 84.895 34.235 86.120 34.405 ;
        RECT 86.750 34.275 87.250 34.885 ;
        RECT 88.545 34.305 89.755 35.055 ;
        RECT 84.290 33.895 84.985 34.065 ;
        RECT 84.815 33.645 84.985 33.895 ;
        RECT 85.160 33.865 85.580 34.065 ;
        RECT 85.750 33.865 86.080 34.065 ;
        RECT 86.250 33.865 86.580 34.065 ;
        RECT 86.750 33.645 86.920 34.275 ;
        RECT 87.105 33.815 87.455 34.065 ;
        RECT 79.025 33.135 79.980 33.355 ;
        RECT 79.255 32.505 79.525 32.965 ;
        RECT 79.695 32.675 79.980 33.135 ;
        RECT 80.265 32.675 80.605 33.645 ;
        RECT 80.775 32.505 80.945 33.645 ;
        RECT 81.135 33.475 83.570 33.645 ;
        RECT 81.215 32.505 81.465 33.305 ;
        RECT 82.110 32.675 82.440 33.475 ;
        RECT 82.740 32.505 83.070 33.305 ;
        RECT 83.240 32.675 83.570 33.475 ;
        RECT 83.945 32.675 84.285 33.645 ;
        RECT 84.455 32.505 84.625 33.645 ;
        RECT 84.815 33.475 87.250 33.645 ;
        RECT 84.895 32.505 85.145 33.305 ;
        RECT 85.790 32.675 86.120 33.475 ;
        RECT 86.420 32.505 86.750 33.305 ;
        RECT 86.920 32.675 87.250 33.475 ;
        RECT 88.545 33.595 89.065 34.135 ;
        RECT 89.235 33.765 89.755 34.305 ;
        RECT 88.545 32.505 89.755 33.595 ;
        RECT 12.100 32.335 89.840 32.505 ;
        RECT 12.185 31.245 13.395 32.335 ;
        RECT 13.565 31.900 18.910 32.335 ;
        RECT 19.085 31.900 24.430 32.335 ;
        RECT 12.185 30.535 12.705 31.075 ;
        RECT 12.875 30.705 13.395 31.245 ;
        RECT 12.185 29.785 13.395 30.535 ;
        RECT 15.150 30.330 15.490 31.160 ;
        RECT 16.970 30.650 17.320 31.900 ;
        RECT 20.670 30.330 21.010 31.160 ;
        RECT 22.490 30.650 22.840 31.900 ;
        RECT 25.065 31.170 25.355 32.335 ;
        RECT 25.525 31.900 30.870 32.335 ;
        RECT 31.045 31.900 36.390 32.335 ;
        RECT 36.565 31.900 41.910 32.335 ;
        RECT 42.085 31.900 47.430 32.335 ;
        RECT 13.565 29.785 18.910 30.330 ;
        RECT 19.085 29.785 24.430 30.330 ;
        RECT 25.065 29.785 25.355 30.510 ;
        RECT 27.110 30.330 27.450 31.160 ;
        RECT 28.930 30.650 29.280 31.900 ;
        RECT 32.630 30.330 32.970 31.160 ;
        RECT 34.450 30.650 34.800 31.900 ;
        RECT 38.150 30.330 38.490 31.160 ;
        RECT 39.970 30.650 40.320 31.900 ;
        RECT 43.670 30.330 44.010 31.160 ;
        RECT 45.490 30.650 45.840 31.900 ;
        RECT 47.605 31.245 50.195 32.335 ;
        RECT 47.605 30.555 48.815 31.075 ;
        RECT 48.985 30.725 50.195 31.245 ;
        RECT 50.825 31.170 51.115 32.335 ;
        RECT 51.290 31.195 51.610 32.335 ;
        RECT 51.790 31.025 51.985 32.075 ;
        RECT 52.165 31.485 52.495 32.165 ;
        RECT 52.695 31.535 52.950 32.335 ;
        RECT 53.325 31.665 53.605 32.335 ;
        RECT 52.165 31.205 52.515 31.485 ;
        RECT 53.775 31.445 54.075 31.995 ;
        RECT 54.275 31.615 54.605 32.335 ;
        RECT 54.795 31.615 55.255 32.165 ;
        RECT 51.350 30.975 51.610 31.025 ;
        RECT 51.345 30.805 51.610 30.975 ;
        RECT 51.350 30.695 51.610 30.805 ;
        RECT 51.790 30.695 52.175 31.025 ;
        RECT 52.345 30.825 52.515 31.205 ;
        RECT 52.705 30.995 52.950 31.355 ;
        RECT 53.140 31.025 53.405 31.385 ;
        RECT 53.775 31.275 54.715 31.445 ;
        RECT 54.545 31.025 54.715 31.275 ;
        RECT 52.345 30.655 52.865 30.825 ;
        RECT 53.140 30.775 53.815 31.025 ;
        RECT 54.035 30.775 54.375 31.025 ;
        RECT 25.525 29.785 30.870 30.330 ;
        RECT 31.045 29.785 36.390 30.330 ;
        RECT 36.565 29.785 41.910 30.330 ;
        RECT 42.085 29.785 47.430 30.330 ;
        RECT 47.605 29.785 50.195 30.555 ;
        RECT 50.825 29.785 51.115 30.510 ;
        RECT 51.290 30.315 52.505 30.485 ;
        RECT 51.290 29.965 51.580 30.315 ;
        RECT 51.775 29.785 52.105 30.145 ;
        RECT 52.275 30.010 52.505 30.315 ;
        RECT 52.695 30.295 52.865 30.655 ;
        RECT 54.545 30.695 54.835 31.025 ;
        RECT 54.545 30.605 54.715 30.695 ;
        RECT 53.325 30.415 54.715 30.605 ;
        RECT 52.695 30.125 52.895 30.295 ;
        RECT 52.695 30.090 52.865 30.125 ;
        RECT 53.325 30.055 53.655 30.415 ;
        RECT 55.005 30.245 55.255 31.615 ;
        RECT 55.515 31.665 55.685 32.165 ;
        RECT 55.855 31.835 56.185 32.335 ;
        RECT 55.515 31.495 56.180 31.665 ;
        RECT 55.430 30.675 55.780 31.325 ;
        RECT 55.950 30.505 56.180 31.495 ;
        RECT 54.275 29.785 54.525 30.245 ;
        RECT 54.695 29.955 55.255 30.245 ;
        RECT 55.515 30.335 56.180 30.505 ;
        RECT 55.515 30.045 55.685 30.335 ;
        RECT 55.855 29.785 56.185 30.165 ;
        RECT 56.355 30.045 56.540 32.165 ;
        RECT 56.780 31.875 57.045 32.335 ;
        RECT 57.215 31.740 57.465 32.165 ;
        RECT 57.675 31.890 58.780 32.060 ;
        RECT 57.160 31.610 57.465 31.740 ;
        RECT 56.710 30.415 56.990 31.365 ;
        RECT 57.160 30.505 57.330 31.610 ;
        RECT 57.500 30.825 57.740 31.420 ;
        RECT 57.910 31.355 58.440 31.720 ;
        RECT 57.910 30.655 58.080 31.355 ;
        RECT 58.610 31.275 58.780 31.890 ;
        RECT 58.950 31.535 59.120 32.335 ;
        RECT 59.290 31.835 59.540 32.165 ;
        RECT 59.765 31.865 60.650 32.035 ;
        RECT 58.610 31.185 59.120 31.275 ;
        RECT 57.160 30.375 57.385 30.505 ;
        RECT 57.555 30.435 58.080 30.655 ;
        RECT 58.250 31.015 59.120 31.185 ;
        RECT 56.795 29.785 57.045 30.245 ;
        RECT 57.215 30.235 57.385 30.375 ;
        RECT 58.250 30.235 58.420 31.015 ;
        RECT 58.950 30.945 59.120 31.015 ;
        RECT 58.630 30.765 58.830 30.795 ;
        RECT 59.290 30.765 59.460 31.835 ;
        RECT 59.630 30.945 59.820 31.665 ;
        RECT 58.630 30.465 59.460 30.765 ;
        RECT 59.990 30.735 60.310 31.695 ;
        RECT 57.215 30.065 57.550 30.235 ;
        RECT 57.745 30.065 58.420 30.235 ;
        RECT 58.740 29.785 59.110 30.285 ;
        RECT 59.290 30.235 59.460 30.465 ;
        RECT 59.845 30.405 60.310 30.735 ;
        RECT 60.480 31.025 60.650 31.865 ;
        RECT 60.830 31.835 61.145 32.335 ;
        RECT 61.375 31.605 61.715 32.165 ;
        RECT 60.820 31.230 61.715 31.605 ;
        RECT 61.885 31.325 62.055 32.335 ;
        RECT 61.525 31.025 61.715 31.230 ;
        RECT 62.225 31.275 62.555 32.120 ;
        RECT 63.795 31.665 63.965 32.165 ;
        RECT 64.135 31.835 64.465 32.335 ;
        RECT 63.795 31.495 64.460 31.665 ;
        RECT 62.225 31.195 62.615 31.275 ;
        RECT 62.400 31.145 62.615 31.195 ;
        RECT 60.480 30.695 61.355 31.025 ;
        RECT 61.525 30.695 62.275 31.025 ;
        RECT 60.480 30.235 60.650 30.695 ;
        RECT 61.525 30.525 61.725 30.695 ;
        RECT 62.445 30.565 62.615 31.145 ;
        RECT 63.710 30.675 64.060 31.325 ;
        RECT 62.390 30.525 62.615 30.565 ;
        RECT 59.290 30.065 59.695 30.235 ;
        RECT 59.865 30.065 60.650 30.235 ;
        RECT 60.925 29.785 61.135 30.315 ;
        RECT 61.395 30.000 61.725 30.525 ;
        RECT 62.235 30.440 62.615 30.525 ;
        RECT 64.230 30.505 64.460 31.495 ;
        RECT 61.895 29.785 62.065 30.395 ;
        RECT 62.235 30.005 62.565 30.440 ;
        RECT 63.795 30.335 64.460 30.505 ;
        RECT 63.795 30.045 63.965 30.335 ;
        RECT 64.135 29.785 64.465 30.165 ;
        RECT 64.635 30.045 64.820 32.165 ;
        RECT 65.060 31.875 65.325 32.335 ;
        RECT 65.495 31.740 65.745 32.165 ;
        RECT 65.955 31.890 67.060 32.060 ;
        RECT 65.440 31.610 65.745 31.740 ;
        RECT 64.990 30.415 65.270 31.365 ;
        RECT 65.440 30.505 65.610 31.610 ;
        RECT 65.780 30.825 66.020 31.420 ;
        RECT 66.190 31.355 66.720 31.720 ;
        RECT 66.190 30.655 66.360 31.355 ;
        RECT 66.890 31.275 67.060 31.890 ;
        RECT 67.230 31.535 67.400 32.335 ;
        RECT 67.570 31.835 67.820 32.165 ;
        RECT 68.045 31.865 68.930 32.035 ;
        RECT 66.890 31.185 67.400 31.275 ;
        RECT 65.440 30.375 65.665 30.505 ;
        RECT 65.835 30.435 66.360 30.655 ;
        RECT 66.530 31.015 67.400 31.185 ;
        RECT 65.075 29.785 65.325 30.245 ;
        RECT 65.495 30.235 65.665 30.375 ;
        RECT 66.530 30.235 66.700 31.015 ;
        RECT 67.230 30.945 67.400 31.015 ;
        RECT 66.910 30.765 67.110 30.795 ;
        RECT 67.570 30.765 67.740 31.835 ;
        RECT 67.910 30.945 68.100 31.665 ;
        RECT 66.910 30.465 67.740 30.765 ;
        RECT 68.270 30.735 68.590 31.695 ;
        RECT 65.495 30.065 65.830 30.235 ;
        RECT 66.025 30.065 66.700 30.235 ;
        RECT 67.020 29.785 67.390 30.285 ;
        RECT 67.570 30.235 67.740 30.465 ;
        RECT 68.125 30.405 68.590 30.735 ;
        RECT 68.760 31.025 68.930 31.865 ;
        RECT 69.110 31.835 69.425 32.335 ;
        RECT 69.655 31.605 69.995 32.165 ;
        RECT 69.100 31.230 69.995 31.605 ;
        RECT 70.165 31.325 70.335 32.335 ;
        RECT 69.805 31.025 69.995 31.230 ;
        RECT 70.505 31.275 70.835 32.120 ;
        RECT 71.005 31.420 71.175 32.335 ;
        RECT 70.505 31.195 70.895 31.275 ;
        RECT 70.680 31.145 70.895 31.195 ;
        RECT 68.760 30.695 69.635 31.025 ;
        RECT 69.805 30.695 70.555 31.025 ;
        RECT 68.760 30.235 68.930 30.695 ;
        RECT 69.805 30.525 70.005 30.695 ;
        RECT 70.725 30.565 70.895 31.145 ;
        RECT 70.670 30.525 70.895 30.565 ;
        RECT 67.570 30.065 67.975 30.235 ;
        RECT 68.145 30.065 68.930 30.235 ;
        RECT 69.205 29.785 69.415 30.315 ;
        RECT 69.675 30.000 70.005 30.525 ;
        RECT 70.515 30.440 70.895 30.525 ;
        RECT 71.530 31.195 71.865 32.165 ;
        RECT 72.035 31.195 72.205 32.335 ;
        RECT 72.375 31.995 74.405 32.165 ;
        RECT 71.530 30.525 71.700 31.195 ;
        RECT 72.375 31.025 72.545 31.995 ;
        RECT 71.870 30.695 72.125 31.025 ;
        RECT 72.350 30.695 72.545 31.025 ;
        RECT 72.715 31.655 73.840 31.825 ;
        RECT 71.955 30.525 72.125 30.695 ;
        RECT 72.715 30.525 72.885 31.655 ;
        RECT 70.175 29.785 70.345 30.395 ;
        RECT 70.515 30.005 70.845 30.440 ;
        RECT 71.015 29.785 71.185 30.300 ;
        RECT 71.530 29.955 71.785 30.525 ;
        RECT 71.955 30.355 72.885 30.525 ;
        RECT 73.055 31.315 74.065 31.485 ;
        RECT 73.055 30.515 73.225 31.315 ;
        RECT 73.430 30.635 73.705 31.115 ;
        RECT 73.425 30.465 73.705 30.635 ;
        RECT 72.710 30.320 72.885 30.355 ;
        RECT 71.955 29.785 72.285 30.185 ;
        RECT 72.710 29.955 73.240 30.320 ;
        RECT 73.430 29.955 73.705 30.465 ;
        RECT 73.875 29.955 74.065 31.315 ;
        RECT 74.235 31.330 74.405 31.995 ;
        RECT 74.575 31.575 74.745 32.335 ;
        RECT 74.980 31.575 75.495 31.985 ;
        RECT 74.235 31.140 74.985 31.330 ;
        RECT 75.155 30.765 75.495 31.575 ;
        RECT 76.585 31.170 76.875 32.335 ;
        RECT 77.105 31.275 77.435 32.120 ;
        RECT 77.605 31.325 77.775 32.335 ;
        RECT 77.945 31.605 78.285 32.165 ;
        RECT 78.515 31.835 78.830 32.335 ;
        RECT 79.010 31.865 79.895 32.035 ;
        RECT 77.045 31.195 77.435 31.275 ;
        RECT 77.945 31.230 78.840 31.605 ;
        RECT 74.265 30.595 75.495 30.765 ;
        RECT 77.045 31.145 77.260 31.195 ;
        RECT 74.245 29.785 74.755 30.320 ;
        RECT 74.975 29.990 75.220 30.595 ;
        RECT 77.045 30.565 77.215 31.145 ;
        RECT 77.945 31.025 78.135 31.230 ;
        RECT 79.010 31.025 79.180 31.865 ;
        RECT 80.120 31.835 80.370 32.165 ;
        RECT 77.385 30.695 78.135 31.025 ;
        RECT 78.305 30.695 79.180 31.025 ;
        RECT 77.045 30.525 77.270 30.565 ;
        RECT 77.935 30.525 78.135 30.695 ;
        RECT 76.585 29.785 76.875 30.510 ;
        RECT 77.045 30.440 77.425 30.525 ;
        RECT 77.095 30.005 77.425 30.440 ;
        RECT 77.595 29.785 77.765 30.395 ;
        RECT 77.935 30.000 78.265 30.525 ;
        RECT 78.525 29.785 78.735 30.315 ;
        RECT 79.010 30.235 79.180 30.695 ;
        RECT 79.350 30.735 79.670 31.695 ;
        RECT 79.840 30.945 80.030 31.665 ;
        RECT 80.200 30.765 80.370 31.835 ;
        RECT 80.540 31.535 80.710 32.335 ;
        RECT 80.880 31.890 81.985 32.060 ;
        RECT 80.880 31.275 81.050 31.890 ;
        RECT 82.195 31.740 82.445 32.165 ;
        RECT 82.615 31.875 82.880 32.335 ;
        RECT 81.220 31.355 81.750 31.720 ;
        RECT 82.195 31.610 82.500 31.740 ;
        RECT 80.540 31.185 81.050 31.275 ;
        RECT 80.540 31.015 81.410 31.185 ;
        RECT 80.540 30.945 80.710 31.015 ;
        RECT 80.830 30.765 81.030 30.795 ;
        RECT 79.350 30.405 79.815 30.735 ;
        RECT 80.200 30.465 81.030 30.765 ;
        RECT 80.200 30.235 80.370 30.465 ;
        RECT 79.010 30.065 79.795 30.235 ;
        RECT 79.965 30.065 80.370 30.235 ;
        RECT 80.550 29.785 80.920 30.285 ;
        RECT 81.240 30.235 81.410 31.015 ;
        RECT 81.580 30.655 81.750 31.355 ;
        RECT 81.920 30.825 82.160 31.420 ;
        RECT 81.580 30.435 82.105 30.655 ;
        RECT 82.330 30.505 82.500 31.610 ;
        RECT 82.275 30.375 82.500 30.505 ;
        RECT 82.670 30.415 82.950 31.365 ;
        RECT 82.275 30.235 82.445 30.375 ;
        RECT 81.240 30.065 81.915 30.235 ;
        RECT 82.110 30.065 82.445 30.235 ;
        RECT 82.615 29.785 82.865 30.245 ;
        RECT 83.120 30.045 83.305 32.165 ;
        RECT 83.475 31.835 83.805 32.335 ;
        RECT 83.975 31.665 84.145 32.165 ;
        RECT 83.480 31.495 84.145 31.665 ;
        RECT 83.480 30.505 83.710 31.495 ;
        RECT 83.880 30.675 84.230 31.325 ;
        RECT 84.405 31.195 84.745 32.165 ;
        RECT 84.915 31.195 85.085 32.335 ;
        RECT 85.355 31.535 85.605 32.335 ;
        RECT 86.250 31.365 86.580 32.165 ;
        RECT 86.880 31.535 87.210 32.335 ;
        RECT 87.380 31.365 87.710 32.165 ;
        RECT 85.275 31.195 87.710 31.365 ;
        RECT 88.545 31.245 89.755 32.335 ;
        RECT 84.405 30.585 84.580 31.195 ;
        RECT 85.275 30.945 85.445 31.195 ;
        RECT 84.750 30.775 85.445 30.945 ;
        RECT 85.620 30.775 86.040 30.975 ;
        RECT 86.210 30.775 86.540 30.975 ;
        RECT 86.710 30.775 87.040 30.975 ;
        RECT 83.480 30.335 84.145 30.505 ;
        RECT 83.475 29.785 83.805 30.165 ;
        RECT 83.975 30.045 84.145 30.335 ;
        RECT 84.405 29.955 84.745 30.585 ;
        RECT 84.915 29.785 85.165 30.585 ;
        RECT 85.355 30.435 86.580 30.605 ;
        RECT 85.355 29.955 85.685 30.435 ;
        RECT 85.855 29.785 86.080 30.245 ;
        RECT 86.250 29.955 86.580 30.435 ;
        RECT 87.210 30.565 87.380 31.195 ;
        RECT 87.565 30.775 87.915 31.025 ;
        RECT 88.545 30.705 89.065 31.245 ;
        RECT 87.210 29.955 87.710 30.565 ;
        RECT 89.235 30.535 89.755 31.075 ;
        RECT 88.545 29.785 89.755 30.535 ;
        RECT 12.100 29.615 89.840 29.785 ;
        RECT 12.185 28.865 13.395 29.615 ;
        RECT 13.565 29.070 18.910 29.615 ;
        RECT 19.085 29.070 24.430 29.615 ;
        RECT 24.605 29.070 29.950 29.615 ;
        RECT 30.125 29.070 35.470 29.615 ;
        RECT 12.185 28.325 12.705 28.865 ;
        RECT 12.875 28.155 13.395 28.695 ;
        RECT 15.150 28.240 15.490 29.070 ;
        RECT 12.185 27.065 13.395 28.155 ;
        RECT 16.970 27.500 17.320 28.750 ;
        RECT 20.670 28.240 21.010 29.070 ;
        RECT 22.490 27.500 22.840 28.750 ;
        RECT 26.190 28.240 26.530 29.070 ;
        RECT 28.010 27.500 28.360 28.750 ;
        RECT 31.710 28.240 32.050 29.070 ;
        RECT 35.645 28.845 37.315 29.615 ;
        RECT 37.945 28.890 38.235 29.615 ;
        RECT 38.405 29.070 43.750 29.615 ;
        RECT 33.530 27.500 33.880 28.750 ;
        RECT 35.645 28.325 36.395 28.845 ;
        RECT 36.565 28.155 37.315 28.675 ;
        RECT 39.990 28.240 40.330 29.070 ;
        RECT 43.925 28.845 46.515 29.615 ;
        RECT 46.720 28.875 47.335 29.445 ;
        RECT 47.505 29.105 47.720 29.615 ;
        RECT 47.950 29.105 48.230 29.435 ;
        RECT 48.410 29.105 48.650 29.615 ;
        RECT 48.985 29.155 49.545 29.445 ;
        RECT 49.715 29.155 49.965 29.615 ;
        RECT 13.565 27.065 18.910 27.500 ;
        RECT 19.085 27.065 24.430 27.500 ;
        RECT 24.605 27.065 29.950 27.500 ;
        RECT 30.125 27.065 35.470 27.500 ;
        RECT 35.645 27.065 37.315 28.155 ;
        RECT 37.945 27.065 38.235 28.230 ;
        RECT 41.810 27.500 42.160 28.750 ;
        RECT 43.925 28.325 45.135 28.845 ;
        RECT 45.305 28.155 46.515 28.675 ;
        RECT 38.405 27.065 43.750 27.500 ;
        RECT 43.925 27.065 46.515 28.155 ;
        RECT 46.720 27.855 47.035 28.875 ;
        RECT 47.205 28.205 47.375 28.705 ;
        RECT 47.625 28.375 47.890 28.935 ;
        RECT 48.060 28.205 48.230 29.105 ;
        RECT 48.400 28.375 48.755 28.935 ;
        RECT 47.205 28.035 48.630 28.205 ;
        RECT 46.720 27.235 47.255 27.855 ;
        RECT 47.425 27.065 47.755 27.865 ;
        RECT 48.240 27.860 48.630 28.035 ;
        RECT 48.985 27.785 49.235 29.155 ;
        RECT 50.585 28.985 50.915 29.345 ;
        RECT 49.525 28.795 50.915 28.985 ;
        RECT 51.290 29.140 51.625 29.400 ;
        RECT 51.795 29.215 52.125 29.615 ;
        RECT 52.295 29.215 53.910 29.385 ;
        RECT 49.525 28.705 49.695 28.795 ;
        RECT 49.405 28.375 49.695 28.705 ;
        RECT 49.865 28.375 50.205 28.625 ;
        RECT 50.425 28.375 51.100 28.625 ;
        RECT 49.525 28.125 49.695 28.375 ;
        RECT 49.525 27.955 50.465 28.125 ;
        RECT 50.835 28.015 51.100 28.375 ;
        RECT 48.985 27.235 49.445 27.785 ;
        RECT 49.635 27.065 49.965 27.785 ;
        RECT 50.165 27.405 50.465 27.955 ;
        RECT 51.290 27.785 51.545 29.140 ;
        RECT 52.295 29.045 52.465 29.215 ;
        RECT 51.905 28.875 52.465 29.045 ;
        RECT 52.730 28.935 53.000 29.035 ;
        RECT 53.190 28.935 53.480 29.035 ;
        RECT 51.905 28.705 52.075 28.875 ;
        RECT 52.725 28.765 53.000 28.935 ;
        RECT 53.185 28.765 53.480 28.935 ;
        RECT 51.770 28.375 52.075 28.705 ;
        RECT 52.270 28.595 52.520 28.705 ;
        RECT 52.265 28.425 52.520 28.595 ;
        RECT 52.270 28.375 52.520 28.425 ;
        RECT 52.730 28.375 53.000 28.765 ;
        RECT 53.190 28.375 53.480 28.765 ;
        RECT 53.650 28.375 54.070 29.040 ;
        RECT 54.455 28.895 54.785 29.615 ;
        RECT 55.975 29.065 56.145 29.355 ;
        RECT 56.315 29.235 56.645 29.615 ;
        RECT 55.975 28.895 56.640 29.065 ;
        RECT 54.380 28.595 54.730 28.705 ;
        RECT 54.380 28.425 54.735 28.595 ;
        RECT 54.380 28.375 54.730 28.425 ;
        RECT 51.905 28.205 52.075 28.375 ;
        RECT 51.905 28.035 54.275 28.205 ;
        RECT 54.525 28.085 54.730 28.375 ;
        RECT 55.890 28.075 56.240 28.725 ;
        RECT 50.635 27.065 50.915 27.735 ;
        RECT 51.290 27.275 51.625 27.785 ;
        RECT 51.875 27.065 52.205 27.865 ;
        RECT 52.450 27.655 53.875 27.825 ;
        RECT 52.450 27.235 52.735 27.655 ;
        RECT 52.990 27.065 53.320 27.485 ;
        RECT 53.545 27.405 53.875 27.655 ;
        RECT 54.105 27.575 54.275 28.035 ;
        RECT 56.410 27.905 56.640 28.895 ;
        RECT 54.535 27.405 54.705 27.905 ;
        RECT 53.545 27.235 54.705 27.405 ;
        RECT 55.975 27.735 56.640 27.905 ;
        RECT 55.975 27.235 56.145 27.735 ;
        RECT 56.315 27.065 56.645 27.565 ;
        RECT 56.815 27.235 57.000 29.355 ;
        RECT 57.255 29.155 57.505 29.615 ;
        RECT 57.675 29.165 58.010 29.335 ;
        RECT 58.205 29.165 58.880 29.335 ;
        RECT 57.675 29.025 57.845 29.165 ;
        RECT 57.170 28.035 57.450 28.985 ;
        RECT 57.620 28.895 57.845 29.025 ;
        RECT 57.620 27.790 57.790 28.895 ;
        RECT 58.015 28.745 58.540 28.965 ;
        RECT 57.960 27.980 58.200 28.575 ;
        RECT 58.370 28.045 58.540 28.745 ;
        RECT 58.710 28.385 58.880 29.165 ;
        RECT 59.200 29.115 59.570 29.615 ;
        RECT 59.750 29.165 60.155 29.335 ;
        RECT 60.325 29.165 61.110 29.335 ;
        RECT 59.750 28.935 59.920 29.165 ;
        RECT 59.090 28.635 59.920 28.935 ;
        RECT 60.305 28.665 60.770 28.995 ;
        RECT 59.090 28.605 59.290 28.635 ;
        RECT 59.410 28.385 59.580 28.455 ;
        RECT 58.710 28.215 59.580 28.385 ;
        RECT 59.070 28.125 59.580 28.215 ;
        RECT 57.620 27.660 57.925 27.790 ;
        RECT 58.370 27.680 58.900 28.045 ;
        RECT 57.240 27.065 57.505 27.525 ;
        RECT 57.675 27.235 57.925 27.660 ;
        RECT 59.070 27.510 59.240 28.125 ;
        RECT 58.135 27.340 59.240 27.510 ;
        RECT 59.410 27.065 59.580 27.865 ;
        RECT 59.750 27.565 59.920 28.635 ;
        RECT 60.090 27.735 60.280 28.455 ;
        RECT 60.450 27.705 60.770 28.665 ;
        RECT 60.940 28.705 61.110 29.165 ;
        RECT 61.385 29.085 61.595 29.615 ;
        RECT 61.855 28.875 62.185 29.400 ;
        RECT 62.355 29.005 62.525 29.615 ;
        RECT 62.695 28.960 63.025 29.395 ;
        RECT 63.195 29.100 63.365 29.615 ;
        RECT 62.695 28.875 63.075 28.960 ;
        RECT 63.705 28.890 63.995 29.615 ;
        RECT 64.335 29.100 64.505 29.615 ;
        RECT 64.675 28.960 65.005 29.395 ;
        RECT 65.175 29.005 65.345 29.615 ;
        RECT 61.985 28.705 62.185 28.875 ;
        RECT 62.850 28.835 63.075 28.875 ;
        RECT 60.940 28.375 61.815 28.705 ;
        RECT 61.985 28.375 62.735 28.705 ;
        RECT 59.750 27.235 60.000 27.565 ;
        RECT 60.940 27.535 61.110 28.375 ;
        RECT 61.985 28.170 62.175 28.375 ;
        RECT 62.905 28.255 63.075 28.835 ;
        RECT 62.860 28.205 63.075 28.255 ;
        RECT 64.625 28.875 65.005 28.960 ;
        RECT 65.515 28.875 65.845 29.400 ;
        RECT 66.105 29.085 66.315 29.615 ;
        RECT 66.590 29.165 67.375 29.335 ;
        RECT 67.545 29.165 67.950 29.335 ;
        RECT 64.625 28.835 64.850 28.875 ;
        RECT 64.625 28.255 64.795 28.835 ;
        RECT 65.515 28.705 65.715 28.875 ;
        RECT 66.590 28.705 66.760 29.165 ;
        RECT 64.965 28.375 65.715 28.705 ;
        RECT 65.885 28.375 66.760 28.705 ;
        RECT 61.280 27.795 62.175 28.170 ;
        RECT 62.685 28.125 63.075 28.205 ;
        RECT 60.225 27.365 61.110 27.535 ;
        RECT 61.290 27.065 61.605 27.565 ;
        RECT 61.835 27.235 62.175 27.795 ;
        RECT 62.345 27.065 62.515 28.075 ;
        RECT 62.685 27.280 63.015 28.125 ;
        RECT 63.185 27.065 63.355 27.980 ;
        RECT 63.705 27.065 63.995 28.230 ;
        RECT 64.625 28.205 64.840 28.255 ;
        RECT 64.625 28.125 65.015 28.205 ;
        RECT 64.345 27.065 64.515 27.980 ;
        RECT 64.685 27.280 65.015 28.125 ;
        RECT 65.525 28.170 65.715 28.375 ;
        RECT 65.185 27.065 65.355 28.075 ;
        RECT 65.525 27.795 66.420 28.170 ;
        RECT 65.525 27.235 65.865 27.795 ;
        RECT 66.095 27.065 66.410 27.565 ;
        RECT 66.590 27.535 66.760 28.375 ;
        RECT 66.930 28.665 67.395 28.995 ;
        RECT 67.780 28.935 67.950 29.165 ;
        RECT 68.130 29.115 68.500 29.615 ;
        RECT 68.820 29.165 69.495 29.335 ;
        RECT 69.690 29.165 70.025 29.335 ;
        RECT 66.930 27.705 67.250 28.665 ;
        RECT 67.780 28.635 68.610 28.935 ;
        RECT 67.420 27.735 67.610 28.455 ;
        RECT 67.780 27.565 67.950 28.635 ;
        RECT 68.410 28.605 68.610 28.635 ;
        RECT 68.120 28.385 68.290 28.455 ;
        RECT 68.820 28.385 68.990 29.165 ;
        RECT 69.855 29.025 70.025 29.165 ;
        RECT 70.195 29.155 70.445 29.615 ;
        RECT 68.120 28.215 68.990 28.385 ;
        RECT 69.160 28.745 69.685 28.965 ;
        RECT 69.855 28.895 70.080 29.025 ;
        RECT 68.120 28.125 68.630 28.215 ;
        RECT 66.590 27.365 67.475 27.535 ;
        RECT 67.700 27.235 67.950 27.565 ;
        RECT 68.120 27.065 68.290 27.865 ;
        RECT 68.460 27.510 68.630 28.125 ;
        RECT 69.160 28.045 69.330 28.745 ;
        RECT 68.800 27.680 69.330 28.045 ;
        RECT 69.500 27.980 69.740 28.575 ;
        RECT 69.910 27.790 70.080 28.895 ;
        RECT 70.250 28.035 70.530 28.985 ;
        RECT 69.775 27.660 70.080 27.790 ;
        RECT 68.460 27.340 69.565 27.510 ;
        RECT 69.775 27.235 70.025 27.660 ;
        RECT 70.195 27.065 70.460 27.525 ;
        RECT 70.700 27.235 70.885 29.355 ;
        RECT 71.055 29.235 71.385 29.615 ;
        RECT 71.555 29.065 71.725 29.355 ;
        RECT 71.060 28.895 71.725 29.065 ;
        RECT 72.075 29.065 72.245 29.355 ;
        RECT 72.415 29.235 72.745 29.615 ;
        RECT 72.075 28.895 72.740 29.065 ;
        RECT 71.060 27.905 71.290 28.895 ;
        RECT 71.460 28.075 71.810 28.725 ;
        RECT 71.990 28.075 72.340 28.725 ;
        RECT 72.510 27.905 72.740 28.895 ;
        RECT 71.060 27.735 71.725 27.905 ;
        RECT 71.055 27.065 71.385 27.565 ;
        RECT 71.555 27.235 71.725 27.735 ;
        RECT 72.075 27.735 72.740 27.905 ;
        RECT 72.075 27.235 72.245 27.735 ;
        RECT 72.415 27.065 72.745 27.565 ;
        RECT 72.915 27.235 73.100 29.355 ;
        RECT 73.355 29.155 73.605 29.615 ;
        RECT 73.775 29.165 74.110 29.335 ;
        RECT 74.305 29.165 74.980 29.335 ;
        RECT 73.775 29.025 73.945 29.165 ;
        RECT 73.270 28.035 73.550 28.985 ;
        RECT 73.720 28.895 73.945 29.025 ;
        RECT 73.720 27.790 73.890 28.895 ;
        RECT 74.115 28.745 74.640 28.965 ;
        RECT 74.060 27.980 74.300 28.575 ;
        RECT 74.470 28.045 74.640 28.745 ;
        RECT 74.810 28.385 74.980 29.165 ;
        RECT 75.300 29.115 75.670 29.615 ;
        RECT 75.850 29.165 76.255 29.335 ;
        RECT 76.425 29.165 77.210 29.335 ;
        RECT 75.850 28.935 76.020 29.165 ;
        RECT 75.190 28.635 76.020 28.935 ;
        RECT 76.405 28.665 76.870 28.995 ;
        RECT 75.190 28.605 75.390 28.635 ;
        RECT 75.510 28.385 75.680 28.455 ;
        RECT 74.810 28.215 75.680 28.385 ;
        RECT 75.170 28.125 75.680 28.215 ;
        RECT 73.720 27.660 74.025 27.790 ;
        RECT 74.470 27.680 75.000 28.045 ;
        RECT 73.340 27.065 73.605 27.525 ;
        RECT 73.775 27.235 74.025 27.660 ;
        RECT 75.170 27.510 75.340 28.125 ;
        RECT 74.235 27.340 75.340 27.510 ;
        RECT 75.510 27.065 75.680 27.865 ;
        RECT 75.850 27.565 76.020 28.635 ;
        RECT 76.190 27.735 76.380 28.455 ;
        RECT 76.550 27.705 76.870 28.665 ;
        RECT 77.040 28.705 77.210 29.165 ;
        RECT 77.485 29.085 77.695 29.615 ;
        RECT 77.955 28.875 78.285 29.400 ;
        RECT 78.455 29.005 78.625 29.615 ;
        RECT 78.795 28.960 79.125 29.395 ;
        RECT 79.855 28.960 80.185 29.395 ;
        RECT 80.355 29.005 80.525 29.615 ;
        RECT 78.795 28.875 79.175 28.960 ;
        RECT 78.085 28.705 78.285 28.875 ;
        RECT 78.950 28.835 79.175 28.875 ;
        RECT 77.040 28.375 77.915 28.705 ;
        RECT 78.085 28.375 78.835 28.705 ;
        RECT 75.850 27.235 76.100 27.565 ;
        RECT 77.040 27.535 77.210 28.375 ;
        RECT 78.085 28.170 78.275 28.375 ;
        RECT 79.005 28.255 79.175 28.835 ;
        RECT 78.960 28.205 79.175 28.255 ;
        RECT 77.380 27.795 78.275 28.170 ;
        RECT 78.785 28.125 79.175 28.205 ;
        RECT 79.805 28.875 80.185 28.960 ;
        RECT 80.695 28.875 81.025 29.400 ;
        RECT 81.285 29.085 81.495 29.615 ;
        RECT 81.770 29.165 82.555 29.335 ;
        RECT 82.725 29.165 83.130 29.335 ;
        RECT 79.805 28.835 80.030 28.875 ;
        RECT 79.805 28.255 79.975 28.835 ;
        RECT 80.695 28.705 80.895 28.875 ;
        RECT 81.770 28.705 81.940 29.165 ;
        RECT 80.145 28.375 80.895 28.705 ;
        RECT 81.065 28.375 81.940 28.705 ;
        RECT 79.805 28.205 80.020 28.255 ;
        RECT 79.805 28.125 80.195 28.205 ;
        RECT 76.325 27.365 77.210 27.535 ;
        RECT 77.390 27.065 77.705 27.565 ;
        RECT 77.935 27.235 78.275 27.795 ;
        RECT 78.445 27.065 78.615 28.075 ;
        RECT 78.785 27.280 79.115 28.125 ;
        RECT 79.865 27.280 80.195 28.125 ;
        RECT 80.705 28.170 80.895 28.375 ;
        RECT 80.365 27.065 80.535 28.075 ;
        RECT 80.705 27.795 81.600 28.170 ;
        RECT 80.705 27.235 81.045 27.795 ;
        RECT 81.275 27.065 81.590 27.565 ;
        RECT 81.770 27.535 81.940 28.375 ;
        RECT 82.110 28.665 82.575 28.995 ;
        RECT 82.960 28.935 83.130 29.165 ;
        RECT 83.310 29.115 83.680 29.615 ;
        RECT 84.000 29.165 84.675 29.335 ;
        RECT 84.870 29.165 85.205 29.335 ;
        RECT 82.110 27.705 82.430 28.665 ;
        RECT 82.960 28.635 83.790 28.935 ;
        RECT 82.600 27.735 82.790 28.455 ;
        RECT 82.960 27.565 83.130 28.635 ;
        RECT 83.590 28.605 83.790 28.635 ;
        RECT 83.300 28.385 83.470 28.455 ;
        RECT 84.000 28.385 84.170 29.165 ;
        RECT 85.035 29.025 85.205 29.165 ;
        RECT 85.375 29.155 85.625 29.615 ;
        RECT 83.300 28.215 84.170 28.385 ;
        RECT 84.340 28.745 84.865 28.965 ;
        RECT 85.035 28.895 85.260 29.025 ;
        RECT 83.300 28.125 83.810 28.215 ;
        RECT 81.770 27.365 82.655 27.535 ;
        RECT 82.880 27.235 83.130 27.565 ;
        RECT 83.300 27.065 83.470 27.865 ;
        RECT 83.640 27.510 83.810 28.125 ;
        RECT 84.340 28.045 84.510 28.745 ;
        RECT 83.980 27.680 84.510 28.045 ;
        RECT 84.680 27.980 84.920 28.575 ;
        RECT 85.090 27.790 85.260 28.895 ;
        RECT 85.430 28.035 85.710 28.985 ;
        RECT 84.955 27.660 85.260 27.790 ;
        RECT 83.640 27.340 84.745 27.510 ;
        RECT 84.955 27.235 85.205 27.660 ;
        RECT 85.375 27.065 85.640 27.525 ;
        RECT 85.880 27.235 86.065 29.355 ;
        RECT 86.235 29.235 86.565 29.615 ;
        RECT 86.735 29.065 86.905 29.355 ;
        RECT 86.240 28.895 86.905 29.065 ;
        RECT 86.240 27.905 86.470 28.895 ;
        RECT 87.165 28.865 88.375 29.615 ;
        RECT 88.545 28.865 89.755 29.615 ;
        RECT 86.640 28.075 86.990 28.725 ;
        RECT 87.165 28.325 87.685 28.865 ;
        RECT 87.855 28.155 88.375 28.695 ;
        RECT 86.240 27.735 86.905 27.905 ;
        RECT 86.235 27.065 86.565 27.565 ;
        RECT 86.735 27.235 86.905 27.735 ;
        RECT 87.165 27.065 88.375 28.155 ;
        RECT 88.545 28.155 89.065 28.695 ;
        RECT 89.235 28.325 89.755 28.865 ;
        RECT 88.545 27.065 89.755 28.155 ;
        RECT 12.100 26.895 89.840 27.065 ;
        RECT 12.185 25.805 13.395 26.895 ;
        RECT 13.565 26.460 18.910 26.895 ;
        RECT 19.085 26.460 24.430 26.895 ;
        RECT 12.185 25.095 12.705 25.635 ;
        RECT 12.875 25.265 13.395 25.805 ;
        RECT 12.185 24.345 13.395 25.095 ;
        RECT 15.150 24.890 15.490 25.720 ;
        RECT 16.970 25.210 17.320 26.460 ;
        RECT 20.670 24.890 21.010 25.720 ;
        RECT 22.490 25.210 22.840 26.460 ;
        RECT 25.065 25.730 25.355 26.895 ;
        RECT 25.525 26.460 30.870 26.895 ;
        RECT 31.045 26.460 36.390 26.895 ;
        RECT 36.565 26.460 41.910 26.895 ;
        RECT 42.085 26.460 47.430 26.895 ;
        RECT 13.565 24.345 18.910 24.890 ;
        RECT 19.085 24.345 24.430 24.890 ;
        RECT 25.065 24.345 25.355 25.070 ;
        RECT 27.110 24.890 27.450 25.720 ;
        RECT 28.930 25.210 29.280 26.460 ;
        RECT 32.630 24.890 32.970 25.720 ;
        RECT 34.450 25.210 34.800 26.460 ;
        RECT 38.150 24.890 38.490 25.720 ;
        RECT 39.970 25.210 40.320 26.460 ;
        RECT 43.670 24.890 44.010 25.720 ;
        RECT 45.490 25.210 45.840 26.460 ;
        RECT 47.605 25.805 49.275 26.895 ;
        RECT 47.605 25.115 48.355 25.635 ;
        RECT 48.525 25.285 49.275 25.805 ;
        RECT 49.445 25.820 49.715 26.725 ;
        RECT 49.885 26.135 50.215 26.895 ;
        RECT 50.395 25.965 50.565 26.725 ;
        RECT 25.525 24.345 30.870 24.890 ;
        RECT 31.045 24.345 36.390 24.890 ;
        RECT 36.565 24.345 41.910 24.890 ;
        RECT 42.085 24.345 47.430 24.890 ;
        RECT 47.605 24.345 49.275 25.115 ;
        RECT 49.445 25.020 49.615 25.820 ;
        RECT 49.900 25.795 50.565 25.965 ;
        RECT 49.900 25.650 50.070 25.795 ;
        RECT 50.825 25.730 51.115 26.895 ;
        RECT 52.320 26.265 52.605 26.725 ;
        RECT 52.775 26.435 53.045 26.895 ;
        RECT 52.320 26.045 53.275 26.265 ;
        RECT 49.785 25.320 50.070 25.650 ;
        RECT 49.900 25.065 50.070 25.320 ;
        RECT 50.305 25.245 50.635 25.615 ;
        RECT 52.205 25.315 52.895 25.875 ;
        RECT 53.065 25.145 53.275 26.045 ;
        RECT 49.445 24.515 49.705 25.020 ;
        RECT 49.900 24.895 50.565 25.065 ;
        RECT 49.885 24.345 50.215 24.725 ;
        RECT 50.395 24.515 50.565 24.895 ;
        RECT 50.825 24.345 51.115 25.070 ;
        RECT 52.320 24.975 53.275 25.145 ;
        RECT 53.445 25.875 53.845 26.725 ;
        RECT 54.035 26.265 54.315 26.725 ;
        RECT 54.835 26.435 55.160 26.895 ;
        RECT 54.035 26.045 55.160 26.265 ;
        RECT 53.445 25.315 54.540 25.875 ;
        RECT 54.710 25.585 55.160 26.045 ;
        RECT 55.330 25.755 55.715 26.725 ;
        RECT 55.975 26.225 56.145 26.725 ;
        RECT 56.315 26.395 56.645 26.895 ;
        RECT 55.975 26.055 56.640 26.225 ;
        RECT 52.320 24.515 52.605 24.975 ;
        RECT 52.775 24.345 53.045 24.805 ;
        RECT 53.445 24.515 53.845 25.315 ;
        RECT 54.710 25.255 55.265 25.585 ;
        RECT 54.710 25.145 55.160 25.255 ;
        RECT 54.035 24.975 55.160 25.145 ;
        RECT 55.435 25.085 55.715 25.755 ;
        RECT 55.890 25.235 56.240 25.885 ;
        RECT 54.035 24.515 54.315 24.975 ;
        RECT 54.835 24.345 55.160 24.805 ;
        RECT 55.330 24.515 55.715 25.085 ;
        RECT 56.410 25.065 56.640 26.055 ;
        RECT 55.975 24.895 56.640 25.065 ;
        RECT 55.975 24.605 56.145 24.895 ;
        RECT 56.315 24.345 56.645 24.725 ;
        RECT 56.815 24.605 57.000 26.725 ;
        RECT 57.240 26.435 57.505 26.895 ;
        RECT 57.675 26.300 57.925 26.725 ;
        RECT 58.135 26.450 59.240 26.620 ;
        RECT 57.620 26.170 57.925 26.300 ;
        RECT 57.170 24.975 57.450 25.925 ;
        RECT 57.620 25.065 57.790 26.170 ;
        RECT 57.960 25.385 58.200 25.980 ;
        RECT 58.370 25.915 58.900 26.280 ;
        RECT 58.370 25.215 58.540 25.915 ;
        RECT 59.070 25.835 59.240 26.450 ;
        RECT 59.410 26.095 59.580 26.895 ;
        RECT 59.750 26.395 60.000 26.725 ;
        RECT 60.225 26.425 61.110 26.595 ;
        RECT 59.070 25.745 59.580 25.835 ;
        RECT 57.620 24.935 57.845 25.065 ;
        RECT 58.015 24.995 58.540 25.215 ;
        RECT 58.710 25.575 59.580 25.745 ;
        RECT 57.255 24.345 57.505 24.805 ;
        RECT 57.675 24.795 57.845 24.935 ;
        RECT 58.710 24.795 58.880 25.575 ;
        RECT 59.410 25.505 59.580 25.575 ;
        RECT 59.090 25.325 59.290 25.355 ;
        RECT 59.750 25.325 59.920 26.395 ;
        RECT 60.090 25.505 60.280 26.225 ;
        RECT 59.090 25.025 59.920 25.325 ;
        RECT 60.450 25.295 60.770 26.255 ;
        RECT 57.675 24.625 58.010 24.795 ;
        RECT 58.205 24.625 58.880 24.795 ;
        RECT 59.200 24.345 59.570 24.845 ;
        RECT 59.750 24.795 59.920 25.025 ;
        RECT 60.305 24.965 60.770 25.295 ;
        RECT 60.940 25.585 61.110 26.425 ;
        RECT 61.290 26.395 61.605 26.895 ;
        RECT 61.835 26.165 62.175 26.725 ;
        RECT 61.280 25.790 62.175 26.165 ;
        RECT 62.345 25.885 62.515 26.895 ;
        RECT 61.985 25.585 62.175 25.790 ;
        RECT 62.685 25.835 63.015 26.680 ;
        RECT 63.245 26.340 63.850 26.895 ;
        RECT 64.025 26.385 64.505 26.725 ;
        RECT 64.675 26.350 64.930 26.895 ;
        RECT 63.245 26.240 63.860 26.340 ;
        RECT 63.675 26.215 63.860 26.240 ;
        RECT 62.685 25.755 63.075 25.835 ;
        RECT 62.860 25.705 63.075 25.755 ;
        RECT 60.940 25.255 61.815 25.585 ;
        RECT 61.985 25.255 62.735 25.585 ;
        RECT 60.940 24.795 61.110 25.255 ;
        RECT 61.985 25.085 62.185 25.255 ;
        RECT 62.905 25.125 63.075 25.705 ;
        RECT 63.245 25.620 63.505 26.070 ;
        RECT 63.675 25.970 64.005 26.215 ;
        RECT 64.175 25.895 64.930 26.145 ;
        RECT 65.100 26.025 65.375 26.725 ;
        RECT 66.555 26.225 66.725 26.725 ;
        RECT 66.895 26.395 67.225 26.895 ;
        RECT 66.555 26.055 67.220 26.225 ;
        RECT 64.160 25.860 64.930 25.895 ;
        RECT 64.145 25.850 64.930 25.860 ;
        RECT 64.140 25.835 65.035 25.850 ;
        RECT 64.120 25.820 65.035 25.835 ;
        RECT 64.100 25.810 65.035 25.820 ;
        RECT 64.075 25.800 65.035 25.810 ;
        RECT 64.005 25.770 65.035 25.800 ;
        RECT 63.985 25.740 65.035 25.770 ;
        RECT 63.965 25.710 65.035 25.740 ;
        RECT 63.935 25.685 65.035 25.710 ;
        RECT 63.900 25.650 65.035 25.685 ;
        RECT 63.870 25.645 65.035 25.650 ;
        RECT 63.870 25.640 64.260 25.645 ;
        RECT 63.870 25.630 64.235 25.640 ;
        RECT 63.870 25.625 64.220 25.630 ;
        RECT 63.870 25.620 64.205 25.625 ;
        RECT 63.245 25.615 64.205 25.620 ;
        RECT 63.245 25.605 64.195 25.615 ;
        RECT 63.245 25.600 64.185 25.605 ;
        RECT 63.245 25.590 64.175 25.600 ;
        RECT 63.245 25.580 64.170 25.590 ;
        RECT 63.245 25.575 64.165 25.580 ;
        RECT 63.245 25.560 64.155 25.575 ;
        RECT 63.245 25.545 64.150 25.560 ;
        RECT 63.245 25.520 64.140 25.545 ;
        RECT 63.245 25.450 64.135 25.520 ;
        RECT 62.850 25.085 63.075 25.125 ;
        RECT 59.750 24.625 60.155 24.795 ;
        RECT 60.325 24.625 61.110 24.795 ;
        RECT 61.385 24.345 61.595 24.875 ;
        RECT 61.855 24.560 62.185 25.085 ;
        RECT 62.695 25.000 63.075 25.085 ;
        RECT 62.355 24.345 62.525 24.955 ;
        RECT 62.695 24.565 63.025 25.000 ;
        RECT 63.245 24.895 63.795 25.280 ;
        RECT 63.965 24.725 64.135 25.450 ;
        RECT 63.245 24.555 64.135 24.725 ;
        RECT 64.305 25.050 64.635 25.475 ;
        RECT 64.805 25.250 65.035 25.645 ;
        RECT 64.305 24.565 64.525 25.050 ;
        RECT 65.205 24.995 65.375 26.025 ;
        RECT 66.470 25.235 66.820 25.885 ;
        RECT 66.990 25.065 67.220 26.055 ;
        RECT 64.695 24.345 64.945 24.885 ;
        RECT 65.115 24.515 65.375 24.995 ;
        RECT 66.555 24.895 67.220 25.065 ;
        RECT 66.555 24.605 66.725 24.895 ;
        RECT 66.895 24.345 67.225 24.725 ;
        RECT 67.395 24.605 67.580 26.725 ;
        RECT 67.820 26.435 68.085 26.895 ;
        RECT 68.255 26.300 68.505 26.725 ;
        RECT 68.715 26.450 69.820 26.620 ;
        RECT 68.200 26.170 68.505 26.300 ;
        RECT 67.750 24.975 68.030 25.925 ;
        RECT 68.200 25.065 68.370 26.170 ;
        RECT 68.540 25.385 68.780 25.980 ;
        RECT 68.950 25.915 69.480 26.280 ;
        RECT 68.950 25.215 69.120 25.915 ;
        RECT 69.650 25.835 69.820 26.450 ;
        RECT 69.990 26.095 70.160 26.895 ;
        RECT 70.330 26.395 70.580 26.725 ;
        RECT 70.805 26.425 71.690 26.595 ;
        RECT 69.650 25.745 70.160 25.835 ;
        RECT 68.200 24.935 68.425 25.065 ;
        RECT 68.595 24.995 69.120 25.215 ;
        RECT 69.290 25.575 70.160 25.745 ;
        RECT 67.835 24.345 68.085 24.805 ;
        RECT 68.255 24.795 68.425 24.935 ;
        RECT 69.290 24.795 69.460 25.575 ;
        RECT 69.990 25.505 70.160 25.575 ;
        RECT 69.670 25.325 69.870 25.355 ;
        RECT 70.330 25.325 70.500 26.395 ;
        RECT 70.670 25.505 70.860 26.225 ;
        RECT 69.670 25.025 70.500 25.325 ;
        RECT 71.030 25.295 71.350 26.255 ;
        RECT 68.255 24.625 68.590 24.795 ;
        RECT 68.785 24.625 69.460 24.795 ;
        RECT 69.780 24.345 70.150 24.845 ;
        RECT 70.330 24.795 70.500 25.025 ;
        RECT 70.885 24.965 71.350 25.295 ;
        RECT 71.520 25.585 71.690 26.425 ;
        RECT 71.870 26.395 72.185 26.895 ;
        RECT 72.415 26.165 72.755 26.725 ;
        RECT 71.860 25.790 72.755 26.165 ;
        RECT 72.925 25.885 73.095 26.895 ;
        RECT 72.565 25.585 72.755 25.790 ;
        RECT 73.265 25.835 73.595 26.680 ;
        RECT 74.010 25.925 74.400 26.100 ;
        RECT 74.885 26.095 75.215 26.895 ;
        RECT 75.385 26.105 75.920 26.725 ;
        RECT 73.265 25.755 73.655 25.835 ;
        RECT 74.010 25.755 75.435 25.925 ;
        RECT 73.440 25.705 73.655 25.755 ;
        RECT 71.520 25.255 72.395 25.585 ;
        RECT 72.565 25.255 73.315 25.585 ;
        RECT 71.520 24.795 71.690 25.255 ;
        RECT 72.565 25.085 72.765 25.255 ;
        RECT 73.485 25.125 73.655 25.705 ;
        RECT 73.430 25.085 73.655 25.125 ;
        RECT 70.330 24.625 70.735 24.795 ;
        RECT 70.905 24.625 71.690 24.795 ;
        RECT 71.965 24.345 72.175 24.875 ;
        RECT 72.435 24.560 72.765 25.085 ;
        RECT 73.275 25.000 73.655 25.085 ;
        RECT 73.885 25.025 74.240 25.585 ;
        RECT 72.935 24.345 73.105 24.955 ;
        RECT 73.275 24.565 73.605 25.000 ;
        RECT 74.410 24.855 74.580 25.755 ;
        RECT 74.750 25.025 75.015 25.585 ;
        RECT 75.265 25.255 75.435 25.755 ;
        RECT 75.605 25.085 75.920 26.105 ;
        RECT 76.585 25.730 76.875 26.895 ;
        RECT 77.045 25.755 77.385 26.725 ;
        RECT 77.555 25.755 77.725 26.895 ;
        RECT 77.995 26.095 78.245 26.895 ;
        RECT 78.890 25.925 79.220 26.725 ;
        RECT 79.520 26.095 79.850 26.895 ;
        RECT 80.020 25.925 80.350 26.725 ;
        RECT 81.275 26.225 81.445 26.725 ;
        RECT 81.615 26.395 81.945 26.895 ;
        RECT 81.275 26.055 81.940 26.225 ;
        RECT 77.915 25.755 80.350 25.925 ;
        RECT 73.990 24.345 74.230 24.855 ;
        RECT 74.410 24.525 74.690 24.855 ;
        RECT 74.920 24.345 75.135 24.855 ;
        RECT 75.305 24.515 75.920 25.085 ;
        RECT 77.045 25.145 77.220 25.755 ;
        RECT 77.915 25.505 78.085 25.755 ;
        RECT 77.390 25.335 78.085 25.505 ;
        RECT 78.260 25.335 78.680 25.535 ;
        RECT 78.850 25.335 79.180 25.535 ;
        RECT 79.350 25.335 79.680 25.535 ;
        RECT 76.585 24.345 76.875 25.070 ;
        RECT 77.045 24.515 77.385 25.145 ;
        RECT 77.555 24.345 77.805 25.145 ;
        RECT 77.995 24.995 79.220 25.165 ;
        RECT 77.995 24.515 78.325 24.995 ;
        RECT 78.495 24.345 78.720 24.805 ;
        RECT 78.890 24.515 79.220 24.995 ;
        RECT 79.850 25.125 80.020 25.755 ;
        RECT 80.205 25.335 80.555 25.585 ;
        RECT 81.190 25.235 81.540 25.885 ;
        RECT 79.850 24.515 80.350 25.125 ;
        RECT 81.710 25.065 81.940 26.055 ;
        RECT 81.275 24.895 81.940 25.065 ;
        RECT 81.275 24.605 81.445 24.895 ;
        RECT 81.615 24.345 81.945 24.725 ;
        RECT 82.115 24.605 82.300 26.725 ;
        RECT 82.540 26.435 82.805 26.895 ;
        RECT 82.975 26.300 83.225 26.725 ;
        RECT 83.435 26.450 84.540 26.620 ;
        RECT 82.920 26.170 83.225 26.300 ;
        RECT 82.470 24.975 82.750 25.925 ;
        RECT 82.920 25.065 83.090 26.170 ;
        RECT 83.260 25.385 83.500 25.980 ;
        RECT 83.670 25.915 84.200 26.280 ;
        RECT 83.670 25.215 83.840 25.915 ;
        RECT 84.370 25.835 84.540 26.450 ;
        RECT 84.710 26.095 84.880 26.895 ;
        RECT 85.050 26.395 85.300 26.725 ;
        RECT 85.525 26.425 86.410 26.595 ;
        RECT 84.370 25.745 84.880 25.835 ;
        RECT 82.920 24.935 83.145 25.065 ;
        RECT 83.315 24.995 83.840 25.215 ;
        RECT 84.010 25.575 84.880 25.745 ;
        RECT 82.555 24.345 82.805 24.805 ;
        RECT 82.975 24.795 83.145 24.935 ;
        RECT 84.010 24.795 84.180 25.575 ;
        RECT 84.710 25.505 84.880 25.575 ;
        RECT 84.390 25.325 84.590 25.355 ;
        RECT 85.050 25.325 85.220 26.395 ;
        RECT 85.390 25.505 85.580 26.225 ;
        RECT 84.390 25.025 85.220 25.325 ;
        RECT 85.750 25.295 86.070 26.255 ;
        RECT 82.975 24.625 83.310 24.795 ;
        RECT 83.505 24.625 84.180 24.795 ;
        RECT 84.500 24.345 84.870 24.845 ;
        RECT 85.050 24.795 85.220 25.025 ;
        RECT 85.605 24.965 86.070 25.295 ;
        RECT 86.240 25.585 86.410 26.425 ;
        RECT 86.590 26.395 86.905 26.895 ;
        RECT 87.135 26.165 87.475 26.725 ;
        RECT 86.580 25.790 87.475 26.165 ;
        RECT 87.645 25.885 87.815 26.895 ;
        RECT 87.285 25.585 87.475 25.790 ;
        RECT 87.985 25.835 88.315 26.680 ;
        RECT 87.985 25.755 88.375 25.835 ;
        RECT 88.160 25.705 88.375 25.755 ;
        RECT 86.240 25.255 87.115 25.585 ;
        RECT 87.285 25.255 88.035 25.585 ;
        RECT 86.240 24.795 86.410 25.255 ;
        RECT 87.285 25.085 87.485 25.255 ;
        RECT 88.205 25.125 88.375 25.705 ;
        RECT 88.545 25.805 89.755 26.895 ;
        RECT 88.545 25.265 89.065 25.805 ;
        RECT 88.150 25.085 88.375 25.125 ;
        RECT 89.235 25.095 89.755 25.635 ;
        RECT 85.050 24.625 85.455 24.795 ;
        RECT 85.625 24.625 86.410 24.795 ;
        RECT 86.685 24.345 86.895 24.875 ;
        RECT 87.155 24.560 87.485 25.085 ;
        RECT 87.995 25.000 88.375 25.085 ;
        RECT 87.655 24.345 87.825 24.955 ;
        RECT 87.995 24.565 88.325 25.000 ;
        RECT 88.545 24.345 89.755 25.095 ;
        RECT 12.100 24.175 89.840 24.345 ;
        RECT 12.185 23.425 13.395 24.175 ;
        RECT 13.565 23.630 18.910 24.175 ;
        RECT 19.085 23.630 24.430 24.175 ;
        RECT 24.605 23.630 29.950 24.175 ;
        RECT 30.125 23.630 35.470 24.175 ;
        RECT 12.185 22.885 12.705 23.425 ;
        RECT 12.875 22.715 13.395 23.255 ;
        RECT 15.150 22.800 15.490 23.630 ;
        RECT 12.185 21.625 13.395 22.715 ;
        RECT 16.970 22.060 17.320 23.310 ;
        RECT 20.670 22.800 21.010 23.630 ;
        RECT 22.490 22.060 22.840 23.310 ;
        RECT 26.190 22.800 26.530 23.630 ;
        RECT 28.010 22.060 28.360 23.310 ;
        RECT 31.710 22.800 32.050 23.630 ;
        RECT 35.645 23.405 37.315 24.175 ;
        RECT 37.945 23.450 38.235 24.175 ;
        RECT 38.405 23.630 43.750 24.175 ;
        RECT 33.530 22.060 33.880 23.310 ;
        RECT 35.645 22.885 36.395 23.405 ;
        RECT 36.565 22.715 37.315 23.235 ;
        RECT 39.990 22.800 40.330 23.630 ;
        RECT 43.925 23.405 46.515 24.175 ;
        RECT 46.775 23.625 46.945 23.915 ;
        RECT 47.115 23.795 47.445 24.175 ;
        RECT 46.775 23.455 47.440 23.625 ;
        RECT 13.565 21.625 18.910 22.060 ;
        RECT 19.085 21.625 24.430 22.060 ;
        RECT 24.605 21.625 29.950 22.060 ;
        RECT 30.125 21.625 35.470 22.060 ;
        RECT 35.645 21.625 37.315 22.715 ;
        RECT 37.945 21.625 38.235 22.790 ;
        RECT 41.810 22.060 42.160 23.310 ;
        RECT 43.925 22.885 45.135 23.405 ;
        RECT 45.305 22.715 46.515 23.235 ;
        RECT 38.405 21.625 43.750 22.060 ;
        RECT 43.925 21.625 46.515 22.715 ;
        RECT 46.690 22.635 47.040 23.285 ;
        RECT 47.210 22.465 47.440 23.455 ;
        RECT 46.775 22.295 47.440 22.465 ;
        RECT 46.775 21.795 46.945 22.295 ;
        RECT 47.115 21.625 47.445 22.125 ;
        RECT 47.615 21.795 47.800 23.915 ;
        RECT 48.055 23.715 48.305 24.175 ;
        RECT 48.475 23.725 48.810 23.895 ;
        RECT 49.005 23.725 49.680 23.895 ;
        RECT 48.475 23.585 48.645 23.725 ;
        RECT 47.970 22.595 48.250 23.545 ;
        RECT 48.420 23.455 48.645 23.585 ;
        RECT 48.420 22.350 48.590 23.455 ;
        RECT 48.815 23.305 49.340 23.525 ;
        RECT 48.760 22.540 49.000 23.135 ;
        RECT 49.170 22.605 49.340 23.305 ;
        RECT 49.510 22.945 49.680 23.725 ;
        RECT 50.000 23.675 50.370 24.175 ;
        RECT 50.550 23.725 50.955 23.895 ;
        RECT 51.125 23.725 51.910 23.895 ;
        RECT 50.550 23.495 50.720 23.725 ;
        RECT 49.890 23.195 50.720 23.495 ;
        RECT 51.105 23.225 51.570 23.555 ;
        RECT 49.890 23.165 50.090 23.195 ;
        RECT 50.210 22.945 50.380 23.015 ;
        RECT 49.510 22.775 50.380 22.945 ;
        RECT 49.870 22.685 50.380 22.775 ;
        RECT 48.420 22.220 48.725 22.350 ;
        RECT 49.170 22.240 49.700 22.605 ;
        RECT 48.040 21.625 48.305 22.085 ;
        RECT 48.475 21.795 48.725 22.220 ;
        RECT 49.870 22.070 50.040 22.685 ;
        RECT 48.935 21.900 50.040 22.070 ;
        RECT 50.210 21.625 50.380 22.425 ;
        RECT 50.550 22.125 50.720 23.195 ;
        RECT 50.890 22.295 51.080 23.015 ;
        RECT 51.250 22.265 51.570 23.225 ;
        RECT 51.740 23.265 51.910 23.725 ;
        RECT 52.185 23.645 52.395 24.175 ;
        RECT 52.655 23.435 52.985 23.960 ;
        RECT 53.155 23.565 53.325 24.175 ;
        RECT 53.495 23.520 53.825 23.955 ;
        RECT 53.495 23.435 53.875 23.520 ;
        RECT 52.785 23.265 52.985 23.435 ;
        RECT 53.650 23.395 53.875 23.435 ;
        RECT 51.740 22.935 52.615 23.265 ;
        RECT 52.785 22.935 53.535 23.265 ;
        RECT 50.550 21.795 50.800 22.125 ;
        RECT 51.740 22.095 51.910 22.935 ;
        RECT 52.785 22.730 52.975 22.935 ;
        RECT 53.705 22.815 53.875 23.395 ;
        RECT 54.045 23.405 57.555 24.175 ;
        RECT 58.650 23.435 58.905 24.005 ;
        RECT 59.075 23.775 59.405 24.175 ;
        RECT 59.830 23.640 60.360 24.005 ;
        RECT 60.550 23.835 60.825 24.005 ;
        RECT 60.545 23.665 60.825 23.835 ;
        RECT 59.830 23.605 60.005 23.640 ;
        RECT 59.075 23.435 60.005 23.605 ;
        RECT 54.045 22.885 55.695 23.405 ;
        RECT 53.660 22.765 53.875 22.815 ;
        RECT 52.080 22.355 52.975 22.730 ;
        RECT 53.485 22.685 53.875 22.765 ;
        RECT 55.865 22.715 57.555 23.235 ;
        RECT 51.025 21.925 51.910 22.095 ;
        RECT 52.090 21.625 52.405 22.125 ;
        RECT 52.635 21.795 52.975 22.355 ;
        RECT 53.145 21.625 53.315 22.635 ;
        RECT 53.485 21.840 53.815 22.685 ;
        RECT 54.045 21.625 57.555 22.715 ;
        RECT 58.650 22.765 58.820 23.435 ;
        RECT 59.075 23.265 59.245 23.435 ;
        RECT 58.990 22.935 59.245 23.265 ;
        RECT 59.470 22.935 59.665 23.265 ;
        RECT 58.650 21.795 58.985 22.765 ;
        RECT 59.155 21.625 59.325 22.765 ;
        RECT 59.495 21.965 59.665 22.935 ;
        RECT 59.835 22.305 60.005 23.435 ;
        RECT 60.175 22.645 60.345 23.445 ;
        RECT 60.550 22.845 60.825 23.665 ;
        RECT 60.995 22.645 61.185 24.005 ;
        RECT 61.365 23.640 61.875 24.175 ;
        RECT 62.095 23.365 62.340 23.970 ;
        RECT 63.705 23.450 63.995 24.175 ;
        RECT 64.165 23.630 69.510 24.175 ;
        RECT 61.385 23.195 62.615 23.365 ;
        RECT 60.175 22.475 61.185 22.645 ;
        RECT 61.355 22.630 62.105 22.820 ;
        RECT 59.835 22.135 60.960 22.305 ;
        RECT 61.355 21.965 61.525 22.630 ;
        RECT 62.275 22.385 62.615 23.195 ;
        RECT 65.750 22.800 66.090 23.630 ;
        RECT 70.235 23.625 70.405 23.915 ;
        RECT 70.575 23.795 70.905 24.175 ;
        RECT 70.235 23.455 70.900 23.625 ;
        RECT 59.495 21.795 61.525 21.965 ;
        RECT 61.695 21.625 61.865 22.385 ;
        RECT 62.100 21.975 62.615 22.385 ;
        RECT 63.705 21.625 63.995 22.790 ;
        RECT 67.570 22.060 67.920 23.310 ;
        RECT 70.150 22.635 70.500 23.285 ;
        RECT 70.670 22.465 70.900 23.455 ;
        RECT 70.235 22.295 70.900 22.465 ;
        RECT 64.165 21.625 69.510 22.060 ;
        RECT 70.235 21.795 70.405 22.295 ;
        RECT 70.575 21.625 70.905 22.125 ;
        RECT 71.075 21.795 71.260 23.915 ;
        RECT 71.515 23.715 71.765 24.175 ;
        RECT 71.935 23.725 72.270 23.895 ;
        RECT 72.465 23.725 73.140 23.895 ;
        RECT 71.935 23.585 72.105 23.725 ;
        RECT 71.430 22.595 71.710 23.545 ;
        RECT 71.880 23.455 72.105 23.585 ;
        RECT 71.880 22.350 72.050 23.455 ;
        RECT 72.275 23.305 72.800 23.525 ;
        RECT 72.220 22.540 72.460 23.135 ;
        RECT 72.630 22.605 72.800 23.305 ;
        RECT 72.970 22.945 73.140 23.725 ;
        RECT 73.460 23.675 73.830 24.175 ;
        RECT 74.010 23.725 74.415 23.895 ;
        RECT 74.585 23.725 75.370 23.895 ;
        RECT 74.010 23.495 74.180 23.725 ;
        RECT 73.350 23.195 74.180 23.495 ;
        RECT 74.565 23.225 75.030 23.555 ;
        RECT 73.350 23.165 73.550 23.195 ;
        RECT 73.670 22.945 73.840 23.015 ;
        RECT 72.970 22.775 73.840 22.945 ;
        RECT 73.330 22.685 73.840 22.775 ;
        RECT 71.880 22.220 72.185 22.350 ;
        RECT 72.630 22.240 73.160 22.605 ;
        RECT 71.500 21.625 71.765 22.085 ;
        RECT 71.935 21.795 72.185 22.220 ;
        RECT 73.330 22.070 73.500 22.685 ;
        RECT 72.395 21.900 73.500 22.070 ;
        RECT 73.670 21.625 73.840 22.425 ;
        RECT 74.010 22.125 74.180 23.195 ;
        RECT 74.350 22.295 74.540 23.015 ;
        RECT 74.710 22.265 75.030 23.225 ;
        RECT 75.200 23.265 75.370 23.725 ;
        RECT 75.645 23.645 75.855 24.175 ;
        RECT 76.115 23.435 76.445 23.960 ;
        RECT 76.615 23.565 76.785 24.175 ;
        RECT 76.955 23.520 77.285 23.955 ;
        RECT 77.595 23.625 77.765 24.005 ;
        RECT 77.945 23.795 78.275 24.175 ;
        RECT 76.955 23.435 77.335 23.520 ;
        RECT 77.595 23.455 78.260 23.625 ;
        RECT 78.455 23.500 78.715 24.005 ;
        RECT 79.050 23.665 79.290 24.175 ;
        RECT 79.470 23.665 79.750 23.995 ;
        RECT 79.980 23.665 80.195 24.175 ;
        RECT 76.245 23.265 76.445 23.435 ;
        RECT 77.110 23.395 77.335 23.435 ;
        RECT 75.200 22.935 76.075 23.265 ;
        RECT 76.245 22.935 76.995 23.265 ;
        RECT 74.010 21.795 74.260 22.125 ;
        RECT 75.200 22.095 75.370 22.935 ;
        RECT 76.245 22.730 76.435 22.935 ;
        RECT 77.165 22.815 77.335 23.395 ;
        RECT 77.525 22.905 77.855 23.275 ;
        RECT 78.090 23.200 78.260 23.455 ;
        RECT 77.120 22.765 77.335 22.815 ;
        RECT 75.540 22.355 76.435 22.730 ;
        RECT 76.945 22.685 77.335 22.765 ;
        RECT 78.090 22.870 78.375 23.200 ;
        RECT 78.090 22.725 78.260 22.870 ;
        RECT 74.485 21.925 75.370 22.095 ;
        RECT 75.550 21.625 75.865 22.125 ;
        RECT 76.095 21.795 76.435 22.355 ;
        RECT 76.605 21.625 76.775 22.635 ;
        RECT 76.945 21.840 77.275 22.685 ;
        RECT 77.595 22.555 78.260 22.725 ;
        RECT 78.545 22.700 78.715 23.500 ;
        RECT 78.945 22.935 79.300 23.495 ;
        RECT 79.470 22.765 79.640 23.665 ;
        RECT 79.810 22.935 80.075 23.495 ;
        RECT 80.365 23.435 80.980 24.005 ;
        RECT 81.275 23.625 81.445 23.915 ;
        RECT 81.615 23.795 81.945 24.175 ;
        RECT 81.275 23.455 81.940 23.625 ;
        RECT 80.325 22.765 80.495 23.265 ;
        RECT 77.595 21.795 77.765 22.555 ;
        RECT 77.945 21.625 78.275 22.385 ;
        RECT 78.445 21.795 78.715 22.700 ;
        RECT 79.070 22.595 80.495 22.765 ;
        RECT 79.070 22.420 79.460 22.595 ;
        RECT 79.945 21.625 80.275 22.425 ;
        RECT 80.665 22.415 80.980 23.435 ;
        RECT 81.190 22.635 81.540 23.285 ;
        RECT 81.710 22.465 81.940 23.455 ;
        RECT 80.445 21.795 80.980 22.415 ;
        RECT 81.275 22.295 81.940 22.465 ;
        RECT 81.275 21.795 81.445 22.295 ;
        RECT 81.615 21.625 81.945 22.125 ;
        RECT 82.115 21.795 82.300 23.915 ;
        RECT 82.555 23.715 82.805 24.175 ;
        RECT 82.975 23.725 83.310 23.895 ;
        RECT 83.505 23.725 84.180 23.895 ;
        RECT 82.975 23.585 83.145 23.725 ;
        RECT 82.470 22.595 82.750 23.545 ;
        RECT 82.920 23.455 83.145 23.585 ;
        RECT 82.920 22.350 83.090 23.455 ;
        RECT 83.315 23.305 83.840 23.525 ;
        RECT 83.260 22.540 83.500 23.135 ;
        RECT 83.670 22.605 83.840 23.305 ;
        RECT 84.010 22.945 84.180 23.725 ;
        RECT 84.500 23.675 84.870 24.175 ;
        RECT 85.050 23.725 85.455 23.895 ;
        RECT 85.625 23.725 86.410 23.895 ;
        RECT 85.050 23.495 85.220 23.725 ;
        RECT 84.390 23.195 85.220 23.495 ;
        RECT 85.605 23.225 86.070 23.555 ;
        RECT 84.390 23.165 84.590 23.195 ;
        RECT 84.710 22.945 84.880 23.015 ;
        RECT 84.010 22.775 84.880 22.945 ;
        RECT 84.370 22.685 84.880 22.775 ;
        RECT 82.920 22.220 83.225 22.350 ;
        RECT 83.670 22.240 84.200 22.605 ;
        RECT 82.540 21.625 82.805 22.085 ;
        RECT 82.975 21.795 83.225 22.220 ;
        RECT 84.370 22.070 84.540 22.685 ;
        RECT 83.435 21.900 84.540 22.070 ;
        RECT 84.710 21.625 84.880 22.425 ;
        RECT 85.050 22.125 85.220 23.195 ;
        RECT 85.390 22.295 85.580 23.015 ;
        RECT 85.750 22.265 86.070 23.225 ;
        RECT 86.240 23.265 86.410 23.725 ;
        RECT 86.685 23.645 86.895 24.175 ;
        RECT 87.155 23.435 87.485 23.960 ;
        RECT 87.655 23.565 87.825 24.175 ;
        RECT 87.995 23.520 88.325 23.955 ;
        RECT 87.995 23.435 88.375 23.520 ;
        RECT 87.285 23.265 87.485 23.435 ;
        RECT 88.150 23.395 88.375 23.435 ;
        RECT 88.545 23.425 89.755 24.175 ;
        RECT 86.240 22.935 87.115 23.265 ;
        RECT 87.285 22.935 88.035 23.265 ;
        RECT 85.050 21.795 85.300 22.125 ;
        RECT 86.240 22.095 86.410 22.935 ;
        RECT 87.285 22.730 87.475 22.935 ;
        RECT 88.205 22.815 88.375 23.395 ;
        RECT 88.160 22.765 88.375 22.815 ;
        RECT 86.580 22.355 87.475 22.730 ;
        RECT 87.985 22.685 88.375 22.765 ;
        RECT 88.545 22.715 89.065 23.255 ;
        RECT 89.235 22.885 89.755 23.425 ;
        RECT 85.525 21.925 86.410 22.095 ;
        RECT 86.590 21.625 86.905 22.125 ;
        RECT 87.135 21.795 87.475 22.355 ;
        RECT 87.645 21.625 87.815 22.635 ;
        RECT 87.985 21.840 88.315 22.685 ;
        RECT 88.545 21.625 89.755 22.715 ;
        RECT 12.100 21.455 89.840 21.625 ;
        RECT 12.185 20.365 13.395 21.455 ;
        RECT 13.565 21.020 18.910 21.455 ;
        RECT 19.085 21.020 24.430 21.455 ;
        RECT 12.185 19.655 12.705 20.195 ;
        RECT 12.875 19.825 13.395 20.365 ;
        RECT 12.185 18.905 13.395 19.655 ;
        RECT 15.150 19.450 15.490 20.280 ;
        RECT 16.970 19.770 17.320 21.020 ;
        RECT 20.670 19.450 21.010 20.280 ;
        RECT 22.490 19.770 22.840 21.020 ;
        RECT 25.065 20.290 25.355 21.455 ;
        RECT 25.525 21.020 30.870 21.455 ;
        RECT 31.045 21.020 36.390 21.455 ;
        RECT 13.565 18.905 18.910 19.450 ;
        RECT 19.085 18.905 24.430 19.450 ;
        RECT 25.065 18.905 25.355 19.630 ;
        RECT 27.110 19.450 27.450 20.280 ;
        RECT 28.930 19.770 29.280 21.020 ;
        RECT 32.630 19.450 32.970 20.280 ;
        RECT 34.450 19.770 34.800 21.020 ;
        RECT 36.565 20.365 37.775 21.455 ;
        RECT 36.565 19.655 37.085 20.195 ;
        RECT 37.255 19.825 37.775 20.365 ;
        RECT 37.945 20.290 38.235 21.455 ;
        RECT 38.405 20.365 41.915 21.455 ;
        RECT 42.545 20.860 42.980 21.285 ;
        RECT 43.150 21.030 43.535 21.455 ;
        RECT 42.545 20.690 43.535 20.860 ;
        RECT 38.405 19.675 40.055 20.195 ;
        RECT 40.225 19.845 41.915 20.365 ;
        RECT 42.545 19.815 43.030 20.520 ;
        RECT 43.200 20.145 43.535 20.690 ;
        RECT 43.705 20.495 44.130 21.285 ;
        RECT 44.300 20.860 44.575 21.285 ;
        RECT 44.745 21.030 45.130 21.455 ;
        RECT 44.300 20.665 45.130 20.860 ;
        RECT 43.705 20.315 44.610 20.495 ;
        RECT 43.200 19.815 43.610 20.145 ;
        RECT 43.780 19.815 44.610 20.315 ;
        RECT 44.780 20.145 45.130 20.665 ;
        RECT 45.300 20.495 45.545 21.285 ;
        RECT 45.735 20.860 45.990 21.285 ;
        RECT 46.160 21.030 46.545 21.455 ;
        RECT 45.735 20.665 46.545 20.860 ;
        RECT 45.300 20.315 46.025 20.495 ;
        RECT 44.780 19.815 45.205 20.145 ;
        RECT 45.375 19.815 46.025 20.315 ;
        RECT 46.195 20.145 46.545 20.665 ;
        RECT 46.715 20.315 46.975 21.285 ;
        RECT 46.195 19.815 46.620 20.145 ;
        RECT 25.525 18.905 30.870 19.450 ;
        RECT 31.045 18.905 36.390 19.450 ;
        RECT 36.565 18.905 37.775 19.655 ;
        RECT 37.945 18.905 38.235 19.630 ;
        RECT 38.405 18.905 41.915 19.675 ;
        RECT 43.200 19.645 43.535 19.815 ;
        RECT 43.780 19.645 44.130 19.815 ;
        RECT 44.780 19.645 45.130 19.815 ;
        RECT 45.375 19.645 45.545 19.815 ;
        RECT 46.195 19.645 46.545 19.815 ;
        RECT 46.790 19.645 46.975 20.315 ;
        RECT 42.545 19.475 43.535 19.645 ;
        RECT 42.545 19.075 42.980 19.475 ;
        RECT 43.150 18.905 43.535 19.305 ;
        RECT 43.705 19.075 44.130 19.645 ;
        RECT 44.320 19.475 45.130 19.645 ;
        RECT 44.320 19.075 44.575 19.475 ;
        RECT 44.745 18.905 45.130 19.305 ;
        RECT 45.300 19.075 45.545 19.645 ;
        RECT 45.735 19.475 46.545 19.645 ;
        RECT 45.735 19.075 45.990 19.475 ;
        RECT 46.160 18.905 46.545 19.305 ;
        RECT 46.715 19.075 46.975 19.645 ;
        RECT 47.145 20.485 47.415 21.255 ;
        RECT 47.585 20.675 47.915 21.455 ;
        RECT 48.120 20.850 48.305 21.255 ;
        RECT 48.475 21.030 48.810 21.455 ;
        RECT 48.120 20.675 48.785 20.850 ;
        RECT 47.145 20.315 48.275 20.485 ;
        RECT 47.145 19.405 47.315 20.315 ;
        RECT 47.485 19.565 47.845 20.145 ;
        RECT 48.025 19.815 48.275 20.315 ;
        RECT 48.445 19.645 48.785 20.675 ;
        RECT 48.990 20.305 49.250 21.455 ;
        RECT 49.425 20.380 49.680 21.285 ;
        RECT 49.850 20.695 50.180 21.455 ;
        RECT 50.395 20.525 50.565 21.285 ;
        RECT 48.100 19.475 48.785 19.645 ;
        RECT 47.145 19.075 47.405 19.405 ;
        RECT 47.615 18.905 47.890 19.385 ;
        RECT 48.100 19.075 48.305 19.475 ;
        RECT 48.475 18.905 48.810 19.305 ;
        RECT 48.990 18.905 49.250 19.745 ;
        RECT 49.425 19.650 49.595 20.380 ;
        RECT 49.850 20.355 50.565 20.525 ;
        RECT 49.850 20.145 50.020 20.355 ;
        RECT 50.825 20.290 51.115 21.455 ;
        RECT 52.210 20.305 52.470 21.455 ;
        RECT 52.645 20.380 52.900 21.285 ;
        RECT 53.070 20.695 53.400 21.455 ;
        RECT 53.615 20.525 53.785 21.285 ;
        RECT 49.765 19.815 50.020 20.145 ;
        RECT 49.425 19.075 49.680 19.650 ;
        RECT 49.850 19.625 50.020 19.815 ;
        RECT 50.300 19.805 50.655 20.175 ;
        RECT 49.850 19.455 50.565 19.625 ;
        RECT 49.850 18.905 50.180 19.285 ;
        RECT 50.395 19.075 50.565 19.455 ;
        RECT 50.825 18.905 51.115 19.630 ;
        RECT 52.210 18.905 52.470 19.745 ;
        RECT 52.645 19.650 52.815 20.380 ;
        RECT 53.070 20.355 53.785 20.525 ;
        RECT 54.045 20.365 55.255 21.455 ;
        RECT 53.070 20.145 53.240 20.355 ;
        RECT 52.985 19.815 53.240 20.145 ;
        RECT 52.645 19.075 52.900 19.650 ;
        RECT 53.070 19.625 53.240 19.815 ;
        RECT 53.520 19.805 53.875 20.175 ;
        RECT 54.045 19.655 54.565 20.195 ;
        RECT 54.735 19.825 55.255 20.365 ;
        RECT 55.425 20.485 55.695 21.255 ;
        RECT 55.865 20.675 56.195 21.455 ;
        RECT 56.400 20.850 56.585 21.255 ;
        RECT 56.755 21.030 57.090 21.455 ;
        RECT 57.265 21.020 62.610 21.455 ;
        RECT 56.400 20.675 57.065 20.850 ;
        RECT 55.425 20.315 56.555 20.485 ;
        RECT 53.070 19.455 53.785 19.625 ;
        RECT 53.070 18.905 53.400 19.285 ;
        RECT 53.615 19.075 53.785 19.455 ;
        RECT 54.045 18.905 55.255 19.655 ;
        RECT 55.425 19.405 55.595 20.315 ;
        RECT 55.765 19.565 56.125 20.145 ;
        RECT 56.305 19.815 56.555 20.315 ;
        RECT 56.725 19.645 57.065 20.675 ;
        RECT 56.380 19.475 57.065 19.645 ;
        RECT 55.425 19.075 55.685 19.405 ;
        RECT 55.895 18.905 56.170 19.385 ;
        RECT 56.380 19.075 56.585 19.475 ;
        RECT 58.850 19.450 59.190 20.280 ;
        RECT 60.670 19.770 61.020 21.020 ;
        RECT 63.705 20.290 63.995 21.455 ;
        RECT 64.165 21.020 69.510 21.455 ;
        RECT 56.755 18.905 57.090 19.305 ;
        RECT 57.265 18.905 62.610 19.450 ;
        RECT 63.705 18.905 63.995 19.630 ;
        RECT 65.750 19.450 66.090 20.280 ;
        RECT 67.570 19.770 67.920 21.020 ;
        RECT 69.685 20.365 71.355 21.455 ;
        RECT 69.685 19.675 70.435 20.195 ;
        RECT 70.605 19.845 71.355 20.365 ;
        RECT 71.530 20.305 71.790 21.455 ;
        RECT 71.965 20.380 72.220 21.285 ;
        RECT 72.390 20.695 72.720 21.455 ;
        RECT 72.935 20.525 73.105 21.285 ;
        RECT 64.165 18.905 69.510 19.450 ;
        RECT 69.685 18.905 71.355 19.675 ;
        RECT 71.530 18.905 71.790 19.745 ;
        RECT 71.965 19.650 72.135 20.380 ;
        RECT 72.390 20.355 73.105 20.525 ;
        RECT 73.365 20.365 74.575 21.455 ;
        RECT 72.390 20.145 72.560 20.355 ;
        RECT 72.305 19.815 72.560 20.145 ;
        RECT 71.965 19.075 72.220 19.650 ;
        RECT 72.390 19.625 72.560 19.815 ;
        RECT 72.840 19.805 73.195 20.175 ;
        RECT 73.365 19.655 73.885 20.195 ;
        RECT 74.055 19.825 74.575 20.365 ;
        RECT 74.750 20.305 75.010 21.455 ;
        RECT 75.185 20.380 75.440 21.285 ;
        RECT 75.610 20.695 75.940 21.455 ;
        RECT 76.155 20.525 76.325 21.285 ;
        RECT 72.390 19.455 73.105 19.625 ;
        RECT 72.390 18.905 72.720 19.285 ;
        RECT 72.935 19.075 73.105 19.455 ;
        RECT 73.365 18.905 74.575 19.655 ;
        RECT 74.750 18.905 75.010 19.745 ;
        RECT 75.185 19.650 75.355 20.380 ;
        RECT 75.610 20.355 76.325 20.525 ;
        RECT 75.610 20.145 75.780 20.355 ;
        RECT 76.585 20.290 76.875 21.455 ;
        RECT 77.970 20.305 78.230 21.455 ;
        RECT 78.405 20.380 78.660 21.285 ;
        RECT 78.830 20.695 79.160 21.455 ;
        RECT 79.375 20.525 79.545 21.285 ;
        RECT 75.525 19.815 75.780 20.145 ;
        RECT 75.185 19.075 75.440 19.650 ;
        RECT 75.610 19.625 75.780 19.815 ;
        RECT 76.060 19.805 76.415 20.175 ;
        RECT 75.610 19.455 76.325 19.625 ;
        RECT 75.610 18.905 75.940 19.285 ;
        RECT 76.155 19.075 76.325 19.455 ;
        RECT 76.585 18.905 76.875 19.630 ;
        RECT 77.970 18.905 78.230 19.745 ;
        RECT 78.405 19.650 78.575 20.380 ;
        RECT 78.830 20.355 79.545 20.525 ;
        RECT 79.895 20.525 80.065 21.285 ;
        RECT 80.280 20.695 80.610 21.455 ;
        RECT 79.895 20.355 80.610 20.525 ;
        RECT 80.780 20.380 81.035 21.285 ;
        RECT 78.830 20.145 79.000 20.355 ;
        RECT 78.745 19.815 79.000 20.145 ;
        RECT 78.405 19.075 78.660 19.650 ;
        RECT 78.830 19.625 79.000 19.815 ;
        RECT 79.280 19.805 79.635 20.175 ;
        RECT 79.805 19.805 80.160 20.175 ;
        RECT 80.440 20.145 80.610 20.355 ;
        RECT 80.440 19.815 80.695 20.145 ;
        RECT 80.440 19.625 80.610 19.815 ;
        RECT 80.865 19.650 81.035 20.380 ;
        RECT 81.210 20.305 81.470 21.455 ;
        RECT 81.735 20.525 81.905 21.285 ;
        RECT 82.120 20.695 82.450 21.455 ;
        RECT 81.735 20.355 82.450 20.525 ;
        RECT 82.620 20.380 82.875 21.285 ;
        RECT 81.645 19.805 82.000 20.175 ;
        RECT 82.280 20.145 82.450 20.355 ;
        RECT 82.280 19.815 82.535 20.145 ;
        RECT 78.830 19.455 79.545 19.625 ;
        RECT 78.830 18.905 79.160 19.285 ;
        RECT 79.375 19.075 79.545 19.455 ;
        RECT 79.895 19.455 80.610 19.625 ;
        RECT 79.895 19.075 80.065 19.455 ;
        RECT 80.280 18.905 80.610 19.285 ;
        RECT 80.780 19.075 81.035 19.650 ;
        RECT 81.210 18.905 81.470 19.745 ;
        RECT 82.280 19.625 82.450 19.815 ;
        RECT 82.705 19.650 82.875 20.380 ;
        RECT 83.050 20.305 83.310 21.455 ;
        RECT 83.670 20.485 84.060 20.660 ;
        RECT 84.545 20.655 84.875 21.455 ;
        RECT 85.045 20.665 85.580 21.285 ;
        RECT 83.670 20.315 85.095 20.485 ;
        RECT 81.735 19.455 82.450 19.625 ;
        RECT 81.735 19.075 81.905 19.455 ;
        RECT 82.120 18.905 82.450 19.285 ;
        RECT 82.620 19.075 82.875 19.650 ;
        RECT 83.050 18.905 83.310 19.745 ;
        RECT 83.545 19.585 83.900 20.145 ;
        RECT 84.070 19.415 84.240 20.315 ;
        RECT 84.410 19.585 84.675 20.145 ;
        RECT 84.925 19.815 85.095 20.315 ;
        RECT 85.265 19.645 85.580 20.665 ;
        RECT 86.795 20.525 86.965 21.285 ;
        RECT 87.180 20.695 87.510 21.455 ;
        RECT 86.795 20.355 87.510 20.525 ;
        RECT 87.680 20.380 87.935 21.285 ;
        RECT 86.705 19.805 87.060 20.175 ;
        RECT 87.340 20.145 87.510 20.355 ;
        RECT 87.340 19.815 87.595 20.145 ;
        RECT 83.650 18.905 83.890 19.415 ;
        RECT 84.070 19.085 84.350 19.415 ;
        RECT 84.580 18.905 84.795 19.415 ;
        RECT 84.965 19.075 85.580 19.645 ;
        RECT 87.340 19.625 87.510 19.815 ;
        RECT 87.765 19.650 87.935 20.380 ;
        RECT 88.110 20.305 88.370 21.455 ;
        RECT 88.545 20.365 89.755 21.455 ;
        RECT 88.545 19.825 89.065 20.365 ;
        RECT 86.795 19.455 87.510 19.625 ;
        RECT 86.795 19.075 86.965 19.455 ;
        RECT 87.180 18.905 87.510 19.285 ;
        RECT 87.680 19.075 87.935 19.650 ;
        RECT 88.110 18.905 88.370 19.745 ;
        RECT 89.235 19.655 89.755 20.195 ;
        RECT 88.545 18.905 89.755 19.655 ;
        RECT 12.100 18.735 89.840 18.905 ;
      LAYER met1 ;
        RECT 118.795 224.800 119.455 225.215 ;
        RECT 121.530 224.805 122.190 225.455 ;
        RECT 124.275 224.945 124.935 225.595 ;
        RECT 127.145 224.965 127.805 225.615 ;
        RECT 95.405 224.565 119.455 224.800 ;
        RECT 95.405 224.555 119.270 224.565 ;
        RECT 95.405 217.665 95.650 224.555 ;
        RECT 121.680 224.145 121.980 224.805 ;
        RECT 96.145 223.845 121.980 224.145 ;
        RECT 95.365 217.405 95.685 217.665 ;
        RECT 96.145 216.895 96.445 223.845 ;
        RECT 124.430 223.590 124.715 224.945 ;
        RECT 96.825 223.305 124.715 223.590 ;
        RECT 96.825 217.525 97.110 223.305 ;
        RECT 127.305 222.970 127.570 224.965 ;
        RECT 129.605 224.960 130.265 225.610 ;
        RECT 97.505 222.705 127.570 222.970 ;
        RECT 96.795 217.240 97.140 217.525 ;
        RECT 97.505 216.905 97.770 222.705 ;
        RECT 129.710 222.425 129.980 224.960 ;
        RECT 132.985 224.945 133.645 225.595 ;
        RECT 134.915 225.075 135.575 225.725 ;
        RECT 137.630 225.315 138.410 225.575 ;
        RECT 98.170 222.155 129.980 222.425 ;
        RECT 98.170 217.640 98.440 222.155 ;
        RECT 133.185 222.000 133.395 224.945 ;
        RECT 98.780 221.790 133.395 222.000 ;
        RECT 98.140 217.370 98.470 217.640 ;
        RECT 98.780 217.055 98.990 221.790 ;
        RECT 135.070 221.535 135.285 225.075 ;
        RECT 137.630 224.895 138.580 225.315 ;
        RECT 99.230 221.320 135.285 221.535 ;
        RECT 99.230 217.630 99.445 221.320 ;
        RECT 138.345 221.075 138.580 224.895 ;
        RECT 149.710 221.830 149.970 222.150 ;
        RECT 99.715 220.840 138.580 221.075 ;
        RECT 99.175 217.370 99.495 217.630 ;
        RECT 99.715 217.080 99.950 220.840 ;
        RECT 149.150 220.770 149.410 221.090 ;
        RECT 115.800 220.285 116.060 220.605 ;
        RECT 96.115 216.595 96.475 216.895 ;
        RECT 97.475 216.640 97.800 216.905 ;
        RECT 98.725 216.795 99.045 217.055 ;
        RECT 99.670 216.820 99.990 217.080 ;
        RECT 110.950 206.310 111.210 206.630 ;
        RECT 109.950 205.860 110.210 206.180 ;
        RECT 110.010 192.545 110.150 205.860 ;
        RECT 111.010 201.530 111.150 206.310 ;
        RECT 111.360 205.830 111.620 206.150 ;
        RECT 111.420 202.635 111.560 205.830 ;
        RECT 111.330 202.375 111.650 202.635 ;
        RECT 111.010 201.390 111.640 201.530 ;
        RECT 111.500 198.530 111.640 201.390 ;
        RECT 111.410 198.200 111.740 198.530 ;
        RECT 109.950 192.225 110.210 192.545 ;
        RECT 100.970 182.410 102.630 184.070 ;
        RECT 112.120 183.415 112.600 219.295 ;
        RECT 113.420 207.865 113.680 208.185 ;
        RECT 112.755 206.960 112.985 207.250 ;
        RECT 112.800 205.425 112.940 206.960 ;
        RECT 112.740 205.105 113.000 205.425 ;
        RECT 112.755 204.660 112.985 204.950 ;
        RECT 112.800 202.665 112.940 204.660 ;
        RECT 113.435 203.955 113.665 204.030 ;
        RECT 113.435 203.815 114.640 203.955 ;
        RECT 113.435 203.740 113.665 203.815 ;
        RECT 113.435 203.280 113.665 203.570 ;
        RECT 113.480 203.125 113.620 203.280 ;
        RECT 113.420 202.805 113.680 203.125 ;
        RECT 114.115 202.795 114.345 203.085 ;
        RECT 112.740 202.345 113.000 202.665 ;
        RECT 113.775 202.400 114.005 202.690 ;
        RECT 113.095 201.945 113.325 202.235 ;
        RECT 113.140 200.825 113.280 201.945 ;
        RECT 113.820 201.500 113.960 202.400 ;
        RECT 113.775 201.210 114.005 201.500 ;
        RECT 113.080 200.505 113.340 200.825 ;
        RECT 113.820 198.980 113.960 201.210 ;
        RECT 114.160 200.985 114.300 202.795 ;
        RECT 114.115 200.695 114.345 200.985 ;
        RECT 114.160 199.415 114.300 200.695 ;
        RECT 114.115 199.125 114.345 199.415 ;
        RECT 113.775 198.690 114.005 198.980 ;
        RECT 112.740 198.435 113.000 198.525 ;
        RECT 112.740 198.295 113.280 198.435 ;
        RECT 112.740 198.205 113.000 198.295 ;
        RECT 112.755 195.675 112.985 195.750 ;
        RECT 113.140 195.675 113.280 198.295 ;
        RECT 114.500 198.065 114.640 203.815 ;
        RECT 114.440 197.745 114.700 198.065 ;
        RECT 114.115 196.380 114.345 196.670 ;
        RECT 112.755 195.535 113.280 195.675 ;
        RECT 112.755 195.460 112.985 195.535 ;
        RECT 114.160 194.845 114.300 196.380 ;
        RECT 113.420 194.525 113.680 194.845 ;
        RECT 114.100 194.525 114.360 194.845 ;
        RECT 112.740 192.225 113.000 192.545 ;
        RECT 112.800 191.150 112.940 192.225 ;
        RECT 113.420 191.765 113.680 192.085 ;
        RECT 112.755 190.860 112.985 191.150 ;
        RECT 114.455 189.940 114.685 190.230 ;
        RECT 113.760 189.465 114.020 189.785 ;
        RECT 113.420 189.005 113.680 189.325 ;
        RECT 113.820 187.930 113.960 189.465 ;
        RECT 114.100 188.545 114.360 188.865 ;
        RECT 113.775 187.640 114.005 187.930 ;
        RECT 114.160 186.550 114.300 188.545 ;
        RECT 114.500 188.405 114.640 189.940 ;
        RECT 114.440 188.085 114.700 188.405 ;
        RECT 114.115 186.260 114.345 186.550 ;
        RECT 114.440 185.785 114.700 186.105 ;
        RECT 114.500 185.630 114.640 185.785 ;
        RECT 114.455 185.340 114.685 185.630 ;
        RECT 114.840 183.415 115.320 219.295 ;
        RECT 115.860 217.370 116.000 220.285 ;
        RECT 148.630 220.050 148.950 220.310 ;
        RECT 148.140 219.570 148.400 219.890 ;
        RECT 116.480 217.525 116.740 217.845 ;
        RECT 115.815 217.080 116.045 217.370 ;
        RECT 116.540 216.450 116.680 217.525 ;
        RECT 116.495 216.160 116.725 216.450 ;
        RECT 117.160 214.765 117.420 215.085 ;
        RECT 117.160 212.925 117.420 213.245 ;
        RECT 117.160 212.465 117.420 212.785 ;
        RECT 116.155 211.560 116.385 211.850 ;
        RECT 116.200 206.345 116.340 211.560 ;
        RECT 117.160 210.165 117.420 210.485 ;
        RECT 117.220 208.185 117.360 210.165 ;
        RECT 117.160 207.865 117.420 208.185 ;
        RECT 116.140 206.025 116.400 206.345 ;
        RECT 117.220 205.870 117.360 207.865 ;
        RECT 117.175 205.580 117.405 205.870 ;
        RECT 116.155 203.270 116.385 203.560 ;
        RECT 115.815 202.835 116.045 203.125 ;
        RECT 115.860 201.555 116.000 202.835 ;
        RECT 115.815 201.265 116.045 201.555 ;
        RECT 115.460 200.505 115.720 200.825 ;
        RECT 115.520 198.510 115.660 200.505 ;
        RECT 115.860 199.455 116.000 201.265 ;
        RECT 116.200 201.040 116.340 203.270 ;
        RECT 117.160 201.655 117.420 201.745 ;
        RECT 116.540 201.515 117.420 201.655 ;
        RECT 116.155 200.750 116.385 201.040 ;
        RECT 116.200 199.850 116.340 200.750 ;
        RECT 116.540 200.305 116.680 201.515 ;
        RECT 117.160 201.425 117.420 201.515 ;
        RECT 116.820 200.505 117.080 200.825 ;
        RECT 116.495 200.015 116.725 200.305 ;
        RECT 116.155 199.560 116.385 199.850 ;
        RECT 115.815 199.165 116.045 199.455 ;
        RECT 116.495 198.895 116.725 198.970 ;
        RECT 116.880 198.895 117.020 200.505 ;
        RECT 116.495 198.755 117.020 198.895 ;
        RECT 116.495 198.680 116.725 198.755 ;
        RECT 115.475 198.220 115.705 198.510 ;
        RECT 116.495 196.380 116.725 196.670 ;
        RECT 116.140 194.985 116.400 195.305 ;
        RECT 116.140 194.525 116.400 194.845 ;
        RECT 116.200 190.230 116.340 194.525 ;
        RECT 116.540 192.990 116.680 196.380 ;
        RECT 117.160 195.905 117.420 196.225 ;
        RECT 116.495 192.700 116.725 192.990 ;
        RECT 116.155 189.940 116.385 190.230 ;
        RECT 116.140 189.465 116.400 189.785 ;
        RECT 116.200 188.390 116.340 189.465 ;
        RECT 116.480 189.005 116.740 189.325 ;
        RECT 116.155 188.100 116.385 188.390 ;
        RECT 116.155 187.640 116.385 187.930 ;
        RECT 116.200 185.185 116.340 187.640 ;
        RECT 116.540 187.010 116.680 189.005 ;
        RECT 116.495 186.720 116.725 187.010 ;
        RECT 117.160 186.245 117.420 186.565 ;
        RECT 117.220 186.090 117.360 186.245 ;
        RECT 117.175 185.800 117.405 186.090 ;
        RECT 116.140 184.865 116.400 185.185 ;
        RECT 117.560 183.415 118.040 219.295 ;
        RECT 119.880 217.525 120.140 217.845 ;
        RECT 119.215 215.230 119.445 215.520 ;
        RECT 118.520 214.765 118.780 215.085 ;
        RECT 118.580 212.265 118.720 214.765 ;
        RECT 119.260 213.000 119.400 215.230 ;
        RECT 119.555 214.795 119.785 215.085 ;
        RECT 119.600 213.515 119.740 214.795 ;
        RECT 119.555 213.225 119.785 213.515 ;
        RECT 119.215 212.710 119.445 213.000 ;
        RECT 118.535 211.975 118.765 212.265 ;
        RECT 119.260 211.810 119.400 212.710 ;
        RECT 119.215 211.520 119.445 211.810 ;
        RECT 119.600 211.415 119.740 213.225 ;
        RECT 119.555 211.125 119.785 211.415 ;
        RECT 119.200 210.625 119.460 210.945 ;
        RECT 118.875 205.580 119.105 205.870 ;
        RECT 118.920 201.285 119.060 205.580 ;
        RECT 118.860 200.965 119.120 201.285 ;
        RECT 119.880 200.505 120.140 200.825 ;
        RECT 119.940 199.430 120.080 200.505 ;
        RECT 119.895 199.140 120.125 199.430 ;
        RECT 118.875 195.215 119.105 195.290 ;
        RECT 118.875 195.075 119.400 195.215 ;
        RECT 118.875 195.000 119.105 195.075 ;
        RECT 118.860 193.605 119.120 193.925 ;
        RECT 118.195 192.915 118.425 192.990 ;
        RECT 118.195 192.775 118.720 192.915 ;
        RECT 118.195 192.700 118.425 192.775 ;
        RECT 118.195 189.940 118.425 190.230 ;
        RECT 118.240 189.785 118.380 189.940 ;
        RECT 118.180 189.465 118.440 189.785 ;
        RECT 118.580 189.695 118.720 192.775 ;
        RECT 118.860 192.225 119.120 192.545 ;
        RECT 118.860 190.845 119.120 191.165 ;
        RECT 118.875 189.695 119.105 189.770 ;
        RECT 118.580 189.555 119.105 189.695 ;
        RECT 118.180 189.005 118.440 189.325 ;
        RECT 118.580 187.395 118.720 189.555 ;
        RECT 118.875 189.480 119.105 189.555 ;
        RECT 118.875 188.560 119.105 188.850 ;
        RECT 118.920 188.405 119.060 188.560 ;
        RECT 118.860 188.085 119.120 188.405 ;
        RECT 118.860 187.395 119.120 187.485 ;
        RECT 118.580 187.255 119.120 187.395 ;
        RECT 118.860 187.165 119.120 187.255 ;
        RECT 118.860 185.785 119.120 186.105 ;
        RECT 119.260 185.645 119.400 195.075 ;
        RECT 119.555 194.080 119.785 194.370 ;
        RECT 119.600 188.865 119.740 194.080 ;
        RECT 119.895 191.320 120.125 191.610 ;
        RECT 119.940 189.325 120.080 191.320 ;
        RECT 119.880 189.005 120.140 189.325 ;
        RECT 119.540 188.545 119.800 188.865 ;
        RECT 119.895 188.100 120.125 188.390 ;
        RECT 119.940 187.945 120.080 188.100 ;
        RECT 119.880 187.625 120.140 187.945 ;
        RECT 119.200 185.325 119.460 185.645 ;
        RECT 118.860 184.865 119.120 185.185 ;
        RECT 120.280 183.415 120.760 219.295 ;
        RECT 121.240 217.985 121.500 218.305 ;
        RECT 121.300 217.370 121.440 217.985 ;
        RECT 121.580 217.525 121.840 217.845 ;
        RECT 121.255 217.080 121.485 217.370 ;
        RECT 121.640 215.070 121.780 217.525 ;
        RECT 121.935 216.160 122.165 216.450 ;
        RECT 121.595 214.780 121.825 215.070 ;
        RECT 120.900 212.925 121.160 213.245 ;
        RECT 120.960 211.850 121.100 212.925 ;
        RECT 121.240 212.465 121.500 212.785 ;
        RECT 120.915 211.560 121.145 211.850 ;
        RECT 120.915 202.820 121.145 203.110 ;
        RECT 120.960 201.745 121.100 202.820 ;
        RECT 120.900 201.425 121.160 201.745 ;
        RECT 121.300 200.735 121.440 212.465 ;
        RECT 121.580 210.165 121.840 210.485 ;
        RECT 121.980 210.025 122.120 216.160 ;
        RECT 121.920 209.705 122.180 210.025 ;
        RECT 121.935 206.960 122.165 207.250 ;
        RECT 121.580 206.025 121.840 206.345 ;
        RECT 121.595 205.120 121.825 205.410 ;
        RECT 121.640 201.195 121.780 205.120 ;
        RECT 121.980 204.950 122.120 206.960 ;
        RECT 121.935 204.660 122.165 204.950 ;
        RECT 121.640 201.055 122.460 201.195 ;
        RECT 120.960 200.595 121.440 200.735 ;
        RECT 120.960 194.385 121.100 200.595 ;
        RECT 121.920 200.505 122.180 200.825 ;
        RECT 121.255 200.035 121.485 200.325 ;
        RECT 121.300 198.225 121.440 200.035 ;
        RECT 121.595 199.640 121.825 199.930 ;
        RECT 121.640 198.740 121.780 199.640 ;
        RECT 121.935 199.185 122.165 199.475 ;
        RECT 121.595 198.450 121.825 198.740 ;
        RECT 121.255 197.935 121.485 198.225 ;
        RECT 121.300 196.655 121.440 197.935 ;
        RECT 121.255 196.365 121.485 196.655 ;
        RECT 121.640 196.220 121.780 198.450 ;
        RECT 121.595 195.930 121.825 196.220 ;
        RECT 121.980 195.675 122.120 199.185 ;
        RECT 122.320 196.225 122.460 201.055 ;
        RECT 122.260 195.905 122.520 196.225 ;
        RECT 121.300 195.535 122.120 195.675 ;
        RECT 120.900 194.065 121.160 194.385 ;
        RECT 120.915 193.620 121.145 193.910 ;
        RECT 120.960 192.085 121.100 193.620 ;
        RECT 121.300 192.990 121.440 195.535 ;
        RECT 121.920 194.985 122.180 195.305 ;
        RECT 121.580 194.065 121.840 194.385 ;
        RECT 121.255 192.700 121.485 192.990 ;
        RECT 120.900 191.765 121.160 192.085 ;
        RECT 121.640 190.690 121.780 194.065 ;
        RECT 121.595 190.400 121.825 190.690 ;
        RECT 121.595 190.155 121.825 190.230 ;
        RECT 121.980 190.155 122.120 194.985 ;
        RECT 122.600 190.845 122.860 191.165 ;
        RECT 121.595 190.015 122.120 190.155 ;
        RECT 121.595 189.940 121.825 190.015 ;
        RECT 121.580 189.005 121.840 189.325 ;
        RECT 120.900 188.085 121.160 188.405 ;
        RECT 120.960 186.550 121.100 188.085 ;
        RECT 121.255 187.640 121.485 187.930 ;
        RECT 120.915 186.260 121.145 186.550 ;
        RECT 121.300 185.185 121.440 187.640 ;
        RECT 121.640 186.105 121.780 189.005 ;
        RECT 121.920 188.545 122.180 188.865 ;
        RECT 121.920 187.165 122.180 187.485 ;
        RECT 122.600 187.165 122.860 187.485 ;
        RECT 121.980 186.550 122.120 187.165 ;
        RECT 122.260 186.705 122.520 187.025 ;
        RECT 121.935 186.260 122.165 186.550 ;
        RECT 121.580 185.785 121.840 186.105 ;
        RECT 121.240 184.865 121.500 185.185 ;
        RECT 122.320 185.170 122.460 186.705 ;
        RECT 122.275 184.880 122.505 185.170 ;
        RECT 123.000 183.415 123.480 219.295 ;
        RECT 124.640 217.755 124.900 217.845 ;
        RECT 124.360 217.615 124.900 217.755 ;
        RECT 123.975 216.205 124.205 216.495 ;
        RECT 124.020 215.545 124.160 216.205 ;
        RECT 123.960 215.225 124.220 215.545 ;
        RECT 124.360 210.945 124.500 217.615 ;
        RECT 124.640 217.525 124.900 217.615 ;
        RECT 124.995 217.055 125.225 217.345 ;
        RECT 124.655 216.660 124.885 216.950 ;
        RECT 124.700 215.760 124.840 216.660 ;
        RECT 124.655 215.470 124.885 215.760 ;
        RECT 124.700 213.240 124.840 215.470 ;
        RECT 125.040 215.245 125.180 217.055 ;
        RECT 124.995 214.955 125.225 215.245 ;
        RECT 125.040 213.675 125.180 214.955 ;
        RECT 124.995 213.385 125.225 213.675 ;
        RECT 124.655 212.950 124.885 213.240 ;
        RECT 124.300 210.625 124.560 210.945 ;
        RECT 125.335 210.640 125.565 210.930 ;
        RECT 124.360 205.870 124.500 210.625 ;
        RECT 125.380 210.025 125.520 210.640 ;
        RECT 125.320 209.705 125.580 210.025 ;
        RECT 124.315 205.795 124.545 205.870 ;
        RECT 123.680 205.655 124.545 205.795 ;
        RECT 123.680 200.825 123.820 205.655 ;
        RECT 124.315 205.580 124.545 205.655 ;
        RECT 124.995 205.095 125.225 205.385 ;
        RECT 123.960 204.645 124.220 204.965 ;
        RECT 124.655 204.700 124.885 204.990 ;
        RECT 124.020 204.415 124.160 204.645 ;
        RECT 124.315 204.415 124.545 204.535 ;
        RECT 124.020 204.275 124.545 204.415 ;
        RECT 124.315 204.245 124.545 204.275 ;
        RECT 124.700 203.800 124.840 204.700 ;
        RECT 124.655 203.510 124.885 203.800 ;
        RECT 124.700 201.280 124.840 203.510 ;
        RECT 125.040 203.285 125.180 205.095 ;
        RECT 124.995 202.995 125.225 203.285 ;
        RECT 125.040 201.715 125.180 202.995 ;
        RECT 124.995 201.425 125.225 201.715 ;
        RECT 124.655 200.990 124.885 201.280 ;
        RECT 123.620 200.505 123.880 200.825 ;
        RECT 123.635 198.680 123.865 198.970 ;
        RECT 123.680 198.065 123.820 198.680 ;
        RECT 124.655 198.220 124.885 198.510 ;
        RECT 123.620 197.745 123.880 198.065 ;
        RECT 124.700 197.605 124.840 198.220 ;
        RECT 124.640 197.285 124.900 197.605 ;
        RECT 124.980 196.365 125.240 196.685 ;
        RECT 125.335 195.920 125.565 196.210 ;
        RECT 125.380 195.305 125.520 195.920 ;
        RECT 125.320 194.985 125.580 195.305 ;
        RECT 124.300 191.765 124.560 192.085 ;
        RECT 123.620 190.845 123.880 191.165 ;
        RECT 123.680 188.850 123.820 190.845 ;
        RECT 124.640 189.465 124.900 189.785 ;
        RECT 124.300 189.005 124.560 189.325 ;
        RECT 123.635 188.560 123.865 188.850 ;
        RECT 124.360 187.470 124.500 189.005 ;
        RECT 124.315 187.180 124.545 187.470 ;
        RECT 124.300 186.705 124.560 187.025 ;
        RECT 124.300 186.245 124.560 186.565 ;
        RECT 124.315 186.015 124.545 186.090 ;
        RECT 124.700 186.015 124.840 189.465 ;
        RECT 125.320 189.005 125.580 189.325 ;
        RECT 125.380 188.390 125.520 189.005 ;
        RECT 125.335 188.100 125.565 188.390 ;
        RECT 124.315 185.875 124.840 186.015 ;
        RECT 124.315 185.800 124.545 185.875 ;
        RECT 125.720 183.415 126.200 219.295 ;
        RECT 128.040 217.985 128.300 218.305 ;
        RECT 126.680 217.525 126.940 217.845 ;
        RECT 127.360 217.525 127.620 217.845 ;
        RECT 126.340 215.225 126.600 215.545 ;
        RECT 126.740 211.315 126.880 217.525 ;
        RECT 127.420 216.450 127.560 217.525 ;
        RECT 128.100 217.370 128.240 217.985 ;
        RECT 128.055 217.080 128.285 217.370 ;
        RECT 127.375 216.160 127.605 216.450 ;
        RECT 128.055 213.400 128.285 213.690 ;
        RECT 127.035 212.940 127.265 213.230 ;
        RECT 127.080 212.785 127.220 212.940 ;
        RECT 128.100 212.785 128.240 213.400 ;
        RECT 127.020 212.465 127.280 212.785 ;
        RECT 128.040 212.465 128.300 212.785 ;
        RECT 127.020 212.005 127.280 212.325 ;
        RECT 127.035 211.315 127.265 211.390 ;
        RECT 126.740 211.175 127.265 211.315 ;
        RECT 127.035 211.100 127.265 211.175 ;
        RECT 126.695 210.615 126.925 210.905 ;
        RECT 126.740 208.805 126.880 210.615 ;
        RECT 127.035 210.220 127.265 210.510 ;
        RECT 127.080 209.320 127.220 210.220 ;
        RECT 127.715 209.765 127.945 210.055 ;
        RECT 127.035 209.030 127.265 209.320 ;
        RECT 126.695 208.515 126.925 208.805 ;
        RECT 126.740 207.235 126.880 208.515 ;
        RECT 126.695 206.945 126.925 207.235 ;
        RECT 127.080 206.800 127.220 209.030 ;
        RECT 127.035 206.510 127.265 206.800 ;
        RECT 127.760 206.345 127.900 209.765 ;
        RECT 127.700 206.025 127.960 206.345 ;
        RECT 127.760 204.965 127.900 206.025 ;
        RECT 126.680 204.645 126.940 204.965 ;
        RECT 127.700 204.645 127.960 204.965 ;
        RECT 126.740 204.030 126.880 204.645 ;
        RECT 128.040 204.185 128.300 204.505 ;
        RECT 126.695 203.740 126.925 204.030 ;
        RECT 127.375 201.900 127.605 202.190 ;
        RECT 127.035 201.655 127.265 201.730 ;
        RECT 126.740 201.515 127.265 201.655 ;
        RECT 126.740 196.225 126.880 201.515 ;
        RECT 127.035 201.440 127.265 201.515 ;
        RECT 127.035 200.520 127.265 200.810 ;
        RECT 127.080 198.525 127.220 200.520 ;
        RECT 127.420 199.890 127.560 201.900 ;
        RECT 127.375 199.600 127.605 199.890 ;
        RECT 127.020 198.205 127.280 198.525 ;
        RECT 127.020 197.745 127.280 198.065 ;
        RECT 127.080 197.130 127.220 197.745 ;
        RECT 128.100 197.605 128.240 204.185 ;
        RECT 128.040 197.285 128.300 197.605 ;
        RECT 127.035 196.840 127.265 197.130 ;
        RECT 126.680 195.905 126.940 196.225 ;
        RECT 126.740 190.230 126.880 195.905 ;
        RECT 127.360 193.605 127.620 193.925 ;
        RECT 127.420 192.530 127.560 193.605 ;
        RECT 127.375 192.240 127.605 192.530 ;
        RECT 127.375 191.995 127.605 192.070 ;
        RECT 127.375 191.855 127.900 191.995 ;
        RECT 127.375 191.780 127.605 191.855 ;
        RECT 127.360 191.305 127.620 191.625 ;
        RECT 127.035 190.860 127.265 191.150 ;
        RECT 126.695 189.940 126.925 190.230 ;
        RECT 127.080 187.485 127.220 190.860 ;
        RECT 127.760 189.785 127.900 191.855 ;
        RECT 127.700 189.465 127.960 189.785 ;
        RECT 127.375 188.560 127.605 188.850 ;
        RECT 127.420 188.405 127.560 188.560 ;
        RECT 127.360 188.085 127.620 188.405 ;
        RECT 127.360 187.625 127.620 187.945 ;
        RECT 128.040 187.625 128.300 187.945 ;
        RECT 127.020 187.165 127.280 187.485 ;
        RECT 127.375 186.260 127.605 186.550 ;
        RECT 127.420 186.105 127.560 186.260 ;
        RECT 127.360 185.785 127.620 186.105 ;
        RECT 128.100 185.630 128.240 187.625 ;
        RECT 128.055 185.340 128.285 185.630 ;
        RECT 128.440 183.415 128.920 219.295 ;
        RECT 130.080 217.525 130.340 217.845 ;
        RECT 130.140 216.450 130.280 217.525 ;
        RECT 130.095 216.160 130.325 216.450 ;
        RECT 130.760 212.925 131.020 213.245 ;
        RECT 129.060 212.465 129.320 212.785 ;
        RECT 129.740 209.705 130.000 210.025 ;
        RECT 129.755 205.795 129.985 205.870 ;
        RECT 129.460 205.655 129.985 205.795 ;
        RECT 129.460 200.350 129.600 205.655 ;
        RECT 129.755 205.580 129.985 205.655 ;
        RECT 129.755 204.875 129.985 204.950 ;
        RECT 129.755 204.735 130.280 204.875 ;
        RECT 129.755 204.660 129.985 204.735 ;
        RECT 129.740 204.185 130.000 204.505 ;
        RECT 130.140 203.495 130.280 204.735 ;
        RECT 130.760 204.645 131.020 204.965 ;
        RECT 130.760 204.185 131.020 204.505 ;
        RECT 130.435 203.495 130.665 203.570 ;
        RECT 130.140 203.355 130.665 203.495 ;
        RECT 130.435 203.280 130.665 203.355 ;
        RECT 130.095 202.820 130.325 203.110 ;
        RECT 129.755 201.900 129.985 202.190 ;
        RECT 129.800 201.745 129.940 201.900 ;
        RECT 129.740 201.425 130.000 201.745 ;
        RECT 129.740 200.505 130.000 200.825 ;
        RECT 129.415 200.060 129.645 200.350 ;
        RECT 130.140 197.515 130.280 202.820 ;
        RECT 130.480 200.365 130.620 203.280 ;
        RECT 130.820 202.650 130.960 204.185 ;
        RECT 130.775 202.360 131.005 202.650 ;
        RECT 130.420 200.045 130.680 200.365 ;
        RECT 130.140 197.375 130.620 197.515 ;
        RECT 130.080 196.825 130.340 197.145 ;
        RECT 130.480 196.225 130.620 197.375 ;
        RECT 130.420 195.905 130.680 196.225 ;
        RECT 129.075 195.000 129.305 195.290 ;
        RECT 129.120 194.385 129.260 195.000 ;
        RECT 129.060 194.065 129.320 194.385 ;
        RECT 129.755 194.295 129.985 194.370 ;
        RECT 129.755 194.155 130.280 194.295 ;
        RECT 129.755 194.080 129.985 194.155 ;
        RECT 129.755 193.160 129.985 193.450 ;
        RECT 129.415 191.780 129.645 192.070 ;
        RECT 129.060 191.305 129.320 191.625 ;
        RECT 129.120 191.150 129.260 191.305 ;
        RECT 129.075 190.860 129.305 191.150 ;
        RECT 129.460 189.785 129.600 191.780 ;
        RECT 129.800 191.610 129.940 193.160 ;
        RECT 129.755 191.320 129.985 191.610 ;
        RECT 129.800 191.165 129.940 191.320 ;
        RECT 129.740 190.845 130.000 191.165 ;
        RECT 129.755 190.615 129.985 190.690 ;
        RECT 130.140 190.615 130.280 194.155 ;
        RECT 130.760 193.605 131.020 193.925 ;
        RECT 129.755 190.475 130.280 190.615 ;
        RECT 129.755 190.400 129.985 190.475 ;
        RECT 129.740 189.925 130.000 190.245 ;
        RECT 129.400 189.465 129.660 189.785 ;
        RECT 129.075 189.235 129.305 189.310 ;
        RECT 129.075 189.095 129.600 189.235 ;
        RECT 129.075 189.020 129.305 189.095 ;
        RECT 129.460 188.775 129.600 189.095 ;
        RECT 129.755 188.775 129.985 188.850 ;
        RECT 129.460 188.635 129.985 188.775 ;
        RECT 129.460 187.025 129.600 188.635 ;
        RECT 129.755 188.560 129.985 188.635 ;
        RECT 129.740 187.625 130.000 187.945 ;
        RECT 130.140 187.855 130.280 190.475 ;
        RECT 130.420 187.855 130.680 187.945 ;
        RECT 130.140 187.715 130.680 187.855 ;
        RECT 130.420 187.625 130.680 187.715 ;
        RECT 129.740 187.165 130.000 187.485 ;
        RECT 129.400 186.705 129.660 187.025 ;
        RECT 129.800 186.550 129.940 187.165 ;
        RECT 129.755 186.260 129.985 186.550 ;
        RECT 130.760 186.245 131.020 186.565 ;
        RECT 130.820 185.630 130.960 186.245 ;
        RECT 130.775 185.340 131.005 185.630 ;
        RECT 131.160 183.415 131.640 219.295 ;
        RECT 131.780 217.525 132.040 217.845 ;
        RECT 133.140 217.525 133.400 217.845 ;
        RECT 132.475 215.230 132.705 215.520 ;
        RECT 132.135 214.795 132.365 215.085 ;
        RECT 132.180 213.515 132.320 214.795 ;
        RECT 132.135 213.225 132.365 213.515 ;
        RECT 132.180 211.415 132.320 213.225 ;
        RECT 132.520 213.000 132.660 215.230 ;
        RECT 132.475 212.710 132.705 213.000 ;
        RECT 132.520 211.810 132.660 212.710 ;
        RECT 133.200 212.265 133.340 217.525 ;
        RECT 133.155 211.975 133.385 212.265 ;
        RECT 132.475 211.520 132.705 211.810 ;
        RECT 132.135 211.125 132.365 211.415 ;
        RECT 132.800 210.625 133.060 210.945 ;
        RECT 133.140 206.945 133.400 207.265 ;
        RECT 131.780 200.965 132.040 201.285 ;
        RECT 131.840 200.810 131.980 200.965 ;
        RECT 131.795 200.520 132.025 200.810 ;
        RECT 132.460 200.505 132.720 200.825 ;
        RECT 131.780 195.905 132.040 196.225 ;
        RECT 131.840 192.990 131.980 195.905 ;
        RECT 132.520 195.290 132.660 200.505 ;
        RECT 133.480 197.745 133.740 198.065 ;
        RECT 133.480 195.445 133.740 195.765 ;
        RECT 132.475 195.000 132.705 195.290 ;
        RECT 131.795 192.700 132.025 192.990 ;
        RECT 132.800 192.685 133.060 193.005 ;
        RECT 132.800 191.765 133.060 192.085 ;
        RECT 133.540 191.150 133.680 195.445 ;
        RECT 133.495 190.860 133.725 191.150 ;
        RECT 131.780 189.465 132.040 189.785 ;
        RECT 131.840 186.550 131.980 189.465 ;
        RECT 132.800 187.395 133.060 187.485 ;
        RECT 132.800 187.255 133.340 187.395 ;
        RECT 132.800 187.165 133.060 187.255 ;
        RECT 131.795 186.260 132.025 186.550 ;
        RECT 132.815 186.260 133.045 186.550 ;
        RECT 132.860 186.105 133.000 186.260 ;
        RECT 132.800 185.785 133.060 186.105 ;
        RECT 133.200 186.015 133.340 187.255 ;
        RECT 133.495 186.015 133.725 186.090 ;
        RECT 133.200 185.875 133.725 186.015 ;
        RECT 133.495 185.800 133.725 185.875 ;
        RECT 132.800 184.865 133.060 185.185 ;
        RECT 133.880 183.415 134.360 219.295 ;
        RECT 134.500 217.525 134.760 217.845 ;
        RECT 134.515 215.700 134.745 215.990 ;
        RECT 134.560 213.245 134.700 215.700 ;
        RECT 135.520 215.225 135.780 215.545 ;
        RECT 135.535 214.320 135.765 214.610 ;
        RECT 135.195 213.400 135.425 213.690 ;
        RECT 135.580 213.615 135.720 214.320 ;
        RECT 135.580 213.475 136.400 213.615 ;
        RECT 134.500 212.925 134.760 213.245 ;
        RECT 134.900 212.355 135.040 212.760 ;
        RECT 134.855 212.325 135.085 212.355 ;
        RECT 134.840 212.005 135.100 212.325 ;
        RECT 134.900 204.875 135.040 212.005 ;
        RECT 135.240 210.945 135.380 213.400 ;
        RECT 135.875 212.915 136.105 213.205 ;
        RECT 135.535 212.520 135.765 212.810 ;
        RECT 135.580 211.620 135.720 212.520 ;
        RECT 135.535 211.330 135.765 211.620 ;
        RECT 135.180 210.625 135.440 210.945 ;
        RECT 135.240 208.185 135.380 210.625 ;
        RECT 135.580 209.100 135.720 211.330 ;
        RECT 135.920 211.105 136.060 212.915 ;
        RECT 135.875 210.815 136.105 211.105 ;
        RECT 135.920 209.535 136.060 210.815 ;
        RECT 135.875 209.245 136.105 209.535 ;
        RECT 135.535 208.810 135.765 209.100 ;
        RECT 135.180 207.865 135.440 208.185 ;
        RECT 135.875 206.715 136.105 206.790 ;
        RECT 134.560 204.735 135.040 204.875 ;
        RECT 135.240 206.575 136.105 206.715 ;
        RECT 134.560 198.525 134.700 204.735 ;
        RECT 134.855 204.245 135.085 204.535 ;
        RECT 134.500 198.205 134.760 198.525 ;
        RECT 134.560 197.590 134.700 198.205 ;
        RECT 134.900 198.065 135.040 204.245 ;
        RECT 134.840 197.745 135.100 198.065 ;
        RECT 135.240 197.605 135.380 206.575 ;
        RECT 135.875 206.500 136.105 206.575 ;
        RECT 135.520 205.565 135.780 205.885 ;
        RECT 135.875 205.095 136.105 205.385 ;
        RECT 135.535 204.700 135.765 204.990 ;
        RECT 135.580 203.800 135.720 204.700 ;
        RECT 135.535 203.510 135.765 203.800 ;
        RECT 135.580 201.280 135.720 203.510 ;
        RECT 135.920 203.285 136.060 205.095 ;
        RECT 136.260 204.965 136.400 213.475 ;
        RECT 136.200 204.645 136.460 204.965 ;
        RECT 135.875 202.995 136.105 203.285 ;
        RECT 135.920 201.715 136.060 202.995 ;
        RECT 135.875 201.425 136.105 201.715 ;
        RECT 135.535 200.990 135.765 201.280 ;
        RECT 136.215 198.680 136.445 198.970 ;
        RECT 136.260 198.525 136.400 198.680 ;
        RECT 136.200 198.205 136.460 198.525 ;
        RECT 134.515 197.300 134.745 197.590 ;
        RECT 135.180 197.285 135.440 197.605 ;
        RECT 134.840 196.595 135.100 196.685 ;
        RECT 135.240 196.595 135.380 197.285 ;
        RECT 135.860 196.825 136.120 197.145 ;
        RECT 134.840 196.455 135.380 196.595 ;
        RECT 134.840 196.365 135.100 196.455 ;
        RECT 134.900 195.290 135.040 196.365 ;
        RECT 134.855 195.000 135.085 195.290 ;
        RECT 134.515 193.620 134.745 193.910 ;
        RECT 134.560 193.005 134.700 193.620 ;
        RECT 134.500 192.685 134.760 193.005 ;
        RECT 135.195 192.915 135.425 192.990 ;
        RECT 134.900 192.775 135.425 192.915 ;
        RECT 134.900 192.455 135.040 192.775 ;
        RECT 135.195 192.700 135.425 192.775 ;
        RECT 134.560 192.315 135.040 192.455 ;
        RECT 135.535 192.455 135.765 192.530 ;
        RECT 135.535 192.315 136.060 192.455 ;
        RECT 134.560 187.855 134.700 192.315 ;
        RECT 135.535 192.240 135.765 192.315 ;
        RECT 135.535 191.780 135.765 192.070 ;
        RECT 135.195 191.535 135.425 191.610 ;
        RECT 134.900 191.395 135.425 191.535 ;
        RECT 134.900 190.230 135.040 191.395 ;
        RECT 135.195 191.320 135.425 191.395 ;
        RECT 135.180 190.845 135.440 191.165 ;
        RECT 135.240 190.690 135.380 190.845 ;
        RECT 135.195 190.400 135.425 190.690 ;
        RECT 134.855 189.940 135.085 190.230 ;
        RECT 135.195 189.480 135.425 189.770 ;
        RECT 135.240 188.405 135.380 189.480 ;
        RECT 135.580 189.325 135.720 191.780 ;
        RECT 135.920 190.245 136.060 192.315 ;
        RECT 135.860 189.925 136.120 190.245 ;
        RECT 135.520 189.005 135.780 189.325 ;
        RECT 135.180 188.085 135.440 188.405 ;
        RECT 135.180 187.855 135.440 187.945 ;
        RECT 134.560 187.715 135.440 187.855 ;
        RECT 135.180 187.625 135.440 187.715 ;
        RECT 135.180 186.245 135.440 186.565 ;
        RECT 135.180 185.785 135.440 186.105 ;
        RECT 135.240 185.630 135.380 185.785 ;
        RECT 135.920 185.645 136.060 189.925 ;
        RECT 136.215 188.560 136.445 188.850 ;
        RECT 136.260 187.025 136.400 188.560 ;
        RECT 136.200 186.705 136.460 187.025 ;
        RECT 135.195 185.340 135.425 185.630 ;
        RECT 135.860 185.325 136.120 185.645 ;
        RECT 136.600 183.415 137.080 219.295 ;
        RECT 138.920 217.985 139.180 218.305 ;
        RECT 138.980 217.370 139.120 217.985 ;
        RECT 138.935 217.080 139.165 217.370 ;
        RECT 138.255 216.160 138.485 216.450 ;
        RECT 137.560 215.225 137.820 215.545 ;
        RECT 137.620 213.615 137.760 215.225 ;
        RECT 137.915 213.615 138.145 213.690 ;
        RECT 137.620 213.475 138.145 213.615 ;
        RECT 137.235 200.980 137.465 201.270 ;
        RECT 137.280 200.825 137.420 200.980 ;
        RECT 137.220 200.505 137.480 200.825 ;
        RECT 137.620 195.765 137.760 213.475 ;
        RECT 137.915 213.400 138.145 213.475 ;
        RECT 137.915 212.480 138.145 212.770 ;
        RECT 137.960 212.325 138.100 212.480 ;
        RECT 137.900 212.005 138.160 212.325 ;
        RECT 138.300 210.945 138.440 216.160 ;
        RECT 138.920 215.685 139.180 216.005 ;
        RECT 138.935 213.860 139.165 214.150 ;
        RECT 138.240 210.625 138.500 210.945 ;
        RECT 138.980 210.485 139.120 213.860 ;
        RECT 138.920 210.165 139.180 210.485 ;
        RECT 138.920 207.865 139.180 208.185 ;
        RECT 138.980 205.885 139.120 207.865 ;
        RECT 138.920 205.565 139.180 205.885 ;
        RECT 138.920 204.645 139.180 204.965 ;
        RECT 138.255 201.440 138.485 201.730 ;
        RECT 138.300 201.285 138.440 201.440 ;
        RECT 138.980 201.285 139.120 204.645 ;
        RECT 138.240 200.965 138.500 201.285 ;
        RECT 138.920 200.965 139.180 201.285 ;
        RECT 137.915 197.760 138.145 198.050 ;
        RECT 137.960 197.605 138.100 197.760 ;
        RECT 137.900 197.285 138.160 197.605 ;
        RECT 138.580 195.905 138.840 196.225 ;
        RECT 137.560 195.445 137.820 195.765 ;
        RECT 137.915 195.000 138.145 195.290 ;
        RECT 137.235 194.755 137.465 194.830 ;
        RECT 137.235 194.615 137.760 194.755 ;
        RECT 137.235 194.540 137.465 194.615 ;
        RECT 137.220 193.605 137.480 193.925 ;
        RECT 137.620 191.165 137.760 194.615 ;
        RECT 137.960 191.995 138.100 195.000 ;
        RECT 138.255 194.755 138.485 194.830 ;
        RECT 138.255 194.615 139.120 194.755 ;
        RECT 138.255 194.540 138.485 194.615 ;
        RECT 138.595 192.700 138.825 192.990 ;
        RECT 138.240 191.995 138.500 192.085 ;
        RECT 137.960 191.855 138.500 191.995 ;
        RECT 138.240 191.765 138.500 191.855 ;
        RECT 138.640 191.625 138.780 192.700 ;
        RECT 138.580 191.305 138.840 191.625 ;
        RECT 137.560 190.845 137.820 191.165 ;
        RECT 138.580 190.845 138.840 191.165 ;
        RECT 138.255 190.615 138.485 190.690 ;
        RECT 137.960 190.475 138.485 190.615 ;
        RECT 137.960 189.310 138.100 190.475 ;
        RECT 138.255 190.400 138.485 190.475 ;
        RECT 138.255 189.695 138.485 189.770 ;
        RECT 138.640 189.695 138.780 190.845 ;
        RECT 138.255 189.555 138.780 189.695 ;
        RECT 138.255 189.480 138.485 189.555 ;
        RECT 137.915 189.020 138.145 189.310 ;
        RECT 138.240 188.085 138.500 188.405 ;
        RECT 138.240 186.705 138.500 187.025 ;
        RECT 138.255 185.800 138.485 186.090 ;
        RECT 138.640 186.015 138.780 189.555 ;
        RECT 138.980 188.405 139.120 194.615 ;
        RECT 138.920 188.085 139.180 188.405 ;
        RECT 138.920 186.015 139.180 186.105 ;
        RECT 138.640 185.875 139.180 186.015 ;
        RECT 138.300 185.645 138.440 185.800 ;
        RECT 138.920 185.785 139.180 185.875 ;
        RECT 138.240 185.325 138.500 185.645 ;
        RECT 139.320 183.415 139.800 219.295 ;
        RECT 140.635 217.540 140.865 217.830 ;
        RECT 140.295 216.205 140.525 216.495 ;
        RECT 140.340 216.005 140.480 216.205 ;
        RECT 140.280 215.685 140.540 216.005 ;
        RECT 139.940 210.855 140.200 210.945 ;
        RECT 139.940 210.715 140.480 210.855 ;
        RECT 139.940 210.625 140.200 210.715 ;
        RECT 139.940 210.165 140.200 210.485 ;
        RECT 140.340 207.635 140.480 210.715 ;
        RECT 140.680 208.185 140.820 217.540 ;
        RECT 141.315 217.055 141.545 217.345 ;
        RECT 140.975 216.660 141.205 216.950 ;
        RECT 141.020 215.760 141.160 216.660 ;
        RECT 140.975 215.470 141.205 215.760 ;
        RECT 141.020 213.240 141.160 215.470 ;
        RECT 141.360 215.245 141.500 217.055 ;
        RECT 141.315 214.955 141.545 215.245 ;
        RECT 141.360 213.675 141.500 214.955 ;
        RECT 141.315 213.385 141.545 213.675 ;
        RECT 140.975 212.950 141.205 213.240 ;
        RECT 140.620 207.865 140.880 208.185 ;
        RECT 140.635 207.635 140.865 207.710 ;
        RECT 140.340 207.495 140.865 207.635 ;
        RECT 140.635 207.420 140.865 207.495 ;
        RECT 141.640 205.565 141.900 205.885 ;
        RECT 140.635 203.740 140.865 204.030 ;
        RECT 140.295 203.280 140.525 203.570 ;
        RECT 139.940 201.425 140.200 201.745 ;
        RECT 140.000 199.430 140.140 201.425 ;
        RECT 139.955 199.140 140.185 199.430 ;
        RECT 140.340 195.765 140.480 203.280 ;
        RECT 140.680 201.745 140.820 203.740 ;
        RECT 140.975 202.575 141.205 202.650 ;
        RECT 140.975 202.435 141.500 202.575 ;
        RECT 140.975 202.360 141.205 202.435 ;
        RECT 140.620 201.425 140.880 201.745 ;
        RECT 140.620 200.965 140.880 201.285 ;
        RECT 140.620 200.045 140.880 200.365 ;
        RECT 140.680 198.525 140.820 200.045 ;
        RECT 140.620 198.205 140.880 198.525 ;
        RECT 140.620 197.745 140.880 198.065 ;
        RECT 140.680 197.145 140.820 197.745 ;
        RECT 140.960 197.285 141.220 197.605 ;
        RECT 141.360 197.515 141.500 202.435 ;
        RECT 141.640 200.505 141.900 200.825 ;
        RECT 141.700 198.510 141.840 200.505 ;
        RECT 141.655 198.220 141.885 198.510 ;
        RECT 141.360 197.375 141.840 197.515 ;
        RECT 140.620 196.825 140.880 197.145 ;
        RECT 141.315 196.815 141.545 197.105 ;
        RECT 140.975 196.420 141.205 196.710 ;
        RECT 140.635 195.965 140.865 196.255 ;
        RECT 140.280 195.445 140.540 195.765 ;
        RECT 140.680 194.845 140.820 195.965 ;
        RECT 141.020 195.520 141.160 196.420 ;
        RECT 140.975 195.230 141.205 195.520 ;
        RECT 140.620 194.525 140.880 194.845 ;
        RECT 141.020 193.000 141.160 195.230 ;
        RECT 141.360 195.005 141.500 196.815 ;
        RECT 141.700 195.765 141.840 197.375 ;
        RECT 141.640 195.445 141.900 195.765 ;
        RECT 141.315 194.715 141.545 195.005 ;
        RECT 141.360 193.435 141.500 194.715 ;
        RECT 141.315 193.145 141.545 193.435 ;
        RECT 140.975 192.710 141.205 193.000 ;
        RECT 141.700 192.455 141.840 195.445 ;
        RECT 140.680 192.315 141.840 192.455 ;
        RECT 140.680 189.770 140.820 192.315 ;
        RECT 141.640 190.385 141.900 190.705 ;
        RECT 140.635 189.480 140.865 189.770 ;
        RECT 140.620 188.545 140.880 188.865 ;
        RECT 141.640 187.625 141.900 187.945 ;
        RECT 140.620 187.165 140.880 187.485 ;
        RECT 139.940 186.245 140.200 186.565 ;
        RECT 139.940 185.785 140.200 186.105 ;
        RECT 140.620 184.865 140.880 185.185 ;
        RECT 142.040 183.415 142.520 219.295 ;
        RECT 144.360 213.385 144.620 213.705 ;
        RECT 143.355 211.090 143.585 211.380 ;
        RECT 143.015 210.655 143.245 210.945 ;
        RECT 143.060 209.375 143.200 210.655 ;
        RECT 143.015 209.085 143.245 209.375 ;
        RECT 142.660 207.865 142.920 208.185 ;
        RECT 142.720 206.255 142.860 207.865 ;
        RECT 143.060 207.275 143.200 209.085 ;
        RECT 143.400 208.860 143.540 211.090 ;
        RECT 143.355 208.570 143.585 208.860 ;
        RECT 144.360 208.785 144.620 209.105 ;
        RECT 143.400 207.670 143.540 208.570 ;
        RECT 143.695 207.780 143.925 208.070 ;
        RECT 143.355 207.380 143.585 207.670 ;
        RECT 143.015 206.985 143.245 207.275 ;
        RECT 143.355 206.500 143.585 206.790 ;
        RECT 143.400 206.330 143.540 206.500 ;
        RECT 143.355 206.255 143.585 206.330 ;
        RECT 142.720 206.115 143.585 206.255 ;
        RECT 142.720 197.605 142.860 206.115 ;
        RECT 143.355 206.040 143.585 206.115 ;
        RECT 143.740 205.885 143.880 207.780 ;
        RECT 144.020 206.485 144.280 206.805 ;
        RECT 143.015 205.555 143.245 205.845 ;
        RECT 143.680 205.565 143.940 205.885 ;
        RECT 143.060 203.745 143.200 205.555 ;
        RECT 143.355 205.160 143.585 205.450 ;
        RECT 143.400 204.260 143.540 205.160 ;
        RECT 144.080 205.105 144.220 206.485 ;
        RECT 144.035 204.815 144.265 205.105 ;
        RECT 143.355 203.970 143.585 204.260 ;
        RECT 143.015 203.455 143.245 203.745 ;
        RECT 143.060 202.175 143.200 203.455 ;
        RECT 143.015 201.885 143.245 202.175 ;
        RECT 143.400 201.740 143.540 203.970 ;
        RECT 144.420 203.955 144.560 208.785 ;
        RECT 144.080 203.815 144.560 203.955 ;
        RECT 143.355 201.450 143.585 201.740 ;
        RECT 143.000 200.965 143.260 201.285 ;
        RECT 142.660 197.285 142.920 197.605 ;
        RECT 143.060 195.750 143.200 200.965 ;
        RECT 143.340 200.045 143.600 200.365 ;
        RECT 143.400 196.595 143.540 200.045 ;
        RECT 144.080 198.970 144.220 203.815 ;
        RECT 144.375 199.140 144.605 199.430 ;
        RECT 144.035 198.680 144.265 198.970 ;
        RECT 144.420 198.525 144.560 199.140 ;
        RECT 144.360 198.205 144.620 198.525 ;
        RECT 144.020 197.745 144.280 198.065 ;
        RECT 143.680 196.825 143.940 197.145 ;
        RECT 143.695 196.595 143.925 196.670 ;
        RECT 143.400 196.455 143.925 196.595 ;
        RECT 143.695 196.380 143.925 196.455 ;
        RECT 143.340 195.905 143.600 196.225 ;
        RECT 143.015 195.460 143.245 195.750 ;
        RECT 142.660 194.525 142.920 194.845 ;
        RECT 142.720 192.990 142.860 194.525 ;
        RECT 143.015 194.080 143.245 194.370 ;
        RECT 142.675 192.700 142.905 192.990 ;
        RECT 143.060 191.610 143.200 194.080 ;
        RECT 143.400 193.835 143.540 195.905 ;
        RECT 143.680 195.445 143.940 195.765 ;
        RECT 143.740 194.830 143.880 195.445 ;
        RECT 143.695 194.540 143.925 194.830 ;
        RECT 143.680 193.835 143.940 193.925 ;
        RECT 143.400 193.695 143.940 193.835 ;
        RECT 143.680 193.605 143.940 193.695 ;
        RECT 143.740 192.070 143.880 193.605 ;
        RECT 143.695 191.780 143.925 192.070 ;
        RECT 143.015 191.320 143.245 191.610 ;
        RECT 143.680 190.845 143.940 191.165 ;
        RECT 143.000 190.385 143.260 190.705 ;
        RECT 143.695 190.400 143.925 190.690 ;
        RECT 143.060 189.695 143.200 190.385 ;
        RECT 143.355 189.695 143.585 189.770 ;
        RECT 143.060 189.555 143.585 189.695 ;
        RECT 143.355 189.480 143.585 189.555 ;
        RECT 142.660 188.545 142.920 188.865 ;
        RECT 142.720 186.550 142.860 188.545 ;
        RECT 143.740 187.945 143.880 190.400 ;
        RECT 143.680 187.625 143.940 187.945 ;
        RECT 143.000 187.165 143.260 187.485 ;
        RECT 142.675 186.260 142.905 186.550 ;
        RECT 143.060 186.090 143.200 187.165 ;
        RECT 143.015 185.800 143.245 186.090 ;
        RECT 143.680 184.865 143.940 185.185 ;
        RECT 144.760 183.415 145.240 219.295 ;
        RECT 146.060 213.385 146.320 213.705 ;
        RECT 146.120 211.390 146.260 213.385 ;
        RECT 146.075 211.315 146.305 211.390 ;
        RECT 146.075 211.175 146.600 211.315 ;
        RECT 146.075 211.100 146.305 211.175 ;
        RECT 146.060 208.785 146.320 209.105 ;
        RECT 146.060 208.325 146.320 208.645 ;
        RECT 146.075 207.420 146.305 207.710 ;
        RECT 145.380 206.485 145.640 206.805 ;
        RECT 145.380 201.425 145.640 201.745 ;
        RECT 146.120 199.355 146.260 207.420 ;
        RECT 146.460 204.950 146.600 211.175 ;
        RECT 147.095 210.180 147.325 210.470 ;
        RECT 146.755 207.880 146.985 208.170 ;
        RECT 146.415 204.660 146.645 204.950 ;
        RECT 146.800 200.825 146.940 207.880 ;
        RECT 147.140 205.425 147.280 210.180 ;
        RECT 147.080 205.105 147.340 205.425 ;
        RECT 146.740 200.505 147.000 200.825 ;
        RECT 147.095 199.600 147.325 199.890 ;
        RECT 146.120 199.215 146.940 199.355 ;
        RECT 146.075 198.680 146.305 198.970 ;
        RECT 146.120 198.525 146.260 198.680 ;
        RECT 146.060 198.205 146.320 198.525 ;
        RECT 145.380 197.745 145.640 198.065 ;
        RECT 145.440 195.290 145.580 197.745 ;
        RECT 146.060 195.445 146.320 195.765 ;
        RECT 145.395 195.000 145.625 195.290 ;
        RECT 146.120 194.830 146.260 195.445 ;
        RECT 146.075 194.540 146.305 194.830 ;
        RECT 146.800 193.925 146.940 199.215 ;
        RECT 147.140 198.985 147.280 199.600 ;
        RECT 147.080 198.665 147.340 198.985 ;
        RECT 146.740 193.605 147.000 193.925 ;
        RECT 147.080 192.225 147.340 192.545 ;
        RECT 145.380 191.765 145.640 192.085 ;
        RECT 145.440 188.850 145.580 191.765 ;
        RECT 147.140 191.610 147.280 192.225 ;
        RECT 147.095 191.320 147.325 191.610 ;
        RECT 146.060 190.385 146.320 190.705 ;
        RECT 145.395 188.560 145.625 188.850 ;
        RECT 145.380 188.085 145.640 188.405 ;
        RECT 145.440 187.470 145.580 188.085 ;
        RECT 146.060 187.625 146.320 187.945 ;
        RECT 145.395 187.180 145.625 187.470 ;
        RECT 146.060 186.245 146.320 186.565 ;
        RECT 145.395 185.800 145.625 186.090 ;
        RECT 145.440 185.645 145.580 185.800 ;
        RECT 145.380 185.325 145.640 185.645 ;
        RECT 146.060 184.865 146.320 185.185 ;
        RECT 147.480 183.415 147.960 219.295 ;
        RECT 148.200 201.290 148.340 219.570 ;
        RECT 148.110 200.960 148.440 201.290 ;
        RECT 148.720 198.955 148.860 220.050 ;
        RECT 148.630 198.695 148.950 198.955 ;
        RECT 149.210 198.060 149.350 220.770 ;
        RECT 149.770 205.430 149.910 221.830 ;
        RECT 149.680 205.100 150.000 205.430 ;
        RECT 148.670 197.920 149.350 198.060 ;
        RECT 148.670 192.550 148.810 197.920 ;
        RECT 148.570 192.220 148.900 192.550 ;
        RECT 101.005 178.120 102.595 182.410 ;
        RECT 100.100 178.100 140.370 178.120 ;
        RECT 100.100 178.080 140.860 178.100 ;
        RECT 99.990 177.050 140.860 178.080 ;
        RECT 99.990 176.770 100.770 177.050 ;
        RECT 99.990 175.260 100.880 176.770 ;
        RECT 106.550 176.380 107.800 176.820 ;
        RECT 117.640 176.640 118.600 176.800 ;
        RECT 120.030 176.750 120.810 177.050 ;
        RECT 140.080 176.800 140.860 177.050 ;
        RECT 104.490 176.370 109.730 176.380 ;
        RECT 101.540 176.270 116.840 176.370 ;
        RECT 101.540 176.260 116.875 176.270 ;
        RECT 101.500 176.140 116.875 176.260 ;
        RECT 101.500 176.030 105.500 176.140 ;
        RECT 106.550 176.060 108.290 176.140 ;
        RECT 108.870 176.060 116.875 176.140 ;
        RECT 106.550 175.980 107.800 176.060 ;
        RECT 108.875 176.040 116.875 176.060 ;
        RECT 100.050 174.670 100.880 175.260 ;
        RECT 101.110 175.730 101.340 175.980 ;
        RECT 105.660 175.840 105.890 175.980 ;
        RECT 108.440 175.840 108.670 175.990 ;
        RECT 105.660 175.730 108.670 175.840 ;
        RECT 117.080 175.730 117.310 175.990 ;
        RECT 101.110 175.290 117.310 175.730 ;
        RECT 101.110 175.020 101.340 175.290 ;
        RECT 105.660 175.260 117.310 175.290 ;
        RECT 105.660 175.170 108.670 175.260 ;
        RECT 105.660 175.020 105.890 175.170 ;
        RECT 108.440 175.030 108.670 175.170 ;
        RECT 117.080 175.030 117.310 175.260 ;
        RECT 101.500 174.740 105.500 174.970 ;
        RECT 108.875 174.760 116.875 174.980 ;
        RECT 117.640 174.760 118.880 176.640 ;
        RECT 108.875 174.750 118.880 174.760 ;
        RECT 101.500 174.670 105.490 174.740 ;
        RECT 100.050 174.560 105.490 174.670 ;
        RECT 108.930 174.620 118.880 174.750 ;
        RECT 119.930 175.260 120.810 176.750 ;
        RECT 126.430 176.330 127.680 176.770 ;
        RECT 137.520 176.620 138.480 176.750 ;
        RECT 124.370 176.320 129.610 176.330 ;
        RECT 121.420 176.220 136.720 176.320 ;
        RECT 121.420 176.210 136.755 176.220 ;
        RECT 121.380 176.090 136.755 176.210 ;
        RECT 121.380 175.980 125.380 176.090 ;
        RECT 126.430 176.010 128.170 176.090 ;
        RECT 128.750 176.010 136.755 176.090 ;
        RECT 126.430 175.930 127.680 176.010 ;
        RECT 128.755 175.990 136.755 176.010 ;
        RECT 120.990 175.680 121.220 175.930 ;
        RECT 125.540 175.790 125.770 175.930 ;
        RECT 128.320 175.790 128.550 175.940 ;
        RECT 125.540 175.680 128.550 175.790 ;
        RECT 136.960 175.680 137.190 175.940 ;
        RECT 119.930 174.620 120.760 175.260 ;
        RECT 120.990 175.240 137.190 175.680 ;
        RECT 120.990 174.970 121.220 175.240 ;
        RECT 125.540 175.210 137.190 175.240 ;
        RECT 125.540 175.120 128.550 175.210 ;
        RECT 125.540 174.970 125.770 175.120 ;
        RECT 128.320 174.980 128.550 175.120 ;
        RECT 136.960 174.980 137.190 175.210 ;
        RECT 121.380 174.690 125.380 174.920 ;
        RECT 128.755 174.710 136.755 174.930 ;
        RECT 137.520 174.710 138.700 176.620 ;
        RECT 128.755 174.700 138.700 174.710 ;
        RECT 121.380 174.620 125.370 174.690 ;
        RECT 108.930 174.590 118.600 174.620 ;
        RECT 100.050 174.470 103.180 174.560 ;
        RECT 116.670 174.540 118.600 174.590 ;
        RECT 12.100 173.620 89.840 174.100 ;
        RECT 45.290 173.420 45.610 173.480 ;
        RECT 46.225 173.420 46.515 173.465 ;
        RECT 45.290 173.280 46.515 173.420 ;
        RECT 45.290 173.220 45.610 173.280 ;
        RECT 46.225 173.235 46.515 173.280 ;
        RECT 65.085 173.420 65.375 173.465 ;
        RECT 71.050 173.420 71.370 173.480 ;
        RECT 65.085 173.280 71.370 173.420 ;
        RECT 65.085 173.235 65.375 173.280 ;
        RECT 71.050 173.220 71.370 173.280 ;
        RECT 71.510 173.420 71.830 173.480 ;
        RECT 75.205 173.420 75.495 173.465 ;
        RECT 80.710 173.420 81.030 173.480 ;
        RECT 71.510 173.280 74.960 173.420 ;
        RECT 71.510 173.220 71.830 173.280 ;
        RECT 62.325 173.080 62.615 173.125 ;
        RECT 74.270 173.080 74.590 173.140 ;
        RECT 62.325 172.940 74.590 173.080 ;
        RECT 74.820 173.080 74.960 173.280 ;
        RECT 75.205 173.280 81.030 173.420 ;
        RECT 75.205 173.235 75.495 173.280 ;
        RECT 80.710 173.220 81.030 173.280 ;
        RECT 83.010 173.420 83.330 173.480 ;
        RECT 88.990 173.420 89.310 173.480 ;
        RECT 83.010 173.280 89.310 173.420 ;
        RECT 83.010 173.220 83.330 173.280 ;
        RECT 88.990 173.220 89.310 173.280 ;
        RECT 74.820 172.940 84.620 173.080 ;
        RECT 62.325 172.895 62.615 172.940 ;
        RECT 74.270 172.880 74.590 172.940 ;
        RECT 83.930 172.740 84.250 172.800 ;
        RECT 67.000 172.600 84.250 172.740 ;
        RECT 47.130 172.200 47.450 172.460 ;
        RECT 59.550 172.200 59.870 172.460 ;
        RECT 60.930 172.400 61.250 172.460 ;
        RECT 61.405 172.400 61.695 172.445 ;
        RECT 60.930 172.260 61.695 172.400 ;
        RECT 60.930 172.200 61.250 172.260 ;
        RECT 61.405 172.215 61.695 172.260 ;
        RECT 63.230 172.200 63.550 172.460 ;
        RECT 64.150 172.200 64.470 172.460 ;
        RECT 58.630 171.520 58.950 171.780 ;
        RECT 60.470 171.520 60.790 171.780 ;
        RECT 66.465 171.720 66.755 171.765 ;
        RECT 67.000 171.720 67.140 172.600 ;
        RECT 83.930 172.540 84.250 172.600 ;
        RECT 67.385 172.215 67.675 172.445 ;
        RECT 70.145 172.400 70.435 172.445 ;
        RECT 70.145 172.260 75.880 172.400 ;
        RECT 70.145 172.215 70.435 172.260 ;
        RECT 67.460 172.060 67.600 172.215 ;
        RECT 68.765 172.060 69.055 172.105 ;
        RECT 69.210 172.060 69.530 172.120 ;
        RECT 67.460 171.920 68.520 172.060 ;
        RECT 66.465 171.580 67.140 171.720 ;
        RECT 66.465 171.535 66.755 171.580 ;
        RECT 67.830 171.520 68.150 171.780 ;
        RECT 68.380 171.720 68.520 171.920 ;
        RECT 68.765 171.920 69.530 172.060 ;
        RECT 68.765 171.875 69.055 171.920 ;
        RECT 69.210 171.860 69.530 171.920 ;
        RECT 69.685 172.060 69.975 172.105 ;
        RECT 70.590 172.060 70.910 172.120 ;
        RECT 69.685 171.920 70.910 172.060 ;
        RECT 69.685 171.875 69.975 171.920 ;
        RECT 70.590 171.860 70.910 171.920 ;
        RECT 71.065 172.060 71.355 172.105 ;
        RECT 71.510 172.060 71.830 172.120 ;
        RECT 71.065 171.920 71.830 172.060 ;
        RECT 71.065 171.875 71.355 171.920 ;
        RECT 71.140 171.720 71.280 171.875 ;
        RECT 71.510 171.860 71.830 171.920 ;
        RECT 71.985 172.060 72.275 172.105 ;
        RECT 71.985 171.920 73.120 172.060 ;
        RECT 71.985 171.875 72.275 171.920 ;
        RECT 68.380 171.580 71.280 171.720 ;
        RECT 72.430 171.520 72.750 171.780 ;
        RECT 72.980 171.720 73.120 171.920 ;
        RECT 73.350 171.860 73.670 172.120 ;
        RECT 73.810 172.060 74.130 172.120 ;
        RECT 74.285 172.060 74.575 172.105 ;
        RECT 73.810 171.920 74.575 172.060 ;
        RECT 75.740 172.060 75.880 172.260 ;
        RECT 76.110 172.200 76.430 172.460 ;
        RECT 81.170 172.400 81.490 172.460 ;
        RECT 76.660 172.260 81.490 172.400 ;
        RECT 76.660 172.060 76.800 172.260 ;
        RECT 81.170 172.200 81.490 172.260 ;
        RECT 81.645 172.400 81.935 172.445 ;
        RECT 83.010 172.400 83.330 172.460 ;
        RECT 81.645 172.260 83.330 172.400 ;
        RECT 81.645 172.215 81.935 172.260 ;
        RECT 83.010 172.200 83.330 172.260 ;
        RECT 83.470 172.400 83.790 172.460 ;
        RECT 84.480 172.445 84.620 172.940 ;
        RECT 84.405 172.400 84.695 172.445 ;
        RECT 83.470 172.260 84.695 172.400 ;
        RECT 83.470 172.200 83.790 172.260 ;
        RECT 84.405 172.215 84.695 172.260 ;
        RECT 86.245 172.400 86.535 172.445 ;
        RECT 87.150 172.400 87.470 172.460 ;
        RECT 86.245 172.260 87.470 172.400 ;
        RECT 86.245 172.215 86.535 172.260 ;
        RECT 87.150 172.200 87.470 172.260 ;
        RECT 75.740 171.920 76.800 172.060 ;
        RECT 77.045 172.060 77.335 172.105 ;
        RECT 77.490 172.060 77.810 172.120 ;
        RECT 77.045 171.920 77.810 172.060 ;
        RECT 73.810 171.860 74.130 171.920 ;
        RECT 74.285 171.875 74.575 171.920 ;
        RECT 77.045 171.875 77.335 171.920 ;
        RECT 77.120 171.720 77.260 171.875 ;
        RECT 77.490 171.860 77.810 171.920 ;
        RECT 77.950 171.860 78.270 172.120 ;
        RECT 78.410 172.060 78.730 172.120 ;
        RECT 79.345 172.060 79.635 172.105 ;
        RECT 78.410 171.920 79.635 172.060 ;
        RECT 78.410 171.860 78.730 171.920 ;
        RECT 79.345 171.875 79.635 171.920 ;
        RECT 79.790 172.060 80.110 172.120 ;
        RECT 80.265 172.060 80.555 172.105 ;
        RECT 79.790 171.920 80.555 172.060 ;
        RECT 79.790 171.860 80.110 171.920 ;
        RECT 80.265 171.875 80.555 171.920 ;
        RECT 82.565 172.060 82.855 172.105 ;
        RECT 84.850 172.060 85.170 172.120 ;
        RECT 82.565 171.920 85.170 172.060 ;
        RECT 82.565 171.875 82.855 171.920 ;
        RECT 84.850 171.860 85.170 171.920 ;
        RECT 85.310 171.860 85.630 172.120 ;
        RECT 85.770 172.060 86.090 172.120 ;
        RECT 87.610 172.060 87.930 172.120 ;
        RECT 85.770 171.920 87.930 172.060 ;
        RECT 85.770 171.860 86.090 171.920 ;
        RECT 87.610 171.860 87.930 171.920 ;
        RECT 72.980 171.580 77.260 171.720 ;
        RECT 78.870 171.520 79.190 171.780 ;
        RECT 80.710 171.720 81.030 171.780 ;
        RECT 81.185 171.720 81.475 171.765 ;
        RECT 80.710 171.580 81.475 171.720 ;
        RECT 80.710 171.520 81.030 171.580 ;
        RECT 81.185 171.535 81.475 171.580 ;
        RECT 83.010 171.720 83.330 171.780 ;
        RECT 83.485 171.720 83.775 171.765 ;
        RECT 83.010 171.580 83.775 171.720 ;
        RECT 83.010 171.520 83.330 171.580 ;
        RECT 83.485 171.535 83.775 171.580 ;
        RECT 83.930 171.720 84.250 171.780 ;
        RECT 87.165 171.720 87.455 171.765 ;
        RECT 83.930 171.580 87.455 171.720 ;
        RECT 83.930 171.520 84.250 171.580 ;
        RECT 87.165 171.535 87.455 171.580 ;
        RECT 12.100 170.900 89.840 171.380 ;
        RECT 100.050 171.200 100.880 174.470 ;
        RECT 104.530 174.010 109.780 174.020 ;
        RECT 104.530 173.900 116.840 174.010 ;
        RECT 101.560 173.840 116.840 173.900 ;
        RECT 101.560 173.830 116.875 173.840 ;
        RECT 101.500 173.700 116.875 173.830 ;
        RECT 101.500 173.690 106.660 173.700 ;
        RECT 101.500 173.600 105.500 173.690 ;
        RECT 108.875 173.610 116.875 173.700 ;
        RECT 108.960 173.600 116.850 173.610 ;
        RECT 101.110 173.240 101.340 173.550 ;
        RECT 101.560 173.240 105.460 173.600 ;
        RECT 105.660 173.240 105.890 173.550 ;
        RECT 101.110 171.900 105.890 173.240 ;
        RECT 101.110 171.590 101.340 171.900 ;
        RECT 105.660 171.590 105.890 171.900 ;
        RECT 108.440 173.020 108.670 173.560 ;
        RECT 109.480 173.020 110.490 173.050 ;
        RECT 117.080 173.020 117.310 173.560 ;
        RECT 108.440 172.120 117.310 173.020 ;
        RECT 108.440 171.600 108.670 172.120 ;
        RECT 109.480 172.050 110.490 172.120 ;
        RECT 117.080 171.600 117.310 172.120 ;
        RECT 101.500 171.310 105.500 171.540 ;
        RECT 108.875 171.320 116.875 171.550 ;
        RECT 100.050 171.160 101.180 171.200 ;
        RECT 100.050 171.080 101.420 171.160 ;
        RECT 101.790 171.090 105.450 171.310 ;
        RECT 101.790 171.080 103.230 171.090 ;
        RECT 100.050 171.040 103.230 171.080 ;
        RECT 100.050 170.950 102.740 171.040 ;
        RECT 108.940 171.030 116.830 171.320 ;
        RECT 100.050 170.890 102.070 170.950 ;
        RECT 100.050 170.840 101.820 170.890 ;
        RECT 63.230 170.700 63.550 170.760 ;
        RECT 68.765 170.700 69.055 170.745 ;
        RECT 73.350 170.700 73.670 170.760 ;
        RECT 63.230 170.560 73.670 170.700 ;
        RECT 63.230 170.500 63.550 170.560 ;
        RECT 68.765 170.515 69.055 170.560 ;
        RECT 73.350 170.500 73.670 170.560 ;
        RECT 73.810 170.700 74.130 170.760 ;
        RECT 78.410 170.700 78.730 170.760 ;
        RECT 73.810 170.560 78.730 170.700 ;
        RECT 73.810 170.500 74.130 170.560 ;
        RECT 78.410 170.500 78.730 170.560 ;
        RECT 78.870 170.500 79.190 170.760 ;
        RECT 80.340 170.560 84.160 170.700 ;
        RECT 60.470 170.160 60.790 170.420 ;
        RECT 76.570 170.360 76.890 170.420 ;
        RECT 78.960 170.360 79.100 170.500 ;
        RECT 76.570 170.220 78.640 170.360 ;
        RECT 78.960 170.220 79.560 170.360 ;
        RECT 76.570 170.160 76.890 170.220 ;
        RECT 41.165 169.835 41.455 170.065 ;
        RECT 41.240 169.680 41.380 169.835 ;
        RECT 42.530 169.820 42.850 170.080 ;
        RECT 43.450 169.820 43.770 170.080 ;
        RECT 43.910 170.020 44.230 170.080 ;
        RECT 51.285 170.020 51.575 170.065 ;
        RECT 43.910 169.880 51.575 170.020 ;
        RECT 43.910 169.820 44.230 169.880 ;
        RECT 51.285 169.835 51.575 169.880 ;
        RECT 52.190 169.820 52.510 170.080 ;
        RECT 59.565 170.020 59.855 170.065 ;
        RECT 60.560 170.020 60.700 170.160 ;
        RECT 74.270 170.065 74.590 170.080 ;
        RECT 59.565 169.880 70.820 170.020 ;
        RECT 59.565 169.835 59.855 169.880 ;
        RECT 44.830 169.680 45.150 169.740 ;
        RECT 41.240 169.540 45.150 169.680 ;
        RECT 44.830 169.480 45.150 169.540 ;
        RECT 60.470 169.480 60.790 169.740 ;
        RECT 61.480 169.540 66.680 169.680 ;
        RECT 41.610 169.140 41.930 169.400 ;
        RECT 42.070 169.140 42.390 169.400 ;
        RECT 58.645 169.340 58.935 169.385 ;
        RECT 61.480 169.340 61.620 169.540 ;
        RECT 58.645 169.200 61.620 169.340 ;
        RECT 61.850 169.340 62.170 169.400 ;
        RECT 64.165 169.340 64.455 169.385 ;
        RECT 61.850 169.200 64.455 169.340 ;
        RECT 66.540 169.340 66.680 169.540 ;
        RECT 66.910 169.480 67.230 169.740 ;
        RECT 69.670 169.340 69.990 169.400 ;
        RECT 66.540 169.200 69.990 169.340 ;
        RECT 58.645 169.155 58.935 169.200 ;
        RECT 61.850 169.140 62.170 169.200 ;
        RECT 64.165 169.155 64.455 169.200 ;
        RECT 69.670 169.140 69.990 169.200 ;
        RECT 40.230 168.800 40.550 169.060 ;
        RECT 48.510 169.000 48.830 169.060 ;
        RECT 51.745 169.000 52.035 169.045 ;
        RECT 48.510 168.860 52.035 169.000 ;
        RECT 48.510 168.800 48.830 168.860 ;
        RECT 51.745 168.815 52.035 168.860 ;
        RECT 63.230 168.800 63.550 169.060 ;
        RECT 70.680 169.000 70.820 169.880 ;
        RECT 74.270 169.835 74.620 170.065 ;
        RECT 75.190 170.020 75.510 170.080 ;
        RECT 78.500 170.065 78.640 170.220 ;
        RECT 75.190 169.880 76.800 170.020 ;
        RECT 74.270 169.820 74.590 169.835 ;
        RECT 75.190 169.820 75.510 169.880 ;
        RECT 71.075 169.680 71.365 169.725 ;
        RECT 73.595 169.680 73.885 169.725 ;
        RECT 74.785 169.680 75.075 169.725 ;
        RECT 71.075 169.540 75.075 169.680 ;
        RECT 71.075 169.495 71.365 169.540 ;
        RECT 73.595 169.495 73.885 169.540 ;
        RECT 74.785 169.495 75.075 169.540 ;
        RECT 75.665 169.680 75.955 169.725 ;
        RECT 76.110 169.680 76.430 169.740 ;
        RECT 75.665 169.540 76.430 169.680 ;
        RECT 76.660 169.680 76.800 169.880 ;
        RECT 78.425 169.835 78.715 170.065 ;
        RECT 78.870 169.820 79.190 170.080 ;
        RECT 79.420 170.065 79.560 170.220 ;
        RECT 80.340 170.065 80.480 170.560 ;
        RECT 81.170 170.360 81.490 170.420 ;
        RECT 81.170 170.220 83.240 170.360 ;
        RECT 81.170 170.160 81.490 170.220 ;
        RECT 79.345 169.835 79.635 170.065 ;
        RECT 80.265 169.835 80.555 170.065 ;
        RECT 81.630 170.020 81.950 170.080 ;
        RECT 83.100 170.065 83.240 170.220 ;
        RECT 84.020 170.065 84.160 170.560 ;
        RECT 84.850 170.360 85.170 170.420 ;
        RECT 85.785 170.360 86.075 170.405 ;
        RECT 84.850 170.220 86.075 170.360 ;
        RECT 84.850 170.160 85.170 170.220 ;
        RECT 85.785 170.175 86.075 170.220 ;
        RECT 82.105 170.020 82.395 170.065 ;
        RECT 81.630 169.880 82.395 170.020 ;
        RECT 79.790 169.680 80.110 169.740 ;
        RECT 76.660 169.540 80.110 169.680 ;
        RECT 75.665 169.495 75.955 169.540 ;
        RECT 76.110 169.480 76.430 169.540 ;
        RECT 79.790 169.480 80.110 169.540 ;
        RECT 80.340 169.680 80.480 169.835 ;
        RECT 81.630 169.820 81.950 169.880 ;
        RECT 82.105 169.835 82.395 169.880 ;
        RECT 82.565 169.835 82.855 170.065 ;
        RECT 83.025 169.835 83.315 170.065 ;
        RECT 83.945 169.835 84.235 170.065 ;
        RECT 85.325 170.020 85.615 170.065 ;
        RECT 84.940 169.880 85.615 170.020 ;
        RECT 80.710 169.680 81.030 169.740 ;
        RECT 80.340 169.540 81.030 169.680 ;
        RECT 71.510 169.340 71.800 169.385 ;
        RECT 73.080 169.340 73.370 169.385 ;
        RECT 75.180 169.340 75.470 169.385 ;
        RECT 80.340 169.340 80.480 169.540 ;
        RECT 80.710 169.480 81.030 169.540 ;
        RECT 71.510 169.200 75.470 169.340 ;
        RECT 71.510 169.155 71.800 169.200 ;
        RECT 73.080 169.155 73.370 169.200 ;
        RECT 75.180 169.155 75.470 169.200 ;
        RECT 76.660 169.200 80.480 169.340 ;
        RECT 82.090 169.340 82.410 169.400 ;
        RECT 82.640 169.340 82.780 169.835 ;
        RECT 84.940 169.740 85.080 169.880 ;
        RECT 85.325 169.835 85.615 169.880 ;
        RECT 85.860 169.740 86.000 170.175 ;
        RECT 86.230 169.820 86.550 170.080 ;
        RECT 87.165 169.835 87.455 170.065 ;
        RECT 84.850 169.480 85.170 169.740 ;
        RECT 85.770 169.480 86.090 169.740 ;
        RECT 87.240 169.340 87.380 169.835 ;
        RECT 82.090 169.200 82.780 169.340 ;
        RECT 83.100 169.200 87.380 169.340 ;
        RECT 76.660 169.000 76.800 169.200 ;
        RECT 82.090 169.140 82.410 169.200 ;
        RECT 70.680 168.860 76.800 169.000 ;
        RECT 77.030 168.800 77.350 169.060 ;
        RECT 78.410 169.000 78.730 169.060 ;
        RECT 80.725 169.000 81.015 169.045 ;
        RECT 78.410 168.860 81.015 169.000 ;
        RECT 78.410 168.800 78.730 168.860 ;
        RECT 80.725 168.815 81.015 168.860 ;
        RECT 81.170 169.000 81.490 169.060 ;
        RECT 83.100 169.000 83.240 169.200 ;
        RECT 81.170 168.860 83.240 169.000 ;
        RECT 81.170 168.800 81.490 168.860 ;
        RECT 84.390 168.800 84.710 169.060 ;
        RECT 12.100 168.180 89.840 168.660 ;
        RECT 45.765 167.980 46.055 168.025 ;
        RECT 47.130 167.980 47.450 168.040 ;
        RECT 45.765 167.840 47.450 167.980 ;
        RECT 45.765 167.795 46.055 167.840 ;
        RECT 47.130 167.780 47.450 167.840 ;
        RECT 51.285 167.980 51.575 168.025 ;
        RECT 52.190 167.980 52.510 168.040 ;
        RECT 51.285 167.840 52.510 167.980 ;
        RECT 51.285 167.795 51.575 167.840 ;
        RECT 39.350 167.640 39.640 167.685 ;
        RECT 41.450 167.640 41.740 167.685 ;
        RECT 43.020 167.640 43.310 167.685 ;
        RECT 39.350 167.500 43.310 167.640 ;
        RECT 39.350 167.455 39.640 167.500 ;
        RECT 41.450 167.455 41.740 167.500 ;
        RECT 43.020 167.455 43.310 167.500 ;
        RECT 39.745 167.300 40.035 167.345 ;
        RECT 40.935 167.300 41.225 167.345 ;
        RECT 43.455 167.300 43.745 167.345 ;
        RECT 39.745 167.160 43.745 167.300 ;
        RECT 39.745 167.115 40.035 167.160 ;
        RECT 40.935 167.115 41.225 167.160 ;
        RECT 43.455 167.115 43.745 167.160 ;
        RECT 48.510 167.100 48.830 167.360 ;
        RECT 38.865 166.960 39.155 167.005 ;
        RECT 38.865 166.820 41.150 166.960 ;
        RECT 38.865 166.775 39.155 166.820 ;
        RECT 41.010 166.680 41.150 166.820 ;
        RECT 47.130 166.760 47.450 167.020 ;
        RECT 48.970 166.960 49.290 167.020 ;
        RECT 49.445 166.960 49.735 167.005 ;
        RECT 48.970 166.820 49.735 166.960 ;
        RECT 48.970 166.760 49.290 166.820 ;
        RECT 49.445 166.775 49.735 166.820 ;
        RECT 49.905 166.960 50.195 167.005 ;
        RECT 51.360 166.960 51.500 167.795 ;
        RECT 52.190 167.780 52.510 167.840 ;
        RECT 64.150 167.980 64.470 168.040 ;
        RECT 67.385 167.980 67.675 168.025 ;
        RECT 75.190 167.980 75.510 168.040 ;
        RECT 64.150 167.840 75.510 167.980 ;
        RECT 64.150 167.780 64.470 167.840 ;
        RECT 67.385 167.795 67.675 167.840 ;
        RECT 75.190 167.780 75.510 167.840 ;
        RECT 75.650 167.780 75.970 168.040 ;
        RECT 83.470 167.980 83.790 168.040 ;
        RECT 83.945 167.980 84.235 168.025 ;
        RECT 83.470 167.840 84.235 167.980 ;
        RECT 83.470 167.780 83.790 167.840 ;
        RECT 83.945 167.795 84.235 167.840 ;
        RECT 55.450 167.640 55.740 167.685 ;
        RECT 57.550 167.640 57.840 167.685 ;
        RECT 59.120 167.640 59.410 167.685 ;
        RECT 55.450 167.500 59.410 167.640 ;
        RECT 55.450 167.455 55.740 167.500 ;
        RECT 57.550 167.455 57.840 167.500 ;
        RECT 59.120 167.455 59.410 167.500 ;
        RECT 60.470 167.640 60.790 167.700 ;
        RECT 61.390 167.640 61.710 167.700 ;
        RECT 61.865 167.640 62.155 167.685 ;
        RECT 60.470 167.500 62.155 167.640 ;
        RECT 60.470 167.440 60.790 167.500 ;
        RECT 61.390 167.440 61.710 167.500 ;
        RECT 61.865 167.455 62.155 167.500 ;
        RECT 62.325 167.455 62.615 167.685 ;
        RECT 70.130 167.640 70.420 167.685 ;
        RECT 71.700 167.640 71.990 167.685 ;
        RECT 73.800 167.640 74.090 167.685 ;
        RECT 70.130 167.500 74.090 167.640 ;
        RECT 70.130 167.455 70.420 167.500 ;
        RECT 71.700 167.455 71.990 167.500 ;
        RECT 73.800 167.455 74.090 167.500 ;
        RECT 77.530 167.640 77.820 167.685 ;
        RECT 79.630 167.640 79.920 167.685 ;
        RECT 81.200 167.640 81.490 167.685 ;
        RECT 77.530 167.500 81.490 167.640 ;
        RECT 77.530 167.455 77.820 167.500 ;
        RECT 79.630 167.455 79.920 167.500 ;
        RECT 81.200 167.455 81.490 167.500 ;
        RECT 86.690 167.640 87.010 167.700 ;
        RECT 87.625 167.640 87.915 167.685 ;
        RECT 86.690 167.500 87.915 167.640 ;
        RECT 55.845 167.300 56.135 167.345 ;
        RECT 57.035 167.300 57.325 167.345 ;
        RECT 59.555 167.300 59.845 167.345 ;
        RECT 55.845 167.160 59.845 167.300 ;
        RECT 55.845 167.115 56.135 167.160 ;
        RECT 57.035 167.115 57.325 167.160 ;
        RECT 59.555 167.115 59.845 167.160 ;
        RECT 49.905 166.820 51.500 166.960 ;
        RECT 53.570 166.960 53.890 167.020 ;
        RECT 54.045 166.960 54.335 167.005 ;
        RECT 53.570 166.820 54.335 166.960 ;
        RECT 49.905 166.775 50.195 166.820 ;
        RECT 53.570 166.760 53.890 166.820 ;
        RECT 54.045 166.775 54.335 166.820 ;
        RECT 54.950 166.760 55.270 167.020 ;
        RECT 56.300 166.960 56.590 167.005 ;
        RECT 62.400 166.960 62.540 167.455 ;
        RECT 86.690 167.440 87.010 167.500 ;
        RECT 87.625 167.455 87.915 167.500 ;
        RECT 100.050 167.500 100.880 170.840 ;
        RECT 108.930 170.540 116.850 170.550 ;
        RECT 105.160 170.530 116.850 170.540 ;
        RECT 101.540 170.410 116.850 170.530 ;
        RECT 101.540 170.400 116.875 170.410 ;
        RECT 101.500 170.280 116.875 170.400 ;
        RECT 101.500 170.170 105.500 170.280 ;
        RECT 101.110 169.830 101.340 170.120 ;
        RECT 101.560 169.830 105.450 170.170 ;
        RECT 105.660 169.830 105.890 170.120 ;
        RECT 101.110 168.460 105.890 169.830 ;
        RECT 101.110 168.160 101.340 168.460 ;
        RECT 105.660 168.160 105.890 168.460 ;
        RECT 101.500 167.880 105.500 168.110 ;
        RECT 101.750 167.650 105.320 167.880 ;
        RECT 101.750 167.500 105.440 167.650 ;
        RECT 63.230 167.300 63.550 167.360 ;
        RECT 64.625 167.300 64.915 167.345 ;
        RECT 63.230 167.160 64.915 167.300 ;
        RECT 63.230 167.100 63.550 167.160 ;
        RECT 64.625 167.115 64.915 167.160 ;
        RECT 65.085 167.115 65.375 167.345 ;
        RECT 69.695 167.300 69.985 167.345 ;
        RECT 72.215 167.300 72.505 167.345 ;
        RECT 73.405 167.300 73.695 167.345 ;
        RECT 77.925 167.300 78.215 167.345 ;
        RECT 79.115 167.300 79.405 167.345 ;
        RECT 81.635 167.300 81.925 167.345 ;
        RECT 86.230 167.300 86.550 167.360 ;
        RECT 88.530 167.300 88.850 167.360 ;
        RECT 69.695 167.160 73.695 167.300 ;
        RECT 69.695 167.115 69.985 167.160 ;
        RECT 72.215 167.115 72.505 167.160 ;
        RECT 73.405 167.115 73.695 167.160 ;
        RECT 74.405 167.160 75.420 167.300 ;
        RECT 65.160 166.960 65.300 167.115 ;
        RECT 74.405 167.005 74.545 167.160 ;
        RECT 75.280 167.020 75.420 167.160 ;
        RECT 77.925 167.160 81.925 167.300 ;
        RECT 77.925 167.115 78.215 167.160 ;
        RECT 79.115 167.115 79.405 167.160 ;
        RECT 81.635 167.115 81.925 167.160 ;
        RECT 85.860 167.160 88.850 167.300 ;
        RECT 100.050 167.240 105.440 167.500 ;
        RECT 106.690 167.330 107.310 170.280 ;
        RECT 108.875 170.180 116.875 170.280 ;
        RECT 108.930 170.170 116.850 170.180 ;
        RECT 108.440 169.470 108.670 170.130 ;
        RECT 109.450 169.470 110.450 169.560 ;
        RECT 117.080 169.470 117.310 170.130 ;
        RECT 108.440 168.650 117.310 169.470 ;
        RECT 108.440 168.170 108.670 168.650 ;
        RECT 109.450 168.560 110.450 168.650 ;
        RECT 117.080 168.170 117.310 168.650 ;
        RECT 108.875 167.890 116.875 168.120 ;
        RECT 56.300 166.820 62.540 166.960 ;
        RECT 62.860 166.820 65.300 166.960 ;
        RECT 56.300 166.775 56.590 166.820 ;
        RECT 40.230 166.665 40.550 166.680 ;
        RECT 40.200 166.435 40.550 166.665 ;
        RECT 41.010 166.480 41.470 166.680 ;
        RECT 40.230 166.420 40.550 166.435 ;
        RECT 41.150 166.420 41.470 166.480 ;
        RECT 48.065 166.620 48.355 166.665 ;
        RECT 50.810 166.620 51.130 166.680 ;
        RECT 48.065 166.480 51.130 166.620 ;
        RECT 48.065 166.435 48.355 166.480 ;
        RECT 50.810 166.420 51.130 166.480 ;
        RECT 60.010 166.620 60.330 166.680 ;
        RECT 62.860 166.620 63.000 166.820 ;
        RECT 74.285 166.775 74.575 167.005 ;
        RECT 74.745 166.775 75.035 167.005 ;
        RECT 75.190 166.960 75.510 167.020 ;
        RECT 76.110 166.960 76.430 167.020 ;
        RECT 77.045 166.960 77.335 167.005 ;
        RECT 81.170 166.960 81.490 167.020 ;
        RECT 82.090 166.960 82.410 167.020 ;
        RECT 75.190 166.820 81.490 166.960 ;
        RECT 60.010 166.480 63.000 166.620 ;
        RECT 71.970 166.620 72.290 166.680 ;
        RECT 72.950 166.620 73.240 166.665 ;
        RECT 71.970 166.480 73.240 166.620 ;
        RECT 60.010 166.420 60.330 166.480 ;
        RECT 71.970 166.420 72.290 166.480 ;
        RECT 72.950 166.435 73.240 166.480 ;
        RECT 74.820 166.340 74.960 166.775 ;
        RECT 75.190 166.760 75.510 166.820 ;
        RECT 76.110 166.760 76.430 166.820 ;
        RECT 77.045 166.775 77.335 166.820 ;
        RECT 81.170 166.760 81.490 166.820 ;
        RECT 81.720 166.820 82.410 166.960 ;
        RECT 78.410 166.665 78.730 166.680 ;
        RECT 78.380 166.435 78.730 166.665 ;
        RECT 78.410 166.420 78.730 166.435 ;
        RECT 78.870 166.620 79.190 166.680 ;
        RECT 81.720 166.620 81.860 166.820 ;
        RECT 82.090 166.760 82.410 166.820 ;
        RECT 82.550 166.960 82.870 167.020 ;
        RECT 85.860 167.005 86.000 167.160 ;
        RECT 86.230 167.100 86.550 167.160 ;
        RECT 88.530 167.100 88.850 167.160 ;
        RECT 100.010 167.220 105.440 167.240 ;
        RECT 84.865 166.960 85.155 167.005 ;
        RECT 82.550 166.820 85.155 166.960 ;
        RECT 82.550 166.760 82.870 166.820 ;
        RECT 84.865 166.775 85.155 166.820 ;
        RECT 85.785 166.775 86.075 167.005 ;
        RECT 86.705 166.960 86.995 167.005 ;
        RECT 87.150 166.960 87.470 167.020 ;
        RECT 86.705 166.820 87.470 166.960 ;
        RECT 86.705 166.775 86.995 166.820 ;
        RECT 87.150 166.760 87.470 166.820 ;
        RECT 100.010 166.760 105.450 167.220 ;
        RECT 78.870 166.480 81.860 166.620 ;
        RECT 78.870 166.420 79.190 166.480 ;
        RECT 86.245 166.435 86.535 166.665 ;
        RECT 46.210 166.080 46.530 166.340 ;
        RECT 48.525 166.280 48.815 166.325 ;
        RECT 48.970 166.280 49.290 166.340 ;
        RECT 48.525 166.140 49.290 166.280 ;
        RECT 48.525 166.095 48.815 166.140 ;
        RECT 48.970 166.080 49.290 166.140 ;
        RECT 64.150 166.080 64.470 166.340 ;
        RECT 74.730 166.080 75.050 166.340 ;
        RECT 86.320 166.280 86.460 166.435 ;
        RECT 87.150 166.280 87.470 166.340 ;
        RECT 86.320 166.140 87.470 166.280 ;
        RECT 87.150 166.080 87.470 166.140 ;
        RECT 12.100 165.460 89.840 165.940 ;
        RECT 100.010 165.410 102.050 166.760 ;
        RECT 103.800 166.750 105.450 166.760 ;
        RECT 102.490 165.480 103.490 166.200 ;
        RECT 103.800 165.940 104.110 166.750 ;
        RECT 104.570 166.470 105.450 166.750 ;
        RECT 105.690 166.930 107.310 167.330 ;
        RECT 108.960 166.980 116.830 167.890 ;
        RECT 104.510 166.240 105.510 166.470 ;
        RECT 105.690 166.280 106.040 166.930 ;
        RECT 106.690 166.920 107.310 166.930 ;
        RECT 108.875 166.750 116.875 166.980 ;
        RECT 108.960 166.740 116.830 166.750 ;
        RECT 104.570 166.030 105.450 166.050 ;
        RECT 103.840 165.650 104.110 165.940 ;
        RECT 104.510 165.800 105.510 166.030 ;
        RECT 105.670 165.990 106.040 166.280 ;
        RECT 105.700 165.930 106.040 165.990 ;
        RECT 106.800 166.600 107.560 166.650 ;
        RECT 108.440 166.600 108.670 166.700 ;
        RECT 106.800 166.390 108.670 166.600 ;
        RECT 117.080 166.390 117.310 166.700 ;
        RECT 106.800 165.970 109.340 166.390 ;
        RECT 116.710 165.970 117.310 166.390 ;
        RECT 104.570 165.650 105.450 165.800 ;
        RECT 104.580 165.480 105.310 165.650 ;
        RECT 43.450 165.260 43.770 165.320 ;
        RECT 43.925 165.260 44.215 165.305 ;
        RECT 43.450 165.120 44.215 165.260 ;
        RECT 43.450 165.060 43.770 165.120 ;
        RECT 43.925 165.075 44.215 165.120 ;
        RECT 61.865 165.260 62.155 165.305 ;
        RECT 62.770 165.260 63.090 165.320 ;
        RECT 66.910 165.260 67.230 165.320 ;
        RECT 61.865 165.120 67.230 165.260 ;
        RECT 61.865 165.075 62.155 165.120 ;
        RECT 62.770 165.060 63.090 165.120 ;
        RECT 66.910 165.060 67.230 165.120 ;
        RECT 77.950 165.260 78.270 165.320 ;
        RECT 81.185 165.260 81.475 165.305 ;
        RECT 77.950 165.120 81.475 165.260 ;
        RECT 77.950 165.060 78.270 165.120 ;
        RECT 81.185 165.075 81.475 165.120 ;
        RECT 46.210 164.920 46.530 164.980 ;
        RECT 47.145 164.920 47.435 164.965 ;
        RECT 75.190 164.920 75.510 164.980 ;
        RECT 46.210 164.780 47.435 164.920 ;
        RECT 46.210 164.720 46.530 164.780 ;
        RECT 47.145 164.735 47.435 164.780 ;
        RECT 71.140 164.780 75.510 164.920 ;
        RECT 42.070 164.580 42.390 164.640 ;
        RECT 44.370 164.580 44.690 164.640 ;
        RECT 48.970 164.625 49.290 164.640 ;
        RECT 45.305 164.580 45.595 164.625 ;
        RECT 48.940 164.580 49.290 164.625 ;
        RECT 42.070 164.440 45.595 164.580 ;
        RECT 48.775 164.440 49.290 164.580 ;
        RECT 42.070 164.380 42.390 164.440 ;
        RECT 44.370 164.380 44.690 164.440 ;
        RECT 45.305 164.395 45.595 164.440 ;
        RECT 48.940 164.395 49.290 164.440 ;
        RECT 48.970 164.380 49.290 164.395 ;
        RECT 54.950 164.380 55.270 164.640 ;
        RECT 56.330 164.625 56.650 164.640 ;
        RECT 56.300 164.395 56.650 164.625 ;
        RECT 56.330 164.380 56.650 164.395 ;
        RECT 68.290 164.580 68.610 164.640 ;
        RECT 71.140 164.625 71.280 164.780 ;
        RECT 69.730 164.580 70.020 164.625 ;
        RECT 68.290 164.440 70.020 164.580 ;
        RECT 68.290 164.380 68.610 164.440 ;
        RECT 69.730 164.395 70.020 164.440 ;
        RECT 71.065 164.395 71.355 164.625 ;
        RECT 71.510 164.380 71.830 164.640 ;
        RECT 74.360 164.625 74.500 164.780 ;
        RECT 75.190 164.720 75.510 164.780 ;
        RECT 77.490 164.920 77.810 164.980 ;
        RECT 81.645 164.920 81.935 164.965 ;
        RECT 77.490 164.780 81.935 164.920 ;
        RECT 77.490 164.720 77.810 164.780 ;
        RECT 81.645 164.735 81.935 164.780 ;
        RECT 73.365 164.395 73.655 164.625 ;
        RECT 74.285 164.395 74.575 164.625 ;
        RECT 37.010 164.240 37.330 164.300 ;
        RECT 43.005 164.240 43.295 164.285 ;
        RECT 37.010 164.100 43.295 164.240 ;
        RECT 37.010 164.040 37.330 164.100 ;
        RECT 43.005 164.055 43.295 164.100 ;
        RECT 44.830 164.040 45.150 164.300 ;
        RECT 46.670 164.040 46.990 164.300 ;
        RECT 47.605 164.055 47.895 164.285 ;
        RECT 48.485 164.240 48.775 164.285 ;
        RECT 49.675 164.240 49.965 164.285 ;
        RECT 52.195 164.240 52.485 164.285 ;
        RECT 48.485 164.100 52.485 164.240 ;
        RECT 48.485 164.055 48.775 164.100 ;
        RECT 49.675 164.055 49.965 164.100 ;
        RECT 52.195 164.055 52.485 164.100 ;
        RECT 55.845 164.240 56.135 164.285 ;
        RECT 57.035 164.240 57.325 164.285 ;
        RECT 59.555 164.240 59.845 164.285 ;
        RECT 55.845 164.100 59.845 164.240 ;
        RECT 55.845 164.055 56.135 164.100 ;
        RECT 57.035 164.055 57.325 164.100 ;
        RECT 59.555 164.055 59.845 164.100 ;
        RECT 66.475 164.240 66.765 164.285 ;
        RECT 68.995 164.240 69.285 164.285 ;
        RECT 70.185 164.240 70.475 164.285 ;
        RECT 66.475 164.100 70.475 164.240 ;
        RECT 73.440 164.240 73.580 164.395 ;
        RECT 74.730 164.380 75.050 164.640 ;
        RECT 75.620 164.580 75.910 164.625 ;
        RECT 77.030 164.580 77.350 164.640 ;
        RECT 75.620 164.440 77.350 164.580 ;
        RECT 75.620 164.395 75.910 164.440 ;
        RECT 77.030 164.380 77.350 164.440 ;
        RECT 82.550 164.380 82.870 164.640 ;
        RECT 88.070 164.380 88.390 164.640 ;
        RECT 74.820 164.240 74.960 164.380 ;
        RECT 73.440 164.100 74.960 164.240 ;
        RECT 75.165 164.240 75.455 164.285 ;
        RECT 76.355 164.240 76.645 164.285 ;
        RECT 78.875 164.240 79.165 164.285 ;
        RECT 75.165 164.100 79.165 164.240 ;
        RECT 66.475 164.055 66.765 164.100 ;
        RECT 68.995 164.055 69.285 164.100 ;
        RECT 70.185 164.055 70.475 164.100 ;
        RECT 75.165 164.055 75.455 164.100 ;
        RECT 76.355 164.055 76.645 164.100 ;
        RECT 78.875 164.055 79.165 164.100 ;
        RECT 83.470 164.240 83.790 164.300 ;
        RECT 86.705 164.240 86.995 164.285 ;
        RECT 83.470 164.100 86.995 164.240 ;
        RECT 41.150 163.900 41.470 163.960 ;
        RECT 47.680 163.900 47.820 164.055 ;
        RECT 83.470 164.040 83.790 164.100 ;
        RECT 86.705 164.055 86.995 164.100 ;
        RECT 41.150 163.760 47.820 163.900 ;
        RECT 48.090 163.900 48.380 163.945 ;
        RECT 50.190 163.900 50.480 163.945 ;
        RECT 51.760 163.900 52.050 163.945 ;
        RECT 48.090 163.760 52.050 163.900 ;
        RECT 41.150 163.700 41.470 163.760 ;
        RECT 48.090 163.715 48.380 163.760 ;
        RECT 50.190 163.715 50.480 163.760 ;
        RECT 51.760 163.715 52.050 163.760 ;
        RECT 55.450 163.900 55.740 163.945 ;
        RECT 57.550 163.900 57.840 163.945 ;
        RECT 59.120 163.900 59.410 163.945 ;
        RECT 55.450 163.760 59.410 163.900 ;
        RECT 55.450 163.715 55.740 163.760 ;
        RECT 57.550 163.715 57.840 163.760 ;
        RECT 59.120 163.715 59.410 163.760 ;
        RECT 66.910 163.900 67.200 163.945 ;
        RECT 68.480 163.900 68.770 163.945 ;
        RECT 70.580 163.900 70.870 163.945 ;
        RECT 74.770 163.900 75.060 163.945 ;
        RECT 76.870 163.900 77.160 163.945 ;
        RECT 78.440 163.900 78.730 163.945 ;
        RECT 85.770 163.900 86.090 163.960 ;
        RECT 88.070 163.900 88.390 163.960 ;
        RECT 66.910 163.760 70.870 163.900 ;
        RECT 66.910 163.715 67.200 163.760 ;
        RECT 68.480 163.715 68.770 163.760 ;
        RECT 70.580 163.715 70.870 163.760 ;
        RECT 71.600 163.760 74.500 163.900 ;
        RECT 40.230 163.360 40.550 163.620 ;
        RECT 53.570 163.560 53.890 163.620 ;
        RECT 54.505 163.560 54.795 163.605 ;
        RECT 53.570 163.420 54.795 163.560 ;
        RECT 53.570 163.360 53.890 163.420 ;
        RECT 54.505 163.375 54.795 163.420 ;
        RECT 64.165 163.560 64.455 163.605 ;
        RECT 65.990 163.560 66.310 163.620 ;
        RECT 64.165 163.420 66.310 163.560 ;
        RECT 64.165 163.375 64.455 163.420 ;
        RECT 65.990 163.360 66.310 163.420 ;
        RECT 66.450 163.560 66.770 163.620 ;
        RECT 71.600 163.560 71.740 163.760 ;
        RECT 66.450 163.420 71.740 163.560 ;
        RECT 74.360 163.560 74.500 163.760 ;
        RECT 74.770 163.760 78.730 163.900 ;
        RECT 74.770 163.715 75.060 163.760 ;
        RECT 76.870 163.715 77.160 163.760 ;
        RECT 78.440 163.715 78.730 163.760 ;
        RECT 83.100 163.760 88.390 163.900 ;
        RECT 83.100 163.560 83.240 163.760 ;
        RECT 85.770 163.700 86.090 163.760 ;
        RECT 88.070 163.700 88.390 163.760 ;
        RECT 74.360 163.420 83.240 163.560 ;
        RECT 83.485 163.560 83.775 163.605 ;
        RECT 85.310 163.560 85.630 163.620 ;
        RECT 83.485 163.420 85.630 163.560 ;
        RECT 66.450 163.360 66.770 163.420 ;
        RECT 83.485 163.375 83.775 163.420 ;
        RECT 85.310 163.360 85.630 163.420 ;
        RECT 12.100 162.740 89.840 163.220 ;
        RECT 37.010 162.340 37.330 162.600 ;
        RECT 46.670 162.540 46.990 162.600 ;
        RECT 51.285 162.540 51.575 162.585 ;
        RECT 46.670 162.400 51.575 162.540 ;
        RECT 46.670 162.340 46.990 162.400 ;
        RECT 51.285 162.355 51.575 162.400 ;
        RECT 55.870 162.340 56.190 162.600 ;
        RECT 56.330 162.540 56.650 162.600 ;
        RECT 57.265 162.540 57.555 162.585 ;
        RECT 56.330 162.400 57.555 162.540 ;
        RECT 56.330 162.340 56.650 162.400 ;
        RECT 57.265 162.355 57.555 162.400 ;
        RECT 65.990 162.540 66.310 162.600 ;
        RECT 65.990 162.400 75.880 162.540 ;
        RECT 65.990 162.340 66.310 162.400 ;
        RECT 39.770 162.200 40.060 162.245 ;
        RECT 41.340 162.200 41.630 162.245 ;
        RECT 43.440 162.200 43.730 162.245 ;
        RECT 48.970 162.200 49.290 162.260 ;
        RECT 39.770 162.060 43.730 162.200 ;
        RECT 39.770 162.015 40.060 162.060 ;
        RECT 41.340 162.015 41.630 162.060 ;
        RECT 43.440 162.015 43.730 162.060 ;
        RECT 45.380 162.060 49.290 162.200 ;
        RECT 39.335 161.860 39.625 161.905 ;
        RECT 41.855 161.860 42.145 161.905 ;
        RECT 43.045 161.860 43.335 161.905 ;
        RECT 39.335 161.720 43.335 161.860 ;
        RECT 39.335 161.675 39.625 161.720 ;
        RECT 41.855 161.675 42.145 161.720 ;
        RECT 43.045 161.675 43.335 161.720 ;
        RECT 38.850 161.520 39.170 161.580 ;
        RECT 41.150 161.520 41.470 161.580 ;
        RECT 43.910 161.520 44.230 161.580 ;
        RECT 45.380 161.565 45.520 162.060 ;
        RECT 48.970 162.000 49.290 162.060 ;
        RECT 54.950 162.200 55.270 162.260 ;
        RECT 61.890 162.200 62.180 162.245 ;
        RECT 63.990 162.200 64.280 162.245 ;
        RECT 65.560 162.200 65.850 162.245 ;
        RECT 54.950 162.060 61.620 162.200 ;
        RECT 54.950 162.000 55.270 162.060 ;
        RECT 48.065 161.860 48.355 161.905 ;
        RECT 48.065 161.720 52.880 161.860 ;
        RECT 48.065 161.675 48.355 161.720 ;
        RECT 52.740 161.580 52.880 161.720 ;
        RECT 56.330 161.660 56.650 161.920 ;
        RECT 57.710 161.860 58.030 161.920 ;
        RECT 60.010 161.860 60.330 161.920 ;
        RECT 61.480 161.905 61.620 162.060 ;
        RECT 61.890 162.060 65.850 162.200 ;
        RECT 61.890 162.015 62.180 162.060 ;
        RECT 63.990 162.015 64.280 162.060 ;
        RECT 65.560 162.015 65.850 162.060 ;
        RECT 68.765 162.015 69.055 162.245 ;
        RECT 57.710 161.720 60.330 161.860 ;
        RECT 57.710 161.660 58.030 161.720 ;
        RECT 60.010 161.660 60.330 161.720 ;
        RECT 61.405 161.675 61.695 161.905 ;
        RECT 62.285 161.860 62.575 161.905 ;
        RECT 63.475 161.860 63.765 161.905 ;
        RECT 65.995 161.860 66.285 161.905 ;
        RECT 62.285 161.720 66.285 161.860 ;
        RECT 62.285 161.675 62.575 161.720 ;
        RECT 63.475 161.675 63.765 161.720 ;
        RECT 65.995 161.675 66.285 161.720 ;
        RECT 38.850 161.380 44.230 161.520 ;
        RECT 38.850 161.320 39.170 161.380 ;
        RECT 41.150 161.320 41.470 161.380 ;
        RECT 43.910 161.320 44.230 161.380 ;
        RECT 44.845 161.335 45.135 161.565 ;
        RECT 45.305 161.335 45.595 161.565 ;
        RECT 46.225 161.520 46.515 161.565 ;
        RECT 47.605 161.520 47.895 161.565 ;
        RECT 46.225 161.380 47.895 161.520 ;
        RECT 46.225 161.335 46.515 161.380 ;
        RECT 47.605 161.335 47.895 161.380 ;
        RECT 41.610 161.180 41.930 161.240 ;
        RECT 42.590 161.180 42.880 161.225 ;
        RECT 41.610 161.040 42.880 161.180 ;
        RECT 44.920 161.180 45.060 161.335 ;
        RECT 48.510 161.320 48.830 161.580 ;
        RECT 48.970 161.320 49.290 161.580 ;
        RECT 49.905 161.520 50.195 161.565 ;
        RECT 50.810 161.520 51.130 161.580 ;
        RECT 49.905 161.380 51.130 161.520 ;
        RECT 49.905 161.335 50.195 161.380 ;
        RECT 50.810 161.320 51.130 161.380 ;
        RECT 52.190 161.320 52.510 161.580 ;
        RECT 52.650 161.320 52.970 161.580 ;
        RECT 53.585 161.335 53.875 161.565 ;
        RECT 48.600 161.180 48.740 161.320 ;
        RECT 53.660 161.180 53.800 161.335 ;
        RECT 54.030 161.320 54.350 161.580 ;
        RECT 55.425 161.520 55.715 161.565 ;
        RECT 57.250 161.520 57.570 161.580 ;
        RECT 55.425 161.380 57.570 161.520 ;
        RECT 55.425 161.335 55.715 161.380 ;
        RECT 57.250 161.320 57.570 161.380 ;
        RECT 59.105 161.520 59.395 161.565 ;
        RECT 68.840 161.520 68.980 162.015 ;
        RECT 70.130 161.860 70.450 161.920 ;
        RECT 75.740 161.905 75.880 162.400 ;
        RECT 88.070 162.340 88.390 162.600 ;
        RECT 79.330 162.000 79.650 162.260 ;
        RECT 81.670 162.200 81.960 162.245 ;
        RECT 83.770 162.200 84.060 162.245 ;
        RECT 85.340 162.200 85.630 162.245 ;
        RECT 81.670 162.060 85.630 162.200 ;
        RECT 81.670 162.015 81.960 162.060 ;
        RECT 83.770 162.015 84.060 162.060 ;
        RECT 85.340 162.015 85.630 162.060 ;
        RECT 71.525 161.860 71.815 161.905 ;
        RECT 70.130 161.720 71.815 161.860 ;
        RECT 70.130 161.660 70.450 161.720 ;
        RECT 71.525 161.675 71.815 161.720 ;
        RECT 75.665 161.675 75.955 161.905 ;
        RECT 79.420 161.860 79.560 162.000 ;
        RECT 82.065 161.860 82.355 161.905 ;
        RECT 83.255 161.860 83.545 161.905 ;
        RECT 85.775 161.860 86.065 161.905 ;
        RECT 76.200 161.720 80.480 161.860 ;
        RECT 59.105 161.380 68.980 161.520 ;
        RECT 69.670 161.520 69.990 161.580 ;
        RECT 76.200 161.520 76.340 161.720 ;
        RECT 69.670 161.380 76.340 161.520 ;
        RECT 76.570 161.520 76.890 161.580 ;
        RECT 78.410 161.520 78.730 161.580 ;
        RECT 76.570 161.380 78.730 161.520 ;
        RECT 59.105 161.335 59.395 161.380 ;
        RECT 69.670 161.320 69.990 161.380 ;
        RECT 76.570 161.320 76.890 161.380 ;
        RECT 78.410 161.320 78.730 161.380 ;
        RECT 78.885 161.335 79.175 161.565 ;
        RECT 79.345 161.520 79.635 161.565 ;
        RECT 79.790 161.520 80.110 161.580 ;
        RECT 80.340 161.565 80.480 161.720 ;
        RECT 82.065 161.720 86.065 161.860 ;
        RECT 82.065 161.675 82.355 161.720 ;
        RECT 83.255 161.675 83.545 161.720 ;
        RECT 85.775 161.675 86.065 161.720 ;
        RECT 100.010 161.770 100.780 165.410 ;
        RECT 102.460 164.360 105.310 165.480 ;
        RECT 105.700 165.180 106.050 165.930 ;
        RECT 106.800 165.810 108.670 165.970 ;
        RECT 106.800 165.760 107.560 165.810 ;
        RECT 108.440 165.740 108.670 165.810 ;
        RECT 117.080 165.740 117.310 165.970 ;
        RECT 108.875 165.460 116.875 165.690 ;
        RECT 105.700 165.120 105.990 165.180 ;
        RECT 105.610 165.000 105.990 165.120 ;
        RECT 108.970 165.060 116.830 165.460 ;
        RECT 117.640 165.060 118.600 174.540 ;
        RECT 119.930 174.510 125.370 174.620 ;
        RECT 128.810 174.600 138.700 174.700 ;
        RECT 139.960 175.280 140.860 176.800 ;
        RECT 146.460 176.380 147.710 176.820 ;
        RECT 144.400 176.370 149.640 176.380 ;
        RECT 141.450 176.270 156.750 176.370 ;
        RECT 141.450 176.260 156.785 176.270 ;
        RECT 141.410 176.140 156.785 176.260 ;
        RECT 141.410 176.030 145.410 176.140 ;
        RECT 146.460 176.060 148.200 176.140 ;
        RECT 148.780 176.060 156.785 176.140 ;
        RECT 146.460 175.980 147.710 176.060 ;
        RECT 148.785 176.040 156.785 176.060 ;
        RECT 141.020 175.730 141.250 175.980 ;
        RECT 145.570 175.840 145.800 175.980 ;
        RECT 148.350 175.840 148.580 175.990 ;
        RECT 145.570 175.730 148.580 175.840 ;
        RECT 156.990 175.730 157.220 175.990 ;
        RECT 141.020 175.290 157.220 175.730 ;
        RECT 139.960 174.670 140.790 175.280 ;
        RECT 141.020 175.020 141.250 175.290 ;
        RECT 145.570 175.260 157.220 175.290 ;
        RECT 145.570 175.170 148.580 175.260 ;
        RECT 145.570 175.020 145.800 175.170 ;
        RECT 148.350 175.030 148.580 175.170 ;
        RECT 156.990 175.030 157.220 175.260 ;
        RECT 141.410 174.740 145.410 174.970 ;
        RECT 148.785 174.760 156.785 174.980 ;
        RECT 157.550 174.760 158.510 176.800 ;
        RECT 148.785 174.750 158.510 174.760 ;
        RECT 141.410 174.670 145.400 174.740 ;
        RECT 128.810 174.540 138.480 174.600 ;
        RECT 119.930 174.420 123.060 174.510 ;
        RECT 136.550 174.490 138.480 174.540 ;
        RECT 119.930 171.150 120.760 174.420 ;
        RECT 124.410 173.960 129.660 173.970 ;
        RECT 124.410 173.850 136.720 173.960 ;
        RECT 121.440 173.790 136.720 173.850 ;
        RECT 121.440 173.780 136.755 173.790 ;
        RECT 121.380 173.650 136.755 173.780 ;
        RECT 121.380 173.640 126.540 173.650 ;
        RECT 121.380 173.550 125.380 173.640 ;
        RECT 128.755 173.560 136.755 173.650 ;
        RECT 128.840 173.550 136.730 173.560 ;
        RECT 120.990 173.190 121.220 173.500 ;
        RECT 121.440 173.190 125.340 173.550 ;
        RECT 125.540 173.190 125.770 173.500 ;
        RECT 120.990 171.850 125.770 173.190 ;
        RECT 120.990 171.540 121.220 171.850 ;
        RECT 125.540 171.540 125.770 171.850 ;
        RECT 128.320 172.970 128.550 173.510 ;
        RECT 129.360 172.970 130.370 173.000 ;
        RECT 136.960 172.970 137.190 173.510 ;
        RECT 128.320 172.070 137.190 172.970 ;
        RECT 128.320 171.550 128.550 172.070 ;
        RECT 129.360 172.000 130.370 172.070 ;
        RECT 136.960 171.550 137.190 172.070 ;
        RECT 121.380 171.260 125.380 171.490 ;
        RECT 128.755 171.270 136.755 171.500 ;
        RECT 119.930 171.110 121.060 171.150 ;
        RECT 119.930 171.030 121.300 171.110 ;
        RECT 121.670 171.040 125.330 171.260 ;
        RECT 121.670 171.030 123.110 171.040 ;
        RECT 119.930 170.990 123.110 171.030 ;
        RECT 119.930 170.900 122.620 170.990 ;
        RECT 128.820 170.980 136.710 171.270 ;
        RECT 119.930 170.840 121.950 170.900 ;
        RECT 119.930 170.790 121.700 170.840 ;
        RECT 119.930 167.450 120.760 170.790 ;
        RECT 128.810 170.490 136.730 170.500 ;
        RECT 125.040 170.480 136.730 170.490 ;
        RECT 121.420 170.360 136.730 170.480 ;
        RECT 121.420 170.350 136.755 170.360 ;
        RECT 121.380 170.230 136.755 170.350 ;
        RECT 121.380 170.120 125.380 170.230 ;
        RECT 120.990 169.780 121.220 170.070 ;
        RECT 121.440 169.780 125.330 170.120 ;
        RECT 125.540 169.780 125.770 170.070 ;
        RECT 120.990 168.410 125.770 169.780 ;
        RECT 120.990 168.110 121.220 168.410 ;
        RECT 125.540 168.110 125.770 168.410 ;
        RECT 121.380 167.830 125.380 168.060 ;
        RECT 121.630 167.600 125.200 167.830 ;
        RECT 121.630 167.450 125.320 167.600 ;
        RECT 119.930 167.170 125.320 167.450 ;
        RECT 126.570 167.280 127.190 170.230 ;
        RECT 128.755 170.130 136.755 170.230 ;
        RECT 128.810 170.120 136.730 170.130 ;
        RECT 128.320 169.420 128.550 170.080 ;
        RECT 129.330 169.420 130.330 169.510 ;
        RECT 136.960 169.420 137.190 170.080 ;
        RECT 128.320 168.600 137.190 169.420 ;
        RECT 128.320 168.120 128.550 168.600 ;
        RECT 129.330 168.510 130.330 168.600 ;
        RECT 136.960 168.120 137.190 168.600 ;
        RECT 128.755 167.840 136.755 168.070 ;
        RECT 119.930 166.710 125.330 167.170 ;
        RECT 119.930 165.370 121.930 166.710 ;
        RECT 123.680 166.700 125.330 166.710 ;
        RECT 122.370 165.430 123.370 166.150 ;
        RECT 123.680 165.890 123.990 166.700 ;
        RECT 124.450 166.420 125.330 166.700 ;
        RECT 125.570 166.880 127.190 167.280 ;
        RECT 128.840 166.930 136.710 167.840 ;
        RECT 124.390 166.190 125.390 166.420 ;
        RECT 125.570 166.230 125.920 166.880 ;
        RECT 126.570 166.870 127.190 166.880 ;
        RECT 128.755 166.700 136.755 166.930 ;
        RECT 128.840 166.690 136.710 166.700 ;
        RECT 124.450 165.980 125.330 166.000 ;
        RECT 123.720 165.600 123.990 165.890 ;
        RECT 124.390 165.750 125.390 165.980 ;
        RECT 125.550 165.940 125.920 166.230 ;
        RECT 125.580 165.880 125.920 165.940 ;
        RECT 126.680 166.550 127.440 166.600 ;
        RECT 128.320 166.550 128.550 166.650 ;
        RECT 126.680 166.340 128.550 166.550 ;
        RECT 136.960 166.340 137.190 166.650 ;
        RECT 126.680 165.920 129.220 166.340 ;
        RECT 136.590 165.920 137.190 166.340 ;
        RECT 124.450 165.600 125.330 165.750 ;
        RECT 124.460 165.430 125.190 165.600 ;
        RECT 102.400 164.130 105.400 164.360 ;
        RECT 105.610 164.170 105.950 165.000 ;
        RECT 107.960 164.990 118.600 165.060 ;
        RECT 102.450 164.100 105.310 164.130 ;
        RECT 102.450 164.080 103.620 164.100 ;
        RECT 104.580 164.090 105.310 164.100 ;
        RECT 102.400 163.690 105.400 163.920 ;
        RECT 105.605 163.880 105.950 164.170 ;
        RECT 106.140 163.950 118.600 164.990 ;
        RECT 120.000 165.360 121.930 165.370 ;
        RECT 106.140 163.930 118.560 163.950 ;
        RECT 105.610 163.770 105.950 163.880 ;
        RECT 106.180 163.920 111.850 163.930 ;
        RECT 112.850 163.920 118.560 163.930 ;
        RECT 102.490 163.520 105.350 163.690 ;
        RECT 106.180 163.520 106.610 163.920 ;
        RECT 102.460 163.150 106.610 163.520 ;
        RECT 79.345 161.380 80.110 161.520 ;
        RECT 79.345 161.335 79.635 161.380 ;
        RECT 44.920 161.040 48.280 161.180 ;
        RECT 48.600 161.040 53.800 161.180 ;
        RECT 56.805 161.180 57.095 161.225 ;
        RECT 58.630 161.180 58.950 161.240 ;
        RECT 56.805 161.040 58.950 161.180 ;
        RECT 41.610 160.980 41.930 161.040 ;
        RECT 42.590 160.995 42.880 161.040 ;
        RECT 46.670 160.640 46.990 160.900 ;
        RECT 48.140 160.840 48.280 161.040 ;
        RECT 56.805 160.995 57.095 161.040 ;
        RECT 58.630 160.980 58.950 161.040 ;
        RECT 59.565 161.180 59.855 161.225 ;
        RECT 61.850 161.180 62.170 161.240 ;
        RECT 59.565 161.040 62.170 161.180 ;
        RECT 59.565 160.995 59.855 161.040 ;
        RECT 61.850 160.980 62.170 161.040 ;
        RECT 62.740 161.180 63.030 161.225 ;
        RECT 65.530 161.180 65.850 161.240 ;
        RECT 70.590 161.180 70.910 161.240 ;
        RECT 62.740 161.040 65.850 161.180 ;
        RECT 62.740 160.995 63.030 161.040 ;
        RECT 65.530 160.980 65.850 161.040 ;
        RECT 68.380 161.040 70.910 161.180 ;
        RECT 53.570 160.840 53.890 160.900 ;
        RECT 48.140 160.700 53.890 160.840 ;
        RECT 53.570 160.640 53.890 160.700 ;
        RECT 54.505 160.840 54.795 160.885 ;
        RECT 55.410 160.840 55.730 160.900 ;
        RECT 68.380 160.885 68.520 161.040 ;
        RECT 70.590 160.980 70.910 161.040 ;
        RECT 71.970 161.180 72.290 161.240 ;
        RECT 77.045 161.180 77.335 161.225 ;
        RECT 71.970 161.040 77.335 161.180 ;
        RECT 71.970 160.980 72.290 161.040 ;
        RECT 77.045 160.995 77.335 161.040 ;
        RECT 77.950 161.180 78.270 161.240 ;
        RECT 78.960 161.180 79.100 161.335 ;
        RECT 79.790 161.320 80.110 161.380 ;
        RECT 80.265 161.335 80.555 161.565 ;
        RECT 81.170 161.320 81.490 161.580 ;
        RECT 77.950 161.040 79.100 161.180 ;
        RECT 80.710 161.180 81.030 161.240 ;
        RECT 82.410 161.180 82.700 161.225 ;
        RECT 80.710 161.040 82.700 161.180 ;
        RECT 77.950 160.980 78.270 161.040 ;
        RECT 80.710 160.980 81.030 161.040 ;
        RECT 82.410 160.995 82.700 161.040 ;
        RECT 54.505 160.700 55.730 160.840 ;
        RECT 54.505 160.655 54.795 160.700 ;
        RECT 55.410 160.640 55.730 160.700 ;
        RECT 68.305 160.655 68.595 160.885 ;
        RECT 68.750 160.840 69.070 160.900 ;
        RECT 71.065 160.840 71.355 160.885 ;
        RECT 68.750 160.700 71.355 160.840 ;
        RECT 68.750 160.640 69.070 160.700 ;
        RECT 71.065 160.655 71.355 160.700 ;
        RECT 72.890 160.640 73.210 160.900 ;
        RECT 12.100 160.020 89.840 160.500 ;
        RECT 37.025 159.820 37.315 159.865 ;
        RECT 40.230 159.820 40.550 159.880 ;
        RECT 37.025 159.680 40.550 159.820 ;
        RECT 37.025 159.635 37.315 159.680 ;
        RECT 40.230 159.620 40.550 159.680 ;
        RECT 40.690 159.620 41.010 159.880 ;
        RECT 48.970 159.820 49.290 159.880 ;
        RECT 53.125 159.820 53.415 159.865 ;
        RECT 54.490 159.820 54.810 159.880 ;
        RECT 48.970 159.680 54.810 159.820 ;
        RECT 48.970 159.620 49.290 159.680 ;
        RECT 53.125 159.635 53.415 159.680 ;
        RECT 54.490 159.620 54.810 159.680 ;
        RECT 55.870 159.820 56.190 159.880 ;
        RECT 60.930 159.820 61.250 159.880 ;
        RECT 55.870 159.680 61.250 159.820 ;
        RECT 55.870 159.620 56.190 159.680 ;
        RECT 60.930 159.620 61.250 159.680 ;
        RECT 64.150 159.620 64.470 159.880 ;
        RECT 65.990 159.620 66.310 159.880 ;
        RECT 68.290 159.620 68.610 159.880 ;
        RECT 70.145 159.820 70.435 159.865 ;
        RECT 72.890 159.820 73.210 159.880 ;
        RECT 70.145 159.680 73.210 159.820 ;
        RECT 70.145 159.635 70.435 159.680 ;
        RECT 72.890 159.620 73.210 159.680 ;
        RECT 87.610 159.820 87.930 159.880 ;
        RECT 88.085 159.820 88.375 159.865 ;
        RECT 87.610 159.680 88.375 159.820 ;
        RECT 87.610 159.620 87.930 159.680 ;
        RECT 88.085 159.635 88.375 159.680 ;
        RECT 100.010 159.670 100.880 161.770 ;
        RECT 106.550 161.380 107.800 161.820 ;
        RECT 117.700 161.800 118.560 163.920 ;
        RECT 120.000 161.800 120.770 165.360 ;
        RECT 122.340 164.310 125.190 165.430 ;
        RECT 125.580 165.130 125.930 165.880 ;
        RECT 126.680 165.760 128.550 165.920 ;
        RECT 126.680 165.710 127.440 165.760 ;
        RECT 128.320 165.690 128.550 165.760 ;
        RECT 136.960 165.690 137.190 165.920 ;
        RECT 128.755 165.410 136.755 165.640 ;
        RECT 125.580 165.070 125.870 165.130 ;
        RECT 125.490 164.950 125.870 165.070 ;
        RECT 128.850 165.010 136.710 165.410 ;
        RECT 137.520 165.010 138.480 174.490 ;
        RECT 139.960 174.560 145.400 174.670 ;
        RECT 148.840 174.590 158.510 174.750 ;
        RECT 139.960 174.470 143.090 174.560 ;
        RECT 156.580 174.540 158.510 174.590 ;
        RECT 139.960 171.200 140.790 174.470 ;
        RECT 144.440 174.010 149.690 174.020 ;
        RECT 144.440 173.900 156.750 174.010 ;
        RECT 141.470 173.840 156.750 173.900 ;
        RECT 141.470 173.830 156.785 173.840 ;
        RECT 141.410 173.700 156.785 173.830 ;
        RECT 141.410 173.690 146.570 173.700 ;
        RECT 141.410 173.600 145.410 173.690 ;
        RECT 148.785 173.610 156.785 173.700 ;
        RECT 148.870 173.600 156.760 173.610 ;
        RECT 141.020 173.240 141.250 173.550 ;
        RECT 141.470 173.240 145.370 173.600 ;
        RECT 145.570 173.240 145.800 173.550 ;
        RECT 141.020 171.900 145.800 173.240 ;
        RECT 141.020 171.590 141.250 171.900 ;
        RECT 145.570 171.590 145.800 171.900 ;
        RECT 148.350 173.020 148.580 173.560 ;
        RECT 149.390 173.020 150.400 173.050 ;
        RECT 156.990 173.020 157.220 173.560 ;
        RECT 148.350 172.120 157.220 173.020 ;
        RECT 148.350 171.600 148.580 172.120 ;
        RECT 149.390 172.050 150.400 172.120 ;
        RECT 156.990 171.600 157.220 172.120 ;
        RECT 141.410 171.310 145.410 171.540 ;
        RECT 148.785 171.320 156.785 171.550 ;
        RECT 139.960 171.160 141.090 171.200 ;
        RECT 139.960 171.080 141.330 171.160 ;
        RECT 141.700 171.090 145.360 171.310 ;
        RECT 141.700 171.080 143.140 171.090 ;
        RECT 139.960 171.040 143.140 171.080 ;
        RECT 139.960 170.950 142.650 171.040 ;
        RECT 148.850 171.030 156.740 171.320 ;
        RECT 139.960 170.890 141.980 170.950 ;
        RECT 139.960 170.840 141.730 170.890 ;
        RECT 139.960 167.500 140.790 170.840 ;
        RECT 148.840 170.540 156.760 170.550 ;
        RECT 145.070 170.530 156.760 170.540 ;
        RECT 141.450 170.410 156.760 170.530 ;
        RECT 141.450 170.400 156.785 170.410 ;
        RECT 141.410 170.280 156.785 170.400 ;
        RECT 141.410 170.170 145.410 170.280 ;
        RECT 141.020 169.830 141.250 170.120 ;
        RECT 141.470 169.830 145.360 170.170 ;
        RECT 145.570 169.830 145.800 170.120 ;
        RECT 141.020 168.460 145.800 169.830 ;
        RECT 141.020 168.160 141.250 168.460 ;
        RECT 145.570 168.160 145.800 168.460 ;
        RECT 141.410 167.880 145.410 168.110 ;
        RECT 141.660 167.650 145.230 167.880 ;
        RECT 141.660 167.500 145.350 167.650 ;
        RECT 139.960 167.270 145.350 167.500 ;
        RECT 146.600 167.330 147.220 170.280 ;
        RECT 148.785 170.180 156.785 170.280 ;
        RECT 148.840 170.170 156.760 170.180 ;
        RECT 148.350 169.470 148.580 170.130 ;
        RECT 149.360 169.470 150.360 169.560 ;
        RECT 156.990 169.470 157.220 170.130 ;
        RECT 148.350 168.650 157.220 169.470 ;
        RECT 148.350 168.170 148.580 168.650 ;
        RECT 149.360 168.560 150.360 168.650 ;
        RECT 156.990 168.170 157.220 168.650 ;
        RECT 148.785 167.890 156.785 168.120 ;
        RECT 122.280 164.080 125.280 164.310 ;
        RECT 125.490 164.120 125.830 164.950 ;
        RECT 127.840 164.940 138.480 165.010 ;
        RECT 122.330 164.050 125.190 164.080 ;
        RECT 122.330 164.030 123.500 164.050 ;
        RECT 124.460 164.040 125.190 164.050 ;
        RECT 122.280 163.640 125.280 163.870 ;
        RECT 125.485 163.830 125.830 164.120 ;
        RECT 126.020 163.900 138.480 164.940 ;
        RECT 139.930 167.220 145.350 167.270 ;
        RECT 139.930 166.760 145.360 167.220 ;
        RECT 139.930 165.410 141.960 166.760 ;
        RECT 143.710 166.750 145.360 166.760 ;
        RECT 142.400 165.480 143.400 166.200 ;
        RECT 143.710 165.940 144.020 166.750 ;
        RECT 144.480 166.470 145.360 166.750 ;
        RECT 145.600 166.930 147.220 167.330 ;
        RECT 148.870 166.980 156.740 167.890 ;
        RECT 144.420 166.240 145.420 166.470 ;
        RECT 145.600 166.280 145.950 166.930 ;
        RECT 146.600 166.920 147.220 166.930 ;
        RECT 148.785 166.750 156.785 166.980 ;
        RECT 148.870 166.740 156.740 166.750 ;
        RECT 144.480 166.030 145.360 166.050 ;
        RECT 143.750 165.650 144.020 165.940 ;
        RECT 144.420 165.800 145.420 166.030 ;
        RECT 145.580 165.990 145.950 166.280 ;
        RECT 145.610 165.930 145.950 165.990 ;
        RECT 146.710 166.600 147.470 166.650 ;
        RECT 148.350 166.600 148.580 166.700 ;
        RECT 146.710 166.390 148.580 166.600 ;
        RECT 156.990 166.390 157.220 166.700 ;
        RECT 146.710 165.970 149.250 166.390 ;
        RECT 156.620 165.970 157.220 166.390 ;
        RECT 144.480 165.650 145.360 165.800 ;
        RECT 144.490 165.480 145.220 165.650 ;
        RECT 126.020 163.880 138.460 163.900 ;
        RECT 125.490 163.720 125.830 163.830 ;
        RECT 126.060 163.870 131.730 163.880 ;
        RECT 132.730 163.870 138.460 163.880 ;
        RECT 122.370 163.470 125.230 163.640 ;
        RECT 126.060 163.470 126.490 163.870 ;
        RECT 122.340 163.100 126.490 163.470 ;
        RECT 104.490 161.370 109.730 161.380 ;
        RECT 101.540 161.270 116.840 161.370 ;
        RECT 101.540 161.260 116.875 161.270 ;
        RECT 101.500 161.140 116.875 161.260 ;
        RECT 101.500 161.030 105.500 161.140 ;
        RECT 106.550 161.060 108.290 161.140 ;
        RECT 108.870 161.060 116.875 161.140 ;
        RECT 106.550 160.980 107.800 161.060 ;
        RECT 108.875 161.040 116.875 161.060 ;
        RECT 101.110 160.730 101.340 160.980 ;
        RECT 105.660 160.840 105.890 160.980 ;
        RECT 108.440 160.840 108.670 160.990 ;
        RECT 105.660 160.730 108.670 160.840 ;
        RECT 117.080 160.730 117.310 160.990 ;
        RECT 101.110 160.290 117.310 160.730 ;
        RECT 101.110 160.020 101.340 160.290 ;
        RECT 105.660 160.260 117.310 160.290 ;
        RECT 105.660 160.170 108.670 160.260 ;
        RECT 105.660 160.020 105.890 160.170 ;
        RECT 108.440 160.030 108.670 160.170 ;
        RECT 117.080 160.030 117.310 160.260 ;
        RECT 101.500 159.740 105.500 159.970 ;
        RECT 108.875 159.760 116.875 159.980 ;
        RECT 117.640 159.760 118.600 161.800 ;
        RECT 108.875 159.750 118.600 159.760 ;
        RECT 101.500 159.670 105.490 159.740 ;
        RECT 38.850 159.480 39.170 159.540 ;
        RECT 33.880 159.340 38.160 159.480 ;
        RECT 33.880 159.185 34.020 159.340 ;
        RECT 33.805 158.955 34.095 159.185 ;
        RECT 34.725 158.955 35.015 159.185 ;
        RECT 34.800 158.800 34.940 158.955 ;
        RECT 36.090 158.940 36.410 159.200 ;
        RECT 37.470 158.940 37.790 159.200 ;
        RECT 37.010 158.800 37.330 158.860 ;
        RECT 34.800 158.660 37.330 158.800 ;
        RECT 38.020 158.800 38.160 159.340 ;
        RECT 38.480 159.340 39.170 159.480 ;
        RECT 38.480 159.185 38.620 159.340 ;
        RECT 38.850 159.280 39.170 159.340 ;
        RECT 39.740 159.480 40.030 159.525 ;
        RECT 40.780 159.480 40.920 159.620 ;
        RECT 100.010 159.560 105.490 159.670 ;
        RECT 108.930 159.590 118.600 159.750 ;
        RECT 39.740 159.340 40.920 159.480 ;
        RECT 46.670 159.480 46.990 159.540 ;
        RECT 47.450 159.480 47.740 159.525 ;
        RECT 46.670 159.340 47.740 159.480 ;
        RECT 39.740 159.295 40.030 159.340 ;
        RECT 46.670 159.280 46.990 159.340 ;
        RECT 47.450 159.295 47.740 159.340 ;
        RECT 53.585 159.480 53.875 159.525 ;
        RECT 57.250 159.480 57.570 159.540 ;
        RECT 53.585 159.340 57.570 159.480 ;
        RECT 53.585 159.295 53.875 159.340 ;
        RECT 57.250 159.280 57.570 159.340 ;
        RECT 58.185 159.480 58.475 159.525 ;
        RECT 60.470 159.480 60.790 159.540 ;
        RECT 58.185 159.340 60.790 159.480 ;
        RECT 58.185 159.295 58.475 159.340 ;
        RECT 60.470 159.280 60.790 159.340 ;
        RECT 70.590 159.480 70.910 159.540 ;
        RECT 74.270 159.480 74.590 159.540 ;
        RECT 76.125 159.480 76.415 159.525 ;
        RECT 70.590 159.340 71.740 159.480 ;
        RECT 70.590 159.280 70.910 159.340 ;
        RECT 38.405 158.955 38.695 159.185 ;
        RECT 43.910 159.140 44.230 159.200 ;
        RECT 46.210 159.140 46.530 159.200 ;
        RECT 38.940 159.000 43.680 159.140 ;
        RECT 38.940 158.800 39.080 159.000 ;
        RECT 38.020 158.660 39.080 158.800 ;
        RECT 39.285 158.800 39.575 158.845 ;
        RECT 40.475 158.800 40.765 158.845 ;
        RECT 42.995 158.800 43.285 158.845 ;
        RECT 39.285 158.660 43.285 158.800 ;
        RECT 43.540 158.800 43.680 159.000 ;
        RECT 43.910 159.000 46.530 159.140 ;
        RECT 43.910 158.940 44.230 159.000 ;
        RECT 46.210 158.940 46.530 159.000 ;
        RECT 55.885 159.140 56.175 159.185 ;
        RECT 56.790 159.140 57.110 159.200 ;
        RECT 55.885 159.000 57.110 159.140 ;
        RECT 55.885 158.955 56.175 159.000 ;
        RECT 56.790 158.940 57.110 159.000 ;
        RECT 59.550 159.140 59.870 159.200 ;
        RECT 71.600 159.140 71.740 159.340 ;
        RECT 74.270 159.340 76.415 159.480 ;
        RECT 74.270 159.280 74.590 159.340 ;
        RECT 76.125 159.295 76.415 159.340 ;
        RECT 100.010 159.470 103.180 159.560 ;
        RECT 116.670 159.540 118.600 159.590 ;
        RECT 75.205 159.140 75.495 159.185 ;
        RECT 59.550 159.000 71.280 159.140 ;
        RECT 71.600 159.000 75.495 159.140 ;
        RECT 59.550 158.940 59.870 159.000 ;
        RECT 47.105 158.800 47.395 158.845 ;
        RECT 48.295 158.800 48.585 158.845 ;
        RECT 50.815 158.800 51.105 158.845 ;
        RECT 43.540 158.660 45.980 158.800 ;
        RECT 37.010 158.600 37.330 158.660 ;
        RECT 39.285 158.615 39.575 158.660 ;
        RECT 40.475 158.615 40.765 158.660 ;
        RECT 42.995 158.615 43.285 158.660 ;
        RECT 38.890 158.460 39.180 158.505 ;
        RECT 40.990 158.460 41.280 158.505 ;
        RECT 42.560 158.460 42.850 158.505 ;
        RECT 38.890 158.320 42.850 158.460 ;
        RECT 38.890 158.275 39.180 158.320 ;
        RECT 40.990 158.275 41.280 158.320 ;
        RECT 42.560 158.275 42.850 158.320 ;
        RECT 34.250 157.920 34.570 158.180 ;
        RECT 35.185 158.120 35.475 158.165 ;
        RECT 41.610 158.120 41.930 158.180 ;
        RECT 35.185 157.980 41.930 158.120 ;
        RECT 35.185 157.935 35.475 157.980 ;
        RECT 41.610 157.920 41.930 157.980 ;
        RECT 45.290 157.920 45.610 158.180 ;
        RECT 45.840 158.120 45.980 158.660 ;
        RECT 47.105 158.660 51.105 158.800 ;
        RECT 47.105 158.615 47.395 158.660 ;
        RECT 48.295 158.615 48.585 158.660 ;
        RECT 50.815 158.615 51.105 158.660 ;
        RECT 55.425 158.800 55.715 158.845 ;
        RECT 60.485 158.800 60.775 158.845 ;
        RECT 62.785 158.800 63.075 158.845 ;
        RECT 55.425 158.660 60.775 158.800 ;
        RECT 55.425 158.615 55.715 158.660 ;
        RECT 60.485 158.615 60.775 158.660 ;
        RECT 61.020 158.660 63.075 158.800 ;
        RECT 46.710 158.460 47.000 158.505 ;
        RECT 48.810 158.460 49.100 158.505 ;
        RECT 50.380 158.460 50.670 158.505 ;
        RECT 57.265 158.460 57.555 158.505 ;
        RECT 46.710 158.320 50.670 158.460 ;
        RECT 46.710 158.275 47.000 158.320 ;
        RECT 48.810 158.275 49.100 158.320 ;
        RECT 50.380 158.275 50.670 158.320 ;
        RECT 55.500 158.320 57.555 158.460 ;
        RECT 50.810 158.120 51.130 158.180 ;
        RECT 55.500 158.165 55.640 158.320 ;
        RECT 57.265 158.275 57.555 158.320 ;
        RECT 60.010 158.260 60.330 158.520 ;
        RECT 45.840 157.980 51.130 158.120 ;
        RECT 50.810 157.920 51.130 157.980 ;
        RECT 55.425 157.935 55.715 158.165 ;
        RECT 55.870 158.120 56.190 158.180 ;
        RECT 56.805 158.120 57.095 158.165 ;
        RECT 55.870 157.980 57.095 158.120 ;
        RECT 55.870 157.920 56.190 157.980 ;
        RECT 56.805 157.935 57.095 157.980 ;
        RECT 58.170 158.120 58.490 158.180 ;
        RECT 61.020 158.120 61.160 158.660 ;
        RECT 62.785 158.615 63.075 158.660 ;
        RECT 63.230 158.800 63.550 158.860 ;
        RECT 66.465 158.800 66.755 158.845 ;
        RECT 63.230 158.660 66.755 158.800 ;
        RECT 63.230 158.600 63.550 158.660 ;
        RECT 66.465 158.615 66.755 158.660 ;
        RECT 66.925 158.800 67.215 158.845 ;
        RECT 70.130 158.800 70.450 158.860 ;
        RECT 66.925 158.660 70.450 158.800 ;
        RECT 66.925 158.615 67.215 158.660 ;
        RECT 61.390 158.260 61.710 158.520 ;
        RECT 61.850 158.460 62.170 158.520 ;
        RECT 67.000 158.460 67.140 158.615 ;
        RECT 70.130 158.600 70.450 158.660 ;
        RECT 70.605 158.615 70.895 158.845 ;
        RECT 61.850 158.320 67.140 158.460 ;
        RECT 68.290 158.460 68.610 158.520 ;
        RECT 70.680 158.460 70.820 158.615 ;
        RECT 68.290 158.320 70.820 158.460 ;
        RECT 71.140 158.460 71.280 159.000 ;
        RECT 75.205 158.955 75.495 159.000 ;
        RECT 77.030 159.140 77.350 159.200 ;
        RECT 77.505 159.140 77.795 159.185 ;
        RECT 77.030 159.000 77.795 159.140 ;
        RECT 77.030 158.940 77.350 159.000 ;
        RECT 77.505 158.955 77.795 159.000 ;
        RECT 77.950 158.940 78.270 159.200 ;
        RECT 78.425 158.955 78.715 159.185 ;
        RECT 71.525 158.800 71.815 158.845 ;
        RECT 71.970 158.800 72.290 158.860 ;
        RECT 71.525 158.660 72.290 158.800 ;
        RECT 71.525 158.615 71.815 158.660 ;
        RECT 71.970 158.600 72.290 158.660 ;
        RECT 72.430 158.800 72.750 158.860 ;
        RECT 78.500 158.800 78.640 158.955 ;
        RECT 79.330 158.940 79.650 159.200 ;
        RECT 80.725 158.955 81.015 159.185 ;
        RECT 72.430 158.660 78.640 158.800 ;
        RECT 78.870 158.800 79.190 158.860 ;
        RECT 80.800 158.800 80.940 158.955 ;
        RECT 81.170 158.940 81.490 159.200 ;
        RECT 81.630 158.940 81.950 159.200 ;
        RECT 82.520 159.140 82.810 159.185 ;
        RECT 84.390 159.140 84.710 159.200 ;
        RECT 82.520 159.000 84.710 159.140 ;
        RECT 82.520 158.955 82.810 159.000 ;
        RECT 84.390 158.940 84.710 159.000 ;
        RECT 81.720 158.800 81.860 158.940 ;
        RECT 78.870 158.660 80.940 158.800 ;
        RECT 81.260 158.660 81.860 158.800 ;
        RECT 82.065 158.800 82.355 158.845 ;
        RECT 83.255 158.800 83.545 158.845 ;
        RECT 85.775 158.800 86.065 158.845 ;
        RECT 82.065 158.660 86.065 158.800 ;
        RECT 72.430 158.600 72.750 158.660 ;
        RECT 78.870 158.600 79.190 158.660 ;
        RECT 79.805 158.460 80.095 158.505 ;
        RECT 71.140 158.320 80.095 158.460 ;
        RECT 61.850 158.260 62.170 158.320 ;
        RECT 68.290 158.260 68.610 158.320 ;
        RECT 79.805 158.275 80.095 158.320 ;
        RECT 58.170 157.980 61.160 158.120 ;
        RECT 67.370 158.120 67.690 158.180 ;
        RECT 72.445 158.120 72.735 158.165 ;
        RECT 67.370 157.980 72.735 158.120 ;
        RECT 58.170 157.920 58.490 157.980 ;
        RECT 67.370 157.920 67.690 157.980 ;
        RECT 72.445 157.935 72.735 157.980 ;
        RECT 77.030 158.120 77.350 158.180 ;
        RECT 81.260 158.120 81.400 158.660 ;
        RECT 82.065 158.615 82.355 158.660 ;
        RECT 83.255 158.615 83.545 158.660 ;
        RECT 85.775 158.615 86.065 158.660 ;
        RECT 81.670 158.460 81.960 158.505 ;
        RECT 83.770 158.460 84.060 158.505 ;
        RECT 85.340 158.460 85.630 158.505 ;
        RECT 81.670 158.320 85.630 158.460 ;
        RECT 81.670 158.275 81.960 158.320 ;
        RECT 83.770 158.275 84.060 158.320 ;
        RECT 85.340 158.275 85.630 158.320 ;
        RECT 85.770 158.120 86.090 158.180 ;
        RECT 77.030 157.980 86.090 158.120 ;
        RECT 77.030 157.920 77.350 157.980 ;
        RECT 85.770 157.920 86.090 157.980 ;
        RECT 12.100 157.300 89.840 157.780 ;
        RECT 37.010 156.900 37.330 157.160 ;
        RECT 42.070 157.100 42.390 157.160 ;
        RECT 43.450 157.100 43.770 157.160 ;
        RECT 45.750 157.100 46.070 157.160 ;
        RECT 42.070 156.960 46.070 157.100 ;
        RECT 42.070 156.900 42.390 156.960 ;
        RECT 43.450 156.900 43.770 156.960 ;
        RECT 45.750 156.900 46.070 156.960 ;
        RECT 52.665 157.100 52.955 157.145 ;
        RECT 54.030 157.100 54.350 157.160 ;
        RECT 52.665 156.960 54.350 157.100 ;
        RECT 52.665 156.915 52.955 156.960 ;
        RECT 54.030 156.900 54.350 156.960 ;
        RECT 56.330 156.900 56.650 157.160 ;
        RECT 57.265 157.100 57.555 157.145 ;
        RECT 58.170 157.100 58.490 157.160 ;
        RECT 57.265 156.960 58.490 157.100 ;
        RECT 57.265 156.915 57.555 156.960 ;
        RECT 39.785 156.760 40.075 156.805 ;
        RECT 42.530 156.760 42.850 156.820 ;
        RECT 36.180 156.620 42.850 156.760 ;
        RECT 36.180 156.080 36.320 156.620 ;
        RECT 39.785 156.575 40.075 156.620 ;
        RECT 42.530 156.560 42.850 156.620 ;
        RECT 54.490 156.760 54.810 156.820 ;
        RECT 57.340 156.760 57.480 156.915 ;
        RECT 58.170 156.900 58.490 156.960 ;
        RECT 58.630 157.100 58.950 157.160 ;
        RECT 59.565 157.100 59.855 157.145 ;
        RECT 71.510 157.100 71.830 157.160 ;
        RECT 77.030 157.100 77.350 157.160 ;
        RECT 58.630 156.960 59.855 157.100 ;
        RECT 58.630 156.900 58.950 156.960 ;
        RECT 59.565 156.915 59.855 156.960 ;
        RECT 63.320 156.960 77.350 157.100 ;
        RECT 60.485 156.760 60.775 156.805 ;
        RECT 62.770 156.760 63.090 156.820 ;
        RECT 54.490 156.620 57.940 156.760 ;
        RECT 54.490 156.560 54.810 156.620 ;
        RECT 36.565 156.420 36.855 156.465 ;
        RECT 45.290 156.420 45.610 156.480 ;
        RECT 45.765 156.420 46.055 156.465 ;
        RECT 36.565 156.280 46.055 156.420 ;
        RECT 36.565 156.235 36.855 156.280 ;
        RECT 45.290 156.220 45.610 156.280 ;
        RECT 45.765 156.235 46.055 156.280 ;
        RECT 47.130 156.420 47.450 156.480 ;
        RECT 56.330 156.420 56.650 156.480 ;
        RECT 57.250 156.420 57.570 156.480 ;
        RECT 47.130 156.280 57.570 156.420 ;
        RECT 57.800 156.420 57.940 156.620 ;
        RECT 60.485 156.620 63.090 156.760 ;
        RECT 60.485 156.575 60.775 156.620 ;
        RECT 62.770 156.560 63.090 156.620 ;
        RECT 61.865 156.420 62.155 156.465 ;
        RECT 62.310 156.420 62.630 156.480 ;
        RECT 57.800 156.280 62.630 156.420 ;
        RECT 47.130 156.220 47.450 156.280 ;
        RECT 56.330 156.220 56.650 156.280 ;
        RECT 57.250 156.220 57.570 156.280 ;
        RECT 61.865 156.235 62.155 156.280 ;
        RECT 62.310 156.220 62.630 156.280 ;
        RECT 37.025 156.080 37.315 156.125 ;
        RECT 36.180 155.940 37.315 156.080 ;
        RECT 37.025 155.895 37.315 155.940 ;
        RECT 37.470 156.080 37.790 156.140 ;
        RECT 37.470 155.940 39.080 156.080 ;
        RECT 37.470 155.880 37.790 155.940 ;
        RECT 38.405 155.555 38.695 155.785 ;
        RECT 38.940 155.740 39.080 155.940 ;
        RECT 41.150 155.880 41.470 156.140 ;
        RECT 42.545 156.130 42.835 156.135 ;
        RECT 42.545 155.990 43.680 156.130 ;
        RECT 42.545 155.905 42.835 155.990 ;
        RECT 42.070 155.740 42.390 155.800 ;
        RECT 38.940 155.600 42.390 155.740 ;
        RECT 43.540 155.740 43.680 155.990 ;
        RECT 50.810 156.080 51.130 156.140 ;
        RECT 51.285 156.080 51.575 156.125 ;
        RECT 50.810 155.940 51.575 156.080 ;
        RECT 50.810 155.880 51.130 155.940 ;
        RECT 51.285 155.895 51.575 155.940 ;
        RECT 52.205 156.080 52.495 156.125 ;
        RECT 52.650 156.080 52.970 156.140 ;
        RECT 52.205 155.940 52.970 156.080 ;
        RECT 52.205 155.895 52.495 155.940 ;
        RECT 52.280 155.740 52.420 155.895 ;
        RECT 52.650 155.880 52.970 155.940 ;
        RECT 53.570 156.080 53.890 156.140 ;
        RECT 54.045 156.080 54.335 156.125 ;
        RECT 53.570 155.940 54.335 156.080 ;
        RECT 53.570 155.880 53.890 155.940 ;
        RECT 54.045 155.895 54.335 155.940 ;
        RECT 43.540 155.600 52.420 155.740 ;
        RECT 54.120 155.740 54.260 155.895 ;
        RECT 54.490 155.880 54.810 156.140 ;
        RECT 54.965 156.080 55.255 156.125 ;
        RECT 55.410 156.080 55.730 156.140 ;
        RECT 54.965 155.940 55.730 156.080 ;
        RECT 54.965 155.895 55.255 155.940 ;
        RECT 55.410 155.880 55.730 155.940 ;
        RECT 55.870 155.880 56.190 156.140 ;
        RECT 59.105 156.080 59.395 156.125 ;
        RECT 60.010 156.080 60.330 156.140 ;
        RECT 63.320 156.125 63.460 156.960 ;
        RECT 71.510 156.900 71.830 156.960 ;
        RECT 77.030 156.900 77.350 156.960 ;
        RECT 80.710 156.900 81.030 157.160 ;
        RECT 84.390 156.900 84.710 157.160 ;
        RECT 65.530 156.560 65.850 156.820 ;
        RECT 67.830 156.760 68.150 156.820 ;
        RECT 67.830 156.620 86.920 156.760 ;
        RECT 67.830 156.560 68.150 156.620 ;
        RECT 68.290 156.420 68.610 156.480 ;
        RECT 65.620 156.280 68.610 156.420 ;
        RECT 59.105 155.940 60.330 156.080 ;
        RECT 59.105 155.895 59.395 155.940 ;
        RECT 59.180 155.740 59.320 155.895 ;
        RECT 60.010 155.880 60.330 155.940 ;
        RECT 63.245 155.895 63.535 156.125 ;
        RECT 63.690 155.880 64.010 156.140 ;
        RECT 64.610 155.880 64.930 156.140 ;
        RECT 65.070 155.880 65.390 156.140 ;
        RECT 54.120 155.600 59.320 155.740 ;
        RECT 62.325 155.740 62.615 155.785 ;
        RECT 65.620 155.740 65.760 156.280 ;
        RECT 68.290 156.220 68.610 156.280 ;
        RECT 68.765 156.420 69.055 156.465 ;
        RECT 70.130 156.420 70.450 156.480 ;
        RECT 71.970 156.420 72.290 156.480 ;
        RECT 72.445 156.420 72.735 156.465 ;
        RECT 68.765 156.280 72.735 156.420 ;
        RECT 68.765 156.235 69.055 156.280 ;
        RECT 70.130 156.220 70.450 156.280 ;
        RECT 71.970 156.220 72.290 156.280 ;
        RECT 72.445 156.235 72.735 156.280 ;
        RECT 72.890 156.420 73.210 156.480 ;
        RECT 78.410 156.420 78.730 156.480 ;
        RECT 84.850 156.420 85.170 156.480 ;
        RECT 72.890 156.280 82.320 156.420 ;
        RECT 72.890 156.220 73.210 156.280 ;
        RECT 78.410 156.220 78.730 156.280 ;
        RECT 67.370 155.880 67.690 156.140 ;
        RECT 71.525 156.080 71.815 156.125 ;
        RECT 77.045 156.080 77.335 156.125 ;
        RECT 71.525 155.940 77.335 156.080 ;
        RECT 71.525 155.895 71.815 155.940 ;
        RECT 77.045 155.895 77.335 155.940 ;
        RECT 80.265 156.080 80.555 156.125 ;
        RECT 80.710 156.080 81.030 156.140 ;
        RECT 82.180 156.125 82.320 156.280 ;
        RECT 82.640 156.280 86.460 156.420 ;
        RECT 82.640 156.125 82.780 156.280 ;
        RECT 84.850 156.220 85.170 156.280 ;
        RECT 80.265 155.940 81.030 156.080 ;
        RECT 80.265 155.895 80.555 155.940 ;
        RECT 62.325 155.600 65.760 155.740 ;
        RECT 67.845 155.740 68.135 155.785 ;
        RECT 73.810 155.740 74.130 155.800 ;
        RECT 67.845 155.600 74.130 155.740 ;
        RECT 35.170 155.200 35.490 155.460 ;
        RECT 37.010 155.400 37.330 155.460 ;
        RECT 38.480 155.400 38.620 155.555 ;
        RECT 42.070 155.540 42.390 155.600 ;
        RECT 62.325 155.555 62.615 155.600 ;
        RECT 67.845 155.555 68.135 155.600 ;
        RECT 73.810 155.540 74.130 155.600 ;
        RECT 74.270 155.540 74.590 155.800 ;
        RECT 75.190 155.540 75.510 155.800 ;
        RECT 80.340 155.740 80.480 155.895 ;
        RECT 80.710 155.880 81.030 155.940 ;
        RECT 82.105 155.895 82.395 156.125 ;
        RECT 82.565 155.895 82.855 156.125 ;
        RECT 83.010 155.880 83.330 156.140 ;
        RECT 83.945 156.080 84.235 156.125 ;
        RECT 83.560 155.940 84.235 156.080 ;
        RECT 75.740 155.600 80.480 155.740 ;
        RECT 83.560 155.740 83.700 155.940 ;
        RECT 83.945 155.895 84.235 155.940 ;
        RECT 85.770 155.880 86.090 156.140 ;
        RECT 86.320 156.125 86.460 156.280 ;
        RECT 86.780 156.125 86.920 156.620 ;
        RECT 100.010 156.200 100.880 159.470 ;
        RECT 104.530 159.010 109.780 159.020 ;
        RECT 104.530 158.900 116.840 159.010 ;
        RECT 101.560 158.840 116.840 158.900 ;
        RECT 101.560 158.830 116.875 158.840 ;
        RECT 101.500 158.700 116.875 158.830 ;
        RECT 101.500 158.690 106.660 158.700 ;
        RECT 101.500 158.600 105.500 158.690 ;
        RECT 108.875 158.610 116.875 158.700 ;
        RECT 108.960 158.600 116.850 158.610 ;
        RECT 101.110 158.240 101.340 158.550 ;
        RECT 101.560 158.240 105.460 158.600 ;
        RECT 105.660 158.240 105.890 158.550 ;
        RECT 101.110 156.900 105.890 158.240 ;
        RECT 101.110 156.590 101.340 156.900 ;
        RECT 105.660 156.590 105.890 156.900 ;
        RECT 108.440 158.020 108.670 158.560 ;
        RECT 109.480 158.020 110.490 158.050 ;
        RECT 117.080 158.020 117.310 158.560 ;
        RECT 108.440 157.120 117.310 158.020 ;
        RECT 108.440 156.600 108.670 157.120 ;
        RECT 109.480 157.050 110.490 157.120 ;
        RECT 117.080 156.600 117.310 157.120 ;
        RECT 101.500 156.310 105.500 156.540 ;
        RECT 108.875 156.320 116.875 156.550 ;
        RECT 100.010 156.160 101.180 156.200 ;
        RECT 86.245 155.895 86.535 156.125 ;
        RECT 86.705 155.895 86.995 156.125 ;
        RECT 87.625 155.895 87.915 156.125 ;
        RECT 100.010 156.080 101.420 156.160 ;
        RECT 101.790 156.090 105.450 156.310 ;
        RECT 101.790 156.080 103.230 156.090 ;
        RECT 100.010 156.040 103.230 156.080 ;
        RECT 100.010 155.950 102.740 156.040 ;
        RECT 108.940 156.030 116.830 156.320 ;
        RECT 87.700 155.740 87.840 155.895 ;
        RECT 83.560 155.600 87.840 155.740 ;
        RECT 100.010 155.890 102.070 155.950 ;
        RECT 100.010 155.840 101.820 155.890 ;
        RECT 37.010 155.260 38.620 155.400 ;
        RECT 39.325 155.400 39.615 155.445 ;
        RECT 40.230 155.400 40.550 155.460 ;
        RECT 39.325 155.260 40.550 155.400 ;
        RECT 37.010 155.200 37.330 155.260 ;
        RECT 39.325 155.215 39.615 155.260 ;
        RECT 40.230 155.200 40.550 155.260 ;
        RECT 41.150 155.400 41.470 155.460 ;
        RECT 43.005 155.400 43.295 155.445 ;
        RECT 41.150 155.260 43.295 155.400 ;
        RECT 41.150 155.200 41.470 155.260 ;
        RECT 43.005 155.215 43.295 155.260 ;
        RECT 49.890 155.200 50.210 155.460 ;
        RECT 51.730 155.200 52.050 155.460 ;
        RECT 57.265 155.400 57.555 155.445 ;
        RECT 58.170 155.400 58.490 155.460 ;
        RECT 57.265 155.260 58.490 155.400 ;
        RECT 57.265 155.215 57.555 155.260 ;
        RECT 58.170 155.200 58.490 155.260 ;
        RECT 59.090 155.400 59.410 155.460 ;
        RECT 69.210 155.400 69.530 155.460 ;
        RECT 59.090 155.260 69.530 155.400 ;
        RECT 59.090 155.200 59.410 155.260 ;
        RECT 69.210 155.200 69.530 155.260 ;
        RECT 69.670 155.200 69.990 155.460 ;
        RECT 71.050 155.400 71.370 155.460 ;
        RECT 71.985 155.400 72.275 155.445 ;
        RECT 72.890 155.400 73.210 155.460 ;
        RECT 71.050 155.260 73.210 155.400 ;
        RECT 71.050 155.200 71.370 155.260 ;
        RECT 71.985 155.215 72.275 155.260 ;
        RECT 72.890 155.200 73.210 155.260 ;
        RECT 74.730 155.400 75.050 155.460 ;
        RECT 75.740 155.400 75.880 155.600 ;
        RECT 74.730 155.260 75.880 155.400 ;
        RECT 76.125 155.400 76.415 155.445 ;
        RECT 77.950 155.400 78.270 155.460 ;
        RECT 76.125 155.260 78.270 155.400 ;
        RECT 74.730 155.200 75.050 155.260 ;
        RECT 76.125 155.215 76.415 155.260 ;
        RECT 77.950 155.200 78.270 155.260 ;
        RECT 79.330 155.400 79.650 155.460 ;
        RECT 83.560 155.400 83.700 155.600 ;
        RECT 79.330 155.260 83.700 155.400 ;
        RECT 79.330 155.200 79.650 155.260 ;
        RECT 12.100 154.580 89.840 155.060 ;
        RECT 39.325 154.380 39.615 154.425 ;
        RECT 39.770 154.380 40.090 154.440 ;
        RECT 39.325 154.240 40.090 154.380 ;
        RECT 39.325 154.195 39.615 154.240 ;
        RECT 39.770 154.180 40.090 154.240 ;
        RECT 40.230 154.380 40.550 154.440 ;
        RECT 48.510 154.380 48.830 154.440 ;
        RECT 40.230 154.240 48.830 154.380 ;
        RECT 40.230 154.180 40.550 154.240 ;
        RECT 48.510 154.180 48.830 154.240 ;
        RECT 49.890 154.380 50.210 154.440 ;
        RECT 52.205 154.380 52.495 154.425 ;
        RECT 49.890 154.240 52.495 154.380 ;
        RECT 49.890 154.180 50.210 154.240 ;
        RECT 52.205 154.195 52.495 154.240 ;
        RECT 60.930 154.380 61.250 154.440 ;
        RECT 61.405 154.380 61.695 154.425 ;
        RECT 60.930 154.240 61.695 154.380 ;
        RECT 60.930 154.180 61.250 154.240 ;
        RECT 61.405 154.195 61.695 154.240 ;
        RECT 62.245 154.380 62.535 154.425 ;
        RECT 64.610 154.380 64.930 154.440 ;
        RECT 62.245 154.240 64.930 154.380 ;
        RECT 62.245 154.195 62.535 154.240 ;
        RECT 64.610 154.180 64.930 154.240 ;
        RECT 74.730 154.180 75.050 154.440 ;
        RECT 77.030 154.380 77.350 154.440 ;
        RECT 79.790 154.380 80.110 154.440 ;
        RECT 86.230 154.380 86.550 154.440 ;
        RECT 87.165 154.380 87.455 154.425 ;
        RECT 77.030 154.240 85.080 154.380 ;
        RECT 77.030 154.180 77.350 154.240 ;
        RECT 79.790 154.180 80.110 154.240 ;
        RECT 36.090 154.040 36.410 154.100 ;
        RECT 40.690 154.040 41.010 154.100 ;
        RECT 46.210 154.040 46.530 154.100 ;
        RECT 51.730 154.040 52.050 154.100 ;
        RECT 60.010 154.040 60.330 154.100 ;
        RECT 63.245 154.040 63.535 154.085 ;
        RECT 36.090 153.900 41.840 154.040 ;
        RECT 36.090 153.840 36.410 153.900 ;
        RECT 40.690 153.840 41.010 153.900 ;
        RECT 34.250 153.700 34.570 153.760 ;
        RECT 39.770 153.700 40.090 153.760 ;
        RECT 34.250 153.560 40.920 153.700 ;
        RECT 34.250 153.500 34.570 153.560 ;
        RECT 39.770 153.500 40.090 153.560 ;
        RECT 40.780 153.405 40.920 153.560 ;
        RECT 41.150 153.500 41.470 153.760 ;
        RECT 41.700 153.745 41.840 153.900 ;
        RECT 46.210 153.900 50.120 154.040 ;
        RECT 46.210 153.840 46.530 153.900 ;
        RECT 49.980 153.745 50.120 153.900 ;
        RECT 51.730 153.900 52.880 154.040 ;
        RECT 51.730 153.840 52.050 153.900 ;
        RECT 41.625 153.515 41.915 153.745 ;
        RECT 48.625 153.700 48.915 153.745 ;
        RECT 48.625 153.560 49.660 153.700 ;
        RECT 48.625 153.515 48.915 153.560 ;
        RECT 40.245 153.175 40.535 153.405 ;
        RECT 40.705 153.175 40.995 153.405 ;
        RECT 45.315 153.360 45.605 153.405 ;
        RECT 47.835 153.360 48.125 153.405 ;
        RECT 49.025 153.360 49.315 153.405 ;
        RECT 45.315 153.220 49.315 153.360 ;
        RECT 49.520 153.360 49.660 153.560 ;
        RECT 49.905 153.515 50.195 153.745 ;
        RECT 51.270 153.500 51.590 153.760 ;
        RECT 52.740 153.745 52.880 153.900 ;
        RECT 60.010 153.900 63.535 154.040 ;
        RECT 60.010 153.840 60.330 153.900 ;
        RECT 63.245 153.855 63.535 153.900 ;
        RECT 69.180 154.040 69.470 154.085 ;
        RECT 69.670 154.040 69.990 154.100 ;
        RECT 69.180 153.900 69.990 154.040 ;
        RECT 69.180 153.855 69.470 153.900 ;
        RECT 69.670 153.840 69.990 153.900 ;
        RECT 73.350 154.040 73.670 154.100 ;
        RECT 83.930 154.040 84.250 154.100 ;
        RECT 73.350 153.900 80.480 154.040 ;
        RECT 73.350 153.840 73.670 153.900 ;
        RECT 52.665 153.515 52.955 153.745 ;
        RECT 54.045 153.700 54.335 153.745 ;
        RECT 54.490 153.700 54.810 153.760 ;
        RECT 54.045 153.560 54.810 153.700 ;
        RECT 54.045 153.515 54.335 153.560 ;
        RECT 54.490 153.500 54.810 153.560 ;
        RECT 55.380 153.700 55.670 153.745 ;
        RECT 57.250 153.700 57.570 153.760 ;
        RECT 55.380 153.560 57.570 153.700 ;
        RECT 55.380 153.515 55.670 153.560 ;
        RECT 57.250 153.500 57.570 153.560 ;
        RECT 78.425 153.700 78.715 153.745 ;
        RECT 78.870 153.700 79.190 153.760 ;
        RECT 78.425 153.560 79.190 153.700 ;
        RECT 78.425 153.515 78.715 153.560 ;
        RECT 78.870 153.500 79.190 153.560 ;
        RECT 79.790 153.500 80.110 153.760 ;
        RECT 80.340 153.745 80.480 153.900 ;
        RECT 81.260 153.900 84.250 154.040 ;
        RECT 81.260 153.745 81.400 153.900 ;
        RECT 83.930 153.840 84.250 153.900 ;
        RECT 80.265 153.515 80.555 153.745 ;
        RECT 81.185 153.515 81.475 153.745 ;
        RECT 81.630 153.500 81.950 153.760 ;
        RECT 82.105 153.720 82.395 153.745 ;
        RECT 83.010 153.720 83.330 153.760 ;
        RECT 84.940 153.745 85.080 154.240 ;
        RECT 86.230 154.240 87.455 154.380 ;
        RECT 86.230 154.180 86.550 154.240 ;
        RECT 87.165 154.195 87.455 154.240 ;
        RECT 82.105 153.580 83.330 153.720 ;
        RECT 82.105 153.515 82.395 153.580 ;
        RECT 83.010 153.500 83.330 153.580 ;
        RECT 84.865 153.515 85.155 153.745 ;
        RECT 85.325 153.515 85.615 153.745 ;
        RECT 50.365 153.360 50.655 153.405 ;
        RECT 49.520 153.220 50.655 153.360 ;
        RECT 45.315 153.175 45.605 153.220 ;
        RECT 47.835 153.175 48.125 153.220 ;
        RECT 49.025 153.175 49.315 153.220 ;
        RECT 50.365 153.175 50.655 153.220 ;
        RECT 54.925 153.360 55.215 153.405 ;
        RECT 56.115 153.360 56.405 153.405 ;
        RECT 58.635 153.360 58.925 153.405 ;
        RECT 54.925 153.220 58.925 153.360 ;
        RECT 54.925 153.175 55.215 153.220 ;
        RECT 56.115 153.175 56.405 153.220 ;
        RECT 58.635 153.175 58.925 153.220 ;
        RECT 66.925 153.175 67.215 153.405 ;
        RECT 40.320 153.020 40.460 153.175 ;
        RECT 42.530 153.020 42.850 153.080 ;
        RECT 40.320 152.880 42.850 153.020 ;
        RECT 42.530 152.820 42.850 152.880 ;
        RECT 42.990 152.820 43.310 153.080 ;
        RECT 45.750 153.020 46.040 153.065 ;
        RECT 47.320 153.020 47.610 153.065 ;
        RECT 49.420 153.020 49.710 153.065 ;
        RECT 45.750 152.880 49.710 153.020 ;
        RECT 45.750 152.835 46.040 152.880 ;
        RECT 47.320 152.835 47.610 152.880 ;
        RECT 49.420 152.835 49.710 152.880 ;
        RECT 54.530 153.020 54.820 153.065 ;
        RECT 56.630 153.020 56.920 153.065 ;
        RECT 58.200 153.020 58.490 153.065 ;
        RECT 54.530 152.880 58.490 153.020 ;
        RECT 54.530 152.835 54.820 152.880 ;
        RECT 56.630 152.835 56.920 152.880 ;
        RECT 58.200 152.835 58.490 152.880 ;
        RECT 60.470 153.020 60.790 153.080 ;
        RECT 60.945 153.020 61.235 153.065 ;
        RECT 67.000 153.020 67.140 153.175 ;
        RECT 67.830 153.160 68.150 153.420 ;
        RECT 68.725 153.360 69.015 153.405 ;
        RECT 69.915 153.360 70.205 153.405 ;
        RECT 72.435 153.360 72.725 153.405 ;
        RECT 68.725 153.220 72.725 153.360 ;
        RECT 68.725 153.175 69.015 153.220 ;
        RECT 69.915 153.175 70.205 153.220 ;
        RECT 72.435 153.175 72.725 153.220 ;
        RECT 75.190 153.360 75.510 153.420 ;
        RECT 83.930 153.360 84.250 153.420 ;
        RECT 85.400 153.360 85.540 153.515 ;
        RECT 86.230 153.500 86.550 153.760 ;
        RECT 86.690 153.500 87.010 153.760 ;
        RECT 88.070 153.500 88.390 153.760 ;
        RECT 75.190 153.220 85.540 153.360 ;
        RECT 75.190 153.160 75.510 153.220 ;
        RECT 83.930 153.160 84.250 153.220 ;
        RECT 60.470 152.880 67.140 153.020 ;
        RECT 68.330 153.020 68.620 153.065 ;
        RECT 70.430 153.020 70.720 153.065 ;
        RECT 72.000 153.020 72.290 153.065 ;
        RECT 68.330 152.880 72.290 153.020 ;
        RECT 60.470 152.820 60.790 152.880 ;
        RECT 60.945 152.835 61.235 152.880 ;
        RECT 68.330 152.835 68.620 152.880 ;
        RECT 70.430 152.835 70.720 152.880 ;
        RECT 72.000 152.835 72.290 152.880 ;
        RECT 73.810 153.020 74.130 153.080 ;
        RECT 80.710 153.020 81.030 153.080 ;
        RECT 82.550 153.020 82.870 153.080 ;
        RECT 73.810 152.880 75.880 153.020 ;
        RECT 73.810 152.820 74.130 152.880 ;
        RECT 51.730 152.680 52.050 152.740 ;
        RECT 54.030 152.680 54.350 152.740 ;
        RECT 51.730 152.540 54.350 152.680 ;
        RECT 51.730 152.480 52.050 152.540 ;
        RECT 54.030 152.480 54.350 152.540 ;
        RECT 62.310 152.480 62.630 152.740 ;
        RECT 64.150 152.480 64.470 152.740 ;
        RECT 75.190 152.480 75.510 152.740 ;
        RECT 75.740 152.680 75.880 152.880 ;
        RECT 80.710 152.880 82.870 153.020 ;
        RECT 80.710 152.820 81.030 152.880 ;
        RECT 82.550 152.820 82.870 152.880 ;
        RECT 83.025 153.020 83.315 153.065 ;
        RECT 83.470 153.020 83.790 153.080 ;
        RECT 83.025 152.880 83.790 153.020 ;
        RECT 83.025 152.835 83.315 152.880 ;
        RECT 83.470 152.820 83.790 152.880 ;
        RECT 78.885 152.680 79.175 152.725 ;
        RECT 75.740 152.540 79.175 152.680 ;
        RECT 78.885 152.495 79.175 152.540 ;
        RECT 79.330 152.680 79.650 152.740 ;
        RECT 83.945 152.680 84.235 152.725 ;
        RECT 79.330 152.540 84.235 152.680 ;
        RECT 79.330 152.480 79.650 152.540 ;
        RECT 83.945 152.495 84.235 152.540 ;
        RECT 100.010 152.500 100.880 155.840 ;
        RECT 108.930 155.540 116.850 155.550 ;
        RECT 105.160 155.530 116.850 155.540 ;
        RECT 101.540 155.410 116.850 155.530 ;
        RECT 101.540 155.400 116.875 155.410 ;
        RECT 101.500 155.280 116.875 155.400 ;
        RECT 101.500 155.170 105.500 155.280 ;
        RECT 101.110 154.830 101.340 155.120 ;
        RECT 101.560 154.830 105.450 155.170 ;
        RECT 105.660 154.830 105.890 155.120 ;
        RECT 101.110 153.460 105.890 154.830 ;
        RECT 101.110 153.160 101.340 153.460 ;
        RECT 105.660 153.160 105.890 153.460 ;
        RECT 101.500 152.880 105.500 153.110 ;
        RECT 101.750 152.650 105.320 152.880 ;
        RECT 101.750 152.500 105.440 152.650 ;
        RECT 12.100 151.860 89.840 152.340 ;
        RECT 100.010 152.220 105.440 152.500 ;
        RECT 106.690 152.330 107.310 155.280 ;
        RECT 108.875 155.180 116.875 155.280 ;
        RECT 108.930 155.170 116.850 155.180 ;
        RECT 108.440 154.470 108.670 155.130 ;
        RECT 109.450 154.470 110.450 154.560 ;
        RECT 117.080 154.470 117.310 155.130 ;
        RECT 108.440 153.650 117.310 154.470 ;
        RECT 108.440 153.170 108.670 153.650 ;
        RECT 109.450 153.560 110.450 153.650 ;
        RECT 117.080 153.170 117.310 153.650 ;
        RECT 108.875 152.890 116.875 153.120 ;
        RECT 100.010 151.760 105.450 152.220 ;
        RECT 40.690 151.460 41.010 151.720 ;
        RECT 42.085 151.660 42.375 151.705 ;
        RECT 51.270 151.660 51.590 151.720 ;
        RECT 42.085 151.520 51.590 151.660 ;
        RECT 42.085 151.475 42.375 151.520 ;
        RECT 51.270 151.460 51.590 151.520 ;
        RECT 51.730 151.660 52.050 151.720 ;
        RECT 52.205 151.660 52.495 151.705 ;
        RECT 51.730 151.520 52.495 151.660 ;
        RECT 51.730 151.460 52.050 151.520 ;
        RECT 52.205 151.475 52.495 151.520 ;
        RECT 53.125 151.660 53.415 151.705 ;
        RECT 56.790 151.660 57.110 151.720 ;
        RECT 53.125 151.520 57.110 151.660 ;
        RECT 53.125 151.475 53.415 151.520 ;
        RECT 56.790 151.460 57.110 151.520 ;
        RECT 57.250 151.460 57.570 151.720 ;
        RECT 75.205 151.660 75.495 151.705 ;
        RECT 78.870 151.660 79.190 151.720 ;
        RECT 75.205 151.520 79.190 151.660 ;
        RECT 75.205 151.475 75.495 151.520 ;
        RECT 78.870 151.460 79.190 151.520 ;
        RECT 83.010 151.660 83.330 151.720 ;
        RECT 88.085 151.660 88.375 151.705 ;
        RECT 83.010 151.520 88.375 151.660 ;
        RECT 83.010 151.460 83.330 151.520 ;
        RECT 88.085 151.475 88.375 151.520 ;
        RECT 50.365 151.320 50.655 151.365 ;
        RECT 52.650 151.320 52.970 151.380 ;
        RECT 50.365 151.180 52.970 151.320 ;
        RECT 50.365 151.135 50.655 151.180 ;
        RECT 52.650 151.120 52.970 151.180 ;
        RECT 55.885 151.320 56.175 151.365 ;
        RECT 68.790 151.320 69.080 151.365 ;
        RECT 70.890 151.320 71.180 151.365 ;
        RECT 72.460 151.320 72.750 151.365 ;
        RECT 55.885 151.180 62.540 151.320 ;
        RECT 55.885 151.135 56.175 151.180 ;
        RECT 44.830 150.980 45.150 151.040 ;
        RECT 47.145 150.980 47.435 151.025 ;
        RECT 44.830 150.840 47.435 150.980 ;
        RECT 44.830 150.780 45.150 150.840 ;
        RECT 47.145 150.795 47.435 150.840 ;
        RECT 57.710 150.980 58.030 151.040 ;
        RECT 60.025 150.980 60.315 151.025 ;
        RECT 57.710 150.840 60.315 150.980 ;
        RECT 62.400 150.980 62.540 151.180 ;
        RECT 68.790 151.180 72.750 151.320 ;
        RECT 68.790 151.135 69.080 151.180 ;
        RECT 70.890 151.135 71.180 151.180 ;
        RECT 72.460 151.135 72.750 151.180 ;
        RECT 73.350 151.320 73.670 151.380 ;
        RECT 79.330 151.320 79.650 151.380 ;
        RECT 73.350 151.180 79.650 151.320 ;
        RECT 73.350 151.120 73.670 151.180 ;
        RECT 79.330 151.120 79.650 151.180 ;
        RECT 81.670 151.320 81.960 151.365 ;
        RECT 83.770 151.320 84.060 151.365 ;
        RECT 85.340 151.320 85.630 151.365 ;
        RECT 81.670 151.180 85.630 151.320 ;
        RECT 81.670 151.135 81.960 151.180 ;
        RECT 83.770 151.135 84.060 151.180 ;
        RECT 85.340 151.135 85.630 151.180 ;
        RECT 69.185 150.980 69.475 151.025 ;
        RECT 70.375 150.980 70.665 151.025 ;
        RECT 72.895 150.980 73.185 151.025 ;
        RECT 79.790 150.980 80.110 151.040 ;
        RECT 80.710 150.980 81.030 151.040 ;
        RECT 62.400 150.840 68.980 150.980 ;
        RECT 57.710 150.780 58.030 150.840 ;
        RECT 60.025 150.795 60.315 150.840 ;
        RECT 35.170 150.640 35.490 150.700 ;
        RECT 40.245 150.640 40.535 150.685 ;
        RECT 35.170 150.500 40.535 150.640 ;
        RECT 35.170 150.440 35.490 150.500 ;
        RECT 40.245 150.455 40.535 150.500 ;
        RECT 40.690 150.640 41.010 150.700 ;
        RECT 41.625 150.640 41.915 150.685 ;
        RECT 40.690 150.500 41.915 150.640 ;
        RECT 40.690 150.440 41.010 150.500 ;
        RECT 41.625 150.455 41.915 150.500 ;
        RECT 42.530 150.440 42.850 150.700 ;
        RECT 49.445 150.455 49.735 150.685 ;
        RECT 50.365 150.640 50.655 150.685 ;
        RECT 51.730 150.640 52.050 150.700 ;
        RECT 50.365 150.500 52.050 150.640 ;
        RECT 50.365 150.455 50.655 150.500 ;
        RECT 21.370 150.300 21.690 150.360 ;
        RECT 23.225 150.300 23.515 150.345 ;
        RECT 21.370 150.160 23.515 150.300 ;
        RECT 21.370 150.100 21.690 150.160 ;
        RECT 23.225 150.115 23.515 150.160 ;
        RECT 24.145 150.300 24.435 150.345 ;
        RECT 47.590 150.300 47.910 150.360 ;
        RECT 24.145 150.160 47.910 150.300 ;
        RECT 49.520 150.300 49.660 150.455 ;
        RECT 51.730 150.440 52.050 150.500 ;
        RECT 56.805 150.640 57.095 150.685 ;
        RECT 59.090 150.640 59.410 150.700 ;
        RECT 56.805 150.500 59.410 150.640 ;
        RECT 56.805 150.455 57.095 150.500 ;
        RECT 59.090 150.440 59.410 150.500 ;
        RECT 59.565 150.640 59.855 150.685 ;
        RECT 64.150 150.640 64.470 150.700 ;
        RECT 59.565 150.500 64.470 150.640 ;
        RECT 59.565 150.455 59.855 150.500 ;
        RECT 64.150 150.440 64.470 150.500 ;
        RECT 64.610 150.440 64.930 150.700 ;
        RECT 67.830 150.640 68.150 150.700 ;
        RECT 68.305 150.640 68.595 150.685 ;
        RECT 67.830 150.500 68.595 150.640 ;
        RECT 68.840 150.640 68.980 150.840 ;
        RECT 69.185 150.840 73.185 150.980 ;
        RECT 69.185 150.795 69.475 150.840 ;
        RECT 70.375 150.795 70.665 150.840 ;
        RECT 72.895 150.795 73.185 150.840 ;
        RECT 77.120 150.840 81.030 150.980 ;
        RECT 77.120 150.685 77.260 150.840 ;
        RECT 79.790 150.780 80.110 150.840 ;
        RECT 80.710 150.780 81.030 150.840 ;
        RECT 81.170 150.780 81.490 151.040 ;
        RECT 82.065 150.980 82.355 151.025 ;
        RECT 83.255 150.980 83.545 151.025 ;
        RECT 85.775 150.980 86.065 151.025 ;
        RECT 82.065 150.840 86.065 150.980 ;
        RECT 82.065 150.795 82.355 150.840 ;
        RECT 83.255 150.795 83.545 150.840 ;
        RECT 85.775 150.795 86.065 150.840 ;
        RECT 68.840 150.500 72.200 150.640 ;
        RECT 67.830 150.440 68.150 150.500 ;
        RECT 68.305 150.455 68.595 150.500 ;
        RECT 51.285 150.300 51.575 150.345 ;
        RECT 53.570 150.300 53.890 150.360 ;
        RECT 49.520 150.160 53.890 150.300 ;
        RECT 24.145 150.115 24.435 150.160 ;
        RECT 47.590 150.100 47.910 150.160 ;
        RECT 51.285 150.115 51.575 150.160 ;
        RECT 53.570 150.100 53.890 150.160 ;
        RECT 54.950 150.300 55.270 150.360 ;
        RECT 61.405 150.300 61.695 150.345 ;
        RECT 68.380 150.300 68.520 150.455 ;
        RECT 54.950 150.160 68.520 150.300 ;
        RECT 69.640 150.300 69.930 150.345 ;
        RECT 71.510 150.300 71.830 150.360 ;
        RECT 69.640 150.160 71.830 150.300 ;
        RECT 72.060 150.300 72.200 150.500 ;
        RECT 77.045 150.455 77.335 150.685 ;
        RECT 77.950 150.440 78.270 150.700 ;
        RECT 78.410 150.440 78.730 150.700 ;
        RECT 78.885 150.640 79.175 150.685 ;
        RECT 84.390 150.640 84.710 150.700 ;
        RECT 78.885 150.500 84.710 150.640 ;
        RECT 78.885 150.455 79.175 150.500 ;
        RECT 84.390 150.440 84.710 150.500 ;
        RECT 100.010 150.410 102.050 151.760 ;
        RECT 103.800 151.750 105.450 151.760 ;
        RECT 102.490 150.480 103.490 151.200 ;
        RECT 103.800 150.940 104.110 151.750 ;
        RECT 104.570 151.470 105.450 151.750 ;
        RECT 105.690 151.930 107.310 152.330 ;
        RECT 108.960 151.980 116.830 152.890 ;
        RECT 104.510 151.240 105.510 151.470 ;
        RECT 105.690 151.280 106.040 151.930 ;
        RECT 106.690 151.920 107.310 151.930 ;
        RECT 108.875 151.750 116.875 151.980 ;
        RECT 108.960 151.740 116.830 151.750 ;
        RECT 104.570 151.030 105.450 151.050 ;
        RECT 103.840 150.650 104.110 150.940 ;
        RECT 104.510 150.800 105.510 151.030 ;
        RECT 105.670 150.990 106.040 151.280 ;
        RECT 105.700 150.930 106.040 150.990 ;
        RECT 106.800 151.600 107.560 151.650 ;
        RECT 108.440 151.600 108.670 151.700 ;
        RECT 106.800 151.390 108.670 151.600 ;
        RECT 117.080 151.390 117.310 151.700 ;
        RECT 106.800 150.970 109.340 151.390 ;
        RECT 116.710 150.970 117.310 151.390 ;
        RECT 104.570 150.650 105.450 150.800 ;
        RECT 104.580 150.480 105.310 150.650 ;
        RECT 82.520 150.300 82.810 150.345 ;
        RECT 83.010 150.300 83.330 150.360 ;
        RECT 72.060 150.160 80.940 150.300 ;
        RECT 54.950 150.100 55.270 150.160 ;
        RECT 61.405 150.115 61.695 150.160 ;
        RECT 69.640 150.115 69.930 150.160 ;
        RECT 71.510 150.100 71.830 150.160 ;
        RECT 44.370 149.760 44.690 150.020 ;
        RECT 50.810 149.960 51.130 150.020 ;
        RECT 52.285 149.960 52.575 150.005 ;
        RECT 50.810 149.820 52.575 149.960 ;
        RECT 50.810 149.760 51.130 149.820 ;
        RECT 52.285 149.775 52.575 149.820 ;
        RECT 59.090 149.760 59.410 150.020 ;
        RECT 67.845 149.960 68.135 150.005 ;
        RECT 70.590 149.960 70.910 150.020 ;
        RECT 67.845 149.820 70.910 149.960 ;
        RECT 67.845 149.775 68.135 149.820 ;
        RECT 70.590 149.760 70.910 149.820 ;
        RECT 80.250 149.760 80.570 150.020 ;
        RECT 80.800 149.960 80.940 150.160 ;
        RECT 82.520 150.160 83.330 150.300 ;
        RECT 82.520 150.115 82.810 150.160 ;
        RECT 83.010 150.100 83.330 150.160 ;
        RECT 83.470 149.960 83.790 150.020 ;
        RECT 80.800 149.820 83.790 149.960 ;
        RECT 83.470 149.760 83.790 149.820 ;
        RECT 12.100 149.140 89.840 149.620 ;
        RECT 45.305 148.940 45.595 148.985 ;
        RECT 45.750 148.940 46.070 149.000 ;
        RECT 45.305 148.800 46.070 148.940 ;
        RECT 45.305 148.755 45.595 148.800 ;
        RECT 45.750 148.740 46.070 148.800 ;
        RECT 50.365 148.940 50.655 148.985 ;
        RECT 52.190 148.940 52.510 149.000 ;
        RECT 50.365 148.800 52.510 148.940 ;
        RECT 50.365 148.755 50.655 148.800 ;
        RECT 52.190 148.740 52.510 148.800 ;
        RECT 59.090 148.940 59.410 149.000 ;
        RECT 59.565 148.940 59.855 148.985 ;
        RECT 59.090 148.800 59.855 148.940 ;
        RECT 59.090 148.740 59.410 148.800 ;
        RECT 59.565 148.755 59.855 148.800 ;
        RECT 61.405 148.940 61.695 148.985 ;
        RECT 64.165 148.940 64.455 148.985 ;
        RECT 61.405 148.800 64.455 148.940 ;
        RECT 61.405 148.755 61.695 148.800 ;
        RECT 64.165 148.755 64.455 148.800 ;
        RECT 66.450 148.940 66.770 149.000 ;
        RECT 66.450 148.800 71.280 148.940 ;
        RECT 40.705 148.600 40.995 148.645 ;
        RECT 41.610 148.600 41.930 148.660 ;
        RECT 47.145 148.600 47.435 148.645 ;
        RECT 40.705 148.460 41.930 148.600 ;
        RECT 40.705 148.415 40.995 148.460 ;
        RECT 41.610 148.400 41.930 148.460 ;
        RECT 43.080 148.460 47.435 148.600 ;
        RECT 43.080 148.320 43.220 148.460 ;
        RECT 47.145 148.415 47.435 148.460 ;
        RECT 19.530 148.260 19.850 148.320 ;
        RECT 21.745 148.260 22.035 148.305 ;
        RECT 19.530 148.120 22.035 148.260 ;
        RECT 19.530 148.060 19.850 148.120 ;
        RECT 21.745 148.075 22.035 148.120 ;
        RECT 23.670 148.260 23.990 148.320 ;
        RECT 27.825 148.260 28.115 148.305 ;
        RECT 23.670 148.120 28.115 148.260 ;
        RECT 23.670 148.060 23.990 148.120 ;
        RECT 27.825 148.075 28.115 148.120 ;
        RECT 28.745 148.260 29.035 148.305 ;
        RECT 30.110 148.260 30.430 148.320 ;
        RECT 28.745 148.120 30.430 148.260 ;
        RECT 28.745 148.075 29.035 148.120 ;
        RECT 30.110 148.060 30.430 148.120 ;
        RECT 40.230 148.060 40.550 148.320 ;
        RECT 41.165 148.260 41.455 148.305 ;
        RECT 42.070 148.260 42.390 148.320 ;
        RECT 41.165 148.120 42.390 148.260 ;
        RECT 41.165 148.075 41.455 148.120 ;
        RECT 42.070 148.060 42.390 148.120 ;
        RECT 42.990 148.060 43.310 148.320 ;
        RECT 44.385 148.260 44.675 148.305 ;
        RECT 45.750 148.260 46.070 148.320 ;
        RECT 46.225 148.260 46.515 148.305 ;
        RECT 44.385 148.120 45.520 148.260 ;
        RECT 44.385 148.075 44.675 148.120 ;
        RECT 20.450 147.720 20.770 147.980 ;
        RECT 21.345 147.920 21.635 147.965 ;
        RECT 22.535 147.920 22.825 147.965 ;
        RECT 25.055 147.920 25.345 147.965 ;
        RECT 21.345 147.780 25.345 147.920 ;
        RECT 21.345 147.735 21.635 147.780 ;
        RECT 22.535 147.735 22.825 147.780 ;
        RECT 25.055 147.735 25.345 147.780 ;
        RECT 42.530 147.720 42.850 147.980 ;
        RECT 20.950 147.580 21.240 147.625 ;
        RECT 23.050 147.580 23.340 147.625 ;
        RECT 24.620 147.580 24.910 147.625 ;
        RECT 20.950 147.440 24.910 147.580 ;
        RECT 20.950 147.395 21.240 147.440 ;
        RECT 23.050 147.395 23.340 147.440 ;
        RECT 24.620 147.395 24.910 147.440 ;
        RECT 25.510 147.580 25.830 147.640 ;
        RECT 27.825 147.580 28.115 147.625 ;
        RECT 25.510 147.440 28.115 147.580 ;
        RECT 25.510 147.380 25.830 147.440 ;
        RECT 27.825 147.395 28.115 147.440 ;
        RECT 35.630 147.580 35.950 147.640 ;
        RECT 44.460 147.580 44.600 148.075 ;
        RECT 44.845 147.735 45.135 147.965 ;
        RECT 45.380 147.920 45.520 148.120 ;
        RECT 45.750 148.120 46.515 148.260 ;
        RECT 45.750 148.060 46.070 148.120 ;
        RECT 46.225 148.075 46.515 148.120 ;
        RECT 47.590 148.260 47.910 148.320 ;
        RECT 48.525 148.260 48.815 148.305 ;
        RECT 47.590 148.120 48.815 148.260 ;
        RECT 47.590 148.060 47.910 148.120 ;
        RECT 48.525 148.075 48.815 148.120 ;
        RECT 50.350 148.260 50.670 148.320 ;
        RECT 52.205 148.260 52.495 148.305 ;
        RECT 50.350 148.120 52.495 148.260 ;
        RECT 50.350 148.060 50.670 148.120 ;
        RECT 52.205 148.075 52.495 148.120 ;
        RECT 45.380 147.780 47.820 147.920 ;
        RECT 35.630 147.440 44.600 147.580 ;
        RECT 35.630 147.380 35.950 147.440 ;
        RECT 26.430 147.240 26.750 147.300 ;
        RECT 27.365 147.240 27.655 147.285 ;
        RECT 26.430 147.100 27.655 147.240 ;
        RECT 26.430 147.040 26.750 147.100 ;
        RECT 27.365 147.055 27.655 147.100 ;
        RECT 41.150 147.240 41.470 147.300 ;
        RECT 41.625 147.240 41.915 147.285 ;
        RECT 41.150 147.100 41.915 147.240 ;
        RECT 44.920 147.240 45.060 147.735 ;
        RECT 47.680 147.625 47.820 147.780 ;
        RECT 52.650 147.720 52.970 147.980 ;
        RECT 53.585 147.920 53.875 147.965 ;
        RECT 56.330 147.920 56.650 147.980 ;
        RECT 53.585 147.780 56.650 147.920 ;
        RECT 53.585 147.735 53.875 147.780 ;
        RECT 56.330 147.720 56.650 147.780 ;
        RECT 60.930 147.920 61.250 147.980 ;
        RECT 61.865 147.920 62.155 147.965 ;
        RECT 60.930 147.780 62.155 147.920 ;
        RECT 60.930 147.720 61.250 147.780 ;
        RECT 61.865 147.735 62.155 147.780 ;
        RECT 62.310 147.720 62.630 147.980 ;
        RECT 47.605 147.395 47.895 147.625 ;
        RECT 57.710 147.240 58.030 147.300 ;
        RECT 44.920 147.100 58.030 147.240 ;
        RECT 64.240 147.240 64.380 148.755 ;
        RECT 66.450 148.740 66.770 148.800 ;
        RECT 67.830 148.600 68.150 148.660 ;
        RECT 71.140 148.600 71.280 148.800 ;
        RECT 71.510 148.740 71.830 149.000 ;
        RECT 73.365 148.940 73.655 148.985 ;
        RECT 75.190 148.940 75.510 149.000 ;
        RECT 73.365 148.800 75.510 148.940 ;
        RECT 73.365 148.755 73.655 148.800 ;
        RECT 75.190 148.740 75.510 148.800 ;
        RECT 83.010 148.740 83.330 149.000 ;
        RECT 82.090 148.600 82.410 148.660 ;
        RECT 67.830 148.460 70.360 148.600 ;
        RECT 71.140 148.460 78.640 148.600 ;
        RECT 67.830 148.400 68.150 148.460 ;
        RECT 69.670 148.305 69.990 148.320 ;
        RECT 69.670 148.075 70.020 148.305 ;
        RECT 70.220 148.260 70.360 148.460 ;
        RECT 71.065 148.260 71.355 148.305 ;
        RECT 70.220 148.120 71.355 148.260 ;
        RECT 71.065 148.075 71.355 148.120 ;
        RECT 71.510 148.260 71.830 148.320 ;
        RECT 78.500 148.305 78.640 148.460 ;
        RECT 82.090 148.460 85.080 148.600 ;
        RECT 82.090 148.400 82.410 148.460 ;
        RECT 71.510 148.120 74.500 148.260 ;
        RECT 69.670 148.060 69.990 148.075 ;
        RECT 71.510 148.060 71.830 148.120 ;
        RECT 66.475 147.920 66.765 147.965 ;
        RECT 68.995 147.920 69.285 147.965 ;
        RECT 70.185 147.920 70.475 147.965 ;
        RECT 66.475 147.780 70.475 147.920 ;
        RECT 66.475 147.735 66.765 147.780 ;
        RECT 68.995 147.735 69.285 147.780 ;
        RECT 70.185 147.735 70.475 147.780 ;
        RECT 71.970 147.920 72.290 147.980 ;
        RECT 74.360 147.965 74.500 148.120 ;
        RECT 78.425 148.075 78.715 148.305 ;
        RECT 84.390 148.060 84.710 148.320 ;
        RECT 84.940 148.305 85.080 148.460 ;
        RECT 84.865 148.075 85.155 148.305 ;
        RECT 85.310 148.060 85.630 148.320 ;
        RECT 85.770 148.260 86.090 148.320 ;
        RECT 86.245 148.260 86.535 148.305 ;
        RECT 85.770 148.120 86.535 148.260 ;
        RECT 85.770 148.060 86.090 148.120 ;
        RECT 86.245 148.075 86.535 148.120 ;
        RECT 86.705 148.260 86.995 148.305 ;
        RECT 87.150 148.260 87.470 148.320 ;
        RECT 88.070 148.260 88.390 148.320 ;
        RECT 86.705 148.120 88.390 148.260 ;
        RECT 86.705 148.075 86.995 148.120 ;
        RECT 87.150 148.060 87.470 148.120 ;
        RECT 88.070 148.060 88.390 148.120 ;
        RECT 73.825 147.920 74.115 147.965 ;
        RECT 71.970 147.780 74.115 147.920 ;
        RECT 71.970 147.720 72.290 147.780 ;
        RECT 73.825 147.735 74.115 147.780 ;
        RECT 74.285 147.735 74.575 147.965 ;
        RECT 82.105 147.735 82.395 147.965 ;
        RECT 84.480 147.920 84.620 148.060 ;
        RECT 84.480 147.780 85.540 147.920 ;
        RECT 66.910 147.580 67.200 147.625 ;
        RECT 68.480 147.580 68.770 147.625 ;
        RECT 70.580 147.580 70.870 147.625 ;
        RECT 82.180 147.580 82.320 147.735 ;
        RECT 85.400 147.640 85.540 147.780 ;
        RECT 66.910 147.440 70.870 147.580 ;
        RECT 66.910 147.395 67.200 147.440 ;
        RECT 68.480 147.395 68.770 147.440 ;
        RECT 70.580 147.395 70.870 147.440 ;
        RECT 73.900 147.440 82.320 147.580 ;
        RECT 73.900 147.240 74.040 147.440 ;
        RECT 85.310 147.380 85.630 147.640 ;
        RECT 64.240 147.100 74.040 147.240 ;
        RECT 74.270 147.240 74.590 147.300 ;
        RECT 75.665 147.240 75.955 147.285 ;
        RECT 74.270 147.100 75.955 147.240 ;
        RECT 41.150 147.040 41.470 147.100 ;
        RECT 41.625 147.055 41.915 147.100 ;
        RECT 57.710 147.040 58.030 147.100 ;
        RECT 74.270 147.040 74.590 147.100 ;
        RECT 75.665 147.055 75.955 147.100 ;
        RECT 79.330 147.040 79.650 147.300 ;
        RECT 87.610 147.040 87.930 147.300 ;
        RECT 12.100 146.420 89.840 146.900 ;
        RECT 100.010 146.720 100.780 150.410 ;
        RECT 102.460 149.360 105.310 150.480 ;
        RECT 105.700 150.180 106.050 150.930 ;
        RECT 106.800 150.810 108.670 150.970 ;
        RECT 106.800 150.760 107.560 150.810 ;
        RECT 108.440 150.740 108.670 150.810 ;
        RECT 117.080 150.740 117.310 150.970 ;
        RECT 108.875 150.460 116.875 150.690 ;
        RECT 105.700 150.120 105.990 150.180 ;
        RECT 105.610 150.000 105.990 150.120 ;
        RECT 108.970 150.060 116.830 150.460 ;
        RECT 117.640 150.060 118.600 159.540 ;
        RECT 119.930 159.670 120.770 161.800 ;
        RECT 126.430 161.380 127.680 161.820 ;
        RECT 137.600 161.800 138.460 163.870 ;
        RECT 124.370 161.370 129.610 161.380 ;
        RECT 121.420 161.270 136.720 161.370 ;
        RECT 121.420 161.260 136.755 161.270 ;
        RECT 121.380 161.140 136.755 161.260 ;
        RECT 121.380 161.030 125.380 161.140 ;
        RECT 126.430 161.060 128.170 161.140 ;
        RECT 128.750 161.060 136.755 161.140 ;
        RECT 126.430 160.980 127.680 161.060 ;
        RECT 128.755 161.040 136.755 161.060 ;
        RECT 120.990 160.730 121.220 160.980 ;
        RECT 125.540 160.840 125.770 160.980 ;
        RECT 128.320 160.840 128.550 160.990 ;
        RECT 125.540 160.730 128.550 160.840 ;
        RECT 136.960 160.730 137.190 160.990 ;
        RECT 120.990 160.290 137.190 160.730 ;
        RECT 120.990 160.020 121.220 160.290 ;
        RECT 125.540 160.260 137.190 160.290 ;
        RECT 125.540 160.170 128.550 160.260 ;
        RECT 125.540 160.020 125.770 160.170 ;
        RECT 128.320 160.030 128.550 160.170 ;
        RECT 136.960 160.030 137.190 160.260 ;
        RECT 121.380 159.740 125.380 159.970 ;
        RECT 128.755 159.760 136.755 159.980 ;
        RECT 137.520 159.760 138.480 161.800 ;
        RECT 128.755 159.750 138.480 159.760 ;
        RECT 121.380 159.670 125.370 159.740 ;
        RECT 119.930 159.560 125.370 159.670 ;
        RECT 128.810 159.590 138.480 159.750 ;
        RECT 119.930 159.470 123.060 159.560 ;
        RECT 136.550 159.540 138.480 159.590 ;
        RECT 119.930 156.200 120.770 159.470 ;
        RECT 124.410 159.010 129.660 159.020 ;
        RECT 124.410 158.900 136.720 159.010 ;
        RECT 121.440 158.840 136.720 158.900 ;
        RECT 121.440 158.830 136.755 158.840 ;
        RECT 121.380 158.700 136.755 158.830 ;
        RECT 121.380 158.690 126.540 158.700 ;
        RECT 121.380 158.600 125.380 158.690 ;
        RECT 128.755 158.610 136.755 158.700 ;
        RECT 128.840 158.600 136.730 158.610 ;
        RECT 120.990 158.240 121.220 158.550 ;
        RECT 121.440 158.240 125.340 158.600 ;
        RECT 125.540 158.240 125.770 158.550 ;
        RECT 120.990 156.900 125.770 158.240 ;
        RECT 120.990 156.590 121.220 156.900 ;
        RECT 125.540 156.590 125.770 156.900 ;
        RECT 128.320 158.020 128.550 158.560 ;
        RECT 129.360 158.020 130.370 158.050 ;
        RECT 136.960 158.020 137.190 158.560 ;
        RECT 128.320 157.120 137.190 158.020 ;
        RECT 128.320 156.600 128.550 157.120 ;
        RECT 129.360 157.050 130.370 157.120 ;
        RECT 136.960 156.600 137.190 157.120 ;
        RECT 121.380 156.310 125.380 156.540 ;
        RECT 128.755 156.320 136.755 156.550 ;
        RECT 119.930 156.160 121.060 156.200 ;
        RECT 119.930 156.080 121.300 156.160 ;
        RECT 121.670 156.090 125.330 156.310 ;
        RECT 121.670 156.080 123.110 156.090 ;
        RECT 119.930 156.040 123.110 156.080 ;
        RECT 119.930 155.950 122.620 156.040 ;
        RECT 128.820 156.030 136.710 156.320 ;
        RECT 119.930 155.890 121.950 155.950 ;
        RECT 119.930 155.840 121.700 155.890 ;
        RECT 119.930 152.500 120.770 155.840 ;
        RECT 128.810 155.540 136.730 155.550 ;
        RECT 125.040 155.530 136.730 155.540 ;
        RECT 121.420 155.410 136.730 155.530 ;
        RECT 121.420 155.400 136.755 155.410 ;
        RECT 121.380 155.280 136.755 155.400 ;
        RECT 121.380 155.170 125.380 155.280 ;
        RECT 120.990 154.830 121.220 155.120 ;
        RECT 121.440 154.830 125.330 155.170 ;
        RECT 125.540 154.830 125.770 155.120 ;
        RECT 120.990 153.460 125.770 154.830 ;
        RECT 120.990 153.160 121.220 153.460 ;
        RECT 125.540 153.160 125.770 153.460 ;
        RECT 121.380 152.880 125.380 153.110 ;
        RECT 121.630 152.650 125.200 152.880 ;
        RECT 121.630 152.500 125.320 152.650 ;
        RECT 119.930 152.220 125.320 152.500 ;
        RECT 126.570 152.330 127.190 155.280 ;
        RECT 128.755 155.180 136.755 155.280 ;
        RECT 128.810 155.170 136.730 155.180 ;
        RECT 128.320 154.470 128.550 155.130 ;
        RECT 129.330 154.470 130.330 154.560 ;
        RECT 136.960 154.470 137.190 155.130 ;
        RECT 128.320 153.650 137.190 154.470 ;
        RECT 128.320 153.170 128.550 153.650 ;
        RECT 129.330 153.560 130.330 153.650 ;
        RECT 136.960 153.170 137.190 153.650 ;
        RECT 128.755 152.890 136.755 153.120 ;
        RECT 119.930 151.760 125.330 152.220 ;
        RECT 119.930 150.420 121.930 151.760 ;
        RECT 123.680 151.750 125.330 151.760 ;
        RECT 122.370 150.480 123.370 151.200 ;
        RECT 123.680 150.940 123.990 151.750 ;
        RECT 124.450 151.470 125.330 151.750 ;
        RECT 125.570 151.930 127.190 152.330 ;
        RECT 128.840 151.980 136.710 152.890 ;
        RECT 124.390 151.240 125.390 151.470 ;
        RECT 125.570 151.280 125.920 151.930 ;
        RECT 126.570 151.920 127.190 151.930 ;
        RECT 128.755 151.750 136.755 151.980 ;
        RECT 128.840 151.740 136.710 151.750 ;
        RECT 124.450 151.030 125.330 151.050 ;
        RECT 123.720 150.650 123.990 150.940 ;
        RECT 124.390 150.800 125.390 151.030 ;
        RECT 125.550 150.990 125.920 151.280 ;
        RECT 125.580 150.930 125.920 150.990 ;
        RECT 126.680 151.600 127.440 151.650 ;
        RECT 128.320 151.600 128.550 151.700 ;
        RECT 126.680 151.390 128.550 151.600 ;
        RECT 136.960 151.390 137.190 151.700 ;
        RECT 126.680 150.970 129.220 151.390 ;
        RECT 136.590 150.970 137.190 151.390 ;
        RECT 124.450 150.650 125.330 150.800 ;
        RECT 124.460 150.480 125.190 150.650 ;
        RECT 102.400 149.130 105.400 149.360 ;
        RECT 105.610 149.170 105.950 150.000 ;
        RECT 107.960 149.990 118.600 150.060 ;
        RECT 102.450 149.100 105.310 149.130 ;
        RECT 102.450 149.080 103.620 149.100 ;
        RECT 104.580 149.090 105.310 149.100 ;
        RECT 102.400 148.690 105.400 148.920 ;
        RECT 105.605 148.880 105.950 149.170 ;
        RECT 106.140 148.950 118.600 149.990 ;
        RECT 120.000 150.410 121.930 150.420 ;
        RECT 106.140 148.930 118.560 148.950 ;
        RECT 105.610 148.770 105.950 148.880 ;
        RECT 106.180 148.920 111.850 148.930 ;
        RECT 112.850 148.920 118.560 148.930 ;
        RECT 102.490 148.520 105.350 148.690 ;
        RECT 106.180 148.520 106.610 148.920 ;
        RECT 102.460 148.150 106.610 148.520 ;
        RECT 41.610 146.220 41.930 146.280 ;
        RECT 43.450 146.220 43.770 146.280 ;
        RECT 41.610 146.080 43.770 146.220 ;
        RECT 41.610 146.020 41.930 146.080 ;
        RECT 43.450 146.020 43.770 146.080 ;
        RECT 61.405 146.220 61.695 146.265 ;
        RECT 64.610 146.220 64.930 146.280 ;
        RECT 61.405 146.080 64.930 146.220 ;
        RECT 61.405 146.035 61.695 146.080 ;
        RECT 64.610 146.020 64.930 146.080 ;
        RECT 67.830 146.220 68.150 146.280 ;
        RECT 77.950 146.220 78.270 146.280 ;
        RECT 80.710 146.220 81.030 146.280 ;
        RECT 67.830 146.080 68.980 146.220 ;
        RECT 67.830 146.020 68.150 146.080 ;
        RECT 17.270 145.880 17.560 145.925 ;
        RECT 19.370 145.880 19.660 145.925 ;
        RECT 20.940 145.880 21.230 145.925 ;
        RECT 17.270 145.740 21.230 145.880 ;
        RECT 17.270 145.695 17.560 145.740 ;
        RECT 19.370 145.695 19.660 145.740 ;
        RECT 20.940 145.695 21.230 145.740 ;
        RECT 27.390 145.880 27.680 145.925 ;
        RECT 29.490 145.880 29.780 145.925 ;
        RECT 31.060 145.880 31.350 145.925 ;
        RECT 27.390 145.740 31.350 145.880 ;
        RECT 27.390 145.695 27.680 145.740 ;
        RECT 29.490 145.695 29.780 145.740 ;
        RECT 31.060 145.695 31.350 145.740 ;
        RECT 34.750 145.880 35.040 145.925 ;
        RECT 36.850 145.880 37.140 145.925 ;
        RECT 38.420 145.880 38.710 145.925 ;
        RECT 34.750 145.740 38.710 145.880 ;
        RECT 34.750 145.695 35.040 145.740 ;
        RECT 36.850 145.695 37.140 145.740 ;
        RECT 38.420 145.695 38.710 145.740 ;
        RECT 42.070 145.880 42.390 145.940 ;
        RECT 45.750 145.880 46.070 145.940 ;
        RECT 42.070 145.740 46.070 145.880 ;
        RECT 42.070 145.680 42.390 145.740 ;
        RECT 45.750 145.680 46.070 145.740 ;
        RECT 51.270 145.680 51.590 145.940 ;
        RECT 54.990 145.880 55.280 145.925 ;
        RECT 57.090 145.880 57.380 145.925 ;
        RECT 58.660 145.880 58.950 145.925 ;
        RECT 68.305 145.880 68.595 145.925 ;
        RECT 54.990 145.740 58.950 145.880 ;
        RECT 54.990 145.695 55.280 145.740 ;
        RECT 57.090 145.695 57.380 145.740 ;
        RECT 58.660 145.695 58.950 145.740 ;
        RECT 61.940 145.740 68.595 145.880 ;
        RECT 68.840 145.880 68.980 146.080 ;
        RECT 77.950 146.080 82.320 146.220 ;
        RECT 77.950 146.020 78.270 146.080 ;
        RECT 80.710 146.020 81.030 146.080 ;
        RECT 77.530 145.880 77.820 145.925 ;
        RECT 79.630 145.880 79.920 145.925 ;
        RECT 81.200 145.880 81.490 145.925 ;
        RECT 68.840 145.740 71.280 145.880 ;
        RECT 17.665 145.540 17.955 145.585 ;
        RECT 18.855 145.540 19.145 145.585 ;
        RECT 21.375 145.540 21.665 145.585 ;
        RECT 26.905 145.540 27.195 145.585 ;
        RECT 27.785 145.540 28.075 145.585 ;
        RECT 28.975 145.540 29.265 145.585 ;
        RECT 31.495 145.540 31.785 145.585 ;
        RECT 17.665 145.400 21.665 145.540 ;
        RECT 17.665 145.355 17.955 145.400 ;
        RECT 18.855 145.355 19.145 145.400 ;
        RECT 21.375 145.355 21.665 145.400 ;
        RECT 25.140 145.400 27.580 145.540 ;
        RECT 16.785 145.200 17.075 145.245 ;
        RECT 20.450 145.200 20.770 145.260 ;
        RECT 25.140 145.200 25.280 145.400 ;
        RECT 26.905 145.355 27.195 145.400 ;
        RECT 27.440 145.260 27.580 145.400 ;
        RECT 27.785 145.400 31.785 145.540 ;
        RECT 27.785 145.355 28.075 145.400 ;
        RECT 28.975 145.355 29.265 145.400 ;
        RECT 31.495 145.355 31.785 145.400 ;
        RECT 35.145 145.540 35.435 145.585 ;
        RECT 36.335 145.540 36.625 145.585 ;
        RECT 38.855 145.540 39.145 145.585 ;
        RECT 35.145 145.400 39.145 145.540 ;
        RECT 45.840 145.540 45.980 145.680 ;
        RECT 55.385 145.540 55.675 145.585 ;
        RECT 56.575 145.540 56.865 145.585 ;
        RECT 59.095 145.540 59.385 145.585 ;
        RECT 45.840 145.400 52.420 145.540 ;
        RECT 35.145 145.355 35.435 145.400 ;
        RECT 36.335 145.355 36.625 145.400 ;
        RECT 38.855 145.355 39.145 145.400 ;
        RECT 16.785 145.060 25.280 145.200 ;
        RECT 16.785 145.015 17.075 145.060 ;
        RECT 20.450 145.000 20.770 145.060 ;
        RECT 25.510 145.000 25.830 145.260 ;
        RECT 26.445 145.200 26.735 145.245 ;
        RECT 26.445 145.060 27.120 145.200 ;
        RECT 26.445 145.015 26.735 145.060 ;
        RECT 26.980 144.920 27.120 145.060 ;
        RECT 27.350 145.000 27.670 145.260 ;
        RECT 34.265 145.200 34.555 145.245 ;
        RECT 34.710 145.200 35.030 145.260 ;
        RECT 44.385 145.200 44.675 145.245 ;
        RECT 34.265 145.060 35.030 145.200 ;
        RECT 34.265 145.015 34.555 145.060 ;
        RECT 34.710 145.000 35.030 145.060 ;
        RECT 41.240 145.060 44.675 145.200 ;
        RECT 18.120 144.860 18.410 144.905 ;
        RECT 18.610 144.860 18.930 144.920 ;
        RECT 18.120 144.720 18.930 144.860 ;
        RECT 18.120 144.675 18.410 144.720 ;
        RECT 18.610 144.660 18.930 144.720 ;
        RECT 26.890 144.660 27.210 144.920 ;
        RECT 28.240 144.860 28.530 144.905 ;
        RECT 29.650 144.860 29.970 144.920 ;
        RECT 28.240 144.720 29.970 144.860 ;
        RECT 28.240 144.675 28.530 144.720 ;
        RECT 29.650 144.660 29.970 144.720 ;
        RECT 35.600 144.860 35.890 144.905 ;
        RECT 36.550 144.860 36.870 144.920 ;
        RECT 35.600 144.720 36.870 144.860 ;
        RECT 35.600 144.675 35.890 144.720 ;
        RECT 36.550 144.660 36.870 144.720 ;
        RECT 23.210 144.520 23.530 144.580 ;
        RECT 23.685 144.520 23.975 144.565 ;
        RECT 23.210 144.380 23.975 144.520 ;
        RECT 23.210 144.320 23.530 144.380 ;
        RECT 23.685 144.335 23.975 144.380 ;
        RECT 25.970 144.320 26.290 144.580 ;
        RECT 32.870 144.520 33.190 144.580 ;
        RECT 33.805 144.520 34.095 144.565 ;
        RECT 32.870 144.380 34.095 144.520 ;
        RECT 32.870 144.320 33.190 144.380 ;
        RECT 33.805 144.335 34.095 144.380 ;
        RECT 37.930 144.520 38.250 144.580 ;
        RECT 40.230 144.520 40.550 144.580 ;
        RECT 41.240 144.565 41.380 145.060 ;
        RECT 44.385 145.015 44.675 145.060 ;
        RECT 50.350 145.000 50.670 145.260 ;
        RECT 52.280 145.245 52.420 145.400 ;
        RECT 55.385 145.400 59.385 145.540 ;
        RECT 55.385 145.355 55.675 145.400 ;
        RECT 56.575 145.355 56.865 145.400 ;
        RECT 59.095 145.355 59.385 145.400 ;
        RECT 51.285 145.015 51.575 145.245 ;
        RECT 52.205 145.015 52.495 145.245 ;
        RECT 54.505 145.200 54.795 145.245 ;
        RECT 54.950 145.200 55.270 145.260 ;
        RECT 54.505 145.060 55.270 145.200 ;
        RECT 54.505 145.015 54.795 145.060 ;
        RECT 42.990 144.860 43.310 144.920 ;
        RECT 51.360 144.860 51.500 145.015 ;
        RECT 54.950 145.000 55.270 145.060 ;
        RECT 55.840 145.200 56.130 145.245 ;
        RECT 61.940 145.200 62.080 145.740 ;
        RECT 68.305 145.695 68.595 145.740 ;
        RECT 62.310 145.540 62.630 145.600 ;
        RECT 64.625 145.540 64.915 145.585 ;
        RECT 65.990 145.540 66.310 145.600 ;
        RECT 62.310 145.400 64.915 145.540 ;
        RECT 62.310 145.340 62.630 145.400 ;
        RECT 64.625 145.355 64.915 145.400 ;
        RECT 65.160 145.400 66.310 145.540 ;
        RECT 55.840 145.060 62.080 145.200 ;
        RECT 55.840 145.015 56.130 145.060 ;
        RECT 42.990 144.720 51.500 144.860 ;
        RECT 59.550 144.860 59.870 144.920 ;
        RECT 62.400 144.860 62.540 145.340 ;
        RECT 63.705 145.200 63.995 145.245 ;
        RECT 65.160 145.200 65.300 145.400 ;
        RECT 65.990 145.340 66.310 145.400 ;
        RECT 70.590 145.340 70.910 145.600 ;
        RECT 71.140 145.585 71.280 145.740 ;
        RECT 77.530 145.740 81.490 145.880 ;
        RECT 77.530 145.695 77.820 145.740 ;
        RECT 79.630 145.695 79.920 145.740 ;
        RECT 81.200 145.695 81.490 145.740 ;
        RECT 71.065 145.355 71.355 145.585 ;
        RECT 73.810 145.540 74.130 145.600 ;
        RECT 75.205 145.540 75.495 145.585 ;
        RECT 73.810 145.400 75.495 145.540 ;
        RECT 73.810 145.340 74.130 145.400 ;
        RECT 75.205 145.355 75.495 145.400 ;
        RECT 77.925 145.540 78.215 145.585 ;
        RECT 79.115 145.540 79.405 145.585 ;
        RECT 81.635 145.540 81.925 145.585 ;
        RECT 77.925 145.400 81.925 145.540 ;
        RECT 82.180 145.540 82.320 146.080 ;
        RECT 82.180 145.400 87.840 145.540 ;
        RECT 77.925 145.355 78.215 145.400 ;
        RECT 79.115 145.355 79.405 145.400 ;
        RECT 81.635 145.355 81.925 145.400 ;
        RECT 63.705 145.060 65.300 145.200 ;
        RECT 65.545 145.200 65.835 145.245 ;
        RECT 71.510 145.200 71.830 145.260 ;
        RECT 65.545 145.060 71.830 145.200 ;
        RECT 63.705 145.015 63.995 145.060 ;
        RECT 65.545 145.015 65.835 145.060 ;
        RECT 71.510 145.000 71.830 145.060 ;
        RECT 74.270 145.000 74.590 145.260 ;
        RECT 77.045 145.200 77.335 145.245 ;
        RECT 81.170 145.200 81.490 145.260 ;
        RECT 77.045 145.060 81.490 145.200 ;
        RECT 77.045 145.015 77.335 145.060 ;
        RECT 81.170 145.000 81.490 145.060 ;
        RECT 85.310 145.200 85.630 145.260 ;
        RECT 85.785 145.200 86.075 145.245 ;
        RECT 85.310 145.060 86.075 145.200 ;
        RECT 85.310 145.000 85.630 145.060 ;
        RECT 85.785 145.015 86.075 145.060 ;
        RECT 86.245 145.015 86.535 145.245 ;
        RECT 70.145 144.860 70.435 144.905 ;
        RECT 59.550 144.720 62.540 144.860 ;
        RECT 67.920 144.720 70.435 144.860 ;
        RECT 42.990 144.660 43.310 144.720 ;
        RECT 59.550 144.660 59.870 144.720 ;
        RECT 41.165 144.520 41.455 144.565 ;
        RECT 37.930 144.380 41.455 144.520 ;
        RECT 37.930 144.320 38.250 144.380 ;
        RECT 40.230 144.320 40.550 144.380 ;
        RECT 41.165 144.335 41.455 144.380 ;
        RECT 41.610 144.320 41.930 144.580 ;
        RECT 47.145 144.520 47.435 144.565 ;
        RECT 48.970 144.520 49.290 144.580 ;
        RECT 47.145 144.380 49.290 144.520 ;
        RECT 47.145 144.335 47.435 144.380 ;
        RECT 48.970 144.320 49.290 144.380 ;
        RECT 62.770 144.320 63.090 144.580 ;
        RECT 65.990 144.320 66.310 144.580 ;
        RECT 67.920 144.565 68.060 144.720 ;
        RECT 70.145 144.675 70.435 144.720 ;
        RECT 78.380 144.860 78.670 144.905 ;
        RECT 80.250 144.860 80.570 144.920 ;
        RECT 78.380 144.720 80.570 144.860 ;
        RECT 78.380 144.675 78.670 144.720 ;
        RECT 80.250 144.660 80.570 144.720 ;
        RECT 83.470 144.860 83.790 144.920 ;
        RECT 84.850 144.860 85.170 144.920 ;
        RECT 86.320 144.860 86.460 145.015 ;
        RECT 86.690 145.000 87.010 145.260 ;
        RECT 87.150 145.200 87.470 145.260 ;
        RECT 87.700 145.245 87.840 145.400 ;
        RECT 87.625 145.200 87.915 145.245 ;
        RECT 87.150 145.060 87.915 145.200 ;
        RECT 87.150 145.000 87.470 145.060 ;
        RECT 87.625 145.015 87.915 145.060 ;
        RECT 83.470 144.720 86.460 144.860 ;
        RECT 83.470 144.660 83.790 144.720 ;
        RECT 84.850 144.660 85.170 144.720 ;
        RECT 100.010 144.620 100.880 146.720 ;
        RECT 106.550 146.330 107.800 146.770 ;
        RECT 117.700 146.750 118.560 148.920 ;
        RECT 120.000 146.750 120.770 150.410 ;
        RECT 122.340 149.360 125.190 150.480 ;
        RECT 125.580 150.180 125.930 150.930 ;
        RECT 126.680 150.810 128.550 150.970 ;
        RECT 126.680 150.760 127.440 150.810 ;
        RECT 128.320 150.740 128.550 150.810 ;
        RECT 136.960 150.740 137.190 150.970 ;
        RECT 128.755 150.460 136.755 150.690 ;
        RECT 125.580 150.120 125.870 150.180 ;
        RECT 125.490 150.000 125.870 150.120 ;
        RECT 128.850 150.060 136.710 150.460 ;
        RECT 137.520 150.060 138.480 159.540 ;
        RECT 122.280 149.130 125.280 149.360 ;
        RECT 125.490 149.170 125.830 150.000 ;
        RECT 127.840 149.990 138.480 150.060 ;
        RECT 122.330 149.100 125.190 149.130 ;
        RECT 122.330 149.080 123.500 149.100 ;
        RECT 124.460 149.090 125.190 149.100 ;
        RECT 122.280 148.690 125.280 148.920 ;
        RECT 125.485 148.880 125.830 149.170 ;
        RECT 126.020 148.950 138.480 149.990 ;
        RECT 139.930 161.720 140.700 165.410 ;
        RECT 142.370 164.360 145.220 165.480 ;
        RECT 145.610 165.180 145.960 165.930 ;
        RECT 146.710 165.810 148.580 165.970 ;
        RECT 146.710 165.760 147.470 165.810 ;
        RECT 148.350 165.740 148.580 165.810 ;
        RECT 156.990 165.740 157.220 165.970 ;
        RECT 148.785 165.460 156.785 165.690 ;
        RECT 145.610 165.120 145.900 165.180 ;
        RECT 145.520 165.000 145.900 165.120 ;
        RECT 148.880 165.060 156.740 165.460 ;
        RECT 157.550 165.060 158.510 174.540 ;
        RECT 142.310 164.130 145.310 164.360 ;
        RECT 145.520 164.170 145.860 165.000 ;
        RECT 147.870 164.990 158.510 165.060 ;
        RECT 142.360 164.100 145.220 164.130 ;
        RECT 142.360 164.080 143.530 164.100 ;
        RECT 144.490 164.090 145.220 164.100 ;
        RECT 142.310 163.690 145.310 163.920 ;
        RECT 145.515 163.880 145.860 164.170 ;
        RECT 146.050 163.950 158.510 164.990 ;
        RECT 146.050 163.930 158.500 163.950 ;
        RECT 145.520 163.770 145.860 163.880 ;
        RECT 146.090 163.920 151.760 163.930 ;
        RECT 152.760 163.920 158.500 163.930 ;
        RECT 142.400 163.520 145.260 163.690 ;
        RECT 146.090 163.520 146.520 163.920 ;
        RECT 142.370 163.150 146.520 163.520 ;
        RECT 139.930 159.620 140.840 161.720 ;
        RECT 146.510 161.330 147.760 161.770 ;
        RECT 157.640 161.750 158.500 163.920 ;
        RECT 144.450 161.320 149.690 161.330 ;
        RECT 141.500 161.220 156.800 161.320 ;
        RECT 141.500 161.210 156.835 161.220 ;
        RECT 141.460 161.090 156.835 161.210 ;
        RECT 141.460 160.980 145.460 161.090 ;
        RECT 146.510 161.010 148.250 161.090 ;
        RECT 148.830 161.010 156.835 161.090 ;
        RECT 146.510 160.930 147.760 161.010 ;
        RECT 148.835 160.990 156.835 161.010 ;
        RECT 141.070 160.680 141.300 160.930 ;
        RECT 145.620 160.790 145.850 160.930 ;
        RECT 148.400 160.790 148.630 160.940 ;
        RECT 145.620 160.680 148.630 160.790 ;
        RECT 157.040 160.680 157.270 160.940 ;
        RECT 141.070 160.240 157.270 160.680 ;
        RECT 141.070 159.970 141.300 160.240 ;
        RECT 145.620 160.210 157.270 160.240 ;
        RECT 145.620 160.120 148.630 160.210 ;
        RECT 145.620 159.970 145.850 160.120 ;
        RECT 148.400 159.980 148.630 160.120 ;
        RECT 157.040 159.980 157.270 160.210 ;
        RECT 141.460 159.690 145.460 159.920 ;
        RECT 148.835 159.710 156.835 159.930 ;
        RECT 157.600 159.710 158.560 161.750 ;
        RECT 148.835 159.700 158.560 159.710 ;
        RECT 141.460 159.620 145.450 159.690 ;
        RECT 139.930 159.510 145.450 159.620 ;
        RECT 148.890 159.540 158.560 159.700 ;
        RECT 139.930 159.420 143.140 159.510 ;
        RECT 156.630 159.490 158.560 159.540 ;
        RECT 139.930 156.150 140.840 159.420 ;
        RECT 144.490 158.960 149.740 158.970 ;
        RECT 144.490 158.850 156.800 158.960 ;
        RECT 141.520 158.790 156.800 158.850 ;
        RECT 141.520 158.780 156.835 158.790 ;
        RECT 141.460 158.650 156.835 158.780 ;
        RECT 141.460 158.640 146.620 158.650 ;
        RECT 141.460 158.550 145.460 158.640 ;
        RECT 148.835 158.560 156.835 158.650 ;
        RECT 148.920 158.550 156.810 158.560 ;
        RECT 141.070 158.190 141.300 158.500 ;
        RECT 141.520 158.190 145.420 158.550 ;
        RECT 145.620 158.190 145.850 158.500 ;
        RECT 141.070 156.850 145.850 158.190 ;
        RECT 141.070 156.540 141.300 156.850 ;
        RECT 145.620 156.540 145.850 156.850 ;
        RECT 148.400 157.970 148.630 158.510 ;
        RECT 149.440 157.970 150.450 158.000 ;
        RECT 157.040 157.970 157.270 158.510 ;
        RECT 148.400 157.070 157.270 157.970 ;
        RECT 148.400 156.550 148.630 157.070 ;
        RECT 149.440 157.000 150.450 157.070 ;
        RECT 157.040 156.550 157.270 157.070 ;
        RECT 141.460 156.260 145.460 156.490 ;
        RECT 148.835 156.270 156.835 156.500 ;
        RECT 139.930 156.110 141.140 156.150 ;
        RECT 139.930 156.030 141.380 156.110 ;
        RECT 141.750 156.040 145.410 156.260 ;
        RECT 141.750 156.030 143.190 156.040 ;
        RECT 139.930 155.990 143.190 156.030 ;
        RECT 139.930 155.900 142.700 155.990 ;
        RECT 148.900 155.980 156.790 156.270 ;
        RECT 139.930 155.840 142.030 155.900 ;
        RECT 139.930 155.790 141.780 155.840 ;
        RECT 139.930 152.450 140.840 155.790 ;
        RECT 148.890 155.490 156.810 155.500 ;
        RECT 145.120 155.480 156.810 155.490 ;
        RECT 141.500 155.360 156.810 155.480 ;
        RECT 141.500 155.350 156.835 155.360 ;
        RECT 141.460 155.230 156.835 155.350 ;
        RECT 141.460 155.120 145.460 155.230 ;
        RECT 141.070 154.780 141.300 155.070 ;
        RECT 141.520 154.780 145.410 155.120 ;
        RECT 145.620 154.780 145.850 155.070 ;
        RECT 141.070 153.410 145.850 154.780 ;
        RECT 141.070 153.110 141.300 153.410 ;
        RECT 145.620 153.110 145.850 153.410 ;
        RECT 141.460 152.830 145.460 153.060 ;
        RECT 141.710 152.600 145.280 152.830 ;
        RECT 141.710 152.450 145.400 152.600 ;
        RECT 139.930 152.170 145.400 152.450 ;
        RECT 146.650 152.280 147.270 155.230 ;
        RECT 148.835 155.130 156.835 155.230 ;
        RECT 148.890 155.120 156.810 155.130 ;
        RECT 148.400 154.420 148.630 155.080 ;
        RECT 149.410 154.420 150.410 154.510 ;
        RECT 157.040 154.420 157.270 155.080 ;
        RECT 148.400 153.600 157.270 154.420 ;
        RECT 148.400 153.120 148.630 153.600 ;
        RECT 149.410 153.510 150.410 153.600 ;
        RECT 157.040 153.120 157.270 153.600 ;
        RECT 148.835 152.840 156.835 153.070 ;
        RECT 139.930 151.710 145.410 152.170 ;
        RECT 139.930 150.360 142.010 151.710 ;
        RECT 143.760 151.700 145.410 151.710 ;
        RECT 142.450 150.430 143.450 151.150 ;
        RECT 143.760 150.890 144.070 151.700 ;
        RECT 144.530 151.420 145.410 151.700 ;
        RECT 145.650 151.880 147.270 152.280 ;
        RECT 148.920 151.930 156.790 152.840 ;
        RECT 144.470 151.190 145.470 151.420 ;
        RECT 145.650 151.230 146.000 151.880 ;
        RECT 146.650 151.870 147.270 151.880 ;
        RECT 148.835 151.700 156.835 151.930 ;
        RECT 148.920 151.690 156.790 151.700 ;
        RECT 144.530 150.980 145.410 151.000 ;
        RECT 143.800 150.600 144.070 150.890 ;
        RECT 144.470 150.750 145.470 150.980 ;
        RECT 145.630 150.940 146.000 151.230 ;
        RECT 145.660 150.880 146.000 150.940 ;
        RECT 146.760 151.550 147.520 151.600 ;
        RECT 148.400 151.550 148.630 151.650 ;
        RECT 146.760 151.340 148.630 151.550 ;
        RECT 157.040 151.340 157.270 151.650 ;
        RECT 146.760 150.920 149.300 151.340 ;
        RECT 156.670 150.920 157.270 151.340 ;
        RECT 144.530 150.600 145.410 150.750 ;
        RECT 144.540 150.430 145.270 150.600 ;
        RECT 126.020 148.930 138.460 148.950 ;
        RECT 125.490 148.770 125.830 148.880 ;
        RECT 126.060 148.920 131.730 148.930 ;
        RECT 132.730 148.920 138.460 148.930 ;
        RECT 122.370 148.520 125.230 148.690 ;
        RECT 126.060 148.520 126.490 148.920 ;
        RECT 122.340 148.150 126.490 148.520 ;
        RECT 104.490 146.320 109.730 146.330 ;
        RECT 101.540 146.220 116.840 146.320 ;
        RECT 101.540 146.210 116.875 146.220 ;
        RECT 101.500 146.090 116.875 146.210 ;
        RECT 101.500 145.980 105.500 146.090 ;
        RECT 106.550 146.010 108.290 146.090 ;
        RECT 108.870 146.010 116.875 146.090 ;
        RECT 106.550 145.930 107.800 146.010 ;
        RECT 108.875 145.990 116.875 146.010 ;
        RECT 101.110 145.680 101.340 145.930 ;
        RECT 105.660 145.790 105.890 145.930 ;
        RECT 108.440 145.790 108.670 145.940 ;
        RECT 105.660 145.680 108.670 145.790 ;
        RECT 117.080 145.680 117.310 145.940 ;
        RECT 101.110 145.240 117.310 145.680 ;
        RECT 101.110 144.970 101.340 145.240 ;
        RECT 105.660 145.210 117.310 145.240 ;
        RECT 105.660 145.120 108.670 145.210 ;
        RECT 105.660 144.970 105.890 145.120 ;
        RECT 108.440 144.980 108.670 145.120 ;
        RECT 117.080 144.980 117.310 145.210 ;
        RECT 101.500 144.690 105.500 144.920 ;
        RECT 108.875 144.710 116.875 144.930 ;
        RECT 117.640 144.710 118.600 146.750 ;
        RECT 108.875 144.700 118.600 144.710 ;
        RECT 101.500 144.620 105.490 144.690 ;
        RECT 67.845 144.335 68.135 144.565 ;
        RECT 72.430 144.320 72.750 144.580 ;
        RECT 74.745 144.520 75.035 144.565 ;
        RECT 82.090 144.520 82.410 144.580 ;
        RECT 74.745 144.380 82.410 144.520 ;
        RECT 74.745 144.335 75.035 144.380 ;
        RECT 82.090 144.320 82.410 144.380 ;
        RECT 83.010 144.520 83.330 144.580 ;
        RECT 83.930 144.520 84.250 144.580 ;
        RECT 83.010 144.380 84.250 144.520 ;
        RECT 83.010 144.320 83.330 144.380 ;
        RECT 83.930 144.320 84.250 144.380 ;
        RECT 84.390 144.320 84.710 144.580 ;
        RECT 100.010 144.510 105.490 144.620 ;
        RECT 108.930 144.540 118.600 144.700 ;
        RECT 100.010 144.420 103.180 144.510 ;
        RECT 116.670 144.490 118.600 144.540 ;
        RECT 12.100 143.700 89.840 144.180 ;
        RECT 17.230 143.500 17.550 143.560 ;
        RECT 20.910 143.500 21.230 143.560 ;
        RECT 25.970 143.500 26.290 143.560 ;
        RECT 17.230 143.360 18.840 143.500 ;
        RECT 17.230 143.300 17.550 143.360 ;
        RECT 14.485 143.160 14.775 143.205 ;
        RECT 18.150 143.160 18.470 143.220 ;
        RECT 14.485 143.020 18.470 143.160 ;
        RECT 18.700 143.160 18.840 143.360 ;
        RECT 20.080 143.360 21.230 143.500 ;
        RECT 20.080 143.160 20.220 143.360 ;
        RECT 20.910 143.300 21.230 143.360 ;
        RECT 22.380 143.360 26.290 143.500 ;
        RECT 18.700 143.020 20.220 143.160 ;
        RECT 14.485 142.975 14.775 143.020 ;
        RECT 18.150 142.960 18.470 143.020 ;
        RECT 20.450 142.960 20.770 143.220 ;
        RECT 21.510 143.160 21.800 143.205 ;
        RECT 22.380 143.160 22.520 143.360 ;
        RECT 25.970 143.300 26.290 143.360 ;
        RECT 29.665 143.500 29.955 143.545 ;
        RECT 30.110 143.500 30.430 143.560 ;
        RECT 29.665 143.360 30.430 143.500 ;
        RECT 29.665 143.315 29.955 143.360 ;
        RECT 30.110 143.300 30.430 143.360 ;
        RECT 45.305 143.500 45.595 143.545 ;
        RECT 47.590 143.500 47.910 143.560 ;
        RECT 45.305 143.360 47.910 143.500 ;
        RECT 45.305 143.315 45.595 143.360 ;
        RECT 47.590 143.300 47.910 143.360 ;
        RECT 50.350 143.500 50.670 143.560 ;
        RECT 53.585 143.500 53.875 143.545 ;
        RECT 50.350 143.360 53.875 143.500 ;
        RECT 50.350 143.300 50.670 143.360 ;
        RECT 53.585 143.315 53.875 143.360 ;
        RECT 57.710 143.500 58.030 143.560 ;
        RECT 67.830 143.500 68.150 143.560 ;
        RECT 57.710 143.360 68.150 143.500 ;
        RECT 57.710 143.300 58.030 143.360 ;
        RECT 67.830 143.300 68.150 143.360 ;
        RECT 69.225 143.500 69.515 143.545 ;
        RECT 69.670 143.500 69.990 143.560 ;
        RECT 69.225 143.360 69.990 143.500 ;
        RECT 69.225 143.315 69.515 143.360 ;
        RECT 69.670 143.300 69.990 143.360 ;
        RECT 71.065 143.500 71.355 143.545 ;
        RECT 79.330 143.500 79.650 143.560 ;
        RECT 71.065 143.360 79.650 143.500 ;
        RECT 71.065 143.315 71.355 143.360 ;
        RECT 79.330 143.300 79.650 143.360 ;
        RECT 27.350 143.160 27.670 143.220 ;
        RECT 42.070 143.160 42.390 143.220 ;
        RECT 46.210 143.160 46.530 143.220 ;
        RECT 54.950 143.160 55.270 143.220 ;
        RECT 64.625 143.160 64.915 143.205 ;
        RECT 21.510 143.020 22.520 143.160 ;
        RECT 23.295 143.020 27.670 143.160 ;
        RECT 21.510 142.975 21.800 143.020 ;
        RECT 14.025 142.635 14.315 142.865 ;
        RECT 14.100 142.140 14.240 142.635 ;
        RECT 14.930 142.620 15.250 142.880 ;
        RECT 15.405 142.820 15.695 142.865 ;
        RECT 22.710 142.820 23.000 142.865 ;
        RECT 23.295 142.820 23.435 143.020 ;
        RECT 27.350 142.960 27.670 143.020 ;
        RECT 38.480 143.020 46.900 143.160 ;
        RECT 24.130 142.865 24.450 142.880 ;
        RECT 31.490 142.865 31.810 142.880 ;
        RECT 38.480 142.865 38.620 143.020 ;
        RECT 42.070 142.960 42.390 143.020 ;
        RECT 46.210 142.960 46.530 143.020 ;
        RECT 24.100 142.820 24.450 142.865 ;
        RECT 15.405 142.680 19.300 142.820 ;
        RECT 15.405 142.635 15.695 142.680 ;
        RECT 16.770 142.280 17.090 142.540 ;
        RECT 17.690 142.525 18.010 142.540 ;
        RECT 19.160 142.525 19.300 142.680 ;
        RECT 22.710 142.680 23.435 142.820 ;
        RECT 23.935 142.680 24.450 142.820 ;
        RECT 22.710 142.635 23.000 142.680 ;
        RECT 24.100 142.635 24.450 142.680 ;
        RECT 31.460 142.635 31.810 142.865 ;
        RECT 38.405 142.635 38.695 142.865 ;
        RECT 39.740 142.820 40.030 142.865 ;
        RECT 41.150 142.820 41.470 142.880 ;
        RECT 46.760 142.865 46.900 143.020 ;
        RECT 54.950 143.020 64.915 143.160 ;
        RECT 54.950 142.960 55.270 143.020 ;
        RECT 64.625 142.975 64.915 143.020 ;
        RECT 68.765 143.160 69.055 143.205 ;
        RECT 72.890 143.160 73.210 143.220 ;
        RECT 68.765 143.020 73.210 143.160 ;
        RECT 68.765 142.975 69.055 143.020 ;
        RECT 72.890 142.960 73.210 143.020 ;
        RECT 82.520 143.160 82.810 143.205 ;
        RECT 84.390 143.160 84.710 143.220 ;
        RECT 82.520 143.020 84.710 143.160 ;
        RECT 82.520 142.975 82.810 143.020 ;
        RECT 84.390 142.960 84.710 143.020 ;
        RECT 39.740 142.680 41.470 142.820 ;
        RECT 39.740 142.635 40.030 142.680 ;
        RECT 24.130 142.620 24.450 142.635 ;
        RECT 31.490 142.620 31.810 142.635 ;
        RECT 41.150 142.620 41.470 142.680 ;
        RECT 46.685 142.635 46.975 142.865 ;
        RECT 47.130 142.820 47.450 142.880 ;
        RECT 47.965 142.820 48.255 142.865 ;
        RECT 47.130 142.680 48.255 142.820 ;
        RECT 47.130 142.620 47.450 142.680 ;
        RECT 47.965 142.635 48.255 142.680 ;
        RECT 56.345 142.635 56.635 142.865 ;
        RECT 56.805 142.820 57.095 142.865 ;
        RECT 58.645 142.820 58.935 142.865 ;
        RECT 56.805 142.680 58.935 142.820 ;
        RECT 56.805 142.635 57.095 142.680 ;
        RECT 58.645 142.635 58.935 142.680 ;
        RECT 71.525 142.820 71.815 142.865 ;
        RECT 73.350 142.820 73.670 142.880 ;
        RECT 71.525 142.680 73.670 142.820 ;
        RECT 71.525 142.635 71.815 142.680 ;
        RECT 17.690 142.295 18.120 142.525 ;
        RECT 19.085 142.480 19.375 142.525 ;
        RECT 21.370 142.480 21.690 142.540 ;
        RECT 19.085 142.340 21.690 142.480 ;
        RECT 19.085 142.295 19.375 142.340 ;
        RECT 17.690 142.280 18.010 142.295 ;
        RECT 21.370 142.280 21.690 142.340 ;
        RECT 23.645 142.480 23.935 142.525 ;
        RECT 24.835 142.480 25.125 142.525 ;
        RECT 27.355 142.480 27.645 142.525 ;
        RECT 23.645 142.340 27.645 142.480 ;
        RECT 23.645 142.295 23.935 142.340 ;
        RECT 24.835 142.295 25.125 142.340 ;
        RECT 27.355 142.295 27.645 142.340 ;
        RECT 30.125 142.295 30.415 142.525 ;
        RECT 31.005 142.480 31.295 142.525 ;
        RECT 32.195 142.480 32.485 142.525 ;
        RECT 34.715 142.480 35.005 142.525 ;
        RECT 31.005 142.340 35.005 142.480 ;
        RECT 31.005 142.295 31.295 142.340 ;
        RECT 32.195 142.295 32.485 142.340 ;
        RECT 34.715 142.295 35.005 142.340 ;
        RECT 39.285 142.480 39.575 142.525 ;
        RECT 40.475 142.480 40.765 142.525 ;
        RECT 42.995 142.480 43.285 142.525 ;
        RECT 39.285 142.340 43.285 142.480 ;
        RECT 39.285 142.295 39.575 142.340 ;
        RECT 40.475 142.295 40.765 142.340 ;
        RECT 42.995 142.295 43.285 142.340 ;
        RECT 47.565 142.480 47.855 142.525 ;
        RECT 48.755 142.480 49.045 142.525 ;
        RECT 51.275 142.480 51.565 142.525 ;
        RECT 47.565 142.340 51.565 142.480 ;
        RECT 47.565 142.295 47.855 142.340 ;
        RECT 48.755 142.295 49.045 142.340 ;
        RECT 51.275 142.295 51.565 142.340 ;
        RECT 14.100 142.000 17.000 142.140 ;
        RECT 16.860 141.800 17.000 142.000 ;
        RECT 18.610 141.940 18.930 142.200 ;
        RECT 21.830 142.140 22.150 142.200 ;
        RECT 22.305 142.140 22.595 142.185 ;
        RECT 21.830 142.000 22.595 142.140 ;
        RECT 21.830 141.940 22.150 142.000 ;
        RECT 22.305 141.955 22.595 142.000 ;
        RECT 23.250 142.140 23.540 142.185 ;
        RECT 25.350 142.140 25.640 142.185 ;
        RECT 26.920 142.140 27.210 142.185 ;
        RECT 23.250 142.000 27.210 142.140 ;
        RECT 23.250 141.955 23.540 142.000 ;
        RECT 25.350 141.955 25.640 142.000 ;
        RECT 26.920 141.955 27.210 142.000 ;
        RECT 23.670 141.800 23.990 141.860 ;
        RECT 16.860 141.660 23.990 141.800 ;
        RECT 23.670 141.600 23.990 141.660 ;
        RECT 27.350 141.800 27.670 141.860 ;
        RECT 30.200 141.800 30.340 142.295 ;
        RECT 30.610 142.140 30.900 142.185 ;
        RECT 32.710 142.140 33.000 142.185 ;
        RECT 34.280 142.140 34.570 142.185 ;
        RECT 30.610 142.000 34.570 142.140 ;
        RECT 30.610 141.955 30.900 142.000 ;
        RECT 32.710 141.955 33.000 142.000 ;
        RECT 34.280 141.955 34.570 142.000 ;
        RECT 38.890 142.140 39.180 142.185 ;
        RECT 40.990 142.140 41.280 142.185 ;
        RECT 42.560 142.140 42.850 142.185 ;
        RECT 38.890 142.000 42.850 142.140 ;
        RECT 38.890 141.955 39.180 142.000 ;
        RECT 40.990 141.955 41.280 142.000 ;
        RECT 42.560 141.955 42.850 142.000 ;
        RECT 47.170 142.140 47.460 142.185 ;
        RECT 49.270 142.140 49.560 142.185 ;
        RECT 50.840 142.140 51.130 142.185 ;
        RECT 56.420 142.140 56.560 142.635 ;
        RECT 73.350 142.620 73.670 142.680 ;
        RECT 79.445 142.820 79.735 142.865 ;
        RECT 80.250 142.820 80.570 142.880 ;
        RECT 79.445 142.680 80.570 142.820 ;
        RECT 79.445 142.635 79.735 142.680 ;
        RECT 80.250 142.620 80.570 142.680 ;
        RECT 80.725 142.820 81.015 142.865 ;
        RECT 81.170 142.820 81.490 142.880 ;
        RECT 80.725 142.680 81.490 142.820 ;
        RECT 80.725 142.635 81.015 142.680 ;
        RECT 81.170 142.620 81.490 142.680 ;
        RECT 57.710 142.280 58.030 142.540 ;
        RECT 58.170 142.480 58.490 142.540 ;
        RECT 61.405 142.480 61.695 142.525 ;
        RECT 58.170 142.340 61.695 142.480 ;
        RECT 58.170 142.280 58.490 142.340 ;
        RECT 61.405 142.295 61.695 142.340 ;
        RECT 69.670 142.480 69.990 142.540 ;
        RECT 71.985 142.480 72.275 142.525 ;
        RECT 69.670 142.340 72.275 142.480 ;
        RECT 69.670 142.280 69.990 142.340 ;
        RECT 71.985 142.295 72.275 142.340 ;
        RECT 76.135 142.480 76.425 142.525 ;
        RECT 78.655 142.480 78.945 142.525 ;
        RECT 79.845 142.480 80.135 142.525 ;
        RECT 76.135 142.340 80.135 142.480 ;
        RECT 76.135 142.295 76.425 142.340 ;
        RECT 78.655 142.295 78.945 142.340 ;
        RECT 79.845 142.295 80.135 142.340 ;
        RECT 82.065 142.480 82.355 142.525 ;
        RECT 83.255 142.480 83.545 142.525 ;
        RECT 85.775 142.480 86.065 142.525 ;
        RECT 82.065 142.340 86.065 142.480 ;
        RECT 82.065 142.295 82.355 142.340 ;
        RECT 83.255 142.295 83.545 142.340 ;
        RECT 85.775 142.295 86.065 142.340 ;
        RECT 47.170 142.000 51.130 142.140 ;
        RECT 47.170 141.955 47.460 142.000 ;
        RECT 49.270 141.955 49.560 142.000 ;
        RECT 50.840 141.955 51.130 142.000 ;
        RECT 51.360 142.000 56.560 142.140 ;
        RECT 62.770 142.140 63.090 142.200 ;
        RECT 76.570 142.140 76.860 142.185 ;
        RECT 78.140 142.140 78.430 142.185 ;
        RECT 80.240 142.140 80.530 142.185 ;
        RECT 62.770 142.000 76.340 142.140 ;
        RECT 34.710 141.800 35.030 141.860 ;
        RECT 27.350 141.660 35.030 141.800 ;
        RECT 27.350 141.600 27.670 141.660 ;
        RECT 34.710 141.600 35.030 141.660 ;
        RECT 37.010 141.600 37.330 141.860 ;
        RECT 43.910 141.800 44.230 141.860 ;
        RECT 51.360 141.800 51.500 142.000 ;
        RECT 62.770 141.940 63.090 142.000 ;
        RECT 43.910 141.660 51.500 141.800 ;
        RECT 43.910 141.600 44.230 141.660 ;
        RECT 54.490 141.600 54.810 141.860 ;
        RECT 73.810 141.600 74.130 141.860 ;
        RECT 76.200 141.800 76.340 142.000 ;
        RECT 76.570 142.000 80.530 142.140 ;
        RECT 76.570 141.955 76.860 142.000 ;
        RECT 78.140 141.955 78.430 142.000 ;
        RECT 80.240 141.955 80.530 142.000 ;
        RECT 81.670 142.140 81.960 142.185 ;
        RECT 83.770 142.140 84.060 142.185 ;
        RECT 85.340 142.140 85.630 142.185 ;
        RECT 81.670 142.000 85.630 142.140 ;
        RECT 81.670 141.955 81.960 142.000 ;
        RECT 83.770 141.955 84.060 142.000 ;
        RECT 85.340 141.955 85.630 142.000 ;
        RECT 83.010 141.800 83.330 141.860 ;
        RECT 76.200 141.660 83.330 141.800 ;
        RECT 83.010 141.600 83.330 141.660 ;
        RECT 88.070 141.600 88.390 141.860 ;
        RECT 12.100 140.980 89.840 141.460 ;
        RECT 100.010 141.150 100.880 144.420 ;
        RECT 104.530 143.960 109.780 143.970 ;
        RECT 104.530 143.850 116.840 143.960 ;
        RECT 101.560 143.790 116.840 143.850 ;
        RECT 101.560 143.780 116.875 143.790 ;
        RECT 101.500 143.650 116.875 143.780 ;
        RECT 101.500 143.640 106.660 143.650 ;
        RECT 101.500 143.550 105.500 143.640 ;
        RECT 108.875 143.560 116.875 143.650 ;
        RECT 108.960 143.550 116.850 143.560 ;
        RECT 101.110 143.190 101.340 143.500 ;
        RECT 101.560 143.190 105.460 143.550 ;
        RECT 105.660 143.190 105.890 143.500 ;
        RECT 101.110 141.850 105.890 143.190 ;
        RECT 101.110 141.540 101.340 141.850 ;
        RECT 105.660 141.540 105.890 141.850 ;
        RECT 108.440 142.970 108.670 143.510 ;
        RECT 109.480 142.970 110.490 143.000 ;
        RECT 117.080 142.970 117.310 143.510 ;
        RECT 108.440 142.070 117.310 142.970 ;
        RECT 108.440 141.550 108.670 142.070 ;
        RECT 109.480 142.000 110.490 142.070 ;
        RECT 117.080 141.550 117.310 142.070 ;
        RECT 101.500 141.260 105.500 141.490 ;
        RECT 108.875 141.270 116.875 141.500 ;
        RECT 100.010 141.110 101.180 141.150 ;
        RECT 100.010 141.030 101.420 141.110 ;
        RECT 101.790 141.040 105.450 141.260 ;
        RECT 101.790 141.030 103.230 141.040 ;
        RECT 100.010 140.990 103.230 141.030 ;
        RECT 100.010 140.900 102.740 140.990 ;
        RECT 108.940 140.980 116.830 141.270 ;
        RECT 100.010 140.840 102.070 140.900 ;
        RECT 16.325 140.780 16.615 140.825 ;
        RECT 17.690 140.780 18.010 140.840 ;
        RECT 16.325 140.640 18.010 140.780 ;
        RECT 16.325 140.595 16.615 140.640 ;
        RECT 17.690 140.580 18.010 140.640 ;
        RECT 19.530 140.580 19.850 140.840 ;
        RECT 20.450 140.780 20.770 140.840 ;
        RECT 25.510 140.780 25.830 140.840 ;
        RECT 38.405 140.780 38.695 140.825 ;
        RECT 42.990 140.780 43.310 140.840 ;
        RECT 20.450 140.640 25.280 140.780 ;
        RECT 20.450 140.580 20.770 140.640 ;
        RECT 14.930 140.440 15.250 140.500 ;
        RECT 24.605 140.440 24.895 140.485 ;
        RECT 14.930 140.300 24.895 140.440 ;
        RECT 25.140 140.440 25.280 140.640 ;
        RECT 25.510 140.640 37.240 140.780 ;
        RECT 25.510 140.580 25.830 140.640 ;
        RECT 25.140 140.300 28.500 140.440 ;
        RECT 14.930 140.240 15.250 140.300 ;
        RECT 24.605 140.255 24.895 140.300 ;
        RECT 18.610 139.900 18.930 140.160 ;
        RECT 19.070 140.100 19.390 140.160 ;
        RECT 20.340 140.100 20.630 140.145 ;
        RECT 19.070 139.960 20.630 140.100 ;
        RECT 19.070 139.900 19.390 139.960 ;
        RECT 20.340 139.915 20.630 139.960 ;
        RECT 21.385 140.100 21.675 140.145 ;
        RECT 27.810 140.100 28.130 140.160 ;
        RECT 21.385 139.960 28.130 140.100 ;
        RECT 21.385 139.915 21.675 139.960 ;
        RECT 27.810 139.900 28.130 139.960 ;
        RECT 18.165 139.760 18.455 139.805 ;
        RECT 22.290 139.760 22.610 139.820 ;
        RECT 22.765 139.760 23.055 139.805 ;
        RECT 18.165 139.620 22.060 139.760 ;
        RECT 18.165 139.575 18.455 139.620 ;
        RECT 20.910 138.880 21.230 139.140 ;
        RECT 21.920 139.080 22.060 139.620 ;
        RECT 22.290 139.620 23.055 139.760 ;
        RECT 22.290 139.560 22.610 139.620 ;
        RECT 22.765 139.575 23.055 139.620 ;
        RECT 23.210 139.560 23.530 139.820 ;
        RECT 24.605 139.760 24.895 139.805 ;
        RECT 25.970 139.760 26.290 139.820 ;
        RECT 24.605 139.620 26.290 139.760 ;
        RECT 24.605 139.575 24.895 139.620 ;
        RECT 25.970 139.560 26.290 139.620 ;
        RECT 26.445 139.760 26.735 139.805 ;
        RECT 28.360 139.760 28.500 140.300 ;
        RECT 29.650 140.240 29.970 140.500 ;
        RECT 35.645 140.440 35.935 140.485 ;
        RECT 36.550 140.440 36.870 140.500 ;
        RECT 30.200 140.300 34.940 140.440 ;
        RECT 30.200 140.145 30.340 140.300 ;
        RECT 30.125 139.915 30.415 140.145 ;
        RECT 30.570 140.100 30.890 140.160 ;
        RECT 31.505 140.100 31.795 140.145 ;
        RECT 30.570 139.960 31.795 140.100 ;
        RECT 30.200 139.760 30.340 139.915 ;
        RECT 30.570 139.900 30.890 139.960 ;
        RECT 31.505 139.915 31.795 139.960 ;
        RECT 31.950 139.900 32.270 140.160 ;
        RECT 32.550 140.100 32.840 140.145 ;
        RECT 34.250 140.100 34.570 140.160 ;
        RECT 32.550 139.960 34.570 140.100 ;
        RECT 32.550 139.915 32.840 139.960 ;
        RECT 34.250 139.900 34.570 139.960 ;
        RECT 26.445 139.620 30.340 139.760 ;
        RECT 33.330 139.760 33.650 139.820 ;
        RECT 33.805 139.760 34.095 139.805 ;
        RECT 33.330 139.620 34.095 139.760 ;
        RECT 26.445 139.575 26.735 139.620 ;
        RECT 33.330 139.560 33.650 139.620 ;
        RECT 33.805 139.575 34.095 139.620 ;
        RECT 24.130 139.420 24.450 139.480 ;
        RECT 25.510 139.420 25.830 139.480 ;
        RECT 28.730 139.465 29.050 139.480 ;
        RECT 28.285 139.420 28.575 139.465 ;
        RECT 24.130 139.280 28.575 139.420 ;
        RECT 24.130 139.220 24.450 139.280 ;
        RECT 25.510 139.220 25.830 139.280 ;
        RECT 28.285 139.235 28.575 139.280 ;
        RECT 28.730 139.235 29.160 139.465 ;
        RECT 30.570 139.420 30.890 139.480 ;
        RECT 32.870 139.420 33.190 139.480 ;
        RECT 34.265 139.420 34.555 139.465 ;
        RECT 30.570 139.280 34.555 139.420 ;
        RECT 34.800 139.420 34.940 140.300 ;
        RECT 35.645 140.300 36.870 140.440 ;
        RECT 35.645 140.255 35.935 140.300 ;
        RECT 36.550 140.240 36.870 140.300 ;
        RECT 35.185 139.760 35.475 139.805 ;
        RECT 36.550 139.760 36.870 139.820 ;
        RECT 37.100 139.805 37.240 140.640 ;
        RECT 38.405 140.640 43.310 140.780 ;
        RECT 38.405 140.595 38.695 140.640 ;
        RECT 42.990 140.580 43.310 140.640 ;
        RECT 46.685 140.780 46.975 140.825 ;
        RECT 47.130 140.780 47.450 140.840 ;
        RECT 53.110 140.780 53.430 140.840 ;
        RECT 57.710 140.780 58.030 140.840 ;
        RECT 46.685 140.640 47.450 140.780 ;
        RECT 46.685 140.595 46.975 140.640 ;
        RECT 47.130 140.580 47.450 140.640 ;
        RECT 51.360 140.640 58.030 140.780 ;
        RECT 39.810 140.440 40.100 140.485 ;
        RECT 41.910 140.440 42.200 140.485 ;
        RECT 43.480 140.440 43.770 140.485 ;
        RECT 39.810 140.300 43.770 140.440 ;
        RECT 39.810 140.255 40.100 140.300 ;
        RECT 41.910 140.255 42.200 140.300 ;
        RECT 43.480 140.255 43.770 140.300 ;
        RECT 40.205 140.100 40.495 140.145 ;
        RECT 41.395 140.100 41.685 140.145 ;
        RECT 43.915 140.100 44.205 140.145 ;
        RECT 40.205 139.960 44.205 140.100 ;
        RECT 40.205 139.915 40.495 139.960 ;
        RECT 41.395 139.915 41.685 139.960 ;
        RECT 43.915 139.915 44.205 139.960 ;
        RECT 48.970 139.900 49.290 140.160 ;
        RECT 49.905 140.100 50.195 140.145 ;
        RECT 51.360 140.100 51.500 140.640 ;
        RECT 53.110 140.580 53.430 140.640 ;
        RECT 57.710 140.580 58.030 140.640 ;
        RECT 58.170 140.580 58.490 140.840 ;
        RECT 60.470 140.780 60.790 140.840 ;
        RECT 77.045 140.780 77.335 140.825 ;
        RECT 60.470 140.640 77.335 140.780 ;
        RECT 60.470 140.580 60.790 140.640 ;
        RECT 77.045 140.595 77.335 140.640 ;
        RECT 80.250 140.780 80.570 140.840 ;
        RECT 84.405 140.780 84.695 140.825 ;
        RECT 80.250 140.640 84.695 140.780 ;
        RECT 80.250 140.580 80.570 140.640 ;
        RECT 84.405 140.595 84.695 140.640 ;
        RECT 100.010 140.790 101.820 140.840 ;
        RECT 51.770 140.440 52.060 140.485 ;
        RECT 53.870 140.440 54.160 140.485 ;
        RECT 55.440 140.440 55.730 140.485 ;
        RECT 51.770 140.300 55.730 140.440 ;
        RECT 51.770 140.255 52.060 140.300 ;
        RECT 53.870 140.255 54.160 140.300 ;
        RECT 55.440 140.255 55.730 140.300 ;
        RECT 59.130 140.440 59.420 140.485 ;
        RECT 61.230 140.440 61.520 140.485 ;
        RECT 62.800 140.440 63.090 140.485 ;
        RECT 59.130 140.300 63.090 140.440 ;
        RECT 59.130 140.255 59.420 140.300 ;
        RECT 61.230 140.255 61.520 140.300 ;
        RECT 62.800 140.255 63.090 140.300 ;
        RECT 66.005 140.440 66.295 140.485 ;
        RECT 66.450 140.440 66.770 140.500 ;
        RECT 66.005 140.300 66.770 140.440 ;
        RECT 66.005 140.255 66.295 140.300 ;
        RECT 66.450 140.240 66.770 140.300 ;
        RECT 68.750 140.440 69.040 140.485 ;
        RECT 70.320 140.440 70.610 140.485 ;
        RECT 72.420 140.440 72.710 140.485 ;
        RECT 68.750 140.300 72.710 140.440 ;
        RECT 68.750 140.255 69.040 140.300 ;
        RECT 70.320 140.255 70.610 140.300 ;
        RECT 72.420 140.255 72.710 140.300 ;
        RECT 79.330 140.440 79.650 140.500 ;
        RECT 79.330 140.300 86.460 140.440 ;
        RECT 79.330 140.240 79.650 140.300 ;
        RECT 49.905 139.960 51.500 140.100 ;
        RECT 52.165 140.100 52.455 140.145 ;
        RECT 53.355 140.100 53.645 140.145 ;
        RECT 55.875 140.100 56.165 140.145 ;
        RECT 52.165 139.960 56.165 140.100 ;
        RECT 49.905 139.915 50.195 139.960 ;
        RECT 52.165 139.915 52.455 139.960 ;
        RECT 53.355 139.915 53.645 139.960 ;
        RECT 55.875 139.915 56.165 139.960 ;
        RECT 59.525 140.100 59.815 140.145 ;
        RECT 60.715 140.100 61.005 140.145 ;
        RECT 63.235 140.100 63.525 140.145 ;
        RECT 59.525 139.960 63.525 140.100 ;
        RECT 59.525 139.915 59.815 139.960 ;
        RECT 60.715 139.915 61.005 139.960 ;
        RECT 63.235 139.915 63.525 139.960 ;
        RECT 68.315 140.100 68.605 140.145 ;
        RECT 70.835 140.100 71.125 140.145 ;
        RECT 72.025 140.100 72.315 140.145 ;
        RECT 74.730 140.100 75.050 140.160 ;
        RECT 68.315 139.960 72.315 140.100 ;
        RECT 68.315 139.915 68.605 139.960 ;
        RECT 70.835 139.915 71.125 139.960 ;
        RECT 72.025 139.915 72.315 139.960 ;
        RECT 74.360 139.960 75.050 140.100 ;
        RECT 35.185 139.620 36.870 139.760 ;
        RECT 35.185 139.575 35.475 139.620 ;
        RECT 36.550 139.560 36.870 139.620 ;
        RECT 37.025 139.575 37.315 139.805 ;
        RECT 37.930 139.560 38.250 139.820 ;
        RECT 38.865 139.575 39.155 139.805 ;
        RECT 39.325 139.760 39.615 139.805 ;
        RECT 42.070 139.760 42.390 139.820 ;
        RECT 46.210 139.760 46.530 139.820 ;
        RECT 51.285 139.760 51.575 139.805 ;
        RECT 39.325 139.620 51.575 139.760 ;
        RECT 39.325 139.575 39.615 139.620 ;
        RECT 35.630 139.420 35.950 139.480 ;
        RECT 34.800 139.280 35.950 139.420 ;
        RECT 38.940 139.420 39.080 139.575 ;
        RECT 42.070 139.560 42.390 139.620 ;
        RECT 46.210 139.560 46.530 139.620 ;
        RECT 51.285 139.575 51.575 139.620 ;
        RECT 52.620 139.760 52.910 139.805 ;
        RECT 54.490 139.760 54.810 139.820 ;
        RECT 52.620 139.620 54.810 139.760 ;
        RECT 52.620 139.575 52.910 139.620 ;
        RECT 54.490 139.560 54.810 139.620 ;
        RECT 54.950 139.760 55.270 139.820 ;
        RECT 58.645 139.760 58.935 139.805 ;
        RECT 54.950 139.620 58.935 139.760 ;
        RECT 54.950 139.560 55.270 139.620 ;
        RECT 58.645 139.575 58.935 139.620 ;
        RECT 71.625 139.760 71.915 139.805 ;
        RECT 72.430 139.760 72.750 139.820 ;
        RECT 71.625 139.620 72.750 139.760 ;
        RECT 71.625 139.575 71.915 139.620 ;
        RECT 72.430 139.560 72.750 139.620 ;
        RECT 72.905 139.760 73.195 139.805 ;
        RECT 72.905 139.620 73.580 139.760 ;
        RECT 72.905 139.575 73.195 139.620 ;
        RECT 40.660 139.420 40.950 139.465 ;
        RECT 41.150 139.420 41.470 139.480 ;
        RECT 38.940 139.280 40.460 139.420 ;
        RECT 28.730 139.220 29.050 139.235 ;
        RECT 30.570 139.220 30.890 139.280 ;
        RECT 32.870 139.220 33.190 139.280 ;
        RECT 34.265 139.235 34.555 139.280 ;
        RECT 35.630 139.220 35.950 139.280 ;
        RECT 22.750 139.080 23.070 139.140 ;
        RECT 23.685 139.080 23.975 139.125 ;
        RECT 21.920 138.940 23.975 139.080 ;
        RECT 22.750 138.880 23.070 138.940 ;
        RECT 23.685 138.895 23.975 138.940 ;
        RECT 27.810 139.080 28.130 139.140 ;
        RECT 29.650 139.080 29.970 139.140 ;
        RECT 27.810 138.940 29.970 139.080 ;
        RECT 27.810 138.880 28.130 138.940 ;
        RECT 29.650 138.880 29.970 138.940 ;
        RECT 31.490 139.080 31.810 139.140 ;
        RECT 33.345 139.080 33.635 139.125 ;
        RECT 31.490 138.940 33.635 139.080 ;
        RECT 31.490 138.880 31.810 138.940 ;
        RECT 33.345 138.895 33.635 138.940 ;
        RECT 34.690 139.080 34.980 139.125 ;
        RECT 35.170 139.080 35.490 139.140 ;
        RECT 34.690 138.940 35.490 139.080 ;
        RECT 34.690 138.895 34.980 138.940 ;
        RECT 35.170 138.880 35.490 138.940 ;
        RECT 36.090 139.080 36.410 139.140 ;
        RECT 36.565 139.080 36.855 139.125 ;
        RECT 36.090 138.940 36.855 139.080 ;
        RECT 40.320 139.080 40.460 139.280 ;
        RECT 40.660 139.280 41.470 139.420 ;
        RECT 40.660 139.235 40.950 139.280 ;
        RECT 41.150 139.220 41.470 139.280 ;
        RECT 48.525 139.420 48.815 139.465 ;
        RECT 55.410 139.420 55.730 139.480 ;
        RECT 60.010 139.465 60.330 139.480 ;
        RECT 48.525 139.280 55.730 139.420 ;
        RECT 48.525 139.235 48.815 139.280 ;
        RECT 55.410 139.220 55.730 139.280 ;
        RECT 59.980 139.235 60.330 139.465 ;
        RECT 60.010 139.220 60.330 139.235 ;
        RECT 73.440 139.140 73.580 139.620 ;
        RECT 74.360 139.465 74.500 139.960 ;
        RECT 74.730 139.900 75.050 139.960 ;
        RECT 76.125 140.100 76.415 140.145 ;
        RECT 76.125 139.960 84.160 140.100 ;
        RECT 76.125 139.915 76.415 139.960 ;
        RECT 75.650 139.760 75.970 139.820 ;
        RECT 79.805 139.760 80.095 139.805 ;
        RECT 75.650 139.620 80.095 139.760 ;
        RECT 75.650 139.560 75.970 139.620 ;
        RECT 79.805 139.575 80.095 139.620 ;
        RECT 83.485 139.575 83.775 139.805 ;
        RECT 74.285 139.235 74.575 139.465 ;
        RECT 75.205 139.235 75.495 139.465 ;
        RECT 76.110 139.420 76.430 139.480 ;
        RECT 83.560 139.420 83.700 139.575 ;
        RECT 76.110 139.280 83.700 139.420 ;
        RECT 84.020 139.420 84.160 139.960 ;
        RECT 85.770 139.560 86.090 139.820 ;
        RECT 86.320 139.805 86.460 140.300 ;
        RECT 86.245 139.575 86.535 139.805 ;
        RECT 86.705 139.575 86.995 139.805 ;
        RECT 87.150 139.760 87.470 139.820 ;
        RECT 87.625 139.760 87.915 139.805 ;
        RECT 87.150 139.620 87.915 139.760 ;
        RECT 86.780 139.420 86.920 139.575 ;
        RECT 87.150 139.560 87.470 139.620 ;
        RECT 87.625 139.575 87.915 139.620 ;
        RECT 84.020 139.280 86.920 139.420 ;
        RECT 44.830 139.080 45.150 139.140 ;
        RECT 40.320 138.940 45.150 139.080 ;
        RECT 36.090 138.880 36.410 138.940 ;
        RECT 36.565 138.895 36.855 138.940 ;
        RECT 44.830 138.880 45.150 138.940 ;
        RECT 45.750 139.080 46.070 139.140 ;
        RECT 46.225 139.080 46.515 139.125 ;
        RECT 45.750 138.940 46.515 139.080 ;
        RECT 45.750 138.880 46.070 138.940 ;
        RECT 46.225 138.895 46.515 138.940 ;
        RECT 65.530 138.880 65.850 139.140 ;
        RECT 73.350 138.880 73.670 139.140 ;
        RECT 73.810 139.080 74.130 139.140 ;
        RECT 75.280 139.080 75.420 139.235 ;
        RECT 76.110 139.220 76.430 139.280 ;
        RECT 73.810 138.940 75.420 139.080 ;
        RECT 73.810 138.880 74.130 138.940 ;
        RECT 80.710 138.880 81.030 139.140 ;
        RECT 12.100 138.260 89.840 138.740 ;
        RECT 26.430 138.060 26.750 138.120 ;
        RECT 24.220 137.920 26.750 138.060 ;
        RECT 18.610 137.720 18.930 137.780 ;
        RECT 22.290 137.720 22.610 137.780 ;
        RECT 23.210 137.765 23.530 137.780 ;
        RECT 24.220 137.765 24.360 137.920 ;
        RECT 26.430 137.860 26.750 137.920 ;
        RECT 33.330 138.105 33.650 138.120 ;
        RECT 33.330 137.875 33.740 138.105 ;
        RECT 34.250 138.060 34.570 138.120 ;
        RECT 35.185 138.060 35.475 138.105 ;
        RECT 34.250 137.920 35.475 138.060 ;
        RECT 33.330 137.860 33.650 137.875 ;
        RECT 34.250 137.860 34.570 137.920 ;
        RECT 35.185 137.875 35.475 137.920 ;
        RECT 41.150 138.060 41.470 138.120 ;
        RECT 42.085 138.060 42.375 138.105 ;
        RECT 41.150 137.920 42.375 138.060 ;
        RECT 41.150 137.860 41.470 137.920 ;
        RECT 42.085 137.875 42.375 137.920 ;
        RECT 52.650 138.060 52.970 138.120 ;
        RECT 54.505 138.060 54.795 138.105 ;
        RECT 52.650 137.920 54.795 138.060 ;
        RECT 52.650 137.860 52.970 137.920 ;
        RECT 54.505 137.875 54.795 137.920 ;
        RECT 54.965 138.060 55.255 138.105 ;
        RECT 55.410 138.060 55.730 138.120 ;
        RECT 54.965 137.920 55.730 138.060 ;
        RECT 54.965 137.875 55.255 137.920 ;
        RECT 55.410 137.860 55.730 137.920 ;
        RECT 59.565 138.060 59.855 138.105 ;
        RECT 60.010 138.060 60.330 138.120 ;
        RECT 59.565 137.920 60.330 138.060 ;
        RECT 59.565 137.875 59.855 137.920 ;
        RECT 60.010 137.860 60.330 137.920 ;
        RECT 60.470 138.060 60.790 138.120 ;
        RECT 61.405 138.060 61.695 138.105 ;
        RECT 77.965 138.060 78.255 138.105 ;
        RECT 60.470 137.920 61.695 138.060 ;
        RECT 60.470 137.860 60.790 137.920 ;
        RECT 61.405 137.875 61.695 137.920 ;
        RECT 72.060 137.920 78.255 138.060 ;
        RECT 23.065 137.720 23.530 137.765 ;
        RECT 18.610 137.580 23.530 137.720 ;
        RECT 18.610 137.520 18.930 137.580 ;
        RECT 22.290 137.520 22.610 137.580 ;
        RECT 23.065 137.535 23.530 137.580 ;
        RECT 24.145 137.535 24.435 137.765 ;
        RECT 27.365 137.720 27.655 137.765 ;
        RECT 30.110 137.720 30.430 137.780 ;
        RECT 27.365 137.580 30.430 137.720 ;
        RECT 27.365 137.535 27.655 137.580 ;
        RECT 23.210 137.520 23.530 137.535 ;
        RECT 30.110 137.520 30.430 137.580 ;
        RECT 32.425 137.720 32.715 137.765 ;
        RECT 37.010 137.720 37.330 137.780 ;
        RECT 32.425 137.580 37.330 137.720 ;
        RECT 32.425 137.535 32.715 137.580 ;
        RECT 37.010 137.520 37.330 137.580 ;
        RECT 42.545 137.720 42.835 137.765 ;
        RECT 47.590 137.720 47.910 137.780 ;
        RECT 42.545 137.580 47.910 137.720 ;
        RECT 42.545 137.535 42.835 137.580 ;
        RECT 47.590 137.520 47.910 137.580 ;
        RECT 56.805 137.720 57.095 137.765 ;
        RECT 66.910 137.720 67.230 137.780 ;
        RECT 56.805 137.580 67.230 137.720 ;
        RECT 56.805 137.535 57.095 137.580 ;
        RECT 66.910 137.520 67.230 137.580 ;
        RECT 71.220 137.720 71.510 137.765 ;
        RECT 72.060 137.720 72.200 137.920 ;
        RECT 77.965 137.875 78.255 137.920 ;
        RECT 79.805 138.060 80.095 138.105 ;
        RECT 80.710 138.060 81.030 138.120 ;
        RECT 79.805 137.920 81.030 138.060 ;
        RECT 79.805 137.875 80.095 137.920 ;
        RECT 80.710 137.860 81.030 137.920 ;
        RECT 82.090 137.860 82.410 138.120 ;
        RECT 73.350 137.720 73.670 137.780 ;
        RECT 77.045 137.720 77.335 137.765 ;
        RECT 81.170 137.720 81.490 137.780 ;
        RECT 87.165 137.720 87.455 137.765 ;
        RECT 71.220 137.580 72.200 137.720 ;
        RECT 72.520 137.580 81.490 137.720 ;
        RECT 71.220 137.535 71.510 137.580 ;
        RECT 23.300 137.380 23.440 137.520 ;
        RECT 25.525 137.380 25.815 137.425 ;
        RECT 23.300 137.240 25.815 137.380 ;
        RECT 25.525 137.195 25.815 137.240 ;
        RECT 25.985 137.195 26.275 137.425 ;
        RECT 29.665 137.380 29.955 137.425 ;
        RECT 30.570 137.380 30.890 137.440 ;
        RECT 29.665 137.240 30.890 137.380 ;
        RECT 29.665 137.195 29.955 137.240 ;
        RECT 26.060 137.040 26.200 137.195 ;
        RECT 30.570 137.180 30.890 137.240 ;
        RECT 34.725 137.380 35.015 137.425 ;
        RECT 35.170 137.380 35.490 137.440 ;
        RECT 34.725 137.240 35.490 137.380 ;
        RECT 34.725 137.195 35.015 137.240 ;
        RECT 35.170 137.180 35.490 137.240 ;
        RECT 35.630 137.180 35.950 137.440 ;
        RECT 37.485 137.380 37.775 137.425 ;
        RECT 45.750 137.380 46.070 137.440 ;
        RECT 37.485 137.240 46.070 137.380 ;
        RECT 37.485 137.195 37.775 137.240 ;
        RECT 45.750 137.180 46.070 137.240 ;
        RECT 46.210 137.380 46.530 137.440 ;
        RECT 48.940 137.380 49.230 137.425 ;
        RECT 51.730 137.380 52.050 137.440 ;
        RECT 46.210 137.240 47.820 137.380 ;
        RECT 46.210 137.180 46.530 137.240 ;
        RECT 24.220 136.900 26.200 137.040 ;
        RECT 27.825 137.040 28.115 137.085 ;
        RECT 28.730 137.040 29.050 137.100 ;
        RECT 27.825 136.900 29.050 137.040 ;
        RECT 22.305 136.700 22.595 136.745 ;
        RECT 23.670 136.700 23.990 136.760 ;
        RECT 22.305 136.560 23.990 136.700 ;
        RECT 22.305 136.515 22.595 136.560 ;
        RECT 23.670 136.500 23.990 136.560 ;
        RECT 22.750 136.360 23.070 136.420 ;
        RECT 23.225 136.360 23.515 136.405 ;
        RECT 24.220 136.360 24.360 136.900 ;
        RECT 27.825 136.855 28.115 136.900 ;
        RECT 28.730 136.840 29.050 136.900 ;
        RECT 30.125 137.040 30.415 137.085 ;
        RECT 33.330 137.040 33.650 137.100 ;
        RECT 30.125 136.900 33.650 137.040 ;
        RECT 30.125 136.855 30.415 136.900 ;
        RECT 24.605 136.700 24.895 136.745 ;
        RECT 26.890 136.700 27.210 136.760 ;
        RECT 30.200 136.700 30.340 136.855 ;
        RECT 33.330 136.840 33.650 136.900 ;
        RECT 39.310 136.840 39.630 137.100 ;
        RECT 47.680 137.085 47.820 137.240 ;
        RECT 48.940 137.240 52.050 137.380 ;
        RECT 48.940 137.195 49.230 137.240 ;
        RECT 51.730 137.180 52.050 137.240 ;
        RECT 57.265 137.380 57.555 137.425 ;
        RECT 58.630 137.380 58.950 137.440 ;
        RECT 57.265 137.240 58.950 137.380 ;
        RECT 57.265 137.195 57.555 137.240 ;
        RECT 58.630 137.180 58.950 137.240 ;
        RECT 61.865 137.380 62.155 137.425 ;
        RECT 65.070 137.380 65.390 137.440 ;
        RECT 72.520 137.425 72.660 137.580 ;
        RECT 73.350 137.520 73.670 137.580 ;
        RECT 77.045 137.535 77.335 137.580 ;
        RECT 81.170 137.520 81.490 137.580 ;
        RECT 82.180 137.580 83.700 137.720 ;
        RECT 61.865 137.240 65.390 137.380 ;
        RECT 61.865 137.195 62.155 137.240 ;
        RECT 65.070 137.180 65.390 137.240 ;
        RECT 72.445 137.195 72.735 137.425 ;
        RECT 72.890 137.180 73.210 137.440 ;
        RECT 73.810 137.380 74.130 137.440 ;
        RECT 82.180 137.380 82.320 137.580 ;
        RECT 73.810 137.240 82.320 137.380 ;
        RECT 82.550 137.380 82.870 137.440 ;
        RECT 83.560 137.425 83.700 137.580 ;
        RECT 85.860 137.580 87.455 137.720 ;
        RECT 83.025 137.380 83.315 137.425 ;
        RECT 82.550 137.240 83.315 137.380 ;
        RECT 73.810 137.180 74.130 137.240 ;
        RECT 82.550 137.180 82.870 137.240 ;
        RECT 83.025 137.195 83.315 137.240 ;
        RECT 83.485 137.195 83.775 137.425 ;
        RECT 84.390 137.180 84.710 137.440 ;
        RECT 84.850 137.180 85.170 137.440 ;
        RECT 47.605 136.855 47.895 137.085 ;
        RECT 48.485 137.040 48.775 137.085 ;
        RECT 49.675 137.040 49.965 137.085 ;
        RECT 52.195 137.040 52.485 137.085 ;
        RECT 48.485 136.900 52.485 137.040 ;
        RECT 48.485 136.855 48.775 136.900 ;
        RECT 49.675 136.855 49.965 136.900 ;
        RECT 52.195 136.855 52.485 136.900 ;
        RECT 57.710 137.040 58.030 137.100 ;
        RECT 59.550 137.040 59.870 137.100 ;
        RECT 57.710 136.900 59.870 137.040 ;
        RECT 57.710 136.840 58.030 136.900 ;
        RECT 59.550 136.840 59.870 136.900 ;
        RECT 62.325 136.855 62.615 137.085 ;
        RECT 67.855 137.040 68.145 137.085 ;
        RECT 70.375 137.040 70.665 137.085 ;
        RECT 71.565 137.040 71.855 137.085 ;
        RECT 67.855 136.900 71.855 137.040 ;
        RECT 67.855 136.855 68.145 136.900 ;
        RECT 70.375 136.855 70.665 136.900 ;
        RECT 71.565 136.855 71.855 136.900 ;
        RECT 78.870 137.040 79.190 137.100 ;
        RECT 80.265 137.040 80.555 137.085 ;
        RECT 78.870 136.900 80.555 137.040 ;
        RECT 24.605 136.560 30.340 136.700 ;
        RECT 37.025 136.700 37.315 136.745 ;
        RECT 42.530 136.700 42.850 136.760 ;
        RECT 37.025 136.560 42.850 136.700 ;
        RECT 24.605 136.515 24.895 136.560 ;
        RECT 26.890 136.500 27.210 136.560 ;
        RECT 37.025 136.515 37.315 136.560 ;
        RECT 42.530 136.500 42.850 136.560 ;
        RECT 48.090 136.700 48.380 136.745 ;
        RECT 50.190 136.700 50.480 136.745 ;
        RECT 51.760 136.700 52.050 136.745 ;
        RECT 48.090 136.560 52.050 136.700 ;
        RECT 48.090 136.515 48.380 136.560 ;
        RECT 50.190 136.515 50.480 136.560 ;
        RECT 51.760 136.515 52.050 136.560 ;
        RECT 61.390 136.700 61.710 136.760 ;
        RECT 62.400 136.700 62.540 136.855 ;
        RECT 78.870 136.840 79.190 136.900 ;
        RECT 80.265 136.855 80.555 136.900 ;
        RECT 80.710 136.840 81.030 137.100 ;
        RECT 61.390 136.560 62.540 136.700 ;
        RECT 68.290 136.700 68.580 136.745 ;
        RECT 69.860 136.700 70.150 136.745 ;
        RECT 71.960 136.700 72.250 136.745 ;
        RECT 68.290 136.560 72.250 136.700 ;
        RECT 61.390 136.500 61.710 136.560 ;
        RECT 68.290 136.515 68.580 136.560 ;
        RECT 69.860 136.515 70.150 136.560 ;
        RECT 71.960 136.515 72.250 136.560 ;
        RECT 78.410 136.700 78.730 136.760 ;
        RECT 85.325 136.700 85.615 136.745 ;
        RECT 78.410 136.560 85.615 136.700 ;
        RECT 78.410 136.500 78.730 136.560 ;
        RECT 85.325 136.515 85.615 136.560 ;
        RECT 85.860 136.420 86.000 137.580 ;
        RECT 87.165 137.535 87.455 137.580 ;
        RECT 100.010 137.450 100.880 140.790 ;
        RECT 108.930 140.490 116.850 140.500 ;
        RECT 105.160 140.480 116.850 140.490 ;
        RECT 101.540 140.360 116.850 140.480 ;
        RECT 101.540 140.350 116.875 140.360 ;
        RECT 101.500 140.230 116.875 140.350 ;
        RECT 101.500 140.120 105.500 140.230 ;
        RECT 101.110 139.780 101.340 140.070 ;
        RECT 101.560 139.780 105.450 140.120 ;
        RECT 105.660 139.780 105.890 140.070 ;
        RECT 101.110 138.410 105.890 139.780 ;
        RECT 101.110 138.110 101.340 138.410 ;
        RECT 105.660 138.110 105.890 138.410 ;
        RECT 101.500 137.830 105.500 138.060 ;
        RECT 101.750 137.600 105.320 137.830 ;
        RECT 101.750 137.450 105.440 137.600 ;
        RECT 86.245 137.195 86.535 137.425 ;
        RECT 86.320 137.040 86.460 137.195 ;
        RECT 100.010 137.170 105.440 137.450 ;
        RECT 106.690 137.280 107.310 140.230 ;
        RECT 108.875 140.130 116.875 140.230 ;
        RECT 108.930 140.120 116.850 140.130 ;
        RECT 108.440 139.420 108.670 140.080 ;
        RECT 109.450 139.420 110.450 139.510 ;
        RECT 117.080 139.420 117.310 140.080 ;
        RECT 108.440 138.600 117.310 139.420 ;
        RECT 108.440 138.120 108.670 138.600 ;
        RECT 109.450 138.510 110.450 138.600 ;
        RECT 117.080 138.120 117.310 138.600 ;
        RECT 108.875 137.840 116.875 138.070 ;
        RECT 87.610 137.040 87.930 137.100 ;
        RECT 86.320 136.900 87.930 137.040 ;
        RECT 87.610 136.840 87.930 136.900 ;
        RECT 100.010 136.710 105.450 137.170 ;
        RECT 22.750 136.220 24.360 136.360 ;
        RECT 30.570 136.360 30.890 136.420 ;
        RECT 33.345 136.360 33.635 136.405 ;
        RECT 30.570 136.220 33.635 136.360 ;
        RECT 22.750 136.160 23.070 136.220 ;
        RECT 23.225 136.175 23.515 136.220 ;
        RECT 30.570 136.160 30.890 136.220 ;
        RECT 33.345 136.175 33.635 136.220 ;
        RECT 34.265 136.360 34.555 136.405 ;
        RECT 35.630 136.360 35.950 136.420 ;
        RECT 34.265 136.220 35.950 136.360 ;
        RECT 34.265 136.175 34.555 136.220 ;
        RECT 35.630 136.160 35.950 136.220 ;
        RECT 65.545 136.360 65.835 136.405 ;
        RECT 65.990 136.360 66.310 136.420 ;
        RECT 76.110 136.360 76.430 136.420 ;
        RECT 65.545 136.220 76.430 136.360 ;
        RECT 65.545 136.175 65.835 136.220 ;
        RECT 65.990 136.160 66.310 136.220 ;
        RECT 76.110 136.160 76.430 136.220 ;
        RECT 77.490 136.360 77.810 136.420 ;
        RECT 85.770 136.360 86.090 136.420 ;
        RECT 77.490 136.220 86.090 136.360 ;
        RECT 77.490 136.160 77.810 136.220 ;
        RECT 85.770 136.160 86.090 136.220 ;
        RECT 12.100 135.540 89.840 136.020 ;
        RECT 39.310 135.340 39.630 135.400 ;
        RECT 39.785 135.340 40.075 135.385 ;
        RECT 39.310 135.200 40.075 135.340 ;
        RECT 39.310 135.140 39.630 135.200 ;
        RECT 39.785 135.155 40.075 135.200 ;
        RECT 41.610 135.140 41.930 135.400 ;
        RECT 44.830 135.140 45.150 135.400 ;
        RECT 45.750 135.140 46.070 135.400 ;
        RECT 47.130 135.140 47.450 135.400 ;
        RECT 51.730 135.140 52.050 135.400 ;
        RECT 61.850 135.140 62.170 135.400 ;
        RECT 69.670 135.340 69.990 135.400 ;
        RECT 80.710 135.340 81.030 135.400 ;
        RECT 69.670 135.200 81.030 135.340 ;
        RECT 69.670 135.140 69.990 135.200 ;
        RECT 80.710 135.140 81.030 135.200 ;
        RECT 100.010 135.360 102.050 136.710 ;
        RECT 103.800 136.700 105.450 136.710 ;
        RECT 102.490 135.430 103.490 136.150 ;
        RECT 103.800 135.890 104.110 136.700 ;
        RECT 104.570 136.420 105.450 136.700 ;
        RECT 105.690 136.880 107.310 137.280 ;
        RECT 108.960 136.930 116.830 137.840 ;
        RECT 104.510 136.190 105.510 136.420 ;
        RECT 105.690 136.230 106.040 136.880 ;
        RECT 106.690 136.870 107.310 136.880 ;
        RECT 108.875 136.700 116.875 136.930 ;
        RECT 108.960 136.690 116.830 136.700 ;
        RECT 104.570 135.980 105.450 136.000 ;
        RECT 103.840 135.600 104.110 135.890 ;
        RECT 104.510 135.750 105.510 135.980 ;
        RECT 105.670 135.940 106.040 136.230 ;
        RECT 105.700 135.880 106.040 135.940 ;
        RECT 106.800 136.550 107.560 136.600 ;
        RECT 108.440 136.550 108.670 136.650 ;
        RECT 106.800 136.340 108.670 136.550 ;
        RECT 117.080 136.340 117.310 136.650 ;
        RECT 106.800 135.920 109.340 136.340 ;
        RECT 116.710 135.920 117.310 136.340 ;
        RECT 104.570 135.600 105.450 135.750 ;
        RECT 104.580 135.430 105.310 135.600 ;
        RECT 40.690 135.000 41.010 135.060 ;
        RECT 48.050 135.000 48.370 135.060 ;
        RECT 81.670 135.000 81.960 135.045 ;
        RECT 83.770 135.000 84.060 135.045 ;
        RECT 85.340 135.000 85.630 135.045 ;
        RECT 40.320 134.860 41.010 135.000 ;
        RECT 29.650 134.660 29.970 134.720 ;
        RECT 39.770 134.660 40.090 134.720 ;
        RECT 40.320 134.705 40.460 134.860 ;
        RECT 40.690 134.800 41.010 134.860 ;
        RECT 44.920 134.860 48.370 135.000 ;
        RECT 29.650 134.520 40.090 134.660 ;
        RECT 29.650 134.460 29.970 134.520 ;
        RECT 39.770 134.460 40.090 134.520 ;
        RECT 40.245 134.475 40.535 134.705 ;
        RECT 44.920 134.660 45.060 134.860 ;
        RECT 48.050 134.800 48.370 134.860 ;
        RECT 48.600 134.860 80.020 135.000 ;
        RECT 40.780 134.520 45.060 134.660 ;
        RECT 45.290 134.660 45.610 134.720 ;
        RECT 46.225 134.660 46.515 134.705 ;
        RECT 45.290 134.520 46.515 134.660 ;
        RECT 10.790 134.320 11.110 134.380 ;
        RECT 40.780 134.365 40.920 134.520 ;
        RECT 45.290 134.460 45.610 134.520 ;
        RECT 46.225 134.475 46.515 134.520 ;
        RECT 13.565 134.320 13.855 134.365 ;
        RECT 10.790 134.180 13.855 134.320 ;
        RECT 10.790 134.120 11.110 134.180 ;
        RECT 13.565 134.135 13.855 134.180 ;
        RECT 40.705 134.135 40.995 134.365 ;
        RECT 42.085 134.320 42.375 134.365 ;
        RECT 42.530 134.320 42.850 134.380 ;
        RECT 42.085 134.180 42.850 134.320 ;
        RECT 42.085 134.135 42.375 134.180 ;
        RECT 42.530 134.120 42.850 134.180 ;
        RECT 43.925 134.320 44.215 134.365 ;
        RECT 45.750 134.320 46.070 134.380 ;
        RECT 43.925 134.180 46.070 134.320 ;
        RECT 43.925 134.135 44.215 134.180 ;
        RECT 45.750 134.120 46.070 134.180 ;
        RECT 46.670 134.120 46.990 134.380 ;
        RECT 34.710 133.780 35.030 134.040 ;
        RECT 38.865 133.980 39.155 134.025 ;
        RECT 47.590 133.980 47.910 134.040 ;
        RECT 38.865 133.840 47.910 133.980 ;
        RECT 38.865 133.795 39.155 133.840 ;
        RECT 47.590 133.780 47.910 133.840 ;
        RECT 14.485 133.640 14.775 133.685 ;
        RECT 24.130 133.640 24.450 133.700 ;
        RECT 14.485 133.500 24.450 133.640 ;
        RECT 14.485 133.455 14.775 133.500 ;
        RECT 24.130 133.440 24.450 133.500 ;
        RECT 46.210 133.640 46.530 133.700 ;
        RECT 48.600 133.640 48.740 134.860 ;
        RECT 50.365 134.660 50.655 134.705 ;
        RECT 50.810 134.660 51.130 134.720 ;
        RECT 50.365 134.520 51.130 134.660 ;
        RECT 50.365 134.475 50.655 134.520 ;
        RECT 50.810 134.460 51.130 134.520 ;
        RECT 53.110 134.660 53.430 134.720 ;
        RECT 54.505 134.660 54.795 134.705 ;
        RECT 53.110 134.520 54.795 134.660 ;
        RECT 53.110 134.460 53.430 134.520 ;
        RECT 54.505 134.475 54.795 134.520 ;
        RECT 63.230 134.460 63.550 134.720 ;
        RECT 66.450 134.660 66.770 134.720 ;
        RECT 72.445 134.660 72.735 134.705 ;
        RECT 66.450 134.520 72.735 134.660 ;
        RECT 66.450 134.460 66.770 134.520 ;
        RECT 72.445 134.475 72.735 134.520 ;
        RECT 75.650 134.660 75.970 134.720 ;
        RECT 75.650 134.520 78.640 134.660 ;
        RECT 75.650 134.460 75.970 134.520 ;
        RECT 52.650 134.320 52.970 134.380 ;
        RECT 58.645 134.320 58.935 134.365 ;
        RECT 52.650 134.180 58.935 134.320 ;
        RECT 52.650 134.120 52.970 134.180 ;
        RECT 58.645 134.135 58.935 134.180 ;
        RECT 62.770 134.120 63.090 134.380 ;
        RECT 68.305 134.135 68.595 134.365 ;
        RECT 53.585 133.980 53.875 134.025 ;
        RECT 57.250 133.980 57.570 134.040 ;
        RECT 53.585 133.840 57.570 133.980 ;
        RECT 68.380 133.980 68.520 134.135 ;
        RECT 71.510 134.120 71.830 134.380 ;
        RECT 77.030 134.320 77.350 134.380 ;
        RECT 78.500 134.365 78.640 134.520 ;
        RECT 78.870 134.460 79.190 134.720 ;
        RECT 77.965 134.320 78.255 134.365 ;
        RECT 77.030 134.180 78.255 134.320 ;
        RECT 77.030 134.120 77.350 134.180 ;
        RECT 77.965 134.135 78.255 134.180 ;
        RECT 78.425 134.135 78.715 134.365 ;
        RECT 76.570 133.980 76.890 134.040 ;
        RECT 68.380 133.840 76.890 133.980 ;
        RECT 53.585 133.795 53.875 133.840 ;
        RECT 57.250 133.780 57.570 133.840 ;
        RECT 76.570 133.780 76.890 133.840 ;
        RECT 46.210 133.500 48.740 133.640 ;
        RECT 54.045 133.640 54.335 133.685 ;
        RECT 55.885 133.640 56.175 133.685 ;
        RECT 54.045 133.500 56.175 133.640 ;
        RECT 46.210 133.440 46.530 133.500 ;
        RECT 54.045 133.455 54.335 133.500 ;
        RECT 55.885 133.455 56.175 133.500 ;
        RECT 66.465 133.640 66.755 133.685 ;
        RECT 66.910 133.640 67.230 133.700 ;
        RECT 66.465 133.500 67.230 133.640 ;
        RECT 66.465 133.455 66.755 133.500 ;
        RECT 66.910 133.440 67.230 133.500 ;
        RECT 67.370 133.440 67.690 133.700 ;
        RECT 67.830 133.640 68.150 133.700 ;
        RECT 68.765 133.640 69.055 133.685 ;
        RECT 67.830 133.500 69.055 133.640 ;
        RECT 67.830 133.440 68.150 133.500 ;
        RECT 68.765 133.455 69.055 133.500 ;
        RECT 73.350 133.640 73.670 133.700 ;
        RECT 75.665 133.640 75.955 133.685 ;
        RECT 73.350 133.500 75.955 133.640 ;
        RECT 73.350 133.440 73.670 133.500 ;
        RECT 75.665 133.455 75.955 133.500 ;
        RECT 77.045 133.640 77.335 133.685 ;
        RECT 78.960 133.640 79.100 134.460 ;
        RECT 79.880 134.365 80.020 134.860 ;
        RECT 81.670 134.860 85.630 135.000 ;
        RECT 81.670 134.815 81.960 134.860 ;
        RECT 83.770 134.815 84.060 134.860 ;
        RECT 85.340 134.815 85.630 134.860 ;
        RECT 81.170 134.460 81.490 134.720 ;
        RECT 82.065 134.660 82.355 134.705 ;
        RECT 83.255 134.660 83.545 134.705 ;
        RECT 85.775 134.660 86.065 134.705 ;
        RECT 82.065 134.520 86.065 134.660 ;
        RECT 82.065 134.475 82.355 134.520 ;
        RECT 83.255 134.475 83.545 134.520 ;
        RECT 85.775 134.475 86.065 134.520 ;
        RECT 79.345 134.135 79.635 134.365 ;
        RECT 79.805 134.135 80.095 134.365 ;
        RECT 77.045 133.500 79.100 133.640 ;
        RECT 79.420 133.640 79.560 134.135 ;
        RECT 82.550 134.025 82.870 134.040 ;
        RECT 82.520 133.795 82.870 134.025 ;
        RECT 82.550 133.780 82.870 133.795 ;
        RECT 84.390 133.640 84.710 133.700 ;
        RECT 79.420 133.500 84.710 133.640 ;
        RECT 77.045 133.455 77.335 133.500 ;
        RECT 84.390 133.440 84.710 133.500 ;
        RECT 87.610 133.640 87.930 133.700 ;
        RECT 88.085 133.640 88.375 133.685 ;
        RECT 87.610 133.500 88.375 133.640 ;
        RECT 87.610 133.440 87.930 133.500 ;
        RECT 88.085 133.455 88.375 133.500 ;
        RECT 12.100 132.820 89.840 133.300 ;
        RECT 16.770 132.620 17.090 132.680 ;
        RECT 29.650 132.620 29.970 132.680 ;
        RECT 16.770 132.480 29.970 132.620 ;
        RECT 16.770 132.420 17.090 132.480 ;
        RECT 29.650 132.420 29.970 132.480 ;
        RECT 44.830 132.620 45.150 132.680 ;
        RECT 47.130 132.620 47.450 132.680 ;
        RECT 50.365 132.620 50.655 132.665 ;
        RECT 44.830 132.480 46.900 132.620 ;
        RECT 44.830 132.420 45.150 132.480 ;
        RECT 24.590 132.280 24.910 132.340 ;
        RECT 30.110 132.280 30.430 132.340 ;
        RECT 45.750 132.280 46.070 132.340 ;
        RECT 24.590 132.140 26.660 132.280 ;
        RECT 24.590 132.080 24.910 132.140 ;
        RECT 26.520 132.000 26.660 132.140 ;
        RECT 27.440 132.140 30.430 132.280 ;
        RECT 16.325 131.940 16.615 131.985 ;
        RECT 20.910 131.940 21.230 132.000 ;
        RECT 23.670 131.940 23.990 132.000 ;
        RECT 16.325 131.800 23.990 131.940 ;
        RECT 16.325 131.755 16.615 131.800 ;
        RECT 20.910 131.740 21.230 131.800 ;
        RECT 23.670 131.740 23.990 131.800 ;
        RECT 24.130 131.740 24.450 132.000 ;
        RECT 26.430 131.740 26.750 132.000 ;
        RECT 27.440 131.985 27.580 132.140 ;
        RECT 30.110 132.080 30.430 132.140 ;
        RECT 41.700 132.140 46.070 132.280 ;
        RECT 46.760 132.280 46.900 132.480 ;
        RECT 47.130 132.480 50.655 132.620 ;
        RECT 47.130 132.420 47.450 132.480 ;
        RECT 50.365 132.435 50.655 132.480 ;
        RECT 53.110 132.420 53.430 132.680 ;
        RECT 63.230 132.420 63.550 132.680 ;
        RECT 71.065 132.620 71.355 132.665 ;
        RECT 71.510 132.620 71.830 132.680 ;
        RECT 71.065 132.480 71.830 132.620 ;
        RECT 71.065 132.435 71.355 132.480 ;
        RECT 71.510 132.420 71.830 132.480 ;
        RECT 73.350 132.420 73.670 132.680 ;
        RECT 74.270 132.620 74.590 132.680 ;
        RECT 85.310 132.620 85.630 132.680 ;
        RECT 74.270 132.480 85.630 132.620 ;
        RECT 74.270 132.420 74.590 132.480 ;
        RECT 85.310 132.420 85.630 132.480 ;
        RECT 46.760 132.140 48.280 132.280 ;
        RECT 27.365 131.755 27.655 131.985 ;
        RECT 29.665 131.940 29.955 131.985 ;
        RECT 27.900 131.800 29.955 131.940 ;
        RECT 15.850 131.645 16.170 131.660 ;
        RECT 15.740 131.415 16.170 131.645 ;
        RECT 18.165 131.600 18.455 131.645 ;
        RECT 19.530 131.600 19.850 131.660 ;
        RECT 18.165 131.460 19.850 131.600 ;
        RECT 18.165 131.415 18.455 131.460 ;
        RECT 15.850 131.400 16.170 131.415 ;
        RECT 19.530 131.400 19.850 131.460 ;
        RECT 25.970 131.400 26.290 131.660 ;
        RECT 25.510 131.260 25.830 131.320 ;
        RECT 27.900 131.260 28.040 131.800 ;
        RECT 29.665 131.755 29.955 131.800 ;
        RECT 32.885 131.755 33.175 131.985 ;
        RECT 33.805 131.755 34.095 131.985 ;
        RECT 30.585 131.600 30.875 131.645 ;
        RECT 31.030 131.600 31.350 131.660 ;
        RECT 30.585 131.460 31.350 131.600 ;
        RECT 30.585 131.415 30.875 131.460 ;
        RECT 31.030 131.400 31.350 131.460 ;
        RECT 25.510 131.120 28.040 131.260 ;
        RECT 28.285 131.260 28.575 131.305 ;
        RECT 29.650 131.260 29.970 131.320 ;
        RECT 28.285 131.120 29.970 131.260 ;
        RECT 32.960 131.260 33.100 131.755 ;
        RECT 33.880 131.600 34.020 131.755 ;
        RECT 34.710 131.740 35.030 132.000 ;
        RECT 35.630 131.940 35.950 132.000 ;
        RECT 38.405 131.940 38.695 131.985 ;
        RECT 35.630 131.800 38.695 131.940 ;
        RECT 35.630 131.740 35.950 131.800 ;
        RECT 38.405 131.755 38.695 131.800 ;
        RECT 39.325 131.755 39.615 131.985 ;
        RECT 40.705 131.940 40.995 131.985 ;
        RECT 41.700 131.940 41.840 132.140 ;
        RECT 45.750 132.080 46.070 132.140 ;
        RECT 42.070 131.985 42.390 132.000 ;
        RECT 40.705 131.800 41.840 131.940 ;
        RECT 40.705 131.755 40.995 131.800 ;
        RECT 42.040 131.755 42.390 131.985 ;
        RECT 48.140 131.940 48.280 132.140 ;
        RECT 49.890 132.080 50.210 132.340 ;
        RECT 81.630 132.280 81.950 132.340 ;
        RECT 87.610 132.280 87.930 132.340 ;
        RECT 78.960 132.140 81.950 132.280 ;
        RECT 52.665 131.940 52.955 131.985 ;
        RECT 48.140 131.800 52.955 131.940 ;
        RECT 52.665 131.755 52.955 131.800 ;
        RECT 54.950 131.940 55.270 132.000 ;
        RECT 56.345 131.940 56.635 131.985 ;
        RECT 54.950 131.800 56.635 131.940 ;
        RECT 38.865 131.600 39.155 131.645 ;
        RECT 33.880 131.460 39.155 131.600 ;
        RECT 38.865 131.415 39.155 131.460 ;
        RECT 35.630 131.260 35.950 131.320 ;
        RECT 37.470 131.260 37.790 131.320 ;
        RECT 32.960 131.120 37.790 131.260 ;
        RECT 25.510 131.060 25.830 131.120 ;
        RECT 28.285 131.075 28.575 131.120 ;
        RECT 29.650 131.060 29.970 131.120 ;
        RECT 35.630 131.060 35.950 131.120 ;
        RECT 37.470 131.060 37.790 131.120 ;
        RECT 37.930 131.260 38.250 131.320 ;
        RECT 39.400 131.260 39.540 131.755 ;
        RECT 42.070 131.740 42.390 131.755 ;
        RECT 54.950 131.740 55.270 131.800 ;
        RECT 56.345 131.755 56.635 131.800 ;
        RECT 57.680 131.940 57.970 131.985 ;
        RECT 62.770 131.940 63.090 132.000 ;
        RECT 57.680 131.800 63.090 131.940 ;
        RECT 57.680 131.755 57.970 131.800 ;
        RECT 62.770 131.740 63.090 131.800 ;
        RECT 64.610 131.940 64.930 132.000 ;
        RECT 65.445 131.940 65.735 131.985 ;
        RECT 64.610 131.800 65.735 131.940 ;
        RECT 64.610 131.740 64.930 131.800 ;
        RECT 65.445 131.755 65.735 131.800 ;
        RECT 68.290 131.940 68.610 132.000 ;
        RECT 73.825 131.940 74.115 131.985 ;
        RECT 75.190 131.940 75.510 132.000 ;
        RECT 68.290 131.800 69.440 131.940 ;
        RECT 68.290 131.740 68.610 131.800 ;
        RECT 41.585 131.600 41.875 131.645 ;
        RECT 42.775 131.600 43.065 131.645 ;
        RECT 45.295 131.600 45.585 131.645 ;
        RECT 41.585 131.460 45.585 131.600 ;
        RECT 41.585 131.415 41.875 131.460 ;
        RECT 42.775 131.415 43.065 131.460 ;
        RECT 45.295 131.415 45.585 131.460 ;
        RECT 48.050 131.600 48.370 131.660 ;
        RECT 51.285 131.600 51.575 131.645 ;
        RECT 53.110 131.600 53.430 131.660 ;
        RECT 48.050 131.460 53.430 131.600 ;
        RECT 48.050 131.400 48.370 131.460 ;
        RECT 51.285 131.415 51.575 131.460 ;
        RECT 53.110 131.400 53.430 131.460 ;
        RECT 57.225 131.600 57.515 131.645 ;
        RECT 58.415 131.600 58.705 131.645 ;
        RECT 60.935 131.600 61.225 131.645 ;
        RECT 57.225 131.460 61.225 131.600 ;
        RECT 57.225 131.415 57.515 131.460 ;
        RECT 58.415 131.415 58.705 131.460 ;
        RECT 60.935 131.415 61.225 131.460 ;
        RECT 64.150 131.400 64.470 131.660 ;
        RECT 65.045 131.600 65.335 131.645 ;
        RECT 66.235 131.600 66.525 131.645 ;
        RECT 68.755 131.600 69.045 131.645 ;
        RECT 65.045 131.460 69.045 131.600 ;
        RECT 65.045 131.415 65.335 131.460 ;
        RECT 66.235 131.415 66.525 131.460 ;
        RECT 68.755 131.415 69.045 131.460 ;
        RECT 37.930 131.120 39.540 131.260 ;
        RECT 41.190 131.260 41.480 131.305 ;
        RECT 43.290 131.260 43.580 131.305 ;
        RECT 44.860 131.260 45.150 131.305 ;
        RECT 41.190 131.120 45.150 131.260 ;
        RECT 37.930 131.060 38.250 131.120 ;
        RECT 41.190 131.075 41.480 131.120 ;
        RECT 43.290 131.075 43.580 131.120 ;
        RECT 44.860 131.075 45.150 131.120 ;
        RECT 56.830 131.260 57.120 131.305 ;
        RECT 58.930 131.260 59.220 131.305 ;
        RECT 60.500 131.260 60.790 131.305 ;
        RECT 56.830 131.120 60.790 131.260 ;
        RECT 56.830 131.075 57.120 131.120 ;
        RECT 58.930 131.075 59.220 131.120 ;
        RECT 60.500 131.075 60.790 131.120 ;
        RECT 64.650 131.260 64.940 131.305 ;
        RECT 66.750 131.260 67.040 131.305 ;
        RECT 68.320 131.260 68.610 131.305 ;
        RECT 64.650 131.120 68.610 131.260 ;
        RECT 69.300 131.260 69.440 131.800 ;
        RECT 73.825 131.800 75.510 131.940 ;
        RECT 73.825 131.755 74.115 131.800 ;
        RECT 75.190 131.740 75.510 131.800 ;
        RECT 77.045 131.755 77.335 131.985 ;
        RECT 77.505 131.940 77.795 131.985 ;
        RECT 77.950 131.940 78.270 132.000 ;
        RECT 77.505 131.800 78.270 131.940 ;
        RECT 77.505 131.755 77.795 131.800 ;
        RECT 69.670 131.600 69.990 131.660 ;
        RECT 74.285 131.600 74.575 131.645 ;
        RECT 69.670 131.460 74.575 131.600 ;
        RECT 77.120 131.600 77.260 131.755 ;
        RECT 77.950 131.740 78.270 131.800 ;
        RECT 78.410 131.740 78.730 132.000 ;
        RECT 78.960 131.985 79.100 132.140 ;
        RECT 81.630 132.080 81.950 132.140 ;
        RECT 82.180 132.140 87.930 132.280 ;
        RECT 78.885 131.755 79.175 131.985 ;
        RECT 79.330 131.740 79.650 132.000 ;
        RECT 81.170 131.740 81.490 132.000 ;
        RECT 82.180 131.940 82.320 132.140 ;
        RECT 87.610 132.080 87.930 132.140 ;
        RECT 81.720 131.800 82.320 131.940 ;
        RECT 82.520 131.940 82.810 131.985 ;
        RECT 83.930 131.940 84.250 132.000 ;
        RECT 82.520 131.800 84.250 131.940 ;
        RECT 81.720 131.600 81.860 131.800 ;
        RECT 82.520 131.755 82.810 131.800 ;
        RECT 83.930 131.740 84.250 131.800 ;
        RECT 100.010 131.720 100.780 135.360 ;
        RECT 102.460 134.310 105.310 135.430 ;
        RECT 105.700 135.130 106.050 135.880 ;
        RECT 106.800 135.760 108.670 135.920 ;
        RECT 106.800 135.710 107.560 135.760 ;
        RECT 108.440 135.690 108.670 135.760 ;
        RECT 117.080 135.690 117.310 135.920 ;
        RECT 108.875 135.410 116.875 135.640 ;
        RECT 105.700 135.070 105.990 135.130 ;
        RECT 105.610 134.950 105.990 135.070 ;
        RECT 108.970 135.010 116.830 135.410 ;
        RECT 117.640 135.010 118.600 144.490 ;
        RECT 119.930 144.620 120.770 146.750 ;
        RECT 126.430 146.330 127.680 146.770 ;
        RECT 137.600 146.750 138.460 148.920 ;
        RECT 124.370 146.320 129.610 146.330 ;
        RECT 121.420 146.220 136.720 146.320 ;
        RECT 121.420 146.210 136.755 146.220 ;
        RECT 121.380 146.090 136.755 146.210 ;
        RECT 121.380 145.980 125.380 146.090 ;
        RECT 126.430 146.010 128.170 146.090 ;
        RECT 128.750 146.010 136.755 146.090 ;
        RECT 126.430 145.930 127.680 146.010 ;
        RECT 128.755 145.990 136.755 146.010 ;
        RECT 120.990 145.680 121.220 145.930 ;
        RECT 125.540 145.790 125.770 145.930 ;
        RECT 128.320 145.790 128.550 145.940 ;
        RECT 125.540 145.680 128.550 145.790 ;
        RECT 136.960 145.680 137.190 145.940 ;
        RECT 120.990 145.240 137.190 145.680 ;
        RECT 120.990 144.970 121.220 145.240 ;
        RECT 125.540 145.210 137.190 145.240 ;
        RECT 125.540 145.120 128.550 145.210 ;
        RECT 125.540 144.970 125.770 145.120 ;
        RECT 128.320 144.980 128.550 145.120 ;
        RECT 136.960 144.980 137.190 145.210 ;
        RECT 121.380 144.690 125.380 144.920 ;
        RECT 128.755 144.710 136.755 144.930 ;
        RECT 137.520 144.710 138.480 146.750 ;
        RECT 128.755 144.700 138.480 144.710 ;
        RECT 121.380 144.620 125.370 144.690 ;
        RECT 119.930 144.510 125.370 144.620 ;
        RECT 128.810 144.540 138.480 144.700 ;
        RECT 119.930 144.420 123.060 144.510 ;
        RECT 136.550 144.490 138.480 144.540 ;
        RECT 119.930 141.150 120.770 144.420 ;
        RECT 124.410 143.960 129.660 143.970 ;
        RECT 124.410 143.850 136.720 143.960 ;
        RECT 121.440 143.790 136.720 143.850 ;
        RECT 121.440 143.780 136.755 143.790 ;
        RECT 121.380 143.650 136.755 143.780 ;
        RECT 121.380 143.640 126.540 143.650 ;
        RECT 121.380 143.550 125.380 143.640 ;
        RECT 128.755 143.560 136.755 143.650 ;
        RECT 128.840 143.550 136.730 143.560 ;
        RECT 120.990 143.190 121.220 143.500 ;
        RECT 121.440 143.190 125.340 143.550 ;
        RECT 125.540 143.190 125.770 143.500 ;
        RECT 120.990 141.850 125.770 143.190 ;
        RECT 120.990 141.540 121.220 141.850 ;
        RECT 125.540 141.540 125.770 141.850 ;
        RECT 128.320 142.970 128.550 143.510 ;
        RECT 129.360 142.970 130.370 143.000 ;
        RECT 136.960 142.970 137.190 143.510 ;
        RECT 128.320 142.070 137.190 142.970 ;
        RECT 128.320 141.550 128.550 142.070 ;
        RECT 129.360 142.000 130.370 142.070 ;
        RECT 136.960 141.550 137.190 142.070 ;
        RECT 121.380 141.260 125.380 141.490 ;
        RECT 128.755 141.270 136.755 141.500 ;
        RECT 119.930 141.110 121.060 141.150 ;
        RECT 119.930 141.030 121.300 141.110 ;
        RECT 121.670 141.040 125.330 141.260 ;
        RECT 121.670 141.030 123.110 141.040 ;
        RECT 119.930 140.990 123.110 141.030 ;
        RECT 119.930 140.900 122.620 140.990 ;
        RECT 128.820 140.980 136.710 141.270 ;
        RECT 119.930 140.840 121.950 140.900 ;
        RECT 119.930 140.790 121.700 140.840 ;
        RECT 119.930 137.450 120.770 140.790 ;
        RECT 128.810 140.490 136.730 140.500 ;
        RECT 125.040 140.480 136.730 140.490 ;
        RECT 121.420 140.360 136.730 140.480 ;
        RECT 121.420 140.350 136.755 140.360 ;
        RECT 121.380 140.230 136.755 140.350 ;
        RECT 121.380 140.120 125.380 140.230 ;
        RECT 120.990 139.780 121.220 140.070 ;
        RECT 121.440 139.780 125.330 140.120 ;
        RECT 125.540 139.780 125.770 140.070 ;
        RECT 120.990 138.410 125.770 139.780 ;
        RECT 120.990 138.110 121.220 138.410 ;
        RECT 125.540 138.110 125.770 138.410 ;
        RECT 121.380 137.830 125.380 138.060 ;
        RECT 121.630 137.600 125.200 137.830 ;
        RECT 121.630 137.450 125.320 137.600 ;
        RECT 119.930 137.170 125.320 137.450 ;
        RECT 126.570 137.280 127.190 140.230 ;
        RECT 128.755 140.130 136.755 140.230 ;
        RECT 128.810 140.120 136.730 140.130 ;
        RECT 128.320 139.420 128.550 140.080 ;
        RECT 129.330 139.420 130.330 139.510 ;
        RECT 136.960 139.420 137.190 140.080 ;
        RECT 128.320 138.600 137.190 139.420 ;
        RECT 128.320 138.120 128.550 138.600 ;
        RECT 129.330 138.510 130.330 138.600 ;
        RECT 136.960 138.120 137.190 138.600 ;
        RECT 128.755 137.840 136.755 138.070 ;
        RECT 119.930 136.710 125.330 137.170 ;
        RECT 119.930 135.370 121.930 136.710 ;
        RECT 123.680 136.700 125.330 136.710 ;
        RECT 122.370 135.430 123.370 136.150 ;
        RECT 123.680 135.890 123.990 136.700 ;
        RECT 124.450 136.420 125.330 136.700 ;
        RECT 125.570 136.880 127.190 137.280 ;
        RECT 128.840 136.930 136.710 137.840 ;
        RECT 124.390 136.190 125.390 136.420 ;
        RECT 125.570 136.230 125.920 136.880 ;
        RECT 126.570 136.870 127.190 136.880 ;
        RECT 128.755 136.700 136.755 136.930 ;
        RECT 128.840 136.690 136.710 136.700 ;
        RECT 124.450 135.980 125.330 136.000 ;
        RECT 123.720 135.600 123.990 135.890 ;
        RECT 124.390 135.750 125.390 135.980 ;
        RECT 125.550 135.940 125.920 136.230 ;
        RECT 125.580 135.880 125.920 135.940 ;
        RECT 126.680 136.550 127.440 136.600 ;
        RECT 128.320 136.550 128.550 136.650 ;
        RECT 126.680 136.340 128.550 136.550 ;
        RECT 136.960 136.340 137.190 136.650 ;
        RECT 126.680 135.920 129.220 136.340 ;
        RECT 136.590 135.920 137.190 136.340 ;
        RECT 124.450 135.600 125.330 135.750 ;
        RECT 124.460 135.430 125.190 135.600 ;
        RECT 102.400 134.080 105.400 134.310 ;
        RECT 105.610 134.120 105.950 134.950 ;
        RECT 107.960 134.940 118.600 135.010 ;
        RECT 102.450 134.050 105.310 134.080 ;
        RECT 102.450 134.030 103.620 134.050 ;
        RECT 104.580 134.040 105.310 134.050 ;
        RECT 102.400 133.640 105.400 133.870 ;
        RECT 105.605 133.830 105.950 134.120 ;
        RECT 106.140 133.900 118.600 134.940 ;
        RECT 120.000 135.360 121.930 135.370 ;
        RECT 106.140 133.880 118.560 133.900 ;
        RECT 105.610 133.720 105.950 133.830 ;
        RECT 106.180 133.870 111.850 133.880 ;
        RECT 112.850 133.870 118.560 133.880 ;
        RECT 102.490 133.470 105.350 133.640 ;
        RECT 106.180 133.470 106.610 133.870 ;
        RECT 102.460 133.100 106.610 133.470 ;
        RECT 77.120 131.460 81.860 131.600 ;
        RECT 82.065 131.600 82.355 131.645 ;
        RECT 83.255 131.600 83.545 131.645 ;
        RECT 85.775 131.600 86.065 131.645 ;
        RECT 82.065 131.460 86.065 131.600 ;
        RECT 69.670 131.400 69.990 131.460 ;
        RECT 74.285 131.415 74.575 131.460 ;
        RECT 82.065 131.415 82.355 131.460 ;
        RECT 83.255 131.415 83.545 131.460 ;
        RECT 85.775 131.415 86.065 131.460 ;
        RECT 69.300 131.120 75.880 131.260 ;
        RECT 64.650 131.075 64.940 131.120 ;
        RECT 66.750 131.075 67.040 131.120 ;
        RECT 68.320 131.075 68.610 131.120 ;
        RECT 14.945 130.920 15.235 130.965 ;
        RECT 15.390 130.920 15.710 130.980 ;
        RECT 14.945 130.780 15.710 130.920 ;
        RECT 14.945 130.735 15.235 130.780 ;
        RECT 15.390 130.720 15.710 130.780 ;
        RECT 23.670 130.920 23.990 130.980 ;
        RECT 25.065 130.920 25.355 130.965 ;
        RECT 26.890 130.920 27.210 130.980 ;
        RECT 23.670 130.780 27.210 130.920 ;
        RECT 23.670 130.720 23.990 130.780 ;
        RECT 25.065 130.735 25.355 130.780 ;
        RECT 26.890 130.720 27.210 130.780 ;
        RECT 28.745 130.920 29.035 130.965 ;
        RECT 30.110 130.920 30.430 130.980 ;
        RECT 28.745 130.780 30.430 130.920 ;
        RECT 28.745 130.735 29.035 130.780 ;
        RECT 30.110 130.720 30.430 130.780 ;
        RECT 33.790 130.720 34.110 130.980 ;
        RECT 45.290 130.920 45.610 130.980 ;
        RECT 47.605 130.920 47.895 130.965 ;
        RECT 45.290 130.780 47.895 130.920 ;
        RECT 45.290 130.720 45.610 130.780 ;
        RECT 47.605 130.735 47.895 130.780 ;
        RECT 48.065 130.920 48.355 130.965 ;
        RECT 48.970 130.920 49.290 130.980 ;
        RECT 48.065 130.780 49.290 130.920 ;
        RECT 48.065 130.735 48.355 130.780 ;
        RECT 48.970 130.720 49.290 130.780 ;
        RECT 63.690 130.920 64.010 130.980 ;
        RECT 70.590 130.920 70.910 130.980 ;
        RECT 63.690 130.780 70.910 130.920 ;
        RECT 63.690 130.720 64.010 130.780 ;
        RECT 70.590 130.720 70.910 130.780 ;
        RECT 71.510 130.720 71.830 130.980 ;
        RECT 75.740 130.920 75.880 131.120 ;
        RECT 76.110 131.060 76.430 131.320 ;
        RECT 77.030 131.260 77.350 131.320 ;
        RECT 78.410 131.260 78.730 131.320 ;
        RECT 77.030 131.120 78.730 131.260 ;
        RECT 77.030 131.060 77.350 131.120 ;
        RECT 78.410 131.060 78.730 131.120 ;
        RECT 80.250 131.260 80.570 131.320 ;
        RECT 81.170 131.260 81.490 131.320 ;
        RECT 80.250 131.120 81.490 131.260 ;
        RECT 80.250 131.060 80.570 131.120 ;
        RECT 81.170 131.060 81.490 131.120 ;
        RECT 81.670 131.260 81.960 131.305 ;
        RECT 83.770 131.260 84.060 131.305 ;
        RECT 85.340 131.260 85.630 131.305 ;
        RECT 81.670 131.120 85.630 131.260 ;
        RECT 81.670 131.075 81.960 131.120 ;
        RECT 83.770 131.075 84.060 131.120 ;
        RECT 85.340 131.075 85.630 131.120 ;
        RECT 79.790 130.920 80.110 130.980 ;
        RECT 75.740 130.780 80.110 130.920 ;
        RECT 79.790 130.720 80.110 130.780 ;
        RECT 80.725 130.920 81.015 130.965 ;
        RECT 82.550 130.920 82.870 130.980 ;
        RECT 80.725 130.780 82.870 130.920 ;
        RECT 80.725 130.735 81.015 130.780 ;
        RECT 82.550 130.720 82.870 130.780 ;
        RECT 83.010 130.920 83.330 130.980 ;
        RECT 84.850 130.920 85.170 130.980 ;
        RECT 83.010 130.780 85.170 130.920 ;
        RECT 83.010 130.720 83.330 130.780 ;
        RECT 84.850 130.720 85.170 130.780 ;
        RECT 85.770 130.920 86.090 130.980 ;
        RECT 88.085 130.920 88.375 130.965 ;
        RECT 85.770 130.780 88.375 130.920 ;
        RECT 85.770 130.720 86.090 130.780 ;
        RECT 88.085 130.735 88.375 130.780 ;
        RECT 12.100 130.100 89.840 130.580 ;
        RECT 15.850 129.900 16.170 129.960 ;
        RECT 21.385 129.900 21.675 129.945 ;
        RECT 15.850 129.760 21.675 129.900 ;
        RECT 15.850 129.700 16.170 129.760 ;
        RECT 21.385 129.715 21.675 129.760 ;
        RECT 27.810 129.900 28.130 129.960 ;
        RECT 31.030 129.900 31.350 129.960 ;
        RECT 27.810 129.760 31.350 129.900 ;
        RECT 27.810 129.700 28.130 129.760 ;
        RECT 31.030 129.700 31.350 129.760 ;
        RECT 33.330 129.900 33.650 129.960 ;
        RECT 37.470 129.900 37.790 129.960 ;
        RECT 39.785 129.900 40.075 129.945 ;
        RECT 33.330 129.760 37.240 129.900 ;
        RECT 33.330 129.700 33.650 129.760 ;
        RECT 14.510 129.560 14.800 129.605 ;
        RECT 16.610 129.560 16.900 129.605 ;
        RECT 18.180 129.560 18.470 129.605 ;
        RECT 14.510 129.420 18.470 129.560 ;
        RECT 14.510 129.375 14.800 129.420 ;
        RECT 16.610 129.375 16.900 129.420 ;
        RECT 18.180 129.375 18.470 129.420 ;
        RECT 25.985 129.560 26.275 129.605 ;
        RECT 26.430 129.560 26.750 129.620 ;
        RECT 25.985 129.420 26.750 129.560 ;
        RECT 31.120 129.560 31.260 129.700 ;
        RECT 37.100 129.560 37.240 129.760 ;
        RECT 37.470 129.760 40.075 129.900 ;
        RECT 37.470 129.700 37.790 129.760 ;
        RECT 39.785 129.715 40.075 129.760 ;
        RECT 42.070 129.900 42.390 129.960 ;
        RECT 42.545 129.900 42.835 129.945 ;
        RECT 42.070 129.760 42.835 129.900 ;
        RECT 42.070 129.700 42.390 129.760 ;
        RECT 42.545 129.715 42.835 129.760 ;
        RECT 43.465 129.900 43.755 129.945 ;
        RECT 50.810 129.900 51.130 129.960 ;
        RECT 43.465 129.760 51.130 129.900 ;
        RECT 43.465 129.715 43.755 129.760 ;
        RECT 50.810 129.700 51.130 129.760 ;
        RECT 57.250 129.700 57.570 129.960 ;
        RECT 57.710 129.900 58.030 129.960 ;
        RECT 60.010 129.900 60.330 129.960 ;
        RECT 67.830 129.900 68.150 129.960 ;
        RECT 57.710 129.760 60.330 129.900 ;
        RECT 57.710 129.700 58.030 129.760 ;
        RECT 60.010 129.700 60.330 129.760 ;
        RECT 61.480 129.760 68.150 129.900 ;
        RECT 46.210 129.560 46.500 129.605 ;
        RECT 47.780 129.560 48.070 129.605 ;
        RECT 49.880 129.560 50.170 129.605 ;
        RECT 61.480 129.560 61.620 129.760 ;
        RECT 67.830 129.700 68.150 129.760 ;
        RECT 72.430 129.900 72.750 129.960 ;
        RECT 77.950 129.900 78.270 129.960 ;
        RECT 81.170 129.900 81.490 129.960 ;
        RECT 72.430 129.760 73.580 129.900 ;
        RECT 72.430 129.700 72.750 129.760 ;
        RECT 31.120 129.420 36.780 129.560 ;
        RECT 37.100 129.420 39.080 129.560 ;
        RECT 25.985 129.375 26.275 129.420 ;
        RECT 26.430 129.360 26.750 129.420 ;
        RECT 14.905 129.220 15.195 129.265 ;
        RECT 16.095 129.220 16.385 129.265 ;
        RECT 18.615 129.220 18.905 129.265 ;
        RECT 21.830 129.220 22.150 129.280 ;
        RECT 29.665 129.220 29.955 129.265 ;
        RECT 14.905 129.080 18.905 129.220 ;
        RECT 14.905 129.035 15.195 129.080 ;
        RECT 16.095 129.035 16.385 129.080 ;
        RECT 18.615 129.035 18.905 129.080 ;
        RECT 21.000 129.080 29.955 129.220 ;
        RECT 13.550 128.880 13.870 128.940 ;
        RECT 15.390 128.925 15.710 128.940 ;
        RECT 14.025 128.880 14.315 128.925 ;
        RECT 15.360 128.880 15.710 128.925 ;
        RECT 13.550 128.740 14.315 128.880 ;
        RECT 15.195 128.740 15.710 128.880 ;
        RECT 13.550 128.680 13.870 128.740 ;
        RECT 14.025 128.695 14.315 128.740 ;
        RECT 15.360 128.695 15.710 128.740 ;
        RECT 15.390 128.680 15.710 128.695 ;
        RECT 16.770 128.880 17.090 128.940 ;
        RECT 21.000 128.880 21.140 129.080 ;
        RECT 21.830 129.020 22.150 129.080 ;
        RECT 29.665 129.035 29.955 129.080 ;
        RECT 16.770 128.740 21.140 128.880 ;
        RECT 16.770 128.680 17.090 128.740 ;
        RECT 21.370 128.680 21.690 128.940 ;
        RECT 22.290 128.680 22.610 128.940 ;
        RECT 23.670 128.925 23.990 128.940 ;
        RECT 23.670 128.695 24.125 128.925 ;
        RECT 23.670 128.680 23.990 128.695 ;
        RECT 24.590 128.680 24.910 128.940 ;
        RECT 25.525 128.695 25.815 128.925 ;
        RECT 26.445 128.695 26.735 128.925 ;
        RECT 26.890 128.880 27.210 128.940 ;
        RECT 27.365 128.880 27.655 128.925 ;
        RECT 26.890 128.740 27.655 128.880 ;
        RECT 29.740 128.880 29.880 129.035 ;
        RECT 31.490 129.020 31.810 129.280 ;
        RECT 32.090 129.220 32.380 129.265 ;
        RECT 33.790 129.220 34.110 129.280 ;
        RECT 32.090 129.080 34.110 129.220 ;
        RECT 32.090 129.035 32.380 129.080 ;
        RECT 33.790 129.020 34.110 129.080 ;
        RECT 34.725 129.220 35.015 129.265 ;
        RECT 36.090 129.220 36.410 129.280 ;
        RECT 34.725 129.080 36.410 129.220 ;
        RECT 34.725 129.035 35.015 129.080 ;
        RECT 33.345 128.880 33.635 128.925 ;
        RECT 34.800 128.880 34.940 129.035 ;
        RECT 36.090 129.020 36.410 129.080 ;
        RECT 29.740 128.740 33.635 128.880 ;
        RECT 19.530 128.540 19.850 128.600 ;
        RECT 22.380 128.540 22.520 128.680 ;
        RECT 19.530 128.400 22.520 128.540 ;
        RECT 22.765 128.540 23.055 128.585 ;
        RECT 23.210 128.540 23.530 128.600 ;
        RECT 25.600 128.540 25.740 128.695 ;
        RECT 22.765 128.400 25.740 128.540 ;
        RECT 19.530 128.340 19.850 128.400 ;
        RECT 22.765 128.355 23.055 128.400 ;
        RECT 23.210 128.340 23.530 128.400 ;
        RECT 20.925 128.200 21.215 128.245 ;
        RECT 21.830 128.200 22.150 128.260 ;
        RECT 20.925 128.060 22.150 128.200 ;
        RECT 20.925 128.015 21.215 128.060 ;
        RECT 21.830 128.000 22.150 128.060 ;
        RECT 22.290 128.200 22.610 128.260 ;
        RECT 26.520 128.200 26.660 128.695 ;
        RECT 26.890 128.680 27.210 128.740 ;
        RECT 27.365 128.695 27.655 128.740 ;
        RECT 33.345 128.695 33.635 128.740 ;
        RECT 33.880 128.740 34.940 128.880 ;
        RECT 36.640 128.880 36.780 129.420 ;
        RECT 38.940 128.925 39.080 129.420 ;
        RECT 46.210 129.420 50.170 129.560 ;
        RECT 46.210 129.375 46.500 129.420 ;
        RECT 47.780 129.375 48.070 129.420 ;
        RECT 49.880 129.375 50.170 129.420 ;
        RECT 55.500 129.420 61.620 129.560 ;
        RECT 61.850 129.560 62.170 129.620 ;
        RECT 66.450 129.560 66.770 129.620 ;
        RECT 61.850 129.420 66.770 129.560 ;
        RECT 41.625 129.220 41.915 129.265 ;
        RECT 43.450 129.220 43.770 129.280 ;
        RECT 41.625 129.080 43.770 129.220 ;
        RECT 41.625 129.035 41.915 129.080 ;
        RECT 43.450 129.020 43.770 129.080 ;
        RECT 45.775 129.220 46.065 129.265 ;
        RECT 48.295 129.220 48.585 129.265 ;
        RECT 49.485 129.220 49.775 129.265 ;
        RECT 45.775 129.080 49.775 129.220 ;
        RECT 45.775 129.035 46.065 129.080 ;
        RECT 48.295 129.035 48.585 129.080 ;
        RECT 49.485 129.035 49.775 129.080 ;
        RECT 38.405 128.880 38.695 128.925 ;
        RECT 36.640 128.740 38.695 128.880 ;
        RECT 31.045 128.540 31.335 128.585 ;
        RECT 32.410 128.540 32.730 128.600 ;
        RECT 33.880 128.540 34.020 128.740 ;
        RECT 38.405 128.695 38.695 128.740 ;
        RECT 38.865 128.695 39.155 128.925 ;
        RECT 41.165 128.880 41.455 128.925 ;
        RECT 44.370 128.880 44.690 128.940 ;
        RECT 41.165 128.740 44.690 128.880 ;
        RECT 41.165 128.695 41.455 128.740 ;
        RECT 44.370 128.680 44.690 128.740 ;
        RECT 48.970 128.925 49.290 128.940 ;
        RECT 48.970 128.880 49.320 128.925 ;
        RECT 50.365 128.880 50.655 128.925 ;
        RECT 52.650 128.880 52.970 128.940 ;
        RECT 55.500 128.925 55.640 129.420 ;
        RECT 61.850 129.360 62.170 129.420 ;
        RECT 66.450 129.360 66.770 129.420 ;
        RECT 69.210 129.560 69.500 129.605 ;
        RECT 70.780 129.560 71.070 129.605 ;
        RECT 72.880 129.560 73.170 129.605 ;
        RECT 69.210 129.420 73.170 129.560 ;
        RECT 69.210 129.375 69.500 129.420 ;
        RECT 70.780 129.375 71.070 129.420 ;
        RECT 72.880 129.375 73.170 129.420 ;
        RECT 59.550 129.020 59.870 129.280 ;
        RECT 60.010 129.020 60.330 129.280 ;
        RECT 63.690 129.220 64.010 129.280 ;
        RECT 67.370 129.220 67.690 129.280 ;
        RECT 73.440 129.265 73.580 129.760 ;
        RECT 77.950 129.760 81.490 129.900 ;
        RECT 77.950 129.700 78.270 129.760 ;
        RECT 81.170 129.700 81.490 129.760 ;
        RECT 83.930 129.700 84.250 129.960 ;
        RECT 84.390 129.700 84.710 129.960 ;
        RECT 100.010 129.620 100.880 131.720 ;
        RECT 106.550 131.330 107.800 131.770 ;
        RECT 117.700 131.750 118.560 133.870 ;
        RECT 120.000 131.810 120.770 135.360 ;
        RECT 122.340 134.310 125.190 135.430 ;
        RECT 125.580 135.130 125.930 135.880 ;
        RECT 126.680 135.760 128.550 135.920 ;
        RECT 126.680 135.710 127.440 135.760 ;
        RECT 128.320 135.690 128.550 135.760 ;
        RECT 136.960 135.690 137.190 135.920 ;
        RECT 128.755 135.410 136.755 135.640 ;
        RECT 125.580 135.070 125.870 135.130 ;
        RECT 125.490 134.950 125.870 135.070 ;
        RECT 128.850 135.010 136.710 135.410 ;
        RECT 137.520 135.010 138.480 144.490 ;
        RECT 122.280 134.080 125.280 134.310 ;
        RECT 125.490 134.120 125.830 134.950 ;
        RECT 127.840 134.940 138.480 135.010 ;
        RECT 122.330 134.050 125.190 134.080 ;
        RECT 122.330 134.030 123.500 134.050 ;
        RECT 124.460 134.040 125.190 134.050 ;
        RECT 122.280 133.640 125.280 133.870 ;
        RECT 125.485 133.830 125.830 134.120 ;
        RECT 126.020 133.900 138.480 134.940 ;
        RECT 139.930 146.720 140.700 150.360 ;
        RECT 142.420 149.310 145.270 150.430 ;
        RECT 145.660 150.130 146.010 150.880 ;
        RECT 146.760 150.760 148.630 150.920 ;
        RECT 146.760 150.710 147.520 150.760 ;
        RECT 148.400 150.690 148.630 150.760 ;
        RECT 157.040 150.690 157.270 150.920 ;
        RECT 148.835 150.410 156.835 150.640 ;
        RECT 145.660 150.070 145.950 150.130 ;
        RECT 145.570 149.950 145.950 150.070 ;
        RECT 148.930 150.010 156.790 150.410 ;
        RECT 157.600 150.010 158.560 159.490 ;
        RECT 142.360 149.080 145.360 149.310 ;
        RECT 145.570 149.120 145.910 149.950 ;
        RECT 147.920 149.940 158.560 150.010 ;
        RECT 142.410 149.050 145.270 149.080 ;
        RECT 142.410 149.030 143.580 149.050 ;
        RECT 144.540 149.040 145.270 149.050 ;
        RECT 142.360 148.640 145.360 148.870 ;
        RECT 145.565 148.830 145.910 149.120 ;
        RECT 146.100 148.900 158.560 149.940 ;
        RECT 146.100 148.880 158.500 148.900 ;
        RECT 145.570 148.720 145.910 148.830 ;
        RECT 146.140 148.870 151.810 148.880 ;
        RECT 152.810 148.870 158.500 148.880 ;
        RECT 142.450 148.470 145.310 148.640 ;
        RECT 146.140 148.470 146.570 148.870 ;
        RECT 142.420 148.100 146.570 148.470 ;
        RECT 139.930 144.620 140.790 146.720 ;
        RECT 146.460 146.330 147.710 146.770 ;
        RECT 157.640 146.750 158.500 148.870 ;
        RECT 144.400 146.320 149.640 146.330 ;
        RECT 141.450 146.220 156.750 146.320 ;
        RECT 141.450 146.210 156.785 146.220 ;
        RECT 141.410 146.090 156.785 146.210 ;
        RECT 141.410 145.980 145.410 146.090 ;
        RECT 146.460 146.010 148.200 146.090 ;
        RECT 148.780 146.010 156.785 146.090 ;
        RECT 146.460 145.930 147.710 146.010 ;
        RECT 148.785 145.990 156.785 146.010 ;
        RECT 141.020 145.680 141.250 145.930 ;
        RECT 145.570 145.790 145.800 145.930 ;
        RECT 148.350 145.790 148.580 145.940 ;
        RECT 145.570 145.680 148.580 145.790 ;
        RECT 156.990 145.680 157.220 145.940 ;
        RECT 141.020 145.240 157.220 145.680 ;
        RECT 141.020 144.970 141.250 145.240 ;
        RECT 145.570 145.210 157.220 145.240 ;
        RECT 145.570 145.120 148.580 145.210 ;
        RECT 145.570 144.970 145.800 145.120 ;
        RECT 148.350 144.980 148.580 145.120 ;
        RECT 156.990 144.980 157.220 145.210 ;
        RECT 141.410 144.690 145.410 144.920 ;
        RECT 148.785 144.710 156.785 144.930 ;
        RECT 157.550 144.710 158.510 146.750 ;
        RECT 148.785 144.700 158.510 144.710 ;
        RECT 141.410 144.620 145.400 144.690 ;
        RECT 139.930 144.510 145.400 144.620 ;
        RECT 148.840 144.540 158.510 144.700 ;
        RECT 139.930 144.420 143.090 144.510 ;
        RECT 156.580 144.490 158.510 144.540 ;
        RECT 139.930 141.150 140.790 144.420 ;
        RECT 144.440 143.960 149.690 143.970 ;
        RECT 144.440 143.850 156.750 143.960 ;
        RECT 141.470 143.790 156.750 143.850 ;
        RECT 141.470 143.780 156.785 143.790 ;
        RECT 141.410 143.650 156.785 143.780 ;
        RECT 141.410 143.640 146.570 143.650 ;
        RECT 141.410 143.550 145.410 143.640 ;
        RECT 148.785 143.560 156.785 143.650 ;
        RECT 148.870 143.550 156.760 143.560 ;
        RECT 141.020 143.190 141.250 143.500 ;
        RECT 141.470 143.190 145.370 143.550 ;
        RECT 145.570 143.190 145.800 143.500 ;
        RECT 141.020 141.850 145.800 143.190 ;
        RECT 141.020 141.540 141.250 141.850 ;
        RECT 145.570 141.540 145.800 141.850 ;
        RECT 148.350 142.970 148.580 143.510 ;
        RECT 149.390 142.970 150.400 143.000 ;
        RECT 156.990 142.970 157.220 143.510 ;
        RECT 148.350 142.070 157.220 142.970 ;
        RECT 148.350 141.550 148.580 142.070 ;
        RECT 149.390 142.000 150.400 142.070 ;
        RECT 156.990 141.550 157.220 142.070 ;
        RECT 141.410 141.260 145.410 141.490 ;
        RECT 148.785 141.270 156.785 141.500 ;
        RECT 139.930 141.110 141.090 141.150 ;
        RECT 139.930 141.030 141.330 141.110 ;
        RECT 141.700 141.040 145.360 141.260 ;
        RECT 141.700 141.030 143.140 141.040 ;
        RECT 139.930 140.990 143.140 141.030 ;
        RECT 139.930 140.900 142.650 140.990 ;
        RECT 148.850 140.980 156.740 141.270 ;
        RECT 139.930 140.840 141.980 140.900 ;
        RECT 139.930 140.790 141.730 140.840 ;
        RECT 139.930 137.450 140.790 140.790 ;
        RECT 148.840 140.490 156.760 140.500 ;
        RECT 145.070 140.480 156.760 140.490 ;
        RECT 141.450 140.360 156.760 140.480 ;
        RECT 141.450 140.350 156.785 140.360 ;
        RECT 141.410 140.230 156.785 140.350 ;
        RECT 141.410 140.120 145.410 140.230 ;
        RECT 141.020 139.780 141.250 140.070 ;
        RECT 141.470 139.780 145.360 140.120 ;
        RECT 145.570 139.780 145.800 140.070 ;
        RECT 141.020 138.410 145.800 139.780 ;
        RECT 141.020 138.110 141.250 138.410 ;
        RECT 145.570 138.110 145.800 138.410 ;
        RECT 141.410 137.830 145.410 138.060 ;
        RECT 141.660 137.600 145.230 137.830 ;
        RECT 141.660 137.450 145.350 137.600 ;
        RECT 139.930 137.170 145.350 137.450 ;
        RECT 146.600 137.280 147.220 140.230 ;
        RECT 148.785 140.130 156.785 140.230 ;
        RECT 148.840 140.120 156.760 140.130 ;
        RECT 148.350 139.420 148.580 140.080 ;
        RECT 149.360 139.420 150.360 139.510 ;
        RECT 156.990 139.420 157.220 140.080 ;
        RECT 148.350 138.600 157.220 139.420 ;
        RECT 148.350 138.120 148.580 138.600 ;
        RECT 149.360 138.510 150.360 138.600 ;
        RECT 156.990 138.120 157.220 138.600 ;
        RECT 148.785 137.840 156.785 138.070 ;
        RECT 139.930 136.710 145.360 137.170 ;
        RECT 139.930 135.360 141.960 136.710 ;
        RECT 143.710 136.700 145.360 136.710 ;
        RECT 142.400 135.430 143.400 136.150 ;
        RECT 143.710 135.890 144.020 136.700 ;
        RECT 144.480 136.420 145.360 136.700 ;
        RECT 145.600 136.880 147.220 137.280 ;
        RECT 148.870 136.930 156.740 137.840 ;
        RECT 144.420 136.190 145.420 136.420 ;
        RECT 145.600 136.230 145.950 136.880 ;
        RECT 146.600 136.870 147.220 136.880 ;
        RECT 148.785 136.700 156.785 136.930 ;
        RECT 148.870 136.690 156.740 136.700 ;
        RECT 144.480 135.980 145.360 136.000 ;
        RECT 143.750 135.600 144.020 135.890 ;
        RECT 144.420 135.750 145.420 135.980 ;
        RECT 145.580 135.940 145.950 136.230 ;
        RECT 145.610 135.880 145.950 135.940 ;
        RECT 146.710 136.550 147.470 136.600 ;
        RECT 148.350 136.550 148.580 136.650 ;
        RECT 146.710 136.340 148.580 136.550 ;
        RECT 156.990 136.340 157.220 136.650 ;
        RECT 146.710 135.920 149.250 136.340 ;
        RECT 156.620 135.920 157.220 136.340 ;
        RECT 144.480 135.600 145.360 135.750 ;
        RECT 144.490 135.430 145.220 135.600 ;
        RECT 126.020 133.880 138.460 133.900 ;
        RECT 125.490 133.720 125.830 133.830 ;
        RECT 126.060 133.870 131.730 133.880 ;
        RECT 132.730 133.870 138.460 133.880 ;
        RECT 122.370 133.470 125.230 133.640 ;
        RECT 126.060 133.470 126.490 133.870 ;
        RECT 122.340 133.100 126.490 133.470 ;
        RECT 104.490 131.320 109.730 131.330 ;
        RECT 101.540 131.220 116.840 131.320 ;
        RECT 101.540 131.210 116.875 131.220 ;
        RECT 101.500 131.090 116.875 131.210 ;
        RECT 101.500 130.980 105.500 131.090 ;
        RECT 106.550 131.010 108.290 131.090 ;
        RECT 108.870 131.010 116.875 131.090 ;
        RECT 106.550 130.930 107.800 131.010 ;
        RECT 108.875 130.990 116.875 131.010 ;
        RECT 101.110 130.680 101.340 130.930 ;
        RECT 105.660 130.790 105.890 130.930 ;
        RECT 108.440 130.790 108.670 130.940 ;
        RECT 105.660 130.680 108.670 130.790 ;
        RECT 117.080 130.680 117.310 130.940 ;
        RECT 101.110 130.240 117.310 130.680 ;
        RECT 101.110 129.970 101.340 130.240 ;
        RECT 105.660 130.210 117.310 130.240 ;
        RECT 105.660 130.120 108.670 130.210 ;
        RECT 105.660 129.970 105.890 130.120 ;
        RECT 108.440 129.980 108.670 130.120 ;
        RECT 117.080 129.980 117.310 130.210 ;
        RECT 101.500 129.690 105.500 129.920 ;
        RECT 108.875 129.710 116.875 129.930 ;
        RECT 117.640 129.710 118.600 131.750 ;
        RECT 108.875 129.700 118.600 129.710 ;
        RECT 101.500 129.620 105.490 129.690 ;
        RECT 74.730 129.560 75.050 129.620 ;
        RECT 76.570 129.560 76.890 129.620 ;
        RECT 74.730 129.420 76.890 129.560 ;
        RECT 74.730 129.360 75.050 129.420 ;
        RECT 76.570 129.360 76.890 129.420 ;
        RECT 79.330 129.360 79.650 129.620 ;
        RECT 82.090 129.560 82.410 129.620 ;
        RECT 82.090 129.420 85.540 129.560 ;
        RECT 82.090 129.360 82.410 129.420 ;
        RECT 62.860 129.080 64.010 129.220 ;
        RECT 48.970 128.740 49.485 128.880 ;
        RECT 50.365 128.740 52.970 128.880 ;
        RECT 48.970 128.695 49.320 128.740 ;
        RECT 50.365 128.695 50.655 128.740 ;
        RECT 48.970 128.680 49.290 128.695 ;
        RECT 52.650 128.680 52.970 128.740 ;
        RECT 55.425 128.695 55.715 128.925 ;
        RECT 55.870 128.680 56.190 128.940 ;
        RECT 62.860 128.925 63.000 129.080 ;
        RECT 63.690 129.020 64.010 129.080 ;
        RECT 64.240 129.080 67.690 129.220 ;
        RECT 56.805 128.880 57.095 128.925 ;
        RECT 62.785 128.880 63.075 128.925 ;
        RECT 56.805 128.740 63.075 128.880 ;
        RECT 56.805 128.695 57.095 128.740 ;
        RECT 62.785 128.695 63.075 128.740 ;
        RECT 63.230 128.680 63.550 128.940 ;
        RECT 64.240 128.925 64.380 129.080 ;
        RECT 67.370 129.020 67.690 129.080 ;
        RECT 68.775 129.220 69.065 129.265 ;
        RECT 71.295 129.220 71.585 129.265 ;
        RECT 72.485 129.220 72.775 129.265 ;
        RECT 68.775 129.080 72.775 129.220 ;
        RECT 68.775 129.035 69.065 129.080 ;
        RECT 71.295 129.035 71.585 129.080 ;
        RECT 72.485 129.035 72.775 129.080 ;
        RECT 73.365 129.035 73.655 129.265 ;
        RECT 75.650 129.220 75.970 129.280 ;
        RECT 75.280 129.080 75.970 129.220 ;
        RECT 64.165 128.695 64.455 128.925 ;
        RECT 64.625 128.880 64.915 128.925 ;
        RECT 65.070 128.880 65.390 128.940 ;
        RECT 64.625 128.740 65.390 128.880 ;
        RECT 64.625 128.695 64.915 128.740 ;
        RECT 65.070 128.680 65.390 128.740 ;
        RECT 65.545 128.880 65.835 128.925 ;
        RECT 67.830 128.880 68.150 128.940 ;
        RECT 65.545 128.740 68.150 128.880 ;
        RECT 65.545 128.695 65.835 128.740 ;
        RECT 67.830 128.680 68.150 128.740 ;
        RECT 74.285 128.880 74.575 128.925 ;
        RECT 74.730 128.880 75.050 128.940 ;
        RECT 75.280 128.925 75.420 129.080 ;
        RECT 75.650 129.020 75.970 129.080 ;
        RECT 76.110 129.220 76.430 129.280 ;
        RECT 79.420 129.220 79.560 129.360 ;
        RECT 76.110 129.080 82.780 129.220 ;
        RECT 76.110 129.020 76.430 129.080 ;
        RECT 78.500 128.925 78.640 129.080 ;
        RECT 74.285 128.740 75.050 128.880 ;
        RECT 74.285 128.695 74.575 128.740 ;
        RECT 74.730 128.680 75.050 128.740 ;
        RECT 75.205 128.695 75.495 128.925 ;
        RECT 78.425 128.695 78.715 128.925 ;
        RECT 78.870 128.680 79.190 128.940 ;
        RECT 79.345 128.680 79.635 128.910 ;
        RECT 80.265 128.880 80.555 128.925 ;
        RECT 80.725 128.880 81.015 128.925 ;
        RECT 81.170 128.880 81.490 128.940 ;
        RECT 80.265 128.740 81.490 128.880 ;
        RECT 80.265 128.695 80.555 128.740 ;
        RECT 80.725 128.695 81.015 128.740 ;
        RECT 81.170 128.680 81.490 128.740 ;
        RECT 81.630 128.680 81.950 128.940 ;
        RECT 82.640 128.925 82.780 129.080 ;
        RECT 82.105 128.695 82.395 128.925 ;
        RECT 82.565 128.695 82.855 128.925 ;
        RECT 84.390 128.880 84.710 128.940 ;
        RECT 85.400 128.925 85.540 129.420 ;
        RECT 100.010 129.510 105.490 129.620 ;
        RECT 108.930 129.540 118.600 129.700 ;
        RECT 100.010 129.420 103.180 129.510 ;
        RECT 116.670 129.490 118.600 129.540 ;
        RECT 85.325 128.880 85.615 128.925 ;
        RECT 84.390 128.740 85.615 128.880 ;
        RECT 31.045 128.400 34.020 128.540 ;
        RECT 34.250 128.540 34.570 128.600 ;
        RECT 35.770 128.540 36.060 128.585 ;
        RECT 34.250 128.400 36.060 128.540 ;
        RECT 31.045 128.355 31.335 128.400 ;
        RECT 32.410 128.340 32.730 128.400 ;
        RECT 34.250 128.340 34.570 128.400 ;
        RECT 35.770 128.355 36.060 128.400 ;
        RECT 37.010 128.340 37.330 128.600 ;
        RECT 56.345 128.540 56.635 128.585 ;
        RECT 69.210 128.540 69.530 128.600 ;
        RECT 56.345 128.400 69.530 128.540 ;
        RECT 56.345 128.355 56.635 128.400 ;
        RECT 69.210 128.340 69.530 128.400 ;
        RECT 71.510 128.540 71.830 128.600 ;
        RECT 72.030 128.540 72.320 128.585 ;
        RECT 71.510 128.400 72.320 128.540 ;
        RECT 71.510 128.340 71.830 128.400 ;
        RECT 72.030 128.355 72.320 128.400 ;
        RECT 76.125 128.540 76.415 128.585 ;
        RECT 79.420 128.540 79.560 128.680 ;
        RECT 76.125 128.400 79.560 128.540 ;
        RECT 82.180 128.540 82.320 128.695 ;
        RECT 84.390 128.680 84.710 128.740 ;
        RECT 85.325 128.695 85.615 128.740 ;
        RECT 87.165 128.880 87.455 128.925 ;
        RECT 87.610 128.880 87.930 128.940 ;
        RECT 87.165 128.740 87.930 128.880 ;
        RECT 87.165 128.695 87.455 128.740 ;
        RECT 87.610 128.680 87.930 128.740 ;
        RECT 83.470 128.540 83.790 128.600 ;
        RECT 82.180 128.400 83.790 128.540 ;
        RECT 76.125 128.355 76.415 128.400 ;
        RECT 83.470 128.340 83.790 128.400 ;
        RECT 85.770 128.340 86.090 128.600 ;
        RECT 86.230 128.540 86.550 128.600 ;
        RECT 88.530 128.540 88.850 128.600 ;
        RECT 86.230 128.400 88.850 128.540 ;
        RECT 86.230 128.340 86.550 128.400 ;
        RECT 88.530 128.340 88.850 128.400 ;
        RECT 22.290 128.060 26.660 128.200 ;
        RECT 26.890 128.200 27.210 128.260 ;
        RECT 27.825 128.200 28.115 128.245 ;
        RECT 26.890 128.060 28.115 128.200 ;
        RECT 22.290 128.000 22.610 128.060 ;
        RECT 26.890 128.000 27.210 128.060 ;
        RECT 27.825 128.015 28.115 128.060 ;
        RECT 32.885 128.200 33.175 128.245 ;
        RECT 33.330 128.200 33.650 128.260 ;
        RECT 32.885 128.060 33.650 128.200 ;
        RECT 32.885 128.015 33.175 128.060 ;
        RECT 33.330 128.000 33.650 128.060 ;
        RECT 33.790 128.200 34.110 128.260 ;
        RECT 35.185 128.200 35.475 128.245 ;
        RECT 33.790 128.060 35.475 128.200 ;
        RECT 33.790 128.000 34.110 128.060 ;
        RECT 35.185 128.015 35.475 128.060 ;
        RECT 36.565 128.200 36.855 128.245 ;
        RECT 37.470 128.200 37.790 128.260 ;
        RECT 36.565 128.060 37.790 128.200 ;
        RECT 36.565 128.015 36.855 128.060 ;
        RECT 37.470 128.000 37.790 128.060 ;
        RECT 37.930 128.000 38.250 128.260 ;
        RECT 54.950 128.000 55.270 128.260 ;
        RECT 59.105 128.200 59.395 128.245 ;
        RECT 61.390 128.200 61.710 128.260 ;
        RECT 59.105 128.060 61.710 128.200 ;
        RECT 59.105 128.015 59.395 128.060 ;
        RECT 61.390 128.000 61.710 128.060 ;
        RECT 61.865 128.200 62.155 128.245 ;
        RECT 62.310 128.200 62.630 128.260 ;
        RECT 63.230 128.200 63.550 128.260 ;
        RECT 61.865 128.060 63.550 128.200 ;
        RECT 61.865 128.015 62.155 128.060 ;
        RECT 62.310 128.000 62.630 128.060 ;
        RECT 63.230 128.000 63.550 128.060 ;
        RECT 63.690 128.000 64.010 128.260 ;
        RECT 65.070 128.000 65.390 128.260 ;
        RECT 77.030 128.000 77.350 128.260 ;
        RECT 77.490 128.200 77.810 128.260 ;
        RECT 85.860 128.200 86.000 128.340 ;
        RECT 77.490 128.060 86.000 128.200 ;
        RECT 77.490 128.000 77.810 128.060 ;
        RECT 12.100 127.380 89.840 127.860 ;
        RECT 21.370 126.980 21.690 127.240 ;
        RECT 59.550 126.980 59.870 127.240 ;
        RECT 70.590 127.180 70.910 127.240 ;
        RECT 71.510 127.180 71.830 127.240 ;
        RECT 64.240 127.040 67.600 127.180 ;
        RECT 64.240 126.900 64.380 127.040 ;
        RECT 34.710 126.840 35.030 126.900 ;
        RECT 13.640 126.700 35.030 126.840 ;
        RECT 13.640 126.560 13.780 126.700 ;
        RECT 13.550 126.300 13.870 126.560 ;
        RECT 14.930 126.545 15.250 126.560 ;
        RECT 14.900 126.315 15.250 126.545 ;
        RECT 14.930 126.300 15.250 126.315 ;
        RECT 20.910 126.300 21.230 126.560 ;
        RECT 21.830 126.300 22.150 126.560 ;
        RECT 22.290 126.300 22.610 126.560 ;
        RECT 23.210 126.300 23.530 126.560 ;
        RECT 23.670 126.300 23.990 126.560 ;
        RECT 24.145 126.315 24.435 126.545 ;
        RECT 25.050 126.500 25.370 126.560 ;
        RECT 27.365 126.500 27.655 126.545 ;
        RECT 25.050 126.360 27.655 126.500 ;
        RECT 14.445 126.160 14.735 126.205 ;
        RECT 15.635 126.160 15.925 126.205 ;
        RECT 18.155 126.160 18.445 126.205 ;
        RECT 14.445 126.020 18.445 126.160 ;
        RECT 21.920 126.160 22.060 126.300 ;
        RECT 24.220 126.160 24.360 126.315 ;
        RECT 25.050 126.300 25.370 126.360 ;
        RECT 27.365 126.315 27.655 126.360 ;
        RECT 27.810 126.300 28.130 126.560 ;
        RECT 30.660 126.545 30.800 126.700 ;
        RECT 34.710 126.640 35.030 126.700 ;
        RECT 52.650 126.840 52.970 126.900 ;
        RECT 64.150 126.840 64.470 126.900 ;
        RECT 52.650 126.700 64.470 126.840 ;
        RECT 52.650 126.640 52.970 126.700 ;
        RECT 64.150 126.640 64.470 126.700 ;
        RECT 65.545 126.840 65.835 126.885 ;
        RECT 66.450 126.840 66.770 126.900 ;
        RECT 65.545 126.700 66.770 126.840 ;
        RECT 65.545 126.655 65.835 126.700 ;
        RECT 66.450 126.640 66.770 126.700 ;
        RECT 29.205 126.315 29.495 126.545 ;
        RECT 30.585 126.315 30.875 126.545 ;
        RECT 31.920 126.500 32.210 126.545 ;
        RECT 33.330 126.500 33.650 126.560 ;
        RECT 31.920 126.360 33.650 126.500 ;
        RECT 31.920 126.315 32.210 126.360 ;
        RECT 21.920 126.020 24.360 126.160 ;
        RECT 24.590 126.160 24.910 126.220 ;
        RECT 26.890 126.160 27.210 126.220 ;
        RECT 29.280 126.160 29.420 126.315 ;
        RECT 33.330 126.300 33.650 126.360 ;
        RECT 54.000 126.500 54.290 126.545 ;
        RECT 59.090 126.500 59.410 126.560 ;
        RECT 54.000 126.360 59.410 126.500 ;
        RECT 54.000 126.315 54.290 126.360 ;
        RECT 59.090 126.300 59.410 126.360 ;
        RECT 59.550 126.500 59.870 126.560 ;
        RECT 60.025 126.500 60.315 126.545 ;
        RECT 59.550 126.360 60.315 126.500 ;
        RECT 59.550 126.300 59.870 126.360 ;
        RECT 60.025 126.315 60.315 126.360 ;
        RECT 63.690 126.500 64.010 126.560 ;
        RECT 65.085 126.500 65.375 126.545 ;
        RECT 63.690 126.360 65.375 126.500 ;
        RECT 63.690 126.300 64.010 126.360 ;
        RECT 65.085 126.315 65.375 126.360 ;
        RECT 24.590 126.020 29.420 126.160 ;
        RECT 31.465 126.160 31.755 126.205 ;
        RECT 32.655 126.160 32.945 126.205 ;
        RECT 35.175 126.160 35.465 126.205 ;
        RECT 31.465 126.020 35.465 126.160 ;
        RECT 14.445 125.975 14.735 126.020 ;
        RECT 15.635 125.975 15.925 126.020 ;
        RECT 18.155 125.975 18.445 126.020 ;
        RECT 24.590 125.960 24.910 126.020 ;
        RECT 26.890 125.960 27.210 126.020 ;
        RECT 31.465 125.975 31.755 126.020 ;
        RECT 32.655 125.975 32.945 126.020 ;
        RECT 35.175 125.975 35.465 126.020 ;
        RECT 52.650 125.960 52.970 126.220 ;
        RECT 53.545 126.160 53.835 126.205 ;
        RECT 54.735 126.160 55.025 126.205 ;
        RECT 57.255 126.160 57.545 126.205 ;
        RECT 53.545 126.020 57.545 126.160 ;
        RECT 53.545 125.975 53.835 126.020 ;
        RECT 54.735 125.975 55.025 126.020 ;
        RECT 57.255 125.975 57.545 126.020 ;
        RECT 61.390 126.160 61.710 126.220 ;
        RECT 63.245 126.160 63.535 126.205 ;
        RECT 61.390 126.020 63.535 126.160 ;
        RECT 61.390 125.960 61.710 126.020 ;
        RECT 63.245 125.975 63.535 126.020 ;
        RECT 14.050 125.820 14.340 125.865 ;
        RECT 16.150 125.820 16.440 125.865 ;
        RECT 17.720 125.820 18.010 125.865 ;
        RECT 14.050 125.680 18.010 125.820 ;
        RECT 14.050 125.635 14.340 125.680 ;
        RECT 16.150 125.635 16.440 125.680 ;
        RECT 17.720 125.635 18.010 125.680 ;
        RECT 28.745 125.820 29.035 125.865 ;
        RECT 30.570 125.820 30.890 125.880 ;
        RECT 28.745 125.680 30.890 125.820 ;
        RECT 28.745 125.635 29.035 125.680 ;
        RECT 30.570 125.620 30.890 125.680 ;
        RECT 31.070 125.820 31.360 125.865 ;
        RECT 33.170 125.820 33.460 125.865 ;
        RECT 34.740 125.820 35.030 125.865 ;
        RECT 31.070 125.680 35.030 125.820 ;
        RECT 31.070 125.635 31.360 125.680 ;
        RECT 33.170 125.635 33.460 125.680 ;
        RECT 34.740 125.635 35.030 125.680 ;
        RECT 53.150 125.820 53.440 125.865 ;
        RECT 55.250 125.820 55.540 125.865 ;
        RECT 56.820 125.820 57.110 125.865 ;
        RECT 53.150 125.680 57.110 125.820 ;
        RECT 53.150 125.635 53.440 125.680 ;
        RECT 55.250 125.635 55.540 125.680 ;
        RECT 56.820 125.635 57.110 125.680 ;
        RECT 62.770 125.820 63.090 125.880 ;
        RECT 62.770 125.680 63.460 125.820 ;
        RECT 62.770 125.620 63.090 125.680 ;
        RECT 20.465 125.480 20.755 125.525 ;
        RECT 21.370 125.480 21.690 125.540 ;
        RECT 20.465 125.340 21.690 125.480 ;
        RECT 20.465 125.295 20.755 125.340 ;
        RECT 21.370 125.280 21.690 125.340 ;
        RECT 25.510 125.280 25.830 125.540 ;
        RECT 26.445 125.480 26.735 125.525 ;
        RECT 26.890 125.480 27.210 125.540 ;
        RECT 26.445 125.340 27.210 125.480 ;
        RECT 26.445 125.295 26.735 125.340 ;
        RECT 26.890 125.280 27.210 125.340 ;
        RECT 36.090 125.480 36.410 125.540 ;
        RECT 37.485 125.480 37.775 125.525 ;
        RECT 37.930 125.480 38.250 125.540 ;
        RECT 36.090 125.340 38.250 125.480 ;
        RECT 36.090 125.280 36.410 125.340 ;
        RECT 37.485 125.295 37.775 125.340 ;
        RECT 37.930 125.280 38.250 125.340 ;
        RECT 55.870 125.480 56.190 125.540 ;
        RECT 61.850 125.480 62.170 125.540 ;
        RECT 55.870 125.340 62.170 125.480 ;
        RECT 63.320 125.480 63.460 125.680 ;
        RECT 64.165 125.635 64.455 125.865 ;
        RECT 65.160 125.820 65.300 126.315 ;
        RECT 65.990 126.300 66.310 126.560 ;
        RECT 66.910 126.300 67.230 126.560 ;
        RECT 67.460 126.160 67.600 127.040 ;
        RECT 70.590 127.040 71.830 127.180 ;
        RECT 70.590 126.980 70.910 127.040 ;
        RECT 71.510 126.980 71.830 127.040 ;
        RECT 71.970 126.980 72.290 127.240 ;
        RECT 75.650 127.180 75.970 127.240 ;
        RECT 79.345 127.180 79.635 127.225 ;
        RECT 73.440 127.040 79.635 127.180 ;
        RECT 73.440 126.840 73.580 127.040 ;
        RECT 75.650 126.980 75.970 127.040 ;
        RECT 79.345 126.995 79.635 127.040 ;
        RECT 81.630 126.980 81.950 127.240 ;
        RECT 83.100 127.040 87.380 127.180 ;
        RECT 68.840 126.700 73.580 126.840 ;
        RECT 73.780 126.840 74.070 126.885 ;
        RECT 77.030 126.840 77.350 126.900 ;
        RECT 73.780 126.700 77.350 126.840 ;
        RECT 68.840 126.545 68.980 126.700 ;
        RECT 73.780 126.655 74.070 126.700 ;
        RECT 77.030 126.640 77.350 126.700 ;
        RECT 77.490 126.840 77.810 126.900 ;
        RECT 80.725 126.840 81.015 126.885 ;
        RECT 83.100 126.840 83.240 127.040 ;
        RECT 87.240 126.885 87.380 127.040 ;
        RECT 86.245 126.840 86.535 126.885 ;
        RECT 77.490 126.700 81.015 126.840 ;
        RECT 77.490 126.640 77.810 126.700 ;
        RECT 80.725 126.655 81.015 126.700 ;
        RECT 81.720 126.700 83.240 126.840 ;
        RECT 83.560 126.700 86.535 126.840 ;
        RECT 68.765 126.315 69.055 126.545 ;
        RECT 69.210 126.300 69.530 126.560 ;
        RECT 70.130 126.300 70.450 126.560 ;
        RECT 70.590 126.300 70.910 126.560 ;
        RECT 71.065 126.500 71.355 126.545 ;
        RECT 71.970 126.500 72.290 126.560 ;
        RECT 71.065 126.360 72.290 126.500 ;
        RECT 71.065 126.315 71.355 126.360 ;
        RECT 71.970 126.300 72.290 126.360 ;
        RECT 79.805 126.500 80.095 126.545 ;
        RECT 81.720 126.500 81.860 126.700 ;
        RECT 83.560 126.560 83.700 126.700 ;
        RECT 86.245 126.655 86.535 126.700 ;
        RECT 87.165 126.840 87.455 126.885 ;
        RECT 88.990 126.840 89.310 126.900 ;
        RECT 87.165 126.700 89.310 126.840 ;
        RECT 87.165 126.655 87.455 126.700 ;
        RECT 88.990 126.640 89.310 126.700 ;
        RECT 79.805 126.360 81.860 126.500 ;
        RECT 79.805 126.315 80.095 126.360 ;
        RECT 82.090 126.300 82.410 126.560 ;
        RECT 83.025 126.315 83.315 126.545 ;
        RECT 72.430 126.160 72.750 126.220 ;
        RECT 67.460 126.020 72.750 126.160 ;
        RECT 72.430 125.960 72.750 126.020 ;
        RECT 73.325 126.160 73.615 126.205 ;
        RECT 74.515 126.160 74.805 126.205 ;
        RECT 77.035 126.160 77.325 126.205 ;
        RECT 82.550 126.160 82.870 126.220 ;
        RECT 73.325 126.020 77.325 126.160 ;
        RECT 73.325 125.975 73.615 126.020 ;
        RECT 74.515 125.975 74.805 126.020 ;
        RECT 77.035 125.975 77.325 126.020 ;
        RECT 77.580 126.020 82.870 126.160 ;
        RECT 83.100 126.160 83.240 126.315 ;
        RECT 83.470 126.300 83.790 126.560 ;
        RECT 83.945 126.500 84.235 126.545 ;
        RECT 84.390 126.500 84.710 126.560 ;
        RECT 83.945 126.360 87.380 126.500 ;
        RECT 83.945 126.315 84.235 126.360 ;
        RECT 84.390 126.300 84.710 126.360 ;
        RECT 87.240 126.220 87.380 126.360 ;
        RECT 84.850 126.160 85.170 126.220 ;
        RECT 86.230 126.160 86.550 126.220 ;
        RECT 83.100 126.020 86.550 126.160 ;
        RECT 66.910 125.820 67.230 125.880 ;
        RECT 65.160 125.680 67.230 125.820 ;
        RECT 64.240 125.480 64.380 125.635 ;
        RECT 66.910 125.620 67.230 125.680 ;
        RECT 72.930 125.820 73.220 125.865 ;
        RECT 75.030 125.820 75.320 125.865 ;
        RECT 76.600 125.820 76.890 125.865 ;
        RECT 72.930 125.680 76.890 125.820 ;
        RECT 72.930 125.635 73.220 125.680 ;
        RECT 75.030 125.635 75.320 125.680 ;
        RECT 76.600 125.635 76.890 125.680 ;
        RECT 63.320 125.340 64.380 125.480 ;
        RECT 67.845 125.480 68.135 125.525 ;
        RECT 77.580 125.480 77.720 126.020 ;
        RECT 82.550 125.960 82.870 126.020 ;
        RECT 84.850 125.960 85.170 126.020 ;
        RECT 86.230 125.960 86.550 126.020 ;
        RECT 87.150 125.960 87.470 126.220 ;
        RECT 100.010 126.150 100.880 129.420 ;
        RECT 104.530 128.960 109.780 128.970 ;
        RECT 104.530 128.850 116.840 128.960 ;
        RECT 101.560 128.790 116.840 128.850 ;
        RECT 101.560 128.780 116.875 128.790 ;
        RECT 101.500 128.650 116.875 128.780 ;
        RECT 101.500 128.640 106.660 128.650 ;
        RECT 101.500 128.550 105.500 128.640 ;
        RECT 108.875 128.560 116.875 128.650 ;
        RECT 108.960 128.550 116.850 128.560 ;
        RECT 101.110 128.190 101.340 128.500 ;
        RECT 101.560 128.190 105.460 128.550 ;
        RECT 105.660 128.190 105.890 128.500 ;
        RECT 101.110 126.850 105.890 128.190 ;
        RECT 101.110 126.540 101.340 126.850 ;
        RECT 105.660 126.540 105.890 126.850 ;
        RECT 108.440 127.970 108.670 128.510 ;
        RECT 109.480 127.970 110.490 128.000 ;
        RECT 117.080 127.970 117.310 128.510 ;
        RECT 108.440 127.070 117.310 127.970 ;
        RECT 108.440 126.550 108.670 127.070 ;
        RECT 109.480 127.000 110.490 127.070 ;
        RECT 117.080 126.550 117.310 127.070 ;
        RECT 101.500 126.260 105.500 126.490 ;
        RECT 108.875 126.270 116.875 126.500 ;
        RECT 100.010 126.110 101.180 126.150 ;
        RECT 100.010 126.030 101.420 126.110 ;
        RECT 101.790 126.040 105.450 126.260 ;
        RECT 101.790 126.030 103.230 126.040 ;
        RECT 100.010 125.990 103.230 126.030 ;
        RECT 100.010 125.900 102.740 125.990 ;
        RECT 108.940 125.980 116.830 126.270 ;
        RECT 77.950 125.820 78.270 125.880 ;
        RECT 85.325 125.820 85.615 125.865 ;
        RECT 77.950 125.680 85.615 125.820 ;
        RECT 77.950 125.620 78.270 125.680 ;
        RECT 85.325 125.635 85.615 125.680 ;
        RECT 100.010 125.840 102.070 125.900 ;
        RECT 100.010 125.790 101.820 125.840 ;
        RECT 67.845 125.340 77.720 125.480 ;
        RECT 83.010 125.480 83.330 125.540 ;
        RECT 84.865 125.480 85.155 125.525 ;
        RECT 83.010 125.340 85.155 125.480 ;
        RECT 55.870 125.280 56.190 125.340 ;
        RECT 61.850 125.280 62.170 125.340 ;
        RECT 67.845 125.295 68.135 125.340 ;
        RECT 83.010 125.280 83.330 125.340 ;
        RECT 84.865 125.295 85.155 125.340 ;
        RECT 12.100 124.660 89.840 125.140 ;
        RECT 14.485 124.460 14.775 124.505 ;
        RECT 14.930 124.460 15.250 124.520 ;
        RECT 14.485 124.320 15.250 124.460 ;
        RECT 14.485 124.275 14.775 124.320 ;
        RECT 14.930 124.260 15.250 124.320 ;
        RECT 19.530 124.260 19.850 124.520 ;
        RECT 21.370 124.460 21.690 124.520 ;
        RECT 22.765 124.460 23.055 124.505 ;
        RECT 21.370 124.320 23.055 124.460 ;
        RECT 21.370 124.260 21.690 124.320 ;
        RECT 22.765 124.275 23.055 124.320 ;
        RECT 46.670 124.260 46.990 124.520 ;
        RECT 49.890 124.460 50.210 124.520 ;
        RECT 52.205 124.460 52.495 124.505 ;
        RECT 57.710 124.460 58.030 124.520 ;
        RECT 49.890 124.320 52.495 124.460 ;
        RECT 49.890 124.260 50.210 124.320 ;
        RECT 52.205 124.275 52.495 124.320 ;
        RECT 55.040 124.320 58.030 124.460 ;
        RECT 19.990 124.120 20.310 124.180 ;
        RECT 16.400 123.980 20.310 124.120 ;
        RECT 16.400 123.825 16.540 123.980 ;
        RECT 19.990 123.920 20.310 123.980 ;
        RECT 21.830 124.120 22.150 124.180 ;
        RECT 22.305 124.120 22.595 124.165 ;
        RECT 34.710 124.120 35.000 124.165 ;
        RECT 36.280 124.120 36.570 124.165 ;
        RECT 38.380 124.120 38.670 124.165 ;
        RECT 21.830 123.980 23.440 124.120 ;
        RECT 21.830 123.920 22.150 123.980 ;
        RECT 22.305 123.935 22.595 123.980 ;
        RECT 23.300 123.840 23.440 123.980 ;
        RECT 34.710 123.980 38.670 124.120 ;
        RECT 34.710 123.935 35.000 123.980 ;
        RECT 36.280 123.935 36.570 123.980 ;
        RECT 38.380 123.935 38.670 123.980 ;
        RECT 42.070 124.120 42.360 124.165 ;
        RECT 43.640 124.120 43.930 124.165 ;
        RECT 45.740 124.120 46.030 124.165 ;
        RECT 42.070 123.980 46.030 124.120 ;
        RECT 42.070 123.935 42.360 123.980 ;
        RECT 43.640 123.935 43.930 123.980 ;
        RECT 45.740 123.935 46.030 123.980 ;
        RECT 16.325 123.595 16.615 123.825 ;
        RECT 16.770 123.780 17.090 123.840 ;
        RECT 17.705 123.780 17.995 123.825 ;
        RECT 16.770 123.640 17.995 123.780 ;
        RECT 16.770 123.580 17.090 123.640 ;
        RECT 17.705 123.595 17.995 123.640 ;
        RECT 23.210 123.580 23.530 123.840 ;
        RECT 34.275 123.780 34.565 123.825 ;
        RECT 36.795 123.780 37.085 123.825 ;
        RECT 37.985 123.780 38.275 123.825 ;
        RECT 34.275 123.640 38.275 123.780 ;
        RECT 34.275 123.595 34.565 123.640 ;
        RECT 36.795 123.595 37.085 123.640 ;
        RECT 37.985 123.595 38.275 123.640 ;
        RECT 41.635 123.780 41.925 123.825 ;
        RECT 44.155 123.780 44.445 123.825 ;
        RECT 45.345 123.780 45.635 123.825 ;
        RECT 41.635 123.640 45.635 123.780 ;
        RECT 41.635 123.595 41.925 123.640 ;
        RECT 44.155 123.595 44.445 123.640 ;
        RECT 45.345 123.595 45.635 123.640 ;
        RECT 46.225 123.780 46.515 123.825 ;
        RECT 48.050 123.780 48.370 123.840 ;
        RECT 46.225 123.640 48.370 123.780 ;
        RECT 46.225 123.595 46.515 123.640 ;
        RECT 48.050 123.580 48.370 123.640 ;
        RECT 54.030 123.780 54.350 123.840 ;
        RECT 55.040 123.825 55.180 124.320 ;
        RECT 57.710 124.260 58.030 124.320 ;
        RECT 59.090 124.460 59.410 124.520 ;
        RECT 60.025 124.460 60.315 124.505 ;
        RECT 59.090 124.320 60.315 124.460 ;
        RECT 59.090 124.260 59.410 124.320 ;
        RECT 60.025 124.275 60.315 124.320 ;
        RECT 61.850 124.460 62.170 124.520 ;
        RECT 62.325 124.460 62.615 124.505 ;
        RECT 61.850 124.320 62.615 124.460 ;
        RECT 61.850 124.260 62.170 124.320 ;
        RECT 62.325 124.275 62.615 124.320 ;
        RECT 62.770 124.460 63.090 124.520 ;
        RECT 63.705 124.460 63.995 124.505 ;
        RECT 62.770 124.320 63.995 124.460 ;
        RECT 62.770 124.260 63.090 124.320 ;
        RECT 63.705 124.275 63.995 124.320 ;
        RECT 64.165 124.460 64.455 124.505 ;
        RECT 64.610 124.460 64.930 124.520 ;
        RECT 64.165 124.320 64.930 124.460 ;
        RECT 64.165 124.275 64.455 124.320 ;
        RECT 64.610 124.260 64.930 124.320 ;
        RECT 65.545 124.460 65.835 124.505 ;
        RECT 65.990 124.460 66.310 124.520 ;
        RECT 65.545 124.320 66.310 124.460 ;
        RECT 65.545 124.275 65.835 124.320 ;
        RECT 65.990 124.260 66.310 124.320 ;
        RECT 66.910 124.260 67.230 124.520 ;
        RECT 73.810 124.460 74.130 124.520 ;
        RECT 74.730 124.460 75.050 124.520 ;
        RECT 83.930 124.460 84.250 124.520 ;
        RECT 73.810 124.320 75.050 124.460 ;
        RECT 73.810 124.260 74.130 124.320 ;
        RECT 74.730 124.260 75.050 124.320 ;
        RECT 78.500 124.320 84.250 124.460 ;
        RECT 67.000 124.120 67.140 124.260 ;
        RECT 76.110 124.120 76.430 124.180 ;
        RECT 66.080 123.980 67.140 124.120 ;
        RECT 68.380 123.980 76.430 124.120 ;
        RECT 54.965 123.780 55.255 123.825 ;
        RECT 54.030 123.640 55.255 123.780 ;
        RECT 54.030 123.580 54.350 123.640 ;
        RECT 54.965 123.595 55.255 123.640 ;
        RECT 57.250 123.780 57.570 123.840 ;
        RECT 57.250 123.640 62.080 123.780 ;
        RECT 57.250 123.580 57.570 123.640 ;
        RECT 15.865 123.440 16.155 123.485 ;
        RECT 17.230 123.440 17.550 123.500 ;
        RECT 15.865 123.300 17.550 123.440 ;
        RECT 15.865 123.255 16.155 123.300 ;
        RECT 17.230 123.240 17.550 123.300 ;
        RECT 18.150 123.240 18.470 123.500 ;
        RECT 19.085 123.440 19.375 123.485 ;
        RECT 20.910 123.440 21.230 123.500 ;
        RECT 19.085 123.300 21.230 123.440 ;
        RECT 19.085 123.255 19.375 123.300 ;
        RECT 20.910 123.240 21.230 123.300 ;
        RECT 21.370 123.240 21.690 123.500 ;
        RECT 22.750 123.240 23.070 123.500 ;
        RECT 25.510 123.240 25.830 123.500 ;
        RECT 26.445 123.255 26.735 123.485 ;
        RECT 26.905 123.255 27.195 123.485 ;
        RECT 27.350 123.440 27.670 123.500 ;
        RECT 37.470 123.485 37.790 123.500 ;
        RECT 30.125 123.440 30.415 123.485 ;
        RECT 27.350 123.300 30.415 123.440 ;
        RECT 15.280 123.100 15.570 123.145 ;
        RECT 18.625 123.100 18.915 123.145 ;
        RECT 21.830 123.100 22.150 123.160 ;
        RECT 26.520 123.100 26.660 123.255 ;
        RECT 15.280 122.960 18.915 123.100 ;
        RECT 15.280 122.915 15.570 122.960 ;
        RECT 18.625 122.915 18.915 122.960 ;
        RECT 21.000 122.960 22.150 123.100 ;
        RECT 19.070 122.760 19.390 122.820 ;
        RECT 21.000 122.805 21.140 122.960 ;
        RECT 21.830 122.900 22.150 122.960 ;
        RECT 24.680 122.960 26.660 123.100 ;
        RECT 26.980 123.100 27.120 123.255 ;
        RECT 27.350 123.240 27.670 123.300 ;
        RECT 30.125 123.255 30.415 123.300 ;
        RECT 37.470 123.440 37.820 123.485 ;
        RECT 38.390 123.440 38.710 123.500 ;
        RECT 38.865 123.440 39.155 123.485 ;
        RECT 37.470 123.300 37.985 123.440 ;
        RECT 38.390 123.300 39.155 123.440 ;
        RECT 37.470 123.255 37.820 123.300 ;
        RECT 37.470 123.240 37.790 123.255 ;
        RECT 38.390 123.240 38.710 123.300 ;
        RECT 38.865 123.255 39.155 123.300 ;
        RECT 46.685 123.255 46.975 123.485 ;
        RECT 47.605 123.440 47.895 123.485 ;
        RECT 49.430 123.440 49.750 123.500 ;
        RECT 47.605 123.300 49.750 123.440 ;
        RECT 47.605 123.255 47.895 123.300 ;
        RECT 27.810 123.100 28.130 123.160 ;
        RECT 29.205 123.100 29.495 123.145 ;
        RECT 45.000 123.100 45.290 123.145 ;
        RECT 46.760 123.100 46.900 123.255 ;
        RECT 49.430 123.240 49.750 123.300 ;
        RECT 54.505 123.440 54.795 123.485 ;
        RECT 55.410 123.440 55.730 123.500 ;
        RECT 56.345 123.440 56.635 123.485 ;
        RECT 54.505 123.300 56.635 123.440 ;
        RECT 54.505 123.255 54.795 123.300 ;
        RECT 55.410 123.240 55.730 123.300 ;
        RECT 56.345 123.255 56.635 123.300 ;
        RECT 60.010 123.440 60.330 123.500 ;
        RECT 60.945 123.440 61.235 123.485 ;
        RECT 60.010 123.300 61.235 123.440 ;
        RECT 60.010 123.240 60.330 123.300 ;
        RECT 60.945 123.255 61.235 123.300 ;
        RECT 61.390 123.240 61.710 123.500 ;
        RECT 61.940 123.440 62.080 123.640 ;
        RECT 64.610 123.620 64.930 123.880 ;
        RECT 65.085 123.820 65.375 123.825 ;
        RECT 65.530 123.820 65.850 123.840 ;
        RECT 66.080 123.825 66.220 123.980 ;
        RECT 65.085 123.680 65.850 123.820 ;
        RECT 65.085 123.595 65.375 123.680 ;
        RECT 65.530 123.580 65.850 123.680 ;
        RECT 66.005 123.595 66.295 123.825 ;
        RECT 66.910 123.780 67.230 123.840 ;
        RECT 68.380 123.780 68.520 123.980 ;
        RECT 76.110 123.920 76.430 123.980 ;
        RECT 66.910 123.640 68.520 123.780 ;
        RECT 66.910 123.580 67.230 123.640 ;
        RECT 62.770 123.440 63.090 123.500 ;
        RECT 61.940 123.300 63.090 123.440 ;
        RECT 62.770 123.240 63.090 123.300 ;
        RECT 63.230 123.240 63.550 123.500 ;
        RECT 66.450 123.240 66.770 123.500 ;
        RECT 67.830 123.240 68.150 123.500 ;
        RECT 68.380 123.485 68.520 123.640 ;
        RECT 68.750 123.780 69.070 123.840 ;
        RECT 70.145 123.780 70.435 123.825 ;
        RECT 68.750 123.640 70.435 123.780 ;
        RECT 68.750 123.580 69.070 123.640 ;
        RECT 70.145 123.595 70.435 123.640 ;
        RECT 71.510 123.780 71.830 123.840 ;
        RECT 73.810 123.780 74.130 123.840 ;
        RECT 71.510 123.640 74.130 123.780 ;
        RECT 71.510 123.580 71.830 123.640 ;
        RECT 73.810 123.580 74.130 123.640 ;
        RECT 68.305 123.255 68.595 123.485 ;
        RECT 69.685 123.440 69.975 123.485 ;
        RECT 70.590 123.440 70.910 123.500 ;
        RECT 69.685 123.300 70.910 123.440 ;
        RECT 69.685 123.255 69.975 123.300 ;
        RECT 70.590 123.240 70.910 123.300 ;
        RECT 77.030 123.240 77.350 123.500 ;
        RECT 77.950 123.240 78.270 123.500 ;
        RECT 78.500 123.485 78.640 124.320 ;
        RECT 83.930 124.260 84.250 124.320 ;
        RECT 81.210 124.120 81.500 124.165 ;
        RECT 83.310 124.120 83.600 124.165 ;
        RECT 84.880 124.120 85.170 124.165 ;
        RECT 81.210 123.980 85.170 124.120 ;
        RECT 81.210 123.935 81.500 123.980 ;
        RECT 83.310 123.935 83.600 123.980 ;
        RECT 84.880 123.935 85.170 123.980 ;
        RECT 81.605 123.780 81.895 123.825 ;
        RECT 82.795 123.780 83.085 123.825 ;
        RECT 85.315 123.780 85.605 123.825 ;
        RECT 81.605 123.640 85.605 123.780 ;
        RECT 81.605 123.595 81.895 123.640 ;
        RECT 82.795 123.595 83.085 123.640 ;
        RECT 85.315 123.595 85.605 123.640 ;
        RECT 78.425 123.255 78.715 123.485 ;
        RECT 78.870 123.240 79.190 123.500 ;
        RECT 80.725 123.440 81.015 123.485 ;
        RECT 79.420 123.300 81.015 123.440 ;
        RECT 48.510 123.100 48.830 123.160 ;
        RECT 67.370 123.100 67.690 123.160 ;
        RECT 26.980 122.960 30.340 123.100 ;
        RECT 24.680 122.805 24.820 122.960 ;
        RECT 27.810 122.900 28.130 122.960 ;
        RECT 29.205 122.915 29.495 122.960 ;
        RECT 30.200 122.820 30.340 122.960 ;
        RECT 45.000 122.960 46.440 123.100 ;
        RECT 46.760 122.960 48.830 123.100 ;
        RECT 45.000 122.915 45.290 122.960 ;
        RECT 20.465 122.760 20.755 122.805 ;
        RECT 19.070 122.620 20.755 122.760 ;
        RECT 19.070 122.560 19.390 122.620 ;
        RECT 20.465 122.575 20.755 122.620 ;
        RECT 20.925 122.575 21.215 122.805 ;
        RECT 24.605 122.575 24.895 122.805 ;
        RECT 28.745 122.760 29.035 122.805 ;
        RECT 29.650 122.760 29.970 122.820 ;
        RECT 28.745 122.620 29.970 122.760 ;
        RECT 28.745 122.575 29.035 122.620 ;
        RECT 29.650 122.560 29.970 122.620 ;
        RECT 30.110 122.560 30.430 122.820 ;
        RECT 30.570 122.760 30.890 122.820 ;
        RECT 31.045 122.760 31.335 122.805 ;
        RECT 30.570 122.620 31.335 122.760 ;
        RECT 30.570 122.560 30.890 122.620 ;
        RECT 31.045 122.575 31.335 122.620 ;
        RECT 31.965 122.760 32.255 122.805 ;
        RECT 33.330 122.760 33.650 122.820 ;
        RECT 31.965 122.620 33.650 122.760 ;
        RECT 31.965 122.575 32.255 122.620 ;
        RECT 33.330 122.560 33.650 122.620 ;
        RECT 39.325 122.760 39.615 122.805 ;
        RECT 41.150 122.760 41.470 122.820 ;
        RECT 39.325 122.620 41.470 122.760 ;
        RECT 46.300 122.760 46.440 122.960 ;
        RECT 48.510 122.900 48.830 122.960 ;
        RECT 53.660 122.960 67.690 123.100 ;
        RECT 53.660 122.760 53.800 122.960 ;
        RECT 67.370 122.900 67.690 122.960 ;
        RECT 68.765 123.100 69.055 123.145 ;
        RECT 70.130 123.100 70.450 123.160 ;
        RECT 68.765 122.960 70.450 123.100 ;
        RECT 68.765 122.915 69.055 122.960 ;
        RECT 70.130 122.900 70.450 122.960 ;
        RECT 73.825 123.100 74.115 123.145 ;
        RECT 76.110 123.100 76.430 123.160 ;
        RECT 79.420 123.100 79.560 123.300 ;
        RECT 80.725 123.255 81.015 123.300 ;
        RECT 73.825 122.960 79.560 123.100 ;
        RECT 80.265 123.100 80.555 123.145 ;
        RECT 81.950 123.100 82.240 123.145 ;
        RECT 80.265 122.960 82.240 123.100 ;
        RECT 73.825 122.915 74.115 122.960 ;
        RECT 76.110 122.900 76.430 122.960 ;
        RECT 80.265 122.915 80.555 122.960 ;
        RECT 81.950 122.915 82.240 122.960 ;
        RECT 46.300 122.620 53.800 122.760 ;
        RECT 39.325 122.575 39.615 122.620 ;
        RECT 41.150 122.560 41.470 122.620 ;
        RECT 54.030 122.560 54.350 122.820 ;
        RECT 59.550 122.560 59.870 122.820 ;
        RECT 62.310 122.760 62.630 122.820 ;
        RECT 66.450 122.760 66.770 122.820 ;
        RECT 62.310 122.620 66.770 122.760 ;
        RECT 62.310 122.560 62.630 122.620 ;
        RECT 66.450 122.560 66.770 122.620 ;
        RECT 66.925 122.760 67.215 122.805 ;
        RECT 72.430 122.760 72.750 122.820 ;
        RECT 66.925 122.620 72.750 122.760 ;
        RECT 66.925 122.575 67.215 122.620 ;
        RECT 72.430 122.560 72.750 122.620 ;
        RECT 73.350 122.560 73.670 122.820 ;
        RECT 77.030 122.760 77.350 122.820 ;
        RECT 80.710 122.760 81.030 122.820 ;
        RECT 77.030 122.620 81.030 122.760 ;
        RECT 77.030 122.560 77.350 122.620 ;
        RECT 80.710 122.560 81.030 122.620 ;
        RECT 83.470 122.760 83.790 122.820 ;
        RECT 87.625 122.760 87.915 122.805 ;
        RECT 83.470 122.620 87.915 122.760 ;
        RECT 83.470 122.560 83.790 122.620 ;
        RECT 87.625 122.575 87.915 122.620 ;
        RECT 100.010 122.450 100.880 125.790 ;
        RECT 108.930 125.490 116.850 125.500 ;
        RECT 105.160 125.480 116.850 125.490 ;
        RECT 101.540 125.360 116.850 125.480 ;
        RECT 101.540 125.350 116.875 125.360 ;
        RECT 101.500 125.230 116.875 125.350 ;
        RECT 101.500 125.120 105.500 125.230 ;
        RECT 101.110 124.780 101.340 125.070 ;
        RECT 101.560 124.780 105.450 125.120 ;
        RECT 105.660 124.780 105.890 125.070 ;
        RECT 101.110 123.410 105.890 124.780 ;
        RECT 101.110 123.110 101.340 123.410 ;
        RECT 105.660 123.110 105.890 123.410 ;
        RECT 101.500 122.830 105.500 123.060 ;
        RECT 101.750 122.600 105.320 122.830 ;
        RECT 101.750 122.450 105.440 122.600 ;
        RECT 12.100 121.940 89.840 122.420 ;
        RECT 100.010 122.170 105.440 122.450 ;
        RECT 106.690 122.280 107.310 125.230 ;
        RECT 108.875 125.130 116.875 125.230 ;
        RECT 108.930 125.120 116.850 125.130 ;
        RECT 108.440 124.420 108.670 125.080 ;
        RECT 109.450 124.420 110.450 124.510 ;
        RECT 117.080 124.420 117.310 125.080 ;
        RECT 108.440 123.600 117.310 124.420 ;
        RECT 108.440 123.120 108.670 123.600 ;
        RECT 109.450 123.510 110.450 123.600 ;
        RECT 117.080 123.120 117.310 123.600 ;
        RECT 108.875 122.840 116.875 123.070 ;
        RECT 17.690 121.740 18.010 121.800 ;
        RECT 19.070 121.785 19.390 121.800 ;
        RECT 19.070 121.740 19.455 121.785 ;
        RECT 16.400 121.600 19.455 121.740 ;
        RECT 16.400 121.105 16.540 121.600 ;
        RECT 17.690 121.540 18.010 121.600 ;
        RECT 19.070 121.555 19.455 121.600 ;
        RECT 20.005 121.740 20.295 121.785 ;
        RECT 20.910 121.740 21.230 121.800 ;
        RECT 20.005 121.600 21.230 121.740 ;
        RECT 20.005 121.555 20.295 121.600 ;
        RECT 19.070 121.540 19.390 121.555 ;
        RECT 20.910 121.540 21.230 121.600 ;
        RECT 24.130 121.740 24.450 121.800 ;
        RECT 25.510 121.740 25.830 121.800 ;
        RECT 24.130 121.600 39.540 121.740 ;
        RECT 24.130 121.540 24.450 121.600 ;
        RECT 25.510 121.540 25.830 121.600 ;
        RECT 18.165 121.215 18.455 121.445 ;
        RECT 33.790 121.400 34.110 121.460 ;
        RECT 39.400 121.445 39.540 121.600 ;
        RECT 55.410 121.540 55.730 121.800 ;
        RECT 62.325 121.740 62.615 121.785 ;
        RECT 61.020 121.600 62.615 121.740 ;
        RECT 38.405 121.400 38.695 121.445 ;
        RECT 33.790 121.260 38.695 121.400 ;
        RECT 16.325 120.875 16.615 121.105 ;
        RECT 16.785 120.875 17.075 121.105 ;
        RECT 17.705 121.060 17.995 121.105 ;
        RECT 18.240 121.060 18.380 121.215 ;
        RECT 33.790 121.200 34.110 121.260 ;
        RECT 38.405 121.215 38.695 121.260 ;
        RECT 39.325 121.215 39.615 121.445 ;
        RECT 48.050 121.400 48.370 121.460 ;
        RECT 41.240 121.260 48.370 121.400 ;
        RECT 21.830 121.060 22.150 121.120 ;
        RECT 17.705 120.920 22.150 121.060 ;
        RECT 17.705 120.875 17.995 120.920 ;
        RECT 16.860 120.040 17.000 120.875 ;
        RECT 21.830 120.860 22.150 120.920 ;
        RECT 25.985 121.060 26.275 121.105 ;
        RECT 26.890 121.060 27.210 121.120 ;
        RECT 25.985 120.920 27.210 121.060 ;
        RECT 25.985 120.875 26.275 120.920 ;
        RECT 26.890 120.860 27.210 120.920 ;
        RECT 27.825 121.060 28.115 121.105 ;
        RECT 28.730 121.060 29.050 121.120 ;
        RECT 27.825 120.920 29.050 121.060 ;
        RECT 27.825 120.875 28.115 120.920 ;
        RECT 28.730 120.860 29.050 120.920 ;
        RECT 29.205 120.875 29.495 121.105 ;
        RECT 18.610 120.720 18.930 120.780 ;
        RECT 22.305 120.720 22.595 120.765 ;
        RECT 22.750 120.720 23.070 120.780 ;
        RECT 29.280 120.720 29.420 120.875 ;
        RECT 30.110 120.860 30.430 121.120 ;
        RECT 32.425 120.875 32.715 121.105 ;
        RECT 35.630 121.060 35.950 121.120 ;
        RECT 32.960 120.920 35.950 121.060 ;
        RECT 31.490 120.720 31.810 120.780 ;
        RECT 18.610 120.580 23.070 120.720 ;
        RECT 18.610 120.520 18.930 120.580 ;
        RECT 22.305 120.535 22.595 120.580 ;
        RECT 22.750 120.520 23.070 120.580 ;
        RECT 23.760 120.580 31.810 120.720 ;
        RECT 17.705 120.380 17.995 120.425 ;
        RECT 18.150 120.380 18.470 120.440 ;
        RECT 23.760 120.425 23.900 120.580 ;
        RECT 31.490 120.520 31.810 120.580 ;
        RECT 17.705 120.240 18.470 120.380 ;
        RECT 17.705 120.195 17.995 120.240 ;
        RECT 18.150 120.180 18.470 120.240 ;
        RECT 23.685 120.195 23.975 120.425 ;
        RECT 27.810 120.380 28.130 120.440 ;
        RECT 26.980 120.240 28.130 120.380 ;
        RECT 19.085 120.040 19.375 120.085 ;
        RECT 22.290 120.040 22.610 120.100 ;
        RECT 26.980 120.085 27.120 120.240 ;
        RECT 27.810 120.180 28.130 120.240 ;
        RECT 28.745 120.380 29.035 120.425 ;
        RECT 30.110 120.380 30.430 120.440 ;
        RECT 31.950 120.380 32.270 120.440 ;
        RECT 28.745 120.240 30.430 120.380 ;
        RECT 28.745 120.195 29.035 120.240 ;
        RECT 30.110 120.180 30.430 120.240 ;
        RECT 30.660 120.240 32.270 120.380 ;
        RECT 32.500 120.380 32.640 120.875 ;
        RECT 32.960 120.765 33.100 120.920 ;
        RECT 35.630 120.860 35.950 120.920 ;
        RECT 36.105 121.060 36.395 121.105 ;
        RECT 38.850 121.060 39.170 121.120 ;
        RECT 41.240 121.105 41.380 121.260 ;
        RECT 48.050 121.200 48.370 121.260 ;
        RECT 49.860 121.400 50.150 121.445 ;
        RECT 61.020 121.400 61.160 121.600 ;
        RECT 62.325 121.555 62.615 121.600 ;
        RECT 67.370 121.740 67.690 121.800 ;
        RECT 82.090 121.740 82.410 121.800 ;
        RECT 83.025 121.740 83.315 121.785 ;
        RECT 67.370 121.600 76.340 121.740 ;
        RECT 67.370 121.540 67.690 121.600 ;
        RECT 49.860 121.260 61.160 121.400 ;
        RECT 61.850 121.400 62.170 121.460 ;
        RECT 75.205 121.400 75.495 121.445 ;
        RECT 61.850 121.260 75.495 121.400 ;
        RECT 49.860 121.215 50.150 121.260 ;
        RECT 61.850 121.200 62.170 121.260 ;
        RECT 75.205 121.215 75.495 121.260 ;
        RECT 36.105 120.920 39.170 121.060 ;
        RECT 36.105 120.875 36.395 120.920 ;
        RECT 38.850 120.860 39.170 120.920 ;
        RECT 41.165 120.875 41.455 121.105 ;
        RECT 42.500 121.060 42.790 121.105 ;
        RECT 48.970 121.060 49.290 121.120 ;
        RECT 42.500 120.920 49.290 121.060 ;
        RECT 42.500 120.875 42.790 120.920 ;
        RECT 48.970 120.860 49.290 120.920 ;
        RECT 58.630 120.860 58.950 121.120 ;
        RECT 59.550 120.860 59.870 121.120 ;
        RECT 60.470 120.860 60.790 121.120 ;
        RECT 60.945 120.875 61.235 121.105 ;
        RECT 32.885 120.535 33.175 120.765 ;
        RECT 34.250 120.520 34.570 120.780 ;
        RECT 36.565 120.535 36.855 120.765 ;
        RECT 37.025 120.720 37.315 120.765 ;
        RECT 37.930 120.720 38.250 120.780 ;
        RECT 37.025 120.580 38.250 120.720 ;
        RECT 37.025 120.535 37.315 120.580 ;
        RECT 33.330 120.380 33.650 120.440 ;
        RECT 36.640 120.380 36.780 120.535 ;
        RECT 37.930 120.520 38.250 120.580 ;
        RECT 42.045 120.720 42.335 120.765 ;
        RECT 43.235 120.720 43.525 120.765 ;
        RECT 45.755 120.720 46.045 120.765 ;
        RECT 42.045 120.580 46.045 120.720 ;
        RECT 42.045 120.535 42.335 120.580 ;
        RECT 43.235 120.535 43.525 120.580 ;
        RECT 45.755 120.535 46.045 120.580 ;
        RECT 48.050 120.720 48.370 120.780 ;
        RECT 48.525 120.720 48.815 120.765 ;
        RECT 48.050 120.580 48.815 120.720 ;
        RECT 48.050 120.520 48.370 120.580 ;
        RECT 48.525 120.535 48.815 120.580 ;
        RECT 49.405 120.720 49.695 120.765 ;
        RECT 50.595 120.720 50.885 120.765 ;
        RECT 53.115 120.720 53.405 120.765 ;
        RECT 58.720 120.720 58.860 120.860 ;
        RECT 49.405 120.580 53.405 120.720 ;
        RECT 49.405 120.535 49.695 120.580 ;
        RECT 50.595 120.535 50.885 120.580 ;
        RECT 53.115 120.535 53.405 120.580 ;
        RECT 53.660 120.580 58.860 120.720 ;
        RECT 59.090 120.720 59.410 120.780 ;
        RECT 61.020 120.720 61.160 120.875 ;
        RECT 61.390 120.860 61.710 121.120 ;
        RECT 64.150 120.860 64.470 121.120 ;
        RECT 71.510 121.060 71.830 121.120 ;
        RECT 72.950 121.060 73.240 121.105 ;
        RECT 71.510 120.920 73.240 121.060 ;
        RECT 71.510 120.860 71.830 120.920 ;
        RECT 72.950 120.875 73.240 120.920 ;
        RECT 74.285 120.875 74.575 121.105 ;
        RECT 74.745 120.875 75.035 121.105 ;
        RECT 75.665 121.060 75.955 121.105 ;
        RECT 76.200 121.060 76.340 121.600 ;
        RECT 82.090 121.600 83.315 121.740 ;
        RECT 82.090 121.540 82.410 121.600 ;
        RECT 83.025 121.555 83.315 121.600 ;
        RECT 86.690 121.740 87.010 121.800 ;
        RECT 87.625 121.740 87.915 121.785 ;
        RECT 86.690 121.600 87.915 121.740 ;
        RECT 83.100 121.400 83.240 121.555 ;
        RECT 86.690 121.540 87.010 121.600 ;
        RECT 87.625 121.555 87.915 121.600 ;
        RECT 100.010 121.710 105.450 122.170 ;
        RECT 84.405 121.400 84.695 121.445 ;
        RECT 83.100 121.260 84.695 121.400 ;
        RECT 84.405 121.215 84.695 121.260 ;
        RECT 85.310 121.200 85.630 121.460 ;
        RECT 85.785 121.400 86.075 121.445 ;
        RECT 88.990 121.400 89.310 121.460 ;
        RECT 85.785 121.260 89.310 121.400 ;
        RECT 85.785 121.215 86.075 121.260 ;
        RECT 88.990 121.200 89.310 121.260 ;
        RECT 75.665 120.920 76.340 121.060 ;
        RECT 77.460 121.060 77.750 121.105 ;
        RECT 79.330 121.060 79.650 121.120 ;
        RECT 77.460 120.920 79.650 121.060 ;
        RECT 75.665 120.875 75.955 120.920 ;
        RECT 77.460 120.875 77.750 120.920 ;
        RECT 59.090 120.580 61.160 120.720 ;
        RECT 69.695 120.720 69.985 120.765 ;
        RECT 72.215 120.720 72.505 120.765 ;
        RECT 73.405 120.720 73.695 120.765 ;
        RECT 69.695 120.580 73.695 120.720 ;
        RECT 37.470 120.380 37.790 120.440 ;
        RECT 32.500 120.240 37.790 120.380 ;
        RECT 16.860 119.900 22.610 120.040 ;
        RECT 19.085 119.855 19.375 119.900 ;
        RECT 22.290 119.840 22.610 119.900 ;
        RECT 26.905 119.855 27.195 120.085 ;
        RECT 29.665 120.040 29.955 120.085 ;
        RECT 30.660 120.040 30.800 120.240 ;
        RECT 31.950 120.180 32.270 120.240 ;
        RECT 33.330 120.180 33.650 120.240 ;
        RECT 37.470 120.180 37.790 120.240 ;
        RECT 41.650 120.380 41.940 120.425 ;
        RECT 43.750 120.380 44.040 120.425 ;
        RECT 45.320 120.380 45.610 120.425 ;
        RECT 41.650 120.240 45.610 120.380 ;
        RECT 41.650 120.195 41.940 120.240 ;
        RECT 43.750 120.195 44.040 120.240 ;
        RECT 45.320 120.195 45.610 120.240 ;
        RECT 49.010 120.380 49.300 120.425 ;
        RECT 51.110 120.380 51.400 120.425 ;
        RECT 52.680 120.380 52.970 120.425 ;
        RECT 49.010 120.240 52.970 120.380 ;
        RECT 49.010 120.195 49.300 120.240 ;
        RECT 51.110 120.195 51.400 120.240 ;
        RECT 52.680 120.195 52.970 120.240 ;
        RECT 29.665 119.900 30.800 120.040 ;
        RECT 29.665 119.855 29.955 119.900 ;
        RECT 31.030 119.840 31.350 120.100 ;
        RECT 34.710 119.840 35.030 120.100 ;
        RECT 48.065 120.040 48.355 120.085 ;
        RECT 53.660 120.040 53.800 120.580 ;
        RECT 59.090 120.520 59.410 120.580 ;
        RECT 69.695 120.535 69.985 120.580 ;
        RECT 72.215 120.535 72.505 120.580 ;
        RECT 73.405 120.535 73.695 120.580 ;
        RECT 54.030 120.380 54.350 120.440 ;
        RECT 67.385 120.380 67.675 120.425 ;
        RECT 68.750 120.380 69.070 120.440 ;
        RECT 54.030 120.240 69.070 120.380 ;
        RECT 54.030 120.180 54.350 120.240 ;
        RECT 67.385 120.195 67.675 120.240 ;
        RECT 68.750 120.180 69.070 120.240 ;
        RECT 70.130 120.380 70.420 120.425 ;
        RECT 71.700 120.380 71.990 120.425 ;
        RECT 73.800 120.380 74.090 120.425 ;
        RECT 70.130 120.240 74.090 120.380 ;
        RECT 70.130 120.195 70.420 120.240 ;
        RECT 71.700 120.195 71.990 120.240 ;
        RECT 73.800 120.195 74.090 120.240 ;
        RECT 48.065 119.900 53.800 120.040 ;
        RECT 48.065 119.855 48.355 119.900 ;
        RECT 55.870 119.840 56.190 120.100 ;
        RECT 56.790 120.040 57.110 120.100 ;
        RECT 65.530 120.040 65.850 120.100 ;
        RECT 56.790 119.900 65.850 120.040 ;
        RECT 74.360 120.040 74.500 120.875 ;
        RECT 74.820 120.720 74.960 120.875 ;
        RECT 79.330 120.860 79.650 120.920 ;
        RECT 86.705 121.060 86.995 121.105 ;
        RECT 88.070 121.060 88.390 121.120 ;
        RECT 86.705 120.920 88.390 121.060 ;
        RECT 86.705 120.875 86.995 120.920 ;
        RECT 88.070 120.860 88.390 120.920 ;
        RECT 74.820 120.580 75.880 120.720 ;
        RECT 75.740 120.440 75.880 120.580 ;
        RECT 76.110 120.520 76.430 120.780 ;
        RECT 77.005 120.720 77.295 120.765 ;
        RECT 78.195 120.720 78.485 120.765 ;
        RECT 80.715 120.720 81.005 120.765 ;
        RECT 77.005 120.580 81.005 120.720 ;
        RECT 77.005 120.535 77.295 120.580 ;
        RECT 78.195 120.535 78.485 120.580 ;
        RECT 80.715 120.535 81.005 120.580 ;
        RECT 75.650 120.180 75.970 120.440 ;
        RECT 76.200 120.040 76.340 120.520 ;
        RECT 76.610 120.380 76.900 120.425 ;
        RECT 78.710 120.380 79.000 120.425 ;
        RECT 80.280 120.380 80.570 120.425 ;
        RECT 76.610 120.240 80.570 120.380 ;
        RECT 76.610 120.195 76.900 120.240 ;
        RECT 78.710 120.195 79.000 120.240 ;
        RECT 80.280 120.195 80.570 120.240 ;
        RECT 81.630 120.380 81.950 120.440 ;
        RECT 83.485 120.380 83.775 120.425 ;
        RECT 81.630 120.240 83.775 120.380 ;
        RECT 81.630 120.180 81.950 120.240 ;
        RECT 83.485 120.195 83.775 120.240 ;
        RECT 100.010 120.360 102.050 121.710 ;
        RECT 103.800 121.700 105.450 121.710 ;
        RECT 102.490 120.430 103.490 121.150 ;
        RECT 103.800 120.890 104.110 121.700 ;
        RECT 104.570 121.420 105.450 121.700 ;
        RECT 105.690 121.880 107.310 122.280 ;
        RECT 108.960 121.930 116.830 122.840 ;
        RECT 104.510 121.190 105.510 121.420 ;
        RECT 105.690 121.230 106.040 121.880 ;
        RECT 106.690 121.870 107.310 121.880 ;
        RECT 108.875 121.700 116.875 121.930 ;
        RECT 108.960 121.690 116.830 121.700 ;
        RECT 104.570 120.980 105.450 121.000 ;
        RECT 103.840 120.600 104.110 120.890 ;
        RECT 104.510 120.750 105.510 120.980 ;
        RECT 105.670 120.940 106.040 121.230 ;
        RECT 105.700 120.880 106.040 120.940 ;
        RECT 106.800 121.550 107.560 121.600 ;
        RECT 108.440 121.550 108.670 121.650 ;
        RECT 106.800 121.340 108.670 121.550 ;
        RECT 117.080 121.340 117.310 121.650 ;
        RECT 106.800 120.920 109.340 121.340 ;
        RECT 116.710 120.920 117.310 121.340 ;
        RECT 104.570 120.600 105.450 120.750 ;
        RECT 104.580 120.430 105.310 120.600 ;
        RECT 77.030 120.040 77.350 120.100 ;
        RECT 74.360 119.900 77.350 120.040 ;
        RECT 56.790 119.840 57.110 119.900 ;
        RECT 65.530 119.840 65.850 119.900 ;
        RECT 77.030 119.840 77.350 119.900 ;
        RECT 12.100 119.220 89.840 119.700 ;
        RECT 23.210 118.820 23.530 119.080 ;
        RECT 28.730 119.020 29.050 119.080 ;
        RECT 31.490 119.020 31.810 119.080 ;
        RECT 28.730 118.880 31.810 119.020 ;
        RECT 28.730 118.820 29.050 118.880 ;
        RECT 31.490 118.820 31.810 118.880 ;
        RECT 48.065 119.020 48.355 119.065 ;
        RECT 48.510 119.020 48.830 119.080 ;
        RECT 48.065 118.880 48.830 119.020 ;
        RECT 48.065 118.835 48.355 118.880 ;
        RECT 48.510 118.820 48.830 118.880 ;
        RECT 48.970 119.020 49.290 119.080 ;
        RECT 51.285 119.020 51.575 119.065 ;
        RECT 48.970 118.880 51.575 119.020 ;
        RECT 48.970 118.820 49.290 118.880 ;
        RECT 51.285 118.835 51.575 118.880 ;
        RECT 58.185 119.020 58.475 119.065 ;
        RECT 60.470 119.020 60.790 119.080 ;
        RECT 58.185 118.880 60.790 119.020 ;
        RECT 58.185 118.835 58.475 118.880 ;
        RECT 60.470 118.820 60.790 118.880 ;
        RECT 64.610 119.020 64.930 119.080 ;
        RECT 66.465 119.020 66.755 119.065 ;
        RECT 64.610 118.880 66.755 119.020 ;
        RECT 64.610 118.820 64.930 118.880 ;
        RECT 66.465 118.835 66.755 118.880 ;
        RECT 73.810 119.020 74.130 119.080 ;
        RECT 74.285 119.020 74.575 119.065 ;
        RECT 73.810 118.880 74.575 119.020 ;
        RECT 73.810 118.820 74.130 118.880 ;
        RECT 74.285 118.835 74.575 118.880 ;
        RECT 74.730 118.820 75.050 119.080 ;
        RECT 78.410 119.020 78.730 119.080 ;
        RECT 81.170 119.020 81.490 119.080 ;
        RECT 78.410 118.880 81.490 119.020 ;
        RECT 78.410 118.820 78.730 118.880 ;
        RECT 81.170 118.820 81.490 118.880 ;
        RECT 23.300 118.680 23.440 118.820 ;
        RECT 22.840 118.540 23.440 118.680 ;
        RECT 24.605 118.680 24.895 118.725 ;
        RECT 28.270 118.680 28.590 118.740 ;
        RECT 31.950 118.680 32.270 118.740 ;
        RECT 24.605 118.540 32.270 118.680 ;
        RECT 22.840 118.045 22.980 118.540 ;
        RECT 24.605 118.495 24.895 118.540 ;
        RECT 28.270 118.480 28.590 118.540 ;
        RECT 31.950 118.480 32.270 118.540 ;
        RECT 38.390 118.680 38.710 118.740 ;
        RECT 41.650 118.680 41.940 118.725 ;
        RECT 43.750 118.680 44.040 118.725 ;
        RECT 45.320 118.680 45.610 118.725 ;
        RECT 38.390 118.540 41.380 118.680 ;
        RECT 38.390 118.480 38.710 118.540 ;
        RECT 23.210 118.140 23.530 118.400 ;
        RECT 29.650 118.340 29.970 118.400 ;
        RECT 28.360 118.200 29.970 118.340 ;
        RECT 22.765 117.815 23.055 118.045 ;
        RECT 26.430 117.800 26.750 118.060 ;
        RECT 27.185 118.000 27.475 118.045 ;
        RECT 28.360 118.000 28.500 118.200 ;
        RECT 29.650 118.140 29.970 118.200 ;
        RECT 35.630 118.340 35.950 118.400 ;
        RECT 41.240 118.385 41.380 118.540 ;
        RECT 41.650 118.540 45.610 118.680 ;
        RECT 41.650 118.495 41.940 118.540 ;
        RECT 43.750 118.495 44.040 118.540 ;
        RECT 45.320 118.495 45.610 118.540 ;
        RECT 59.550 118.680 59.870 118.740 ;
        RECT 65.990 118.680 66.310 118.740 ;
        RECT 71.510 118.680 71.830 118.740 ;
        RECT 74.820 118.680 74.960 118.820 ;
        RECT 59.550 118.540 68.520 118.680 ;
        RECT 59.550 118.480 59.870 118.540 ;
        RECT 65.990 118.480 66.310 118.540 ;
        RECT 35.630 118.200 40.000 118.340 ;
        RECT 35.630 118.140 35.950 118.200 ;
        RECT 27.185 117.860 28.500 118.000 ;
        RECT 28.975 118.000 29.265 118.045 ;
        RECT 30.570 118.000 30.890 118.060 ;
        RECT 28.975 117.860 30.890 118.000 ;
        RECT 27.185 117.815 27.475 117.860 ;
        RECT 28.975 117.815 29.265 117.860 ;
        RECT 30.570 117.800 30.890 117.860 ;
        RECT 33.790 118.000 34.110 118.060 ;
        RECT 38.390 118.000 38.710 118.060 ;
        RECT 39.860 118.045 40.000 118.200 ;
        RECT 41.165 118.155 41.455 118.385 ;
        RECT 42.045 118.340 42.335 118.385 ;
        RECT 43.235 118.340 43.525 118.385 ;
        RECT 45.755 118.340 46.045 118.385 ;
        RECT 42.045 118.200 46.045 118.340 ;
        RECT 42.045 118.155 42.335 118.200 ;
        RECT 43.235 118.155 43.525 118.200 ;
        RECT 45.755 118.155 46.045 118.200 ;
        RECT 53.570 118.340 53.890 118.400 ;
        RECT 54.045 118.340 54.335 118.385 ;
        RECT 53.570 118.200 54.335 118.340 ;
        RECT 53.570 118.140 53.890 118.200 ;
        RECT 54.045 118.155 54.335 118.200 ;
        RECT 58.630 118.340 58.950 118.400 ;
        RECT 59.105 118.340 59.395 118.385 ;
        RECT 66.910 118.340 67.230 118.400 ;
        RECT 68.380 118.385 68.520 118.540 ;
        RECT 71.140 118.540 74.960 118.680 ;
        RECT 58.630 118.200 59.395 118.340 ;
        RECT 58.630 118.140 58.950 118.200 ;
        RECT 59.105 118.155 59.395 118.200 ;
        RECT 60.100 118.200 67.230 118.340 ;
        RECT 33.790 117.860 38.710 118.000 ;
        RECT 33.790 117.800 34.110 117.860 ;
        RECT 38.390 117.800 38.710 117.860 ;
        RECT 39.785 117.815 40.075 118.045 ;
        RECT 40.690 118.000 41.010 118.060 ;
        RECT 53.110 118.000 53.430 118.060 ;
        RECT 55.425 118.000 55.715 118.045 ;
        RECT 40.690 117.860 45.520 118.000 ;
        RECT 40.690 117.800 41.010 117.860 ;
        RECT 25.970 117.660 26.290 117.720 ;
        RECT 27.825 117.660 28.115 117.705 ;
        RECT 25.970 117.520 28.115 117.660 ;
        RECT 25.970 117.460 26.290 117.520 ;
        RECT 27.825 117.475 28.115 117.520 ;
        RECT 28.285 117.660 28.575 117.705 ;
        RECT 30.110 117.660 30.430 117.720 ;
        RECT 28.285 117.520 30.430 117.660 ;
        RECT 28.285 117.475 28.575 117.520 ;
        RECT 30.110 117.460 30.430 117.520 ;
        RECT 34.725 117.660 35.015 117.705 ;
        RECT 41.610 117.660 41.930 117.720 ;
        RECT 34.725 117.520 41.930 117.660 ;
        RECT 34.725 117.475 35.015 117.520 ;
        RECT 41.610 117.460 41.930 117.520 ;
        RECT 42.500 117.660 42.790 117.705 ;
        RECT 44.370 117.660 44.690 117.720 ;
        RECT 42.500 117.520 44.690 117.660 ;
        RECT 45.380 117.660 45.520 117.860 ;
        RECT 53.110 117.860 55.715 118.000 ;
        RECT 53.110 117.800 53.430 117.860 ;
        RECT 55.425 117.815 55.715 117.860 ;
        RECT 55.885 117.815 56.175 118.045 ;
        RECT 56.330 118.000 56.650 118.060 ;
        RECT 56.805 118.000 57.095 118.045 ;
        RECT 56.330 117.860 57.095 118.000 ;
        RECT 45.750 117.660 46.070 117.720 ;
        RECT 45.380 117.520 46.070 117.660 ;
        RECT 42.500 117.475 42.790 117.520 ;
        RECT 44.370 117.460 44.690 117.520 ;
        RECT 45.750 117.460 46.070 117.520 ;
        RECT 54.030 117.660 54.350 117.720 ;
        RECT 55.960 117.660 56.100 117.815 ;
        RECT 56.330 117.800 56.650 117.860 ;
        RECT 56.805 117.815 57.095 117.860 ;
        RECT 57.265 118.000 57.555 118.045 ;
        RECT 58.170 118.000 58.490 118.060 ;
        RECT 60.100 118.045 60.240 118.200 ;
        RECT 66.910 118.140 67.230 118.200 ;
        RECT 68.305 118.155 68.595 118.385 ;
        RECT 68.750 118.140 69.070 118.400 ;
        RECT 71.140 118.385 71.280 118.540 ;
        RECT 71.510 118.480 71.830 118.540 ;
        RECT 71.065 118.155 71.355 118.385 ;
        RECT 71.985 118.340 72.275 118.385 ;
        RECT 77.490 118.340 77.810 118.400 ;
        RECT 71.985 118.200 77.810 118.340 ;
        RECT 71.985 118.155 72.275 118.200 ;
        RECT 77.490 118.140 77.810 118.200 ;
        RECT 77.950 118.340 78.270 118.400 ;
        RECT 80.250 118.340 80.570 118.400 ;
        RECT 77.950 118.200 80.570 118.340 ;
        RECT 77.950 118.140 78.270 118.200 ;
        RECT 80.250 118.140 80.570 118.200 ;
        RECT 57.265 117.860 58.490 118.000 ;
        RECT 57.265 117.815 57.555 117.860 ;
        RECT 58.170 117.800 58.490 117.860 ;
        RECT 60.025 117.815 60.315 118.045 ;
        RECT 65.070 118.000 65.390 118.060 ;
        RECT 67.385 118.000 67.675 118.045 ;
        RECT 65.070 117.860 67.675 118.000 ;
        RECT 65.070 117.800 65.390 117.860 ;
        RECT 67.385 117.815 67.675 117.860 ;
        RECT 67.830 117.800 68.150 118.060 ;
        RECT 72.445 118.000 72.735 118.045 ;
        RECT 73.350 118.000 73.670 118.060 ;
        RECT 72.445 117.860 73.670 118.000 ;
        RECT 72.445 117.815 72.735 117.860 ;
        RECT 73.350 117.800 73.670 117.860 ;
        RECT 76.125 118.000 76.415 118.045 ;
        RECT 82.090 118.000 82.410 118.060 ;
        RECT 76.125 117.860 82.410 118.000 ;
        RECT 76.125 117.815 76.415 117.860 ;
        RECT 82.090 117.800 82.410 117.860 ;
        RECT 83.470 117.800 83.790 118.060 ;
        RECT 84.865 118.000 85.155 118.045 ;
        RECT 86.230 118.000 86.550 118.060 ;
        RECT 84.865 117.860 86.550 118.000 ;
        RECT 84.865 117.815 85.155 117.860 ;
        RECT 86.230 117.800 86.550 117.860 ;
        RECT 86.690 117.800 87.010 118.060 ;
        RECT 54.030 117.520 56.100 117.660 ;
        RECT 57.710 117.660 58.030 117.720 ;
        RECT 61.405 117.660 61.695 117.705 ;
        RECT 57.710 117.520 61.695 117.660 ;
        RECT 54.030 117.460 54.350 117.520 ;
        RECT 57.710 117.460 58.030 117.520 ;
        RECT 61.405 117.475 61.695 117.520 ;
        RECT 64.150 117.660 64.470 117.720 ;
        RECT 65.545 117.660 65.835 117.705 ;
        RECT 66.450 117.660 66.770 117.720 ;
        RECT 72.890 117.660 73.210 117.720 ;
        RECT 77.045 117.660 77.335 117.705 ;
        RECT 64.150 117.520 66.770 117.660 ;
        RECT 29.650 117.120 29.970 117.380 ;
        RECT 40.230 117.120 40.550 117.380 ;
        RECT 52.190 117.320 52.510 117.380 ;
        RECT 53.125 117.320 53.415 117.365 ;
        RECT 52.190 117.180 53.415 117.320 ;
        RECT 52.190 117.120 52.510 117.180 ;
        RECT 53.125 117.135 53.415 117.180 ;
        RECT 53.585 117.320 53.875 117.365 ;
        RECT 55.870 117.320 56.190 117.380 ;
        RECT 53.585 117.180 56.190 117.320 ;
        RECT 53.585 117.135 53.875 117.180 ;
        RECT 55.870 117.120 56.190 117.180 ;
        RECT 60.470 117.320 60.790 117.380 ;
        RECT 60.945 117.320 61.235 117.365 ;
        RECT 60.470 117.180 61.235 117.320 ;
        RECT 61.480 117.320 61.620 117.475 ;
        RECT 64.150 117.460 64.470 117.520 ;
        RECT 65.545 117.475 65.835 117.520 ;
        RECT 66.450 117.460 66.770 117.520 ;
        RECT 68.610 117.520 77.335 117.660 ;
        RECT 68.610 117.320 68.750 117.520 ;
        RECT 72.890 117.460 73.210 117.520 ;
        RECT 77.045 117.475 77.335 117.520 ;
        RECT 78.870 117.660 79.190 117.720 ;
        RECT 80.725 117.660 81.015 117.705 ;
        RECT 83.010 117.660 83.330 117.720 ;
        RECT 78.870 117.520 81.015 117.660 ;
        RECT 78.870 117.460 79.190 117.520 ;
        RECT 80.725 117.475 81.015 117.520 ;
        RECT 81.260 117.520 83.330 117.660 ;
        RECT 61.480 117.180 68.750 117.320 ;
        RECT 75.205 117.320 75.495 117.365 ;
        RECT 81.260 117.320 81.400 117.520 ;
        RECT 83.010 117.460 83.330 117.520 ;
        RECT 75.205 117.180 81.400 117.320 ;
        RECT 60.470 117.120 60.790 117.180 ;
        RECT 60.945 117.135 61.235 117.180 ;
        RECT 75.205 117.135 75.495 117.180 ;
        RECT 82.550 117.120 82.870 117.380 ;
        RECT 85.770 117.120 86.090 117.380 ;
        RECT 87.610 117.120 87.930 117.380 ;
        RECT 12.100 116.500 89.840 116.980 ;
        RECT 100.010 116.810 100.780 120.360 ;
        RECT 102.460 119.310 105.310 120.430 ;
        RECT 105.700 120.130 106.050 120.880 ;
        RECT 106.800 120.760 108.670 120.920 ;
        RECT 106.800 120.710 107.560 120.760 ;
        RECT 108.440 120.690 108.670 120.760 ;
        RECT 117.080 120.690 117.310 120.920 ;
        RECT 108.875 120.410 116.875 120.640 ;
        RECT 105.700 120.070 105.990 120.130 ;
        RECT 105.610 119.950 105.990 120.070 ;
        RECT 108.970 120.010 116.830 120.410 ;
        RECT 117.640 120.010 118.600 129.490 ;
        RECT 119.930 129.680 120.770 131.810 ;
        RECT 126.430 131.390 127.680 131.830 ;
        RECT 137.600 131.810 138.460 133.870 ;
        RECT 124.370 131.380 129.610 131.390 ;
        RECT 121.420 131.280 136.720 131.380 ;
        RECT 121.420 131.270 136.755 131.280 ;
        RECT 121.380 131.150 136.755 131.270 ;
        RECT 121.380 131.040 125.380 131.150 ;
        RECT 126.430 131.070 128.170 131.150 ;
        RECT 128.750 131.070 136.755 131.150 ;
        RECT 126.430 130.990 127.680 131.070 ;
        RECT 128.755 131.050 136.755 131.070 ;
        RECT 120.990 130.740 121.220 130.990 ;
        RECT 125.540 130.850 125.770 130.990 ;
        RECT 128.320 130.850 128.550 131.000 ;
        RECT 125.540 130.740 128.550 130.850 ;
        RECT 136.960 130.740 137.190 131.000 ;
        RECT 120.990 130.300 137.190 130.740 ;
        RECT 120.990 130.030 121.220 130.300 ;
        RECT 125.540 130.270 137.190 130.300 ;
        RECT 125.540 130.180 128.550 130.270 ;
        RECT 125.540 130.030 125.770 130.180 ;
        RECT 128.320 130.040 128.550 130.180 ;
        RECT 136.960 130.040 137.190 130.270 ;
        RECT 121.380 129.750 125.380 129.980 ;
        RECT 128.755 129.770 136.755 129.990 ;
        RECT 137.520 129.770 138.480 131.810 ;
        RECT 128.755 129.760 138.480 129.770 ;
        RECT 121.380 129.680 125.370 129.750 ;
        RECT 119.930 129.570 125.370 129.680 ;
        RECT 128.810 129.600 138.480 129.760 ;
        RECT 119.930 129.480 123.060 129.570 ;
        RECT 136.550 129.550 138.480 129.600 ;
        RECT 119.930 126.210 120.770 129.480 ;
        RECT 124.410 129.020 129.660 129.030 ;
        RECT 124.410 128.910 136.720 129.020 ;
        RECT 121.440 128.850 136.720 128.910 ;
        RECT 121.440 128.840 136.755 128.850 ;
        RECT 121.380 128.710 136.755 128.840 ;
        RECT 121.380 128.700 126.540 128.710 ;
        RECT 121.380 128.610 125.380 128.700 ;
        RECT 128.755 128.620 136.755 128.710 ;
        RECT 128.840 128.610 136.730 128.620 ;
        RECT 120.990 128.250 121.220 128.560 ;
        RECT 121.440 128.250 125.340 128.610 ;
        RECT 125.540 128.250 125.770 128.560 ;
        RECT 120.990 126.910 125.770 128.250 ;
        RECT 120.990 126.600 121.220 126.910 ;
        RECT 125.540 126.600 125.770 126.910 ;
        RECT 128.320 128.030 128.550 128.570 ;
        RECT 129.360 128.030 130.370 128.060 ;
        RECT 136.960 128.030 137.190 128.570 ;
        RECT 128.320 127.130 137.190 128.030 ;
        RECT 128.320 126.610 128.550 127.130 ;
        RECT 129.360 127.060 130.370 127.130 ;
        RECT 136.960 126.610 137.190 127.130 ;
        RECT 121.380 126.320 125.380 126.550 ;
        RECT 128.755 126.330 136.755 126.560 ;
        RECT 119.930 126.170 121.060 126.210 ;
        RECT 119.930 126.090 121.300 126.170 ;
        RECT 121.670 126.100 125.330 126.320 ;
        RECT 121.670 126.090 123.110 126.100 ;
        RECT 119.930 126.050 123.110 126.090 ;
        RECT 119.930 125.960 122.620 126.050 ;
        RECT 128.820 126.040 136.710 126.330 ;
        RECT 119.930 125.900 121.950 125.960 ;
        RECT 119.930 125.850 121.700 125.900 ;
        RECT 119.930 122.510 120.770 125.850 ;
        RECT 128.810 125.550 136.730 125.560 ;
        RECT 125.040 125.540 136.730 125.550 ;
        RECT 121.420 125.420 136.730 125.540 ;
        RECT 121.420 125.410 136.755 125.420 ;
        RECT 121.380 125.290 136.755 125.410 ;
        RECT 121.380 125.180 125.380 125.290 ;
        RECT 120.990 124.840 121.220 125.130 ;
        RECT 121.440 124.840 125.330 125.180 ;
        RECT 125.540 124.840 125.770 125.130 ;
        RECT 120.990 123.470 125.770 124.840 ;
        RECT 120.990 123.170 121.220 123.470 ;
        RECT 125.540 123.170 125.770 123.470 ;
        RECT 121.380 122.890 125.380 123.120 ;
        RECT 121.630 122.660 125.200 122.890 ;
        RECT 121.630 122.510 125.320 122.660 ;
        RECT 119.930 122.230 125.320 122.510 ;
        RECT 126.570 122.340 127.190 125.290 ;
        RECT 128.755 125.190 136.755 125.290 ;
        RECT 128.810 125.180 136.730 125.190 ;
        RECT 128.320 124.480 128.550 125.140 ;
        RECT 129.330 124.480 130.330 124.570 ;
        RECT 136.960 124.480 137.190 125.140 ;
        RECT 128.320 123.660 137.190 124.480 ;
        RECT 128.320 123.180 128.550 123.660 ;
        RECT 129.330 123.570 130.330 123.660 ;
        RECT 136.960 123.180 137.190 123.660 ;
        RECT 128.755 122.900 136.755 123.130 ;
        RECT 119.930 121.770 125.330 122.230 ;
        RECT 119.930 120.430 121.930 121.770 ;
        RECT 123.680 121.760 125.330 121.770 ;
        RECT 122.370 120.490 123.370 121.210 ;
        RECT 123.680 120.950 123.990 121.760 ;
        RECT 124.450 121.480 125.330 121.760 ;
        RECT 125.570 121.940 127.190 122.340 ;
        RECT 128.840 121.990 136.710 122.900 ;
        RECT 124.390 121.250 125.390 121.480 ;
        RECT 125.570 121.290 125.920 121.940 ;
        RECT 126.570 121.930 127.190 121.940 ;
        RECT 128.755 121.760 136.755 121.990 ;
        RECT 128.840 121.750 136.710 121.760 ;
        RECT 124.450 121.040 125.330 121.060 ;
        RECT 123.720 120.660 123.990 120.950 ;
        RECT 124.390 120.810 125.390 121.040 ;
        RECT 125.550 121.000 125.920 121.290 ;
        RECT 125.580 120.940 125.920 121.000 ;
        RECT 126.680 121.610 127.440 121.660 ;
        RECT 128.320 121.610 128.550 121.710 ;
        RECT 126.680 121.400 128.550 121.610 ;
        RECT 136.960 121.400 137.190 121.710 ;
        RECT 126.680 120.980 129.220 121.400 ;
        RECT 136.590 120.980 137.190 121.400 ;
        RECT 124.450 120.660 125.330 120.810 ;
        RECT 124.460 120.490 125.190 120.660 ;
        RECT 102.400 119.080 105.400 119.310 ;
        RECT 105.610 119.120 105.950 119.950 ;
        RECT 107.960 119.940 118.600 120.010 ;
        RECT 102.450 119.050 105.310 119.080 ;
        RECT 102.450 119.030 103.620 119.050 ;
        RECT 104.580 119.040 105.310 119.050 ;
        RECT 102.400 118.640 105.400 118.870 ;
        RECT 105.605 118.830 105.950 119.120 ;
        RECT 106.140 118.900 118.600 119.940 ;
        RECT 120.000 120.420 121.930 120.430 ;
        RECT 106.140 118.880 118.560 118.900 ;
        RECT 105.610 118.720 105.950 118.830 ;
        RECT 106.180 118.870 111.850 118.880 ;
        RECT 112.850 118.870 118.560 118.880 ;
        RECT 102.490 118.470 105.350 118.640 ;
        RECT 106.180 118.470 106.610 118.870 ;
        RECT 102.460 118.100 106.610 118.470 ;
        RECT 100.000 116.780 100.780 116.810 ;
        RECT 24.590 116.300 24.910 116.360 ;
        RECT 21.460 116.160 24.910 116.300 ;
        RECT 10.790 115.620 11.110 115.680 ;
        RECT 13.565 115.620 13.855 115.665 ;
        RECT 10.790 115.480 13.855 115.620 ;
        RECT 10.790 115.420 11.110 115.480 ;
        RECT 13.565 115.435 13.855 115.480 ;
        RECT 20.925 115.620 21.215 115.665 ;
        RECT 21.460 115.620 21.600 116.160 ;
        RECT 24.590 116.100 24.910 116.160 ;
        RECT 25.970 116.100 26.290 116.360 ;
        RECT 32.870 116.100 33.190 116.360 ;
        RECT 33.330 116.100 33.650 116.360 ;
        RECT 44.370 116.100 44.690 116.360 ;
        RECT 60.930 116.100 61.250 116.360 ;
        RECT 66.910 116.300 67.230 116.360 ;
        RECT 68.290 116.300 68.610 116.360 ;
        RECT 66.910 116.160 68.610 116.300 ;
        RECT 66.910 116.100 67.230 116.160 ;
        RECT 68.290 116.100 68.610 116.160 ;
        RECT 77.030 116.300 77.350 116.360 ;
        RECT 78.870 116.300 79.190 116.360 ;
        RECT 77.030 116.160 79.190 116.300 ;
        RECT 77.030 116.100 77.350 116.160 ;
        RECT 78.870 116.100 79.190 116.160 ;
        RECT 79.330 116.100 79.650 116.360 ;
        RECT 83.945 116.300 84.235 116.345 ;
        RECT 86.690 116.300 87.010 116.360 ;
        RECT 83.945 116.160 87.010 116.300 ;
        RECT 83.945 116.115 84.235 116.160 ;
        RECT 86.690 116.100 87.010 116.160 ;
        RECT 24.145 115.960 24.435 116.005 ;
        RECT 22.380 115.820 24.435 115.960 ;
        RECT 22.380 115.680 22.520 115.820 ;
        RECT 24.145 115.775 24.435 115.820 ;
        RECT 30.125 115.960 30.415 116.005 ;
        RECT 31.490 115.960 31.810 116.020 ;
        RECT 30.125 115.820 31.810 115.960 ;
        RECT 30.125 115.775 30.415 115.820 ;
        RECT 31.490 115.760 31.810 115.820 ;
        RECT 33.930 115.960 34.220 116.005 ;
        RECT 34.710 115.960 35.030 116.020 ;
        RECT 33.930 115.820 35.030 115.960 ;
        RECT 33.930 115.775 34.220 115.820 ;
        RECT 34.710 115.760 35.030 115.820 ;
        RECT 35.630 115.960 35.950 116.020 ;
        RECT 37.025 115.960 37.315 116.005 ;
        RECT 37.470 115.960 37.790 116.020 ;
        RECT 40.690 115.960 41.010 116.020 ;
        RECT 35.630 115.820 41.010 115.960 ;
        RECT 35.630 115.760 35.950 115.820 ;
        RECT 37.025 115.775 37.315 115.820 ;
        RECT 37.470 115.760 37.790 115.820 ;
        RECT 40.690 115.760 41.010 115.820 ;
        RECT 41.610 115.960 41.930 116.020 ;
        RECT 47.590 115.960 47.910 116.020 ;
        RECT 57.710 115.960 58.030 116.020 ;
        RECT 41.610 115.820 58.030 115.960 ;
        RECT 41.610 115.760 41.930 115.820 ;
        RECT 47.590 115.760 47.910 115.820 ;
        RECT 57.710 115.760 58.030 115.820 ;
        RECT 58.630 115.960 58.950 116.020 ;
        RECT 62.770 115.960 63.090 116.020 ;
        RECT 67.830 115.960 68.150 116.020 ;
        RECT 58.630 115.820 63.090 115.960 ;
        RECT 58.630 115.760 58.950 115.820 ;
        RECT 62.770 115.760 63.090 115.820 ;
        RECT 66.080 115.820 68.150 115.960 ;
        RECT 20.925 115.480 21.600 115.620 ;
        RECT 21.845 115.620 22.135 115.665 ;
        RECT 22.290 115.620 22.610 115.680 ;
        RECT 21.845 115.480 22.610 115.620 ;
        RECT 20.925 115.435 21.215 115.480 ;
        RECT 21.845 115.435 22.135 115.480 ;
        RECT 22.290 115.420 22.610 115.480 ;
        RECT 22.765 115.435 23.055 115.665 ;
        RECT 23.210 115.620 23.530 115.680 ;
        RECT 23.685 115.620 23.975 115.665 ;
        RECT 23.210 115.480 23.975 115.620 ;
        RECT 21.385 115.280 21.675 115.325 ;
        RECT 22.840 115.280 22.980 115.435 ;
        RECT 23.210 115.420 23.530 115.480 ;
        RECT 23.685 115.435 23.975 115.480 ;
        RECT 24.605 115.435 24.895 115.665 ;
        RECT 25.970 115.620 26.290 115.680 ;
        RECT 26.905 115.620 27.195 115.665 ;
        RECT 25.970 115.480 27.195 115.620 ;
        RECT 21.385 115.140 22.980 115.280 ;
        RECT 24.680 115.280 24.820 115.435 ;
        RECT 25.970 115.420 26.290 115.480 ;
        RECT 26.905 115.435 27.195 115.480 ;
        RECT 27.365 115.435 27.655 115.665 ;
        RECT 27.440 115.280 27.580 115.435 ;
        RECT 28.270 115.420 28.590 115.680 ;
        RECT 28.730 115.420 29.050 115.680 ;
        RECT 31.030 115.620 31.350 115.680 ;
        RECT 31.030 115.480 32.640 115.620 ;
        RECT 31.030 115.420 31.350 115.480 ;
        RECT 31.120 115.280 31.260 115.420 ;
        RECT 24.680 115.140 31.260 115.280 ;
        RECT 31.505 115.280 31.795 115.325 ;
        RECT 31.950 115.280 32.270 115.340 ;
        RECT 31.505 115.140 32.270 115.280 ;
        RECT 32.500 115.280 32.640 115.480 ;
        RECT 36.090 115.420 36.410 115.680 ;
        RECT 39.325 115.620 39.615 115.665 ;
        RECT 39.770 115.620 40.090 115.680 ;
        RECT 36.640 115.480 38.160 115.620 ;
        RECT 36.640 115.280 36.780 115.480 ;
        RECT 37.470 115.385 37.760 115.480 ;
        RECT 32.500 115.140 36.780 115.280 ;
        RECT 38.020 115.280 38.160 115.480 ;
        RECT 39.325 115.480 40.090 115.620 ;
        RECT 39.325 115.435 39.615 115.480 ;
        RECT 39.770 115.420 40.090 115.480 ;
        RECT 41.150 115.420 41.470 115.680 ;
        RECT 44.845 115.435 45.135 115.665 ;
        RECT 44.920 115.280 45.060 115.435 ;
        RECT 45.750 115.420 46.070 115.680 ;
        RECT 52.650 115.620 52.970 115.680 ;
        RECT 55.410 115.665 55.730 115.680 ;
        RECT 54.045 115.620 54.335 115.665 ;
        RECT 52.650 115.480 54.335 115.620 ;
        RECT 52.650 115.420 52.970 115.480 ;
        RECT 54.045 115.435 54.335 115.480 ;
        RECT 55.380 115.435 55.730 115.665 ;
        RECT 55.410 115.420 55.730 115.435 ;
        RECT 60.470 115.620 60.790 115.680 ;
        RECT 61.405 115.620 61.695 115.665 ;
        RECT 63.690 115.620 64.010 115.680 ;
        RECT 60.470 115.480 64.010 115.620 ;
        RECT 60.470 115.420 60.790 115.480 ;
        RECT 61.405 115.435 61.695 115.480 ;
        RECT 63.690 115.420 64.010 115.480 ;
        RECT 64.150 115.420 64.470 115.680 ;
        RECT 65.070 115.420 65.390 115.680 ;
        RECT 66.080 115.340 66.220 115.820 ;
        RECT 67.830 115.760 68.150 115.820 ;
        RECT 78.410 115.760 78.730 116.020 ;
        RECT 80.250 115.960 80.570 116.020 ;
        RECT 84.390 115.960 84.710 116.020 ;
        RECT 80.250 115.820 84.710 115.960 ;
        RECT 80.250 115.760 80.570 115.820 ;
        RECT 66.925 115.620 67.215 115.665 ;
        RECT 68.290 115.620 68.610 115.730 ;
        RECT 69.670 115.665 69.990 115.680 ;
        RECT 66.925 115.480 68.610 115.620 ;
        RECT 66.925 115.435 67.215 115.480 ;
        RECT 68.290 115.470 68.610 115.480 ;
        RECT 69.640 115.435 69.990 115.665 ;
        RECT 78.500 115.620 78.640 115.760 ;
        RECT 80.725 115.620 81.015 115.665 ;
        RECT 78.500 115.480 81.015 115.620 ;
        RECT 80.725 115.435 81.015 115.480 ;
        RECT 69.670 115.420 69.990 115.435 ;
        RECT 81.170 115.420 81.490 115.680 ;
        RECT 81.630 115.420 81.950 115.680 ;
        RECT 82.640 115.665 82.780 115.820 ;
        RECT 84.390 115.760 84.710 115.820 ;
        RECT 82.565 115.435 82.855 115.665 ;
        RECT 83.025 115.435 83.315 115.665 ;
        RECT 85.325 115.620 85.615 115.665 ;
        RECT 85.770 115.620 86.090 115.680 ;
        RECT 85.325 115.480 86.090 115.620 ;
        RECT 85.325 115.435 85.615 115.480 ;
        RECT 38.020 115.140 45.060 115.280 ;
        RECT 21.385 115.095 21.675 115.140 ;
        RECT 31.505 115.095 31.795 115.140 ;
        RECT 31.950 115.080 32.270 115.140 ;
        RECT 51.270 115.080 51.590 115.340 ;
        RECT 54.925 115.280 55.215 115.325 ;
        RECT 56.115 115.280 56.405 115.325 ;
        RECT 58.635 115.280 58.925 115.325 ;
        RECT 54.925 115.140 58.925 115.280 ;
        RECT 54.925 115.095 55.215 115.140 ;
        RECT 56.115 115.095 56.405 115.140 ;
        RECT 58.635 115.095 58.925 115.140 ;
        RECT 61.865 115.280 62.155 115.325 ;
        RECT 62.310 115.280 62.630 115.340 ;
        RECT 61.865 115.140 62.630 115.280 ;
        RECT 61.865 115.095 62.155 115.140 ;
        RECT 62.310 115.080 62.630 115.140 ;
        RECT 63.230 115.080 63.550 115.340 ;
        RECT 65.545 115.095 65.835 115.325 ;
        RECT 32.870 114.940 33.190 115.000 ;
        RECT 38.405 114.940 38.695 114.985 ;
        RECT 32.870 114.800 38.695 114.940 ;
        RECT 32.870 114.740 33.190 114.800 ;
        RECT 38.405 114.755 38.695 114.800 ;
        RECT 54.530 114.940 54.820 114.985 ;
        RECT 56.630 114.940 56.920 114.985 ;
        RECT 58.200 114.940 58.490 114.985 ;
        RECT 63.320 114.940 63.460 115.080 ;
        RECT 65.620 114.940 65.760 115.095 ;
        RECT 65.990 115.080 66.310 115.340 ;
        RECT 66.450 115.280 66.770 115.340 ;
        RECT 68.305 115.280 68.595 115.325 ;
        RECT 66.450 115.140 68.595 115.280 ;
        RECT 66.450 115.080 66.770 115.140 ;
        RECT 68.305 115.095 68.595 115.140 ;
        RECT 69.185 115.280 69.475 115.325 ;
        RECT 70.375 115.280 70.665 115.325 ;
        RECT 72.895 115.280 73.185 115.325 ;
        RECT 69.185 115.140 73.185 115.280 ;
        RECT 69.185 115.095 69.475 115.140 ;
        RECT 70.375 115.095 70.665 115.140 ;
        RECT 72.895 115.095 73.185 115.140 ;
        RECT 78.425 115.280 78.715 115.325 ;
        RECT 83.100 115.280 83.240 115.435 ;
        RECT 85.770 115.420 86.090 115.480 ;
        RECT 86.245 115.435 86.535 115.665 ;
        RECT 86.320 115.280 86.460 115.435 ;
        RECT 86.690 115.420 87.010 115.680 ;
        RECT 88.990 115.280 89.310 115.340 ;
        RECT 78.425 115.140 83.240 115.280 ;
        RECT 85.860 115.140 89.310 115.280 ;
        RECT 78.425 115.095 78.715 115.140 ;
        RECT 54.530 114.800 58.490 114.940 ;
        RECT 54.530 114.755 54.820 114.800 ;
        RECT 56.630 114.755 56.920 114.800 ;
        RECT 58.200 114.755 58.490 114.800 ;
        RECT 61.480 114.800 65.760 114.940 ;
        RECT 68.790 114.940 69.080 114.985 ;
        RECT 70.890 114.940 71.180 114.985 ;
        RECT 72.460 114.940 72.750 114.985 ;
        RECT 68.790 114.800 72.750 114.940 ;
        RECT 14.485 114.600 14.775 114.645 ;
        RECT 23.670 114.600 23.990 114.660 ;
        RECT 14.485 114.460 23.990 114.600 ;
        RECT 14.485 114.415 14.775 114.460 ;
        RECT 23.670 114.400 23.990 114.460 ;
        RECT 25.525 114.600 25.815 114.645 ;
        RECT 25.970 114.600 26.290 114.660 ;
        RECT 25.525 114.460 26.290 114.600 ;
        RECT 25.525 114.415 25.815 114.460 ;
        RECT 25.970 114.400 26.290 114.460 ;
        RECT 29.205 114.600 29.495 114.645 ;
        RECT 30.110 114.600 30.430 114.660 ;
        RECT 29.205 114.460 30.430 114.600 ;
        RECT 29.205 114.415 29.495 114.460 ;
        RECT 30.110 114.400 30.430 114.460 ;
        RECT 34.710 114.400 35.030 114.660 ;
        RECT 35.185 114.600 35.475 114.645 ;
        RECT 35.630 114.600 35.950 114.660 ;
        RECT 35.185 114.460 35.950 114.600 ;
        RECT 35.185 114.415 35.475 114.460 ;
        RECT 35.630 114.400 35.950 114.460 ;
        RECT 39.310 114.600 39.630 114.660 ;
        RECT 44.845 114.600 45.135 114.645 ;
        RECT 39.310 114.460 45.135 114.600 ;
        RECT 39.310 114.400 39.630 114.460 ;
        RECT 44.845 114.415 45.135 114.460 ;
        RECT 49.890 114.600 50.210 114.660 ;
        RECT 54.030 114.600 54.350 114.660 ;
        RECT 61.480 114.645 61.620 114.800 ;
        RECT 68.790 114.755 69.080 114.800 ;
        RECT 70.890 114.755 71.180 114.800 ;
        RECT 72.460 114.755 72.750 114.800 ;
        RECT 75.205 114.940 75.495 114.985 ;
        RECT 78.500 114.940 78.640 115.095 ;
        RECT 85.860 115.000 86.000 115.140 ;
        RECT 88.990 115.080 89.310 115.140 ;
        RECT 75.205 114.800 78.640 114.940 ;
        RECT 83.470 114.940 83.790 115.000 ;
        RECT 84.405 114.940 84.695 114.985 ;
        RECT 83.470 114.800 84.695 114.940 ;
        RECT 75.205 114.755 75.495 114.800 ;
        RECT 83.470 114.740 83.790 114.800 ;
        RECT 84.405 114.755 84.695 114.800 ;
        RECT 85.770 114.740 86.090 115.000 ;
        RECT 100.000 114.680 100.830 116.780 ;
        RECT 106.500 116.390 107.750 116.830 ;
        RECT 117.700 116.810 118.560 118.870 ;
        RECT 120.000 116.810 120.770 120.420 ;
        RECT 122.340 119.370 125.190 120.490 ;
        RECT 125.580 120.190 125.930 120.940 ;
        RECT 126.680 120.820 128.550 120.980 ;
        RECT 126.680 120.770 127.440 120.820 ;
        RECT 128.320 120.750 128.550 120.820 ;
        RECT 136.960 120.750 137.190 120.980 ;
        RECT 128.755 120.470 136.755 120.700 ;
        RECT 125.580 120.130 125.870 120.190 ;
        RECT 125.490 120.010 125.870 120.130 ;
        RECT 128.850 120.070 136.710 120.470 ;
        RECT 137.520 120.070 138.480 129.550 ;
        RECT 122.280 119.140 125.280 119.370 ;
        RECT 125.490 119.180 125.830 120.010 ;
        RECT 127.840 120.000 138.480 120.070 ;
        RECT 122.330 119.110 125.190 119.140 ;
        RECT 122.330 119.090 123.500 119.110 ;
        RECT 124.460 119.100 125.190 119.110 ;
        RECT 122.280 118.700 125.280 118.930 ;
        RECT 125.485 118.890 125.830 119.180 ;
        RECT 126.020 118.960 138.480 120.000 ;
        RECT 139.930 131.780 140.700 135.360 ;
        RECT 142.370 134.310 145.220 135.430 ;
        RECT 145.610 135.130 145.960 135.880 ;
        RECT 146.710 135.760 148.580 135.920 ;
        RECT 146.710 135.710 147.470 135.760 ;
        RECT 148.350 135.690 148.580 135.760 ;
        RECT 156.990 135.690 157.220 135.920 ;
        RECT 148.785 135.410 156.785 135.640 ;
        RECT 145.610 135.070 145.900 135.130 ;
        RECT 145.520 134.950 145.900 135.070 ;
        RECT 148.880 135.010 156.740 135.410 ;
        RECT 157.550 135.010 158.510 144.490 ;
        RECT 142.310 134.080 145.310 134.310 ;
        RECT 145.520 134.120 145.860 134.950 ;
        RECT 147.870 134.940 158.510 135.010 ;
        RECT 142.360 134.050 145.220 134.080 ;
        RECT 142.360 134.030 143.530 134.050 ;
        RECT 144.490 134.040 145.220 134.050 ;
        RECT 142.310 133.640 145.310 133.870 ;
        RECT 145.515 133.830 145.860 134.120 ;
        RECT 146.050 133.900 158.510 134.940 ;
        RECT 146.050 133.880 158.500 133.900 ;
        RECT 145.520 133.720 145.860 133.830 ;
        RECT 146.090 133.870 151.760 133.880 ;
        RECT 152.760 133.870 158.500 133.880 ;
        RECT 142.400 133.470 145.260 133.640 ;
        RECT 146.090 133.470 146.520 133.870 ;
        RECT 142.370 133.100 146.520 133.470 ;
        RECT 139.930 129.680 140.790 131.780 ;
        RECT 146.460 131.390 147.710 131.830 ;
        RECT 157.640 131.810 158.500 133.870 ;
        RECT 144.400 131.380 149.640 131.390 ;
        RECT 141.450 131.280 156.750 131.380 ;
        RECT 141.450 131.270 156.785 131.280 ;
        RECT 141.410 131.150 156.785 131.270 ;
        RECT 141.410 131.040 145.410 131.150 ;
        RECT 146.460 131.070 148.200 131.150 ;
        RECT 148.780 131.070 156.785 131.150 ;
        RECT 146.460 130.990 147.710 131.070 ;
        RECT 148.785 131.050 156.785 131.070 ;
        RECT 141.020 130.740 141.250 130.990 ;
        RECT 145.570 130.850 145.800 130.990 ;
        RECT 148.350 130.850 148.580 131.000 ;
        RECT 145.570 130.740 148.580 130.850 ;
        RECT 156.990 130.740 157.220 131.000 ;
        RECT 141.020 130.300 157.220 130.740 ;
        RECT 141.020 130.030 141.250 130.300 ;
        RECT 145.570 130.270 157.220 130.300 ;
        RECT 145.570 130.180 148.580 130.270 ;
        RECT 145.570 130.030 145.800 130.180 ;
        RECT 148.350 130.040 148.580 130.180 ;
        RECT 156.990 130.040 157.220 130.270 ;
        RECT 141.410 129.750 145.410 129.980 ;
        RECT 148.785 129.770 156.785 129.990 ;
        RECT 157.550 129.770 158.510 131.810 ;
        RECT 148.785 129.760 158.510 129.770 ;
        RECT 141.410 129.680 145.400 129.750 ;
        RECT 139.930 129.570 145.400 129.680 ;
        RECT 148.840 129.600 158.510 129.760 ;
        RECT 139.930 129.480 143.090 129.570 ;
        RECT 156.580 129.550 158.510 129.600 ;
        RECT 139.930 126.210 140.790 129.480 ;
        RECT 144.440 129.020 149.690 129.030 ;
        RECT 144.440 128.910 156.750 129.020 ;
        RECT 141.470 128.850 156.750 128.910 ;
        RECT 141.470 128.840 156.785 128.850 ;
        RECT 141.410 128.710 156.785 128.840 ;
        RECT 141.410 128.700 146.570 128.710 ;
        RECT 141.410 128.610 145.410 128.700 ;
        RECT 148.785 128.620 156.785 128.710 ;
        RECT 148.870 128.610 156.760 128.620 ;
        RECT 141.020 128.250 141.250 128.560 ;
        RECT 141.470 128.250 145.370 128.610 ;
        RECT 145.570 128.250 145.800 128.560 ;
        RECT 141.020 126.910 145.800 128.250 ;
        RECT 141.020 126.600 141.250 126.910 ;
        RECT 145.570 126.600 145.800 126.910 ;
        RECT 148.350 128.030 148.580 128.570 ;
        RECT 149.390 128.030 150.400 128.060 ;
        RECT 156.990 128.030 157.220 128.570 ;
        RECT 148.350 127.130 157.220 128.030 ;
        RECT 148.350 126.610 148.580 127.130 ;
        RECT 149.390 127.060 150.400 127.130 ;
        RECT 156.990 126.610 157.220 127.130 ;
        RECT 141.410 126.320 145.410 126.550 ;
        RECT 148.785 126.330 156.785 126.560 ;
        RECT 139.930 126.170 141.090 126.210 ;
        RECT 139.930 126.090 141.330 126.170 ;
        RECT 141.700 126.100 145.360 126.320 ;
        RECT 141.700 126.090 143.140 126.100 ;
        RECT 139.930 126.050 143.140 126.090 ;
        RECT 139.930 125.960 142.650 126.050 ;
        RECT 148.850 126.040 156.740 126.330 ;
        RECT 139.930 125.900 141.980 125.960 ;
        RECT 139.930 125.850 141.730 125.900 ;
        RECT 139.930 122.510 140.790 125.850 ;
        RECT 148.840 125.550 156.760 125.560 ;
        RECT 145.070 125.540 156.760 125.550 ;
        RECT 141.450 125.420 156.760 125.540 ;
        RECT 141.450 125.410 156.785 125.420 ;
        RECT 141.410 125.290 156.785 125.410 ;
        RECT 141.410 125.180 145.410 125.290 ;
        RECT 141.020 124.840 141.250 125.130 ;
        RECT 141.470 124.840 145.360 125.180 ;
        RECT 145.570 124.840 145.800 125.130 ;
        RECT 141.020 123.470 145.800 124.840 ;
        RECT 141.020 123.170 141.250 123.470 ;
        RECT 145.570 123.170 145.800 123.470 ;
        RECT 141.410 122.890 145.410 123.120 ;
        RECT 141.660 122.660 145.230 122.890 ;
        RECT 141.660 122.510 145.350 122.660 ;
        RECT 139.930 122.230 145.350 122.510 ;
        RECT 146.600 122.340 147.220 125.290 ;
        RECT 148.785 125.190 156.785 125.290 ;
        RECT 148.840 125.180 156.760 125.190 ;
        RECT 148.350 124.480 148.580 125.140 ;
        RECT 149.360 124.480 150.360 124.570 ;
        RECT 156.990 124.480 157.220 125.140 ;
        RECT 148.350 123.660 157.220 124.480 ;
        RECT 148.350 123.180 148.580 123.660 ;
        RECT 149.360 123.570 150.360 123.660 ;
        RECT 156.990 123.180 157.220 123.660 ;
        RECT 148.785 122.900 156.785 123.130 ;
        RECT 139.930 121.770 145.360 122.230 ;
        RECT 139.930 120.420 141.960 121.770 ;
        RECT 143.710 121.760 145.360 121.770 ;
        RECT 142.400 120.490 143.400 121.210 ;
        RECT 143.710 120.950 144.020 121.760 ;
        RECT 144.480 121.480 145.360 121.760 ;
        RECT 145.600 121.940 147.220 122.340 ;
        RECT 148.870 121.990 156.740 122.900 ;
        RECT 144.420 121.250 145.420 121.480 ;
        RECT 145.600 121.290 145.950 121.940 ;
        RECT 146.600 121.930 147.220 121.940 ;
        RECT 148.785 121.760 156.785 121.990 ;
        RECT 148.870 121.750 156.740 121.760 ;
        RECT 144.480 121.040 145.360 121.060 ;
        RECT 143.750 120.660 144.020 120.950 ;
        RECT 144.420 120.810 145.420 121.040 ;
        RECT 145.580 121.000 145.950 121.290 ;
        RECT 145.610 120.940 145.950 121.000 ;
        RECT 146.710 121.610 147.470 121.660 ;
        RECT 148.350 121.610 148.580 121.710 ;
        RECT 146.710 121.400 148.580 121.610 ;
        RECT 156.990 121.400 157.220 121.710 ;
        RECT 146.710 120.980 149.250 121.400 ;
        RECT 156.620 120.980 157.220 121.400 ;
        RECT 144.480 120.660 145.360 120.810 ;
        RECT 144.490 120.490 145.220 120.660 ;
        RECT 126.020 118.940 138.460 118.960 ;
        RECT 125.490 118.780 125.830 118.890 ;
        RECT 126.060 118.930 131.730 118.940 ;
        RECT 132.730 118.930 138.460 118.940 ;
        RECT 122.370 118.530 125.230 118.700 ;
        RECT 126.060 118.530 126.490 118.930 ;
        RECT 122.340 118.160 126.490 118.530 ;
        RECT 104.440 116.380 109.680 116.390 ;
        RECT 101.490 116.280 116.790 116.380 ;
        RECT 101.490 116.270 116.825 116.280 ;
        RECT 101.450 116.150 116.825 116.270 ;
        RECT 101.450 116.040 105.450 116.150 ;
        RECT 106.500 116.070 108.240 116.150 ;
        RECT 108.820 116.070 116.825 116.150 ;
        RECT 106.500 115.990 107.750 116.070 ;
        RECT 108.825 116.050 116.825 116.070 ;
        RECT 101.060 115.740 101.290 115.990 ;
        RECT 105.610 115.850 105.840 115.990 ;
        RECT 108.390 115.850 108.620 116.000 ;
        RECT 105.610 115.740 108.620 115.850 ;
        RECT 117.030 115.740 117.260 116.000 ;
        RECT 101.060 115.300 117.260 115.740 ;
        RECT 101.060 115.030 101.290 115.300 ;
        RECT 105.610 115.270 117.260 115.300 ;
        RECT 105.610 115.180 108.620 115.270 ;
        RECT 105.610 115.030 105.840 115.180 ;
        RECT 108.390 115.040 108.620 115.180 ;
        RECT 117.030 115.040 117.260 115.270 ;
        RECT 101.450 114.750 105.450 114.980 ;
        RECT 108.825 114.770 116.825 114.990 ;
        RECT 117.590 114.770 118.560 116.810 ;
        RECT 108.825 114.760 118.560 114.770 ;
        RECT 101.450 114.680 105.440 114.750 ;
        RECT 61.405 114.600 61.695 114.645 ;
        RECT 49.890 114.460 61.695 114.600 ;
        RECT 49.890 114.400 50.210 114.460 ;
        RECT 54.030 114.400 54.350 114.460 ;
        RECT 61.405 114.415 61.695 114.460 ;
        RECT 63.245 114.600 63.535 114.645 ;
        RECT 65.990 114.600 66.310 114.660 ;
        RECT 63.245 114.460 66.310 114.600 ;
        RECT 63.245 114.415 63.535 114.460 ;
        RECT 65.990 114.400 66.310 114.460 ;
        RECT 67.845 114.600 68.135 114.645 ;
        RECT 72.890 114.600 73.210 114.660 ;
        RECT 67.845 114.460 73.210 114.600 ;
        RECT 67.845 114.415 68.135 114.460 ;
        RECT 72.890 114.400 73.210 114.460 ;
        RECT 75.650 114.400 75.970 114.660 ;
        RECT 77.950 114.600 78.270 114.660 ;
        RECT 81.170 114.600 81.490 114.660 ;
        RECT 77.950 114.460 81.490 114.600 ;
        RECT 77.950 114.400 78.270 114.460 ;
        RECT 81.170 114.400 81.490 114.460 ;
        RECT 87.625 114.600 87.915 114.645 ;
        RECT 88.070 114.600 88.390 114.660 ;
        RECT 87.625 114.460 88.390 114.600 ;
        RECT 87.625 114.415 87.915 114.460 ;
        RECT 88.070 114.400 88.390 114.460 ;
        RECT 100.000 114.570 105.440 114.680 ;
        RECT 108.880 114.600 118.560 114.760 ;
        RECT 100.000 114.480 103.130 114.570 ;
        RECT 116.620 114.550 118.560 114.600 ;
        RECT 12.100 113.780 89.840 114.260 ;
        RECT 23.210 113.380 23.530 113.640 ;
        RECT 25.510 113.380 25.830 113.640 ;
        RECT 37.485 113.580 37.775 113.625 ;
        RECT 42.990 113.580 43.310 113.640 ;
        RECT 27.900 113.440 31.720 113.580 ;
        RECT 16.770 113.240 17.090 113.300 ;
        RECT 17.705 113.240 17.995 113.285 ;
        RECT 16.770 113.100 22.060 113.240 ;
        RECT 16.770 113.040 17.090 113.100 ;
        RECT 17.705 113.055 17.995 113.100 ;
        RECT 14.945 112.900 15.235 112.945 ;
        RECT 17.230 112.900 17.550 112.960 ;
        RECT 20.005 112.900 20.295 112.945 ;
        RECT 14.945 112.760 20.295 112.900 ;
        RECT 14.945 112.715 15.235 112.760 ;
        RECT 17.230 112.700 17.550 112.760 ;
        RECT 20.005 112.715 20.295 112.760 ;
        RECT 20.450 112.700 20.770 112.960 ;
        RECT 21.920 112.945 22.060 113.100 ;
        RECT 21.845 112.900 22.135 112.945 ;
        RECT 21.845 112.760 24.360 112.900 ;
        RECT 21.845 112.715 22.135 112.760 ;
        RECT 15.405 112.560 15.695 112.605 ;
        RECT 18.610 112.560 18.930 112.620 ;
        RECT 15.405 112.420 18.930 112.560 ;
        RECT 15.405 112.375 15.695 112.420 ;
        RECT 18.610 112.360 18.930 112.420 ;
        RECT 19.420 112.375 19.710 112.605 ;
        RECT 20.910 112.560 21.230 112.620 ;
        RECT 22.305 112.560 22.595 112.605 ;
        RECT 20.910 112.420 22.595 112.560 ;
        RECT 17.690 112.020 18.010 112.280 ;
        RECT 19.495 112.220 19.635 112.375 ;
        RECT 20.910 112.360 21.230 112.420 ;
        RECT 22.305 112.375 22.595 112.420 ;
        RECT 23.075 112.560 23.365 112.605 ;
        RECT 23.670 112.560 23.990 112.620 ;
        RECT 23.075 112.420 23.990 112.560 ;
        RECT 23.075 112.375 23.365 112.420 ;
        RECT 23.670 112.360 23.990 112.420 ;
        RECT 21.370 112.220 21.690 112.280 ;
        RECT 19.495 112.080 21.690 112.220 ;
        RECT 24.220 112.220 24.360 112.760 ;
        RECT 26.430 112.560 26.720 112.605 ;
        RECT 27.900 112.560 28.040 113.440 ;
        RECT 31.580 113.300 31.720 113.440 ;
        RECT 37.485 113.440 43.310 113.580 ;
        RECT 37.485 113.395 37.775 113.440 ;
        RECT 42.990 113.380 43.310 113.440 ;
        RECT 48.065 113.580 48.355 113.625 ;
        RECT 48.970 113.580 49.290 113.640 ;
        RECT 48.065 113.440 49.290 113.580 ;
        RECT 48.065 113.395 48.355 113.440 ;
        RECT 48.970 113.380 49.290 113.440 ;
        RECT 55.410 113.380 55.730 113.640 ;
        RECT 60.485 113.580 60.775 113.625 ;
        RECT 65.070 113.580 65.390 113.640 ;
        RECT 60.485 113.440 65.390 113.580 ;
        RECT 60.485 113.395 60.775 113.440 ;
        RECT 65.070 113.380 65.390 113.440 ;
        RECT 68.290 113.380 68.610 113.640 ;
        RECT 69.670 113.580 69.990 113.640 ;
        RECT 70.145 113.580 70.435 113.625 ;
        RECT 69.670 113.440 70.435 113.580 ;
        RECT 69.670 113.380 69.990 113.440 ;
        RECT 70.145 113.395 70.435 113.440 ;
        RECT 75.190 113.580 75.510 113.640 ;
        RECT 82.090 113.580 82.410 113.640 ;
        RECT 75.190 113.440 82.410 113.580 ;
        RECT 75.190 113.380 75.510 113.440 ;
        RECT 82.090 113.380 82.410 113.440 ;
        RECT 30.570 113.240 30.890 113.300 ;
        RECT 28.820 113.100 30.890 113.240 ;
        RECT 28.820 112.945 28.960 113.100 ;
        RECT 30.570 113.040 30.890 113.100 ;
        RECT 31.490 113.240 31.810 113.300 ;
        RECT 37.930 113.240 38.250 113.300 ;
        RECT 31.490 113.100 38.250 113.240 ;
        RECT 31.490 113.040 31.810 113.100 ;
        RECT 37.930 113.040 38.250 113.100 ;
        RECT 38.390 113.240 38.710 113.300 ;
        RECT 41.650 113.240 41.940 113.285 ;
        RECT 43.750 113.240 44.040 113.285 ;
        RECT 45.320 113.240 45.610 113.285 ;
        RECT 38.390 113.100 41.380 113.240 ;
        RECT 38.390 113.040 38.710 113.100 ;
        RECT 28.745 112.715 29.035 112.945 ;
        RECT 31.950 112.900 32.270 112.960 ;
        RECT 34.265 112.900 34.555 112.945 ;
        RECT 29.740 112.760 34.555 112.900 ;
        RECT 26.430 112.420 28.040 112.560 ;
        RECT 26.430 112.375 26.720 112.420 ;
        RECT 28.270 112.360 28.590 112.620 ;
        RECT 29.190 112.360 29.510 112.620 ;
        RECT 29.740 112.220 29.880 112.760 ;
        RECT 31.950 112.700 32.270 112.760 ;
        RECT 34.265 112.715 34.555 112.760 ;
        RECT 40.230 112.700 40.550 112.960 ;
        RECT 41.240 112.945 41.380 113.100 ;
        RECT 41.650 113.100 45.610 113.240 ;
        RECT 41.650 113.055 41.940 113.100 ;
        RECT 43.750 113.055 44.040 113.100 ;
        RECT 45.320 113.055 45.610 113.100 ;
        RECT 57.250 113.040 57.570 113.300 ;
        RECT 58.170 113.240 58.490 113.300 ;
        RECT 60.930 113.240 61.250 113.300 ;
        RECT 64.610 113.240 64.930 113.300 ;
        RECT 69.225 113.240 69.515 113.285 ;
        RECT 70.590 113.240 70.910 113.300 ;
        RECT 58.170 113.100 60.240 113.240 ;
        RECT 58.170 113.040 58.490 113.100 ;
        RECT 41.165 112.715 41.455 112.945 ;
        RECT 42.045 112.900 42.335 112.945 ;
        RECT 43.235 112.900 43.525 112.945 ;
        RECT 45.755 112.900 46.045 112.945 ;
        RECT 42.045 112.760 46.045 112.900 ;
        RECT 42.045 112.715 42.335 112.760 ;
        RECT 43.235 112.715 43.525 112.760 ;
        RECT 45.755 112.715 46.045 112.760 ;
        RECT 53.110 112.900 53.430 112.960 ;
        RECT 56.805 112.900 57.095 112.945 ;
        RECT 53.110 112.760 58.860 112.900 ;
        RECT 53.110 112.700 53.430 112.760 ;
        RECT 56.805 112.715 57.095 112.760 ;
        RECT 30.585 112.560 30.875 112.605 ;
        RECT 31.030 112.560 31.350 112.620 ;
        RECT 30.585 112.420 31.350 112.560 ;
        RECT 30.585 112.375 30.875 112.420 ;
        RECT 24.220 112.080 29.880 112.220 ;
        RECT 21.370 112.020 21.690 112.080 ;
        RECT 30.660 111.940 30.800 112.375 ;
        RECT 31.030 112.360 31.350 112.420 ;
        RECT 32.870 112.560 33.190 112.620 ;
        RECT 35.645 112.560 35.935 112.605 ;
        RECT 32.870 112.420 35.935 112.560 ;
        RECT 32.870 112.360 33.190 112.420 ;
        RECT 35.645 112.375 35.935 112.420 ;
        RECT 38.850 112.560 39.170 112.620 ;
        RECT 39.785 112.560 40.075 112.605 ;
        RECT 38.850 112.420 40.075 112.560 ;
        RECT 38.850 112.360 39.170 112.420 ;
        RECT 39.785 112.375 40.075 112.420 ;
        RECT 48.050 112.560 48.370 112.620 ;
        RECT 51.270 112.560 51.590 112.620 ;
        RECT 48.050 112.420 51.590 112.560 ;
        RECT 48.050 112.360 48.370 112.420 ;
        RECT 51.270 112.360 51.590 112.420 ;
        RECT 56.330 112.360 56.650 112.620 ;
        RECT 57.725 112.560 58.015 112.605 ;
        RECT 58.170 112.560 58.490 112.620 ;
        RECT 58.720 112.605 58.860 112.760 ;
        RECT 57.725 112.420 58.490 112.560 ;
        RECT 57.725 112.375 58.015 112.420 ;
        RECT 58.170 112.360 58.490 112.420 ;
        RECT 58.645 112.375 58.935 112.605 ;
        RECT 59.550 112.360 59.870 112.620 ;
        RECT 60.100 112.605 60.240 113.100 ;
        RECT 60.930 113.100 61.620 113.240 ;
        RECT 60.930 113.040 61.250 113.100 ;
        RECT 61.480 112.945 61.620 113.100 ;
        RECT 64.610 113.100 68.980 113.240 ;
        RECT 64.610 113.040 64.930 113.100 ;
        RECT 61.405 112.715 61.695 112.945 ;
        RECT 60.025 112.560 60.315 112.605 ;
        RECT 60.470 112.560 60.790 112.620 ;
        RECT 60.025 112.420 60.790 112.560 ;
        RECT 60.025 112.375 60.315 112.420 ;
        RECT 60.470 112.360 60.790 112.420 ;
        RECT 60.945 112.560 61.235 112.605 ;
        RECT 64.700 112.560 64.840 113.040 ;
        RECT 67.370 112.900 67.690 112.960 ;
        RECT 66.540 112.760 67.690 112.900 ;
        RECT 60.945 112.420 64.840 112.560 ;
        RECT 60.945 112.375 61.235 112.420 ;
        RECT 65.070 112.360 65.390 112.620 ;
        RECT 65.990 112.360 66.310 112.620 ;
        RECT 66.540 112.605 66.680 112.760 ;
        RECT 67.370 112.700 67.690 112.760 ;
        RECT 66.465 112.375 66.755 112.605 ;
        RECT 66.925 112.560 67.215 112.605 ;
        RECT 67.830 112.560 68.150 112.620 ;
        RECT 68.840 112.605 68.980 113.100 ;
        RECT 69.225 113.100 70.910 113.240 ;
        RECT 69.225 113.055 69.515 113.100 ;
        RECT 70.590 113.040 70.910 113.100 ;
        RECT 71.510 113.240 71.830 113.300 ;
        RECT 78.410 113.240 78.730 113.300 ;
        RECT 71.510 113.100 78.730 113.240 ;
        RECT 71.510 113.040 71.830 113.100 ;
        RECT 78.410 113.040 78.730 113.100 ;
        RECT 81.670 113.240 81.960 113.285 ;
        RECT 83.770 113.240 84.060 113.285 ;
        RECT 85.340 113.240 85.630 113.285 ;
        RECT 81.670 113.100 85.630 113.240 ;
        RECT 81.670 113.055 81.960 113.100 ;
        RECT 83.770 113.055 84.060 113.100 ;
        RECT 85.340 113.055 85.630 113.100 ;
        RECT 72.430 112.700 72.750 112.960 ;
        RECT 72.890 112.700 73.210 112.960 ;
        RECT 82.065 112.900 82.355 112.945 ;
        RECT 83.255 112.900 83.545 112.945 ;
        RECT 85.775 112.900 86.065 112.945 ;
        RECT 82.065 112.760 86.065 112.900 ;
        RECT 82.065 112.715 82.355 112.760 ;
        RECT 83.255 112.715 83.545 112.760 ;
        RECT 85.775 112.715 86.065 112.760 ;
        RECT 66.925 112.420 68.150 112.560 ;
        RECT 66.925 112.375 67.215 112.420 ;
        RECT 67.830 112.360 68.150 112.420 ;
        RECT 68.765 112.375 69.055 112.605 ;
        RECT 69.670 112.560 69.990 112.620 ;
        RECT 71.050 112.560 71.370 112.620 ;
        RECT 69.670 112.420 71.370 112.560 ;
        RECT 69.670 112.360 69.990 112.420 ;
        RECT 71.050 112.360 71.370 112.420 ;
        RECT 71.985 112.560 72.275 112.605 ;
        RECT 75.650 112.560 75.970 112.620 ;
        RECT 71.985 112.420 75.970 112.560 ;
        RECT 71.985 112.375 72.275 112.420 ;
        RECT 75.650 112.360 75.970 112.420 ;
        RECT 77.490 112.560 77.810 112.620 ;
        RECT 78.870 112.560 79.190 112.620 ;
        RECT 81.185 112.560 81.475 112.605 ;
        RECT 77.490 112.420 81.475 112.560 ;
        RECT 77.490 112.360 77.810 112.420 ;
        RECT 78.870 112.360 79.190 112.420 ;
        RECT 81.185 112.375 81.475 112.420 ;
        RECT 33.330 112.220 33.650 112.280 ;
        RECT 36.105 112.220 36.395 112.265 ;
        RECT 33.330 112.080 36.395 112.220 ;
        RECT 33.330 112.020 33.650 112.080 ;
        RECT 36.105 112.035 36.395 112.080 ;
        RECT 36.690 112.220 36.980 112.265 ;
        RECT 42.500 112.220 42.790 112.265 ;
        RECT 50.810 112.220 51.130 112.280 ;
        RECT 36.690 112.080 38.160 112.220 ;
        RECT 36.690 112.035 36.980 112.080 ;
        RECT 14.010 111.680 14.330 111.940 ;
        RECT 18.610 111.680 18.930 111.940 ;
        RECT 26.445 111.880 26.735 111.925 ;
        RECT 30.570 111.880 30.890 111.940 ;
        RECT 38.020 111.925 38.160 112.080 ;
        RECT 42.500 112.080 51.130 112.220 ;
        RECT 42.500 112.035 42.790 112.080 ;
        RECT 50.810 112.020 51.130 112.080 ;
        RECT 59.105 112.220 59.395 112.265 ;
        RECT 61.390 112.220 61.710 112.280 ;
        RECT 76.570 112.220 76.890 112.280 ;
        RECT 59.105 112.080 68.980 112.220 ;
        RECT 59.105 112.035 59.395 112.080 ;
        RECT 61.390 112.020 61.710 112.080 ;
        RECT 68.840 111.940 68.980 112.080 ;
        RECT 76.570 112.080 78.180 112.220 ;
        RECT 76.570 112.020 76.890 112.080 ;
        RECT 26.445 111.740 30.890 111.880 ;
        RECT 26.445 111.695 26.735 111.740 ;
        RECT 30.570 111.680 30.890 111.740 ;
        RECT 37.945 111.695 38.235 111.925 ;
        RECT 61.850 111.880 62.170 111.940 ;
        RECT 64.625 111.880 64.915 111.925 ;
        RECT 61.850 111.740 64.915 111.880 ;
        RECT 61.850 111.680 62.170 111.740 ;
        RECT 64.625 111.695 64.915 111.740 ;
        RECT 68.750 111.680 69.070 111.940 ;
        RECT 71.050 111.880 71.370 111.940 ;
        RECT 77.505 111.880 77.795 111.925 ;
        RECT 71.050 111.740 77.795 111.880 ;
        RECT 78.040 111.880 78.180 112.080 ;
        RECT 78.410 112.020 78.730 112.280 ;
        RECT 79.345 112.035 79.635 112.265 ;
        RECT 81.630 112.220 81.950 112.280 ;
        RECT 82.410 112.220 82.700 112.265 ;
        RECT 81.630 112.080 82.700 112.220 ;
        RECT 79.420 111.880 79.560 112.035 ;
        RECT 81.630 112.020 81.950 112.080 ;
        RECT 82.410 112.035 82.700 112.080 ;
        RECT 78.040 111.740 79.560 111.880 ;
        RECT 86.230 111.880 86.550 111.940 ;
        RECT 88.085 111.880 88.375 111.925 ;
        RECT 86.230 111.740 88.375 111.880 ;
        RECT 71.050 111.680 71.370 111.740 ;
        RECT 77.505 111.695 77.795 111.740 ;
        RECT 86.230 111.680 86.550 111.740 ;
        RECT 88.085 111.695 88.375 111.740 ;
        RECT 12.100 111.060 89.840 111.540 ;
        RECT 100.000 111.210 100.830 114.480 ;
        RECT 104.480 114.020 109.730 114.030 ;
        RECT 104.480 113.910 116.790 114.020 ;
        RECT 101.510 113.850 116.790 113.910 ;
        RECT 101.510 113.840 116.825 113.850 ;
        RECT 101.450 113.710 116.825 113.840 ;
        RECT 101.450 113.700 106.610 113.710 ;
        RECT 101.450 113.610 105.450 113.700 ;
        RECT 108.825 113.620 116.825 113.710 ;
        RECT 108.910 113.610 116.800 113.620 ;
        RECT 101.060 113.250 101.290 113.560 ;
        RECT 101.510 113.250 105.410 113.610 ;
        RECT 105.610 113.250 105.840 113.560 ;
        RECT 101.060 111.910 105.840 113.250 ;
        RECT 101.060 111.600 101.290 111.910 ;
        RECT 105.610 111.600 105.840 111.910 ;
        RECT 108.390 113.030 108.620 113.570 ;
        RECT 109.430 113.030 110.440 113.060 ;
        RECT 117.030 113.030 117.260 113.570 ;
        RECT 108.390 112.130 117.260 113.030 ;
        RECT 108.390 111.610 108.620 112.130 ;
        RECT 109.430 112.060 110.440 112.130 ;
        RECT 117.030 111.610 117.260 112.130 ;
        RECT 101.450 111.320 105.450 111.550 ;
        RECT 108.825 111.330 116.825 111.560 ;
        RECT 100.000 111.170 101.130 111.210 ;
        RECT 100.000 111.090 101.370 111.170 ;
        RECT 101.740 111.100 105.400 111.320 ;
        RECT 101.740 111.090 103.180 111.100 ;
        RECT 100.000 111.050 103.180 111.090 ;
        RECT 100.000 110.960 102.690 111.050 ;
        RECT 108.890 111.040 116.780 111.330 ;
        RECT 20.925 110.860 21.215 110.905 ;
        RECT 22.290 110.860 22.610 110.920 ;
        RECT 20.925 110.720 22.610 110.860 ;
        RECT 20.925 110.675 21.215 110.720 ;
        RECT 22.290 110.660 22.610 110.720 ;
        RECT 28.270 110.860 28.590 110.920 ;
        RECT 28.745 110.860 29.035 110.905 ;
        RECT 28.270 110.720 29.035 110.860 ;
        RECT 28.270 110.660 28.590 110.720 ;
        RECT 28.745 110.675 29.035 110.720 ;
        RECT 30.120 110.860 30.410 110.905 ;
        RECT 36.560 110.860 36.850 110.905 ;
        RECT 30.120 110.720 36.850 110.860 ;
        RECT 30.120 110.675 30.410 110.720 ;
        RECT 36.560 110.675 36.850 110.720 ;
        RECT 38.405 110.860 38.695 110.905 ;
        RECT 38.850 110.860 39.170 110.920 ;
        RECT 38.405 110.720 39.170 110.860 ;
        RECT 38.405 110.675 38.695 110.720 ;
        RECT 38.850 110.660 39.170 110.720 ;
        RECT 50.810 110.660 51.130 110.920 ;
        RECT 58.170 110.860 58.490 110.920 ;
        RECT 59.565 110.860 59.855 110.905 ;
        RECT 58.170 110.720 59.855 110.860 ;
        RECT 58.170 110.660 58.490 110.720 ;
        RECT 59.565 110.675 59.855 110.720 ;
        RECT 62.770 110.860 63.090 110.920 ;
        RECT 64.625 110.860 64.915 110.905 ;
        RECT 78.410 110.860 78.730 110.920 ;
        RECT 80.710 110.860 81.030 110.920 ;
        RECT 62.770 110.720 64.915 110.860 ;
        RECT 62.770 110.660 63.090 110.720 ;
        RECT 64.625 110.675 64.915 110.720 ;
        RECT 70.680 110.720 75.880 110.860 ;
        RECT 15.360 110.520 15.650 110.565 ;
        RECT 18.610 110.520 18.930 110.580 ;
        RECT 15.360 110.380 18.930 110.520 ;
        RECT 15.360 110.335 15.650 110.380 ;
        RECT 18.610 110.320 18.930 110.380 ;
        RECT 26.430 110.520 26.750 110.580 ;
        RECT 42.990 110.520 43.310 110.580 ;
        RECT 43.970 110.520 44.260 110.565 ;
        RECT 26.430 110.380 28.040 110.520 ;
        RECT 26.430 110.320 26.750 110.380 ;
        RECT 20.910 110.180 21.230 110.240 ;
        RECT 22.290 110.180 22.610 110.240 ;
        RECT 23.225 110.180 23.515 110.225 ;
        RECT 20.910 110.040 22.060 110.180 ;
        RECT 20.910 109.980 21.230 110.040 ;
        RECT 13.550 109.840 13.870 109.900 ;
        RECT 14.025 109.840 14.315 109.885 ;
        RECT 13.550 109.700 14.315 109.840 ;
        RECT 13.550 109.640 13.870 109.700 ;
        RECT 14.025 109.655 14.315 109.700 ;
        RECT 14.905 109.840 15.195 109.885 ;
        RECT 16.095 109.840 16.385 109.885 ;
        RECT 18.615 109.840 18.905 109.885 ;
        RECT 14.905 109.700 18.905 109.840 ;
        RECT 14.905 109.655 15.195 109.700 ;
        RECT 16.095 109.655 16.385 109.700 ;
        RECT 18.615 109.655 18.905 109.700 ;
        RECT 21.370 109.640 21.690 109.900 ;
        RECT 21.920 109.840 22.060 110.040 ;
        RECT 22.290 110.040 23.515 110.180 ;
        RECT 22.290 109.980 22.610 110.040 ;
        RECT 23.225 109.995 23.515 110.040 ;
        RECT 24.590 110.180 24.910 110.240 ;
        RECT 25.525 110.180 25.815 110.225 ;
        RECT 24.590 110.040 25.815 110.180 ;
        RECT 24.590 109.980 24.910 110.040 ;
        RECT 25.525 109.995 25.815 110.040 ;
        RECT 27.350 109.980 27.670 110.240 ;
        RECT 27.900 110.225 28.040 110.380 ;
        RECT 42.990 110.380 44.260 110.520 ;
        RECT 42.990 110.320 43.310 110.380 ;
        RECT 43.970 110.335 44.260 110.380 ;
        RECT 56.330 110.520 56.650 110.580 ;
        RECT 59.090 110.520 59.410 110.580 ;
        RECT 63.230 110.520 63.550 110.580 ;
        RECT 67.370 110.520 67.690 110.580 ;
        RECT 56.330 110.380 62.540 110.520 ;
        RECT 56.330 110.320 56.650 110.380 ;
        RECT 59.090 110.320 59.410 110.380 ;
        RECT 27.825 109.995 28.115 110.225 ;
        RECT 29.650 110.180 29.970 110.240 ;
        RECT 31.505 110.180 31.795 110.225 ;
        RECT 34.725 110.180 35.015 110.225 ;
        RECT 29.650 110.040 31.795 110.180 ;
        RECT 29.650 109.980 29.970 110.040 ;
        RECT 31.505 109.995 31.795 110.040 ;
        RECT 31.995 110.040 35.015 110.180 ;
        RECT 22.765 109.840 23.055 109.885 ;
        RECT 21.920 109.700 23.055 109.840 ;
        RECT 22.765 109.655 23.055 109.700 ;
        RECT 26.890 109.840 27.210 109.900 ;
        RECT 31.995 109.840 32.135 110.040 ;
        RECT 34.725 109.995 35.015 110.040 ;
        RECT 48.970 110.180 49.290 110.240 ;
        RECT 49.905 110.180 50.195 110.225 ;
        RECT 48.970 110.040 50.195 110.180 ;
        RECT 48.970 109.980 49.290 110.040 ;
        RECT 49.905 109.995 50.195 110.040 ;
        RECT 58.630 110.180 58.950 110.240 ;
        RECT 58.630 110.040 61.620 110.180 ;
        RECT 58.630 109.980 58.950 110.040 ;
        RECT 26.890 109.700 32.135 109.840 ;
        RECT 26.890 109.640 27.210 109.700 ;
        RECT 32.870 109.640 33.190 109.900 ;
        RECT 34.265 109.840 34.555 109.885 ;
        RECT 37.010 109.840 37.330 109.900 ;
        RECT 33.500 109.700 37.330 109.840 ;
        RECT 14.510 109.500 14.800 109.545 ;
        RECT 16.610 109.500 16.900 109.545 ;
        RECT 18.180 109.500 18.470 109.545 ;
        RECT 14.510 109.360 18.470 109.500 ;
        RECT 14.510 109.315 14.800 109.360 ;
        RECT 16.610 109.315 16.900 109.360 ;
        RECT 18.180 109.315 18.470 109.360 ;
        RECT 31.030 109.500 31.350 109.560 ;
        RECT 33.500 109.500 33.640 109.700 ;
        RECT 34.265 109.655 34.555 109.700 ;
        RECT 37.010 109.640 37.330 109.700 ;
        RECT 40.715 109.840 41.005 109.885 ;
        RECT 43.235 109.840 43.525 109.885 ;
        RECT 44.425 109.840 44.715 109.885 ;
        RECT 40.715 109.700 44.715 109.840 ;
        RECT 40.715 109.655 41.005 109.700 ;
        RECT 43.235 109.655 43.525 109.700 ;
        RECT 44.425 109.655 44.715 109.700 ;
        RECT 45.305 109.840 45.595 109.885 ;
        RECT 48.050 109.840 48.370 109.900 ;
        RECT 45.305 109.700 48.370 109.840 ;
        RECT 45.305 109.655 45.595 109.700 ;
        RECT 48.050 109.640 48.370 109.700 ;
        RECT 48.510 109.840 48.830 109.900 ;
        RECT 53.585 109.840 53.875 109.885 ;
        RECT 48.510 109.700 53.875 109.840 ;
        RECT 48.510 109.640 48.830 109.700 ;
        RECT 53.585 109.655 53.875 109.700 ;
        RECT 60.485 109.655 60.775 109.885 ;
        RECT 31.030 109.360 33.640 109.500 ;
        RECT 33.805 109.500 34.095 109.545 ;
        RECT 39.770 109.500 40.090 109.560 ;
        RECT 33.805 109.360 40.090 109.500 ;
        RECT 31.030 109.300 31.350 109.360 ;
        RECT 33.805 109.315 34.095 109.360 ;
        RECT 39.770 109.300 40.090 109.360 ;
        RECT 41.150 109.500 41.440 109.545 ;
        RECT 42.720 109.500 43.010 109.545 ;
        RECT 44.820 109.500 45.110 109.545 ;
        RECT 41.150 109.360 45.110 109.500 ;
        RECT 60.560 109.500 60.700 109.655 ;
        RECT 60.930 109.640 61.250 109.900 ;
        RECT 61.480 109.885 61.620 110.040 ;
        RECT 61.850 109.980 62.170 110.240 ;
        RECT 62.400 110.180 62.540 110.380 ;
        RECT 63.230 110.380 67.690 110.520 ;
        RECT 63.230 110.320 63.550 110.380 ;
        RECT 67.370 110.320 67.690 110.380 ;
        RECT 64.165 110.180 64.455 110.225 ;
        RECT 62.400 110.040 64.455 110.180 ;
        RECT 64.165 109.995 64.455 110.040 ;
        RECT 70.145 110.180 70.435 110.225 ;
        RECT 70.680 110.180 70.820 110.720 ;
        RECT 72.430 110.520 72.750 110.580 ;
        RECT 71.600 110.380 72.750 110.520 ;
        RECT 70.145 110.040 70.820 110.180 ;
        RECT 70.145 109.995 70.435 110.040 ;
        RECT 71.050 109.980 71.370 110.240 ;
        RECT 71.600 110.225 71.740 110.380 ;
        RECT 72.430 110.320 72.750 110.380 ;
        RECT 73.365 110.520 73.655 110.565 ;
        RECT 75.050 110.520 75.340 110.565 ;
        RECT 73.365 110.380 75.340 110.520 ;
        RECT 75.740 110.520 75.880 110.720 ;
        RECT 78.410 110.720 81.030 110.860 ;
        RECT 78.410 110.660 78.730 110.720 ;
        RECT 80.710 110.660 81.030 110.720 ;
        RECT 81.185 110.860 81.475 110.905 ;
        RECT 81.630 110.860 81.950 110.920 ;
        RECT 81.185 110.720 81.950 110.860 ;
        RECT 81.185 110.675 81.475 110.720 ;
        RECT 81.630 110.660 81.950 110.720 ;
        RECT 82.090 110.860 82.410 110.920 ;
        RECT 84.865 110.860 85.155 110.905 ;
        RECT 82.090 110.720 85.155 110.860 ;
        RECT 82.090 110.660 82.410 110.720 ;
        RECT 84.865 110.675 85.155 110.720 ;
        RECT 100.000 110.900 102.020 110.960 ;
        RECT 100.000 110.850 101.770 110.900 ;
        RECT 79.790 110.520 80.110 110.580 ;
        RECT 75.740 110.380 80.110 110.520 ;
        RECT 73.365 110.335 73.655 110.380 ;
        RECT 75.050 110.335 75.340 110.380 ;
        RECT 79.790 110.320 80.110 110.380 ;
        RECT 80.250 110.520 80.570 110.580 ;
        RECT 80.250 110.380 86.000 110.520 ;
        RECT 80.250 110.320 80.570 110.380 ;
        RECT 71.525 109.995 71.815 110.225 ;
        RECT 71.985 110.180 72.275 110.225 ;
        RECT 82.565 110.180 82.855 110.225 ;
        RECT 71.985 110.040 82.855 110.180 ;
        RECT 71.985 109.995 72.275 110.040 ;
        RECT 82.565 109.995 82.855 110.040 ;
        RECT 83.025 109.995 83.315 110.225 ;
        RECT 61.405 109.840 61.695 109.885 ;
        RECT 67.370 109.840 67.690 109.900 ;
        RECT 72.060 109.840 72.200 109.995 ;
        RECT 61.405 109.700 62.080 109.840 ;
        RECT 61.405 109.655 61.695 109.700 ;
        RECT 61.940 109.560 62.080 109.700 ;
        RECT 67.370 109.700 72.200 109.840 ;
        RECT 67.370 109.640 67.690 109.700 ;
        RECT 73.825 109.655 74.115 109.885 ;
        RECT 74.705 109.840 74.995 109.885 ;
        RECT 75.895 109.840 76.185 109.885 ;
        RECT 78.415 109.840 78.705 109.885 ;
        RECT 74.705 109.700 78.705 109.840 ;
        RECT 83.100 109.840 83.240 109.995 ;
        RECT 83.470 109.980 83.790 110.240 ;
        RECT 84.390 109.980 84.710 110.240 ;
        RECT 85.860 110.225 86.000 110.380 ;
        RECT 85.785 109.995 86.075 110.225 ;
        RECT 86.245 110.180 86.535 110.225 ;
        RECT 86.690 110.180 87.010 110.240 ;
        RECT 86.245 110.040 87.010 110.180 ;
        RECT 86.245 109.995 86.535 110.040 ;
        RECT 83.930 109.840 84.250 109.900 ;
        RECT 83.100 109.700 84.250 109.840 ;
        RECT 74.705 109.655 74.995 109.700 ;
        RECT 75.895 109.655 76.185 109.700 ;
        RECT 78.415 109.655 78.705 109.700 ;
        RECT 60.560 109.360 61.620 109.500 ;
        RECT 41.150 109.315 41.440 109.360 ;
        RECT 42.720 109.315 43.010 109.360 ;
        RECT 44.820 109.315 45.110 109.360 ;
        RECT 61.480 109.220 61.620 109.360 ;
        RECT 61.850 109.300 62.170 109.560 ;
        RECT 25.970 108.960 26.290 109.220 ;
        RECT 46.210 109.160 46.530 109.220 ;
        RECT 47.145 109.160 47.435 109.205 ;
        RECT 46.210 109.020 47.435 109.160 ;
        RECT 46.210 108.960 46.530 109.020 ;
        RECT 47.145 108.975 47.435 109.020 ;
        RECT 61.390 108.960 61.710 109.220 ;
        RECT 73.900 109.160 74.040 109.655 ;
        RECT 83.930 109.640 84.250 109.700 ;
        RECT 74.310 109.500 74.600 109.545 ;
        RECT 76.410 109.500 76.700 109.545 ;
        RECT 77.980 109.500 78.270 109.545 ;
        RECT 74.310 109.360 78.270 109.500 ;
        RECT 74.310 109.315 74.600 109.360 ;
        RECT 76.410 109.315 76.700 109.360 ;
        RECT 77.980 109.315 78.270 109.360 ;
        RECT 83.470 109.500 83.790 109.560 ;
        RECT 85.860 109.500 86.000 109.995 ;
        RECT 86.690 109.980 87.010 110.040 ;
        RECT 87.150 109.980 87.470 110.240 ;
        RECT 87.625 110.180 87.915 110.225 ;
        RECT 87.625 110.040 88.300 110.180 ;
        RECT 87.625 109.995 87.915 110.040 ;
        RECT 88.160 109.900 88.300 110.040 ;
        RECT 88.070 109.640 88.390 109.900 ;
        RECT 83.470 109.360 86.000 109.500 ;
        RECT 83.470 109.300 83.790 109.360 ;
        RECT 77.490 109.160 77.810 109.220 ;
        RECT 73.900 109.020 77.810 109.160 ;
        RECT 77.490 108.960 77.810 109.020 ;
        RECT 12.100 108.340 89.840 108.820 ;
        RECT 13.550 108.140 13.870 108.200 ;
        RECT 13.550 108.000 24.360 108.140 ;
        RECT 13.550 107.940 13.870 108.000 ;
        RECT 14.050 107.800 14.340 107.845 ;
        RECT 16.150 107.800 16.440 107.845 ;
        RECT 17.720 107.800 18.010 107.845 ;
        RECT 14.050 107.660 18.010 107.800 ;
        RECT 14.050 107.615 14.340 107.660 ;
        RECT 16.150 107.615 16.440 107.660 ;
        RECT 17.720 107.615 18.010 107.660 ;
        RECT 20.465 107.800 20.755 107.845 ;
        RECT 20.910 107.800 21.230 107.860 ;
        RECT 20.465 107.660 21.230 107.800 ;
        RECT 24.220 107.800 24.360 108.000 ;
        RECT 24.590 107.940 24.910 108.200 ;
        RECT 27.350 107.940 27.670 108.200 ;
        RECT 28.270 107.940 28.590 108.200 ;
        RECT 29.190 108.140 29.510 108.200 ;
        RECT 30.570 108.140 30.890 108.200 ;
        RECT 29.190 108.000 30.890 108.140 ;
        RECT 29.190 107.940 29.510 108.000 ;
        RECT 30.570 107.940 30.890 108.000 ;
        RECT 37.930 108.140 38.250 108.200 ;
        RECT 40.245 108.140 40.535 108.185 ;
        RECT 37.930 108.000 40.535 108.140 ;
        RECT 37.930 107.940 38.250 108.000 ;
        RECT 40.245 107.955 40.535 108.000 ;
        RECT 47.590 108.140 47.910 108.200 ;
        RECT 48.985 108.140 49.275 108.185 ;
        RECT 47.590 108.000 49.275 108.140 ;
        RECT 47.590 107.940 47.910 108.000 ;
        RECT 48.985 107.955 49.275 108.000 ;
        RECT 60.470 107.940 60.790 108.200 ;
        RECT 64.150 108.140 64.470 108.200 ;
        RECT 68.290 108.140 68.610 108.200 ;
        RECT 80.250 108.140 80.570 108.200 ;
        RECT 83.945 108.140 84.235 108.185 ;
        RECT 62.400 108.000 64.470 108.140 ;
        RECT 33.830 107.800 34.120 107.845 ;
        RECT 35.930 107.800 36.220 107.845 ;
        RECT 37.500 107.800 37.790 107.845 ;
        RECT 50.350 107.800 50.670 107.860 ;
        RECT 24.220 107.660 33.100 107.800 ;
        RECT 20.465 107.615 20.755 107.660 ;
        RECT 20.910 107.600 21.230 107.660 ;
        RECT 13.550 107.260 13.870 107.520 ;
        RECT 14.445 107.460 14.735 107.505 ;
        RECT 15.635 107.460 15.925 107.505 ;
        RECT 18.155 107.460 18.445 107.505 ;
        RECT 14.445 107.320 18.445 107.460 ;
        RECT 21.000 107.460 21.140 107.600 ;
        RECT 22.305 107.460 22.595 107.505 ;
        RECT 30.110 107.460 30.430 107.520 ;
        RECT 21.000 107.320 22.595 107.460 ;
        RECT 14.445 107.275 14.735 107.320 ;
        RECT 15.635 107.275 15.925 107.320 ;
        RECT 18.155 107.275 18.445 107.320 ;
        RECT 22.305 107.275 22.595 107.320 ;
        RECT 23.760 107.320 30.430 107.460 ;
        RECT 14.010 107.120 14.330 107.180 ;
        RECT 23.760 107.165 23.900 107.320 ;
        RECT 30.110 107.260 30.430 107.320 ;
        RECT 31.505 107.460 31.795 107.505 ;
        RECT 32.410 107.460 32.730 107.520 ;
        RECT 31.505 107.320 32.730 107.460 ;
        RECT 31.505 107.275 31.795 107.320 ;
        RECT 32.410 107.260 32.730 107.320 ;
        RECT 14.845 107.120 15.135 107.165 ;
        RECT 14.010 106.980 15.135 107.120 ;
        RECT 14.010 106.920 14.330 106.980 ;
        RECT 14.845 106.935 15.135 106.980 ;
        RECT 22.765 106.935 23.055 107.165 ;
        RECT 23.685 106.935 23.975 107.165 ;
        RECT 27.810 107.120 28.130 107.180 ;
        RECT 28.285 107.120 28.575 107.165 ;
        RECT 27.810 106.980 28.575 107.120 ;
        RECT 22.840 106.780 22.980 106.935 ;
        RECT 27.810 106.920 28.130 106.980 ;
        RECT 28.285 106.935 28.575 106.980 ;
        RECT 28.730 106.920 29.050 107.180 ;
        RECT 31.030 106.920 31.350 107.180 ;
        RECT 32.960 107.120 33.100 107.660 ;
        RECT 33.830 107.660 37.790 107.800 ;
        RECT 33.830 107.615 34.120 107.660 ;
        RECT 35.930 107.615 36.220 107.660 ;
        RECT 37.500 107.615 37.790 107.660 ;
        RECT 49.060 107.660 50.670 107.800 ;
        RECT 34.225 107.460 34.515 107.505 ;
        RECT 35.415 107.460 35.705 107.505 ;
        RECT 37.935 107.460 38.225 107.505 ;
        RECT 34.225 107.320 38.225 107.460 ;
        RECT 34.225 107.275 34.515 107.320 ;
        RECT 35.415 107.275 35.705 107.320 ;
        RECT 37.935 107.275 38.225 107.320 ;
        RECT 47.605 107.460 47.895 107.505 ;
        RECT 48.510 107.460 48.830 107.520 ;
        RECT 49.060 107.505 49.200 107.660 ;
        RECT 50.350 107.600 50.670 107.660 ;
        RECT 51.745 107.800 52.035 107.845 ;
        RECT 53.110 107.800 53.430 107.860 ;
        RECT 51.745 107.660 53.430 107.800 ;
        RECT 60.560 107.800 60.700 107.940 ;
        RECT 62.400 107.800 62.540 108.000 ;
        RECT 64.150 107.940 64.470 108.000 ;
        RECT 64.700 108.000 68.610 108.140 ;
        RECT 60.560 107.660 62.540 107.800 ;
        RECT 51.745 107.615 52.035 107.660 ;
        RECT 47.605 107.320 48.830 107.460 ;
        RECT 47.605 107.275 47.895 107.320 ;
        RECT 48.510 107.260 48.830 107.320 ;
        RECT 48.985 107.275 49.275 107.505 ;
        RECT 49.445 107.460 49.735 107.505 ;
        RECT 51.820 107.460 51.960 107.615 ;
        RECT 53.110 107.600 53.430 107.660 ;
        RECT 49.445 107.320 51.960 107.460 ;
        RECT 52.665 107.460 52.955 107.505 ;
        RECT 53.570 107.460 53.890 107.520 ;
        RECT 62.400 107.505 62.540 107.660 ;
        RECT 52.665 107.320 53.890 107.460 ;
        RECT 49.445 107.275 49.735 107.320 ;
        RECT 52.665 107.275 52.955 107.320 ;
        RECT 53.570 107.260 53.890 107.320 ;
        RECT 62.325 107.275 62.615 107.505 ;
        RECT 62.770 107.460 63.090 107.520 ;
        RECT 64.165 107.460 64.455 107.505 ;
        RECT 64.700 107.460 64.840 108.000 ;
        RECT 68.290 107.940 68.610 108.000 ;
        RECT 76.660 108.000 84.235 108.140 ;
        RECT 65.085 107.615 65.375 107.845 ;
        RECT 67.830 107.800 68.150 107.860 ;
        RECT 71.050 107.800 71.370 107.860 ;
        RECT 71.970 107.800 72.290 107.860 ;
        RECT 67.830 107.660 72.290 107.800 ;
        RECT 62.770 107.320 64.840 107.460 ;
        RECT 62.770 107.260 63.090 107.320 ;
        RECT 64.165 107.275 64.455 107.320 ;
        RECT 33.345 107.120 33.635 107.165 ;
        RECT 33.790 107.120 34.110 107.180 ;
        RECT 34.710 107.165 35.030 107.180 ;
        RECT 34.680 107.120 35.030 107.165 ;
        RECT 32.960 106.980 34.110 107.120 ;
        RECT 34.515 106.980 35.030 107.120 ;
        RECT 33.345 106.935 33.635 106.980 ;
        RECT 33.790 106.920 34.110 106.980 ;
        RECT 34.680 106.935 35.030 106.980 ;
        RECT 44.385 106.935 44.675 107.165 ;
        RECT 45.305 106.935 45.595 107.165 ;
        RECT 34.710 106.920 35.030 106.935 ;
        RECT 27.350 106.780 27.670 106.840 ;
        RECT 22.840 106.640 27.670 106.780 ;
        RECT 27.350 106.580 27.670 106.640 ;
        RECT 29.665 106.780 29.955 106.825 ;
        RECT 35.630 106.780 35.950 106.840 ;
        RECT 29.665 106.640 35.950 106.780 ;
        RECT 29.665 106.595 29.955 106.640 ;
        RECT 35.630 106.580 35.950 106.640 ;
        RECT 23.670 106.440 23.990 106.500 ;
        RECT 28.270 106.440 28.590 106.500 ;
        RECT 23.670 106.300 28.590 106.440 ;
        RECT 23.670 106.240 23.990 106.300 ;
        RECT 28.270 106.240 28.590 106.300 ;
        RECT 32.885 106.440 33.175 106.485 ;
        RECT 36.090 106.440 36.410 106.500 ;
        RECT 32.885 106.300 36.410 106.440 ;
        RECT 44.460 106.440 44.600 106.935 ;
        RECT 45.380 106.780 45.520 106.935 ;
        RECT 45.750 106.920 46.070 107.180 ;
        RECT 46.210 106.920 46.530 107.180 ;
        RECT 49.890 106.920 50.210 107.180 ;
        RECT 51.270 106.920 51.590 107.180 ;
        RECT 54.965 107.120 55.255 107.165 ;
        RECT 52.740 106.980 55.255 107.120 ;
        RECT 52.740 106.840 52.880 106.980 ;
        RECT 54.965 106.935 55.255 106.980 ;
        RECT 55.425 107.120 55.715 107.165 ;
        RECT 55.870 107.120 56.190 107.180 ;
        RECT 55.425 106.980 56.190 107.120 ;
        RECT 55.425 106.935 55.715 106.980 ;
        RECT 55.870 106.920 56.190 106.980 ;
        RECT 56.345 106.935 56.635 107.165 ;
        RECT 47.130 106.780 47.450 106.840 ;
        RECT 45.380 106.640 47.450 106.780 ;
        RECT 47.130 106.580 47.450 106.640 ;
        RECT 48.065 106.780 48.355 106.825 ;
        RECT 50.810 106.780 51.130 106.840 ;
        RECT 48.065 106.640 51.130 106.780 ;
        RECT 48.065 106.595 48.355 106.640 ;
        RECT 50.810 106.580 51.130 106.640 ;
        RECT 52.650 106.580 52.970 106.840 ;
        RECT 56.420 106.780 56.560 106.935 ;
        RECT 56.790 106.920 57.110 107.180 ;
        RECT 60.470 107.120 60.790 107.180 ;
        RECT 61.850 107.120 62.170 107.180 ;
        RECT 60.470 106.980 62.170 107.120 ;
        RECT 60.470 106.920 60.790 106.980 ;
        RECT 61.850 106.920 62.170 106.980 ;
        RECT 63.690 106.920 64.010 107.180 ;
        RECT 65.160 107.120 65.300 107.615 ;
        RECT 67.830 107.600 68.150 107.660 ;
        RECT 71.050 107.600 71.370 107.660 ;
        RECT 71.970 107.600 72.290 107.660 ;
        RECT 65.545 107.120 65.835 107.165 ;
        RECT 65.160 106.980 65.835 107.120 ;
        RECT 65.545 106.935 65.835 106.980 ;
        RECT 67.845 106.935 68.135 107.165 ;
        RECT 76.125 107.120 76.415 107.165 ;
        RECT 76.660 107.120 76.800 108.000 ;
        RECT 80.250 107.940 80.570 108.000 ;
        RECT 83.945 107.955 84.235 108.000 ;
        RECT 87.150 108.140 87.470 108.200 ;
        RECT 87.625 108.140 87.915 108.185 ;
        RECT 87.150 108.000 87.915 108.140 ;
        RECT 87.150 107.940 87.470 108.000 ;
        RECT 87.625 107.955 87.915 108.000 ;
        RECT 77.530 107.800 77.820 107.845 ;
        RECT 79.630 107.800 79.920 107.845 ;
        RECT 81.200 107.800 81.490 107.845 ;
        RECT 77.530 107.660 81.490 107.800 ;
        RECT 77.530 107.615 77.820 107.660 ;
        RECT 79.630 107.615 79.920 107.660 ;
        RECT 81.200 107.615 81.490 107.660 ;
        RECT 77.925 107.460 78.215 107.505 ;
        RECT 79.115 107.460 79.405 107.505 ;
        RECT 81.635 107.460 81.925 107.505 ;
        RECT 88.070 107.460 88.390 107.520 ;
        RECT 77.925 107.320 81.925 107.460 ;
        RECT 77.925 107.275 78.215 107.320 ;
        RECT 79.115 107.275 79.405 107.320 ;
        RECT 81.635 107.275 81.925 107.320 ;
        RECT 82.180 107.320 88.390 107.460 ;
        RECT 76.125 106.980 76.800 107.120 ;
        RECT 77.045 107.120 77.335 107.165 ;
        RECT 77.490 107.120 77.810 107.180 ;
        RECT 82.180 107.120 82.320 107.320 ;
        RECT 88.070 107.260 88.390 107.320 ;
        RECT 100.000 107.510 100.830 110.850 ;
        RECT 108.880 110.550 116.800 110.560 ;
        RECT 105.110 110.540 116.800 110.550 ;
        RECT 101.490 110.420 116.800 110.540 ;
        RECT 101.490 110.410 116.825 110.420 ;
        RECT 101.450 110.290 116.825 110.410 ;
        RECT 101.450 110.180 105.450 110.290 ;
        RECT 101.060 109.840 101.290 110.130 ;
        RECT 101.510 109.840 105.400 110.180 ;
        RECT 105.610 109.840 105.840 110.130 ;
        RECT 101.060 108.470 105.840 109.840 ;
        RECT 101.060 108.170 101.290 108.470 ;
        RECT 105.610 108.170 105.840 108.470 ;
        RECT 101.450 107.890 105.450 108.120 ;
        RECT 101.700 107.660 105.270 107.890 ;
        RECT 101.700 107.510 105.390 107.660 ;
        RECT 100.000 107.230 105.390 107.510 ;
        RECT 106.640 107.340 107.260 110.290 ;
        RECT 108.825 110.190 116.825 110.290 ;
        RECT 108.880 110.180 116.800 110.190 ;
        RECT 108.390 109.480 108.620 110.140 ;
        RECT 109.400 109.480 110.400 109.570 ;
        RECT 117.030 109.480 117.260 110.140 ;
        RECT 108.390 108.660 117.260 109.480 ;
        RECT 108.390 108.180 108.620 108.660 ;
        RECT 109.400 108.570 110.400 108.660 ;
        RECT 117.030 108.180 117.260 108.660 ;
        RECT 108.825 107.900 116.825 108.130 ;
        RECT 77.045 106.980 77.810 107.120 ;
        RECT 76.125 106.935 76.415 106.980 ;
        RECT 77.045 106.935 77.335 106.980 ;
        RECT 60.010 106.780 60.330 106.840 ;
        RECT 65.070 106.780 65.390 106.840 ;
        RECT 67.920 106.780 68.060 106.935 ;
        RECT 77.490 106.920 77.810 106.980 ;
        RECT 78.040 106.980 82.320 107.120 ;
        RECT 56.420 106.640 60.330 106.780 ;
        RECT 60.010 106.580 60.330 106.640 ;
        RECT 63.780 106.640 68.060 106.780 ;
        RECT 74.270 106.780 74.590 106.840 ;
        RECT 78.040 106.780 78.180 106.980 ;
        RECT 84.850 106.920 85.170 107.180 ;
        RECT 86.230 106.920 86.550 107.180 ;
        RECT 86.705 107.120 86.995 107.165 ;
        RECT 87.610 107.120 87.930 107.180 ;
        RECT 86.705 106.980 87.930 107.120 ;
        RECT 86.705 106.935 86.995 106.980 ;
        RECT 87.610 106.920 87.930 106.980 ;
        RECT 78.410 106.825 78.730 106.840 ;
        RECT 74.270 106.640 78.180 106.780 ;
        RECT 63.780 106.500 63.920 106.640 ;
        RECT 65.070 106.580 65.390 106.640 ;
        RECT 74.270 106.580 74.590 106.640 ;
        RECT 78.380 106.595 78.730 106.825 ;
        RECT 85.785 106.595 86.075 106.825 ;
        RECT 100.000 106.770 105.400 107.230 ;
        RECT 78.410 106.580 78.730 106.595 ;
        RECT 48.510 106.440 48.830 106.500 ;
        RECT 44.460 106.300 48.830 106.440 ;
        RECT 32.885 106.255 33.175 106.300 ;
        RECT 36.090 106.240 36.410 106.300 ;
        RECT 48.510 106.240 48.830 106.300 ;
        RECT 54.030 106.240 54.350 106.500 ;
        RECT 59.090 106.440 59.410 106.500 ;
        RECT 61.850 106.440 62.170 106.500 ;
        RECT 59.090 106.300 62.170 106.440 ;
        RECT 59.090 106.240 59.410 106.300 ;
        RECT 61.850 106.240 62.170 106.300 ;
        RECT 63.690 106.240 64.010 106.500 ;
        RECT 64.610 106.440 64.930 106.500 ;
        RECT 66.005 106.440 66.295 106.485 ;
        RECT 64.610 106.300 66.295 106.440 ;
        RECT 64.610 106.240 64.930 106.300 ;
        RECT 66.005 106.255 66.295 106.300 ;
        RECT 66.465 106.440 66.755 106.485 ;
        RECT 71.970 106.440 72.290 106.500 ;
        RECT 66.465 106.300 72.290 106.440 ;
        RECT 66.465 106.255 66.755 106.300 ;
        RECT 71.970 106.240 72.290 106.300 ;
        RECT 75.205 106.440 75.495 106.485 ;
        RECT 82.550 106.440 82.870 106.500 ;
        RECT 75.205 106.300 82.870 106.440 ;
        RECT 85.860 106.440 86.000 106.595 ;
        RECT 86.690 106.440 87.010 106.500 ;
        RECT 85.860 106.300 87.010 106.440 ;
        RECT 75.205 106.255 75.495 106.300 ;
        RECT 82.550 106.240 82.870 106.300 ;
        RECT 86.690 106.240 87.010 106.300 ;
        RECT 12.100 105.620 89.840 106.100 ;
        RECT 23.670 105.420 23.990 105.480 ;
        RECT 19.160 105.280 23.990 105.420 ;
        RECT 19.160 105.125 19.300 105.280 ;
        RECT 23.670 105.220 23.990 105.280 ;
        RECT 26.905 105.420 27.195 105.465 ;
        RECT 27.350 105.420 27.670 105.480 ;
        RECT 30.570 105.420 30.890 105.480 ;
        RECT 26.905 105.280 30.890 105.420 ;
        RECT 26.905 105.235 27.195 105.280 ;
        RECT 27.350 105.220 27.670 105.280 ;
        RECT 30.570 105.220 30.890 105.280 ;
        RECT 32.870 105.420 33.190 105.480 ;
        RECT 33.345 105.420 33.635 105.465 ;
        RECT 32.870 105.280 33.635 105.420 ;
        RECT 32.870 105.220 33.190 105.280 ;
        RECT 33.345 105.235 33.635 105.280 ;
        RECT 33.805 105.235 34.095 105.465 ;
        RECT 38.850 105.420 39.170 105.480 ;
        RECT 35.260 105.280 39.170 105.420 ;
        RECT 19.085 104.895 19.375 105.125 ;
        RECT 24.605 105.080 24.895 105.125 ;
        RECT 25.050 105.080 25.370 105.140 ;
        RECT 20.310 104.940 25.370 105.080 ;
        RECT 16.325 104.740 16.615 104.785 ;
        RECT 20.310 104.740 20.450 104.940 ;
        RECT 24.605 104.895 24.895 104.940 ;
        RECT 16.325 104.600 20.450 104.740 ;
        RECT 20.925 104.740 21.215 104.785 ;
        RECT 23.220 104.740 23.510 104.785 ;
        RECT 20.925 104.600 23.510 104.740 ;
        RECT 16.325 104.555 16.615 104.600 ;
        RECT 20.925 104.555 21.215 104.600 ;
        RECT 23.220 104.555 23.510 104.600 ;
        RECT 23.685 104.740 23.975 104.785 ;
        RECT 24.680 104.740 24.820 104.895 ;
        RECT 25.050 104.880 25.370 104.940 ;
        RECT 26.430 105.080 26.750 105.140 ;
        RECT 33.880 105.080 34.020 105.235 ;
        RECT 35.260 105.080 35.400 105.280 ;
        RECT 38.850 105.220 39.170 105.280 ;
        RECT 48.065 105.420 48.355 105.465 ;
        RECT 48.510 105.420 48.830 105.480 ;
        RECT 48.065 105.280 48.830 105.420 ;
        RECT 48.065 105.235 48.355 105.280 ;
        RECT 48.510 105.220 48.830 105.280 ;
        RECT 60.010 105.220 60.330 105.480 ;
        RECT 60.930 105.220 61.250 105.480 ;
        RECT 61.850 105.420 62.170 105.480 ;
        RECT 62.785 105.420 63.075 105.465 ;
        RECT 61.850 105.280 63.075 105.420 ;
        RECT 61.850 105.220 62.170 105.280 ;
        RECT 62.785 105.235 63.075 105.280 ;
        RECT 64.610 105.220 64.930 105.480 ;
        RECT 68.765 105.420 69.055 105.465 ;
        RECT 71.525 105.420 71.815 105.465 ;
        RECT 68.765 105.280 71.815 105.420 ;
        RECT 68.765 105.235 69.055 105.280 ;
        RECT 71.525 105.235 71.815 105.280 ;
        RECT 77.045 105.420 77.335 105.465 ;
        RECT 78.410 105.420 78.730 105.480 ;
        RECT 79.330 105.420 79.650 105.480 ;
        RECT 100.000 105.430 102.000 106.770 ;
        RECT 103.750 106.760 105.400 106.770 ;
        RECT 102.440 105.490 103.440 106.210 ;
        RECT 103.750 105.950 104.060 106.760 ;
        RECT 104.520 106.480 105.400 106.760 ;
        RECT 105.640 106.940 107.260 107.340 ;
        RECT 108.910 106.990 116.780 107.900 ;
        RECT 104.460 106.250 105.460 106.480 ;
        RECT 105.640 106.290 105.990 106.940 ;
        RECT 106.640 106.930 107.260 106.940 ;
        RECT 108.825 106.760 116.825 106.990 ;
        RECT 108.910 106.750 116.780 106.760 ;
        RECT 104.520 106.040 105.400 106.060 ;
        RECT 103.790 105.660 104.060 105.950 ;
        RECT 104.460 105.810 105.460 106.040 ;
        RECT 105.620 106.000 105.990 106.290 ;
        RECT 105.650 105.940 105.990 106.000 ;
        RECT 106.750 106.610 107.510 106.660 ;
        RECT 108.390 106.610 108.620 106.710 ;
        RECT 106.750 106.400 108.620 106.610 ;
        RECT 117.030 106.400 117.260 106.710 ;
        RECT 106.750 105.980 109.290 106.400 ;
        RECT 116.660 105.980 117.260 106.400 ;
        RECT 104.520 105.660 105.400 105.810 ;
        RECT 104.530 105.490 105.260 105.660 ;
        RECT 100.080 105.420 102.000 105.430 ;
        RECT 77.045 105.280 78.730 105.420 ;
        RECT 77.045 105.235 77.335 105.280 ;
        RECT 78.410 105.220 78.730 105.280 ;
        RECT 78.960 105.280 79.650 105.420 ;
        RECT 26.430 104.940 34.020 105.080 ;
        RECT 34.800 104.940 35.400 105.080 ;
        RECT 26.430 104.880 26.750 104.940 ;
        RECT 26.890 104.740 27.210 104.800 ;
        RECT 27.365 104.740 27.655 104.785 ;
        RECT 23.685 104.600 27.655 104.740 ;
        RECT 23.685 104.555 23.975 104.600 ;
        RECT 16.785 104.400 17.075 104.445 ;
        RECT 21.000 104.400 21.140 104.555 ;
        RECT 16.785 104.260 21.140 104.400 ;
        RECT 23.300 104.400 23.440 104.555 ;
        RECT 26.890 104.540 27.210 104.600 ;
        RECT 27.365 104.555 27.655 104.600 ;
        RECT 27.810 104.540 28.130 104.800 ;
        RECT 30.110 104.740 30.430 104.800 ;
        RECT 31.045 104.740 31.335 104.785 ;
        RECT 30.110 104.600 31.335 104.740 ;
        RECT 30.110 104.540 30.430 104.600 ;
        RECT 31.045 104.555 31.335 104.600 ;
        RECT 32.410 104.540 32.730 104.800 ;
        RECT 34.800 104.785 34.940 104.940 ;
        RECT 36.090 104.880 36.410 105.140 ;
        RECT 34.725 104.740 35.015 104.785 ;
        RECT 33.880 104.600 35.015 104.740 ;
        RECT 28.730 104.400 29.050 104.460 ;
        RECT 31.965 104.400 32.255 104.445 ;
        RECT 33.880 104.400 34.020 104.600 ;
        RECT 34.725 104.555 35.015 104.600 ;
        RECT 35.185 104.740 35.475 104.785 ;
        RECT 35.630 104.740 35.950 104.800 ;
        RECT 35.185 104.600 35.950 104.740 ;
        RECT 35.185 104.555 35.475 104.600 ;
        RECT 35.630 104.540 35.950 104.600 ;
        RECT 42.500 104.740 42.790 104.785 ;
        RECT 44.370 104.740 44.690 104.800 ;
        RECT 48.600 104.785 48.740 105.220 ;
        RECT 49.890 105.080 50.210 105.140 ;
        RECT 50.365 105.080 50.655 105.125 ;
        RECT 49.890 104.940 50.655 105.080 ;
        RECT 49.890 104.880 50.210 104.940 ;
        RECT 50.365 104.895 50.655 104.940 ;
        RECT 53.080 105.080 53.370 105.125 ;
        RECT 54.030 105.080 54.350 105.140 ;
        RECT 64.700 105.080 64.840 105.220 ;
        RECT 53.080 104.940 54.350 105.080 ;
        RECT 53.080 104.895 53.370 104.940 ;
        RECT 54.030 104.880 54.350 104.940 ;
        RECT 60.560 104.940 64.840 105.080 ;
        RECT 66.925 105.080 67.215 105.125 ;
        RECT 68.290 105.080 68.610 105.140 ;
        RECT 72.430 105.080 72.750 105.140 ;
        RECT 75.190 105.080 75.510 105.140 ;
        RECT 78.960 105.080 79.100 105.280 ;
        RECT 79.330 105.220 79.650 105.280 ;
        RECT 81.170 105.080 81.490 105.140 ;
        RECT 84.390 105.080 84.710 105.140 ;
        RECT 66.925 104.940 68.750 105.080 ;
        RECT 42.500 104.600 44.690 104.740 ;
        RECT 42.500 104.555 42.790 104.600 ;
        RECT 44.370 104.540 44.690 104.600 ;
        RECT 48.525 104.555 48.815 104.785 ;
        RECT 59.565 104.740 59.855 104.785 ;
        RECT 60.010 104.740 60.330 104.800 ;
        RECT 60.560 104.785 60.700 104.940 ;
        RECT 66.925 104.895 67.215 104.940 ;
        RECT 68.290 104.880 68.750 104.940 ;
        RECT 72.430 104.940 79.100 105.080 ;
        RECT 72.430 104.880 72.750 104.940 ;
        RECT 75.190 104.880 75.510 104.940 ;
        RECT 59.565 104.600 60.330 104.740 ;
        RECT 59.565 104.555 59.855 104.600 ;
        RECT 60.010 104.540 60.330 104.600 ;
        RECT 60.485 104.555 60.775 104.785 ;
        RECT 61.865 104.740 62.155 104.785 ;
        RECT 62.310 104.740 62.630 104.800 ;
        RECT 63.230 104.740 63.550 104.800 ;
        RECT 61.865 104.600 62.630 104.740 ;
        RECT 63.135 104.600 63.550 104.740 ;
        RECT 64.165 104.730 64.455 104.785 ;
        RECT 61.865 104.555 62.155 104.600 ;
        RECT 62.310 104.540 62.630 104.600 ;
        RECT 63.230 104.540 63.550 104.600 ;
        RECT 63.780 104.590 64.455 104.730 ;
        RECT 23.300 104.260 26.660 104.400 ;
        RECT 16.785 104.215 17.075 104.260 ;
        RECT 26.520 104.120 26.660 104.260 ;
        RECT 28.730 104.260 34.020 104.400 ;
        RECT 28.730 104.200 29.050 104.260 ;
        RECT 31.965 104.215 32.255 104.260 ;
        RECT 41.150 104.200 41.470 104.460 ;
        RECT 42.045 104.400 42.335 104.445 ;
        RECT 43.235 104.400 43.525 104.445 ;
        RECT 45.755 104.400 46.045 104.445 ;
        RECT 42.045 104.260 46.045 104.400 ;
        RECT 42.045 104.215 42.335 104.260 ;
        RECT 43.235 104.215 43.525 104.260 ;
        RECT 45.755 104.215 46.045 104.260 ;
        RECT 48.050 104.400 48.370 104.460 ;
        RECT 51.745 104.400 52.035 104.445 ;
        RECT 48.050 104.260 52.035 104.400 ;
        RECT 48.050 104.200 48.370 104.260 ;
        RECT 51.745 104.215 52.035 104.260 ;
        RECT 52.625 104.400 52.915 104.445 ;
        RECT 53.815 104.400 54.105 104.445 ;
        RECT 56.335 104.400 56.625 104.445 ;
        RECT 52.625 104.260 56.625 104.400 ;
        RECT 52.625 104.215 52.915 104.260 ;
        RECT 53.815 104.215 54.105 104.260 ;
        RECT 56.335 104.215 56.625 104.260 ;
        RECT 58.170 104.400 58.490 104.460 ;
        RECT 63.320 104.400 63.460 104.540 ;
        RECT 58.170 104.260 63.460 104.400 ;
        RECT 58.170 104.200 58.490 104.260 ;
        RECT 26.430 103.860 26.750 104.120 ;
        RECT 29.190 104.060 29.510 104.120 ;
        RECT 31.505 104.060 31.795 104.105 ;
        RECT 29.190 103.920 31.795 104.060 ;
        RECT 29.190 103.860 29.510 103.920 ;
        RECT 31.505 103.875 31.795 103.920 ;
        RECT 41.650 104.060 41.940 104.105 ;
        RECT 43.750 104.060 44.040 104.105 ;
        RECT 45.320 104.060 45.610 104.105 ;
        RECT 41.650 103.920 45.610 104.060 ;
        RECT 41.650 103.875 41.940 103.920 ;
        RECT 43.750 103.875 44.040 103.920 ;
        RECT 45.320 103.875 45.610 103.920 ;
        RECT 52.230 104.060 52.520 104.105 ;
        RECT 54.330 104.060 54.620 104.105 ;
        RECT 55.900 104.060 56.190 104.105 ;
        RECT 52.230 103.920 56.190 104.060 ;
        RECT 52.230 103.875 52.520 103.920 ;
        RECT 54.330 103.875 54.620 103.920 ;
        RECT 55.900 103.875 56.190 103.920 ;
        RECT 56.790 104.060 57.110 104.120 ;
        RECT 59.550 104.060 59.870 104.120 ;
        RECT 63.780 104.060 63.920 104.590 ;
        RECT 64.165 104.555 64.455 104.590 ;
        RECT 65.070 104.540 65.390 104.800 ;
        RECT 65.990 104.540 66.310 104.800 ;
        RECT 67.370 104.540 67.690 104.800 ;
        RECT 67.830 104.540 68.150 104.800 ;
        RECT 68.610 104.740 68.750 104.880 ;
        RECT 70.130 104.740 70.450 104.800 ;
        RECT 78.960 104.785 79.100 104.940 ;
        RECT 80.340 104.940 84.710 105.080 ;
        RECT 68.610 104.600 70.450 104.740 ;
        RECT 70.130 104.540 70.450 104.600 ;
        RECT 71.065 104.740 71.355 104.785 ;
        RECT 73.365 104.740 73.655 104.785 ;
        RECT 78.425 104.740 78.715 104.785 ;
        RECT 71.065 104.600 73.655 104.740 ;
        RECT 71.065 104.555 71.355 104.600 ;
        RECT 73.365 104.555 73.655 104.600 ;
        RECT 77.580 104.600 78.715 104.740 ;
        RECT 71.970 104.200 72.290 104.460 ;
        RECT 76.110 104.200 76.430 104.460 ;
        RECT 56.790 103.920 63.920 104.060 ;
        RECT 77.580 104.060 77.720 104.600 ;
        RECT 78.425 104.555 78.715 104.600 ;
        RECT 78.885 104.555 79.175 104.785 ;
        RECT 79.330 104.540 79.650 104.800 ;
        RECT 80.340 104.785 80.480 104.940 ;
        RECT 81.170 104.880 81.490 104.940 ;
        RECT 84.390 104.880 84.710 104.940 ;
        RECT 80.265 104.555 80.555 104.785 ;
        RECT 81.630 104.740 81.950 104.800 ;
        RECT 82.465 104.740 82.755 104.785 ;
        RECT 81.630 104.600 82.755 104.740 ;
        RECT 81.630 104.540 81.950 104.600 ;
        RECT 82.465 104.555 82.755 104.600 ;
        RECT 77.950 104.400 78.270 104.460 ;
        RECT 81.185 104.400 81.475 104.445 ;
        RECT 77.950 104.260 81.475 104.400 ;
        RECT 77.950 104.200 78.270 104.260 ;
        RECT 81.185 104.215 81.475 104.260 ;
        RECT 82.065 104.400 82.355 104.445 ;
        RECT 83.255 104.400 83.545 104.445 ;
        RECT 85.775 104.400 86.065 104.445 ;
        RECT 82.065 104.260 86.065 104.400 ;
        RECT 102.410 104.370 105.260 105.490 ;
        RECT 105.650 105.190 106.000 105.940 ;
        RECT 106.750 105.820 108.620 105.980 ;
        RECT 106.750 105.770 107.510 105.820 ;
        RECT 108.390 105.750 108.620 105.820 ;
        RECT 117.030 105.750 117.260 105.980 ;
        RECT 108.825 105.470 116.825 105.700 ;
        RECT 105.650 105.130 105.940 105.190 ;
        RECT 105.560 105.010 105.940 105.130 ;
        RECT 108.920 105.070 116.780 105.470 ;
        RECT 117.590 105.070 118.560 114.550 ;
        RECT 119.930 114.680 120.770 116.810 ;
        RECT 126.430 116.390 127.680 116.830 ;
        RECT 137.600 116.810 138.460 118.930 ;
        RECT 124.370 116.380 129.610 116.390 ;
        RECT 121.420 116.280 136.720 116.380 ;
        RECT 121.420 116.270 136.755 116.280 ;
        RECT 121.380 116.150 136.755 116.270 ;
        RECT 121.380 116.040 125.380 116.150 ;
        RECT 126.430 116.070 128.170 116.150 ;
        RECT 128.750 116.070 136.755 116.150 ;
        RECT 126.430 115.990 127.680 116.070 ;
        RECT 128.755 116.050 136.755 116.070 ;
        RECT 120.990 115.740 121.220 115.990 ;
        RECT 125.540 115.850 125.770 115.990 ;
        RECT 128.320 115.850 128.550 116.000 ;
        RECT 125.540 115.740 128.550 115.850 ;
        RECT 136.960 115.740 137.190 116.000 ;
        RECT 120.990 115.300 137.190 115.740 ;
        RECT 120.990 115.030 121.220 115.300 ;
        RECT 125.540 115.270 137.190 115.300 ;
        RECT 125.540 115.180 128.550 115.270 ;
        RECT 125.540 115.030 125.770 115.180 ;
        RECT 128.320 115.040 128.550 115.180 ;
        RECT 136.960 115.040 137.190 115.270 ;
        RECT 121.380 114.750 125.380 114.980 ;
        RECT 128.755 114.770 136.755 114.990 ;
        RECT 137.520 114.770 138.480 116.810 ;
        RECT 128.755 114.760 138.480 114.770 ;
        RECT 121.380 114.680 125.370 114.750 ;
        RECT 119.930 114.570 125.370 114.680 ;
        RECT 128.810 114.600 138.480 114.760 ;
        RECT 119.930 114.480 123.060 114.570 ;
        RECT 136.550 114.550 138.480 114.600 ;
        RECT 119.930 111.210 120.770 114.480 ;
        RECT 124.410 114.020 129.660 114.030 ;
        RECT 124.410 113.910 136.720 114.020 ;
        RECT 121.440 113.850 136.720 113.910 ;
        RECT 121.440 113.840 136.755 113.850 ;
        RECT 121.380 113.710 136.755 113.840 ;
        RECT 121.380 113.700 126.540 113.710 ;
        RECT 121.380 113.610 125.380 113.700 ;
        RECT 128.755 113.620 136.755 113.710 ;
        RECT 128.840 113.610 136.730 113.620 ;
        RECT 120.990 113.250 121.220 113.560 ;
        RECT 121.440 113.250 125.340 113.610 ;
        RECT 125.540 113.250 125.770 113.560 ;
        RECT 120.990 111.910 125.770 113.250 ;
        RECT 120.990 111.600 121.220 111.910 ;
        RECT 125.540 111.600 125.770 111.910 ;
        RECT 128.320 113.030 128.550 113.570 ;
        RECT 129.360 113.030 130.370 113.060 ;
        RECT 136.960 113.030 137.190 113.570 ;
        RECT 128.320 112.130 137.190 113.030 ;
        RECT 128.320 111.610 128.550 112.130 ;
        RECT 129.360 112.060 130.370 112.130 ;
        RECT 136.960 111.610 137.190 112.130 ;
        RECT 121.380 111.320 125.380 111.550 ;
        RECT 128.755 111.330 136.755 111.560 ;
        RECT 119.930 111.170 121.060 111.210 ;
        RECT 119.930 111.090 121.300 111.170 ;
        RECT 121.670 111.100 125.330 111.320 ;
        RECT 121.670 111.090 123.110 111.100 ;
        RECT 119.930 111.050 123.110 111.090 ;
        RECT 119.930 110.960 122.620 111.050 ;
        RECT 128.820 111.040 136.710 111.330 ;
        RECT 119.930 110.900 121.950 110.960 ;
        RECT 119.930 110.850 121.700 110.900 ;
        RECT 119.930 107.510 120.770 110.850 ;
        RECT 128.810 110.550 136.730 110.560 ;
        RECT 125.040 110.540 136.730 110.550 ;
        RECT 121.420 110.420 136.730 110.540 ;
        RECT 121.420 110.410 136.755 110.420 ;
        RECT 121.380 110.290 136.755 110.410 ;
        RECT 121.380 110.180 125.380 110.290 ;
        RECT 120.990 109.840 121.220 110.130 ;
        RECT 121.440 109.840 125.330 110.180 ;
        RECT 125.540 109.840 125.770 110.130 ;
        RECT 120.990 108.470 125.770 109.840 ;
        RECT 120.990 108.170 121.220 108.470 ;
        RECT 125.540 108.170 125.770 108.470 ;
        RECT 121.380 107.890 125.380 108.120 ;
        RECT 121.630 107.660 125.200 107.890 ;
        RECT 121.630 107.510 125.320 107.660 ;
        RECT 119.930 107.230 125.320 107.510 ;
        RECT 126.570 107.340 127.190 110.290 ;
        RECT 128.755 110.190 136.755 110.290 ;
        RECT 128.810 110.180 136.730 110.190 ;
        RECT 128.320 109.480 128.550 110.140 ;
        RECT 129.330 109.480 130.330 109.570 ;
        RECT 136.960 109.480 137.190 110.140 ;
        RECT 128.320 108.660 137.190 109.480 ;
        RECT 128.320 108.180 128.550 108.660 ;
        RECT 129.330 108.570 130.330 108.660 ;
        RECT 136.960 108.180 137.190 108.660 ;
        RECT 128.755 107.900 136.755 108.130 ;
        RECT 119.930 106.770 125.330 107.230 ;
        RECT 119.930 105.880 121.930 106.770 ;
        RECT 123.680 106.760 125.330 106.770 ;
        RECT 82.065 104.215 82.355 104.260 ;
        RECT 83.255 104.215 83.545 104.260 ;
        RECT 85.775 104.215 86.065 104.260 ;
        RECT 102.350 104.140 105.350 104.370 ;
        RECT 105.560 104.180 105.900 105.010 ;
        RECT 107.910 105.000 118.560 105.070 ;
        RECT 102.400 104.110 105.260 104.140 ;
        RECT 81.670 104.060 81.960 104.105 ;
        RECT 83.770 104.060 84.060 104.105 ;
        RECT 85.340 104.060 85.630 104.105 ;
        RECT 102.400 104.090 103.570 104.110 ;
        RECT 104.530 104.100 105.260 104.110 ;
        RECT 77.580 103.920 78.180 104.060 ;
        RECT 56.790 103.860 57.110 103.920 ;
        RECT 59.550 103.860 59.870 103.920 ;
        RECT 18.150 103.720 18.470 103.780 ;
        RECT 19.990 103.720 20.310 103.780 ;
        RECT 18.150 103.580 20.310 103.720 ;
        RECT 18.150 103.520 18.470 103.580 ;
        RECT 19.990 103.520 20.310 103.580 ;
        RECT 22.290 103.720 22.610 103.780 ;
        RECT 22.765 103.720 23.055 103.765 ;
        RECT 22.290 103.580 23.055 103.720 ;
        RECT 22.290 103.520 22.610 103.580 ;
        RECT 22.765 103.535 23.055 103.580 ;
        RECT 28.270 103.720 28.590 103.780 ;
        RECT 30.110 103.720 30.430 103.780 ;
        RECT 28.270 103.580 30.430 103.720 ;
        RECT 28.270 103.520 28.590 103.580 ;
        RECT 30.110 103.520 30.430 103.580 ;
        RECT 36.105 103.720 36.395 103.765 ;
        RECT 39.310 103.720 39.630 103.780 ;
        RECT 36.105 103.580 39.630 103.720 ;
        RECT 36.105 103.535 36.395 103.580 ;
        RECT 39.310 103.520 39.630 103.580 ;
        RECT 39.770 103.720 40.090 103.780 ;
        RECT 47.130 103.720 47.450 103.780 ;
        RECT 39.770 103.580 47.450 103.720 ;
        RECT 39.770 103.520 40.090 103.580 ;
        RECT 47.130 103.520 47.450 103.580 ;
        RECT 50.350 103.520 50.670 103.780 ;
        RECT 51.285 103.720 51.575 103.765 ;
        RECT 53.570 103.720 53.890 103.780 ;
        RECT 51.285 103.580 53.890 103.720 ;
        RECT 51.285 103.535 51.575 103.580 ;
        RECT 53.570 103.520 53.890 103.580 ;
        RECT 56.330 103.720 56.650 103.780 ;
        RECT 58.645 103.720 58.935 103.765 ;
        RECT 56.330 103.580 58.935 103.720 ;
        RECT 56.330 103.520 56.650 103.580 ;
        RECT 58.645 103.535 58.935 103.580 ;
        RECT 69.210 103.520 69.530 103.780 ;
        RECT 78.040 103.720 78.180 103.920 ;
        RECT 81.670 103.920 85.630 104.060 ;
        RECT 81.670 103.875 81.960 103.920 ;
        RECT 83.770 103.875 84.060 103.920 ;
        RECT 85.340 103.875 85.630 103.920 ;
        RECT 82.090 103.720 82.410 103.780 ;
        RECT 78.040 103.580 82.410 103.720 ;
        RECT 82.090 103.520 82.410 103.580 ;
        RECT 86.230 103.720 86.550 103.780 ;
        RECT 88.085 103.720 88.375 103.765 ;
        RECT 86.230 103.580 88.375 103.720 ;
        RECT 102.350 103.700 105.350 103.930 ;
        RECT 105.555 103.890 105.900 104.180 ;
        RECT 106.090 104.040 118.560 105.000 ;
        RECT 119.900 105.420 121.930 105.880 ;
        RECT 122.370 105.490 123.370 106.210 ;
        RECT 123.680 105.950 123.990 106.760 ;
        RECT 124.450 106.480 125.330 106.760 ;
        RECT 125.570 106.940 127.190 107.340 ;
        RECT 128.840 106.990 136.710 107.900 ;
        RECT 124.390 106.250 125.390 106.480 ;
        RECT 125.570 106.290 125.920 106.940 ;
        RECT 126.570 106.930 127.190 106.940 ;
        RECT 128.755 106.760 136.755 106.990 ;
        RECT 128.840 106.750 136.710 106.760 ;
        RECT 124.450 106.040 125.330 106.060 ;
        RECT 123.720 105.660 123.990 105.950 ;
        RECT 124.390 105.810 125.390 106.040 ;
        RECT 125.550 106.000 125.920 106.290 ;
        RECT 125.580 105.940 125.920 106.000 ;
        RECT 126.680 106.610 127.440 106.660 ;
        RECT 128.320 106.610 128.550 106.710 ;
        RECT 126.680 106.400 128.550 106.610 ;
        RECT 136.960 106.400 137.190 106.710 ;
        RECT 126.680 105.980 129.220 106.400 ;
        RECT 136.590 105.980 137.190 106.400 ;
        RECT 124.450 105.660 125.330 105.810 ;
        RECT 124.460 105.490 125.190 105.660 ;
        RECT 106.090 103.960 118.550 104.040 ;
        RECT 106.090 103.940 118.420 103.960 ;
        RECT 105.560 103.780 105.900 103.890 ;
        RECT 106.130 103.930 111.800 103.940 ;
        RECT 112.800 103.930 118.420 103.940 ;
        RECT 86.230 103.520 86.550 103.580 ;
        RECT 88.085 103.535 88.375 103.580 ;
        RECT 102.440 103.530 105.300 103.700 ;
        RECT 106.130 103.530 107.465 103.930 ;
        RECT 12.100 102.900 89.840 103.380 ;
        RECT 102.410 103.160 107.465 103.530 ;
        RECT 106.195 102.975 107.465 103.160 ;
        RECT 50.810 102.700 51.130 102.760 ;
        RECT 51.285 102.700 51.575 102.745 ;
        RECT 37.100 102.560 49.200 102.700 ;
        RECT 37.100 101.725 37.240 102.560 ;
        RECT 43.910 102.360 44.200 102.405 ;
        RECT 45.480 102.360 45.770 102.405 ;
        RECT 47.580 102.360 47.870 102.405 ;
        RECT 43.910 102.220 47.870 102.360 ;
        RECT 43.910 102.175 44.200 102.220 ;
        RECT 45.480 102.175 45.770 102.220 ;
        RECT 47.580 102.175 47.870 102.220 ;
        RECT 43.475 102.020 43.765 102.065 ;
        RECT 45.995 102.020 46.285 102.065 ;
        RECT 47.185 102.020 47.475 102.065 ;
        RECT 43.475 101.880 47.475 102.020 ;
        RECT 43.475 101.835 43.765 101.880 ;
        RECT 45.995 101.835 46.285 101.880 ;
        RECT 47.185 101.835 47.475 101.880 ;
        RECT 49.060 102.020 49.200 102.560 ;
        RECT 50.810 102.560 51.575 102.700 ;
        RECT 50.810 102.500 51.130 102.560 ;
        RECT 51.285 102.515 51.575 102.560 ;
        RECT 51.730 102.700 52.050 102.760 ;
        RECT 56.790 102.700 57.110 102.760 ;
        RECT 51.730 102.560 57.110 102.700 ;
        RECT 51.730 102.500 52.050 102.560 ;
        RECT 56.790 102.500 57.110 102.560 ;
        RECT 57.265 102.700 57.555 102.745 ;
        RECT 58.170 102.700 58.490 102.760 ;
        RECT 57.265 102.560 58.490 102.700 ;
        RECT 57.265 102.515 57.555 102.560 ;
        RECT 58.170 102.500 58.490 102.560 ;
        RECT 60.025 102.700 60.315 102.745 ;
        RECT 65.070 102.700 65.390 102.760 ;
        RECT 60.025 102.560 65.390 102.700 ;
        RECT 60.025 102.515 60.315 102.560 ;
        RECT 65.070 102.500 65.390 102.560 ;
        RECT 65.990 102.500 66.310 102.760 ;
        RECT 69.670 102.700 69.990 102.760 ;
        RECT 66.540 102.560 69.990 102.700 ;
        RECT 49.430 102.360 49.750 102.420 ;
        RECT 49.905 102.360 50.195 102.405 ;
        RECT 55.410 102.360 55.730 102.420 ;
        RECT 49.430 102.220 55.730 102.360 ;
        RECT 49.430 102.160 49.750 102.220 ;
        RECT 49.905 102.175 50.195 102.220 ;
        RECT 55.410 102.160 55.730 102.220 ;
        RECT 56.330 102.160 56.650 102.420 ;
        RECT 59.105 102.175 59.395 102.405 ;
        RECT 62.310 102.360 62.630 102.420 ;
        RECT 60.560 102.220 62.630 102.360 ;
        RECT 53.125 102.020 53.415 102.065 ;
        RECT 49.060 101.880 53.415 102.020 ;
        RECT 49.060 101.740 49.200 101.880 ;
        RECT 53.125 101.835 53.415 101.880 ;
        RECT 54.950 102.020 55.270 102.080 ;
        RECT 59.180 102.020 59.320 102.175 ;
        RECT 54.950 101.880 59.320 102.020 ;
        RECT 54.950 101.820 55.270 101.880 ;
        RECT 36.105 101.495 36.395 101.725 ;
        RECT 37.025 101.495 37.315 101.725 ;
        RECT 37.945 101.495 38.235 101.725 ;
        RECT 41.150 101.680 41.470 101.740 ;
        RECT 48.050 101.680 48.370 101.740 ;
        RECT 41.150 101.540 48.370 101.680 ;
        RECT 36.180 101.340 36.320 101.495 ;
        RECT 38.020 101.340 38.160 101.495 ;
        RECT 41.150 101.480 41.470 101.540 ;
        RECT 48.050 101.480 48.370 101.540 ;
        RECT 48.970 101.480 49.290 101.740 ;
        RECT 50.365 101.680 50.655 101.725 ;
        RECT 54.030 101.680 54.350 101.740 ;
        RECT 50.365 101.540 54.350 101.680 ;
        RECT 50.365 101.495 50.655 101.540 ;
        RECT 54.030 101.480 54.350 101.540 ;
        RECT 54.490 101.480 54.810 101.740 ;
        RECT 58.630 101.680 58.950 101.740 ;
        RECT 60.560 101.680 60.700 102.220 ;
        RECT 62.310 102.160 62.630 102.220 ;
        RECT 60.930 102.020 61.250 102.080 ;
        RECT 63.245 102.020 63.535 102.065 ;
        RECT 60.930 101.880 63.535 102.020 ;
        RECT 60.930 101.820 61.250 101.880 ;
        RECT 63.245 101.835 63.535 101.880 ;
        RECT 58.630 101.540 60.700 101.680 ;
        RECT 58.630 101.480 58.950 101.540 ;
        RECT 61.405 101.495 61.695 101.725 ;
        RECT 61.850 101.680 62.170 101.740 ;
        RECT 62.325 101.680 62.615 101.725 ;
        RECT 61.850 101.540 62.615 101.680 ;
        RECT 36.180 101.200 38.160 101.340 ;
        RECT 36.550 100.800 36.870 101.060 ;
        RECT 38.020 101.000 38.160 101.200 ;
        RECT 40.705 101.340 40.995 101.385 ;
        RECT 41.610 101.340 41.930 101.400 ;
        RECT 46.840 101.340 47.130 101.385 ;
        RECT 47.590 101.340 47.910 101.400 ;
        RECT 52.190 101.385 52.510 101.400 ;
        RECT 40.705 101.200 45.980 101.340 ;
        RECT 40.705 101.155 40.995 101.200 ;
        RECT 41.610 101.140 41.930 101.200 ;
        RECT 45.840 101.060 45.980 101.200 ;
        RECT 46.840 101.200 47.910 101.340 ;
        RECT 46.840 101.155 47.130 101.200 ;
        RECT 47.590 101.140 47.910 101.200 ;
        RECT 52.080 101.340 52.510 101.385 ;
        RECT 53.110 101.340 53.430 101.400 ;
        RECT 52.080 101.200 53.430 101.340 ;
        RECT 52.080 101.155 52.510 101.200 ;
        RECT 52.190 101.140 52.510 101.155 ;
        RECT 53.110 101.140 53.430 101.200 ;
        RECT 56.330 101.340 56.650 101.400 ;
        RECT 57.725 101.340 58.015 101.385 ;
        RECT 56.330 101.200 58.015 101.340 ;
        RECT 56.330 101.140 56.650 101.200 ;
        RECT 57.725 101.155 58.015 101.200 ;
        RECT 59.550 101.340 59.870 101.400 ;
        RECT 61.480 101.340 61.620 101.495 ;
        RECT 61.850 101.480 62.170 101.540 ;
        RECT 62.325 101.495 62.615 101.540 ;
        RECT 62.770 101.480 63.090 101.740 ;
        RECT 64.165 101.495 64.455 101.725 ;
        RECT 64.610 101.680 64.930 101.740 ;
        RECT 66.540 101.725 66.680 102.560 ;
        RECT 69.670 102.500 69.990 102.560 ;
        RECT 77.030 102.700 77.350 102.760 ;
        RECT 77.965 102.700 78.255 102.745 ;
        RECT 77.030 102.560 78.255 102.700 ;
        RECT 77.030 102.500 77.350 102.560 ;
        RECT 77.965 102.515 78.255 102.560 ;
        RECT 81.185 102.700 81.475 102.745 ;
        RECT 81.630 102.700 81.950 102.760 ;
        RECT 83.470 102.700 83.790 102.760 ;
        RECT 81.185 102.560 81.950 102.700 ;
        RECT 81.185 102.515 81.475 102.560 ;
        RECT 81.630 102.500 81.950 102.560 ;
        RECT 82.180 102.560 83.790 102.700 ;
        RECT 68.330 102.360 68.620 102.405 ;
        RECT 70.430 102.360 70.720 102.405 ;
        RECT 72.000 102.360 72.290 102.405 ;
        RECT 68.330 102.220 72.290 102.360 ;
        RECT 68.330 102.175 68.620 102.220 ;
        RECT 70.430 102.175 70.720 102.220 ;
        RECT 72.000 102.175 72.290 102.220 ;
        RECT 74.745 102.360 75.035 102.405 ;
        RECT 76.110 102.360 76.430 102.420 ;
        RECT 74.745 102.220 76.430 102.360 ;
        RECT 74.745 102.175 75.035 102.220 ;
        RECT 76.110 102.160 76.430 102.220 ;
        RECT 68.725 102.020 69.015 102.065 ;
        RECT 69.915 102.020 70.205 102.065 ;
        RECT 72.435 102.020 72.725 102.065 ;
        RECT 82.180 102.020 82.320 102.560 ;
        RECT 83.470 102.500 83.790 102.560 ;
        RECT 82.550 102.360 82.870 102.420 ;
        RECT 82.550 102.220 86.000 102.360 ;
        RECT 82.550 102.160 82.870 102.220 ;
        RECT 83.930 102.020 84.250 102.080 ;
        RECT 68.725 101.880 72.725 102.020 ;
        RECT 68.725 101.835 69.015 101.880 ;
        RECT 69.915 101.835 70.205 101.880 ;
        RECT 72.435 101.835 72.725 101.880 ;
        RECT 78.960 101.880 82.320 102.020 ;
        RECT 83.100 101.880 84.250 102.020 ;
        RECT 65.545 101.680 65.835 101.725 ;
        RECT 64.610 101.540 65.835 101.680 ;
        RECT 63.690 101.340 64.010 101.400 ;
        RECT 59.550 101.200 64.010 101.340 ;
        RECT 59.550 101.140 59.870 101.200 ;
        RECT 63.690 101.140 64.010 101.200 ;
        RECT 41.165 101.000 41.455 101.045 ;
        RECT 42.070 101.000 42.390 101.060 ;
        RECT 38.020 100.860 42.390 101.000 ;
        RECT 41.165 100.815 41.455 100.860 ;
        RECT 42.070 100.800 42.390 100.860 ;
        RECT 45.750 100.800 46.070 101.060 ;
        RECT 48.050 101.000 48.370 101.060 ;
        RECT 49.890 101.000 50.210 101.060 ;
        RECT 52.665 101.000 52.955 101.045 ;
        RECT 48.050 100.860 52.955 101.000 ;
        RECT 48.050 100.800 48.370 100.860 ;
        RECT 49.890 100.800 50.210 100.860 ;
        RECT 52.665 100.815 52.955 100.860 ;
        RECT 55.410 101.000 55.730 101.060 ;
        RECT 60.010 101.000 60.330 101.060 ;
        RECT 60.930 101.000 61.250 101.060 ;
        RECT 64.240 101.000 64.380 101.495 ;
        RECT 64.610 101.480 64.930 101.540 ;
        RECT 65.545 101.495 65.835 101.540 ;
        RECT 66.465 101.495 66.755 101.725 ;
        RECT 67.830 101.480 68.150 101.740 ;
        RECT 69.210 101.725 69.530 101.740 ;
        RECT 69.180 101.680 69.530 101.725 ;
        RECT 69.015 101.540 69.530 101.680 ;
        RECT 69.180 101.495 69.530 101.540 ;
        RECT 69.210 101.480 69.530 101.495 ;
        RECT 76.110 101.480 76.430 101.740 ;
        RECT 78.960 101.725 79.100 101.880 ;
        RECT 78.885 101.495 79.175 101.725 ;
        RECT 79.345 101.680 79.635 101.725 ;
        RECT 79.790 101.680 80.110 101.740 ;
        RECT 79.345 101.540 80.110 101.680 ;
        RECT 79.345 101.495 79.635 101.540 ;
        RECT 79.790 101.480 80.110 101.540 ;
        RECT 80.250 101.480 80.570 101.740 ;
        RECT 80.725 101.495 81.015 101.725 ;
        RECT 82.090 101.680 82.410 101.740 ;
        RECT 83.100 101.725 83.240 101.880 ;
        RECT 83.930 101.820 84.250 101.880 ;
        RECT 82.565 101.680 82.855 101.725 ;
        RECT 82.090 101.540 82.855 101.680 ;
        RECT 80.800 101.340 80.940 101.495 ;
        RECT 82.090 101.480 82.410 101.540 ;
        RECT 82.565 101.495 82.855 101.540 ;
        RECT 83.025 101.495 83.315 101.725 ;
        RECT 83.470 101.480 83.790 101.740 ;
        RECT 84.390 101.480 84.710 101.740 ;
        RECT 85.860 101.725 86.000 102.220 ;
        RECT 85.785 101.680 86.075 101.725 ;
        RECT 87.150 101.680 87.470 101.740 ;
        RECT 85.785 101.540 87.470 101.680 ;
        RECT 85.785 101.495 86.075 101.540 ;
        RECT 87.150 101.480 87.470 101.540 ;
        RECT 87.625 101.680 87.915 101.725 ;
        RECT 88.070 101.680 88.390 101.740 ;
        RECT 87.625 101.540 88.390 101.680 ;
        RECT 87.625 101.495 87.915 101.540 ;
        RECT 88.070 101.480 88.390 101.540 ;
        RECT 85.310 101.340 85.630 101.400 ;
        RECT 86.230 101.340 86.550 101.400 ;
        RECT 80.800 101.200 85.080 101.340 ;
        RECT 55.410 100.860 64.380 101.000 ;
        RECT 55.410 100.800 55.730 100.860 ;
        RECT 60.010 100.800 60.330 100.860 ;
        RECT 60.930 100.800 61.250 100.860 ;
        RECT 65.070 100.800 65.390 101.060 ;
        RECT 72.890 101.000 73.210 101.060 ;
        RECT 84.940 101.045 85.080 101.200 ;
        RECT 85.310 101.200 86.550 101.340 ;
        RECT 85.310 101.140 85.630 101.200 ;
        RECT 86.230 101.140 86.550 101.200 ;
        RECT 86.690 101.140 87.010 101.400 ;
        RECT 106.195 101.085 107.455 102.975 ;
        RECT 119.900 102.760 120.990 105.420 ;
        RECT 122.340 104.370 125.190 105.490 ;
        RECT 125.580 105.190 125.930 105.940 ;
        RECT 126.680 105.820 128.550 105.980 ;
        RECT 126.680 105.770 127.440 105.820 ;
        RECT 128.320 105.750 128.550 105.820 ;
        RECT 136.960 105.750 137.190 105.980 ;
        RECT 128.755 105.470 136.755 105.700 ;
        RECT 125.580 105.130 125.870 105.190 ;
        RECT 125.490 105.010 125.870 105.130 ;
        RECT 128.850 105.070 136.710 105.470 ;
        RECT 137.520 105.070 138.480 114.550 ;
        RECT 139.930 116.780 140.700 120.420 ;
        RECT 142.370 119.370 145.220 120.490 ;
        RECT 145.610 120.190 145.960 120.940 ;
        RECT 146.710 120.820 148.580 120.980 ;
        RECT 146.710 120.770 147.470 120.820 ;
        RECT 148.350 120.750 148.580 120.820 ;
        RECT 156.990 120.750 157.220 120.980 ;
        RECT 148.785 120.470 156.785 120.700 ;
        RECT 145.610 120.130 145.900 120.190 ;
        RECT 145.520 120.010 145.900 120.130 ;
        RECT 148.880 120.070 156.740 120.470 ;
        RECT 157.550 120.070 158.510 129.550 ;
        RECT 142.310 119.140 145.310 119.370 ;
        RECT 145.520 119.180 145.860 120.010 ;
        RECT 147.870 120.000 158.510 120.070 ;
        RECT 142.360 119.110 145.220 119.140 ;
        RECT 142.360 119.090 143.530 119.110 ;
        RECT 144.490 119.100 145.220 119.110 ;
        RECT 142.310 118.700 145.310 118.930 ;
        RECT 145.515 118.890 145.860 119.180 ;
        RECT 146.050 118.960 158.510 120.000 ;
        RECT 146.050 118.940 158.500 118.960 ;
        RECT 145.520 118.780 145.860 118.890 ;
        RECT 146.090 118.930 151.760 118.940 ;
        RECT 152.760 118.930 158.500 118.940 ;
        RECT 142.400 118.530 145.260 118.700 ;
        RECT 146.090 118.530 146.520 118.930 ;
        RECT 142.370 118.160 146.520 118.530 ;
        RECT 139.930 114.680 140.790 116.780 ;
        RECT 146.460 116.390 147.710 116.830 ;
        RECT 157.640 116.810 158.500 118.930 ;
        RECT 144.400 116.380 149.640 116.390 ;
        RECT 141.450 116.280 156.750 116.380 ;
        RECT 141.450 116.270 156.785 116.280 ;
        RECT 141.410 116.150 156.785 116.270 ;
        RECT 141.410 116.040 145.410 116.150 ;
        RECT 146.460 116.070 148.200 116.150 ;
        RECT 148.780 116.070 156.785 116.150 ;
        RECT 146.460 115.990 147.710 116.070 ;
        RECT 148.785 116.050 156.785 116.070 ;
        RECT 141.020 115.740 141.250 115.990 ;
        RECT 145.570 115.850 145.800 115.990 ;
        RECT 148.350 115.850 148.580 116.000 ;
        RECT 145.570 115.740 148.580 115.850 ;
        RECT 156.990 115.740 157.220 116.000 ;
        RECT 141.020 115.300 157.220 115.740 ;
        RECT 141.020 115.030 141.250 115.300 ;
        RECT 145.570 115.270 157.220 115.300 ;
        RECT 145.570 115.180 148.580 115.270 ;
        RECT 145.570 115.030 145.800 115.180 ;
        RECT 148.350 115.040 148.580 115.180 ;
        RECT 156.990 115.040 157.220 115.270 ;
        RECT 141.410 114.750 145.410 114.980 ;
        RECT 148.785 114.770 156.785 114.990 ;
        RECT 157.550 114.770 158.510 116.810 ;
        RECT 148.785 114.760 158.510 114.770 ;
        RECT 141.410 114.680 145.400 114.750 ;
        RECT 139.930 114.570 145.400 114.680 ;
        RECT 148.840 114.600 158.510 114.760 ;
        RECT 139.930 114.480 143.090 114.570 ;
        RECT 156.580 114.550 158.510 114.600 ;
        RECT 139.930 111.210 140.790 114.480 ;
        RECT 144.440 114.020 149.690 114.030 ;
        RECT 144.440 113.910 156.750 114.020 ;
        RECT 141.470 113.850 156.750 113.910 ;
        RECT 141.470 113.840 156.785 113.850 ;
        RECT 141.410 113.710 156.785 113.840 ;
        RECT 141.410 113.700 146.570 113.710 ;
        RECT 141.410 113.610 145.410 113.700 ;
        RECT 148.785 113.620 156.785 113.710 ;
        RECT 148.870 113.610 156.760 113.620 ;
        RECT 141.020 113.250 141.250 113.560 ;
        RECT 141.470 113.250 145.370 113.610 ;
        RECT 145.570 113.250 145.800 113.560 ;
        RECT 141.020 111.910 145.800 113.250 ;
        RECT 141.020 111.600 141.250 111.910 ;
        RECT 145.570 111.600 145.800 111.910 ;
        RECT 148.350 113.030 148.580 113.570 ;
        RECT 149.390 113.030 150.400 113.060 ;
        RECT 156.990 113.030 157.220 113.570 ;
        RECT 148.350 112.130 157.220 113.030 ;
        RECT 148.350 111.610 148.580 112.130 ;
        RECT 149.390 112.060 150.400 112.130 ;
        RECT 156.990 111.610 157.220 112.130 ;
        RECT 141.410 111.320 145.410 111.550 ;
        RECT 148.785 111.330 156.785 111.560 ;
        RECT 139.930 111.170 141.090 111.210 ;
        RECT 139.930 111.090 141.330 111.170 ;
        RECT 141.700 111.100 145.360 111.320 ;
        RECT 141.700 111.090 143.140 111.100 ;
        RECT 139.930 111.050 143.140 111.090 ;
        RECT 139.930 110.960 142.650 111.050 ;
        RECT 148.850 111.040 156.740 111.330 ;
        RECT 139.930 110.900 141.980 110.960 ;
        RECT 139.930 110.850 141.730 110.900 ;
        RECT 139.930 107.510 140.790 110.850 ;
        RECT 148.840 110.550 156.760 110.560 ;
        RECT 145.070 110.540 156.760 110.550 ;
        RECT 141.450 110.420 156.760 110.540 ;
        RECT 141.450 110.410 156.785 110.420 ;
        RECT 141.410 110.290 156.785 110.410 ;
        RECT 141.410 110.180 145.410 110.290 ;
        RECT 141.020 109.840 141.250 110.130 ;
        RECT 141.470 109.840 145.360 110.180 ;
        RECT 145.570 109.840 145.800 110.130 ;
        RECT 141.020 108.470 145.800 109.840 ;
        RECT 141.020 108.170 141.250 108.470 ;
        RECT 145.570 108.170 145.800 108.470 ;
        RECT 141.410 107.890 145.410 108.120 ;
        RECT 141.660 107.660 145.230 107.890 ;
        RECT 141.660 107.510 145.350 107.660 ;
        RECT 139.930 107.230 145.350 107.510 ;
        RECT 146.600 107.340 147.220 110.290 ;
        RECT 148.785 110.190 156.785 110.290 ;
        RECT 148.840 110.180 156.760 110.190 ;
        RECT 148.350 109.480 148.580 110.140 ;
        RECT 149.360 109.480 150.360 109.570 ;
        RECT 156.990 109.480 157.220 110.140 ;
        RECT 148.350 108.660 157.220 109.480 ;
        RECT 148.350 108.180 148.580 108.660 ;
        RECT 149.360 108.570 150.360 108.660 ;
        RECT 156.990 108.180 157.220 108.660 ;
        RECT 148.785 107.900 156.785 108.130 ;
        RECT 139.930 106.770 145.360 107.230 ;
        RECT 139.930 106.630 141.960 106.770 ;
        RECT 139.960 105.430 141.960 106.630 ;
        RECT 143.710 106.760 145.360 106.770 ;
        RECT 142.400 105.490 143.400 106.210 ;
        RECT 143.710 105.950 144.020 106.760 ;
        RECT 144.480 106.480 145.360 106.760 ;
        RECT 145.600 106.940 147.220 107.340 ;
        RECT 148.870 106.990 156.740 107.900 ;
        RECT 144.420 106.250 145.420 106.480 ;
        RECT 145.600 106.290 145.950 106.940 ;
        RECT 146.600 106.930 147.220 106.940 ;
        RECT 148.785 106.760 156.785 106.990 ;
        RECT 148.870 106.750 156.740 106.760 ;
        RECT 144.480 106.040 145.360 106.060 ;
        RECT 143.750 105.660 144.020 105.950 ;
        RECT 144.420 105.810 145.420 106.040 ;
        RECT 145.580 106.000 145.950 106.290 ;
        RECT 145.610 105.940 145.950 106.000 ;
        RECT 146.710 106.610 147.470 106.660 ;
        RECT 148.350 106.610 148.580 106.710 ;
        RECT 146.710 106.400 148.580 106.610 ;
        RECT 156.990 106.400 157.220 106.710 ;
        RECT 146.710 105.980 149.250 106.400 ;
        RECT 156.620 105.980 157.220 106.400 ;
        RECT 144.480 105.660 145.360 105.810 ;
        RECT 144.490 105.490 145.220 105.660 ;
        RECT 140.040 105.420 141.960 105.430 ;
        RECT 122.280 104.140 125.280 104.370 ;
        RECT 125.490 104.180 125.830 105.010 ;
        RECT 127.840 105.000 138.480 105.070 ;
        RECT 122.330 104.110 125.190 104.140 ;
        RECT 122.330 104.090 123.500 104.110 ;
        RECT 124.460 104.100 125.190 104.110 ;
        RECT 122.280 103.700 125.280 103.930 ;
        RECT 125.485 103.890 125.830 104.180 ;
        RECT 126.020 103.960 138.480 105.000 ;
        RECT 142.370 104.370 145.220 105.490 ;
        RECT 145.610 105.190 145.960 105.940 ;
        RECT 146.710 105.820 148.580 105.980 ;
        RECT 146.710 105.770 147.470 105.820 ;
        RECT 148.350 105.750 148.580 105.820 ;
        RECT 156.990 105.750 157.220 105.980 ;
        RECT 148.785 105.470 156.785 105.700 ;
        RECT 145.610 105.130 145.900 105.190 ;
        RECT 145.520 105.010 145.900 105.130 ;
        RECT 148.880 105.070 156.740 105.470 ;
        RECT 157.550 105.070 158.510 114.550 ;
        RECT 142.310 104.140 145.310 104.370 ;
        RECT 145.520 104.180 145.860 105.010 ;
        RECT 147.870 105.000 158.510 105.070 ;
        RECT 142.360 104.110 145.220 104.140 ;
        RECT 142.360 104.090 143.530 104.110 ;
        RECT 144.490 104.100 145.220 104.110 ;
        RECT 126.020 103.940 138.350 103.960 ;
        RECT 125.490 103.780 125.830 103.890 ;
        RECT 126.060 103.930 131.730 103.940 ;
        RECT 132.730 103.930 138.350 103.940 ;
        RECT 122.370 103.530 125.230 103.700 ;
        RECT 126.060 103.530 126.490 103.930 ;
        RECT 142.310 103.700 145.310 103.930 ;
        RECT 145.515 103.890 145.860 104.180 ;
        RECT 146.050 103.960 158.510 105.000 ;
        RECT 146.050 103.940 158.460 103.960 ;
        RECT 145.520 103.780 145.860 103.890 ;
        RECT 146.090 103.930 151.760 103.940 ;
        RECT 152.760 103.930 158.460 103.940 ;
        RECT 142.400 103.530 145.260 103.700 ;
        RECT 146.090 103.530 146.520 103.930 ;
        RECT 122.340 103.160 126.490 103.530 ;
        RECT 142.370 103.160 146.520 103.530 ;
        RECT 113.040 102.695 116.730 102.710 ;
        RECT 119.900 102.695 135.450 102.760 ;
        RECT 113.040 101.710 135.450 102.695 ;
        RECT 113.040 101.690 132.370 101.710 ;
        RECT 113.040 101.675 123.360 101.690 ;
        RECT 113.040 101.660 116.730 101.675 ;
        RECT 99.990 101.065 112.800 101.085 ;
        RECT 75.205 101.000 75.495 101.045 ;
        RECT 72.890 100.860 75.495 101.000 ;
        RECT 72.890 100.800 73.210 100.860 ;
        RECT 75.205 100.815 75.495 100.860 ;
        RECT 84.865 100.815 85.155 101.045 ;
        RECT 12.100 100.180 89.840 100.660 ;
        RECT 99.970 100.255 112.810 101.065 ;
        RECT 99.990 100.195 112.800 100.255 ;
        RECT 26.430 99.980 26.750 100.040 ;
        RECT 39.325 99.980 39.615 100.025 ;
        RECT 46.210 99.980 46.530 100.040 ;
        RECT 26.430 99.840 32.640 99.980 ;
        RECT 26.430 99.780 26.750 99.840 ;
        RECT 22.750 99.640 23.070 99.700 ;
        RECT 25.510 99.640 25.830 99.700 ;
        RECT 25.985 99.640 26.275 99.685 ;
        RECT 22.750 99.500 26.275 99.640 ;
        RECT 22.750 99.440 23.070 99.500 ;
        RECT 25.510 99.440 25.830 99.500 ;
        RECT 25.985 99.455 26.275 99.500 ;
        RECT 27.350 99.640 27.670 99.700 ;
        RECT 27.350 99.500 30.800 99.640 ;
        RECT 27.350 99.440 27.670 99.500 ;
        RECT 18.165 99.300 18.455 99.345 ;
        RECT 18.610 99.300 18.930 99.360 ;
        RECT 18.165 99.160 18.930 99.300 ;
        RECT 18.165 99.115 18.455 99.160 ;
        RECT 18.610 99.100 18.930 99.160 ;
        RECT 19.085 99.300 19.375 99.345 ;
        RECT 21.830 99.300 22.150 99.360 ;
        RECT 30.660 99.345 30.800 99.500 ;
        RECT 32.500 99.360 32.640 99.840 ;
        RECT 39.325 99.840 46.530 99.980 ;
        RECT 39.325 99.795 39.615 99.840 ;
        RECT 46.210 99.780 46.530 99.840 ;
        RECT 48.970 99.980 49.290 100.040 ;
        RECT 52.190 99.980 52.510 100.040 ;
        RECT 48.970 99.840 55.640 99.980 ;
        RECT 48.970 99.780 49.290 99.840 ;
        RECT 52.190 99.780 52.510 99.840 ;
        RECT 41.610 99.640 41.930 99.700 ;
        RECT 43.450 99.685 43.770 99.700 ;
        RECT 40.780 99.500 41.930 99.640 ;
        RECT 19.085 99.160 22.150 99.300 ;
        RECT 19.085 99.115 19.375 99.160 ;
        RECT 21.830 99.100 22.150 99.160 ;
        RECT 30.585 99.300 30.875 99.345 ;
        RECT 31.490 99.300 31.810 99.360 ;
        RECT 30.585 99.160 31.810 99.300 ;
        RECT 30.585 99.115 30.875 99.160 ;
        RECT 31.490 99.100 31.810 99.160 ;
        RECT 32.410 99.300 32.730 99.360 ;
        RECT 34.265 99.300 34.555 99.345 ;
        RECT 32.410 99.160 34.555 99.300 ;
        RECT 32.410 99.100 32.730 99.160 ;
        RECT 34.265 99.115 34.555 99.160 ;
        RECT 36.550 99.300 36.870 99.360 ;
        RECT 38.405 99.300 38.695 99.345 ;
        RECT 36.550 99.160 38.695 99.300 ;
        RECT 36.550 99.100 36.870 99.160 ;
        RECT 38.405 99.115 38.695 99.160 ;
        RECT 39.325 99.300 39.615 99.345 ;
        RECT 39.770 99.300 40.090 99.360 ;
        RECT 40.780 99.345 40.920 99.500 ;
        RECT 41.610 99.440 41.930 99.500 ;
        RECT 43.420 99.455 43.770 99.685 ;
        RECT 43.450 99.440 43.770 99.455 ;
        RECT 48.510 99.640 48.830 99.700 ;
        RECT 49.445 99.640 49.735 99.685 ;
        RECT 54.490 99.640 54.810 99.700 ;
        RECT 55.500 99.685 55.640 99.840 ;
        RECT 57.250 99.780 57.570 100.040 ;
        RECT 59.090 99.980 59.410 100.040 ;
        RECT 61.405 99.980 61.695 100.025 ;
        RECT 59.090 99.840 61.695 99.980 ;
        RECT 59.090 99.780 59.410 99.840 ;
        RECT 61.405 99.795 61.695 99.840 ;
        RECT 63.245 99.980 63.535 100.025 ;
        RECT 76.110 99.980 76.430 100.040 ;
        RECT 63.245 99.840 76.430 99.980 ;
        RECT 63.245 99.795 63.535 99.840 ;
        RECT 76.110 99.780 76.430 99.840 ;
        RECT 77.490 99.780 77.810 100.040 ;
        RECT 83.470 99.980 83.790 100.040 ;
        RECT 88.085 99.980 88.375 100.025 ;
        RECT 83.470 99.840 88.375 99.980 ;
        RECT 83.470 99.780 83.790 99.840 ;
        RECT 88.085 99.795 88.375 99.840 ;
        RECT 100.990 99.835 101.430 100.195 ;
        RECT 102.570 100.085 103.730 100.195 ;
        RECT 102.570 99.835 103.010 100.085 ;
        RECT 104.160 99.835 104.600 100.195 ;
        RECT 105.750 99.835 106.190 100.195 ;
        RECT 100.130 99.785 100.360 99.815 ;
        RECT 100.520 99.785 100.750 99.835 ;
        RECT 48.510 99.500 54.810 99.640 ;
        RECT 48.510 99.440 48.830 99.500 ;
        RECT 49.445 99.455 49.735 99.500 ;
        RECT 54.490 99.440 54.810 99.500 ;
        RECT 55.425 99.455 55.715 99.685 ;
        RECT 56.505 99.640 56.795 99.685 ;
        RECT 58.170 99.640 58.490 99.700 ;
        RECT 67.830 99.640 68.150 99.700 ;
        RECT 85.310 99.640 85.630 99.700 ;
        RECT 87.165 99.640 87.455 99.685 ;
        RECT 56.505 99.500 61.160 99.640 ;
        RECT 56.505 99.455 56.795 99.500 ;
        RECT 58.170 99.440 58.490 99.500 ;
        RECT 39.325 99.160 40.090 99.300 ;
        RECT 39.325 99.115 39.615 99.160 ;
        RECT 29.665 98.960 29.955 99.005 ;
        RECT 34.725 98.960 35.015 99.005 ;
        RECT 29.665 98.820 35.015 98.960 ;
        RECT 38.480 98.960 38.620 99.115 ;
        RECT 39.770 99.100 40.090 99.160 ;
        RECT 40.705 99.115 40.995 99.345 ;
        RECT 41.150 99.300 41.470 99.360 ;
        RECT 42.085 99.300 42.375 99.345 ;
        RECT 45.290 99.300 45.610 99.360 ;
        RECT 41.150 99.160 42.375 99.300 ;
        RECT 41.150 99.100 41.470 99.160 ;
        RECT 42.085 99.115 42.375 99.160 ;
        RECT 42.620 99.290 43.680 99.300 ;
        RECT 44.000 99.290 51.040 99.300 ;
        RECT 42.620 99.160 51.040 99.290 ;
        RECT 42.620 98.960 42.760 99.160 ;
        RECT 43.540 99.150 44.140 99.160 ;
        RECT 45.290 99.100 45.610 99.160 ;
        RECT 38.480 98.820 42.760 98.960 ;
        RECT 42.965 98.960 43.255 99.005 ;
        RECT 44.155 98.960 44.445 99.005 ;
        RECT 46.675 98.960 46.965 99.005 ;
        RECT 42.965 98.820 46.965 98.960 ;
        RECT 29.665 98.775 29.955 98.820 ;
        RECT 34.725 98.775 35.015 98.820 ;
        RECT 42.965 98.775 43.255 98.820 ;
        RECT 44.155 98.775 44.445 98.820 ;
        RECT 46.675 98.775 46.965 98.820 ;
        RECT 42.570 98.620 42.860 98.665 ;
        RECT 44.670 98.620 44.960 98.665 ;
        RECT 46.240 98.620 46.530 98.665 ;
        RECT 50.350 98.620 50.670 98.680 ;
        RECT 50.900 98.665 51.040 99.160 ;
        RECT 53.585 99.115 53.875 99.345 ;
        RECT 54.045 99.300 54.335 99.345 ;
        RECT 54.950 99.300 55.270 99.360 ;
        RECT 54.045 99.160 55.270 99.300 ;
        RECT 54.045 99.115 54.335 99.160 ;
        RECT 53.660 98.960 53.800 99.115 ;
        RECT 54.950 99.100 55.270 99.160 ;
        RECT 55.870 99.100 56.190 99.360 ;
        RECT 57.725 99.300 58.015 99.345 ;
        RECT 56.420 99.160 58.015 99.300 ;
        RECT 55.960 98.960 56.100 99.100 ;
        RECT 53.660 98.820 56.100 98.960 ;
        RECT 42.570 98.480 46.530 98.620 ;
        RECT 42.570 98.435 42.860 98.480 ;
        RECT 44.670 98.435 44.960 98.480 ;
        RECT 46.240 98.435 46.530 98.480 ;
        RECT 48.600 98.480 50.670 98.620 ;
        RECT 17.230 98.280 17.550 98.340 ;
        RECT 18.165 98.280 18.455 98.325 ;
        RECT 17.230 98.140 18.455 98.280 ;
        RECT 17.230 98.080 17.550 98.140 ;
        RECT 18.165 98.095 18.455 98.140 ;
        RECT 40.245 98.280 40.535 98.325 ;
        RECT 48.600 98.280 48.740 98.480 ;
        RECT 50.350 98.420 50.670 98.480 ;
        RECT 50.825 98.435 51.115 98.665 ;
        RECT 51.745 98.620 52.035 98.665 ;
        RECT 55.870 98.620 56.190 98.680 ;
        RECT 51.745 98.480 56.190 98.620 ;
        RECT 51.745 98.435 52.035 98.480 ;
        RECT 55.870 98.420 56.190 98.480 ;
        RECT 40.245 98.140 48.740 98.280 ;
        RECT 40.245 98.095 40.535 98.140 ;
        RECT 53.570 98.080 53.890 98.340 ;
        RECT 54.490 98.280 54.810 98.340 ;
        RECT 56.420 98.325 56.560 99.160 ;
        RECT 57.725 99.115 58.015 99.160 ;
        RECT 58.645 99.115 58.935 99.345 ;
        RECT 58.720 98.960 58.860 99.115 ;
        RECT 59.550 99.100 59.870 99.360 ;
        RECT 61.020 99.345 61.160 99.500 ;
        RECT 66.080 99.500 68.750 99.640 ;
        RECT 60.945 99.115 61.235 99.345 ;
        RECT 62.325 99.300 62.615 99.345 ;
        RECT 64.150 99.300 64.470 99.360 ;
        RECT 66.080 99.345 66.220 99.500 ;
        RECT 67.830 99.440 68.150 99.500 ;
        RECT 67.370 99.345 67.690 99.360 ;
        RECT 62.325 99.160 64.470 99.300 ;
        RECT 62.325 99.115 62.615 99.160 ;
        RECT 64.150 99.100 64.470 99.160 ;
        RECT 66.005 99.115 66.295 99.345 ;
        RECT 67.340 99.115 67.690 99.345 ;
        RECT 68.610 99.300 68.750 99.500 ;
        RECT 78.500 99.500 87.455 99.640 ;
        RECT 77.950 99.300 78.270 99.360 ;
        RECT 78.500 99.345 78.640 99.500 ;
        RECT 85.310 99.440 85.630 99.500 ;
        RECT 87.165 99.455 87.455 99.500 ;
        RECT 68.610 99.160 78.270 99.300 ;
        RECT 67.370 99.100 67.690 99.115 ;
        RECT 77.950 99.100 78.270 99.160 ;
        RECT 78.425 99.115 78.715 99.345 ;
        RECT 79.330 99.300 79.650 99.360 ;
        RECT 80.165 99.300 80.455 99.345 ;
        RECT 79.330 99.160 80.455 99.300 ;
        RECT 79.330 99.100 79.650 99.160 ;
        RECT 80.165 99.115 80.455 99.160 ;
        RECT 84.850 99.300 85.170 99.360 ;
        RECT 85.770 99.300 86.090 99.360 ;
        RECT 86.245 99.300 86.535 99.345 ;
        RECT 84.850 99.160 86.535 99.300 ;
        RECT 84.850 99.100 85.170 99.160 ;
        RECT 85.770 99.100 86.090 99.160 ;
        RECT 86.245 99.115 86.535 99.160 ;
        RECT 60.010 98.960 60.330 99.020 ;
        RECT 58.720 98.820 60.330 98.960 ;
        RECT 60.010 98.760 60.330 98.820 ;
        RECT 66.885 98.960 67.175 99.005 ;
        RECT 68.075 98.960 68.365 99.005 ;
        RECT 70.595 98.960 70.885 99.005 ;
        RECT 66.885 98.820 70.885 98.960 ;
        RECT 66.885 98.775 67.175 98.820 ;
        RECT 68.075 98.775 68.365 98.820 ;
        RECT 70.595 98.775 70.885 98.820 ;
        RECT 76.125 98.775 76.415 99.005 ;
        RECT 78.040 98.960 78.180 99.100 ;
        RECT 78.885 98.960 79.175 99.005 ;
        RECT 78.040 98.820 79.175 98.960 ;
        RECT 78.885 98.775 79.175 98.820 ;
        RECT 79.765 98.960 80.055 99.005 ;
        RECT 80.955 98.960 81.245 99.005 ;
        RECT 83.475 98.960 83.765 99.005 ;
        RECT 79.765 98.820 83.765 98.960 ;
        RECT 79.765 98.775 80.055 98.820 ;
        RECT 80.955 98.775 81.245 98.820 ;
        RECT 83.475 98.775 83.765 98.820 ;
        RECT 66.490 98.620 66.780 98.665 ;
        RECT 68.590 98.620 68.880 98.665 ;
        RECT 70.160 98.620 70.450 98.665 ;
        RECT 66.490 98.480 70.450 98.620 ;
        RECT 66.490 98.435 66.780 98.480 ;
        RECT 68.590 98.435 68.880 98.480 ;
        RECT 70.160 98.435 70.450 98.480 ;
        RECT 72.905 98.620 73.195 98.665 ;
        RECT 76.200 98.620 76.340 98.775 ;
        RECT 77.030 98.620 77.350 98.680 ;
        RECT 72.905 98.480 77.350 98.620 ;
        RECT 72.905 98.435 73.195 98.480 ;
        RECT 77.030 98.420 77.350 98.480 ;
        RECT 79.370 98.620 79.660 98.665 ;
        RECT 81.470 98.620 81.760 98.665 ;
        RECT 83.040 98.620 83.330 98.665 ;
        RECT 79.370 98.480 83.330 98.620 ;
        RECT 79.370 98.435 79.660 98.480 ;
        RECT 81.470 98.435 81.760 98.480 ;
        RECT 83.040 98.435 83.330 98.480 ;
        RECT 56.345 98.280 56.635 98.325 ;
        RECT 54.490 98.140 56.635 98.280 ;
        RECT 54.490 98.080 54.810 98.140 ;
        RECT 56.345 98.095 56.635 98.140 ;
        RECT 59.550 98.280 59.870 98.340 ;
        RECT 61.390 98.280 61.710 98.340 ;
        RECT 59.550 98.140 61.710 98.280 ;
        RECT 59.550 98.080 59.870 98.140 ;
        RECT 61.390 98.080 61.710 98.140 ;
        RECT 73.350 98.080 73.670 98.340 ;
        RECT 83.470 98.280 83.790 98.340 ;
        RECT 85.785 98.280 86.075 98.325 ;
        RECT 83.470 98.140 86.075 98.280 ;
        RECT 83.470 98.080 83.790 98.140 ;
        RECT 85.785 98.095 86.075 98.140 ;
        RECT 12.100 97.460 89.840 97.940 ;
        RECT 14.485 97.260 14.775 97.305 ;
        RECT 16.310 97.260 16.630 97.320 ;
        RECT 14.485 97.120 16.630 97.260 ;
        RECT 14.485 97.075 14.775 97.120 ;
        RECT 16.310 97.060 16.630 97.120 ;
        RECT 16.785 97.260 17.075 97.305 ;
        RECT 20.910 97.260 21.230 97.320 ;
        RECT 16.785 97.120 21.230 97.260 ;
        RECT 16.785 97.075 17.075 97.120 ;
        RECT 20.910 97.060 21.230 97.120 ;
        RECT 23.210 97.260 23.530 97.320 ;
        RECT 24.145 97.260 24.435 97.305 ;
        RECT 23.210 97.120 24.435 97.260 ;
        RECT 23.210 97.060 23.530 97.120 ;
        RECT 24.145 97.075 24.435 97.120 ;
        RECT 29.205 97.260 29.495 97.305 ;
        RECT 29.650 97.260 29.970 97.320 ;
        RECT 29.205 97.120 29.970 97.260 ;
        RECT 29.205 97.075 29.495 97.120 ;
        RECT 29.650 97.060 29.970 97.120 ;
        RECT 33.330 97.060 33.650 97.320 ;
        RECT 43.005 97.260 43.295 97.305 ;
        RECT 43.450 97.260 43.770 97.320 ;
        RECT 43.005 97.120 43.770 97.260 ;
        RECT 43.005 97.075 43.295 97.120 ;
        RECT 43.450 97.060 43.770 97.120 ;
        RECT 44.370 97.060 44.690 97.320 ;
        RECT 57.710 97.060 58.030 97.320 ;
        RECT 67.370 97.260 67.690 97.320 ;
        RECT 67.845 97.260 68.135 97.305 ;
        RECT 67.370 97.120 68.135 97.260 ;
        RECT 67.370 97.060 67.690 97.120 ;
        RECT 67.845 97.075 68.135 97.120 ;
        RECT 68.290 97.260 68.610 97.320 ;
        RECT 78.425 97.260 78.715 97.305 ;
        RECT 79.330 97.260 79.650 97.320 ;
        RECT 82.090 97.260 82.410 97.320 ;
        RECT 68.290 97.120 74.960 97.260 ;
        RECT 68.290 97.060 68.610 97.120 ;
        RECT 20.465 96.920 20.755 96.965 ;
        RECT 21.370 96.920 21.690 96.980 ;
        RECT 25.510 96.920 25.830 96.980 ;
        RECT 20.465 96.780 25.830 96.920 ;
        RECT 20.465 96.735 20.755 96.780 ;
        RECT 21.370 96.720 21.690 96.780 ;
        RECT 25.510 96.720 25.830 96.780 ;
        RECT 49.445 96.920 49.735 96.965 ;
        RECT 50.350 96.920 50.670 96.980 ;
        RECT 49.445 96.780 50.670 96.920 ;
        RECT 74.820 96.920 74.960 97.120 ;
        RECT 78.425 97.120 79.650 97.260 ;
        RECT 78.425 97.075 78.715 97.120 ;
        RECT 79.330 97.060 79.650 97.120 ;
        RECT 79.880 97.120 82.410 97.260 ;
        RECT 74.820 96.780 75.420 96.920 ;
        RECT 49.445 96.735 49.735 96.780 ;
        RECT 50.350 96.720 50.670 96.780 ;
        RECT 7.110 96.580 7.430 96.640 ;
        RECT 65.070 96.580 65.390 96.640 ;
        RECT 70.605 96.580 70.895 96.625 ;
        RECT 7.110 96.440 51.500 96.580 ;
        RECT 7.110 96.380 7.430 96.440 ;
        RECT 18.610 96.040 18.930 96.300 ;
        RECT 19.545 96.250 19.835 96.285 ;
        RECT 19.260 96.110 19.835 96.250 ;
        RECT 15.390 95.700 15.710 95.960 ;
        RECT 17.705 95.900 17.995 95.945 ;
        RECT 18.150 95.900 18.470 95.960 ;
        RECT 17.705 95.760 18.470 95.900 ;
        RECT 19.260 95.900 19.400 96.110 ;
        RECT 19.545 96.055 19.835 96.110 ;
        RECT 19.990 96.040 20.310 96.300 ;
        RECT 21.830 96.240 22.150 96.300 ;
        RECT 22.320 96.240 22.610 96.285 ;
        RECT 21.830 96.100 22.610 96.240 ;
        RECT 21.830 96.040 22.150 96.100 ;
        RECT 22.320 96.055 22.610 96.100 ;
        RECT 23.210 96.040 23.530 96.300 ;
        RECT 23.670 96.040 23.990 96.300 ;
        RECT 24.605 96.055 24.895 96.285 ;
        RECT 23.300 95.900 23.440 96.040 ;
        RECT 19.260 95.760 23.440 95.900 ;
        RECT 24.130 95.900 24.450 95.960 ;
        RECT 24.680 95.900 24.820 96.055 ;
        RECT 25.510 96.040 25.830 96.300 ;
        RECT 25.970 96.040 26.290 96.300 ;
        RECT 30.125 96.240 30.415 96.285 ;
        RECT 31.490 96.240 31.810 96.300 ;
        RECT 30.125 96.100 31.810 96.240 ;
        RECT 30.125 96.055 30.415 96.100 ;
        RECT 31.490 96.040 31.810 96.100 ;
        RECT 32.410 96.040 32.730 96.300 ;
        RECT 32.890 96.055 33.180 96.285 ;
        RECT 43.005 96.055 43.295 96.285 ;
        RECT 43.925 96.240 44.215 96.285 ;
        RECT 45.305 96.240 45.595 96.285 ;
        RECT 43.925 96.100 45.595 96.240 ;
        RECT 43.925 96.055 44.215 96.100 ;
        RECT 45.305 96.055 45.595 96.100 ;
        RECT 26.890 95.900 27.210 95.960 ;
        RECT 24.130 95.760 27.210 95.900 ;
        RECT 17.705 95.715 17.995 95.760 ;
        RECT 18.150 95.700 18.470 95.760 ;
        RECT 24.130 95.700 24.450 95.760 ;
        RECT 26.890 95.700 27.210 95.760 ;
        RECT 31.045 95.715 31.335 95.945 ;
        RECT 31.580 95.900 31.720 96.040 ;
        RECT 32.960 95.900 33.100 96.055 ;
        RECT 31.580 95.760 33.100 95.900 ;
        RECT 13.550 95.360 13.870 95.620 ;
        RECT 14.470 95.605 14.790 95.620 ;
        RECT 14.405 95.375 14.790 95.605 ;
        RECT 14.470 95.360 14.790 95.375 ;
        RECT 15.850 95.360 16.170 95.620 ;
        RECT 16.705 95.560 16.995 95.605 ;
        RECT 18.610 95.560 18.930 95.620 ;
        RECT 16.705 95.420 18.930 95.560 ;
        RECT 16.705 95.375 16.995 95.420 ;
        RECT 18.610 95.360 18.930 95.420 ;
        RECT 19.070 95.360 19.390 95.620 ;
        RECT 22.290 95.360 22.610 95.620 ;
        RECT 23.225 95.560 23.515 95.605 ;
        RECT 23.670 95.560 23.990 95.620 ;
        RECT 23.225 95.420 23.990 95.560 ;
        RECT 31.120 95.560 31.260 95.715 ;
        RECT 32.410 95.560 32.730 95.620 ;
        RECT 37.010 95.560 37.330 95.620 ;
        RECT 31.120 95.420 37.330 95.560 ;
        RECT 43.080 95.560 43.220 96.055 ;
        RECT 45.380 95.900 45.520 96.055 ;
        RECT 45.750 96.040 46.070 96.300 ;
        RECT 46.210 96.040 46.530 96.300 ;
        RECT 47.145 96.240 47.435 96.285 ;
        RECT 48.050 96.240 48.370 96.300 ;
        RECT 47.145 96.100 48.370 96.240 ;
        RECT 47.145 96.055 47.435 96.100 ;
        RECT 48.050 96.040 48.370 96.100 ;
        RECT 48.510 96.040 48.830 96.300 ;
        RECT 49.890 96.040 50.210 96.300 ;
        RECT 51.360 96.285 51.500 96.440 ;
        RECT 65.070 96.440 70.895 96.580 ;
        RECT 65.070 96.380 65.390 96.440 ;
        RECT 70.605 96.395 70.895 96.440 ;
        RECT 51.285 96.055 51.575 96.285 ;
        RECT 69.685 96.240 69.975 96.285 ;
        RECT 73.350 96.240 73.670 96.300 ;
        RECT 69.685 96.100 73.670 96.240 ;
        RECT 69.685 96.055 69.975 96.100 ;
        RECT 73.350 96.040 73.670 96.100 ;
        RECT 74.285 96.055 74.575 96.285 ;
        RECT 50.810 95.900 51.130 95.960 ;
        RECT 45.380 95.760 51.130 95.900 ;
        RECT 50.810 95.700 51.130 95.760 ;
        RECT 71.050 95.900 71.370 95.960 ;
        RECT 74.360 95.900 74.500 96.055 ;
        RECT 74.730 96.040 75.050 96.300 ;
        RECT 75.280 96.285 75.420 96.780 ;
        RECT 75.205 96.055 75.495 96.285 ;
        RECT 76.110 96.040 76.430 96.300 ;
        RECT 77.030 96.040 77.350 96.300 ;
        RECT 77.950 96.240 78.270 96.300 ;
        RECT 79.880 96.285 80.020 97.120 ;
        RECT 82.090 97.060 82.410 97.120 ;
        RECT 80.710 96.920 81.030 96.980 ;
        RECT 80.340 96.780 81.030 96.920 ;
        RECT 80.340 96.285 80.480 96.780 ;
        RECT 80.710 96.720 81.030 96.780 ;
        RECT 82.105 96.580 82.395 96.625 ;
        RECT 84.390 96.580 84.710 96.640 ;
        RECT 87.610 96.580 87.930 96.640 ;
        RECT 80.800 96.440 82.395 96.580 ;
        RECT 80.800 96.285 80.940 96.440 ;
        RECT 82.105 96.395 82.395 96.440 ;
        RECT 84.020 96.440 87.930 96.580 ;
        RECT 79.805 96.240 80.095 96.285 ;
        RECT 77.950 96.100 80.095 96.240 ;
        RECT 77.950 96.040 78.270 96.100 ;
        RECT 79.805 96.055 80.095 96.100 ;
        RECT 80.265 96.055 80.555 96.285 ;
        RECT 80.725 96.055 81.015 96.285 ;
        RECT 81.170 96.240 81.490 96.300 ;
        RECT 84.020 96.285 84.160 96.440 ;
        RECT 84.390 96.380 84.710 96.440 ;
        RECT 87.610 96.380 87.930 96.440 ;
        RECT 81.645 96.240 81.935 96.285 ;
        RECT 81.170 96.100 81.935 96.240 ;
        RECT 81.170 96.040 81.490 96.100 ;
        RECT 81.645 96.055 81.935 96.100 ;
        RECT 83.945 96.055 84.235 96.285 ;
        RECT 88.070 96.040 88.390 96.300 ;
        RECT 71.050 95.760 74.500 95.900 ;
        RECT 71.050 95.700 71.370 95.760 ;
        RECT 83.010 95.700 83.330 95.960 ;
        RECT 84.405 95.900 84.695 95.945 ;
        RECT 84.850 95.900 85.170 95.960 ;
        RECT 84.405 95.760 85.170 95.900 ;
        RECT 84.405 95.715 84.695 95.760 ;
        RECT 84.850 95.700 85.170 95.760 ;
        RECT 85.325 95.900 85.615 95.945 ;
        RECT 85.770 95.900 86.090 95.960 ;
        RECT 85.325 95.760 86.090 95.900 ;
        RECT 85.325 95.715 85.615 95.760 ;
        RECT 85.770 95.700 86.090 95.760 ;
        RECT 47.605 95.560 47.895 95.605 ;
        RECT 43.080 95.420 47.895 95.560 ;
        RECT 23.225 95.375 23.515 95.420 ;
        RECT 23.670 95.360 23.990 95.420 ;
        RECT 32.410 95.360 32.730 95.420 ;
        RECT 37.010 95.360 37.330 95.420 ;
        RECT 47.605 95.375 47.895 95.420 ;
        RECT 70.145 95.560 70.435 95.605 ;
        RECT 73.365 95.560 73.655 95.605 ;
        RECT 70.145 95.420 73.655 95.560 ;
        RECT 70.145 95.375 70.435 95.420 ;
        RECT 73.365 95.375 73.655 95.420 ;
        RECT 77.965 95.560 78.255 95.605 ;
        RECT 81.630 95.560 81.950 95.620 ;
        RECT 77.965 95.420 81.950 95.560 ;
        RECT 77.965 95.375 78.255 95.420 ;
        RECT 81.630 95.360 81.950 95.420 ;
        RECT 86.245 95.560 86.535 95.605 ;
        RECT 86.690 95.560 87.010 95.620 ;
        RECT 86.245 95.420 87.010 95.560 ;
        RECT 86.245 95.375 86.535 95.420 ;
        RECT 86.690 95.360 87.010 95.420 ;
        RECT 87.165 95.560 87.455 95.605 ;
        RECT 88.070 95.560 88.390 95.620 ;
        RECT 87.165 95.420 88.390 95.560 ;
        RECT 87.165 95.375 87.455 95.420 ;
        RECT 88.070 95.360 88.390 95.420 ;
        RECT 12.100 94.740 89.840 95.220 ;
        RECT 21.370 94.340 21.690 94.600 ;
        RECT 48.510 94.540 48.830 94.600 ;
        RECT 51.270 94.540 51.590 94.600 ;
        RECT 51.745 94.540 52.035 94.585 ;
        RECT 48.510 94.400 52.035 94.540 ;
        RECT 48.510 94.340 48.830 94.400 ;
        RECT 31.950 94.200 32.270 94.260 ;
        RECT 33.330 94.245 33.650 94.260 ;
        RECT 14.560 94.060 20.450 94.200 ;
        RECT 13.550 93.860 13.870 93.920 ;
        RECT 14.560 93.905 14.700 94.060 ;
        RECT 15.850 93.905 16.170 93.920 ;
        RECT 14.485 93.860 14.775 93.905 ;
        RECT 15.820 93.860 16.170 93.905 ;
        RECT 13.550 93.720 14.775 93.860 ;
        RECT 15.655 93.720 16.170 93.860 ;
        RECT 13.550 93.660 13.870 93.720 ;
        RECT 14.485 93.675 14.775 93.720 ;
        RECT 15.820 93.675 16.170 93.720 ;
        RECT 15.850 93.660 16.170 93.675 ;
        RECT 15.365 93.520 15.655 93.565 ;
        RECT 16.555 93.520 16.845 93.565 ;
        RECT 19.075 93.520 19.365 93.565 ;
        RECT 15.365 93.380 19.365 93.520 ;
        RECT 20.310 93.520 20.450 94.060 ;
        RECT 22.840 94.060 32.270 94.200 ;
        RECT 22.290 93.660 22.610 93.920 ;
        RECT 22.840 93.520 22.980 94.060 ;
        RECT 23.760 93.905 23.900 94.060 ;
        RECT 31.950 94.000 32.270 94.060 ;
        RECT 32.425 94.015 32.715 94.245 ;
        RECT 33.330 94.015 33.715 94.245 ;
        RECT 35.185 94.200 35.475 94.245 ;
        RECT 37.930 94.200 38.250 94.260 ;
        RECT 35.185 94.060 38.250 94.200 ;
        RECT 35.185 94.015 35.475 94.060 ;
        RECT 23.225 93.675 23.515 93.905 ;
        RECT 23.685 93.675 23.975 93.905 ;
        RECT 20.310 93.380 22.980 93.520 ;
        RECT 23.300 93.520 23.440 93.675 ;
        RECT 24.130 93.660 24.450 93.920 ;
        RECT 25.050 93.905 25.370 93.920 ;
        RECT 25.020 93.675 25.370 93.905 ;
        RECT 25.050 93.660 25.370 93.675 ;
        RECT 24.220 93.520 24.360 93.660 ;
        RECT 23.300 93.380 24.360 93.520 ;
        RECT 24.565 93.520 24.855 93.565 ;
        RECT 25.755 93.520 26.045 93.565 ;
        RECT 28.275 93.520 28.565 93.565 ;
        RECT 24.565 93.380 28.565 93.520 ;
        RECT 32.500 93.520 32.640 94.015 ;
        RECT 33.330 94.000 33.650 94.015 ;
        RECT 37.930 94.000 38.250 94.060 ;
        RECT 34.710 93.660 35.030 93.920 ;
        RECT 36.090 93.660 36.410 93.920 ;
        RECT 49.060 93.905 49.200 94.400 ;
        RECT 51.270 94.340 51.590 94.400 ;
        RECT 51.745 94.355 52.035 94.400 ;
        RECT 52.665 94.540 52.955 94.585 ;
        RECT 53.110 94.540 53.430 94.600 ;
        RECT 52.665 94.400 53.430 94.540 ;
        RECT 52.665 94.355 52.955 94.400 ;
        RECT 53.110 94.340 53.430 94.400 ;
        RECT 60.025 94.540 60.315 94.585 ;
        RECT 60.470 94.540 60.790 94.600 ;
        RECT 63.690 94.540 64.010 94.600 ;
        RECT 60.025 94.400 64.010 94.540 ;
        RECT 60.025 94.355 60.315 94.400 ;
        RECT 60.470 94.340 60.790 94.400 ;
        RECT 63.690 94.340 64.010 94.400 ;
        RECT 71.970 94.340 72.290 94.600 ;
        RECT 75.650 94.340 75.970 94.600 ;
        RECT 78.870 94.340 79.190 94.600 ;
        RECT 80.250 94.540 80.570 94.600 ;
        RECT 83.945 94.540 84.235 94.585 ;
        RECT 80.250 94.400 84.235 94.540 ;
        RECT 80.250 94.340 80.570 94.400 ;
        RECT 83.945 94.355 84.235 94.400 ;
        RECT 50.350 94.200 50.670 94.260 ;
        RECT 55.870 94.200 56.190 94.260 ;
        RECT 56.345 94.200 56.635 94.245 ;
        RECT 58.170 94.200 58.490 94.260 ;
        RECT 83.010 94.200 83.330 94.260 ;
        RECT 50.350 94.060 55.180 94.200 ;
        RECT 50.350 94.000 50.670 94.060 ;
        RECT 48.985 93.675 49.275 93.905 ;
        RECT 52.190 93.660 52.510 93.920 ;
        RECT 53.570 93.905 53.890 93.920 ;
        RECT 53.570 93.675 54.025 93.905 ;
        RECT 54.505 93.675 54.795 93.905 ;
        RECT 55.040 93.860 55.180 94.060 ;
        RECT 55.870 94.060 61.160 94.200 ;
        RECT 55.870 94.000 56.190 94.060 ;
        RECT 56.345 94.015 56.635 94.060 ;
        RECT 58.170 94.000 58.490 94.060 ;
        RECT 61.020 93.905 61.160 94.060 ;
        RECT 76.660 94.060 86.920 94.200 ;
        RECT 57.265 93.860 57.555 93.905 ;
        RECT 58.645 93.860 58.935 93.905 ;
        RECT 55.040 93.720 58.935 93.860 ;
        RECT 57.265 93.675 57.555 93.720 ;
        RECT 58.645 93.675 58.935 93.720 ;
        RECT 59.565 93.675 59.855 93.905 ;
        RECT 60.945 93.675 61.235 93.905 ;
        RECT 62.325 93.860 62.615 93.905 ;
        RECT 67.830 93.860 68.150 93.920 ;
        RECT 71.050 93.860 71.370 93.920 ;
        RECT 62.325 93.720 71.370 93.860 ;
        RECT 62.325 93.675 62.615 93.720 ;
        RECT 53.570 93.660 53.890 93.675 ;
        RECT 35.170 93.520 35.490 93.580 ;
        RECT 32.500 93.380 35.490 93.520 ;
        RECT 15.365 93.335 15.655 93.380 ;
        RECT 16.555 93.335 16.845 93.380 ;
        RECT 19.075 93.335 19.365 93.380 ;
        RECT 24.565 93.335 24.855 93.380 ;
        RECT 25.755 93.335 26.045 93.380 ;
        RECT 28.275 93.335 28.565 93.380 ;
        RECT 35.170 93.320 35.490 93.380 ;
        RECT 49.445 93.520 49.735 93.565 ;
        RECT 49.890 93.520 50.210 93.580 ;
        RECT 54.580 93.520 54.720 93.675 ;
        RECT 54.950 93.520 55.270 93.580 ;
        RECT 59.640 93.520 59.780 93.675 ;
        RECT 49.445 93.380 50.210 93.520 ;
        RECT 49.445 93.335 49.735 93.380 ;
        RECT 49.890 93.320 50.210 93.380 ;
        RECT 50.900 93.380 59.780 93.520 ;
        RECT 60.010 93.520 60.330 93.580 ;
        RECT 62.400 93.520 62.540 93.675 ;
        RECT 67.830 93.660 68.150 93.720 ;
        RECT 71.050 93.660 71.370 93.720 ;
        RECT 72.890 93.660 73.210 93.920 ;
        RECT 74.745 93.860 75.035 93.905 ;
        RECT 76.110 93.860 76.430 93.920 ;
        RECT 76.660 93.905 76.800 94.060 ;
        RECT 83.010 94.000 83.330 94.060 ;
        RECT 74.745 93.720 76.430 93.860 ;
        RECT 74.745 93.675 75.035 93.720 ;
        RECT 76.110 93.660 76.430 93.720 ;
        RECT 76.585 93.675 76.875 93.905 ;
        RECT 77.030 93.660 77.350 93.920 ;
        RECT 77.965 93.860 78.255 93.905 ;
        RECT 79.330 93.860 79.650 93.920 ;
        RECT 77.965 93.720 79.650 93.860 ;
        RECT 77.965 93.675 78.255 93.720 ;
        RECT 79.330 93.660 79.650 93.720 ;
        RECT 79.805 93.675 80.095 93.905 ;
        RECT 60.010 93.380 62.540 93.520 ;
        RECT 62.785 93.520 63.075 93.565 ;
        RECT 64.610 93.520 64.930 93.580 ;
        RECT 68.290 93.520 68.610 93.580 ;
        RECT 62.785 93.380 68.610 93.520 ;
        RECT 79.880 93.520 80.020 93.675 ;
        RECT 80.710 93.660 81.030 93.920 ;
        RECT 81.630 93.660 81.950 93.920 ;
        RECT 83.470 93.860 83.790 93.920 ;
        RECT 84.865 93.860 85.155 93.905 ;
        RECT 83.470 93.720 85.155 93.860 ;
        RECT 83.470 93.660 83.790 93.720 ;
        RECT 84.865 93.675 85.155 93.720 ;
        RECT 85.310 93.660 85.630 93.920 ;
        RECT 86.780 93.905 86.920 94.060 ;
        RECT 85.785 93.675 86.075 93.905 ;
        RECT 86.705 93.675 86.995 93.905 ;
        RECT 100.130 93.895 100.750 99.785 ;
        RECT 80.250 93.520 80.570 93.580 ;
        RECT 79.880 93.380 80.570 93.520 ;
        RECT 50.900 93.225 51.040 93.380 ;
        RECT 54.950 93.320 55.270 93.380 ;
        RECT 60.010 93.320 60.330 93.380 ;
        RECT 62.785 93.335 63.075 93.380 ;
        RECT 64.610 93.320 64.930 93.380 ;
        RECT 68.290 93.320 68.610 93.380 ;
        RECT 80.250 93.320 80.570 93.380 ;
        RECT 84.390 93.520 84.710 93.580 ;
        RECT 85.860 93.520 86.000 93.675 ;
        RECT 100.130 93.615 100.370 93.895 ;
        RECT 100.520 93.835 100.750 93.895 ;
        RECT 100.960 93.895 101.430 99.835 ;
        RECT 102.100 99.765 102.330 99.835 ;
        RECT 101.800 93.915 102.330 99.765 ;
        RECT 101.800 93.895 101.960 93.915 ;
        RECT 100.960 93.835 101.190 93.895 ;
        RECT 101.810 93.655 101.960 93.895 ;
        RECT 102.100 93.835 102.330 93.915 ;
        RECT 102.540 93.915 103.010 99.835 ;
        RECT 103.680 99.765 103.910 99.835 ;
        RECT 103.310 95.175 103.920 99.765 ;
        RECT 102.540 93.835 102.770 93.915 ;
        RECT 103.290 93.885 103.920 95.175 ;
        RECT 104.120 93.925 104.600 99.835 ;
        RECT 105.260 99.785 105.490 99.835 ;
        RECT 88.530 93.520 88.850 93.580 ;
        RECT 84.390 93.380 88.850 93.520 ;
        RECT 84.390 93.320 84.710 93.380 ;
        RECT 88.530 93.320 88.850 93.380 ;
        RECT 14.970 93.180 15.260 93.225 ;
        RECT 17.070 93.180 17.360 93.225 ;
        RECT 18.640 93.180 18.930 93.225 ;
        RECT 14.970 93.040 18.930 93.180 ;
        RECT 14.970 92.995 15.260 93.040 ;
        RECT 17.070 92.995 17.360 93.040 ;
        RECT 18.640 92.995 18.930 93.040 ;
        RECT 24.170 93.180 24.460 93.225 ;
        RECT 26.270 93.180 26.560 93.225 ;
        RECT 27.840 93.180 28.130 93.225 ;
        RECT 24.170 93.040 28.130 93.180 ;
        RECT 24.170 92.995 24.460 93.040 ;
        RECT 26.270 92.995 26.560 93.040 ;
        RECT 27.840 92.995 28.130 93.040 ;
        RECT 50.825 92.995 51.115 93.225 ;
        RECT 58.185 93.180 58.475 93.225 ;
        RECT 62.310 93.180 62.630 93.240 ;
        RECT 65.530 93.180 65.850 93.240 ;
        RECT 58.185 93.040 65.850 93.180 ;
        RECT 58.185 92.995 58.475 93.040 ;
        RECT 62.310 92.980 62.630 93.040 ;
        RECT 65.530 92.980 65.850 93.040 ;
        RECT 73.825 93.180 74.115 93.225 ;
        RECT 81.630 93.180 81.950 93.240 ;
        RECT 73.825 93.040 81.950 93.180 ;
        RECT 73.825 92.995 74.115 93.040 ;
        RECT 81.630 92.980 81.950 93.040 ;
        RECT 82.550 92.980 82.870 93.240 ;
        RECT 23.225 92.840 23.515 92.885 ;
        RECT 25.510 92.840 25.830 92.900 ;
        RECT 23.225 92.700 25.830 92.840 ;
        RECT 23.225 92.655 23.515 92.700 ;
        RECT 25.510 92.640 25.830 92.700 ;
        RECT 26.890 92.840 27.210 92.900 ;
        RECT 30.585 92.840 30.875 92.885 ;
        RECT 26.890 92.700 30.875 92.840 ;
        RECT 26.890 92.640 27.210 92.700 ;
        RECT 30.585 92.655 30.875 92.700 ;
        RECT 32.870 92.840 33.190 92.900 ;
        RECT 33.345 92.840 33.635 92.885 ;
        RECT 32.870 92.700 33.635 92.840 ;
        RECT 32.870 92.640 33.190 92.700 ;
        RECT 33.345 92.655 33.635 92.700 ;
        RECT 34.250 92.640 34.570 92.900 ;
        RECT 35.630 92.840 35.950 92.900 ;
        RECT 37.025 92.840 37.315 92.885 ;
        RECT 35.630 92.700 37.315 92.840 ;
        RECT 35.630 92.640 35.950 92.700 ;
        RECT 37.025 92.655 37.315 92.700 ;
        RECT 42.070 92.840 42.390 92.900 ;
        RECT 48.985 92.840 49.275 92.885 ;
        RECT 42.070 92.700 49.275 92.840 ;
        RECT 42.070 92.640 42.390 92.700 ;
        RECT 48.985 92.655 49.275 92.700 ;
        RECT 69.670 92.840 69.990 92.900 ;
        RECT 77.950 92.840 78.270 92.900 ;
        RECT 69.670 92.700 78.270 92.840 ;
        RECT 69.670 92.640 69.990 92.700 ;
        RECT 77.950 92.640 78.270 92.700 ;
        RECT 80.725 92.840 81.015 92.885 ;
        RECT 83.930 92.840 84.250 92.900 ;
        RECT 80.725 92.700 84.250 92.840 ;
        RECT 80.725 92.655 81.015 92.700 ;
        RECT 83.930 92.640 84.250 92.700 ;
        RECT 12.100 92.020 89.840 92.500 ;
        RECT 18.150 91.820 18.470 91.880 ;
        RECT 24.605 91.820 24.895 91.865 ;
        RECT 25.050 91.820 25.370 91.880 ;
        RECT 18.150 91.680 22.060 91.820 ;
        RECT 18.150 91.620 18.470 91.680 ;
        RECT 21.920 91.525 22.060 91.680 ;
        RECT 24.605 91.680 25.370 91.820 ;
        RECT 24.605 91.635 24.895 91.680 ;
        RECT 25.050 91.620 25.370 91.680 ;
        RECT 31.965 91.820 32.255 91.865 ;
        RECT 32.870 91.820 33.190 91.880 ;
        RECT 31.965 91.680 33.190 91.820 ;
        RECT 31.965 91.635 32.255 91.680 ;
        RECT 32.870 91.620 33.190 91.680 ;
        RECT 36.090 91.820 36.410 91.880 ;
        RECT 40.245 91.820 40.535 91.865 ;
        RECT 36.090 91.680 40.535 91.820 ;
        RECT 36.090 91.620 36.410 91.680 ;
        RECT 40.245 91.635 40.535 91.680 ;
        RECT 51.270 91.820 51.590 91.880 ;
        RECT 53.110 91.820 53.430 91.880 ;
        RECT 51.270 91.680 53.430 91.820 ;
        RECT 51.270 91.620 51.590 91.680 ;
        RECT 53.110 91.620 53.430 91.680 ;
        RECT 55.410 91.620 55.730 91.880 ;
        RECT 58.645 91.820 58.935 91.865 ;
        RECT 60.930 91.820 61.250 91.880 ;
        RECT 58.645 91.680 61.250 91.820 ;
        RECT 58.645 91.635 58.935 91.680 ;
        RECT 60.930 91.620 61.250 91.680 ;
        RECT 71.510 91.820 71.830 91.880 ;
        RECT 83.470 91.820 83.790 91.880 ;
        RECT 71.510 91.680 83.790 91.820 ;
        RECT 71.510 91.620 71.830 91.680 ;
        RECT 83.470 91.620 83.790 91.680 ;
        RECT 14.050 91.480 14.340 91.525 ;
        RECT 16.150 91.480 16.440 91.525 ;
        RECT 17.720 91.480 18.010 91.525 ;
        RECT 14.050 91.340 18.010 91.480 ;
        RECT 14.050 91.295 14.340 91.340 ;
        RECT 16.150 91.295 16.440 91.340 ;
        RECT 17.720 91.295 18.010 91.340 ;
        RECT 21.845 91.295 22.135 91.525 ;
        RECT 33.370 91.480 33.660 91.525 ;
        RECT 35.470 91.480 35.760 91.525 ;
        RECT 37.040 91.480 37.330 91.525 ;
        RECT 33.370 91.340 37.330 91.480 ;
        RECT 33.370 91.295 33.660 91.340 ;
        RECT 35.470 91.295 35.760 91.340 ;
        RECT 37.040 91.295 37.330 91.340 ;
        RECT 42.990 91.480 43.280 91.525 ;
        RECT 44.560 91.480 44.850 91.525 ;
        RECT 46.660 91.480 46.950 91.525 ;
        RECT 59.090 91.480 59.410 91.540 ;
        RECT 42.990 91.340 46.950 91.480 ;
        RECT 42.990 91.295 43.280 91.340 ;
        RECT 44.560 91.295 44.850 91.340 ;
        RECT 46.660 91.295 46.950 91.340 ;
        RECT 55.960 91.340 59.410 91.480 ;
        RECT 13.550 90.940 13.870 91.200 ;
        RECT 14.445 91.140 14.735 91.185 ;
        RECT 15.635 91.140 15.925 91.185 ;
        RECT 18.155 91.140 18.445 91.185 ;
        RECT 30.110 91.140 30.430 91.200 ;
        RECT 14.445 91.000 18.445 91.140 ;
        RECT 14.445 90.955 14.735 91.000 ;
        RECT 15.635 90.955 15.925 91.000 ;
        RECT 18.155 90.955 18.445 91.000 ;
        RECT 29.280 91.000 30.430 91.140 ;
        RECT 14.010 90.800 14.330 90.860 ;
        RECT 14.845 90.800 15.135 90.845 ;
        RECT 14.010 90.660 15.135 90.800 ;
        RECT 14.010 90.600 14.330 90.660 ;
        RECT 14.845 90.615 15.135 90.660 ;
        RECT 25.510 90.600 25.830 90.860 ;
        RECT 26.890 90.600 27.210 90.860 ;
        RECT 27.365 90.615 27.655 90.845 ;
        RECT 27.810 90.800 28.130 90.860 ;
        RECT 29.280 90.800 29.420 91.000 ;
        RECT 30.110 90.940 30.430 91.000 ;
        RECT 31.950 91.140 32.270 91.200 ;
        RECT 32.870 91.140 33.190 91.200 ;
        RECT 31.950 91.000 33.190 91.140 ;
        RECT 31.950 90.940 32.270 91.000 ;
        RECT 32.870 90.940 33.190 91.000 ;
        RECT 33.765 91.140 34.055 91.185 ;
        RECT 34.955 91.140 35.245 91.185 ;
        RECT 37.475 91.140 37.765 91.185 ;
        RECT 33.765 91.000 37.765 91.140 ;
        RECT 33.765 90.955 34.055 91.000 ;
        RECT 34.955 90.955 35.245 91.000 ;
        RECT 37.475 90.955 37.765 91.000 ;
        RECT 42.555 91.140 42.845 91.185 ;
        RECT 45.075 91.140 45.365 91.185 ;
        RECT 46.265 91.140 46.555 91.185 ;
        RECT 55.410 91.140 55.730 91.200 ;
        RECT 42.555 91.000 46.555 91.140 ;
        RECT 42.555 90.955 42.845 91.000 ;
        RECT 45.075 90.955 45.365 91.000 ;
        RECT 46.265 90.955 46.555 91.000 ;
        RECT 54.120 91.000 55.730 91.140 ;
        RECT 27.810 90.660 29.420 90.800 ;
        RECT 29.650 90.800 29.970 90.860 ;
        RECT 34.250 90.845 34.570 90.860 ;
        RECT 30.585 90.800 30.875 90.845 ;
        RECT 29.650 90.660 30.875 90.800 ;
        RECT 20.910 90.460 21.230 90.520 ;
        RECT 22.765 90.460 23.055 90.505 ;
        RECT 20.910 90.320 23.055 90.460 ;
        RECT 20.910 90.260 21.230 90.320 ;
        RECT 22.765 90.275 23.055 90.320 ;
        RECT 26.430 90.260 26.750 90.520 ;
        RECT 27.440 90.460 27.580 90.615 ;
        RECT 27.810 90.600 28.130 90.660 ;
        RECT 29.650 90.600 29.970 90.660 ;
        RECT 30.585 90.615 30.875 90.660 ;
        RECT 31.505 90.615 31.795 90.845 ;
        RECT 32.425 90.615 32.715 90.845 ;
        RECT 34.220 90.800 34.570 90.845 ;
        RECT 34.055 90.660 34.570 90.800 ;
        RECT 34.220 90.615 34.570 90.660 ;
        RECT 30.110 90.460 30.430 90.520 ;
        RECT 31.580 90.460 31.720 90.615 ;
        RECT 27.440 90.320 29.420 90.460 ;
        RECT 29.280 90.180 29.420 90.320 ;
        RECT 30.110 90.320 31.720 90.460 ;
        RECT 30.110 90.260 30.430 90.320 ;
        RECT 20.465 90.120 20.755 90.165 ;
        RECT 21.830 90.120 22.150 90.180 ;
        RECT 20.465 89.980 22.150 90.120 ;
        RECT 20.465 89.935 20.755 89.980 ;
        RECT 21.830 89.920 22.150 89.980 ;
        RECT 23.210 89.920 23.530 90.180 ;
        RECT 23.685 90.120 23.975 90.165 ;
        RECT 24.130 90.120 24.450 90.180 ;
        RECT 23.685 89.980 24.450 90.120 ;
        RECT 23.685 89.935 23.975 89.980 ;
        RECT 24.130 89.920 24.450 89.980 ;
        RECT 27.350 90.120 27.670 90.180 ;
        RECT 28.285 90.120 28.575 90.165 ;
        RECT 27.350 89.980 28.575 90.120 ;
        RECT 27.350 89.920 27.670 89.980 ;
        RECT 28.285 89.935 28.575 89.980 ;
        RECT 29.190 89.920 29.510 90.180 ;
        RECT 32.500 90.120 32.640 90.615 ;
        RECT 34.250 90.600 34.570 90.615 ;
        RECT 47.130 90.600 47.450 90.860 ;
        RECT 53.125 90.800 53.415 90.845 ;
        RECT 53.570 90.800 53.890 90.860 ;
        RECT 54.120 90.845 54.260 91.000 ;
        RECT 55.410 90.940 55.730 91.000 ;
        RECT 53.125 90.660 53.890 90.800 ;
        RECT 53.125 90.615 53.415 90.660 ;
        RECT 53.570 90.600 53.890 90.660 ;
        RECT 54.045 90.615 54.335 90.845 ;
        RECT 55.960 90.800 56.100 91.340 ;
        RECT 59.090 91.280 59.410 91.340 ;
        RECT 60.485 91.480 60.775 91.525 ;
        RECT 65.070 91.480 65.390 91.540 ;
        RECT 75.650 91.480 75.970 91.540 ;
        RECT 60.485 91.340 65.390 91.480 ;
        RECT 60.485 91.295 60.775 91.340 ;
        RECT 65.070 91.280 65.390 91.340 ;
        RECT 72.520 91.340 75.970 91.480 ;
        RECT 57.250 91.140 57.570 91.200 ;
        RECT 60.945 91.140 61.235 91.185 ;
        RECT 63.230 91.140 63.550 91.200 ;
        RECT 57.250 91.000 59.780 91.140 ;
        RECT 57.250 90.940 57.570 91.000 ;
        RECT 54.580 90.660 56.100 90.800 ;
        RECT 56.330 90.800 56.650 90.860 ;
        RECT 57.340 90.800 57.480 90.940 ;
        RECT 56.330 90.660 57.480 90.800 ;
        RECT 36.550 90.460 36.870 90.520 ;
        RECT 45.810 90.460 46.100 90.505 ;
        RECT 36.550 90.320 46.100 90.460 ;
        RECT 36.550 90.260 36.870 90.320 ;
        RECT 45.810 90.275 46.100 90.320 ;
        RECT 51.730 90.460 52.050 90.520 ;
        RECT 54.580 90.505 54.720 90.660 ;
        RECT 56.330 90.600 56.650 90.660 ;
        RECT 58.630 90.600 58.950 90.860 ;
        RECT 59.640 90.845 59.780 91.000 ;
        RECT 60.945 91.000 63.550 91.140 ;
        RECT 60.945 90.955 61.235 91.000 ;
        RECT 63.230 90.940 63.550 91.000 ;
        RECT 59.105 90.615 59.395 90.845 ;
        RECT 59.565 90.615 59.855 90.845 ;
        RECT 60.025 90.800 60.315 90.845 ;
        RECT 60.470 90.800 60.790 90.860 ;
        RECT 68.750 90.800 69.070 90.860 ;
        RECT 60.025 90.660 60.790 90.800 ;
        RECT 60.025 90.615 60.315 90.660 ;
        RECT 54.505 90.460 54.795 90.505 ;
        RECT 55.585 90.460 55.875 90.505 ;
        RECT 56.420 90.460 56.560 90.600 ;
        RECT 51.730 90.320 54.795 90.460 ;
        RECT 55.375 90.320 56.560 90.460 ;
        RECT 56.790 90.460 57.110 90.520 ;
        RECT 58.720 90.460 58.860 90.600 ;
        RECT 56.790 90.320 58.860 90.460 ;
        RECT 59.180 90.460 59.320 90.615 ;
        RECT 60.470 90.600 60.790 90.660 ;
        RECT 61.020 90.660 69.070 90.800 ;
        RECT 61.020 90.460 61.160 90.660 ;
        RECT 68.750 90.600 69.070 90.660 ;
        RECT 71.970 90.600 72.290 90.860 ;
        RECT 72.520 90.845 72.660 91.340 ;
        RECT 75.650 91.280 75.970 91.340 ;
        RECT 77.530 91.480 77.820 91.525 ;
        RECT 79.630 91.480 79.920 91.525 ;
        RECT 81.200 91.480 81.490 91.525 ;
        RECT 77.530 91.340 81.490 91.480 ;
        RECT 77.530 91.295 77.820 91.340 ;
        RECT 79.630 91.295 79.920 91.340 ;
        RECT 81.200 91.295 81.490 91.340 ;
        RECT 77.925 91.140 78.215 91.185 ;
        RECT 79.115 91.140 79.405 91.185 ;
        RECT 81.635 91.140 81.925 91.185 ;
        RECT 77.925 91.000 81.925 91.140 ;
        RECT 77.925 90.955 78.215 91.000 ;
        RECT 79.115 90.955 79.405 91.000 ;
        RECT 81.635 90.955 81.925 91.000 ;
        RECT 83.930 91.140 84.250 91.200 ;
        RECT 100.130 91.185 100.510 93.615 ;
        RECT 100.710 93.605 101.000 93.630 ;
        RECT 100.700 92.905 101.020 93.605 ;
        RECT 100.650 91.875 101.650 92.905 ;
        RECT 100.700 91.185 101.020 91.875 ;
        RECT 83.930 91.000 86.460 91.140 ;
        RECT 83.930 90.940 84.250 91.000 ;
        RECT 72.445 90.615 72.735 90.845 ;
        RECT 72.890 90.600 73.210 90.860 ;
        RECT 73.810 90.600 74.130 90.860 ;
        RECT 74.285 90.615 74.575 90.845 ;
        RECT 74.745 90.800 75.035 90.845 ;
        RECT 76.570 90.800 76.890 90.860 ;
        RECT 74.745 90.660 76.890 90.800 ;
        RECT 74.745 90.615 75.035 90.660 ;
        RECT 59.180 90.320 61.160 90.460 ;
        RECT 51.730 90.260 52.050 90.320 ;
        RECT 54.505 90.275 54.795 90.320 ;
        RECT 55.500 90.275 55.875 90.320 ;
        RECT 37.930 90.120 38.250 90.180 ;
        RECT 39.785 90.120 40.075 90.165 ;
        RECT 32.500 89.980 40.075 90.120 ;
        RECT 37.930 89.920 38.250 89.980 ;
        RECT 39.785 89.935 40.075 89.980 ;
        RECT 53.110 90.120 53.430 90.180 ;
        RECT 53.585 90.120 53.875 90.165 ;
        RECT 53.110 89.980 53.875 90.120 ;
        RECT 53.110 89.920 53.430 89.980 ;
        RECT 53.585 89.935 53.875 89.980 ;
        RECT 54.030 90.120 54.350 90.180 ;
        RECT 55.500 90.120 55.640 90.275 ;
        RECT 56.790 90.260 57.110 90.320 ;
        RECT 61.405 90.275 61.695 90.505 ;
        RECT 54.030 89.980 55.640 90.120 ;
        RECT 54.030 89.920 54.350 89.980 ;
        RECT 56.330 89.920 56.650 90.180 ;
        RECT 57.265 90.120 57.555 90.165 ;
        RECT 58.630 90.120 58.950 90.180 ;
        RECT 57.265 89.980 58.950 90.120 ;
        RECT 57.265 89.935 57.555 89.980 ;
        RECT 58.630 89.920 58.950 89.980 ;
        RECT 59.550 90.120 59.870 90.180 ;
        RECT 61.480 90.120 61.620 90.275 ;
        RECT 62.310 90.260 62.630 90.520 ;
        RECT 72.060 90.460 72.200 90.600 ;
        RECT 74.360 90.460 74.500 90.615 ;
        RECT 76.570 90.600 76.890 90.660 ;
        RECT 77.045 90.800 77.335 90.845 ;
        RECT 80.250 90.800 80.570 90.860 ;
        RECT 86.320 90.845 86.460 91.000 ;
        RECT 100.130 90.875 100.370 91.185 ;
        RECT 100.720 91.145 101.020 91.185 ;
        RECT 100.720 91.135 101.010 91.145 ;
        RECT 101.810 91.125 102.010 93.655 ;
        RECT 102.290 93.625 102.580 93.630 ;
        RECT 102.280 92.955 102.620 93.625 ;
        RECT 102.150 91.925 103.150 92.955 ;
        RECT 102.280 91.155 102.620 91.925 ;
        RECT 102.300 91.135 102.590 91.155 ;
        RECT 100.530 90.875 100.760 90.975 ;
        RECT 100.130 90.865 100.760 90.875 ;
        RECT 85.785 90.800 86.075 90.845 ;
        RECT 77.045 90.660 79.560 90.800 ;
        RECT 77.045 90.615 77.335 90.660 ;
        RECT 79.420 90.520 79.560 90.660 ;
        RECT 80.250 90.660 86.075 90.800 ;
        RECT 80.250 90.600 80.570 90.660 ;
        RECT 85.785 90.615 86.075 90.660 ;
        RECT 86.245 90.615 86.535 90.845 ;
        RECT 86.690 90.600 87.010 90.860 ;
        RECT 87.625 90.800 87.915 90.845 ;
        RECT 88.070 90.800 88.390 90.860 ;
        RECT 87.625 90.660 88.390 90.800 ;
        RECT 87.625 90.615 87.915 90.660 ;
        RECT 75.190 90.460 75.510 90.520 ;
        RECT 72.060 90.320 75.510 90.460 ;
        RECT 75.190 90.260 75.510 90.320 ;
        RECT 76.125 90.460 76.415 90.505 ;
        RECT 78.270 90.460 78.560 90.505 ;
        RECT 76.125 90.320 78.560 90.460 ;
        RECT 76.125 90.275 76.415 90.320 ;
        RECT 78.270 90.275 78.560 90.320 ;
        RECT 79.330 90.260 79.650 90.520 ;
        RECT 80.710 90.460 81.030 90.520 ;
        RECT 82.090 90.460 82.410 90.520 ;
        RECT 80.710 90.320 82.410 90.460 ;
        RECT 80.710 90.260 81.030 90.320 ;
        RECT 82.090 90.260 82.410 90.320 ;
        RECT 85.310 90.460 85.630 90.520 ;
        RECT 87.700 90.460 87.840 90.615 ;
        RECT 88.070 90.600 88.390 90.660 ;
        RECT 85.310 90.320 87.840 90.460 ;
        RECT 85.310 90.260 85.630 90.320 ;
        RECT 59.550 89.980 61.620 90.120 ;
        RECT 63.245 90.120 63.535 90.165 ;
        RECT 65.990 90.120 66.310 90.180 ;
        RECT 63.245 89.980 66.310 90.120 ;
        RECT 59.550 89.920 59.870 89.980 ;
        RECT 63.245 89.935 63.535 89.980 ;
        RECT 65.990 89.920 66.310 89.980 ;
        RECT 69.210 90.120 69.530 90.180 ;
        RECT 71.050 90.120 71.370 90.180 ;
        RECT 69.210 89.980 71.370 90.120 ;
        RECT 69.210 89.920 69.530 89.980 ;
        RECT 71.050 89.920 71.370 89.980 ;
        RECT 71.985 90.120 72.275 90.165 ;
        RECT 73.350 90.120 73.670 90.180 ;
        RECT 71.985 89.980 73.670 90.120 ;
        RECT 71.985 89.935 72.275 89.980 ;
        RECT 73.350 89.920 73.670 89.980 ;
        RECT 76.570 90.120 76.890 90.180 ;
        RECT 81.630 90.120 81.950 90.180 ;
        RECT 83.945 90.120 84.235 90.165 ;
        RECT 76.570 89.980 84.235 90.120 ;
        RECT 76.570 89.920 76.890 89.980 ;
        RECT 81.630 89.920 81.950 89.980 ;
        RECT 83.945 89.935 84.235 89.980 ;
        RECT 84.390 89.920 84.710 90.180 ;
        RECT 12.100 89.300 89.840 89.780 ;
        RECT 21.370 89.100 21.690 89.160 ;
        RECT 22.305 89.100 22.595 89.145 ;
        RECT 21.370 88.960 22.595 89.100 ;
        RECT 21.370 88.900 21.690 88.960 ;
        RECT 22.305 88.915 22.595 88.960 ;
        RECT 24.130 88.900 24.450 89.160 ;
        RECT 26.430 88.900 26.750 89.160 ;
        RECT 28.745 89.100 29.035 89.145 ;
        RECT 29.650 89.100 29.970 89.160 ;
        RECT 36.090 89.100 36.410 89.160 ;
        RECT 28.745 88.960 29.970 89.100 ;
        RECT 28.745 88.915 29.035 88.960 ;
        RECT 29.650 88.900 29.970 88.960 ;
        RECT 31.580 88.960 36.410 89.100 ;
        RECT 23.210 88.760 23.530 88.820 ;
        RECT 31.580 88.805 31.720 88.960 ;
        RECT 36.090 88.900 36.410 88.960 ;
        RECT 36.550 88.900 36.870 89.160 ;
        RECT 51.730 89.100 52.050 89.160 ;
        RECT 52.205 89.100 52.495 89.145 ;
        RECT 51.730 88.960 52.495 89.100 ;
        RECT 51.730 88.900 52.050 88.960 ;
        RECT 52.205 88.915 52.495 88.960 ;
        RECT 53.570 88.900 53.890 89.160 ;
        RECT 54.490 88.900 54.810 89.160 ;
        RECT 55.410 89.100 55.730 89.160 ;
        RECT 60.945 89.100 61.235 89.145 ;
        RECT 55.410 88.960 61.235 89.100 ;
        RECT 55.410 88.900 55.730 88.960 ;
        RECT 60.945 88.915 61.235 88.960 ;
        RECT 61.850 89.100 62.170 89.160 ;
        RECT 63.245 89.100 63.535 89.145 ;
        RECT 61.850 88.960 63.535 89.100 ;
        RECT 61.850 88.900 62.170 88.960 ;
        RECT 63.245 88.915 63.535 88.960 ;
        RECT 64.150 88.900 64.470 89.160 ;
        RECT 69.685 89.100 69.975 89.145 ;
        RECT 83.010 89.100 83.330 89.160 ;
        RECT 69.685 88.960 83.330 89.100 ;
        RECT 100.100 89.065 100.760 90.865 ;
        RECT 100.130 89.045 100.360 89.065 ;
        RECT 100.530 88.975 100.760 89.065 ;
        RECT 100.970 90.905 101.200 90.975 ;
        RECT 100.970 89.095 101.530 90.905 ;
        RECT 101.810 90.865 101.960 91.125 ;
        RECT 102.110 90.865 102.340 90.975 ;
        RECT 101.810 90.855 102.340 90.865 ;
        RECT 100.970 88.975 101.200 89.095 ;
        RECT 69.685 88.915 69.975 88.960 ;
        RECT 83.010 88.900 83.330 88.960 ;
        RECT 23.210 88.620 29.880 88.760 ;
        RECT 23.210 88.560 23.530 88.620 ;
        RECT 13.550 88.220 13.870 88.480 ;
        RECT 14.930 88.465 15.250 88.480 ;
        RECT 14.900 88.235 15.250 88.465 ;
        RECT 14.930 88.220 15.250 88.235 ;
        RECT 16.770 88.420 17.090 88.480 ;
        RECT 20.925 88.420 21.215 88.465 ;
        RECT 16.770 88.280 21.215 88.420 ;
        RECT 16.770 88.220 17.090 88.280 ;
        RECT 20.925 88.235 21.215 88.280 ;
        RECT 21.845 88.235 22.135 88.465 ;
        RECT 22.290 88.420 22.610 88.480 ;
        RECT 22.765 88.420 23.055 88.465 ;
        RECT 22.290 88.280 23.055 88.420 ;
        RECT 14.445 88.080 14.735 88.125 ;
        RECT 15.635 88.080 15.925 88.125 ;
        RECT 18.155 88.080 18.445 88.125 ;
        RECT 14.445 87.940 18.445 88.080 ;
        RECT 21.920 88.080 22.060 88.235 ;
        RECT 22.290 88.220 22.610 88.280 ;
        RECT 22.765 88.235 23.055 88.280 ;
        RECT 23.685 88.420 23.975 88.465 ;
        RECT 24.590 88.420 24.910 88.480 ;
        RECT 25.065 88.420 25.355 88.465 ;
        RECT 23.685 88.280 25.355 88.420 ;
        RECT 23.685 88.235 23.975 88.280 ;
        RECT 24.590 88.220 24.910 88.280 ;
        RECT 25.065 88.235 25.355 88.280 ;
        RECT 25.985 88.420 26.275 88.465 ;
        RECT 26.890 88.420 27.210 88.480 ;
        RECT 25.985 88.280 27.210 88.420 ;
        RECT 25.985 88.235 26.275 88.280 ;
        RECT 26.060 88.080 26.200 88.235 ;
        RECT 26.890 88.220 27.210 88.280 ;
        RECT 27.810 88.220 28.130 88.480 ;
        RECT 28.270 88.220 28.590 88.480 ;
        RECT 29.740 88.465 29.880 88.620 ;
        RECT 31.505 88.575 31.795 88.805 ;
        RECT 31.950 88.760 32.270 88.820 ;
        RECT 32.505 88.760 32.795 88.805 ;
        RECT 34.710 88.760 35.030 88.820 ;
        RECT 31.950 88.620 35.030 88.760 ;
        RECT 31.950 88.560 32.270 88.620 ;
        RECT 32.505 88.575 32.795 88.620 ;
        RECT 34.710 88.560 35.030 88.620 ;
        RECT 35.170 88.760 35.490 88.820 ;
        RECT 35.645 88.760 35.935 88.805 ;
        RECT 38.850 88.760 39.170 88.820 ;
        RECT 41.625 88.760 41.915 88.805 ;
        RECT 35.170 88.620 41.915 88.760 ;
        RECT 54.580 88.760 54.720 88.900 ;
        RECT 57.250 88.760 57.570 88.820 ;
        RECT 61.405 88.760 61.695 88.805 ;
        RECT 54.580 88.620 56.100 88.760 ;
        RECT 35.170 88.560 35.490 88.620 ;
        RECT 35.645 88.575 35.935 88.620 ;
        RECT 38.850 88.560 39.170 88.620 ;
        RECT 41.625 88.575 41.915 88.620 ;
        RECT 29.665 88.235 29.955 88.465 ;
        RECT 30.110 88.420 30.430 88.480 ;
        RECT 32.040 88.420 32.180 88.560 ;
        RECT 30.110 88.280 32.180 88.420 ;
        RECT 33.805 88.420 34.095 88.465 ;
        RECT 43.005 88.420 43.295 88.465 ;
        RECT 33.805 88.280 43.295 88.420 ;
        RECT 30.110 88.220 30.430 88.280 ;
        RECT 33.805 88.235 34.095 88.280 ;
        RECT 43.005 88.235 43.295 88.280 ;
        RECT 43.450 88.420 43.770 88.480 ;
        RECT 43.925 88.420 44.215 88.465 ;
        RECT 43.450 88.280 44.215 88.420 ;
        RECT 21.920 87.940 26.200 88.080 ;
        RECT 26.430 88.080 26.750 88.140 ;
        RECT 30.585 88.080 30.875 88.125 ;
        RECT 26.430 87.940 30.875 88.080 ;
        RECT 14.445 87.895 14.735 87.940 ;
        RECT 15.635 87.895 15.925 87.940 ;
        RECT 18.155 87.895 18.445 87.940 ;
        RECT 26.430 87.880 26.750 87.940 ;
        RECT 30.585 87.895 30.875 87.940 ;
        RECT 14.050 87.740 14.340 87.785 ;
        RECT 16.150 87.740 16.440 87.785 ;
        RECT 17.720 87.740 18.010 87.785 ;
        RECT 14.050 87.600 18.010 87.740 ;
        RECT 14.050 87.555 14.340 87.600 ;
        RECT 16.150 87.555 16.440 87.600 ;
        RECT 17.720 87.555 18.010 87.600 ;
        RECT 20.450 87.740 20.770 87.800 ;
        RECT 24.590 87.740 24.910 87.800 ;
        RECT 28.270 87.740 28.590 87.800 ;
        RECT 31.490 87.740 31.810 87.800 ;
        RECT 20.450 87.600 28.590 87.740 ;
        RECT 20.450 87.540 20.770 87.600 ;
        RECT 24.590 87.540 24.910 87.600 ;
        RECT 28.270 87.540 28.590 87.600 ;
        RECT 28.820 87.600 31.810 87.740 ;
        RECT 21.370 87.400 21.690 87.460 ;
        RECT 28.820 87.400 28.960 87.600 ;
        RECT 31.490 87.540 31.810 87.600 ;
        RECT 33.345 87.740 33.635 87.785 ;
        RECT 33.880 87.740 34.020 88.235 ;
        RECT 43.450 88.220 43.770 88.280 ;
        RECT 43.925 88.235 44.215 88.280 ;
        RECT 50.350 88.220 50.670 88.480 ;
        RECT 51.270 88.220 51.590 88.480 ;
        RECT 52.190 88.420 52.510 88.480 ;
        RECT 53.125 88.420 53.415 88.465 ;
        RECT 52.190 88.280 53.415 88.420 ;
        RECT 52.190 88.220 52.510 88.280 ;
        RECT 53.125 88.235 53.415 88.280 ;
        RECT 54.490 88.220 54.810 88.480 ;
        RECT 54.950 88.220 55.270 88.480 ;
        RECT 55.960 88.465 56.100 88.620 ;
        RECT 57.250 88.620 61.695 88.760 ;
        RECT 63.690 88.760 64.010 88.820 ;
        RECT 64.925 88.760 65.215 88.805 ;
        RECT 57.250 88.560 57.570 88.620 ;
        RECT 61.405 88.575 61.695 88.620 ;
        RECT 62.555 88.590 62.845 88.635 ;
        RECT 55.885 88.235 56.175 88.465 ;
        RECT 58.645 88.420 58.935 88.465 ;
        RECT 59.105 88.420 59.395 88.465 ;
        RECT 56.420 88.280 59.395 88.420 ;
        RECT 34.250 87.740 34.570 87.800 ;
        RECT 33.345 87.600 34.570 87.740 ;
        RECT 33.345 87.555 33.635 87.600 ;
        RECT 34.250 87.540 34.570 87.600 ;
        RECT 35.170 87.740 35.490 87.800 ;
        RECT 39.785 87.740 40.075 87.785 ;
        RECT 44.845 87.740 45.135 87.785 ;
        RECT 35.170 87.600 40.075 87.740 ;
        RECT 35.170 87.540 35.490 87.600 ;
        RECT 39.785 87.555 40.075 87.600 ;
        RECT 41.700 87.600 45.135 87.740 ;
        RECT 51.360 87.740 51.500 88.220 ;
        RECT 55.040 87.740 55.180 88.220 ;
        RECT 56.420 88.140 56.560 88.280 ;
        RECT 58.645 88.235 58.935 88.280 ;
        RECT 59.105 88.235 59.395 88.280 ;
        RECT 60.010 88.420 60.330 88.480 ;
        RECT 62.500 88.420 62.845 88.590 ;
        RECT 63.690 88.620 65.215 88.760 ;
        RECT 63.690 88.560 64.010 88.620 ;
        RECT 64.925 88.575 65.215 88.620 ;
        RECT 65.990 88.560 66.310 88.820 ;
        RECT 68.305 88.760 68.595 88.805 ;
        RECT 71.985 88.760 72.275 88.805 ;
        RECT 73.810 88.760 74.130 88.820 ;
        RECT 76.585 88.760 76.875 88.805 ;
        RECT 68.305 88.620 73.580 88.760 ;
        RECT 68.305 88.575 68.595 88.620 ;
        RECT 71.985 88.575 72.275 88.620 ;
        RECT 60.010 88.405 62.845 88.420 ;
        RECT 60.010 88.280 62.640 88.405 ;
        RECT 60.010 88.220 60.330 88.280 ;
        RECT 67.830 88.220 68.150 88.480 ;
        RECT 70.605 88.235 70.895 88.465 ;
        RECT 71.065 88.235 71.355 88.465 ;
        RECT 72.890 88.420 73.210 88.480 ;
        RECT 73.440 88.465 73.580 88.620 ;
        RECT 73.810 88.620 76.875 88.760 ;
        RECT 73.810 88.560 74.130 88.620 ;
        RECT 76.585 88.575 76.875 88.620 ;
        RECT 77.030 88.760 77.350 88.820 ;
        RECT 78.425 88.760 78.715 88.805 ;
        RECT 81.170 88.760 81.490 88.820 ;
        RECT 77.030 88.620 78.715 88.760 ;
        RECT 77.030 88.560 77.350 88.620 ;
        RECT 78.425 88.575 78.715 88.620 ;
        RECT 80.340 88.620 81.490 88.760 ;
        RECT 73.365 88.420 73.655 88.465 ;
        RECT 72.890 88.280 73.655 88.420 ;
        RECT 55.425 88.080 55.715 88.125 ;
        RECT 56.330 88.080 56.650 88.140 ;
        RECT 55.425 87.940 56.650 88.080 ;
        RECT 55.425 87.895 55.715 87.940 ;
        RECT 56.330 87.880 56.650 87.940 ;
        RECT 57.250 88.080 57.570 88.140 ;
        RECT 58.185 88.080 58.475 88.125 ;
        RECT 57.250 87.940 59.320 88.080 ;
        RECT 57.250 87.880 57.570 87.940 ;
        RECT 58.185 87.895 58.475 87.940 ;
        RECT 59.180 87.740 59.320 87.940 ;
        RECT 59.550 87.880 59.870 88.140 ;
        RECT 60.930 88.080 61.250 88.140 ;
        RECT 64.150 88.080 64.470 88.140 ;
        RECT 69.210 88.080 69.530 88.140 ;
        RECT 60.930 87.940 64.470 88.080 ;
        RECT 60.930 87.880 61.250 87.940 ;
        RECT 64.150 87.880 64.470 87.940 ;
        RECT 68.610 87.940 69.530 88.080 ;
        RECT 63.230 87.740 63.550 87.800 ;
        RECT 68.610 87.740 68.750 87.940 ;
        RECT 69.210 87.880 69.530 87.940 ;
        RECT 51.360 87.600 54.720 87.740 ;
        RECT 55.040 87.600 58.860 87.740 ;
        RECT 59.180 87.600 68.750 87.740 ;
        RECT 70.680 87.740 70.820 88.235 ;
        RECT 71.140 88.080 71.280 88.235 ;
        RECT 72.890 88.220 73.210 88.280 ;
        RECT 73.365 88.235 73.655 88.280 ;
        RECT 74.285 88.235 74.575 88.465 ;
        RECT 76.110 88.420 76.430 88.480 ;
        RECT 77.505 88.420 77.795 88.465 ;
        RECT 76.110 88.280 77.795 88.420 ;
        RECT 73.810 88.080 74.130 88.140 ;
        RECT 74.360 88.080 74.500 88.235 ;
        RECT 76.110 88.220 76.430 88.280 ;
        RECT 77.505 88.235 77.795 88.280 ;
        RECT 79.790 88.220 80.110 88.480 ;
        RECT 80.340 88.465 80.480 88.620 ;
        RECT 81.170 88.560 81.490 88.620 ;
        RECT 82.520 88.760 82.810 88.805 ;
        RECT 84.390 88.760 84.710 88.820 ;
        RECT 101.360 88.775 101.530 89.095 ;
        RECT 101.770 89.055 102.340 90.855 ;
        RECT 101.820 89.045 102.340 89.055 ;
        RECT 102.110 88.975 102.340 89.045 ;
        RECT 102.550 90.925 102.780 90.975 ;
        RECT 102.550 90.895 103.060 90.925 ;
        RECT 102.550 89.085 103.090 90.895 ;
        RECT 103.290 90.875 103.480 93.885 ;
        RECT 103.680 93.835 103.910 93.885 ;
        RECT 104.120 93.835 104.350 93.925 ;
        RECT 104.870 93.885 105.490 99.785 ;
        RECT 103.840 92.955 104.200 93.635 ;
        RECT 103.660 91.925 104.660 92.955 ;
        RECT 103.840 91.135 104.200 91.925 ;
        RECT 103.690 90.875 103.920 90.975 ;
        RECT 103.290 90.205 103.920 90.875 ;
        RECT 102.550 88.975 102.780 89.085 ;
        RECT 102.920 88.855 103.090 89.085 ;
        RECT 103.310 89.005 103.920 90.205 ;
        RECT 103.690 88.975 103.920 89.005 ;
        RECT 104.130 90.925 104.360 90.975 ;
        RECT 104.130 89.045 104.670 90.925 ;
        RECT 104.890 90.905 105.060 93.885 ;
        RECT 105.260 93.835 105.490 93.885 ;
        RECT 105.700 93.915 106.190 99.835 ;
        RECT 106.840 99.755 107.070 99.835 ;
        RECT 105.700 93.835 105.930 93.915 ;
        RECT 106.430 93.875 107.070 99.755 ;
        RECT 105.450 93.625 105.740 93.630 ;
        RECT 105.440 92.985 105.780 93.625 ;
        RECT 105.270 91.955 106.270 92.985 ;
        RECT 105.440 91.145 105.780 91.955 ;
        RECT 105.460 91.135 105.750 91.145 ;
        RECT 105.270 90.905 105.500 90.975 ;
        RECT 104.890 90.865 105.500 90.905 ;
        RECT 104.870 89.065 105.500 90.865 ;
        RECT 104.900 89.045 105.500 89.065 ;
        RECT 104.130 88.975 104.360 89.045 ;
        RECT 82.520 88.620 84.710 88.760 ;
        RECT 82.520 88.575 82.810 88.620 ;
        RECT 84.390 88.560 84.710 88.620 ;
        RECT 100.000 88.635 101.000 88.645 ;
        RECT 101.280 88.635 101.530 88.775 ;
        RECT 102.910 88.635 103.090 88.855 ;
        RECT 104.500 88.805 104.670 89.045 ;
        RECT 105.270 88.975 105.500 89.045 ;
        RECT 105.710 90.905 105.940 90.975 ;
        RECT 105.710 89.025 106.250 90.905 ;
        RECT 106.440 90.895 106.630 93.875 ;
        RECT 106.840 93.835 107.070 93.875 ;
        RECT 107.270 93.865 107.710 100.195 ;
        RECT 108.890 99.835 109.330 100.195 ;
        RECT 110.480 99.835 110.920 100.195 ;
        RECT 112.060 99.835 112.500 100.195 ;
        RECT 108.420 99.815 108.650 99.835 ;
        RECT 107.970 93.885 108.650 99.815 ;
        RECT 107.280 93.835 107.510 93.865 ;
        RECT 107.030 93.625 107.320 93.630 ;
        RECT 107.010 92.955 107.370 93.625 ;
        RECT 106.820 91.925 107.820 92.955 ;
        RECT 107.010 91.135 107.370 91.925 ;
        RECT 106.850 90.895 107.080 90.975 ;
        RECT 106.440 89.045 107.080 90.895 ;
        RECT 105.710 88.975 105.940 89.025 ;
        RECT 104.490 88.635 104.670 88.805 ;
        RECT 106.080 88.635 106.250 89.025 ;
        RECT 106.850 88.975 107.080 89.045 ;
        RECT 107.290 90.925 107.520 90.975 ;
        RECT 107.980 90.935 108.240 93.885 ;
        RECT 108.420 93.835 108.650 93.885 ;
        RECT 108.860 93.895 109.330 99.835 ;
        RECT 110.000 99.795 110.230 99.835 ;
        RECT 108.860 93.835 109.090 93.895 ;
        RECT 109.550 93.885 110.230 99.795 ;
        RECT 108.610 93.625 108.900 93.630 ;
        RECT 108.580 92.985 108.920 93.625 ;
        RECT 108.440 91.955 109.440 92.985 ;
        RECT 108.580 91.135 108.920 91.955 ;
        RECT 108.430 90.935 108.660 90.975 ;
        RECT 107.290 89.045 107.830 90.925 ;
        RECT 107.290 88.975 107.520 89.045 ;
        RECT 107.660 88.635 107.830 89.045 ;
        RECT 107.980 89.015 108.660 90.935 ;
        RECT 108.430 88.975 108.660 89.015 ;
        RECT 108.870 90.915 109.100 90.975 ;
        RECT 108.870 89.035 109.420 90.915 ;
        RECT 109.600 90.895 109.860 93.885 ;
        RECT 110.000 93.835 110.230 93.885 ;
        RECT 110.440 93.875 110.920 99.835 ;
        RECT 111.580 99.795 111.810 99.835 ;
        RECT 111.150 93.905 111.810 99.795 ;
        RECT 111.150 93.885 111.410 93.905 ;
        RECT 110.440 93.835 110.670 93.875 ;
        RECT 111.160 93.675 111.410 93.885 ;
        RECT 111.580 93.835 111.810 93.905 ;
        RECT 112.020 93.925 112.500 99.835 ;
        RECT 112.020 93.835 112.250 93.925 ;
        RECT 110.190 93.625 110.480 93.630 ;
        RECT 110.180 92.955 110.510 93.625 ;
        RECT 110.010 91.925 111.010 92.955 ;
        RECT 110.180 91.135 110.510 91.925 ;
        RECT 111.160 91.575 111.460 93.675 ;
        RECT 111.770 93.625 112.060 93.630 ;
        RECT 111.750 92.975 112.110 93.625 ;
        RECT 111.670 91.945 112.670 92.975 ;
        RECT 111.240 91.125 111.460 91.575 ;
        RECT 111.750 91.135 112.110 91.945 ;
        RECT 110.010 90.895 110.240 90.975 ;
        RECT 109.580 89.045 110.240 90.895 ;
        RECT 108.870 88.975 109.100 89.035 ;
        RECT 109.260 88.635 109.420 89.035 ;
        RECT 110.010 88.975 110.240 89.045 ;
        RECT 110.450 90.915 110.680 90.975 ;
        RECT 110.450 89.025 111.000 90.915 ;
        RECT 111.240 90.885 111.420 91.125 ;
        RECT 111.590 90.885 111.820 90.975 ;
        RECT 111.240 90.735 111.820 90.885 ;
        RECT 111.210 89.065 111.820 90.735 ;
        RECT 111.220 89.035 111.820 89.065 ;
        RECT 110.450 88.975 110.680 89.025 ;
        RECT 110.830 88.635 111.000 89.025 ;
        RECT 111.590 88.975 111.820 89.035 ;
        RECT 112.030 90.915 112.260 90.975 ;
        RECT 112.030 89.065 112.720 90.915 ;
        RECT 112.030 88.975 112.260 89.065 ;
        RECT 112.410 88.815 112.720 89.065 ;
        RECT 112.390 88.775 112.720 88.815 ;
        RECT 112.390 88.635 112.880 88.775 ;
        RECT 100.000 88.605 112.880 88.635 ;
        RECT 99.980 88.550 112.880 88.605 ;
        RECT 113.070 88.550 113.700 101.660 ;
        RECT 119.900 101.650 120.990 101.675 ;
        RECT 134.480 99.950 135.430 101.710 ;
        RECT 136.630 99.960 138.450 102.060 ;
        RECT 139.570 99.960 141.390 102.060 ;
        RECT 142.470 99.960 144.300 102.090 ;
        RECT 145.440 99.960 147.270 102.090 ;
        RECT 148.420 99.970 150.250 102.100 ;
        RECT 136.630 99.955 136.880 99.960 ;
        RECT 138.110 99.955 138.360 99.960 ;
        RECT 139.590 99.955 139.840 99.960 ;
        RECT 141.070 99.955 141.320 99.960 ;
        RECT 142.550 99.955 142.800 99.960 ;
        RECT 144.030 99.955 144.280 99.960 ;
        RECT 145.510 99.955 145.760 99.960 ;
        RECT 146.990 99.955 147.240 99.960 ;
        RECT 148.470 99.955 148.720 99.970 ;
        RECT 149.950 99.955 150.200 99.970 ;
        RECT 151.370 99.960 153.200 102.090 ;
        RECT 151.430 99.955 151.680 99.960 ;
        RECT 152.910 99.955 153.160 99.960 ;
        RECT 154.340 99.950 156.170 102.080 ;
        RECT 157.270 99.980 158.460 103.930 ;
        RECT 157.350 99.955 157.600 99.980 ;
        RECT 135.150 99.340 135.400 99.365 ;
        RECT 136.630 99.340 136.880 99.365 ;
        RECT 135.100 99.300 136.910 99.340 ;
        RECT 135.100 97.270 136.940 99.300 ;
        RECT 138.090 97.270 139.910 99.370 ;
        RECT 141.030 97.280 142.850 99.380 ;
        RECT 144.030 99.360 144.280 99.365 ;
        RECT 145.510 99.360 145.760 99.365 ;
        RECT 135.100 97.240 136.910 97.270 ;
        RECT 138.110 97.260 138.360 97.270 ;
        RECT 139.590 97.260 139.840 97.270 ;
        RECT 141.070 97.260 141.320 97.280 ;
        RECT 142.550 97.260 142.800 97.280 ;
        RECT 143.960 97.230 145.790 99.360 ;
        RECT 146.940 97.240 148.770 99.370 ;
        RECT 149.930 97.240 151.760 99.370 ;
        RECT 152.910 99.360 153.160 99.365 ;
        RECT 154.390 99.360 154.640 99.365 ;
        RECT 152.850 97.230 154.680 99.360 ;
        RECT 155.820 97.240 157.650 99.370 ;
        RECT 80.265 88.235 80.555 88.465 ;
        RECT 84.850 88.420 85.170 88.480 ;
        RECT 80.800 88.280 85.170 88.420 ;
        RECT 71.140 87.940 74.500 88.080 ;
        RECT 78.885 88.080 79.175 88.125 ;
        RECT 80.800 88.080 80.940 88.280 ;
        RECT 84.850 88.220 85.170 88.280 ;
        RECT 78.885 87.940 80.940 88.080 ;
        RECT 73.810 87.880 74.130 87.940 ;
        RECT 78.885 87.895 79.175 87.940 ;
        RECT 81.185 87.895 81.475 88.125 ;
        RECT 82.065 88.080 82.355 88.125 ;
        RECT 83.255 88.080 83.545 88.125 ;
        RECT 85.775 88.080 86.065 88.125 ;
        RECT 82.065 87.940 86.065 88.080 ;
        RECT 82.065 87.895 82.355 87.940 ;
        RECT 83.255 87.895 83.545 87.940 ;
        RECT 85.775 87.895 86.065 87.940 ;
        RECT 74.745 87.740 75.035 87.785 ;
        RECT 77.030 87.740 77.350 87.800 ;
        RECT 70.680 87.600 74.500 87.740 ;
        RECT 21.370 87.260 28.960 87.400 ;
        RECT 29.190 87.400 29.510 87.460 ;
        RECT 31.030 87.400 31.350 87.460 ;
        RECT 29.190 87.260 31.350 87.400 ;
        RECT 21.370 87.200 21.690 87.260 ;
        RECT 29.190 87.200 29.510 87.260 ;
        RECT 31.030 87.200 31.350 87.260 ;
        RECT 32.425 87.400 32.715 87.445 ;
        RECT 34.710 87.400 35.030 87.460 ;
        RECT 32.425 87.260 35.030 87.400 ;
        RECT 32.425 87.215 32.715 87.260 ;
        RECT 34.710 87.200 35.030 87.260 ;
        RECT 35.630 87.200 35.950 87.460 ;
        RECT 41.700 87.445 41.840 87.600 ;
        RECT 44.845 87.555 45.135 87.600 ;
        RECT 41.625 87.215 41.915 87.445 ;
        RECT 42.530 87.200 42.850 87.460 ;
        RECT 51.270 87.200 51.590 87.460 ;
        RECT 54.580 87.400 54.720 87.600 ;
        RECT 56.330 87.400 56.650 87.460 ;
        RECT 54.580 87.260 56.650 87.400 ;
        RECT 56.330 87.200 56.650 87.260 ;
        RECT 56.790 87.200 57.110 87.460 ;
        RECT 58.170 87.200 58.490 87.460 ;
        RECT 58.720 87.400 58.860 87.600 ;
        RECT 63.230 87.540 63.550 87.600 ;
        RECT 59.105 87.400 59.395 87.445 ;
        RECT 58.720 87.260 59.395 87.400 ;
        RECT 59.105 87.215 59.395 87.260 ;
        RECT 60.470 87.400 60.790 87.460 ;
        RECT 62.325 87.400 62.615 87.445 ;
        RECT 60.470 87.260 62.615 87.400 ;
        RECT 60.470 87.200 60.790 87.260 ;
        RECT 62.325 87.215 62.615 87.260 ;
        RECT 65.070 87.200 65.390 87.460 ;
        RECT 72.430 87.200 72.750 87.460 ;
        RECT 74.360 87.400 74.500 87.600 ;
        RECT 74.745 87.600 77.350 87.740 ;
        RECT 74.745 87.555 75.035 87.600 ;
        RECT 77.030 87.540 77.350 87.600 ;
        RECT 79.330 87.740 79.650 87.800 ;
        RECT 81.260 87.740 81.400 87.895 ;
        RECT 79.330 87.600 81.400 87.740 ;
        RECT 81.670 87.740 81.960 87.785 ;
        RECT 83.770 87.740 84.060 87.785 ;
        RECT 85.340 87.740 85.630 87.785 ;
        RECT 81.670 87.600 85.630 87.740 ;
        RECT 99.980 87.685 113.700 88.550 ;
        RECT 99.980 87.645 113.630 87.685 ;
        RECT 99.980 87.615 112.880 87.645 ;
        RECT 79.330 87.540 79.650 87.600 ;
        RECT 81.670 87.555 81.960 87.600 ;
        RECT 83.770 87.555 84.060 87.600 ;
        RECT 85.340 87.555 85.630 87.600 ;
        RECT 100.000 87.575 112.880 87.615 ;
        RECT 85.770 87.400 86.090 87.460 ;
        RECT 86.690 87.400 87.010 87.460 ;
        RECT 88.085 87.400 88.375 87.445 ;
        RECT 74.360 87.260 88.375 87.400 ;
        RECT 85.770 87.200 86.090 87.260 ;
        RECT 86.690 87.200 87.010 87.260 ;
        RECT 88.085 87.215 88.375 87.260 ;
        RECT 12.100 86.580 89.840 87.060 ;
        RECT 14.485 86.380 14.775 86.425 ;
        RECT 14.930 86.380 15.250 86.440 ;
        RECT 14.485 86.240 15.250 86.380 ;
        RECT 14.485 86.195 14.775 86.240 ;
        RECT 14.930 86.180 15.250 86.240 ;
        RECT 15.390 86.380 15.710 86.440 ;
        RECT 19.990 86.380 20.310 86.440 ;
        RECT 15.390 86.240 20.310 86.380 ;
        RECT 15.390 86.180 15.710 86.240 ;
        RECT 19.990 86.180 20.310 86.240 ;
        RECT 20.465 86.380 20.755 86.425 ;
        RECT 23.685 86.380 23.975 86.425 ;
        RECT 25.970 86.380 26.290 86.440 ;
        RECT 20.465 86.240 21.980 86.380 ;
        RECT 20.465 86.195 20.755 86.240 ;
        RECT 21.840 86.100 21.980 86.240 ;
        RECT 23.685 86.240 26.290 86.380 ;
        RECT 23.685 86.195 23.975 86.240 ;
        RECT 25.970 86.180 26.290 86.240 ;
        RECT 29.650 86.380 29.970 86.440 ;
        RECT 30.125 86.380 30.415 86.425 ;
        RECT 29.650 86.240 30.415 86.380 ;
        RECT 29.650 86.180 29.970 86.240 ;
        RECT 30.125 86.195 30.415 86.240 ;
        RECT 30.570 86.180 30.890 86.440 ;
        RECT 33.330 86.380 33.650 86.440 ;
        RECT 33.805 86.380 34.095 86.425 ;
        RECT 33.330 86.240 34.095 86.380 ;
        RECT 33.330 86.180 33.650 86.240 ;
        RECT 33.805 86.195 34.095 86.240 ;
        RECT 34.710 86.380 35.030 86.440 ;
        RECT 37.930 86.380 38.250 86.440 ;
        RECT 34.710 86.240 38.250 86.380 ;
        RECT 34.710 86.180 35.030 86.240 ;
        RECT 37.930 86.180 38.250 86.240 ;
        RECT 39.785 86.380 40.075 86.425 ;
        RECT 41.150 86.380 41.470 86.440 ;
        RECT 43.450 86.380 43.770 86.440 ;
        RECT 39.785 86.240 43.770 86.380 ;
        RECT 39.785 86.195 40.075 86.240 ;
        RECT 41.150 86.180 41.470 86.240 ;
        RECT 43.450 86.180 43.770 86.240 ;
        RECT 47.145 86.380 47.435 86.425 ;
        RECT 47.590 86.380 47.910 86.440 ;
        RECT 47.145 86.240 47.910 86.380 ;
        RECT 47.145 86.195 47.435 86.240 ;
        RECT 47.590 86.180 47.910 86.240 ;
        RECT 48.065 86.380 48.355 86.425 ;
        RECT 49.430 86.380 49.750 86.440 ;
        RECT 54.950 86.380 55.270 86.440 ;
        RECT 48.065 86.240 49.750 86.380 ;
        RECT 48.065 86.195 48.355 86.240 ;
        RECT 49.430 86.180 49.750 86.240 ;
        RECT 50.440 86.240 55.270 86.380 ;
        RECT 21.385 85.855 21.675 86.085 ;
        RECT 17.245 85.700 17.535 85.745 ;
        RECT 20.450 85.700 20.770 85.760 ;
        RECT 17.245 85.560 20.770 85.700 ;
        RECT 21.460 85.700 21.600 85.855 ;
        RECT 21.830 85.840 22.150 86.100 ;
        RECT 24.590 86.040 24.910 86.100 ;
        RECT 29.205 86.040 29.495 86.085 ;
        RECT 30.660 86.040 30.800 86.180 ;
        RECT 42.530 86.040 42.820 86.085 ;
        RECT 44.100 86.040 44.390 86.085 ;
        RECT 46.200 86.040 46.490 86.085 ;
        RECT 24.590 85.900 27.120 86.040 ;
        RECT 24.590 85.840 24.910 85.900 ;
        RECT 23.210 85.700 23.530 85.760 ;
        RECT 26.980 85.700 27.120 85.900 ;
        RECT 29.205 85.900 30.800 86.040 ;
        RECT 33.880 85.900 38.620 86.040 ;
        RECT 29.205 85.855 29.495 85.900 ;
        RECT 33.880 85.760 34.020 85.900 ;
        RECT 30.125 85.700 30.415 85.745 ;
        RECT 21.460 85.560 26.660 85.700 ;
        RECT 26.980 85.560 30.415 85.700 ;
        RECT 17.245 85.515 17.535 85.560 ;
        RECT 20.450 85.500 20.770 85.560 ;
        RECT 23.210 85.500 23.530 85.560 ;
        RECT 18.625 85.175 18.915 85.405 ;
        RECT 20.005 85.360 20.295 85.405 ;
        RECT 20.910 85.360 21.230 85.420 ;
        RECT 20.005 85.220 21.230 85.360 ;
        RECT 20.005 85.175 20.295 85.220 ;
        RECT 15.405 85.020 15.695 85.065 ;
        RECT 16.310 85.020 16.630 85.080 ;
        RECT 15.405 84.880 16.630 85.020 ;
        RECT 18.700 85.020 18.840 85.175 ;
        RECT 20.910 85.160 21.230 85.220 ;
        RECT 23.670 85.360 23.990 85.420 ;
        RECT 25.525 85.360 25.815 85.405 ;
        RECT 23.670 85.220 25.815 85.360 ;
        RECT 23.670 85.160 23.990 85.220 ;
        RECT 25.525 85.175 25.815 85.220 ;
        RECT 25.970 85.160 26.290 85.420 ;
        RECT 26.520 85.405 26.660 85.560 ;
        RECT 30.125 85.515 30.415 85.560 ;
        RECT 30.570 85.700 30.890 85.760 ;
        RECT 30.570 85.560 33.100 85.700 ;
        RECT 30.570 85.500 30.890 85.560 ;
        RECT 26.445 85.175 26.735 85.405 ;
        RECT 26.890 85.160 27.210 85.420 ;
        RECT 27.365 85.175 27.655 85.405 ;
        RECT 25.050 85.020 25.370 85.080 ;
        RECT 18.700 84.880 25.370 85.020 ;
        RECT 26.060 85.020 26.200 85.160 ;
        RECT 27.440 85.020 27.580 85.175 ;
        RECT 31.030 85.160 31.350 85.420 ;
        RECT 31.490 85.160 31.810 85.420 ;
        RECT 32.410 85.160 32.730 85.420 ;
        RECT 32.960 85.360 33.100 85.560 ;
        RECT 33.790 85.500 34.110 85.760 ;
        RECT 34.340 85.700 35.400 85.740 ;
        RECT 34.340 85.600 36.785 85.700 ;
        RECT 34.340 85.360 34.480 85.600 ;
        RECT 35.260 85.560 36.785 85.600 ;
        RECT 32.960 85.220 34.480 85.360 ;
        RECT 34.710 85.160 35.030 85.420 ;
        RECT 36.090 85.160 36.410 85.420 ;
        RECT 36.645 85.405 36.785 85.560 ;
        RECT 36.570 85.175 36.860 85.405 ;
        RECT 37.930 85.160 38.250 85.420 ;
        RECT 38.480 85.405 38.620 85.900 ;
        RECT 42.530 85.900 46.490 86.040 ;
        RECT 42.530 85.855 42.820 85.900 ;
        RECT 44.100 85.855 44.390 85.900 ;
        RECT 46.200 85.855 46.490 85.900 ;
        RECT 42.095 85.700 42.385 85.745 ;
        RECT 44.615 85.700 44.905 85.745 ;
        RECT 45.805 85.700 46.095 85.745 ;
        RECT 42.095 85.560 46.095 85.700 ;
        RECT 42.095 85.515 42.385 85.560 ;
        RECT 44.615 85.515 44.905 85.560 ;
        RECT 45.805 85.515 46.095 85.560 ;
        RECT 46.685 85.700 46.975 85.745 ;
        RECT 47.130 85.700 47.450 85.760 ;
        RECT 46.685 85.560 47.450 85.700 ;
        RECT 46.685 85.515 46.975 85.560 ;
        RECT 47.130 85.500 47.450 85.560 ;
        RECT 38.430 85.175 38.720 85.405 ;
        RECT 42.530 85.360 42.850 85.420 ;
        RECT 45.350 85.360 45.640 85.405 ;
        RECT 42.530 85.220 45.640 85.360 ;
        RECT 42.530 85.160 42.850 85.220 ;
        RECT 45.350 85.175 45.640 85.220 ;
        RECT 48.510 85.360 48.830 85.420 ;
        RECT 49.905 85.360 50.195 85.405 ;
        RECT 48.510 85.220 50.195 85.360 ;
        RECT 50.440 85.360 50.580 86.240 ;
        RECT 54.950 86.180 55.270 86.240 ;
        RECT 55.410 86.180 55.730 86.440 ;
        RECT 56.330 86.380 56.650 86.440 ;
        RECT 59.090 86.380 59.410 86.440 ;
        RECT 71.525 86.380 71.815 86.425 ;
        RECT 56.330 86.240 59.410 86.380 ;
        RECT 56.330 86.180 56.650 86.240 ;
        RECT 59.090 86.180 59.410 86.240 ;
        RECT 67.000 86.240 71.815 86.380 ;
        RECT 52.205 86.040 52.495 86.085 ;
        RECT 59.550 86.040 59.870 86.100 ;
        RECT 60.930 86.040 61.250 86.100 ;
        RECT 65.070 86.040 65.390 86.100 ;
        RECT 52.205 85.900 61.250 86.040 ;
        RECT 52.205 85.855 52.495 85.900 ;
        RECT 59.550 85.840 59.870 85.900 ;
        RECT 60.930 85.840 61.250 85.900 ;
        RECT 63.320 85.900 65.390 86.040 ;
        RECT 50.810 85.700 51.130 85.760 ;
        RECT 50.810 85.645 52.420 85.700 ;
        RECT 52.665 85.645 52.955 85.745 ;
        RECT 53.810 85.700 54.720 85.740 ;
        RECT 60.470 85.700 60.790 85.760 ;
        RECT 50.810 85.560 52.955 85.645 ;
        RECT 50.810 85.500 51.130 85.560 ;
        RECT 52.280 85.515 52.955 85.560 ;
        RECT 53.330 85.600 60.790 85.700 ;
        RECT 53.330 85.560 53.950 85.600 ;
        RECT 54.580 85.560 60.790 85.600 ;
        RECT 52.280 85.505 52.880 85.515 ;
        RECT 51.285 85.360 51.575 85.405 ;
        RECT 50.440 85.220 51.575 85.360 ;
        RECT 48.510 85.160 48.830 85.220 ;
        RECT 49.905 85.175 50.195 85.220 ;
        RECT 51.285 85.175 51.575 85.220 ;
        RECT 51.745 85.360 52.035 85.405 ;
        RECT 53.330 85.360 53.470 85.560 ;
        RECT 60.470 85.500 60.790 85.560 ;
        RECT 54.030 85.360 54.350 85.420 ;
        RECT 51.745 85.220 53.470 85.360 ;
        RECT 53.840 85.220 54.350 85.360 ;
        RECT 51.745 85.175 52.035 85.220 ;
        RECT 54.030 85.160 54.350 85.220 ;
        RECT 54.735 85.175 55.025 85.405 ;
        RECT 55.410 85.360 55.730 85.420 ;
        RECT 55.885 85.360 56.175 85.405 ;
        RECT 55.410 85.220 56.175 85.360 ;
        RECT 26.060 84.880 27.580 85.020 ;
        RECT 15.405 84.835 15.695 84.880 ;
        RECT 16.310 84.820 16.630 84.880 ;
        RECT 25.050 84.820 25.370 84.880 ;
        RECT 35.630 84.820 35.950 85.080 ;
        RECT 37.470 84.820 37.790 85.080 ;
        RECT 54.810 85.020 54.950 85.175 ;
        RECT 55.410 85.160 55.730 85.220 ;
        RECT 55.885 85.175 56.175 85.220 ;
        RECT 56.330 85.160 56.650 85.420 ;
        RECT 56.805 85.360 57.095 85.405 ;
        RECT 57.250 85.360 57.570 85.420 ;
        RECT 56.805 85.220 57.570 85.360 ;
        RECT 56.805 85.175 57.095 85.220 ;
        RECT 57.250 85.160 57.570 85.220 ;
        RECT 57.725 85.360 58.015 85.405 ;
        RECT 58.170 85.360 58.490 85.420 ;
        RECT 57.725 85.220 58.490 85.360 ;
        RECT 57.725 85.175 58.015 85.220 ;
        RECT 58.170 85.160 58.490 85.220 ;
        RECT 58.630 85.160 58.950 85.420 ;
        RECT 59.090 85.160 59.410 85.420 ;
        RECT 59.550 85.160 59.870 85.420 ;
        RECT 61.390 85.360 61.710 85.420 ;
        RECT 63.320 85.405 63.460 85.900 ;
        RECT 65.070 85.840 65.390 85.900 ;
        RECT 64.165 85.700 64.455 85.745 ;
        RECT 65.990 85.700 66.310 85.760 ;
        RECT 64.165 85.560 66.310 85.700 ;
        RECT 64.165 85.515 64.455 85.560 ;
        RECT 65.990 85.500 66.310 85.560 ;
        RECT 62.325 85.360 62.615 85.405 ;
        RECT 61.390 85.220 62.615 85.360 ;
        RECT 61.390 85.160 61.710 85.220 ;
        RECT 62.325 85.175 62.615 85.220 ;
        RECT 63.245 85.175 63.535 85.405 ;
        RECT 63.705 85.175 63.995 85.405 ;
        RECT 65.085 85.360 65.375 85.405 ;
        RECT 65.530 85.360 65.850 85.420 ;
        RECT 65.085 85.220 65.850 85.360 ;
        RECT 65.085 85.175 65.375 85.220 ;
        RECT 61.480 85.020 61.620 85.160 ;
        RECT 54.810 84.880 55.640 85.020 ;
        RECT 55.500 84.740 55.640 84.880 ;
        RECT 60.100 84.880 61.620 85.020 ;
        RECT 22.290 84.680 22.610 84.740 ;
        RECT 23.685 84.680 23.975 84.725 ;
        RECT 22.290 84.540 23.975 84.680 ;
        RECT 22.290 84.480 22.610 84.540 ;
        RECT 23.685 84.495 23.975 84.540 ;
        RECT 24.605 84.680 24.895 84.725 ;
        RECT 25.970 84.680 26.290 84.740 ;
        RECT 24.605 84.540 26.290 84.680 ;
        RECT 24.605 84.495 24.895 84.540 ;
        RECT 25.970 84.480 26.290 84.540 ;
        RECT 26.430 84.680 26.750 84.740 ;
        RECT 28.745 84.680 29.035 84.725 ;
        RECT 26.430 84.540 29.035 84.680 ;
        RECT 26.430 84.480 26.750 84.540 ;
        RECT 28.745 84.495 29.035 84.540 ;
        RECT 32.425 84.680 32.715 84.725 ;
        RECT 38.390 84.680 38.710 84.740 ;
        RECT 32.425 84.540 38.710 84.680 ;
        RECT 32.425 84.495 32.715 84.540 ;
        RECT 38.390 84.480 38.710 84.540 ;
        RECT 39.310 84.480 39.630 84.740 ;
        RECT 48.050 84.480 48.370 84.740 ;
        RECT 53.110 84.480 53.430 84.740 ;
        RECT 55.410 84.480 55.730 84.740 ;
        RECT 58.170 84.680 58.490 84.740 ;
        RECT 60.100 84.680 60.240 84.880 ;
        RECT 58.170 84.540 60.240 84.680 ;
        RECT 60.945 84.680 61.235 84.725 ;
        RECT 61.390 84.680 61.710 84.740 ;
        RECT 60.945 84.540 61.710 84.680 ;
        RECT 58.170 84.480 58.490 84.540 ;
        RECT 60.945 84.495 61.235 84.540 ;
        RECT 61.390 84.480 61.710 84.540 ;
        RECT 63.230 84.680 63.550 84.740 ;
        RECT 63.780 84.680 63.920 85.175 ;
        RECT 65.530 85.160 65.850 85.220 ;
        RECT 66.465 85.360 66.755 85.405 ;
        RECT 67.000 85.360 67.140 86.240 ;
        RECT 71.525 86.195 71.815 86.240 ;
        RECT 73.825 86.380 74.115 86.425 ;
        RECT 76.570 86.380 76.890 86.440 ;
        RECT 77.965 86.380 78.255 86.425 ;
        RECT 73.825 86.240 78.255 86.380 ;
        RECT 73.825 86.195 74.115 86.240 ;
        RECT 76.570 86.180 76.890 86.240 ;
        RECT 77.965 86.195 78.255 86.240 ;
        RECT 78.885 86.380 79.175 86.425 ;
        RECT 79.790 86.380 80.110 86.440 ;
        RECT 78.885 86.240 80.110 86.380 ;
        RECT 78.885 86.195 79.175 86.240 ;
        RECT 79.790 86.180 80.110 86.240 ;
        RECT 80.265 86.380 80.555 86.425 ;
        RECT 80.710 86.380 81.030 86.440 ;
        RECT 80.265 86.240 81.030 86.380 ;
        RECT 80.265 86.195 80.555 86.240 ;
        RECT 80.710 86.180 81.030 86.240 ;
        RECT 75.190 86.040 75.510 86.100 ;
        RECT 82.105 86.040 82.395 86.085 ;
        RECT 75.190 85.900 82.395 86.040 ;
        RECT 75.190 85.840 75.510 85.900 ;
        RECT 82.105 85.855 82.395 85.900 ;
        RECT 85.325 85.855 85.615 86.085 ;
        RECT 81.630 85.700 81.950 85.760 ;
        RECT 81.630 85.560 83.700 85.700 ;
        RECT 81.630 85.500 81.950 85.560 ;
        RECT 66.465 85.220 67.140 85.360 ;
        RECT 66.465 85.175 66.755 85.220 ;
        RECT 68.290 85.160 68.610 85.420 ;
        RECT 69.210 85.360 69.530 85.420 ;
        RECT 69.685 85.360 69.975 85.405 ;
        RECT 77.490 85.360 77.810 85.420 ;
        RECT 79.805 85.360 80.095 85.405 ;
        RECT 69.210 85.220 69.975 85.360 ;
        RECT 69.210 85.160 69.530 85.220 ;
        RECT 69.685 85.175 69.975 85.220 ;
        RECT 72.980 85.220 77.260 85.360 ;
        RECT 72.980 85.080 73.120 85.220 ;
        RECT 64.610 85.020 64.930 85.080 ;
        RECT 67.385 85.020 67.675 85.065 ;
        RECT 64.610 84.880 67.675 85.020 ;
        RECT 64.610 84.820 64.930 84.880 ;
        RECT 67.385 84.835 67.675 84.880 ;
        RECT 67.845 85.020 68.135 85.065 ;
        RECT 70.605 85.020 70.895 85.065 ;
        RECT 71.050 85.020 71.370 85.080 ;
        RECT 67.845 84.880 69.900 85.020 ;
        RECT 67.845 84.835 68.135 84.880 ;
        RECT 69.760 84.740 69.900 84.880 ;
        RECT 70.605 84.880 71.370 85.020 ;
        RECT 70.605 84.835 70.895 84.880 ;
        RECT 71.050 84.820 71.370 84.880 ;
        RECT 72.890 84.820 73.210 85.080 ;
        RECT 73.350 85.020 73.670 85.080 ;
        RECT 77.120 85.065 77.260 85.220 ;
        RECT 77.490 85.220 80.095 85.360 ;
        RECT 77.490 85.160 77.810 85.220 ;
        RECT 79.805 85.175 80.095 85.220 ;
        RECT 81.170 85.160 81.490 85.420 ;
        RECT 83.010 85.160 83.330 85.420 ;
        RECT 83.560 85.405 83.700 85.560 ;
        RECT 83.485 85.175 83.775 85.405 ;
        RECT 84.390 85.160 84.710 85.420 ;
        RECT 84.865 85.360 85.155 85.405 ;
        RECT 85.400 85.360 85.540 85.855 ;
        RECT 84.865 85.220 85.540 85.360 ;
        RECT 84.865 85.175 85.155 85.220 ;
        RECT 86.245 85.175 86.535 85.405 ;
        RECT 73.825 85.020 74.115 85.065 ;
        RECT 73.350 84.880 74.115 85.020 ;
        RECT 73.350 84.820 73.670 84.880 ;
        RECT 73.825 84.835 74.115 84.880 ;
        RECT 77.045 84.835 77.335 85.065 ;
        RECT 86.320 85.020 86.460 85.175 ;
        RECT 86.690 85.160 87.010 85.420 ;
        RECT 87.150 85.160 87.470 85.420 ;
        RECT 88.085 85.360 88.375 85.405 ;
        RECT 88.530 85.360 88.850 85.420 ;
        RECT 88.085 85.220 88.850 85.360 ;
        RECT 88.085 85.175 88.375 85.220 ;
        RECT 88.530 85.160 88.850 85.220 ;
        RECT 79.880 84.880 86.460 85.020 ;
        RECT 100.540 84.895 101.150 87.235 ;
        RECT 101.980 87.045 102.640 87.365 ;
        RECT 102.030 84.925 102.640 87.045 ;
        RECT 102.480 84.895 102.640 84.925 ;
        RECT 103.500 84.885 104.050 87.235 ;
        RECT 79.880 84.740 80.020 84.880 ;
        RECT 105.010 84.865 105.560 87.215 ;
        RECT 106.470 84.895 107.020 87.245 ;
        RECT 107.950 84.925 108.500 87.275 ;
        RECT 109.400 84.915 109.950 87.265 ;
        RECT 110.900 84.925 111.450 87.275 ;
        RECT 112.320 87.135 112.880 87.575 ;
        RECT 112.320 84.975 112.890 87.135 ;
        RECT 112.320 84.965 112.880 84.975 ;
        RECT 64.150 84.680 64.470 84.740 ;
        RECT 63.230 84.540 64.470 84.680 ;
        RECT 63.230 84.480 63.550 84.540 ;
        RECT 64.150 84.480 64.470 84.540 ;
        RECT 66.005 84.680 66.295 84.725 ;
        RECT 66.910 84.680 67.230 84.740 ;
        RECT 66.005 84.540 67.230 84.680 ;
        RECT 66.005 84.495 66.295 84.540 ;
        RECT 66.910 84.480 67.230 84.540 ;
        RECT 69.210 84.480 69.530 84.740 ;
        RECT 69.670 84.480 69.990 84.740 ;
        RECT 71.510 84.680 71.830 84.740 ;
        RECT 74.745 84.680 75.035 84.725 ;
        RECT 71.510 84.540 75.035 84.680 ;
        RECT 71.510 84.480 71.830 84.540 ;
        RECT 74.745 84.495 75.035 84.540 ;
        RECT 75.650 84.680 75.970 84.740 ;
        RECT 77.965 84.680 78.255 84.725 ;
        RECT 78.410 84.680 78.730 84.740 ;
        RECT 75.650 84.540 78.730 84.680 ;
        RECT 75.650 84.480 75.970 84.540 ;
        RECT 77.965 84.495 78.255 84.540 ;
        RECT 78.410 84.480 78.730 84.540 ;
        RECT 79.790 84.480 80.110 84.740 ;
        RECT 12.100 83.860 89.840 84.340 ;
        RECT 14.470 83.660 14.790 83.720 ;
        RECT 16.785 83.660 17.075 83.705 ;
        RECT 14.470 83.520 17.075 83.660 ;
        RECT 14.470 83.460 14.790 83.520 ;
        RECT 16.785 83.475 17.075 83.520 ;
        RECT 18.610 83.660 18.930 83.720 ;
        RECT 19.545 83.660 19.835 83.705 ;
        RECT 18.610 83.520 19.835 83.660 ;
        RECT 18.610 83.460 18.930 83.520 ;
        RECT 19.545 83.475 19.835 83.520 ;
        RECT 25.050 83.660 25.370 83.720 ;
        RECT 31.030 83.660 31.350 83.720 ;
        RECT 25.050 83.520 31.350 83.660 ;
        RECT 25.050 83.460 25.370 83.520 ;
        RECT 31.030 83.460 31.350 83.520 ;
        RECT 35.170 83.460 35.490 83.720 ;
        RECT 37.470 83.460 37.790 83.720 ;
        RECT 41.150 83.660 41.470 83.720 ;
        RECT 38.480 83.520 41.470 83.660 ;
        RECT 31.965 83.320 32.255 83.365 ;
        RECT 33.790 83.320 34.110 83.380 ;
        RECT 31.965 83.180 34.110 83.320 ;
        RECT 31.965 83.135 32.255 83.180 ;
        RECT 33.790 83.120 34.110 83.180 ;
        RECT 35.645 83.320 35.935 83.365 ;
        RECT 38.480 83.320 38.620 83.520 ;
        RECT 41.150 83.460 41.470 83.520 ;
        RECT 45.765 83.660 46.055 83.705 ;
        RECT 48.050 83.660 48.370 83.720 ;
        RECT 45.765 83.520 48.370 83.660 ;
        RECT 45.765 83.475 46.055 83.520 ;
        RECT 48.050 83.460 48.370 83.520 ;
        RECT 54.505 83.660 54.795 83.705 ;
        RECT 55.870 83.660 56.190 83.720 ;
        RECT 59.565 83.660 59.855 83.705 ;
        RECT 60.010 83.660 60.330 83.720 ;
        RECT 54.505 83.520 56.190 83.660 ;
        RECT 54.505 83.475 54.795 83.520 ;
        RECT 55.870 83.460 56.190 83.520 ;
        RECT 56.420 83.520 60.330 83.660 ;
        RECT 51.270 83.320 51.590 83.380 ;
        RECT 56.420 83.365 56.560 83.520 ;
        RECT 59.565 83.475 59.855 83.520 ;
        RECT 60.010 83.460 60.330 83.520 ;
        RECT 60.470 83.460 60.790 83.720 ;
        RECT 60.930 83.460 61.250 83.720 ;
        RECT 61.850 83.660 62.170 83.720 ;
        RECT 65.530 83.660 65.850 83.720 ;
        RECT 99.980 83.715 100.370 83.725 ;
        RECT 61.850 83.520 65.850 83.660 ;
        RECT 61.850 83.460 62.170 83.520 ;
        RECT 65.530 83.460 65.850 83.520 ;
        RECT 66.925 83.660 67.215 83.705 ;
        RECT 69.685 83.660 69.975 83.705 ;
        RECT 66.925 83.520 69.975 83.660 ;
        RECT 66.925 83.475 67.215 83.520 ;
        RECT 69.685 83.475 69.975 83.520 ;
        RECT 77.505 83.660 77.795 83.705 ;
        RECT 77.505 83.520 87.840 83.660 ;
        RECT 77.505 83.475 77.795 83.520 ;
        RECT 35.645 83.180 38.620 83.320 ;
        RECT 38.940 83.180 47.360 83.320 ;
        RECT 35.645 83.135 35.935 83.180 ;
        RECT 16.325 82.980 16.615 83.025 ;
        RECT 16.770 82.980 17.090 83.040 ;
        RECT 16.325 82.840 17.090 82.980 ;
        RECT 16.325 82.795 16.615 82.840 ;
        RECT 16.770 82.780 17.090 82.840 ;
        RECT 17.230 82.780 17.550 83.040 ;
        RECT 19.070 82.780 19.390 83.040 ;
        RECT 20.005 82.980 20.295 83.025 ;
        RECT 30.110 82.980 30.430 83.040 ;
        RECT 20.005 82.840 30.430 82.980 ;
        RECT 20.005 82.795 20.295 82.840 ;
        RECT 30.110 82.780 30.430 82.840 ;
        RECT 32.410 82.980 32.730 83.040 ;
        RECT 32.885 82.980 33.175 83.025 ;
        RECT 32.410 82.840 33.175 82.980 ;
        RECT 32.410 82.780 32.730 82.840 ;
        RECT 32.885 82.795 33.175 82.840 ;
        RECT 34.250 82.780 34.570 83.040 ;
        RECT 33.345 82.640 33.635 82.685 ;
        RECT 35.720 82.640 35.860 83.135 ;
        RECT 36.550 82.780 36.870 83.040 ;
        RECT 38.940 83.025 39.080 83.180 ;
        RECT 47.220 83.040 47.360 83.180 ;
        RECT 51.270 83.180 56.100 83.320 ;
        RECT 51.270 83.120 51.590 83.180 ;
        RECT 38.865 82.795 39.155 83.025 ;
        RECT 40.145 82.980 40.435 83.025 ;
        RECT 39.400 82.840 40.435 82.980 ;
        RECT 33.345 82.500 35.860 82.640 ;
        RECT 38.390 82.640 38.710 82.700 ;
        RECT 39.400 82.640 39.540 82.840 ;
        RECT 40.145 82.795 40.435 82.840 ;
        RECT 47.130 82.980 47.450 83.040 ;
        RECT 55.960 83.025 56.100 83.180 ;
        RECT 56.345 83.135 56.635 83.365 ;
        RECT 56.805 83.320 57.095 83.365 ;
        RECT 59.090 83.320 59.410 83.380 ;
        RECT 60.560 83.320 60.700 83.460 ;
        RECT 56.805 83.180 60.700 83.320 ;
        RECT 61.020 83.320 61.160 83.460 ;
        RECT 87.700 83.380 87.840 83.520 ;
        RECT 63.690 83.320 64.010 83.380 ;
        RECT 61.020 83.180 62.540 83.320 ;
        RECT 56.805 83.135 57.095 83.180 ;
        RECT 59.090 83.120 59.410 83.180 ;
        RECT 47.605 82.980 47.895 83.025 ;
        RECT 47.130 82.840 47.895 82.980 ;
        RECT 47.130 82.780 47.450 82.840 ;
        RECT 47.605 82.795 47.895 82.840 ;
        RECT 48.940 82.980 49.230 83.025 ;
        RECT 54.965 82.980 55.255 83.025 ;
        RECT 48.940 82.840 55.255 82.980 ;
        RECT 48.940 82.795 49.230 82.840 ;
        RECT 54.965 82.795 55.255 82.840 ;
        RECT 55.885 82.795 56.175 83.025 ;
        RECT 57.395 82.980 57.685 83.025 ;
        RECT 57.340 82.795 57.685 82.980 ;
        RECT 58.645 82.795 58.935 83.025 ;
        RECT 38.390 82.500 39.540 82.640 ;
        RECT 39.745 82.640 40.035 82.685 ;
        RECT 40.935 82.640 41.225 82.685 ;
        RECT 43.455 82.640 43.745 82.685 ;
        RECT 39.745 82.500 43.745 82.640 ;
        RECT 33.345 82.455 33.635 82.500 ;
        RECT 38.390 82.440 38.710 82.500 ;
        RECT 39.745 82.455 40.035 82.500 ;
        RECT 40.935 82.455 41.225 82.500 ;
        RECT 43.455 82.455 43.745 82.500 ;
        RECT 48.485 82.640 48.775 82.685 ;
        RECT 49.675 82.640 49.965 82.685 ;
        RECT 52.195 82.640 52.485 82.685 ;
        RECT 48.485 82.500 52.485 82.640 ;
        RECT 48.485 82.455 48.775 82.500 ;
        RECT 49.675 82.455 49.965 82.500 ;
        RECT 52.195 82.455 52.485 82.500 ;
        RECT 52.650 82.640 52.970 82.700 ;
        RECT 57.340 82.640 57.480 82.795 ;
        RECT 52.650 82.500 57.480 82.640 ;
        RECT 58.185 82.640 58.475 82.685 ;
        RECT 58.720 82.640 58.860 82.795 ;
        RECT 59.550 82.780 59.870 83.040 ;
        RECT 60.025 82.980 60.315 83.025 ;
        RECT 60.470 82.980 60.790 83.040 ;
        RECT 60.025 82.840 60.790 82.980 ;
        RECT 60.025 82.795 60.315 82.840 ;
        RECT 60.470 82.780 60.790 82.840 ;
        RECT 60.945 82.795 61.235 83.025 ;
        RECT 61.405 82.795 61.695 83.025 ;
        RECT 61.020 82.640 61.160 82.795 ;
        RECT 58.185 82.500 58.860 82.640 ;
        RECT 59.180 82.500 61.160 82.640 ;
        RECT 52.650 82.440 52.970 82.500 ;
        RECT 58.185 82.455 58.475 82.500 ;
        RECT 39.350 82.300 39.640 82.345 ;
        RECT 41.450 82.300 41.740 82.345 ;
        RECT 43.020 82.300 43.310 82.345 ;
        RECT 39.350 82.160 43.310 82.300 ;
        RECT 39.350 82.115 39.640 82.160 ;
        RECT 41.450 82.115 41.740 82.160 ;
        RECT 43.020 82.115 43.310 82.160 ;
        RECT 48.090 82.300 48.380 82.345 ;
        RECT 50.190 82.300 50.480 82.345 ;
        RECT 51.760 82.300 52.050 82.345 ;
        RECT 48.090 82.160 52.050 82.300 ;
        RECT 48.090 82.115 48.380 82.160 ;
        RECT 50.190 82.115 50.480 82.160 ;
        RECT 51.760 82.115 52.050 82.160 ;
        RECT 55.870 82.300 56.190 82.360 ;
        RECT 57.250 82.300 57.570 82.360 ;
        RECT 58.260 82.300 58.400 82.455 ;
        RECT 55.870 82.160 58.400 82.300 ;
        RECT 58.630 82.300 58.950 82.360 ;
        RECT 59.180 82.300 59.320 82.500 ;
        RECT 58.630 82.160 59.320 82.300 ;
        RECT 60.930 82.300 61.250 82.360 ;
        RECT 61.480 82.300 61.620 82.795 ;
        RECT 61.850 82.780 62.170 83.040 ;
        RECT 62.400 82.980 62.540 83.180 ;
        RECT 63.690 83.180 79.100 83.320 ;
        RECT 63.690 83.120 64.010 83.180 ;
        RECT 78.960 83.040 79.100 83.180 ;
        RECT 80.340 83.180 84.160 83.320 ;
        RECT 80.340 83.040 80.480 83.180 ;
        RECT 64.165 82.980 64.455 83.025 ;
        RECT 62.400 82.840 64.455 82.980 ;
        RECT 64.165 82.795 64.455 82.840 ;
        RECT 65.070 82.780 65.390 83.040 ;
        RECT 65.530 82.780 65.850 83.040 ;
        RECT 66.005 82.980 66.295 83.025 ;
        RECT 68.290 82.980 68.610 83.040 ;
        RECT 66.005 82.840 68.610 82.980 ;
        RECT 66.005 82.795 66.295 82.840 ;
        RECT 64.610 82.640 64.930 82.700 ;
        RECT 66.080 82.640 66.220 82.795 ;
        RECT 68.290 82.780 68.610 82.840 ;
        RECT 69.225 82.980 69.515 83.025 ;
        RECT 71.525 82.980 71.815 83.025 ;
        RECT 69.225 82.840 71.815 82.980 ;
        RECT 69.225 82.795 69.515 82.840 ;
        RECT 71.525 82.795 71.815 82.840 ;
        RECT 76.585 82.980 76.875 83.025 ;
        RECT 77.030 82.980 77.350 83.040 ;
        RECT 76.585 82.840 77.350 82.980 ;
        RECT 76.585 82.795 76.875 82.840 ;
        RECT 77.030 82.780 77.350 82.840 ;
        RECT 78.870 82.980 79.190 83.040 ;
        RECT 79.805 82.980 80.095 83.025 ;
        RECT 78.870 82.840 80.095 82.980 ;
        RECT 78.870 82.780 79.190 82.840 ;
        RECT 79.805 82.795 80.095 82.840 ;
        RECT 64.610 82.500 66.220 82.640 ;
        RECT 66.910 82.640 67.230 82.700 ;
        RECT 66.910 82.500 69.440 82.640 ;
        RECT 64.610 82.440 64.930 82.500 ;
        RECT 66.910 82.440 67.230 82.500 ;
        RECT 60.930 82.160 61.620 82.300 ;
        RECT 63.245 82.300 63.535 82.345 ;
        RECT 68.750 82.300 69.070 82.360 ;
        RECT 63.245 82.160 69.070 82.300 ;
        RECT 69.300 82.300 69.440 82.500 ;
        RECT 70.145 82.455 70.435 82.685 ;
        RECT 72.890 82.640 73.210 82.700 ;
        RECT 74.285 82.640 74.575 82.685 ;
        RECT 72.890 82.500 74.575 82.640 ;
        RECT 70.220 82.300 70.360 82.455 ;
        RECT 72.890 82.440 73.210 82.500 ;
        RECT 74.285 82.455 74.575 82.500 ;
        RECT 75.650 82.440 75.970 82.700 ;
        RECT 69.300 82.160 70.360 82.300 ;
        RECT 79.880 82.300 80.020 82.795 ;
        RECT 80.250 82.780 80.570 83.040 ;
        RECT 80.725 82.795 81.015 83.025 ;
        RECT 80.800 82.640 80.940 82.795 ;
        RECT 81.630 82.780 81.950 83.040 ;
        RECT 83.470 82.780 83.790 83.040 ;
        RECT 84.020 83.025 84.160 83.180 ;
        RECT 87.610 83.120 87.930 83.380 ;
        RECT 83.945 82.795 84.235 83.025 ;
        RECT 84.405 82.980 84.695 83.025 ;
        RECT 84.850 82.980 85.170 83.040 ;
        RECT 84.405 82.840 85.170 82.980 ;
        RECT 84.405 82.795 84.695 82.840 ;
        RECT 84.850 82.780 85.170 82.840 ;
        RECT 85.325 82.980 85.615 83.025 ;
        RECT 86.230 82.980 86.550 83.040 ;
        RECT 85.325 82.840 86.550 82.980 ;
        RECT 85.325 82.795 85.615 82.840 ;
        RECT 86.230 82.780 86.550 82.840 ;
        RECT 86.690 82.780 87.010 83.040 ;
        RECT 85.785 82.640 86.075 82.685 ;
        RECT 80.800 82.500 86.075 82.640 ;
        RECT 85.785 82.455 86.075 82.500 ;
        RECT 80.710 82.300 81.030 82.360 ;
        RECT 79.880 82.160 81.030 82.300 ;
        RECT 55.870 82.100 56.190 82.160 ;
        RECT 57.250 82.100 57.570 82.160 ;
        RECT 58.630 82.100 58.950 82.160 ;
        RECT 60.930 82.100 61.250 82.160 ;
        RECT 63.245 82.115 63.535 82.160 ;
        RECT 68.750 82.100 69.070 82.160 ;
        RECT 80.710 82.100 81.030 82.160 ;
        RECT 81.630 82.300 81.950 82.360 ;
        RECT 86.230 82.300 86.550 82.360 ;
        RECT 81.630 82.160 86.550 82.300 ;
        RECT 81.630 82.100 81.950 82.160 ;
        RECT 86.230 82.100 86.550 82.160 ;
        RECT 30.110 81.960 30.430 82.020 ;
        RECT 31.045 81.960 31.335 82.005 ;
        RECT 30.110 81.820 31.335 81.960 ;
        RECT 30.110 81.760 30.430 81.820 ;
        RECT 31.045 81.775 31.335 81.820 ;
        RECT 54.030 81.960 54.350 82.020 ;
        RECT 59.550 81.960 59.870 82.020 ;
        RECT 54.030 81.820 59.870 81.960 ;
        RECT 54.030 81.760 54.350 81.820 ;
        RECT 59.550 81.760 59.870 81.820 ;
        RECT 67.370 81.760 67.690 82.020 ;
        RECT 68.290 81.960 68.610 82.020 ;
        RECT 75.190 81.960 75.510 82.020 ;
        RECT 68.290 81.820 75.510 81.960 ;
        RECT 68.290 81.760 68.610 81.820 ;
        RECT 75.190 81.760 75.510 81.820 ;
        RECT 78.425 81.960 78.715 82.005 ;
        RECT 80.250 81.960 80.570 82.020 ;
        RECT 78.425 81.820 80.570 81.960 ;
        RECT 78.425 81.775 78.715 81.820 ;
        RECT 80.250 81.760 80.570 81.820 ;
        RECT 82.090 81.760 82.410 82.020 ;
        RECT 12.100 81.140 89.840 81.620 ;
        RECT 99.980 81.555 101.000 83.715 ;
        RECT 34.710 80.740 35.030 81.000 ;
        RECT 58.645 80.940 58.935 80.985 ;
        RECT 59.090 80.940 59.410 81.000 ;
        RECT 58.645 80.800 59.410 80.940 ;
        RECT 58.645 80.755 58.935 80.800 ;
        RECT 59.090 80.740 59.410 80.800 ;
        RECT 60.025 80.755 60.315 80.985 ;
        RECT 60.470 80.940 60.790 81.000 ;
        RECT 61.865 80.940 62.155 80.985 ;
        RECT 74.745 80.940 75.035 80.985 ;
        RECT 60.470 80.800 62.155 80.940 ;
        RECT 37.930 80.400 38.250 80.660 ;
        RECT 50.350 80.400 50.670 80.660 ;
        RECT 51.730 80.600 52.050 80.660 ;
        RECT 54.030 80.600 54.350 80.660 ;
        RECT 54.950 80.600 55.270 80.660 ;
        RECT 56.805 80.600 57.095 80.645 ;
        RECT 51.730 80.460 54.720 80.600 ;
        RECT 51.730 80.400 52.050 80.460 ;
        RECT 54.030 80.400 54.350 80.460 ;
        RECT 26.890 80.260 27.210 80.320 ;
        RECT 27.825 80.260 28.115 80.305 ;
        RECT 26.890 80.120 28.115 80.260 ;
        RECT 26.890 80.060 27.210 80.120 ;
        RECT 27.825 80.075 28.115 80.120 ;
        RECT 31.030 80.260 31.350 80.320 ;
        RECT 35.185 80.260 35.475 80.305 ;
        RECT 38.020 80.260 38.160 80.400 ;
        RECT 41.150 80.260 41.470 80.320 ;
        RECT 42.530 80.260 42.850 80.320 ;
        RECT 31.030 80.120 38.160 80.260 ;
        RECT 38.940 80.120 42.850 80.260 ;
        RECT 31.030 80.060 31.350 80.120 ;
        RECT 35.185 80.075 35.475 80.120 ;
        RECT 23.210 79.720 23.530 79.980 ;
        RECT 28.270 79.920 28.590 79.980 ;
        RECT 28.745 79.920 29.035 79.965 ;
        RECT 28.270 79.780 29.035 79.920 ;
        RECT 28.270 79.720 28.590 79.780 ;
        RECT 28.745 79.735 29.035 79.780 ;
        RECT 29.205 79.920 29.495 79.965 ;
        RECT 29.650 79.920 29.970 79.980 ;
        RECT 29.205 79.780 29.970 79.920 ;
        RECT 29.205 79.735 29.495 79.780 ;
        RECT 29.650 79.720 29.970 79.780 ;
        RECT 31.965 79.920 32.255 79.965 ;
        RECT 32.870 79.920 33.190 79.980 ;
        RECT 31.965 79.780 33.190 79.920 ;
        RECT 31.965 79.735 32.255 79.780 ;
        RECT 32.870 79.720 33.190 79.780 ;
        RECT 33.790 79.720 34.110 79.980 ;
        RECT 36.565 79.920 36.855 79.965 ;
        RECT 37.010 79.920 37.330 79.980 ;
        RECT 36.565 79.780 37.330 79.920 ;
        RECT 36.565 79.735 36.855 79.780 ;
        RECT 37.010 79.720 37.330 79.780 ;
        RECT 37.470 79.720 37.790 79.980 ;
        RECT 37.945 79.920 38.235 79.965 ;
        RECT 38.390 79.920 38.710 79.980 ;
        RECT 38.940 79.965 39.080 80.120 ;
        RECT 41.150 80.060 41.470 80.120 ;
        RECT 42.530 80.060 42.850 80.120 ;
        RECT 52.650 80.260 52.970 80.320 ;
        RECT 54.580 80.305 54.720 80.460 ;
        RECT 54.950 80.460 57.095 80.600 ;
        RECT 54.950 80.400 55.270 80.460 ;
        RECT 56.805 80.415 57.095 80.460 ;
        RECT 59.550 80.400 59.870 80.660 ;
        RECT 60.100 80.600 60.240 80.755 ;
        RECT 60.470 80.740 60.790 80.800 ;
        RECT 61.865 80.755 62.155 80.800 ;
        RECT 62.400 80.800 75.035 80.940 ;
        RECT 60.100 80.460 62.080 80.600 ;
        RECT 61.940 80.320 62.080 80.460 ;
        RECT 53.585 80.260 53.875 80.305 ;
        RECT 52.650 80.120 53.875 80.260 ;
        RECT 52.650 80.060 52.970 80.120 ;
        RECT 53.585 80.075 53.875 80.120 ;
        RECT 54.505 80.075 54.795 80.305 ;
        RECT 56.330 80.260 56.650 80.320 ;
        RECT 60.485 80.260 60.775 80.305 ;
        RECT 56.330 80.120 60.775 80.260 ;
        RECT 56.330 80.060 56.650 80.120 ;
        RECT 60.485 80.075 60.775 80.120 ;
        RECT 61.850 80.060 62.170 80.320 ;
        RECT 37.945 79.780 38.710 79.920 ;
        RECT 37.945 79.735 38.235 79.780 ;
        RECT 38.390 79.720 38.710 79.780 ;
        RECT 38.865 79.735 39.155 79.965 ;
        RECT 40.245 79.735 40.535 79.965 ;
        RECT 45.765 79.920 46.055 79.965 ;
        RECT 46.670 79.920 46.990 79.980 ;
        RECT 45.765 79.780 46.990 79.920 ;
        RECT 45.765 79.735 46.055 79.780 ;
        RECT 30.570 79.580 30.890 79.640 ;
        RECT 40.320 79.580 40.460 79.735 ;
        RECT 46.670 79.720 46.990 79.780 ;
        RECT 47.145 79.735 47.435 79.965 ;
        RECT 42.990 79.580 43.310 79.640 ;
        RECT 30.570 79.440 43.310 79.580 ;
        RECT 47.220 79.580 47.360 79.735 ;
        RECT 48.050 79.720 48.370 79.980 ;
        RECT 49.430 79.720 49.750 79.980 ;
        RECT 51.270 79.920 51.590 79.980 ;
        RECT 62.400 79.965 62.540 80.800 ;
        RECT 74.745 80.755 75.035 80.800 ;
        RECT 77.965 80.940 78.255 80.985 ;
        RECT 82.550 80.940 82.870 81.000 ;
        RECT 84.850 80.940 85.170 81.000 ;
        RECT 88.085 80.940 88.375 80.985 ;
        RECT 77.965 80.800 83.700 80.940 ;
        RECT 77.965 80.755 78.255 80.800 ;
        RECT 82.550 80.740 82.870 80.800 ;
        RECT 63.230 80.600 63.550 80.660 ;
        RECT 62.860 80.460 63.550 80.600 ;
        RECT 53.125 79.920 53.415 79.965 ;
        RECT 51.270 79.780 53.415 79.920 ;
        RECT 51.270 79.720 51.590 79.780 ;
        RECT 53.125 79.735 53.415 79.780 ;
        RECT 60.025 79.735 60.315 79.965 ;
        RECT 62.325 79.735 62.615 79.965 ;
        RECT 48.510 79.580 48.830 79.640 ;
        RECT 47.220 79.440 48.830 79.580 ;
        RECT 60.100 79.580 60.240 79.735 ;
        RECT 62.860 79.580 63.000 80.460 ;
        RECT 63.230 80.400 63.550 80.460 ;
        RECT 66.030 80.600 66.320 80.645 ;
        RECT 68.130 80.600 68.420 80.645 ;
        RECT 69.700 80.600 69.990 80.645 ;
        RECT 66.030 80.460 69.990 80.600 ;
        RECT 66.030 80.415 66.320 80.460 ;
        RECT 68.130 80.415 68.420 80.460 ;
        RECT 69.700 80.415 69.990 80.460 ;
        RECT 76.570 80.600 76.890 80.660 ;
        RECT 77.505 80.600 77.795 80.645 ;
        RECT 76.570 80.460 77.795 80.600 ;
        RECT 76.570 80.400 76.890 80.460 ;
        RECT 77.505 80.415 77.795 80.460 ;
        RECT 79.370 80.600 79.660 80.645 ;
        RECT 81.470 80.600 81.760 80.645 ;
        RECT 83.040 80.600 83.330 80.645 ;
        RECT 79.370 80.460 83.330 80.600 ;
        RECT 83.560 80.600 83.700 80.800 ;
        RECT 84.850 80.800 88.375 80.940 ;
        RECT 84.850 80.740 85.170 80.800 ;
        RECT 88.085 80.755 88.375 80.800 ;
        RECT 87.150 80.600 87.470 80.660 ;
        RECT 83.560 80.460 87.470 80.600 ;
        RECT 79.370 80.415 79.660 80.460 ;
        RECT 81.470 80.415 81.760 80.460 ;
        RECT 83.040 80.415 83.330 80.460 ;
        RECT 87.150 80.400 87.470 80.460 ;
        RECT 65.070 80.260 65.390 80.320 ;
        RECT 63.320 80.120 65.390 80.260 ;
        RECT 63.320 79.965 63.460 80.120 ;
        RECT 65.070 80.060 65.390 80.120 ;
        RECT 66.425 80.260 66.715 80.305 ;
        RECT 67.615 80.260 67.905 80.305 ;
        RECT 70.135 80.260 70.425 80.305 ;
        RECT 66.425 80.120 70.425 80.260 ;
        RECT 66.425 80.075 66.715 80.120 ;
        RECT 67.615 80.075 67.905 80.120 ;
        RECT 70.135 80.075 70.425 80.120 ;
        RECT 73.350 80.260 73.670 80.320 ;
        RECT 76.110 80.260 76.430 80.320 ;
        RECT 79.765 80.260 80.055 80.305 ;
        RECT 80.955 80.260 81.245 80.305 ;
        RECT 83.475 80.260 83.765 80.305 ;
        RECT 73.350 80.120 75.880 80.260 ;
        RECT 73.350 80.060 73.670 80.120 ;
        RECT 63.245 79.735 63.535 79.965 ;
        RECT 63.690 79.720 64.010 79.980 ;
        RECT 64.165 79.920 64.455 79.965 ;
        RECT 64.610 79.920 64.930 79.980 ;
        RECT 64.165 79.780 64.930 79.920 ;
        RECT 64.165 79.735 64.455 79.780 ;
        RECT 64.610 79.720 64.930 79.780 ;
        RECT 65.545 79.920 65.835 79.965 ;
        RECT 65.990 79.920 66.310 79.980 ;
        RECT 72.905 79.920 73.195 79.965 ;
        RECT 75.205 79.920 75.495 79.965 ;
        RECT 65.545 79.780 66.310 79.920 ;
        RECT 65.545 79.735 65.835 79.780 ;
        RECT 65.990 79.720 66.310 79.780 ;
        RECT 66.540 79.780 73.195 79.920 ;
        RECT 66.540 79.580 66.680 79.780 ;
        RECT 72.905 79.735 73.195 79.780 ;
        RECT 74.360 79.780 75.495 79.920 ;
        RECT 75.740 79.920 75.880 80.120 ;
        RECT 76.110 80.120 78.640 80.260 ;
        RECT 76.110 80.060 76.430 80.120 ;
        RECT 75.740 79.890 76.800 79.920 ;
        RECT 76.990 79.890 77.280 79.935 ;
        RECT 75.740 79.780 77.280 79.890 ;
        RECT 60.100 79.440 63.000 79.580 ;
        RECT 64.700 79.440 66.680 79.580 ;
        RECT 66.880 79.580 67.170 79.625 ;
        RECT 67.370 79.580 67.690 79.640 ;
        RECT 66.880 79.440 67.690 79.580 ;
        RECT 30.570 79.380 30.890 79.440 ;
        RECT 42.990 79.380 43.310 79.440 ;
        RECT 48.510 79.380 48.830 79.440 ;
        RECT 23.670 79.040 23.990 79.300 ;
        RECT 27.810 79.240 28.130 79.300 ;
        RECT 29.205 79.240 29.495 79.285 ;
        RECT 27.810 79.100 29.495 79.240 ;
        RECT 27.810 79.040 28.130 79.100 ;
        RECT 29.205 79.055 29.495 79.100 ;
        RECT 29.650 79.240 29.970 79.300 ;
        RECT 32.410 79.240 32.730 79.300 ;
        RECT 29.650 79.100 32.730 79.240 ;
        RECT 29.650 79.040 29.970 79.100 ;
        RECT 32.410 79.040 32.730 79.100 ;
        RECT 32.885 79.240 33.175 79.285 ;
        RECT 34.250 79.240 34.570 79.300 ;
        RECT 32.885 79.100 34.570 79.240 ;
        RECT 32.885 79.055 33.175 79.100 ;
        RECT 34.250 79.040 34.570 79.100 ;
        RECT 34.710 79.240 35.030 79.300 ;
        RECT 35.645 79.240 35.935 79.285 ;
        RECT 34.710 79.100 35.935 79.240 ;
        RECT 34.710 79.040 35.030 79.100 ;
        RECT 35.645 79.055 35.935 79.100 ;
        RECT 36.550 79.240 36.870 79.300 ;
        RECT 39.325 79.240 39.615 79.285 ;
        RECT 36.550 79.100 39.615 79.240 ;
        RECT 36.550 79.040 36.870 79.100 ;
        RECT 39.325 79.055 39.615 79.100 ;
        RECT 41.150 79.040 41.470 79.300 ;
        RECT 48.050 79.240 48.370 79.300 ;
        RECT 51.285 79.240 51.575 79.285 ;
        RECT 48.050 79.100 51.575 79.240 ;
        RECT 48.050 79.040 48.370 79.100 ;
        RECT 51.285 79.055 51.575 79.100 ;
        RECT 58.645 79.240 58.935 79.285 ;
        RECT 60.010 79.240 60.330 79.300 ;
        RECT 58.645 79.100 60.330 79.240 ;
        RECT 58.645 79.055 58.935 79.100 ;
        RECT 60.010 79.040 60.330 79.100 ;
        RECT 61.850 79.240 62.170 79.300 ;
        RECT 64.700 79.240 64.840 79.440 ;
        RECT 66.880 79.395 67.170 79.440 ;
        RECT 67.370 79.380 67.690 79.440 ;
        RECT 71.050 79.580 71.370 79.640 ;
        RECT 73.825 79.580 74.115 79.625 ;
        RECT 71.050 79.440 74.115 79.580 ;
        RECT 71.050 79.380 71.370 79.440 ;
        RECT 73.825 79.395 74.115 79.440 ;
        RECT 61.850 79.100 64.840 79.240 ;
        RECT 65.085 79.240 65.375 79.285 ;
        RECT 70.590 79.240 70.910 79.300 ;
        RECT 65.085 79.100 70.910 79.240 ;
        RECT 61.850 79.040 62.170 79.100 ;
        RECT 65.085 79.055 65.375 79.100 ;
        RECT 70.590 79.040 70.910 79.100 ;
        RECT 72.445 79.240 72.735 79.285 ;
        RECT 72.890 79.240 73.210 79.300 ;
        RECT 72.445 79.100 73.210 79.240 ;
        RECT 72.445 79.055 72.735 79.100 ;
        RECT 72.890 79.040 73.210 79.100 ;
        RECT 73.350 79.240 73.670 79.300 ;
        RECT 74.360 79.240 74.500 79.780 ;
        RECT 75.205 79.735 75.495 79.780 ;
        RECT 76.660 79.750 77.280 79.780 ;
        RECT 76.990 79.705 77.280 79.750 ;
        RECT 78.500 79.625 78.640 80.120 ;
        RECT 79.765 80.120 83.765 80.260 ;
        RECT 79.765 80.075 80.055 80.120 ;
        RECT 80.955 80.075 81.245 80.120 ;
        RECT 83.475 80.075 83.765 80.120 ;
        RECT 78.885 79.920 79.175 79.965 ;
        RECT 79.330 79.920 79.650 79.980 ;
        RECT 80.250 79.965 80.570 79.980 ;
        RECT 80.220 79.920 80.570 79.965 ;
        RECT 78.885 79.780 79.650 79.920 ;
        RECT 80.055 79.780 80.570 79.920 ;
        RECT 78.885 79.735 79.175 79.780 ;
        RECT 79.330 79.720 79.650 79.780 ;
        RECT 80.220 79.735 80.570 79.780 ;
        RECT 80.250 79.720 80.570 79.735 ;
        RECT 84.850 79.920 85.170 79.980 ;
        RECT 87.165 79.920 87.455 79.965 ;
        RECT 84.850 79.780 87.455 79.920 ;
        RECT 84.850 79.720 85.170 79.780 ;
        RECT 87.165 79.735 87.455 79.780 ;
        RECT 78.425 79.580 78.715 79.625 ;
        RECT 83.010 79.580 83.330 79.640 ;
        RECT 78.425 79.440 83.330 79.580 ;
        RECT 78.425 79.395 78.715 79.440 ;
        RECT 83.010 79.380 83.330 79.440 ;
        RECT 86.245 79.580 86.535 79.625 ;
        RECT 87.610 79.580 87.930 79.640 ;
        RECT 86.245 79.440 87.930 79.580 ;
        RECT 86.245 79.395 86.535 79.440 ;
        RECT 87.610 79.380 87.930 79.440 ;
        RECT 73.350 79.100 74.500 79.240 ;
        RECT 75.650 79.240 75.970 79.300 ;
        RECT 81.170 79.240 81.490 79.300 ;
        RECT 75.650 79.100 81.490 79.240 ;
        RECT 73.350 79.040 73.670 79.100 ;
        RECT 75.650 79.040 75.970 79.100 ;
        RECT 81.170 79.040 81.490 79.100 ;
        RECT 85.785 79.240 86.075 79.285 ;
        RECT 86.690 79.240 87.010 79.300 ;
        RECT 85.785 79.100 87.010 79.240 ;
        RECT 85.785 79.055 86.075 79.100 ;
        RECT 86.690 79.040 87.010 79.100 ;
        RECT 12.100 78.420 89.840 78.900 ;
        RECT 20.910 78.220 21.230 78.280 ;
        RECT 22.290 78.220 22.610 78.280 ;
        RECT 29.665 78.220 29.955 78.265 ;
        RECT 32.410 78.220 32.730 78.280 ;
        RECT 33.790 78.220 34.110 78.280 ;
        RECT 20.910 78.080 28.500 78.220 ;
        RECT 20.910 78.020 21.230 78.080 ;
        RECT 22.290 78.020 22.610 78.080 ;
        RECT 25.065 77.880 25.355 77.925 ;
        RECT 25.510 77.880 25.830 77.940 ;
        RECT 25.065 77.740 25.830 77.880 ;
        RECT 25.065 77.695 25.355 77.740 ;
        RECT 25.510 77.680 25.830 77.740 ;
        RECT 26.215 77.710 26.505 77.755 ;
        RECT 15.865 77.355 16.155 77.585 ;
        RECT 15.940 77.200 16.080 77.355 ;
        RECT 16.770 77.340 17.090 77.600 ;
        RECT 23.685 77.355 23.975 77.585 ;
        RECT 18.610 77.200 18.930 77.260 ;
        RECT 15.940 77.060 18.930 77.200 ;
        RECT 23.760 77.200 23.900 77.355 ;
        RECT 24.590 77.340 24.910 77.600 ;
        RECT 26.190 77.540 26.505 77.710 ;
        RECT 27.810 77.540 28.130 77.600 ;
        RECT 28.360 77.585 28.500 78.080 ;
        RECT 29.665 78.080 34.110 78.220 ;
        RECT 29.665 78.035 29.955 78.080 ;
        RECT 32.410 78.020 32.730 78.080 ;
        RECT 33.790 78.020 34.110 78.080 ;
        RECT 41.165 78.220 41.455 78.265 ;
        RECT 42.070 78.220 42.390 78.280 ;
        RECT 41.165 78.080 42.390 78.220 ;
        RECT 41.165 78.035 41.455 78.080 ;
        RECT 42.070 78.020 42.390 78.080 ;
        RECT 52.190 78.220 52.510 78.280 ;
        RECT 53.585 78.220 53.875 78.265 ;
        RECT 52.190 78.080 53.875 78.220 ;
        RECT 52.190 78.020 52.510 78.080 ;
        RECT 53.585 78.035 53.875 78.080 ;
        RECT 55.425 78.220 55.715 78.265 ;
        RECT 59.090 78.220 59.410 78.280 ;
        RECT 55.425 78.080 59.410 78.220 ;
        RECT 55.425 78.035 55.715 78.080 ;
        RECT 59.090 78.020 59.410 78.080 ;
        RECT 60.485 78.220 60.775 78.265 ;
        RECT 61.850 78.220 62.170 78.280 ;
        RECT 60.485 78.080 62.170 78.220 ;
        RECT 60.485 78.035 60.775 78.080 ;
        RECT 61.850 78.020 62.170 78.080 ;
        RECT 70.590 78.020 70.910 78.280 ;
        RECT 77.490 78.020 77.810 78.280 ;
        RECT 78.885 78.220 79.175 78.265 ;
        RECT 82.550 78.220 82.870 78.280 ;
        RECT 78.885 78.080 82.870 78.220 ;
        RECT 78.885 78.035 79.175 78.080 ;
        RECT 82.550 78.020 82.870 78.080 ;
        RECT 87.610 78.020 87.930 78.280 ;
        RECT 47.130 77.880 47.450 77.940 ;
        RECT 57.710 77.880 58.030 77.940 ;
        RECT 29.280 77.740 35.860 77.880 ;
        RECT 26.190 77.400 28.130 77.540 ;
        RECT 27.810 77.340 28.130 77.400 ;
        RECT 28.285 77.540 28.575 77.585 ;
        RECT 28.730 77.540 29.050 77.600 ;
        RECT 29.280 77.585 29.420 77.740 ;
        RECT 28.285 77.400 29.050 77.540 ;
        RECT 28.285 77.355 28.575 77.400 ;
        RECT 28.730 77.340 29.050 77.400 ;
        RECT 29.205 77.355 29.495 77.585 ;
        RECT 32.410 77.540 32.730 77.600 ;
        RECT 30.200 77.400 32.730 77.540 ;
        RECT 26.890 77.200 27.210 77.260 ;
        RECT 23.760 77.060 27.210 77.200 ;
        RECT 18.610 77.000 18.930 77.060 ;
        RECT 26.890 77.000 27.210 77.060 ;
        RECT 27.365 77.200 27.655 77.245 ;
        RECT 30.200 77.200 30.340 77.400 ;
        RECT 32.410 77.340 32.730 77.400 ;
        RECT 35.170 77.585 35.490 77.600 ;
        RECT 35.170 77.355 35.520 77.585 ;
        RECT 35.720 77.540 35.860 77.740 ;
        RECT 36.640 77.740 45.980 77.880 ;
        RECT 36.640 77.585 36.780 77.740 ;
        RECT 35.720 77.400 36.320 77.540 ;
        RECT 35.170 77.340 35.490 77.355 ;
        RECT 27.365 77.060 30.340 77.200 ;
        RECT 31.975 77.200 32.265 77.245 ;
        RECT 34.495 77.200 34.785 77.245 ;
        RECT 35.685 77.200 35.975 77.245 ;
        RECT 31.975 77.060 35.975 77.200 ;
        RECT 36.180 77.200 36.320 77.400 ;
        RECT 36.565 77.355 36.855 77.585 ;
        RECT 38.405 77.540 38.695 77.585 ;
        RECT 40.690 77.540 41.010 77.600 ;
        RECT 38.405 77.400 41.010 77.540 ;
        RECT 38.405 77.355 38.695 77.400 ;
        RECT 40.690 77.340 41.010 77.400 ;
        RECT 41.150 77.340 41.470 77.600 ;
        RECT 41.610 77.340 41.930 77.600 ;
        RECT 45.840 77.585 45.980 77.740 ;
        RECT 47.130 77.740 58.030 77.880 ;
        RECT 47.130 77.680 47.450 77.740 ;
        RECT 57.710 77.680 58.030 77.740 ;
        RECT 72.890 77.880 73.210 77.940 ;
        RECT 80.680 77.880 80.970 77.925 ;
        RECT 82.090 77.880 82.410 77.940 ;
        RECT 72.890 77.740 78.180 77.880 ;
        RECT 72.890 77.680 73.210 77.740 ;
        RECT 45.765 77.540 46.055 77.585 ;
        RECT 46.670 77.540 46.990 77.600 ;
        RECT 48.050 77.585 48.370 77.600 ;
        RECT 48.020 77.540 48.370 77.585 ;
        RECT 45.765 77.400 46.990 77.540 ;
        RECT 47.855 77.400 48.370 77.540 ;
        RECT 45.765 77.355 46.055 77.400 ;
        RECT 46.670 77.340 46.990 77.400 ;
        RECT 48.020 77.355 48.370 77.400 ;
        RECT 48.050 77.340 48.370 77.355 ;
        RECT 54.030 77.540 54.350 77.600 ;
        RECT 56.345 77.540 56.635 77.585 ;
        RECT 54.030 77.400 56.635 77.540 ;
        RECT 54.030 77.340 54.350 77.400 ;
        RECT 56.345 77.355 56.635 77.400 ;
        RECT 47.565 77.200 47.855 77.245 ;
        RECT 48.755 77.200 49.045 77.245 ;
        RECT 51.275 77.200 51.565 77.245 ;
        RECT 36.180 77.060 40.460 77.200 ;
        RECT 27.365 77.015 27.655 77.060 ;
        RECT 31.975 77.015 32.265 77.060 ;
        RECT 34.495 77.015 34.785 77.060 ;
        RECT 35.685 77.015 35.975 77.060 ;
        RECT 24.590 76.860 24.910 76.920 ;
        RECT 28.270 76.860 28.590 76.920 ;
        RECT 31.030 76.860 31.350 76.920 ;
        RECT 24.590 76.720 31.350 76.860 ;
        RECT 24.590 76.660 24.910 76.720 ;
        RECT 28.270 76.660 28.590 76.720 ;
        RECT 31.030 76.660 31.350 76.720 ;
        RECT 32.410 76.860 32.700 76.905 ;
        RECT 33.980 76.860 34.270 76.905 ;
        RECT 36.080 76.860 36.370 76.905 ;
        RECT 32.410 76.720 36.370 76.860 ;
        RECT 32.410 76.675 32.700 76.720 ;
        RECT 33.980 76.675 34.270 76.720 ;
        RECT 36.080 76.675 36.370 76.720 ;
        RECT 39.770 76.660 40.090 76.920 ;
        RECT 40.320 76.905 40.460 77.060 ;
        RECT 47.565 77.060 51.565 77.200 ;
        RECT 56.420 77.200 56.560 77.355 ;
        RECT 57.250 77.340 57.570 77.600 ;
        RECT 59.550 77.340 59.870 77.600 ;
        RECT 61.405 77.540 61.695 77.585 ;
        RECT 62.770 77.540 63.090 77.600 ;
        RECT 60.100 77.400 63.090 77.540 ;
        RECT 58.645 77.200 58.935 77.245 ;
        RECT 56.420 77.060 58.935 77.200 ;
        RECT 47.565 77.015 47.855 77.060 ;
        RECT 48.755 77.015 49.045 77.060 ;
        RECT 51.275 77.015 51.565 77.060 ;
        RECT 58.645 77.015 58.935 77.060 ;
        RECT 59.090 77.200 59.410 77.260 ;
        RECT 60.100 77.200 60.240 77.400 ;
        RECT 61.405 77.355 61.695 77.400 ;
        RECT 62.770 77.340 63.090 77.400 ;
        RECT 63.245 77.540 63.535 77.585 ;
        RECT 66.910 77.540 67.230 77.600 ;
        RECT 63.245 77.400 67.230 77.540 ;
        RECT 63.245 77.355 63.535 77.400 ;
        RECT 66.910 77.340 67.230 77.400 ;
        RECT 70.145 77.540 70.435 77.585 ;
        RECT 72.445 77.540 72.735 77.585 ;
        RECT 70.145 77.400 72.735 77.540 ;
        RECT 70.145 77.355 70.435 77.400 ;
        RECT 72.445 77.355 72.735 77.400 ;
        RECT 76.110 77.340 76.430 77.600 ;
        RECT 78.040 77.585 78.180 77.740 ;
        RECT 80.680 77.740 82.410 77.880 ;
        RECT 80.680 77.695 80.970 77.740 ;
        RECT 82.090 77.680 82.410 77.740 ;
        RECT 99.980 77.735 100.370 81.555 ;
        RECT 101.460 81.315 102.460 83.715 ;
        RECT 102.950 81.585 103.950 83.735 ;
        RECT 101.210 81.085 102.460 81.315 ;
        RECT 100.650 80.925 102.460 81.085 ;
        RECT 102.720 80.945 103.950 81.585 ;
        RECT 104.430 81.575 105.430 83.725 ;
        RECT 105.890 81.575 106.890 83.715 ;
        RECT 100.650 80.625 101.930 80.925 ;
        RECT 100.650 78.745 101.650 80.625 ;
        RECT 102.720 80.475 103.400 80.945 ;
        RECT 104.210 80.935 105.430 81.575 ;
        RECT 104.210 80.475 104.890 80.935 ;
        RECT 105.700 80.925 106.890 81.575 ;
        RECT 107.390 81.545 108.390 83.735 ;
        RECT 110.330 83.715 112.640 83.725 ;
        RECT 107.150 80.945 108.390 81.545 ;
        RECT 108.900 81.535 109.900 83.715 ;
        RECT 110.330 81.545 112.810 83.715 ;
        RECT 105.700 80.475 106.380 80.925 ;
        RECT 107.150 80.475 107.830 80.945 ;
        RECT 102.100 80.005 103.400 80.475 ;
        RECT 102.100 78.835 103.140 80.005 ;
        RECT 103.610 79.995 104.890 80.475 ;
        RECT 105.080 79.995 106.380 80.475 ;
        RECT 103.610 78.835 104.650 79.995 ;
        RECT 105.080 78.835 106.120 79.995 ;
        RECT 106.570 79.965 107.830 80.475 ;
        RECT 108.650 80.925 109.900 81.535 ;
        RECT 110.160 80.935 112.810 81.545 ;
        RECT 108.650 80.465 109.330 80.925 ;
        RECT 110.160 80.475 110.840 80.935 ;
        RECT 111.810 80.925 112.810 80.935 ;
        RECT 100.650 78.295 101.880 78.745 ;
        RECT 102.100 78.295 103.430 78.835 ;
        RECT 103.610 78.295 104.920 78.835 ;
        RECT 105.080 78.295 106.410 78.835 ;
        RECT 106.570 78.825 107.610 79.965 ;
        RECT 108.050 79.955 109.330 80.465 ;
        RECT 109.530 79.965 110.840 80.475 ;
        RECT 108.050 78.825 109.090 79.955 ;
        RECT 106.570 78.295 107.840 78.825 ;
        RECT 101.200 77.735 101.880 78.295 ;
        RECT 102.750 77.745 103.430 78.295 ;
        RECT 104.240 77.755 104.920 78.295 ;
        RECT 105.730 77.755 106.410 78.295 ;
        RECT 107.160 77.755 107.840 78.295 ;
        RECT 108.050 78.285 109.350 78.825 ;
        RECT 109.530 78.295 110.570 79.965 ;
        RECT 108.670 77.755 109.350 78.285 ;
        RECT 77.505 77.355 77.795 77.585 ;
        RECT 77.965 77.355 78.255 77.585 ;
        RECT 59.090 77.060 60.240 77.200 ;
        RECT 60.470 77.200 60.790 77.260 ;
        RECT 64.165 77.200 64.455 77.245 ;
        RECT 60.470 77.060 64.455 77.200 ;
        RECT 59.090 77.000 59.410 77.060 ;
        RECT 60.470 77.000 60.790 77.060 ;
        RECT 64.165 77.015 64.455 77.060 ;
        RECT 68.750 77.200 69.070 77.260 ;
        RECT 71.065 77.200 71.355 77.245 ;
        RECT 68.750 77.060 71.355 77.200 ;
        RECT 68.750 77.000 69.070 77.060 ;
        RECT 71.065 77.015 71.355 77.060 ;
        RECT 75.650 77.000 75.970 77.260 ;
        RECT 77.580 77.200 77.720 77.355 ;
        RECT 86.690 77.340 87.010 77.600 ;
        RECT 78.410 77.200 78.730 77.260 ;
        RECT 77.580 77.060 78.730 77.200 ;
        RECT 78.410 77.000 78.730 77.060 ;
        RECT 79.330 77.000 79.650 77.260 ;
        RECT 80.225 77.200 80.515 77.245 ;
        RECT 81.415 77.200 81.705 77.245 ;
        RECT 83.935 77.200 84.225 77.245 ;
        RECT 80.225 77.060 84.225 77.200 ;
        RECT 80.225 77.015 80.515 77.060 ;
        RECT 81.415 77.015 81.705 77.060 ;
        RECT 83.935 77.015 84.225 77.060 ;
        RECT 40.245 76.675 40.535 76.905 ;
        RECT 47.170 76.860 47.460 76.905 ;
        RECT 49.270 76.860 49.560 76.905 ;
        RECT 50.840 76.860 51.130 76.905 ;
        RECT 47.170 76.720 51.130 76.860 ;
        RECT 47.170 76.675 47.460 76.720 ;
        RECT 49.270 76.675 49.560 76.720 ;
        RECT 50.840 76.675 51.130 76.720 ;
        RECT 76.570 76.860 76.890 76.920 ;
        RECT 77.045 76.860 77.335 76.905 ;
        RECT 76.570 76.720 77.335 76.860 ;
        RECT 76.570 76.660 76.890 76.720 ;
        RECT 77.045 76.675 77.335 76.720 ;
        RECT 79.830 76.860 80.120 76.905 ;
        RECT 81.930 76.860 82.220 76.905 ;
        RECT 83.500 76.860 83.790 76.905 ;
        RECT 79.830 76.720 83.790 76.860 ;
        RECT 79.830 76.675 80.120 76.720 ;
        RECT 81.930 76.675 82.220 76.720 ;
        RECT 83.500 76.675 83.790 76.720 ;
        RECT 16.310 76.320 16.630 76.580 ;
        RECT 24.145 76.520 24.435 76.565 ;
        RECT 25.050 76.520 25.370 76.580 ;
        RECT 24.145 76.380 25.370 76.520 ;
        RECT 24.145 76.335 24.435 76.380 ;
        RECT 25.050 76.320 25.370 76.380 ;
        RECT 25.985 76.520 26.275 76.565 ;
        RECT 26.430 76.520 26.750 76.580 ;
        RECT 25.985 76.380 26.750 76.520 ;
        RECT 25.985 76.335 26.275 76.380 ;
        RECT 26.430 76.320 26.750 76.380 ;
        RECT 26.890 76.320 27.210 76.580 ;
        RECT 28.730 76.520 29.050 76.580 ;
        RECT 33.330 76.520 33.650 76.580 ;
        RECT 28.730 76.380 33.650 76.520 ;
        RECT 28.730 76.320 29.050 76.380 ;
        RECT 33.330 76.320 33.650 76.380 ;
        RECT 35.630 76.520 35.950 76.580 ;
        RECT 39.095 76.520 39.385 76.565 ;
        RECT 35.630 76.380 39.385 76.520 ;
        RECT 35.630 76.320 35.950 76.380 ;
        RECT 39.095 76.335 39.385 76.380 ;
        RECT 67.370 76.320 67.690 76.580 ;
        RECT 67.830 76.520 68.150 76.580 ;
        RECT 68.305 76.520 68.595 76.565 ;
        RECT 67.830 76.380 68.595 76.520 ;
        RECT 67.830 76.320 68.150 76.380 ;
        RECT 68.305 76.335 68.595 76.380 ;
        RECT 84.850 76.520 85.170 76.580 ;
        RECT 86.245 76.520 86.535 76.565 ;
        RECT 84.850 76.380 86.535 76.520 ;
        RECT 84.850 76.320 85.170 76.380 ;
        RECT 86.245 76.335 86.535 76.380 ;
        RECT 12.100 75.700 89.840 76.180 ;
        RECT 99.980 75.585 101.000 77.735 ;
        RECT 101.200 77.165 102.510 77.735 ;
        RECT 102.750 77.255 103.960 77.745 ;
        RECT 104.240 77.255 105.470 77.755 ;
        RECT 105.730 77.255 106.940 77.755 ;
        RECT 101.470 75.575 102.510 77.165 ;
        RECT 102.920 75.565 103.960 77.255 ;
        RECT 104.430 75.575 105.470 77.255 ;
        RECT 105.900 75.575 106.940 77.255 ;
        RECT 107.160 77.245 108.430 77.755 ;
        RECT 108.670 77.245 109.900 77.755 ;
        RECT 107.390 75.575 108.430 77.245 ;
        RECT 108.860 75.575 109.900 77.245 ;
        RECT 30.570 75.500 30.890 75.560 ;
        RECT 32.870 75.500 33.190 75.560 ;
        RECT 13.640 75.360 33.190 75.500 ;
        RECT 13.640 74.865 13.780 75.360 ;
        RECT 30.570 75.300 30.890 75.360 ;
        RECT 32.870 75.300 33.190 75.360 ;
        RECT 42.530 75.300 42.850 75.560 ;
        RECT 71.510 75.500 71.830 75.560 ;
        RECT 76.110 75.500 76.430 75.560 ;
        RECT 82.090 75.500 82.410 75.560 ;
        RECT 71.510 75.360 83.240 75.500 ;
        RECT 71.510 75.300 71.830 75.360 ;
        RECT 76.110 75.300 76.430 75.360 ;
        RECT 82.090 75.300 82.410 75.360 ;
        RECT 14.050 75.160 14.340 75.205 ;
        RECT 16.150 75.160 16.440 75.205 ;
        RECT 17.720 75.160 18.010 75.205 ;
        RECT 14.050 75.020 18.010 75.160 ;
        RECT 14.050 74.975 14.340 75.020 ;
        RECT 16.150 74.975 16.440 75.020 ;
        RECT 17.720 74.975 18.010 75.020 ;
        RECT 18.610 75.160 18.930 75.220 ;
        RECT 20.465 75.160 20.755 75.205 ;
        RECT 18.610 75.020 20.755 75.160 ;
        RECT 18.610 74.960 18.930 75.020 ;
        RECT 20.465 74.975 20.755 75.020 ;
        RECT 22.290 75.160 22.610 75.220 ;
        RECT 22.765 75.160 23.055 75.205 ;
        RECT 27.365 75.160 27.655 75.205 ;
        RECT 27.810 75.160 28.130 75.220 ;
        RECT 42.990 75.160 43.310 75.220 ;
        RECT 64.150 75.160 64.470 75.220 ;
        RECT 66.950 75.160 67.240 75.205 ;
        RECT 69.050 75.160 69.340 75.205 ;
        RECT 70.620 75.160 70.910 75.205 ;
        RECT 22.290 75.020 26.660 75.160 ;
        RECT 13.565 74.635 13.855 74.865 ;
        RECT 14.445 74.820 14.735 74.865 ;
        RECT 15.635 74.820 15.925 74.865 ;
        RECT 18.155 74.820 18.445 74.865 ;
        RECT 14.445 74.680 18.445 74.820 ;
        RECT 20.540 74.820 20.680 74.975 ;
        RECT 22.290 74.960 22.610 75.020 ;
        RECT 22.765 74.975 23.055 75.020 ;
        RECT 23.225 74.820 23.515 74.865 ;
        RECT 20.540 74.680 23.515 74.820 ;
        RECT 14.445 74.635 14.735 74.680 ;
        RECT 15.635 74.635 15.925 74.680 ;
        RECT 18.155 74.635 18.445 74.680 ;
        RECT 23.225 74.635 23.515 74.680 ;
        RECT 20.910 74.480 21.230 74.540 ;
        RECT 21.385 74.480 21.675 74.525 ;
        RECT 20.910 74.340 21.675 74.480 ;
        RECT 20.910 74.280 21.230 74.340 ;
        RECT 21.385 74.295 21.675 74.340 ;
        RECT 21.830 74.480 22.150 74.540 ;
        RECT 24.145 74.480 24.435 74.525 ;
        RECT 21.830 74.340 24.435 74.480 ;
        RECT 21.830 74.280 22.150 74.340 ;
        RECT 24.145 74.295 24.435 74.340 ;
        RECT 24.590 74.280 24.910 74.540 ;
        RECT 26.520 74.525 26.660 75.020 ;
        RECT 27.365 75.020 28.130 75.160 ;
        RECT 27.365 74.975 27.655 75.020 ;
        RECT 27.810 74.960 28.130 75.020 ;
        RECT 42.620 75.020 43.310 75.160 ;
        RECT 26.905 74.820 27.195 74.865 ;
        RECT 31.030 74.820 31.350 74.880 ;
        RECT 26.905 74.680 31.350 74.820 ;
        RECT 26.905 74.635 27.195 74.680 ;
        RECT 31.030 74.620 31.350 74.680 ;
        RECT 32.870 74.820 33.190 74.880 ;
        RECT 33.345 74.820 33.635 74.865 ;
        RECT 32.870 74.680 33.635 74.820 ;
        RECT 32.870 74.620 33.190 74.680 ;
        RECT 33.345 74.635 33.635 74.680 ;
        RECT 36.550 74.820 36.870 74.880 ;
        RECT 42.620 74.865 42.760 75.020 ;
        RECT 42.990 74.960 43.310 75.020 ;
        RECT 61.480 75.020 65.300 75.160 ;
        RECT 37.025 74.820 37.315 74.865 ;
        RECT 36.550 74.680 37.315 74.820 ;
        RECT 36.550 74.620 36.870 74.680 ;
        RECT 37.025 74.635 37.315 74.680 ;
        RECT 42.545 74.635 42.835 74.865 ;
        RECT 25.525 74.480 25.815 74.525 ;
        RECT 25.095 74.340 25.815 74.480 ;
        RECT 14.930 74.185 15.250 74.200 ;
        RECT 14.900 73.955 15.250 74.185 ;
        RECT 14.930 73.940 15.250 73.955 ;
        RECT 22.750 73.940 23.070 74.200 ;
        RECT 23.225 74.140 23.515 74.185 ;
        RECT 23.670 74.140 23.990 74.200 ;
        RECT 23.225 74.000 23.990 74.140 ;
        RECT 23.225 73.955 23.515 74.000 ;
        RECT 23.670 73.940 23.990 74.000 ;
        RECT 20.910 73.800 21.230 73.860 ;
        RECT 21.845 73.800 22.135 73.845 ;
        RECT 20.910 73.660 22.135 73.800 ;
        RECT 20.910 73.600 21.230 73.660 ;
        RECT 21.845 73.615 22.135 73.660 ;
        RECT 24.130 73.800 24.450 73.860 ;
        RECT 25.095 73.800 25.235 74.340 ;
        RECT 25.525 74.295 25.815 74.340 ;
        RECT 26.445 74.295 26.735 74.525 ;
        RECT 27.810 74.280 28.130 74.540 ;
        RECT 29.665 74.480 29.955 74.525 ;
        RECT 41.610 74.480 41.930 74.540 ;
        RECT 29.665 74.340 41.930 74.480 ;
        RECT 29.665 74.295 29.955 74.340 ;
        RECT 41.610 74.280 41.930 74.340 ;
        RECT 42.990 74.280 43.310 74.540 ;
        RECT 43.910 74.480 44.230 74.540 ;
        RECT 47.590 74.480 47.910 74.540 ;
        RECT 43.910 74.340 47.910 74.480 ;
        RECT 43.910 74.280 44.230 74.340 ;
        RECT 47.590 74.280 47.910 74.340 ;
        RECT 48.050 74.480 48.370 74.540 ;
        RECT 48.525 74.480 48.815 74.525 ;
        RECT 48.050 74.340 48.815 74.480 ;
        RECT 48.050 74.280 48.370 74.340 ;
        RECT 48.525 74.295 48.815 74.340 ;
        RECT 54.950 74.480 55.270 74.540 ;
        RECT 55.870 74.480 56.190 74.540 ;
        RECT 54.950 74.340 56.190 74.480 ;
        RECT 54.950 74.280 55.270 74.340 ;
        RECT 55.870 74.280 56.190 74.340 ;
        RECT 56.330 74.480 56.650 74.540 ;
        RECT 57.725 74.480 58.015 74.525 ;
        RECT 56.330 74.340 58.015 74.480 ;
        RECT 56.330 74.280 56.650 74.340 ;
        RECT 57.725 74.295 58.015 74.340 ;
        RECT 58.185 74.480 58.475 74.525 ;
        RECT 59.550 74.480 59.870 74.540 ;
        RECT 58.185 74.340 59.870 74.480 ;
        RECT 58.185 74.295 58.475 74.340 ;
        RECT 59.550 74.280 59.870 74.340 ;
        RECT 60.010 74.280 60.330 74.540 ;
        RECT 40.690 73.940 41.010 74.200 ;
        RECT 59.105 74.140 59.395 74.185 ;
        RECT 61.480 74.140 61.620 75.020 ;
        RECT 64.150 74.960 64.470 75.020 ;
        RECT 61.850 74.820 62.170 74.880 ;
        RECT 61.850 74.680 64.840 74.820 ;
        RECT 61.850 74.620 62.170 74.680 ;
        RECT 64.700 74.525 64.840 74.680 ;
        RECT 65.160 74.525 65.300 75.020 ;
        RECT 66.950 75.020 70.910 75.160 ;
        RECT 66.950 74.975 67.240 75.020 ;
        RECT 69.050 74.975 69.340 75.020 ;
        RECT 70.620 74.975 70.910 75.020 ;
        RECT 73.365 75.160 73.655 75.205 ;
        RECT 75.650 75.160 75.970 75.220 ;
        RECT 77.490 75.160 77.810 75.220 ;
        RECT 73.365 75.020 77.810 75.160 ;
        RECT 83.100 75.160 83.240 75.360 ;
        RECT 83.470 75.300 83.790 75.560 ;
        RECT 84.390 75.300 84.710 75.560 ;
        RECT 83.100 75.020 83.700 75.160 ;
        RECT 73.365 74.975 73.655 75.020 ;
        RECT 75.650 74.960 75.970 75.020 ;
        RECT 77.490 74.960 77.810 75.020 ;
        RECT 67.345 74.820 67.635 74.865 ;
        RECT 68.535 74.820 68.825 74.865 ;
        RECT 71.055 74.820 71.345 74.865 ;
        RECT 67.345 74.680 71.345 74.820 ;
        RECT 67.345 74.635 67.635 74.680 ;
        RECT 68.535 74.635 68.825 74.680 ;
        RECT 71.055 74.635 71.345 74.680 ;
        RECT 78.410 74.820 78.730 74.880 ;
        RECT 79.805 74.820 80.095 74.865 ;
        RECT 83.010 74.820 83.330 74.880 ;
        RECT 78.410 74.680 80.095 74.820 ;
        RECT 78.410 74.620 78.730 74.680 ;
        RECT 79.805 74.635 80.095 74.680 ;
        RECT 81.720 74.680 83.330 74.820 ;
        RECT 62.785 74.480 63.075 74.525 ;
        RECT 63.245 74.480 63.535 74.525 ;
        RECT 62.785 74.340 63.535 74.480 ;
        RECT 62.785 74.295 63.075 74.340 ;
        RECT 63.245 74.295 63.535 74.340 ;
        RECT 64.625 74.295 64.915 74.525 ;
        RECT 65.085 74.295 65.375 74.525 ;
        RECT 66.450 74.280 66.770 74.540 ;
        RECT 67.830 74.525 68.150 74.540 ;
        RECT 67.800 74.480 68.150 74.525 ;
        RECT 67.635 74.340 68.150 74.480 ;
        RECT 67.800 74.295 68.150 74.340 ;
        RECT 76.125 74.480 76.415 74.525 ;
        RECT 77.030 74.480 77.350 74.540 ;
        RECT 81.720 74.525 81.860 74.680 ;
        RECT 83.010 74.620 83.330 74.680 ;
        RECT 76.125 74.340 77.350 74.480 ;
        RECT 76.125 74.295 76.415 74.340 ;
        RECT 67.830 74.280 68.150 74.295 ;
        RECT 77.030 74.280 77.350 74.340 ;
        RECT 81.645 74.295 81.935 74.525 ;
        RECT 82.550 74.280 82.870 74.540 ;
        RECT 83.560 74.480 83.700 75.020 ;
        RECT 85.325 74.480 85.615 74.525 ;
        RECT 83.560 74.340 85.615 74.480 ;
        RECT 85.325 74.295 85.615 74.340 ;
        RECT 87.150 74.280 87.470 74.540 ;
        RECT 59.105 74.000 61.620 74.140 ;
        RECT 59.105 73.955 59.395 74.000 ;
        RECT 64.165 73.955 64.455 74.185 ;
        RECT 80.250 74.140 80.570 74.200 ;
        RECT 80.725 74.140 81.015 74.185 ;
        RECT 75.280 74.000 80.020 74.140 ;
        RECT 24.130 73.660 25.235 73.800 ;
        RECT 27.350 73.800 27.670 73.860 ;
        RECT 28.745 73.800 29.035 73.845 ;
        RECT 27.350 73.660 29.035 73.800 ;
        RECT 24.130 73.600 24.450 73.660 ;
        RECT 27.350 73.600 27.670 73.660 ;
        RECT 28.745 73.615 29.035 73.660 ;
        RECT 39.310 73.800 39.630 73.860 ;
        RECT 40.245 73.800 40.535 73.845 ;
        RECT 39.310 73.660 40.535 73.800 ;
        RECT 39.310 73.600 39.630 73.660 ;
        RECT 40.245 73.615 40.535 73.660 ;
        RECT 43.450 73.800 43.770 73.860 ;
        RECT 43.925 73.800 44.215 73.845 ;
        RECT 43.450 73.660 44.215 73.800 ;
        RECT 43.450 73.600 43.770 73.660 ;
        RECT 43.925 73.615 44.215 73.660 ;
        RECT 45.290 73.800 45.610 73.860 ;
        RECT 45.765 73.800 46.055 73.845 ;
        RECT 45.290 73.660 46.055 73.800 ;
        RECT 45.290 73.600 45.610 73.660 ;
        RECT 45.765 73.615 46.055 73.660 ;
        RECT 55.410 73.800 55.730 73.860 ;
        RECT 56.805 73.800 57.095 73.845 ;
        RECT 55.410 73.660 57.095 73.800 ;
        RECT 55.410 73.600 55.730 73.660 ;
        RECT 56.805 73.615 57.095 73.660 ;
        RECT 58.645 73.800 58.935 73.845 ;
        RECT 64.240 73.800 64.380 73.955 ;
        RECT 58.645 73.660 64.380 73.800 ;
        RECT 65.530 73.800 65.850 73.860 ;
        RECT 75.280 73.845 75.420 74.000 ;
        RECT 79.880 73.860 80.020 74.000 ;
        RECT 80.250 74.000 81.015 74.140 ;
        RECT 80.250 73.940 80.570 74.000 ;
        RECT 80.725 73.955 81.015 74.000 ;
        RECT 83.010 74.140 83.330 74.200 ;
        RECT 85.785 74.140 86.075 74.185 ;
        RECT 83.010 74.000 86.075 74.140 ;
        RECT 83.010 73.940 83.330 74.000 ;
        RECT 85.785 73.955 86.075 74.000 ;
        RECT 86.245 73.955 86.535 74.185 ;
        RECT 66.005 73.800 66.295 73.845 ;
        RECT 65.530 73.660 66.295 73.800 ;
        RECT 58.645 73.615 58.935 73.660 ;
        RECT 65.530 73.600 65.850 73.660 ;
        RECT 66.005 73.615 66.295 73.660 ;
        RECT 75.205 73.615 75.495 73.845 ;
        RECT 77.030 73.600 77.350 73.860 ;
        RECT 79.790 73.800 80.110 73.860 ;
        RECT 85.310 73.800 85.630 73.860 ;
        RECT 86.320 73.800 86.460 73.955 ;
        RECT 79.790 73.660 86.460 73.800 ;
        RECT 79.790 73.600 80.110 73.660 ;
        RECT 85.310 73.600 85.630 73.660 ;
        RECT 12.100 72.980 89.840 73.460 ;
        RECT 14.485 72.780 14.775 72.825 ;
        RECT 14.930 72.780 15.250 72.840 ;
        RECT 14.485 72.640 15.250 72.780 ;
        RECT 14.485 72.595 14.775 72.640 ;
        RECT 14.930 72.580 15.250 72.640 ;
        RECT 15.865 72.780 16.155 72.825 ;
        RECT 16.310 72.780 16.630 72.840 ;
        RECT 15.865 72.640 16.630 72.780 ;
        RECT 15.865 72.595 16.155 72.640 ;
        RECT 16.310 72.580 16.630 72.640 ;
        RECT 23.685 72.780 23.975 72.825 ;
        RECT 25.510 72.780 25.830 72.840 ;
        RECT 31.505 72.780 31.795 72.825 ;
        RECT 35.170 72.780 35.490 72.840 ;
        RECT 23.685 72.640 26.200 72.780 ;
        RECT 23.685 72.595 23.975 72.640 ;
        RECT 25.510 72.580 25.830 72.640 ;
        RECT 15.405 72.440 15.695 72.485 ;
        RECT 17.705 72.440 17.995 72.485 ;
        RECT 15.405 72.300 17.995 72.440 ;
        RECT 15.405 72.255 15.695 72.300 ;
        RECT 17.705 72.255 17.995 72.300 ;
        RECT 18.610 72.240 18.930 72.500 ;
        RECT 20.465 72.440 20.755 72.485 ;
        RECT 20.910 72.440 21.230 72.500 ;
        RECT 26.060 72.485 26.200 72.640 ;
        RECT 31.505 72.640 35.490 72.780 ;
        RECT 31.505 72.595 31.795 72.640 ;
        RECT 35.170 72.580 35.490 72.640 ;
        RECT 35.630 72.580 35.950 72.840 ;
        RECT 38.865 72.780 39.155 72.825 ;
        RECT 42.990 72.780 43.310 72.840 ;
        RECT 47.605 72.780 47.895 72.825 ;
        RECT 38.865 72.640 47.895 72.780 ;
        RECT 38.865 72.595 39.155 72.640 ;
        RECT 42.990 72.580 43.310 72.640 ;
        RECT 47.605 72.595 47.895 72.640 ;
        RECT 48.050 72.580 48.370 72.840 ;
        RECT 58.645 72.595 58.935 72.825 ;
        RECT 60.010 72.780 60.330 72.840 ;
        RECT 60.945 72.780 61.235 72.825 ;
        RECT 60.010 72.640 61.235 72.780 ;
        RECT 20.465 72.300 23.440 72.440 ;
        RECT 20.465 72.255 20.755 72.300 ;
        RECT 20.910 72.240 21.230 72.300 ;
        RECT 15.850 72.100 16.170 72.160 ;
        RECT 16.325 72.100 16.615 72.145 ;
        RECT 15.850 71.960 16.615 72.100 ;
        RECT 15.850 71.900 16.170 71.960 ;
        RECT 16.325 71.915 16.615 71.960 ;
        RECT 16.770 72.100 17.090 72.160 ;
        RECT 19.545 72.100 19.835 72.145 ;
        RECT 16.770 71.960 19.835 72.100 ;
        RECT 16.770 71.900 17.090 71.960 ;
        RECT 19.160 71.820 19.300 71.960 ;
        RECT 19.545 71.915 19.835 71.960 ;
        RECT 20.005 72.100 20.295 72.145 ;
        RECT 21.385 72.100 21.675 72.145 ;
        RECT 22.290 72.100 22.610 72.160 ;
        RECT 22.765 72.100 23.055 72.145 ;
        RECT 20.005 71.960 20.680 72.100 ;
        RECT 20.005 71.915 20.295 71.960 ;
        RECT 20.540 71.820 20.680 71.960 ;
        RECT 21.385 71.960 21.785 72.100 ;
        RECT 22.290 71.960 23.055 72.100 ;
        RECT 21.385 71.915 21.675 71.960 ;
        RECT 17.245 71.760 17.535 71.805 ;
        RECT 18.150 71.760 18.470 71.820 ;
        RECT 17.245 71.620 18.470 71.760 ;
        RECT 17.245 71.575 17.535 71.620 ;
        RECT 18.150 71.560 18.470 71.620 ;
        RECT 19.070 71.560 19.390 71.820 ;
        RECT 20.450 71.560 20.770 71.820 ;
        RECT 21.460 71.760 21.600 71.915 ;
        RECT 22.290 71.900 22.610 71.960 ;
        RECT 22.765 71.915 23.055 71.960 ;
        RECT 21.845 71.760 22.135 71.805 ;
        RECT 21.000 71.620 22.135 71.760 ;
        RECT 23.300 71.760 23.440 72.300 ;
        RECT 25.985 72.255 26.275 72.485 ;
        RECT 30.585 72.440 30.875 72.485 ;
        RECT 40.690 72.440 41.010 72.500 ;
        RECT 58.720 72.440 58.860 72.595 ;
        RECT 60.010 72.580 60.330 72.640 ;
        RECT 60.945 72.595 61.235 72.640 ;
        RECT 66.005 72.780 66.295 72.825 ;
        RECT 67.370 72.780 67.690 72.840 ;
        RECT 66.005 72.640 67.690 72.780 ;
        RECT 66.005 72.595 66.295 72.640 ;
        RECT 67.370 72.580 67.690 72.640 ;
        RECT 70.605 72.780 70.895 72.825 ;
        RECT 74.745 72.780 75.035 72.825 ;
        RECT 77.030 72.780 77.350 72.840 ;
        RECT 70.605 72.640 74.040 72.780 ;
        RECT 70.605 72.595 70.895 72.640 ;
        RECT 30.585 72.300 31.720 72.440 ;
        RECT 30.585 72.255 30.875 72.300 ;
        RECT 31.580 72.160 31.720 72.300 ;
        RECT 32.040 72.300 35.400 72.440 ;
        RECT 25.050 71.900 25.370 72.160 ;
        RECT 25.525 72.100 25.815 72.145 ;
        RECT 26.430 72.100 26.750 72.160 ;
        RECT 25.525 71.960 26.750 72.100 ;
        RECT 25.525 71.915 25.815 71.960 ;
        RECT 26.430 71.900 26.750 71.960 ;
        RECT 26.905 71.915 27.195 72.145 ;
        RECT 25.970 71.760 26.290 71.820 ;
        RECT 23.300 71.620 26.290 71.760 ;
        RECT 18.240 71.420 18.380 71.560 ;
        RECT 19.530 71.420 19.850 71.480 ;
        RECT 18.240 71.280 19.850 71.420 ;
        RECT 19.530 71.220 19.850 71.280 ;
        RECT 21.000 71.080 21.140 71.620 ;
        RECT 21.845 71.575 22.135 71.620 ;
        RECT 25.970 71.560 26.290 71.620 ;
        RECT 21.385 71.420 21.675 71.465 ;
        RECT 26.980 71.420 27.120 71.915 ;
        RECT 27.350 71.900 27.670 72.160 ;
        RECT 31.490 71.900 31.810 72.160 ;
        RECT 32.040 72.145 32.180 72.300 ;
        RECT 35.260 72.160 35.400 72.300 ;
        RECT 37.560 72.300 41.010 72.440 ;
        RECT 31.965 71.915 32.255 72.145 ;
        RECT 32.885 72.100 33.175 72.145 ;
        RECT 34.250 72.100 34.570 72.160 ;
        RECT 32.885 71.960 34.570 72.100 ;
        RECT 32.885 71.915 33.175 71.960 ;
        RECT 34.250 71.900 34.570 71.960 ;
        RECT 34.710 71.900 35.030 72.160 ;
        RECT 35.170 71.900 35.490 72.160 ;
        RECT 36.090 72.100 36.410 72.160 ;
        RECT 37.560 72.145 37.700 72.300 ;
        RECT 40.690 72.240 41.010 72.300 ;
        RECT 41.700 72.300 47.360 72.440 ;
        RECT 36.565 72.100 36.855 72.145 ;
        RECT 36.090 71.960 36.855 72.100 ;
        RECT 36.090 71.900 36.410 71.960 ;
        RECT 36.565 71.915 36.855 71.960 ;
        RECT 37.485 71.915 37.775 72.145 ;
        RECT 39.310 71.900 39.630 72.160 ;
        RECT 33.330 71.560 33.650 71.820 ;
        RECT 33.805 71.575 34.095 71.805 ;
        RECT 37.025 71.760 37.315 71.805 ;
        RECT 41.150 71.760 41.470 71.820 ;
        RECT 41.700 71.760 41.840 72.300 ;
        RECT 45.290 72.145 45.610 72.160 ;
        RECT 45.290 72.100 45.640 72.145 ;
        RECT 45.290 71.960 45.805 72.100 ;
        RECT 45.290 71.915 45.640 71.960 ;
        RECT 45.290 71.900 45.610 71.915 ;
        RECT 46.670 71.900 46.990 72.160 ;
        RECT 47.220 72.145 47.360 72.300 ;
        RECT 47.680 72.300 58.860 72.440 ;
        RECT 47.680 72.160 47.820 72.300 ;
        RECT 60.470 72.240 60.790 72.500 ;
        RECT 66.910 72.440 67.230 72.500 ;
        RECT 73.900 72.440 74.040 72.640 ;
        RECT 74.745 72.640 77.350 72.780 ;
        RECT 74.745 72.595 75.035 72.640 ;
        RECT 77.030 72.580 77.350 72.640 ;
        RECT 82.090 72.780 82.410 72.840 ;
        RECT 83.945 72.780 84.235 72.825 ;
        RECT 86.690 72.780 87.010 72.840 ;
        RECT 82.090 72.640 83.700 72.780 ;
        RECT 82.090 72.580 82.410 72.640 ;
        RECT 77.490 72.440 77.810 72.500 ;
        RECT 83.560 72.440 83.700 72.640 ;
        RECT 83.945 72.640 87.010 72.780 ;
        RECT 83.945 72.595 84.235 72.640 ;
        RECT 86.690 72.580 87.010 72.640 ;
        RECT 66.910 72.300 72.200 72.440 ;
        RECT 73.900 72.300 77.260 72.440 ;
        RECT 66.910 72.240 67.230 72.300 ;
        RECT 47.145 71.915 47.435 72.145 ;
        RECT 47.590 71.900 47.910 72.160 ;
        RECT 51.745 72.100 52.035 72.145 ;
        RECT 54.045 72.100 54.335 72.145 ;
        RECT 51.745 71.960 54.335 72.100 ;
        RECT 51.745 71.915 52.035 71.960 ;
        RECT 54.045 71.915 54.335 71.960 ;
        RECT 66.465 72.100 66.755 72.145 ;
        RECT 68.290 72.100 68.610 72.160 ;
        RECT 66.465 71.960 68.610 72.100 ;
        RECT 66.465 71.915 66.755 71.960 ;
        RECT 68.290 71.900 68.610 71.960 ;
        RECT 72.060 72.100 72.200 72.300 ;
        RECT 77.120 72.145 77.260 72.300 ;
        RECT 77.490 72.300 83.240 72.440 ;
        RECT 83.560 72.300 86.460 72.440 ;
        RECT 77.490 72.240 77.810 72.300 ;
        RECT 72.060 71.960 75.880 72.100 ;
        RECT 37.025 71.620 41.840 71.760 ;
        RECT 42.095 71.760 42.385 71.805 ;
        RECT 44.615 71.760 44.905 71.805 ;
        RECT 45.805 71.760 46.095 71.805 ;
        RECT 49.445 71.760 49.735 71.805 ;
        RECT 42.095 71.620 46.095 71.760 ;
        RECT 37.025 71.575 37.315 71.620 ;
        RECT 21.385 71.280 27.120 71.420 ;
        RECT 28.745 71.420 29.035 71.465 ;
        RECT 31.030 71.420 31.350 71.480 ;
        RECT 28.745 71.280 31.350 71.420 ;
        RECT 21.385 71.235 21.675 71.280 ;
        RECT 28.745 71.235 29.035 71.280 ;
        RECT 31.030 71.220 31.350 71.280 ;
        RECT 22.290 71.080 22.610 71.140 ;
        RECT 23.670 71.080 23.990 71.140 ;
        RECT 21.000 70.940 23.990 71.080 ;
        RECT 22.290 70.880 22.610 70.940 ;
        RECT 23.670 70.880 23.990 70.940 ;
        RECT 24.145 71.080 24.435 71.125 ;
        RECT 24.590 71.080 24.910 71.140 ;
        RECT 24.145 70.940 24.910 71.080 ;
        RECT 24.145 70.895 24.435 70.940 ;
        RECT 24.590 70.880 24.910 70.940 ;
        RECT 30.110 71.080 30.430 71.140 ;
        RECT 30.585 71.080 30.875 71.125 ;
        RECT 30.110 70.940 30.875 71.080 ;
        RECT 30.110 70.880 30.430 70.940 ;
        RECT 30.585 70.895 30.875 70.940 ;
        RECT 33.330 71.080 33.650 71.140 ;
        RECT 33.880 71.080 34.020 71.575 ;
        RECT 41.150 71.560 41.470 71.620 ;
        RECT 42.095 71.575 42.385 71.620 ;
        RECT 44.615 71.575 44.905 71.620 ;
        RECT 45.805 71.575 46.095 71.620 ;
        RECT 47.680 71.620 49.735 71.760 ;
        RECT 47.680 71.480 47.820 71.620 ;
        RECT 49.445 71.575 49.735 71.620 ;
        RECT 52.190 71.560 52.510 71.820 ;
        RECT 53.110 71.560 53.430 71.820 ;
        RECT 56.330 71.760 56.650 71.820 ;
        RECT 56.805 71.760 57.095 71.805 ;
        RECT 56.330 71.620 57.095 71.760 ;
        RECT 56.330 71.560 56.650 71.620 ;
        RECT 56.805 71.575 57.095 71.620 ;
        RECT 61.405 71.575 61.695 71.805 ;
        RECT 36.550 71.420 36.870 71.480 ;
        RECT 39.785 71.420 40.075 71.465 ;
        RECT 36.550 71.280 40.075 71.420 ;
        RECT 36.550 71.220 36.870 71.280 ;
        RECT 39.785 71.235 40.075 71.280 ;
        RECT 42.530 71.420 42.820 71.465 ;
        RECT 44.100 71.420 44.390 71.465 ;
        RECT 46.200 71.420 46.490 71.465 ;
        RECT 42.530 71.280 46.490 71.420 ;
        RECT 42.530 71.235 42.820 71.280 ;
        RECT 44.100 71.235 44.390 71.280 ;
        RECT 46.200 71.235 46.490 71.280 ;
        RECT 47.590 71.220 47.910 71.480 ;
        RECT 55.870 71.420 56.190 71.480 ;
        RECT 61.480 71.420 61.620 71.575 ;
        RECT 66.910 71.560 67.230 71.820 ;
        RECT 69.670 71.760 69.990 71.820 ;
        RECT 72.060 71.805 72.200 71.960 ;
        RECT 71.065 71.760 71.355 71.805 ;
        RECT 69.670 71.620 71.355 71.760 ;
        RECT 69.670 71.560 69.990 71.620 ;
        RECT 71.065 71.575 71.355 71.620 ;
        RECT 71.985 71.575 72.275 71.805 ;
        RECT 74.730 71.760 75.050 71.820 ;
        RECT 75.740 71.805 75.880 71.960 ;
        RECT 77.045 71.915 77.335 72.145 ;
        RECT 78.410 72.100 78.730 72.160 ;
        RECT 80.725 72.100 81.015 72.145 ;
        RECT 78.410 71.960 81.015 72.100 ;
        RECT 78.410 71.900 78.730 71.960 ;
        RECT 80.725 71.915 81.015 71.960 ;
        RECT 81.170 71.900 81.490 72.160 ;
        RECT 83.100 72.145 83.240 72.300 ;
        RECT 82.105 71.915 82.395 72.145 ;
        RECT 83.025 71.915 83.315 72.145 ;
        RECT 84.405 72.100 84.695 72.145 ;
        RECT 84.850 72.100 85.170 72.160 ;
        RECT 84.405 71.960 85.170 72.100 ;
        RECT 84.405 71.915 84.695 71.960 ;
        RECT 75.205 71.760 75.495 71.805 ;
        RECT 74.730 71.620 75.495 71.760 ;
        RECT 74.730 71.560 75.050 71.620 ;
        RECT 75.205 71.575 75.495 71.620 ;
        RECT 75.665 71.575 75.955 71.805 ;
        RECT 79.790 71.560 80.110 71.820 ;
        RECT 80.250 71.760 80.570 71.820 ;
        RECT 82.180 71.760 82.320 71.915 ;
        RECT 80.250 71.620 82.320 71.760 ;
        RECT 82.550 71.760 82.870 71.820 ;
        RECT 84.480 71.760 84.620 71.915 ;
        RECT 84.850 71.900 85.170 71.960 ;
        RECT 85.310 71.900 85.630 72.160 ;
        RECT 85.770 71.900 86.090 72.160 ;
        RECT 86.320 72.145 86.460 72.300 ;
        RECT 86.245 71.915 86.535 72.145 ;
        RECT 82.550 71.620 84.620 71.760 ;
        RECT 80.250 71.560 80.570 71.620 ;
        RECT 82.550 71.560 82.870 71.620 ;
        RECT 55.870 71.280 61.620 71.420 ;
        RECT 68.290 71.420 68.610 71.480 ;
        RECT 72.905 71.420 73.195 71.465 ;
        RECT 68.290 71.280 73.195 71.420 ;
        RECT 55.870 71.220 56.190 71.280 ;
        RECT 68.290 71.220 68.610 71.280 ;
        RECT 72.905 71.235 73.195 71.280 ;
        RECT 74.270 71.420 74.590 71.480 ;
        RECT 87.165 71.420 87.455 71.465 ;
        RECT 74.270 71.280 87.455 71.420 ;
        RECT 74.270 71.220 74.590 71.280 ;
        RECT 87.165 71.235 87.455 71.280 ;
        RECT 33.330 70.940 34.020 71.080 ;
        RECT 34.250 71.080 34.570 71.140 ;
        RECT 41.610 71.080 41.930 71.140 ;
        RECT 47.130 71.080 47.450 71.140 ;
        RECT 34.250 70.940 47.450 71.080 ;
        RECT 33.330 70.880 33.650 70.940 ;
        RECT 34.250 70.880 34.570 70.940 ;
        RECT 41.610 70.880 41.930 70.940 ;
        RECT 47.130 70.880 47.450 70.940 ;
        RECT 48.050 71.080 48.370 71.140 ;
        RECT 49.905 71.080 50.195 71.125 ;
        RECT 48.050 70.940 50.195 71.080 ;
        RECT 48.050 70.880 48.370 70.940 ;
        RECT 49.905 70.895 50.195 70.940 ;
        RECT 64.150 70.880 64.470 71.140 ;
        RECT 67.830 71.080 68.150 71.140 ;
        RECT 68.765 71.080 69.055 71.125 ;
        RECT 67.830 70.940 69.055 71.080 ;
        RECT 67.830 70.880 68.150 70.940 ;
        RECT 68.765 70.895 69.055 70.940 ;
        RECT 77.490 71.080 77.810 71.140 ;
        RECT 80.710 71.080 81.030 71.140 ;
        RECT 77.490 70.940 81.030 71.080 ;
        RECT 77.490 70.880 77.810 70.940 ;
        RECT 80.710 70.880 81.030 70.940 ;
        RECT 12.100 70.260 89.840 70.740 ;
        RECT 16.785 70.060 17.075 70.105 ;
        RECT 22.305 70.060 22.595 70.105 ;
        RECT 22.750 70.060 23.070 70.120 ;
        RECT 32.410 70.060 32.730 70.120 ;
        RECT 16.785 69.920 19.760 70.060 ;
        RECT 16.785 69.875 17.075 69.920 ;
        RECT 16.860 69.380 17.000 69.875 ;
        RECT 15.020 69.240 17.000 69.380 ;
        RECT 19.620 69.380 19.760 69.920 ;
        RECT 22.305 69.920 23.070 70.060 ;
        RECT 22.305 69.875 22.595 69.920 ;
        RECT 22.750 69.860 23.070 69.920 ;
        RECT 30.660 69.920 32.730 70.060 ;
        RECT 21.830 69.720 22.150 69.780 ;
        RECT 24.145 69.720 24.435 69.765 ;
        RECT 21.830 69.580 24.435 69.720 ;
        RECT 21.830 69.520 22.150 69.580 ;
        RECT 24.145 69.535 24.435 69.580 ;
        RECT 27.365 69.720 27.655 69.765 ;
        RECT 30.660 69.720 30.800 69.920 ;
        RECT 32.410 69.860 32.730 69.920 ;
        RECT 35.170 70.060 35.490 70.120 ;
        RECT 37.945 70.060 38.235 70.105 ;
        RECT 35.170 69.920 38.235 70.060 ;
        RECT 35.170 69.860 35.490 69.920 ;
        RECT 37.945 69.875 38.235 69.920 ;
        RECT 40.690 70.060 41.010 70.120 ;
        RECT 47.605 70.060 47.895 70.105 ;
        RECT 40.690 69.920 47.895 70.060 ;
        RECT 40.690 69.860 41.010 69.920 ;
        RECT 47.605 69.875 47.895 69.920 ;
        RECT 52.190 70.060 52.510 70.120 ;
        RECT 52.665 70.060 52.955 70.105 ;
        RECT 52.190 69.920 52.955 70.060 ;
        RECT 27.365 69.580 30.800 69.720 ;
        RECT 31.070 69.720 31.360 69.765 ;
        RECT 33.170 69.720 33.460 69.765 ;
        RECT 34.740 69.720 35.030 69.765 ;
        RECT 31.070 69.580 35.030 69.720 ;
        RECT 27.365 69.535 27.655 69.580 ;
        RECT 31.070 69.535 31.360 69.580 ;
        RECT 33.170 69.535 33.460 69.580 ;
        RECT 34.740 69.535 35.030 69.580 ;
        RECT 41.190 69.720 41.480 69.765 ;
        RECT 43.290 69.720 43.580 69.765 ;
        RECT 44.860 69.720 45.150 69.765 ;
        RECT 41.190 69.580 45.150 69.720 ;
        RECT 41.190 69.535 41.480 69.580 ;
        RECT 43.290 69.535 43.580 69.580 ;
        RECT 44.860 69.535 45.150 69.580 ;
        RECT 19.990 69.380 20.310 69.440 ;
        RECT 19.620 69.240 20.310 69.380 ;
        RECT 15.020 69.085 15.160 69.240 ;
        RECT 14.945 68.855 15.235 69.085 ;
        RECT 15.405 69.040 15.695 69.085 ;
        RECT 19.070 69.040 19.390 69.100 ;
        RECT 19.620 69.085 19.760 69.240 ;
        RECT 19.990 69.180 20.310 69.240 ;
        RECT 15.405 68.900 19.390 69.040 ;
        RECT 15.405 68.855 15.695 68.900 ;
        RECT 14.010 68.700 14.330 68.760 ;
        RECT 16.860 68.745 17.000 68.900 ;
        RECT 19.070 68.840 19.390 68.900 ;
        RECT 19.545 68.855 19.835 69.085 ;
        RECT 21.920 69.040 22.060 69.520 ;
        RECT 23.670 69.380 23.990 69.440 ;
        RECT 24.605 69.380 24.895 69.425 ;
        RECT 23.670 69.240 24.895 69.380 ;
        RECT 23.670 69.180 23.990 69.240 ;
        RECT 24.605 69.195 24.895 69.240 ;
        RECT 31.465 69.380 31.755 69.425 ;
        RECT 32.655 69.380 32.945 69.425 ;
        RECT 35.175 69.380 35.465 69.425 ;
        RECT 31.465 69.240 35.465 69.380 ;
        RECT 31.465 69.195 31.755 69.240 ;
        RECT 32.655 69.195 32.945 69.240 ;
        RECT 35.175 69.195 35.465 69.240 ;
        RECT 37.470 69.380 37.790 69.440 ;
        RECT 41.585 69.380 41.875 69.425 ;
        RECT 42.775 69.380 43.065 69.425 ;
        RECT 45.295 69.380 45.585 69.425 ;
        RECT 37.470 69.240 40.460 69.380 ;
        RECT 37.470 69.180 37.790 69.240 ;
        RECT 20.080 68.900 22.060 69.040 ;
        RECT 20.080 68.745 20.220 68.900 ;
        RECT 23.225 68.855 23.515 69.085 ;
        RECT 29.205 69.040 29.495 69.085 ;
        RECT 29.650 69.040 29.970 69.100 ;
        RECT 29.205 68.900 29.970 69.040 ;
        RECT 29.205 68.855 29.495 68.900 ;
        RECT 15.865 68.700 16.155 68.745 ;
        RECT 14.010 68.560 16.155 68.700 ;
        RECT 16.860 68.560 17.155 68.745 ;
        RECT 20.005 68.700 20.295 68.745 ;
        RECT 14.010 68.500 14.330 68.560 ;
        RECT 15.865 68.515 16.155 68.560 ;
        RECT 16.865 68.515 17.155 68.560 ;
        RECT 17.320 68.560 20.295 68.700 ;
        RECT 14.515 68.360 14.805 68.405 ;
        RECT 15.390 68.360 15.710 68.420 ;
        RECT 14.515 68.220 15.710 68.360 ;
        RECT 15.940 68.360 16.080 68.515 ;
        RECT 17.320 68.360 17.460 68.560 ;
        RECT 20.005 68.515 20.295 68.560 ;
        RECT 20.450 68.700 20.770 68.760 ;
        RECT 20.925 68.700 21.215 68.745 ;
        RECT 23.300 68.700 23.440 68.855 ;
        RECT 29.650 68.840 29.970 68.900 ;
        RECT 30.570 68.840 30.890 69.100 ;
        RECT 37.010 69.040 37.330 69.100 ;
        RECT 40.320 69.085 40.460 69.240 ;
        RECT 41.585 69.240 45.585 69.380 ;
        RECT 41.585 69.195 41.875 69.240 ;
        RECT 42.775 69.195 43.065 69.240 ;
        RECT 45.295 69.195 45.585 69.240 ;
        RECT 38.865 69.040 39.155 69.085 ;
        RECT 36.180 68.900 39.155 69.040 ;
        RECT 25.970 68.700 26.290 68.760 ;
        RECT 20.450 68.560 26.290 68.700 ;
        RECT 20.450 68.500 20.770 68.560 ;
        RECT 20.925 68.515 21.215 68.560 ;
        RECT 25.970 68.500 26.290 68.560 ;
        RECT 28.285 68.700 28.575 68.745 ;
        RECT 30.125 68.700 30.415 68.745 ;
        RECT 31.030 68.700 31.350 68.760 ;
        RECT 28.285 68.560 29.880 68.700 ;
        RECT 28.285 68.515 28.575 68.560 ;
        RECT 15.940 68.220 17.460 68.360 ;
        RECT 14.515 68.175 14.805 68.220 ;
        RECT 15.390 68.160 15.710 68.220 ;
        RECT 17.690 68.160 18.010 68.420 ;
        RECT 18.150 68.160 18.470 68.420 ;
        RECT 22.290 68.360 22.610 68.420 ;
        RECT 26.430 68.360 26.750 68.420 ;
        RECT 22.290 68.220 26.750 68.360 ;
        RECT 22.290 68.160 22.610 68.220 ;
        RECT 26.430 68.160 26.750 68.220 ;
        RECT 28.730 68.160 29.050 68.420 ;
        RECT 29.740 68.360 29.880 68.560 ;
        RECT 30.125 68.560 31.350 68.700 ;
        RECT 30.125 68.515 30.415 68.560 ;
        RECT 31.030 68.500 31.350 68.560 ;
        RECT 31.920 68.700 32.210 68.745 ;
        RECT 32.870 68.700 33.190 68.760 ;
        RECT 31.920 68.560 33.190 68.700 ;
        RECT 31.920 68.515 32.210 68.560 ;
        RECT 32.870 68.500 33.190 68.560 ;
        RECT 35.630 68.360 35.950 68.420 ;
        RECT 36.180 68.360 36.320 68.900 ;
        RECT 37.010 68.840 37.330 68.900 ;
        RECT 38.865 68.855 39.155 68.900 ;
        RECT 40.245 68.855 40.535 69.085 ;
        RECT 40.705 69.040 40.995 69.085 ;
        RECT 46.670 69.040 46.990 69.100 ;
        RECT 40.705 68.900 46.990 69.040 ;
        RECT 47.680 69.040 47.820 69.875 ;
        RECT 52.190 69.860 52.510 69.920 ;
        RECT 52.665 69.875 52.955 69.920 ;
        RECT 56.805 70.060 57.095 70.105 ;
        RECT 60.010 70.060 60.330 70.120 ;
        RECT 56.805 69.920 60.330 70.060 ;
        RECT 56.805 69.875 57.095 69.920 ;
        RECT 60.010 69.860 60.330 69.920 ;
        RECT 65.085 70.060 65.375 70.105 ;
        RECT 81.630 70.060 81.950 70.120 ;
        RECT 65.085 69.920 81.950 70.060 ;
        RECT 65.085 69.875 65.375 69.920 ;
        RECT 81.630 69.860 81.950 69.920 ;
        RECT 59.550 69.720 59.840 69.765 ;
        RECT 61.120 69.720 61.410 69.765 ;
        RECT 63.220 69.720 63.510 69.765 ;
        RECT 59.550 69.580 63.510 69.720 ;
        RECT 59.550 69.535 59.840 69.580 ;
        RECT 61.120 69.535 61.410 69.580 ;
        RECT 63.220 69.535 63.510 69.580 ;
        RECT 66.950 69.720 67.240 69.765 ;
        RECT 69.050 69.720 69.340 69.765 ;
        RECT 70.620 69.720 70.910 69.765 ;
        RECT 66.950 69.580 70.910 69.720 ;
        RECT 66.950 69.535 67.240 69.580 ;
        RECT 69.050 69.535 69.340 69.580 ;
        RECT 70.620 69.535 70.910 69.580 ;
        RECT 73.365 69.720 73.655 69.765 ;
        RECT 76.570 69.720 76.890 69.780 ;
        RECT 79.790 69.720 80.110 69.780 ;
        RECT 73.365 69.580 80.110 69.720 ;
        RECT 73.365 69.535 73.655 69.580 ;
        RECT 76.570 69.520 76.890 69.580 ;
        RECT 79.790 69.520 80.110 69.580 ;
        RECT 55.410 69.180 55.730 69.440 ;
        RECT 59.115 69.380 59.405 69.425 ;
        RECT 61.635 69.380 61.925 69.425 ;
        RECT 62.825 69.380 63.115 69.425 ;
        RECT 65.530 69.380 65.850 69.440 ;
        RECT 59.115 69.240 63.115 69.380 ;
        RECT 59.115 69.195 59.405 69.240 ;
        RECT 61.635 69.195 61.925 69.240 ;
        RECT 62.825 69.195 63.115 69.240 ;
        RECT 63.320 69.240 65.850 69.380 ;
        RECT 48.985 69.040 49.275 69.085 ;
        RECT 47.680 68.900 49.275 69.040 ;
        RECT 40.705 68.855 40.995 68.900 ;
        RECT 46.670 68.840 46.990 68.900 ;
        RECT 48.985 68.855 49.275 68.900 ;
        RECT 52.190 68.840 52.510 69.100 ;
        RECT 54.505 69.040 54.795 69.085 ;
        RECT 56.790 69.040 57.110 69.100 ;
        RECT 54.505 68.900 57.110 69.040 ;
        RECT 54.505 68.855 54.795 68.900 ;
        RECT 56.790 68.840 57.110 68.900 ;
        RECT 62.425 69.040 62.715 69.085 ;
        RECT 63.320 69.040 63.460 69.240 ;
        RECT 65.530 69.180 65.850 69.240 ;
        RECT 66.450 69.180 66.770 69.440 ;
        RECT 67.345 69.380 67.635 69.425 ;
        RECT 68.535 69.380 68.825 69.425 ;
        RECT 71.055 69.380 71.345 69.425 ;
        RECT 67.345 69.240 71.345 69.380 ;
        RECT 67.345 69.195 67.635 69.240 ;
        RECT 68.535 69.195 68.825 69.240 ;
        RECT 71.055 69.195 71.345 69.240 ;
        RECT 74.270 69.380 74.590 69.440 ;
        RECT 83.010 69.380 83.330 69.440 ;
        RECT 86.230 69.380 86.550 69.440 ;
        RECT 74.270 69.240 86.550 69.380 ;
        RECT 74.270 69.180 74.590 69.240 ;
        RECT 83.010 69.180 83.330 69.240 ;
        RECT 86.230 69.180 86.550 69.240 ;
        RECT 62.425 68.900 63.460 69.040 ;
        RECT 62.425 68.855 62.715 68.900 ;
        RECT 63.690 68.840 64.010 69.100 ;
        RECT 65.990 68.840 66.310 69.100 ;
        RECT 66.540 69.040 66.680 69.180 ;
        RECT 73.825 69.040 74.115 69.085 ;
        RECT 76.110 69.040 76.430 69.100 ;
        RECT 77.045 69.040 77.335 69.085 ;
        RECT 66.540 68.900 75.420 69.040 ;
        RECT 73.825 68.855 74.115 68.900 ;
        RECT 36.550 68.700 36.870 68.760 ;
        RECT 42.040 68.700 42.330 68.745 ;
        RECT 42.990 68.700 43.310 68.760 ;
        RECT 67.830 68.745 68.150 68.760 ;
        RECT 36.550 68.560 40.460 68.700 ;
        RECT 36.550 68.500 36.870 68.560 ;
        RECT 37.485 68.360 37.775 68.405 ;
        RECT 29.740 68.220 37.775 68.360 ;
        RECT 35.630 68.160 35.950 68.220 ;
        RECT 37.485 68.175 37.775 68.220 ;
        RECT 39.770 68.160 40.090 68.420 ;
        RECT 40.320 68.360 40.460 68.560 ;
        RECT 42.040 68.560 43.310 68.700 ;
        RECT 42.040 68.515 42.330 68.560 ;
        RECT 42.990 68.500 43.310 68.560 ;
        RECT 48.065 68.515 48.355 68.745 ;
        RECT 67.800 68.515 68.150 68.745 ;
        RECT 75.280 68.700 75.420 68.900 ;
        RECT 76.110 68.900 77.335 69.040 ;
        RECT 76.110 68.840 76.430 68.900 ;
        RECT 77.045 68.855 77.335 68.900 ;
        RECT 77.490 69.040 77.810 69.100 ;
        RECT 83.485 69.040 83.775 69.085 ;
        RECT 77.490 68.900 83.775 69.040 ;
        RECT 77.490 68.840 77.810 68.900 ;
        RECT 83.485 68.855 83.775 68.900 ;
        RECT 83.930 68.840 84.250 69.100 ;
        RECT 84.405 69.040 84.695 69.085 ;
        RECT 84.850 69.040 85.170 69.100 ;
        RECT 84.405 68.900 85.170 69.040 ;
        RECT 84.405 68.855 84.695 68.900 ;
        RECT 84.850 68.840 85.170 68.900 ;
        RECT 85.310 68.840 85.630 69.100 ;
        RECT 79.330 68.700 79.650 68.760 ;
        RECT 80.725 68.700 81.015 68.745 ;
        RECT 81.170 68.700 81.490 68.760 ;
        RECT 75.280 68.560 81.490 68.700 ;
        RECT 48.140 68.360 48.280 68.515 ;
        RECT 67.830 68.500 68.150 68.515 ;
        RECT 79.330 68.500 79.650 68.560 ;
        RECT 80.725 68.515 81.015 68.560 ;
        RECT 81.170 68.500 81.490 68.560 ;
        RECT 85.785 68.515 86.075 68.745 ;
        RECT 86.690 68.700 87.010 68.760 ;
        RECT 88.530 68.700 88.850 68.760 ;
        RECT 86.690 68.560 88.850 68.700 ;
        RECT 40.320 68.220 48.280 68.360 ;
        RECT 49.890 68.160 50.210 68.420 ;
        RECT 51.730 68.160 52.050 68.420 ;
        RECT 54.965 68.360 55.255 68.405 ;
        RECT 60.010 68.360 60.330 68.420 ;
        RECT 54.965 68.220 60.330 68.360 ;
        RECT 54.965 68.175 55.255 68.220 ;
        RECT 60.010 68.160 60.330 68.220 ;
        RECT 65.070 68.360 65.390 68.420 ;
        RECT 76.110 68.360 76.430 68.420 ;
        RECT 65.070 68.220 76.430 68.360 ;
        RECT 65.070 68.160 65.390 68.220 ;
        RECT 76.110 68.160 76.430 68.220 ;
        RECT 77.030 68.360 77.350 68.420 ;
        RECT 80.250 68.360 80.570 68.420 ;
        RECT 77.030 68.220 80.570 68.360 ;
        RECT 77.030 68.160 77.350 68.220 ;
        RECT 80.250 68.160 80.570 68.220 ;
        RECT 82.105 68.360 82.395 68.405 ;
        RECT 82.550 68.360 82.870 68.420 ;
        RECT 82.105 68.220 82.870 68.360 ;
        RECT 82.105 68.175 82.395 68.220 ;
        RECT 82.550 68.160 82.870 68.220 ;
        RECT 84.390 68.360 84.710 68.420 ;
        RECT 85.860 68.360 86.000 68.515 ;
        RECT 86.690 68.500 87.010 68.560 ;
        RECT 88.530 68.500 88.850 68.560 ;
        RECT 84.390 68.220 86.000 68.360 ;
        RECT 84.390 68.160 84.710 68.220 ;
        RECT 87.610 68.160 87.930 68.420 ;
        RECT 12.100 67.540 89.840 68.020 ;
        RECT 13.565 67.340 13.855 67.385 ;
        RECT 14.010 67.340 14.330 67.400 ;
        RECT 13.565 67.200 14.330 67.340 ;
        RECT 13.565 67.155 13.855 67.200 ;
        RECT 14.010 67.140 14.330 67.200 ;
        RECT 17.690 67.340 18.010 67.400 ;
        RECT 20.910 67.340 21.230 67.400 ;
        RECT 24.145 67.340 24.435 67.385 ;
        RECT 17.690 67.200 21.230 67.340 ;
        RECT 17.690 67.140 18.010 67.200 ;
        RECT 20.910 67.140 21.230 67.200 ;
        RECT 21.460 67.200 24.435 67.340 ;
        RECT 15.850 67.000 16.170 67.060 ;
        RECT 21.460 67.000 21.600 67.200 ;
        RECT 24.145 67.155 24.435 67.200 ;
        RECT 26.430 67.340 26.750 67.400 ;
        RECT 28.285 67.340 28.575 67.385 ;
        RECT 26.430 67.200 28.575 67.340 ;
        RECT 26.430 67.140 26.750 67.200 ;
        RECT 28.285 67.155 28.575 67.200 ;
        RECT 28.730 67.340 29.050 67.400 ;
        RECT 31.030 67.340 31.350 67.400 ;
        RECT 28.730 67.200 31.350 67.340 ;
        RECT 28.730 67.140 29.050 67.200 ;
        RECT 31.030 67.140 31.350 67.200 ;
        RECT 31.505 67.340 31.795 67.385 ;
        RECT 32.870 67.340 33.190 67.400 ;
        RECT 31.505 67.200 33.190 67.340 ;
        RECT 31.505 67.155 31.795 67.200 ;
        RECT 32.870 67.140 33.190 67.200 ;
        RECT 36.565 67.340 36.855 67.385 ;
        RECT 37.470 67.340 37.790 67.400 ;
        RECT 36.565 67.200 37.790 67.340 ;
        RECT 36.565 67.155 36.855 67.200 ;
        RECT 37.470 67.140 37.790 67.200 ;
        RECT 42.215 67.340 42.505 67.385 ;
        RECT 49.890 67.340 50.210 67.400 ;
        RECT 42.215 67.200 50.210 67.340 ;
        RECT 42.215 67.155 42.505 67.200 ;
        RECT 49.890 67.140 50.210 67.200 ;
        RECT 56.345 67.340 56.635 67.385 ;
        RECT 60.470 67.340 60.790 67.400 ;
        RECT 56.345 67.200 60.790 67.340 ;
        RECT 56.345 67.155 56.635 67.200 ;
        RECT 60.470 67.140 60.790 67.200 ;
        RECT 65.990 67.340 66.310 67.400 ;
        RECT 74.270 67.340 74.590 67.400 ;
        RECT 65.990 67.200 74.590 67.340 ;
        RECT 65.990 67.140 66.310 67.200 ;
        RECT 74.270 67.140 74.590 67.200 ;
        RECT 74.745 67.340 75.035 67.385 ;
        RECT 75.190 67.340 75.510 67.400 ;
        RECT 82.090 67.340 82.410 67.400 ;
        RECT 74.745 67.200 75.510 67.340 ;
        RECT 74.745 67.155 75.035 67.200 ;
        RECT 75.190 67.140 75.510 67.200 ;
        RECT 75.740 67.200 82.410 67.340 ;
        RECT 15.850 66.860 21.600 67.000 ;
        RECT 21.765 67.000 22.055 67.045 ;
        RECT 22.290 67.000 22.610 67.060 ;
        RECT 21.765 66.860 22.610 67.000 ;
        RECT 15.850 66.800 16.170 66.860 ;
        RECT 21.765 66.815 22.055 66.860 ;
        RECT 22.290 66.800 22.610 66.860 ;
        RECT 22.750 66.800 23.070 67.060 ;
        RECT 30.570 67.000 30.890 67.060 ;
        RECT 23.300 66.860 30.890 67.000 ;
        RECT 19.185 66.660 19.475 66.705 ;
        RECT 20.465 66.680 20.755 66.705 ;
        RECT 20.465 66.660 21.600 66.680 ;
        RECT 23.300 66.660 23.440 66.860 ;
        RECT 30.570 66.800 30.890 66.860 ;
        RECT 31.950 67.000 32.270 67.060 ;
        RECT 32.425 67.000 32.715 67.045 ;
        RECT 31.950 66.860 32.715 67.000 ;
        RECT 31.950 66.800 32.270 66.860 ;
        RECT 32.425 66.815 32.715 66.860 ;
        RECT 38.850 67.000 39.170 67.060 ;
        RECT 41.165 67.000 41.455 67.045 ;
        RECT 38.850 66.860 41.455 67.000 ;
        RECT 38.850 66.800 39.170 66.860 ;
        RECT 41.165 66.815 41.455 66.860 ;
        RECT 47.100 67.000 47.390 67.045 ;
        RECT 48.050 67.000 48.370 67.060 ;
        RECT 47.100 66.860 48.370 67.000 ;
        RECT 47.100 66.815 47.390 66.860 ;
        RECT 48.050 66.800 48.370 66.860 ;
        RECT 55.870 66.800 56.190 67.060 ;
        RECT 62.020 67.000 62.310 67.045 ;
        RECT 64.150 67.000 64.470 67.060 ;
        RECT 68.290 67.045 68.610 67.060 ;
        RECT 68.260 67.000 68.610 67.045 ;
        RECT 62.020 66.860 64.470 67.000 ;
        RECT 68.095 66.860 68.610 67.000 ;
        RECT 62.020 66.815 62.310 66.860 ;
        RECT 64.150 66.800 64.470 66.860 ;
        RECT 68.260 66.815 68.610 66.860 ;
        RECT 68.290 66.800 68.610 66.815 ;
        RECT 19.185 66.520 20.220 66.660 ;
        RECT 19.185 66.475 19.475 66.520 ;
        RECT 15.875 66.320 16.165 66.365 ;
        RECT 18.395 66.320 18.685 66.365 ;
        RECT 19.585 66.320 19.875 66.365 ;
        RECT 15.875 66.180 19.875 66.320 ;
        RECT 20.080 66.320 20.220 66.520 ;
        RECT 20.465 66.540 23.440 66.660 ;
        RECT 20.465 66.475 20.755 66.540 ;
        RECT 21.460 66.520 23.440 66.540 ;
        RECT 23.670 66.460 23.990 66.720 ;
        RECT 24.130 66.660 24.450 66.720 ;
        RECT 25.525 66.660 25.815 66.705 ;
        RECT 24.130 66.520 25.815 66.660 ;
        RECT 24.130 66.460 24.450 66.520 ;
        RECT 25.525 66.475 25.815 66.520 ;
        RECT 26.430 66.660 26.750 66.720 ;
        RECT 26.905 66.660 27.195 66.705 ;
        RECT 26.430 66.520 27.195 66.660 ;
        RECT 26.430 66.460 26.750 66.520 ;
        RECT 26.905 66.475 27.195 66.520 ;
        RECT 27.350 66.460 27.670 66.720 ;
        RECT 28.745 66.475 29.035 66.705 ;
        RECT 29.665 66.660 29.955 66.705 ;
        RECT 29.280 66.520 29.955 66.660 ;
        RECT 28.820 66.320 28.960 66.475 ;
        RECT 20.080 66.180 21.140 66.320 ;
        RECT 15.875 66.135 16.165 66.180 ;
        RECT 18.395 66.135 18.685 66.180 ;
        RECT 19.585 66.135 19.875 66.180 ;
        RECT 21.000 66.025 21.140 66.180 ;
        RECT 21.460 66.180 28.960 66.320 ;
        RECT 16.310 65.980 16.600 66.025 ;
        RECT 17.880 65.980 18.170 66.025 ;
        RECT 19.980 65.980 20.270 66.025 ;
        RECT 16.310 65.840 20.270 65.980 ;
        RECT 16.310 65.795 16.600 65.840 ;
        RECT 17.880 65.795 18.170 65.840 ;
        RECT 19.980 65.795 20.270 65.840 ;
        RECT 20.925 65.795 21.215 66.025 ;
        RECT 21.460 65.700 21.600 66.180 ;
        RECT 25.970 65.980 26.290 66.040 ;
        RECT 29.280 65.980 29.420 66.520 ;
        RECT 29.665 66.475 29.955 66.520 ;
        RECT 30.110 66.460 30.430 66.720 ;
        RECT 34.265 66.660 34.555 66.705 ;
        RECT 32.960 66.520 34.555 66.660 ;
        RECT 25.970 65.840 29.420 65.980 ;
        RECT 30.200 65.980 30.340 66.460 ;
        RECT 32.960 66.040 33.100 66.520 ;
        RECT 34.265 66.475 34.555 66.520 ;
        RECT 35.630 66.460 35.950 66.720 ;
        RECT 37.025 66.475 37.315 66.705 ;
        RECT 39.785 66.660 40.075 66.705 ;
        RECT 42.070 66.660 42.390 66.720 ;
        RECT 39.785 66.520 42.390 66.660 ;
        RECT 39.785 66.475 40.075 66.520 ;
        RECT 34.710 66.320 35.030 66.380 ;
        RECT 37.100 66.320 37.240 66.475 ;
        RECT 42.070 66.460 42.390 66.520 ;
        RECT 45.765 66.660 46.055 66.705 ;
        RECT 46.210 66.660 46.530 66.720 ;
        RECT 45.765 66.520 46.530 66.660 ;
        RECT 45.765 66.475 46.055 66.520 ;
        RECT 46.210 66.460 46.530 66.520 ;
        RECT 48.510 66.660 48.830 66.720 ;
        RECT 48.510 66.520 51.040 66.660 ;
        RECT 48.510 66.460 48.830 66.520 ;
        RECT 50.900 66.380 51.040 66.520 ;
        RECT 53.110 66.460 53.430 66.720 ;
        RECT 54.030 66.460 54.350 66.720 ;
        RECT 63.245 66.660 63.535 66.705 ;
        RECT 63.690 66.660 64.010 66.720 ;
        RECT 66.910 66.660 67.230 66.720 ;
        RECT 75.740 66.705 75.880 67.200 ;
        RECT 82.090 67.140 82.410 67.200 ;
        RECT 80.710 67.000 81.030 67.060 ;
        RECT 76.660 66.860 81.030 67.000 ;
        RECT 63.245 66.520 67.230 66.660 ;
        RECT 63.245 66.475 63.535 66.520 ;
        RECT 63.690 66.460 64.010 66.520 ;
        RECT 66.910 66.460 67.230 66.520 ;
        RECT 75.665 66.475 75.955 66.705 ;
        RECT 76.110 66.660 76.430 66.720 ;
        RECT 76.660 66.705 76.800 66.860 ;
        RECT 80.710 66.800 81.030 66.860 ;
        RECT 76.585 66.660 76.875 66.705 ;
        RECT 76.110 66.520 76.875 66.660 ;
        RECT 76.110 66.460 76.430 66.520 ;
        RECT 76.585 66.475 76.875 66.520 ;
        RECT 77.030 66.460 77.350 66.720 ;
        RECT 78.410 66.660 78.730 66.720 ;
        RECT 77.580 66.520 78.730 66.660 ;
        RECT 34.710 66.180 37.240 66.320 ;
        RECT 46.645 66.320 46.935 66.365 ;
        RECT 47.835 66.320 48.125 66.365 ;
        RECT 50.355 66.320 50.645 66.365 ;
        RECT 46.645 66.180 50.645 66.320 ;
        RECT 34.710 66.120 35.030 66.180 ;
        RECT 46.645 66.135 46.935 66.180 ;
        RECT 47.835 66.135 48.125 66.180 ;
        RECT 50.355 66.135 50.645 66.180 ;
        RECT 50.810 66.320 51.130 66.380 ;
        RECT 54.120 66.320 54.260 66.460 ;
        RECT 50.810 66.180 54.260 66.320 ;
        RECT 58.655 66.320 58.945 66.365 ;
        RECT 61.175 66.320 61.465 66.365 ;
        RECT 62.365 66.320 62.655 66.365 ;
        RECT 58.655 66.180 62.655 66.320 ;
        RECT 50.810 66.120 51.130 66.180 ;
        RECT 58.655 66.135 58.945 66.180 ;
        RECT 61.175 66.135 61.465 66.180 ;
        RECT 62.365 66.135 62.655 66.180 ;
        RECT 67.805 66.320 68.095 66.365 ;
        RECT 68.995 66.320 69.285 66.365 ;
        RECT 71.515 66.320 71.805 66.365 ;
        RECT 67.805 66.180 71.805 66.320 ;
        RECT 67.805 66.135 68.095 66.180 ;
        RECT 68.995 66.135 69.285 66.180 ;
        RECT 71.515 66.135 71.805 66.180 ;
        RECT 32.870 65.980 33.190 66.040 ;
        RECT 30.200 65.840 33.190 65.980 ;
        RECT 25.970 65.780 26.290 65.840 ;
        RECT 32.870 65.780 33.190 65.840 ;
        RECT 40.705 65.980 40.995 66.025 ;
        RECT 42.530 65.980 42.850 66.040 ;
        RECT 40.705 65.840 42.850 65.980 ;
        RECT 40.705 65.795 40.995 65.840 ;
        RECT 42.530 65.780 42.850 65.840 ;
        RECT 42.990 65.780 43.310 66.040 ;
        RECT 46.250 65.980 46.540 66.025 ;
        RECT 48.350 65.980 48.640 66.025 ;
        RECT 49.920 65.980 50.210 66.025 ;
        RECT 46.250 65.840 50.210 65.980 ;
        RECT 46.250 65.795 46.540 65.840 ;
        RECT 48.350 65.795 48.640 65.840 ;
        RECT 49.920 65.795 50.210 65.840 ;
        RECT 59.090 65.980 59.380 66.025 ;
        RECT 60.660 65.980 60.950 66.025 ;
        RECT 62.760 65.980 63.050 66.025 ;
        RECT 59.090 65.840 63.050 65.980 ;
        RECT 59.090 65.795 59.380 65.840 ;
        RECT 60.660 65.795 60.950 65.840 ;
        RECT 62.760 65.795 63.050 65.840 ;
        RECT 67.410 65.980 67.700 66.025 ;
        RECT 69.510 65.980 69.800 66.025 ;
        RECT 71.080 65.980 71.370 66.025 ;
        RECT 67.410 65.840 71.370 65.980 ;
        RECT 67.410 65.795 67.700 65.840 ;
        RECT 69.510 65.795 69.800 65.840 ;
        RECT 71.080 65.795 71.370 65.840 ;
        RECT 73.825 65.980 74.115 66.025 ;
        RECT 76.570 65.980 76.890 66.040 ;
        RECT 73.825 65.840 76.890 65.980 ;
        RECT 73.825 65.795 74.115 65.840 ;
        RECT 76.570 65.780 76.890 65.840 ;
        RECT 21.370 65.440 21.690 65.700 ;
        RECT 21.830 65.640 22.150 65.700 ;
        RECT 23.670 65.640 23.990 65.700 ;
        RECT 21.830 65.500 23.990 65.640 ;
        RECT 21.830 65.440 22.150 65.500 ;
        RECT 23.670 65.440 23.990 65.500 ;
        RECT 24.130 65.640 24.450 65.700 ;
        RECT 28.745 65.640 29.035 65.685 ;
        RECT 24.130 65.500 29.035 65.640 ;
        RECT 24.130 65.440 24.450 65.500 ;
        RECT 28.745 65.455 29.035 65.500 ;
        RECT 32.425 65.640 32.715 65.685 ;
        RECT 34.725 65.640 35.015 65.685 ;
        RECT 32.425 65.500 35.015 65.640 ;
        RECT 32.425 65.455 32.715 65.500 ;
        RECT 34.725 65.455 35.015 65.500 ;
        RECT 41.150 65.640 41.470 65.700 ;
        RECT 42.085 65.640 42.375 65.685 ;
        RECT 41.150 65.500 42.375 65.640 ;
        RECT 41.150 65.440 41.470 65.500 ;
        RECT 42.085 65.455 42.375 65.500 ;
        RECT 52.650 65.640 52.970 65.700 ;
        RECT 56.330 65.640 56.650 65.700 ;
        RECT 52.650 65.500 56.650 65.640 ;
        RECT 77.580 65.640 77.720 66.520 ;
        RECT 78.410 66.460 78.730 66.520 ;
        RECT 79.345 66.475 79.635 66.705 ;
        RECT 77.950 66.320 78.270 66.380 ;
        RECT 79.420 66.320 79.560 66.475 ;
        RECT 81.170 66.460 81.490 66.720 ;
        RECT 82.465 66.660 82.755 66.705 ;
        RECT 81.720 66.520 82.755 66.660 ;
        RECT 77.950 66.180 79.560 66.320 ;
        RECT 80.710 66.320 81.030 66.380 ;
        RECT 81.720 66.320 81.860 66.520 ;
        RECT 82.465 66.475 82.755 66.520 ;
        RECT 80.710 66.180 81.860 66.320 ;
        RECT 82.065 66.320 82.355 66.365 ;
        RECT 83.255 66.320 83.545 66.365 ;
        RECT 85.775 66.320 86.065 66.365 ;
        RECT 82.065 66.180 86.065 66.320 ;
        RECT 77.950 66.120 78.270 66.180 ;
        RECT 80.710 66.120 81.030 66.180 ;
        RECT 82.065 66.135 82.355 66.180 ;
        RECT 83.255 66.135 83.545 66.180 ;
        RECT 85.775 66.135 86.065 66.180 ;
        RECT 81.670 65.980 81.960 66.025 ;
        RECT 83.770 65.980 84.060 66.025 ;
        RECT 85.340 65.980 85.630 66.025 ;
        RECT 81.670 65.840 85.630 65.980 ;
        RECT 81.670 65.795 81.960 65.840 ;
        RECT 83.770 65.795 84.060 65.840 ;
        RECT 85.340 65.795 85.630 65.840 ;
        RECT 77.965 65.640 78.255 65.685 ;
        RECT 77.580 65.500 78.255 65.640 ;
        RECT 52.650 65.440 52.970 65.500 ;
        RECT 56.330 65.440 56.650 65.500 ;
        RECT 77.965 65.455 78.255 65.500 ;
        RECT 78.410 65.640 78.730 65.700 ;
        RECT 80.265 65.640 80.555 65.685 ;
        RECT 78.410 65.500 80.555 65.640 ;
        RECT 78.410 65.440 78.730 65.500 ;
        RECT 80.265 65.455 80.555 65.500 ;
        RECT 82.090 65.640 82.410 65.700 ;
        RECT 86.690 65.640 87.010 65.700 ;
        RECT 88.085 65.640 88.375 65.685 ;
        RECT 82.090 65.500 88.375 65.640 ;
        RECT 82.090 65.440 82.410 65.500 ;
        RECT 86.690 65.440 87.010 65.500 ;
        RECT 88.085 65.455 88.375 65.500 ;
        RECT 12.100 64.820 89.840 65.300 ;
        RECT 15.390 64.620 15.710 64.680 ;
        RECT 15.390 64.480 18.840 64.620 ;
        RECT 15.390 64.420 15.710 64.480 ;
        RECT 14.050 64.280 14.340 64.325 ;
        RECT 16.150 64.280 16.440 64.325 ;
        RECT 17.720 64.280 18.010 64.325 ;
        RECT 14.050 64.140 18.010 64.280 ;
        RECT 14.050 64.095 14.340 64.140 ;
        RECT 16.150 64.095 16.440 64.140 ;
        RECT 17.720 64.095 18.010 64.140 ;
        RECT 14.445 63.940 14.735 63.985 ;
        RECT 15.635 63.940 15.925 63.985 ;
        RECT 18.155 63.940 18.445 63.985 ;
        RECT 14.445 63.800 18.445 63.940 ;
        RECT 18.700 63.940 18.840 64.480 ;
        RECT 20.450 64.420 20.770 64.680 ;
        RECT 20.925 64.620 21.215 64.665 ;
        RECT 22.290 64.620 22.610 64.680 ;
        RECT 20.925 64.480 22.610 64.620 ;
        RECT 20.925 64.435 21.215 64.480 ;
        RECT 22.290 64.420 22.610 64.480 ;
        RECT 32.870 64.420 33.190 64.680 ;
        RECT 33.805 64.620 34.095 64.665 ;
        RECT 35.170 64.620 35.490 64.680 ;
        RECT 37.470 64.620 37.790 64.680 ;
        RECT 33.805 64.480 37.790 64.620 ;
        RECT 33.805 64.435 34.095 64.480 ;
        RECT 35.170 64.420 35.490 64.480 ;
        RECT 37.470 64.420 37.790 64.480 ;
        RECT 49.430 64.620 49.750 64.680 ;
        RECT 49.430 64.480 50.120 64.620 ;
        RECT 49.430 64.420 49.750 64.480 ;
        RECT 28.745 64.280 29.035 64.325 ;
        RECT 29.650 64.280 29.970 64.340 ;
        RECT 28.745 64.140 29.970 64.280 ;
        RECT 28.745 64.095 29.035 64.140 ;
        RECT 29.650 64.080 29.970 64.140 ;
        RECT 30.125 63.940 30.415 63.985 ;
        RECT 39.310 63.940 39.630 64.000 ;
        RECT 18.700 63.800 21.140 63.940 ;
        RECT 14.445 63.755 14.735 63.800 ;
        RECT 15.635 63.755 15.925 63.800 ;
        RECT 18.155 63.755 18.445 63.800 ;
        RECT 13.565 63.600 13.855 63.645 ;
        RECT 20.450 63.600 20.770 63.660 ;
        RECT 21.000 63.645 21.140 63.800 ;
        RECT 30.125 63.800 39.630 63.940 ;
        RECT 49.980 63.940 50.120 64.480 ;
        RECT 51.270 64.420 51.590 64.680 ;
        RECT 52.190 64.620 52.510 64.680 ;
        RECT 55.425 64.620 55.715 64.665 ;
        RECT 52.190 64.480 55.715 64.620 ;
        RECT 52.190 64.420 52.510 64.480 ;
        RECT 55.425 64.435 55.715 64.480 ;
        RECT 56.345 64.620 56.635 64.665 ;
        RECT 59.090 64.620 59.410 64.680 ;
        RECT 72.890 64.620 73.210 64.680 ;
        RECT 56.345 64.480 59.410 64.620 ;
        RECT 56.345 64.435 56.635 64.480 ;
        RECT 59.090 64.420 59.410 64.480 ;
        RECT 61.020 64.480 73.210 64.620 ;
        RECT 50.365 64.280 50.655 64.325 ;
        RECT 54.950 64.280 55.270 64.340 ;
        RECT 50.365 64.140 55.270 64.280 ;
        RECT 50.365 64.095 50.655 64.140 ;
        RECT 54.950 64.080 55.270 64.140 ;
        RECT 53.255 63.940 53.545 63.985 ;
        RECT 61.020 63.940 61.160 64.480 ;
        RECT 72.890 64.420 73.210 64.480 ;
        RECT 73.365 64.620 73.655 64.665 ;
        RECT 73.810 64.620 74.130 64.680 ;
        RECT 73.365 64.480 74.130 64.620 ;
        RECT 73.365 64.435 73.655 64.480 ;
        RECT 73.810 64.420 74.130 64.480 ;
        RECT 77.490 64.620 77.810 64.680 ;
        RECT 79.330 64.620 79.650 64.680 ;
        RECT 77.490 64.480 79.650 64.620 ;
        RECT 77.490 64.420 77.810 64.480 ;
        RECT 79.330 64.420 79.650 64.480 ;
        RECT 80.710 64.420 81.030 64.680 ;
        RECT 87.610 64.620 87.930 64.680 ;
        RECT 81.260 64.480 87.930 64.620 ;
        RECT 81.260 64.280 81.400 64.480 ;
        RECT 87.610 64.420 87.930 64.480 ;
        RECT 78.500 64.140 81.400 64.280 ;
        RECT 81.670 64.280 81.960 64.325 ;
        RECT 83.770 64.280 84.060 64.325 ;
        RECT 85.340 64.280 85.630 64.325 ;
        RECT 81.670 64.140 85.630 64.280 ;
        RECT 76.110 63.940 76.430 64.000 ;
        RECT 49.980 63.800 52.420 63.940 ;
        RECT 30.125 63.755 30.415 63.800 ;
        RECT 39.310 63.740 39.630 63.800 ;
        RECT 13.565 63.460 20.770 63.600 ;
        RECT 13.565 63.415 13.855 63.460 ;
        RECT 20.450 63.400 20.770 63.460 ;
        RECT 20.925 63.415 21.215 63.645 ;
        RECT 21.845 63.415 22.135 63.645 ;
        RECT 27.350 63.600 27.670 63.660 ;
        RECT 28.285 63.600 28.575 63.645 ;
        RECT 27.350 63.460 28.575 63.600 ;
        RECT 14.930 63.305 15.250 63.320 ;
        RECT 14.900 63.075 15.250 63.305 ;
        RECT 14.930 63.060 15.250 63.075 ;
        RECT 17.690 63.260 18.010 63.320 ;
        RECT 21.920 63.260 22.060 63.415 ;
        RECT 27.350 63.400 27.670 63.460 ;
        RECT 28.285 63.415 28.575 63.460 ;
        RECT 29.190 63.400 29.510 63.660 ;
        RECT 29.665 63.415 29.955 63.645 ;
        RECT 30.585 63.600 30.875 63.645 ;
        RECT 31.030 63.600 31.350 63.660 ;
        RECT 35.170 63.600 35.490 63.660 ;
        RECT 52.280 63.645 52.420 63.800 ;
        RECT 53.255 63.800 61.160 63.940 ;
        RECT 72.980 63.800 76.430 63.940 ;
        RECT 53.255 63.755 53.545 63.800 ;
        RECT 30.585 63.460 35.490 63.600 ;
        RECT 30.585 63.415 30.875 63.460 ;
        RECT 17.690 63.120 22.060 63.260 ;
        RECT 22.290 63.260 22.610 63.320 ;
        RECT 25.510 63.260 25.830 63.320 ;
        RECT 22.290 63.120 25.830 63.260 ;
        RECT 29.740 63.260 29.880 63.415 ;
        RECT 31.030 63.400 31.350 63.460 ;
        RECT 35.170 63.400 35.490 63.460 ;
        RECT 52.205 63.600 52.495 63.645 ;
        RECT 52.650 63.600 52.970 63.660 ;
        RECT 52.205 63.460 52.970 63.600 ;
        RECT 52.205 63.415 52.495 63.460 ;
        RECT 52.650 63.400 52.970 63.460 ;
        RECT 54.030 63.400 54.350 63.660 ;
        RECT 57.710 63.600 58.030 63.660 ;
        RECT 65.070 63.600 65.390 63.660 ;
        RECT 72.980 63.645 73.120 63.800 ;
        RECT 76.110 63.740 76.430 63.800 ;
        RECT 57.710 63.460 65.390 63.600 ;
        RECT 57.710 63.400 58.030 63.460 ;
        RECT 65.070 63.400 65.390 63.460 ;
        RECT 72.905 63.415 73.195 63.645 ;
        RECT 73.825 63.600 74.115 63.645 ;
        RECT 75.205 63.600 75.495 63.645 ;
        RECT 75.650 63.600 75.970 63.660 ;
        RECT 78.500 63.645 78.640 64.140 ;
        RECT 81.670 64.095 81.960 64.140 ;
        RECT 83.770 64.095 84.060 64.140 ;
        RECT 85.340 64.095 85.630 64.140 ;
        RECT 86.230 64.280 86.550 64.340 ;
        RECT 88.085 64.280 88.375 64.325 ;
        RECT 86.230 64.140 88.375 64.280 ;
        RECT 86.230 64.080 86.550 64.140 ;
        RECT 88.085 64.095 88.375 64.140 ;
        RECT 81.170 63.740 81.490 64.000 ;
        RECT 82.065 63.940 82.355 63.985 ;
        RECT 83.255 63.940 83.545 63.985 ;
        RECT 85.775 63.940 86.065 63.985 ;
        RECT 82.065 63.800 86.065 63.940 ;
        RECT 82.065 63.755 82.355 63.800 ;
        RECT 83.255 63.755 83.545 63.800 ;
        RECT 85.775 63.755 86.065 63.800 ;
        RECT 73.825 63.460 75.970 63.600 ;
        RECT 73.825 63.415 74.115 63.460 ;
        RECT 75.205 63.415 75.495 63.460 ;
        RECT 75.650 63.400 75.970 63.460 ;
        RECT 77.505 63.415 77.795 63.645 ;
        RECT 78.425 63.415 78.715 63.645 ;
        RECT 30.110 63.260 30.430 63.320 ;
        RECT 33.725 63.260 34.015 63.305 ;
        RECT 34.250 63.260 34.570 63.320 ;
        RECT 29.740 63.120 34.570 63.260 ;
        RECT 17.690 63.060 18.010 63.120 ;
        RECT 22.290 63.060 22.610 63.120 ;
        RECT 25.510 63.060 25.830 63.120 ;
        RECT 30.110 63.060 30.430 63.120 ;
        RECT 33.725 63.075 34.015 63.120 ;
        RECT 34.250 63.060 34.570 63.120 ;
        RECT 34.725 63.260 35.015 63.305 ;
        RECT 35.630 63.260 35.950 63.320 ;
        RECT 34.725 63.120 35.950 63.260 ;
        RECT 34.725 63.075 35.015 63.120 ;
        RECT 35.630 63.060 35.950 63.120 ;
        RECT 48.525 63.260 48.815 63.305 ;
        RECT 50.810 63.260 51.130 63.320 ;
        RECT 48.525 63.120 51.130 63.260 ;
        RECT 48.525 63.075 48.815 63.120 ;
        RECT 50.810 63.060 51.130 63.120 ;
        RECT 51.730 63.260 52.050 63.320 ;
        RECT 54.505 63.260 54.795 63.305 ;
        RECT 66.910 63.260 67.230 63.320 ;
        RECT 68.765 63.260 69.055 63.305 ;
        RECT 51.730 63.120 54.260 63.260 ;
        RECT 51.730 63.060 52.050 63.120 ;
        RECT 16.770 62.920 17.090 62.980 ;
        RECT 19.530 62.920 19.850 62.980 ;
        RECT 16.770 62.780 19.850 62.920 ;
        RECT 16.770 62.720 17.090 62.780 ;
        RECT 19.530 62.720 19.850 62.780 ;
        RECT 30.570 62.920 30.890 62.980 ;
        RECT 31.950 62.920 32.270 62.980 ;
        RECT 47.130 62.920 47.450 62.980 ;
        RECT 30.570 62.780 47.450 62.920 ;
        RECT 30.570 62.720 30.890 62.780 ;
        RECT 31.950 62.720 32.270 62.780 ;
        RECT 47.130 62.720 47.450 62.780 ;
        RECT 49.575 62.920 49.865 62.965 ;
        RECT 50.350 62.920 50.670 62.980 ;
        RECT 52.190 62.920 52.510 62.980 ;
        RECT 49.575 62.780 52.510 62.920 ;
        RECT 54.120 62.920 54.260 63.120 ;
        RECT 54.505 63.120 64.840 63.260 ;
        RECT 54.505 63.075 54.795 63.120 ;
        RECT 55.505 62.920 55.795 62.965 ;
        RECT 54.120 62.780 55.795 62.920 ;
        RECT 64.700 62.920 64.840 63.120 ;
        RECT 66.910 63.120 69.055 63.260 ;
        RECT 66.910 63.060 67.230 63.120 ;
        RECT 68.765 63.075 69.055 63.120 ;
        RECT 74.285 63.260 74.575 63.305 ;
        RECT 76.110 63.260 76.430 63.320 ;
        RECT 74.285 63.120 76.430 63.260 ;
        RECT 74.285 63.075 74.575 63.120 ;
        RECT 76.110 63.060 76.430 63.120 ;
        RECT 70.130 62.920 70.450 62.980 ;
        RECT 77.030 62.920 77.350 62.980 ;
        RECT 77.580 62.920 77.720 63.415 ;
        RECT 78.870 63.400 79.190 63.660 ;
        RECT 79.330 63.400 79.650 63.660 ;
        RECT 82.550 63.645 82.870 63.660 ;
        RECT 82.520 63.600 82.870 63.645 ;
        RECT 82.355 63.460 82.870 63.600 ;
        RECT 82.520 63.415 82.870 63.460 ;
        RECT 82.550 63.400 82.870 63.415 ;
        RECT 77.950 63.260 78.270 63.320 ;
        RECT 83.010 63.260 83.330 63.320 ;
        RECT 77.950 63.120 83.330 63.260 ;
        RECT 77.950 63.060 78.270 63.120 ;
        RECT 83.010 63.060 83.330 63.120 ;
        RECT 85.310 62.920 85.630 62.980 ;
        RECT 64.700 62.780 85.630 62.920 ;
        RECT 49.575 62.735 49.865 62.780 ;
        RECT 50.350 62.720 50.670 62.780 ;
        RECT 52.190 62.720 52.510 62.780 ;
        RECT 55.505 62.735 55.795 62.780 ;
        RECT 70.130 62.720 70.450 62.780 ;
        RECT 77.030 62.720 77.350 62.780 ;
        RECT 85.310 62.720 85.630 62.780 ;
        RECT 12.100 62.100 89.840 62.580 ;
        RECT 14.930 61.700 15.250 61.960 ;
        RECT 22.750 61.900 23.070 61.960 ;
        RECT 17.780 61.760 23.070 61.900 ;
        RECT 15.785 61.560 16.075 61.605 ;
        RECT 15.785 61.420 16.540 61.560 ;
        RECT 15.785 61.375 16.075 61.420 ;
        RECT 16.400 60.880 16.540 61.420 ;
        RECT 16.770 61.360 17.090 61.620 ;
        RECT 17.780 61.265 17.920 61.760 ;
        RECT 22.750 61.700 23.070 61.760 ;
        RECT 42.530 61.900 42.850 61.960 ;
        RECT 43.925 61.900 44.215 61.945 ;
        RECT 42.530 61.760 44.215 61.900 ;
        RECT 42.530 61.700 42.850 61.760 ;
        RECT 43.925 61.715 44.215 61.760 ;
        RECT 74.730 61.700 75.050 61.960 ;
        RECT 81.630 61.900 81.950 61.960 ;
        RECT 75.740 61.760 81.950 61.900 ;
        RECT 18.625 61.560 18.915 61.605 ;
        RECT 19.530 61.560 19.850 61.620 ;
        RECT 18.625 61.420 19.850 61.560 ;
        RECT 18.625 61.375 18.915 61.420 ;
        RECT 19.530 61.360 19.850 61.420 ;
        RECT 35.170 61.360 35.490 61.620 ;
        RECT 44.845 61.560 45.135 61.605 ;
        RECT 49.890 61.560 50.210 61.620 ;
        RECT 44.845 61.420 50.210 61.560 ;
        RECT 44.845 61.375 45.135 61.420 ;
        RECT 49.890 61.360 50.210 61.420 ;
        RECT 52.205 61.560 52.495 61.605 ;
        RECT 52.205 61.420 55.180 61.560 ;
        RECT 52.205 61.375 52.495 61.420 ;
        RECT 17.705 61.035 17.995 61.265 ;
        RECT 18.150 61.220 18.470 61.280 ;
        RECT 19.085 61.220 19.375 61.265 ;
        RECT 18.150 61.080 19.375 61.220 ;
        RECT 18.150 61.020 18.470 61.080 ;
        RECT 19.085 61.035 19.375 61.080 ;
        RECT 20.005 61.220 20.295 61.265 ;
        RECT 24.130 61.220 24.450 61.280 ;
        RECT 20.005 61.080 24.450 61.220 ;
        RECT 20.005 61.035 20.295 61.080 ;
        RECT 24.130 61.020 24.450 61.080 ;
        RECT 26.890 61.020 27.210 61.280 ;
        RECT 30.110 61.020 30.430 61.280 ;
        RECT 31.490 61.020 31.810 61.280 ;
        RECT 33.345 61.035 33.635 61.265 ;
        RECT 34.265 61.220 34.555 61.265 ;
        RECT 34.710 61.220 35.030 61.280 ;
        RECT 34.265 61.080 35.030 61.220 ;
        RECT 34.265 61.035 34.555 61.080 ;
        RECT 19.545 60.880 19.835 60.925 ;
        RECT 16.400 60.740 19.835 60.880 ;
        RECT 31.580 60.880 31.720 61.020 ;
        RECT 32.870 60.880 33.190 60.940 ;
        RECT 31.580 60.740 33.190 60.880 ;
        RECT 19.545 60.695 19.835 60.740 ;
        RECT 32.870 60.680 33.190 60.740 ;
        RECT 23.670 60.540 23.990 60.600 ;
        RECT 26.905 60.540 27.195 60.585 ;
        RECT 23.670 60.400 27.195 60.540 ;
        RECT 23.670 60.340 23.990 60.400 ;
        RECT 26.905 60.355 27.195 60.400 ;
        RECT 29.190 60.540 29.510 60.600 ;
        RECT 30.570 60.540 30.890 60.600 ;
        RECT 33.420 60.540 33.560 61.035 ;
        RECT 34.710 61.020 35.030 61.080 ;
        RECT 43.450 61.020 43.770 61.280 ;
        RECT 48.065 61.035 48.355 61.265 ;
        RECT 48.985 61.220 49.275 61.265 ;
        RECT 51.730 61.220 52.050 61.280 ;
        RECT 55.040 61.265 55.180 61.420 ;
        RECT 48.985 61.080 52.050 61.220 ;
        RECT 48.985 61.035 49.275 61.080 ;
        RECT 48.140 60.880 48.280 61.035 ;
        RECT 51.730 61.020 52.050 61.080 ;
        RECT 53.125 61.220 53.415 61.265 ;
        RECT 54.965 61.220 55.255 61.265 ;
        RECT 55.410 61.220 55.730 61.280 ;
        RECT 53.125 61.080 54.720 61.220 ;
        RECT 53.125 61.035 53.415 61.080 ;
        RECT 49.430 60.880 49.750 60.940 ;
        RECT 48.140 60.740 49.750 60.880 ;
        RECT 49.430 60.680 49.750 60.740 ;
        RECT 50.810 60.880 51.130 60.940 ;
        RECT 53.585 60.880 53.875 60.925 ;
        RECT 50.810 60.740 53.875 60.880 ;
        RECT 54.580 60.880 54.720 61.080 ;
        RECT 54.965 61.080 55.730 61.220 ;
        RECT 54.965 61.035 55.255 61.080 ;
        RECT 55.410 61.020 55.730 61.080 ;
        RECT 66.910 61.020 67.230 61.280 ;
        RECT 75.740 61.265 75.880 61.760 ;
        RECT 81.630 61.700 81.950 61.760 ;
        RECT 83.010 61.900 83.330 61.960 ;
        RECT 85.770 61.900 86.090 61.960 ;
        RECT 88.085 61.900 88.375 61.945 ;
        RECT 83.010 61.760 88.375 61.900 ;
        RECT 83.010 61.700 83.330 61.760 ;
        RECT 85.770 61.700 86.090 61.760 ;
        RECT 88.085 61.715 88.375 61.760 ;
        RECT 80.725 61.560 81.015 61.605 ;
        RECT 82.410 61.560 82.700 61.605 ;
        RECT 80.725 61.420 82.700 61.560 ;
        RECT 80.725 61.375 81.015 61.420 ;
        RECT 82.410 61.375 82.700 61.420 ;
        RECT 73.825 61.035 74.115 61.265 ;
        RECT 75.665 61.035 75.955 61.265 ;
        RECT 77.030 61.220 77.350 61.280 ;
        RECT 77.505 61.220 77.795 61.265 ;
        RECT 77.030 61.080 77.795 61.220 ;
        RECT 59.090 60.880 59.410 60.940 ;
        RECT 54.580 60.740 59.410 60.880 ;
        RECT 73.900 60.880 74.040 61.035 ;
        RECT 77.030 61.020 77.350 61.080 ;
        RECT 77.505 61.035 77.795 61.080 ;
        RECT 78.410 61.020 78.730 61.280 ;
        RECT 78.870 61.020 79.190 61.280 ;
        RECT 79.345 61.220 79.635 61.265 ;
        RECT 83.930 61.220 84.250 61.280 ;
        RECT 79.345 61.080 84.250 61.220 ;
        RECT 79.345 61.035 79.635 61.080 ;
        RECT 83.930 61.020 84.250 61.080 ;
        RECT 80.710 60.880 81.030 60.940 ;
        RECT 73.900 60.740 81.030 60.880 ;
        RECT 50.810 60.680 51.130 60.740 ;
        RECT 53.585 60.695 53.875 60.740 ;
        RECT 59.090 60.680 59.410 60.740 ;
        RECT 80.710 60.680 81.030 60.740 ;
        RECT 81.170 60.680 81.490 60.940 ;
        RECT 82.065 60.880 82.355 60.925 ;
        RECT 83.255 60.880 83.545 60.925 ;
        RECT 85.775 60.880 86.065 60.925 ;
        RECT 82.065 60.740 86.065 60.880 ;
        RECT 82.065 60.695 82.355 60.740 ;
        RECT 83.255 60.695 83.545 60.740 ;
        RECT 85.775 60.695 86.065 60.740 ;
        RECT 29.190 60.400 33.560 60.540 ;
        RECT 47.590 60.540 47.910 60.600 ;
        RECT 54.045 60.540 54.335 60.585 ;
        RECT 47.590 60.400 54.335 60.540 ;
        RECT 29.190 60.340 29.510 60.400 ;
        RECT 30.570 60.340 30.890 60.400 ;
        RECT 47.590 60.340 47.910 60.400 ;
        RECT 54.045 60.355 54.335 60.400 ;
        RECT 72.905 60.540 73.195 60.585 ;
        RECT 81.670 60.540 81.960 60.585 ;
        RECT 83.770 60.540 84.060 60.585 ;
        RECT 85.340 60.540 85.630 60.585 ;
        RECT 72.905 60.400 81.400 60.540 ;
        RECT 72.905 60.355 73.195 60.400 ;
        RECT 15.850 60.000 16.170 60.260 ;
        RECT 36.090 60.000 36.410 60.260 ;
        RECT 44.830 60.000 45.150 60.260 ;
        RECT 48.970 60.000 49.290 60.260 ;
        RECT 51.285 60.200 51.575 60.245 ;
        RECT 52.190 60.200 52.510 60.260 ;
        RECT 51.285 60.060 52.510 60.200 ;
        RECT 51.285 60.015 51.575 60.060 ;
        RECT 52.190 60.000 52.510 60.060 ;
        RECT 54.505 60.200 54.795 60.245 ;
        RECT 61.390 60.200 61.710 60.260 ;
        RECT 54.505 60.060 61.710 60.200 ;
        RECT 54.505 60.015 54.795 60.060 ;
        RECT 61.390 60.000 61.710 60.060 ;
        RECT 76.125 60.200 76.415 60.245 ;
        RECT 76.570 60.200 76.890 60.260 ;
        RECT 76.125 60.060 76.890 60.200 ;
        RECT 81.260 60.200 81.400 60.400 ;
        RECT 81.670 60.400 85.630 60.540 ;
        RECT 81.670 60.355 81.960 60.400 ;
        RECT 83.770 60.355 84.060 60.400 ;
        RECT 85.340 60.355 85.630 60.400 ;
        RECT 82.550 60.200 82.870 60.260 ;
        RECT 81.260 60.060 82.870 60.200 ;
        RECT 76.125 60.015 76.415 60.060 ;
        RECT 76.570 60.000 76.890 60.060 ;
        RECT 82.550 60.000 82.870 60.060 ;
        RECT 12.100 59.380 89.840 59.860 ;
        RECT 22.305 59.180 22.595 59.225 ;
        RECT 22.750 59.180 23.070 59.240 ;
        RECT 22.305 59.040 23.070 59.180 ;
        RECT 22.305 58.995 22.595 59.040 ;
        RECT 22.750 58.980 23.070 59.040 ;
        RECT 32.885 59.180 33.175 59.225 ;
        RECT 35.170 59.180 35.490 59.240 ;
        RECT 32.885 59.040 35.490 59.180 ;
        RECT 32.885 58.995 33.175 59.040 ;
        RECT 35.170 58.980 35.490 59.040 ;
        RECT 42.085 59.180 42.375 59.225 ;
        RECT 42.530 59.180 42.850 59.240 ;
        RECT 42.085 59.040 42.850 59.180 ;
        RECT 42.085 58.995 42.375 59.040 ;
        RECT 42.530 58.980 42.850 59.040 ;
        RECT 43.005 59.180 43.295 59.225 ;
        RECT 46.210 59.180 46.530 59.240 ;
        RECT 43.005 59.040 46.530 59.180 ;
        RECT 43.005 58.995 43.295 59.040 ;
        RECT 46.210 58.980 46.530 59.040 ;
        RECT 46.685 59.180 46.975 59.225 ;
        RECT 49.890 59.180 50.210 59.240 ;
        RECT 46.685 59.040 50.210 59.180 ;
        RECT 46.685 58.995 46.975 59.040 ;
        RECT 49.890 58.980 50.210 59.040 ;
        RECT 50.350 58.980 50.670 59.240 ;
        RECT 71.525 59.180 71.815 59.225 ;
        RECT 83.010 59.180 83.330 59.240 ;
        RECT 71.525 59.040 83.330 59.180 ;
        RECT 71.525 58.995 71.815 59.040 ;
        RECT 83.010 58.980 83.330 59.040 ;
        RECT 87.625 59.180 87.915 59.225 ;
        RECT 88.070 59.180 88.390 59.240 ;
        RECT 87.625 59.040 88.390 59.180 ;
        RECT 87.625 58.995 87.915 59.040 ;
        RECT 88.070 58.980 88.390 59.040 ;
        RECT 35.630 58.840 35.920 58.885 ;
        RECT 37.200 58.840 37.490 58.885 ;
        RECT 39.300 58.840 39.590 58.885 ;
        RECT 35.630 58.700 39.590 58.840 ;
        RECT 35.630 58.655 35.920 58.700 ;
        RECT 37.200 58.655 37.490 58.700 ;
        RECT 39.300 58.655 39.590 58.700 ;
        RECT 47.130 58.640 47.450 58.900 ;
        RECT 51.285 58.840 51.575 58.885 ;
        RECT 48.600 58.700 51.575 58.840 ;
        RECT 20.450 58.500 20.770 58.560 ;
        RECT 26.430 58.500 26.750 58.560 ;
        RECT 28.285 58.500 28.575 58.545 ;
        RECT 20.450 58.360 28.575 58.500 ;
        RECT 20.450 58.300 20.770 58.360 ;
        RECT 26.430 58.300 26.750 58.360 ;
        RECT 28.285 58.315 28.575 58.360 ;
        RECT 35.195 58.500 35.485 58.545 ;
        RECT 37.715 58.500 38.005 58.545 ;
        RECT 38.905 58.500 39.195 58.545 ;
        RECT 35.195 58.360 39.195 58.500 ;
        RECT 35.195 58.315 35.485 58.360 ;
        RECT 37.715 58.315 38.005 58.360 ;
        RECT 38.905 58.315 39.195 58.360 ;
        RECT 23.210 57.960 23.530 58.220 ;
        RECT 24.590 57.960 24.910 58.220 ;
        RECT 30.110 58.160 30.430 58.220 ;
        RECT 26.060 58.020 30.430 58.160 ;
        RECT 24.145 57.820 24.435 57.865 ;
        RECT 26.060 57.820 26.200 58.020 ;
        RECT 30.110 57.960 30.430 58.020 ;
        RECT 32.425 58.160 32.715 58.205 ;
        RECT 33.790 58.160 34.110 58.220 ;
        RECT 32.425 58.020 34.110 58.160 ;
        RECT 32.425 57.975 32.715 58.020 ;
        RECT 33.790 57.960 34.110 58.020 ;
        RECT 39.770 57.960 40.090 58.220 ;
        RECT 40.245 58.160 40.535 58.205 ;
        RECT 41.150 58.160 41.470 58.220 ;
        RECT 43.465 58.160 43.755 58.205 ;
        RECT 40.245 58.020 43.755 58.160 ;
        RECT 40.245 57.975 40.535 58.020 ;
        RECT 41.150 57.960 41.470 58.020 ;
        RECT 43.465 57.975 43.755 58.020 ;
        RECT 47.145 58.160 47.435 58.205 ;
        RECT 48.050 58.160 48.370 58.220 ;
        RECT 48.600 58.205 48.740 58.700 ;
        RECT 51.285 58.655 51.575 58.700 ;
        RECT 62.810 58.840 63.100 58.885 ;
        RECT 64.910 58.840 65.200 58.885 ;
        RECT 66.480 58.840 66.770 58.885 ;
        RECT 77.030 58.840 77.350 58.900 ;
        RECT 62.810 58.700 66.770 58.840 ;
        RECT 62.810 58.655 63.100 58.700 ;
        RECT 64.910 58.655 65.200 58.700 ;
        RECT 66.480 58.655 66.770 58.700 ;
        RECT 74.820 58.700 77.350 58.840 ;
        RECT 48.970 58.500 49.290 58.560 ;
        RECT 54.045 58.500 54.335 58.545 ;
        RECT 48.970 58.360 54.335 58.500 ;
        RECT 48.970 58.300 49.290 58.360 ;
        RECT 54.045 58.315 54.335 58.360 ;
        RECT 63.205 58.500 63.495 58.545 ;
        RECT 64.395 58.500 64.685 58.545 ;
        RECT 66.915 58.500 67.205 58.545 ;
        RECT 63.205 58.360 67.205 58.500 ;
        RECT 63.205 58.315 63.495 58.360 ;
        RECT 64.395 58.315 64.685 58.360 ;
        RECT 66.915 58.315 67.205 58.360 ;
        RECT 71.050 58.500 71.370 58.560 ;
        RECT 71.050 58.360 74.500 58.500 ;
        RECT 71.050 58.300 71.370 58.360 ;
        RECT 47.145 58.020 48.370 58.160 ;
        RECT 47.145 57.975 47.435 58.020 ;
        RECT 48.050 57.960 48.370 58.020 ;
        RECT 48.525 57.975 48.815 58.205 ;
        RECT 49.430 57.960 49.750 58.220 ;
        RECT 50.365 58.160 50.655 58.205 ;
        RECT 52.190 58.160 52.510 58.220 ;
        RECT 49.980 58.020 52.510 58.160 ;
        RECT 24.145 57.680 26.200 57.820 ;
        RECT 26.445 57.820 26.735 57.865 ;
        RECT 31.030 57.820 31.350 57.880 ;
        RECT 26.445 57.680 31.350 57.820 ;
        RECT 24.145 57.635 24.435 57.680 ;
        RECT 26.445 57.635 26.735 57.680 ;
        RECT 31.030 57.620 31.350 57.680 ;
        RECT 38.390 57.865 38.710 57.880 ;
        RECT 38.390 57.635 38.740 57.865 ;
        RECT 42.085 57.820 42.375 57.865 ;
        RECT 42.085 57.680 43.680 57.820 ;
        RECT 42.085 57.635 42.375 57.680 ;
        RECT 38.390 57.620 38.710 57.635 ;
        RECT 43.540 57.540 43.680 57.680 ;
        RECT 26.905 57.480 27.195 57.525 ;
        RECT 29.190 57.480 29.510 57.540 ;
        RECT 38.850 57.480 39.170 57.540 ;
        RECT 26.905 57.340 39.170 57.480 ;
        RECT 26.905 57.295 27.195 57.340 ;
        RECT 29.190 57.280 29.510 57.340 ;
        RECT 38.850 57.280 39.170 57.340 ;
        RECT 43.450 57.280 43.770 57.540 ;
        RECT 48.065 57.480 48.355 57.525 ;
        RECT 49.980 57.480 50.120 58.020 ;
        RECT 50.365 57.975 50.655 58.020 ;
        RECT 52.190 57.960 52.510 58.020 ;
        RECT 59.090 57.960 59.410 58.220 ;
        RECT 62.325 58.160 62.615 58.205 ;
        RECT 62.325 58.020 67.140 58.160 ;
        RECT 62.325 57.975 62.615 58.020 ;
        RECT 64.240 57.880 64.380 58.020 ;
        RECT 67.000 57.880 67.140 58.020 ;
        RECT 72.430 57.960 72.750 58.220 ;
        RECT 74.360 58.205 74.500 58.360 ;
        RECT 74.820 58.205 74.960 58.700 ;
        RECT 77.030 58.640 77.350 58.700 ;
        RECT 77.530 58.840 77.820 58.885 ;
        RECT 79.630 58.840 79.920 58.885 ;
        RECT 81.200 58.840 81.490 58.885 ;
        RECT 77.530 58.700 81.490 58.840 ;
        RECT 77.530 58.655 77.820 58.700 ;
        RECT 79.630 58.655 79.920 58.700 ;
        RECT 81.200 58.655 81.490 58.700 ;
        RECT 77.925 58.500 78.215 58.545 ;
        RECT 79.115 58.500 79.405 58.545 ;
        RECT 81.635 58.500 81.925 58.545 ;
        RECT 75.280 58.360 77.720 58.500 ;
        RECT 75.280 58.205 75.420 58.360 ;
        RECT 74.285 57.975 74.575 58.205 ;
        RECT 74.745 57.975 75.035 58.205 ;
        RECT 75.205 57.975 75.495 58.205 ;
        RECT 76.125 58.160 76.415 58.205 ;
        RECT 76.570 58.160 76.890 58.220 ;
        RECT 76.125 58.020 76.890 58.160 ;
        RECT 76.125 57.975 76.415 58.020 ;
        RECT 76.570 57.960 76.890 58.020 ;
        RECT 77.045 57.975 77.335 58.205 ;
        RECT 77.580 58.160 77.720 58.360 ;
        RECT 77.925 58.360 81.925 58.500 ;
        RECT 77.925 58.315 78.215 58.360 ;
        RECT 79.115 58.315 79.405 58.360 ;
        RECT 81.635 58.315 81.925 58.360 ;
        RECT 84.405 58.160 84.695 58.205 ;
        RECT 77.580 58.020 84.695 58.160 ;
        RECT 84.405 57.975 84.695 58.020 ;
        RECT 86.705 58.160 86.995 58.205 ;
        RECT 87.150 58.160 87.470 58.220 ;
        RECT 86.705 58.020 87.470 58.160 ;
        RECT 86.705 57.975 86.995 58.020 ;
        RECT 63.690 57.865 64.010 57.880 ;
        RECT 63.660 57.635 64.010 57.865 ;
        RECT 63.690 57.620 64.010 57.635 ;
        RECT 64.150 57.620 64.470 57.880 ;
        RECT 66.910 57.820 67.230 57.880 ;
        RECT 71.970 57.820 72.290 57.880 ;
        RECT 77.120 57.820 77.260 57.975 ;
        RECT 87.150 57.960 87.470 58.020 ;
        RECT 78.270 57.820 78.560 57.865 ;
        RECT 85.325 57.820 85.615 57.865 ;
        RECT 66.910 57.680 77.260 57.820 ;
        RECT 77.580 57.680 78.560 57.820 ;
        RECT 66.910 57.620 67.230 57.680 ;
        RECT 71.970 57.620 72.290 57.680 ;
        RECT 48.065 57.340 50.120 57.480 ;
        RECT 50.350 57.480 50.670 57.540 ;
        RECT 55.885 57.480 56.175 57.525 ;
        RECT 50.350 57.340 56.175 57.480 ;
        RECT 48.065 57.295 48.355 57.340 ;
        RECT 50.350 57.280 50.670 57.340 ;
        RECT 55.885 57.295 56.175 57.340 ;
        RECT 68.750 57.480 69.070 57.540 ;
        RECT 69.225 57.480 69.515 57.525 ;
        RECT 68.750 57.340 69.515 57.480 ;
        RECT 68.750 57.280 69.070 57.340 ;
        RECT 69.225 57.295 69.515 57.340 ;
        RECT 72.905 57.480 73.195 57.525 ;
        RECT 77.580 57.480 77.720 57.680 ;
        RECT 78.270 57.635 78.560 57.680 ;
        RECT 84.020 57.680 85.615 57.820 ;
        RECT 72.905 57.340 77.720 57.480 ;
        RECT 80.710 57.480 81.030 57.540 ;
        RECT 84.020 57.525 84.160 57.680 ;
        RECT 85.325 57.635 85.615 57.680 ;
        RECT 86.245 57.635 86.535 57.865 ;
        RECT 83.945 57.480 84.235 57.525 ;
        RECT 80.710 57.340 84.235 57.480 ;
        RECT 72.905 57.295 73.195 57.340 ;
        RECT 80.710 57.280 81.030 57.340 ;
        RECT 83.945 57.295 84.235 57.340 ;
        RECT 84.390 57.480 84.710 57.540 ;
        RECT 86.320 57.480 86.460 57.635 ;
        RECT 87.150 57.480 87.470 57.540 ;
        RECT 84.390 57.340 87.470 57.480 ;
        RECT 84.390 57.280 84.710 57.340 ;
        RECT 87.150 57.280 87.470 57.340 ;
        RECT 12.100 56.660 89.840 57.140 ;
        RECT 21.845 56.460 22.135 56.505 ;
        RECT 23.210 56.460 23.530 56.520 ;
        RECT 21.845 56.320 23.530 56.460 ;
        RECT 21.845 56.275 22.135 56.320 ;
        RECT 23.210 56.260 23.530 56.320 ;
        RECT 25.065 56.460 25.355 56.505 ;
        RECT 27.365 56.460 27.655 56.505 ;
        RECT 25.065 56.320 27.655 56.460 ;
        RECT 25.065 56.275 25.355 56.320 ;
        RECT 27.365 56.275 27.655 56.320 ;
        RECT 28.745 56.460 29.035 56.505 ;
        RECT 30.110 56.460 30.430 56.520 ;
        RECT 28.745 56.320 30.430 56.460 ;
        RECT 28.745 56.275 29.035 56.320 ;
        RECT 30.110 56.260 30.430 56.320 ;
        RECT 38.390 56.260 38.710 56.520 ;
        RECT 41.150 56.260 41.470 56.520 ;
        RECT 49.430 56.460 49.750 56.520 ;
        RECT 51.730 56.460 52.050 56.520 ;
        RECT 49.430 56.320 52.050 56.460 ;
        RECT 49.430 56.260 49.750 56.320 ;
        RECT 51.730 56.260 52.050 56.320 ;
        RECT 71.050 56.260 71.370 56.520 ;
        RECT 79.330 56.460 79.650 56.520 ;
        RECT 75.280 56.320 79.650 56.460 ;
        RECT 25.970 56.120 26.290 56.180 ;
        RECT 26.905 56.120 27.195 56.165 ;
        RECT 21.000 55.980 27.195 56.120 ;
        RECT 21.000 55.825 21.140 55.980 ;
        RECT 25.970 55.920 26.290 55.980 ;
        RECT 26.905 55.935 27.195 55.980 ;
        RECT 27.950 56.120 28.240 56.165 ;
        RECT 29.650 56.120 29.970 56.180 ;
        RECT 27.950 55.980 29.970 56.120 ;
        RECT 27.950 55.935 28.240 55.980 ;
        RECT 29.650 55.920 29.970 55.980 ;
        RECT 36.090 56.120 36.410 56.180 ;
        RECT 39.165 56.120 39.455 56.165 ;
        RECT 36.090 55.980 39.455 56.120 ;
        RECT 36.090 55.920 36.410 55.980 ;
        RECT 39.165 55.935 39.455 55.980 ;
        RECT 40.245 55.935 40.535 56.165 ;
        RECT 68.750 56.120 69.070 56.180 ;
        RECT 75.280 56.120 75.420 56.320 ;
        RECT 79.330 56.260 79.650 56.320 ;
        RECT 80.340 56.320 81.400 56.460 ;
        RECT 48.140 55.980 55.640 56.120 ;
        RECT 20.465 55.595 20.755 55.825 ;
        RECT 20.925 55.595 21.215 55.825 ;
        RECT 20.540 55.440 20.680 55.595 ;
        RECT 23.210 55.580 23.530 55.840 ;
        RECT 26.430 55.780 26.750 55.840 ;
        RECT 30.585 55.780 30.875 55.825 ;
        RECT 23.760 55.640 26.200 55.780 ;
        RECT 21.370 55.440 21.690 55.500 ;
        RECT 23.760 55.485 23.900 55.640 ;
        RECT 20.540 55.300 21.690 55.440 ;
        RECT 21.370 55.240 21.690 55.300 ;
        RECT 21.845 55.255 22.135 55.485 ;
        RECT 23.685 55.255 23.975 55.485 ;
        RECT 24.590 55.440 24.910 55.500 ;
        RECT 25.525 55.440 25.815 55.485 ;
        RECT 24.590 55.300 25.815 55.440 ;
        RECT 26.060 55.440 26.200 55.640 ;
        RECT 26.430 55.640 30.875 55.780 ;
        RECT 26.430 55.580 26.750 55.640 ;
        RECT 30.585 55.595 30.875 55.640 ;
        RECT 36.565 55.780 36.855 55.825 ;
        RECT 37.930 55.780 38.250 55.840 ;
        RECT 40.320 55.780 40.460 55.935 ;
        RECT 48.140 55.825 48.280 55.980 ;
        RECT 36.565 55.640 38.250 55.780 ;
        RECT 36.565 55.595 36.855 55.640 ;
        RECT 37.930 55.580 38.250 55.640 ;
        RECT 38.940 55.640 40.460 55.780 ;
        RECT 46.785 55.780 47.075 55.825 ;
        RECT 46.785 55.640 47.820 55.780 ;
        RECT 38.940 55.500 39.080 55.640 ;
        RECT 46.785 55.595 47.075 55.640 ;
        RECT 33.790 55.440 34.110 55.500 ;
        RECT 34.265 55.440 34.555 55.485 ;
        RECT 26.060 55.300 34.555 55.440 ;
        RECT 21.920 54.760 22.060 55.255 ;
        RECT 24.590 55.240 24.910 55.300 ;
        RECT 25.525 55.255 25.815 55.300 ;
        RECT 33.790 55.240 34.110 55.300 ;
        RECT 34.265 55.255 34.555 55.300 ;
        RECT 38.850 55.240 39.170 55.500 ;
        RECT 43.475 55.440 43.765 55.485 ;
        RECT 45.995 55.440 46.285 55.485 ;
        RECT 47.185 55.440 47.475 55.485 ;
        RECT 43.475 55.300 47.475 55.440 ;
        RECT 47.680 55.440 47.820 55.640 ;
        RECT 48.065 55.595 48.355 55.825 ;
        RECT 49.890 55.780 50.210 55.840 ;
        RECT 55.500 55.825 55.640 55.980 ;
        RECT 68.750 55.980 75.420 56.120 ;
        RECT 75.650 56.120 75.970 56.180 ;
        RECT 77.490 56.120 77.810 56.180 ;
        RECT 80.340 56.120 80.480 56.320 ;
        RECT 75.650 55.980 80.480 56.120 ;
        RECT 68.750 55.920 69.070 55.980 ;
        RECT 75.650 55.920 75.970 55.980 ;
        RECT 77.490 55.920 77.810 55.980 ;
        RECT 80.710 55.920 81.030 56.180 ;
        RECT 81.260 56.120 81.400 56.320 ;
        RECT 83.485 56.120 83.775 56.165 ;
        RECT 81.260 55.980 81.430 56.120 ;
        RECT 53.125 55.780 53.415 55.825 ;
        RECT 49.890 55.640 53.415 55.780 ;
        RECT 49.890 55.580 50.210 55.640 ;
        RECT 53.125 55.595 53.415 55.640 ;
        RECT 55.425 55.780 55.715 55.825 ;
        RECT 55.870 55.780 56.190 55.840 ;
        RECT 55.425 55.640 56.190 55.780 ;
        RECT 55.425 55.595 55.715 55.640 ;
        RECT 55.870 55.580 56.190 55.640 ;
        RECT 56.760 55.780 57.050 55.825 ;
        RECT 58.630 55.780 58.950 55.840 ;
        RECT 56.760 55.640 58.950 55.780 ;
        RECT 56.760 55.595 57.050 55.640 ;
        RECT 58.630 55.580 58.950 55.640 ;
        RECT 64.150 55.580 64.470 55.840 ;
        RECT 65.500 55.780 65.790 55.825 ;
        RECT 69.670 55.780 69.990 55.840 ;
        RECT 65.500 55.640 69.990 55.780 ;
        RECT 65.500 55.595 65.790 55.640 ;
        RECT 69.670 55.580 69.990 55.640 ;
        RECT 71.970 55.580 72.290 55.840 ;
        RECT 73.350 55.825 73.670 55.840 ;
        RECT 73.320 55.595 73.670 55.825 ;
        RECT 73.350 55.580 73.670 55.595 ;
        RECT 80.250 55.580 80.570 55.840 ;
        RECT 81.290 55.825 81.430 55.980 ;
        RECT 81.720 55.980 83.775 56.120 ;
        RECT 81.720 55.840 81.860 55.980 ;
        RECT 83.485 55.935 83.775 55.980 ;
        RECT 84.850 56.120 85.170 56.180 ;
        RECT 85.325 56.120 85.615 56.165 ;
        RECT 84.850 55.980 85.615 56.120 ;
        RECT 84.850 55.920 85.170 55.980 ;
        RECT 85.325 55.935 85.615 55.980 ;
        RECT 85.785 56.120 86.075 56.165 ;
        RECT 87.150 56.120 87.470 56.180 ;
        RECT 85.785 55.980 87.470 56.120 ;
        RECT 85.785 55.935 86.075 55.980 ;
        RECT 87.150 55.920 87.470 55.980 ;
        RECT 81.185 55.595 81.475 55.825 ;
        RECT 81.630 55.580 81.950 55.840 ;
        RECT 82.105 55.595 82.395 55.825 ;
        RECT 84.405 55.595 84.695 55.825 ;
        RECT 47.680 55.300 48.280 55.440 ;
        RECT 43.475 55.255 43.765 55.300 ;
        RECT 45.995 55.255 46.285 55.300 ;
        RECT 47.185 55.255 47.475 55.300 ;
        RECT 35.185 55.100 35.475 55.145 ;
        RECT 40.230 55.100 40.550 55.160 ;
        RECT 35.185 54.960 40.550 55.100 ;
        RECT 35.185 54.915 35.475 54.960 ;
        RECT 40.230 54.900 40.550 54.960 ;
        RECT 43.910 55.100 44.200 55.145 ;
        RECT 45.480 55.100 45.770 55.145 ;
        RECT 47.580 55.100 47.870 55.145 ;
        RECT 43.910 54.960 47.870 55.100 ;
        RECT 48.140 55.100 48.280 55.300 ;
        RECT 48.510 55.240 48.830 55.500 ;
        RECT 54.490 55.240 54.810 55.500 ;
        RECT 56.305 55.440 56.595 55.485 ;
        RECT 57.495 55.440 57.785 55.485 ;
        RECT 60.015 55.440 60.305 55.485 ;
        RECT 56.305 55.300 60.305 55.440 ;
        RECT 56.305 55.255 56.595 55.300 ;
        RECT 57.495 55.255 57.785 55.300 ;
        RECT 60.015 55.255 60.305 55.300 ;
        RECT 65.045 55.440 65.335 55.485 ;
        RECT 66.235 55.440 66.525 55.485 ;
        RECT 68.755 55.440 69.045 55.485 ;
        RECT 65.045 55.300 69.045 55.440 ;
        RECT 65.045 55.255 65.335 55.300 ;
        RECT 66.235 55.255 66.525 55.300 ;
        RECT 68.755 55.255 69.045 55.300 ;
        RECT 72.865 55.440 73.155 55.485 ;
        RECT 74.055 55.440 74.345 55.485 ;
        RECT 76.575 55.440 76.865 55.485 ;
        RECT 82.180 55.440 82.320 55.595 ;
        RECT 72.865 55.300 76.865 55.440 ;
        RECT 72.865 55.255 73.155 55.300 ;
        RECT 74.055 55.255 74.345 55.300 ;
        RECT 76.575 55.255 76.865 55.300 ;
        RECT 78.960 55.300 82.320 55.440 ;
        RECT 84.480 55.440 84.620 55.595 ;
        RECT 86.690 55.580 87.010 55.840 ;
        RECT 86.230 55.440 86.550 55.500 ;
        RECT 84.480 55.300 86.550 55.440 ;
        RECT 52.205 55.100 52.495 55.145 ;
        RECT 48.140 54.960 52.495 55.100 ;
        RECT 43.910 54.915 44.200 54.960 ;
        RECT 45.480 54.915 45.770 54.960 ;
        RECT 47.580 54.915 47.870 54.960 ;
        RECT 52.205 54.915 52.495 54.960 ;
        RECT 55.910 55.100 56.200 55.145 ;
        RECT 58.010 55.100 58.300 55.145 ;
        RECT 59.580 55.100 59.870 55.145 ;
        RECT 55.910 54.960 59.870 55.100 ;
        RECT 55.910 54.915 56.200 54.960 ;
        RECT 58.010 54.915 58.300 54.960 ;
        RECT 59.580 54.915 59.870 54.960 ;
        RECT 64.650 55.100 64.940 55.145 ;
        RECT 66.750 55.100 67.040 55.145 ;
        RECT 68.320 55.100 68.610 55.145 ;
        RECT 64.650 54.960 68.610 55.100 ;
        RECT 64.650 54.915 64.940 54.960 ;
        RECT 66.750 54.915 67.040 54.960 ;
        RECT 68.320 54.915 68.610 54.960 ;
        RECT 72.470 55.100 72.760 55.145 ;
        RECT 74.570 55.100 74.860 55.145 ;
        RECT 76.140 55.100 76.430 55.145 ;
        RECT 72.470 54.960 76.430 55.100 ;
        RECT 72.470 54.915 72.760 54.960 ;
        RECT 74.570 54.915 74.860 54.960 ;
        RECT 76.140 54.915 76.430 54.960 ;
        RECT 78.960 54.820 79.100 55.300 ;
        RECT 86.230 55.240 86.550 55.300 ;
        RECT 79.330 54.900 79.650 55.160 ;
        RECT 26.890 54.760 27.210 54.820 ;
        RECT 21.920 54.620 27.210 54.760 ;
        RECT 26.890 54.560 27.210 54.620 ;
        RECT 39.310 54.560 39.630 54.820 ;
        RECT 52.650 54.760 52.970 54.820 ;
        RECT 54.045 54.760 54.335 54.805 ;
        RECT 52.650 54.620 54.335 54.760 ;
        RECT 52.650 54.560 52.970 54.620 ;
        RECT 54.045 54.575 54.335 54.620 ;
        RECT 60.470 54.760 60.790 54.820 ;
        RECT 62.325 54.760 62.615 54.805 ;
        RECT 67.830 54.760 68.150 54.820 ;
        RECT 72.890 54.760 73.210 54.820 ;
        RECT 60.470 54.620 73.210 54.760 ;
        RECT 60.470 54.560 60.790 54.620 ;
        RECT 62.325 54.575 62.615 54.620 ;
        RECT 67.830 54.560 68.150 54.620 ;
        RECT 72.890 54.560 73.210 54.620 ;
        RECT 78.870 54.560 79.190 54.820 ;
        RECT 79.790 54.760 80.110 54.820 ;
        RECT 87.625 54.760 87.915 54.805 ;
        RECT 79.790 54.620 87.915 54.760 ;
        RECT 79.790 54.560 80.110 54.620 ;
        RECT 87.625 54.575 87.915 54.620 ;
        RECT 12.100 53.940 89.840 54.420 ;
        RECT 15.850 53.740 16.170 53.800 ;
        RECT 16.325 53.740 16.615 53.785 ;
        RECT 15.850 53.600 16.615 53.740 ;
        RECT 15.850 53.540 16.170 53.600 ;
        RECT 16.325 53.555 16.615 53.600 ;
        RECT 24.590 53.540 24.910 53.800 ;
        RECT 26.445 53.555 26.735 53.785 ;
        RECT 26.890 53.740 27.210 53.800 ;
        RECT 29.205 53.740 29.495 53.785 ;
        RECT 26.890 53.600 29.495 53.740 ;
        RECT 14.470 53.400 14.790 53.460 ;
        RECT 19.085 53.400 19.375 53.445 ;
        RECT 14.470 53.260 19.375 53.400 ;
        RECT 14.470 53.200 14.790 53.260 ;
        RECT 19.085 53.215 19.375 53.260 ;
        RECT 18.150 53.060 18.470 53.120 ;
        RECT 17.780 52.920 18.470 53.060 ;
        RECT 17.780 52.765 17.920 52.920 ;
        RECT 18.150 52.860 18.470 52.920 ;
        RECT 17.705 52.535 17.995 52.765 ;
        RECT 22.290 52.720 22.610 52.780 ;
        RECT 18.240 52.580 22.610 52.720 ;
        RECT 14.010 52.380 14.330 52.440 ;
        RECT 16.165 52.380 16.455 52.425 ;
        RECT 14.010 52.240 16.455 52.380 ;
        RECT 14.010 52.180 14.330 52.240 ;
        RECT 16.165 52.195 16.455 52.240 ;
        RECT 16.770 52.380 17.090 52.440 ;
        RECT 17.245 52.380 17.535 52.425 ;
        RECT 16.770 52.240 17.535 52.380 ;
        RECT 16.770 52.180 17.090 52.240 ;
        RECT 17.245 52.195 17.535 52.240 ;
        RECT 18.240 52.100 18.380 52.580 ;
        RECT 22.290 52.520 22.610 52.580 ;
        RECT 22.765 52.720 23.055 52.765 ;
        RECT 24.130 52.720 24.450 52.780 ;
        RECT 22.765 52.580 24.450 52.720 ;
        RECT 24.680 52.720 24.820 53.540 ;
        RECT 26.520 53.400 26.660 53.555 ;
        RECT 26.890 53.540 27.210 53.600 ;
        RECT 29.205 53.555 29.495 53.600 ;
        RECT 30.570 53.740 30.890 53.800 ;
        RECT 31.505 53.740 31.795 53.785 ;
        RECT 30.570 53.600 31.795 53.740 ;
        RECT 30.570 53.540 30.890 53.600 ;
        RECT 31.505 53.555 31.795 53.600 ;
        RECT 48.065 53.740 48.355 53.785 ;
        RECT 48.510 53.740 48.830 53.800 ;
        RECT 48.065 53.600 48.830 53.740 ;
        RECT 48.065 53.555 48.355 53.600 ;
        RECT 48.510 53.540 48.830 53.600 ;
        RECT 49.430 53.540 49.750 53.800 ;
        RECT 63.690 53.540 64.010 53.800 ;
        RECT 73.810 53.540 74.130 53.800 ;
        RECT 87.610 53.540 87.930 53.800 ;
        RECT 37.930 53.400 38.250 53.460 ;
        RECT 26.520 53.260 38.250 53.400 ;
        RECT 37.930 53.200 38.250 53.260 ;
        RECT 41.650 53.400 41.940 53.445 ;
        RECT 43.750 53.400 44.040 53.445 ;
        RECT 45.320 53.400 45.610 53.445 ;
        RECT 41.650 53.260 45.610 53.400 ;
        RECT 41.650 53.215 41.940 53.260 ;
        RECT 43.750 53.215 44.040 53.260 ;
        RECT 45.320 53.215 45.610 53.260 ;
        RECT 50.365 53.215 50.655 53.445 ;
        RECT 51.770 53.400 52.060 53.445 ;
        RECT 53.870 53.400 54.160 53.445 ;
        RECT 55.440 53.400 55.730 53.445 ;
        RECT 51.770 53.260 55.730 53.400 ;
        RECT 51.770 53.215 52.060 53.260 ;
        RECT 53.870 53.215 54.160 53.260 ;
        RECT 55.440 53.215 55.730 53.260 ;
        RECT 67.830 53.400 68.150 53.460 ;
        RECT 78.870 53.400 79.190 53.460 ;
        RECT 67.830 53.260 79.190 53.400 ;
        RECT 25.050 53.060 25.370 53.120 ;
        RECT 25.050 52.920 26.200 53.060 ;
        RECT 25.050 52.860 25.370 52.920 ;
        RECT 25.525 52.720 25.815 52.765 ;
        RECT 24.680 52.580 25.815 52.720 ;
        RECT 26.060 52.720 26.200 52.920 ;
        RECT 26.430 52.860 26.750 53.120 ;
        RECT 42.045 53.060 42.335 53.105 ;
        RECT 43.235 53.060 43.525 53.105 ;
        RECT 45.755 53.060 46.045 53.105 ;
        RECT 27.440 52.920 30.800 53.060 ;
        RECT 26.905 52.720 27.195 52.765 ;
        RECT 26.060 52.580 27.195 52.720 ;
        RECT 22.765 52.535 23.055 52.580 ;
        RECT 24.130 52.520 24.450 52.580 ;
        RECT 25.525 52.535 25.815 52.580 ;
        RECT 26.905 52.535 27.195 52.580 ;
        RECT 19.085 52.380 19.375 52.425 ;
        RECT 21.370 52.380 21.690 52.440 ;
        RECT 23.670 52.380 23.990 52.440 ;
        RECT 19.085 52.240 20.450 52.380 ;
        RECT 19.085 52.195 19.375 52.240 ;
        RECT 15.390 51.840 15.710 52.100 ;
        RECT 18.150 51.840 18.470 52.100 ;
        RECT 20.310 52.040 20.450 52.240 ;
        RECT 21.370 52.240 23.990 52.380 ;
        RECT 21.370 52.180 21.690 52.240 ;
        RECT 23.670 52.180 23.990 52.240 ;
        RECT 20.910 52.040 21.230 52.100 ;
        RECT 23.210 52.040 23.530 52.100 ;
        RECT 27.440 52.040 27.580 52.920 ;
        RECT 30.660 52.765 30.800 52.920 ;
        RECT 42.045 52.920 46.045 53.060 ;
        RECT 42.045 52.875 42.335 52.920 ;
        RECT 43.235 52.875 43.525 52.920 ;
        RECT 45.755 52.875 46.045 52.920 ;
        RECT 48.050 53.060 48.370 53.120 ;
        RECT 50.440 53.060 50.580 53.215 ;
        RECT 67.830 53.200 68.150 53.260 ;
        RECT 48.050 52.920 50.580 53.060 ;
        RECT 48.050 52.860 48.370 52.920 ;
        RECT 30.125 52.720 30.415 52.765 ;
        RECT 27.900 52.580 30.415 52.720 ;
        RECT 27.900 52.085 28.040 52.580 ;
        RECT 30.125 52.535 30.415 52.580 ;
        RECT 30.585 52.535 30.875 52.765 ;
        RECT 31.965 52.720 32.255 52.765 ;
        RECT 32.870 52.720 33.190 52.780 ;
        RECT 31.965 52.580 33.190 52.720 ;
        RECT 31.965 52.535 32.255 52.580 ;
        RECT 32.870 52.520 33.190 52.580 ;
        RECT 33.805 52.535 34.095 52.765 ;
        RECT 34.250 52.720 34.570 52.780 ;
        RECT 40.705 52.720 40.995 52.765 ;
        RECT 34.250 52.580 40.995 52.720 ;
        RECT 33.880 52.380 34.020 52.535 ;
        RECT 34.250 52.520 34.570 52.580 ;
        RECT 40.705 52.535 40.995 52.580 ;
        RECT 41.165 52.535 41.455 52.765 ;
        RECT 42.500 52.720 42.790 52.765 ;
        RECT 44.830 52.720 45.150 52.780 ;
        RECT 42.500 52.580 45.150 52.720 ;
        RECT 42.500 52.535 42.790 52.580 ;
        RECT 37.025 52.380 37.315 52.425 ;
        RECT 38.390 52.380 38.710 52.440 ;
        RECT 39.770 52.380 40.090 52.440 ;
        RECT 41.240 52.380 41.380 52.535 ;
        RECT 44.830 52.520 45.150 52.580 ;
        RECT 33.880 52.240 41.380 52.380 ;
        RECT 37.025 52.195 37.315 52.240 ;
        RECT 38.390 52.180 38.710 52.240 ;
        RECT 39.770 52.180 40.090 52.240 ;
        RECT 48.510 52.180 48.830 52.440 ;
        RECT 50.440 52.380 50.580 52.920 ;
        RECT 52.165 53.060 52.455 53.105 ;
        RECT 53.355 53.060 53.645 53.105 ;
        RECT 55.875 53.060 56.165 53.105 ;
        RECT 52.165 52.920 56.165 53.060 ;
        RECT 52.165 52.875 52.455 52.920 ;
        RECT 53.355 52.875 53.645 52.920 ;
        RECT 55.875 52.875 56.165 52.920 ;
        RECT 66.450 52.860 66.770 53.120 ;
        RECT 67.370 53.060 67.690 53.120 ;
        RECT 67.370 52.920 74.040 53.060 ;
        RECT 67.370 52.860 67.690 52.920 ;
        RECT 51.285 52.720 51.575 52.765 ;
        RECT 63.245 52.720 63.535 52.765 ;
        RECT 65.070 52.720 65.390 52.780 ;
        RECT 73.900 52.765 74.040 52.920 ;
        RECT 73.365 52.720 73.655 52.765 ;
        RECT 51.285 52.580 56.100 52.720 ;
        RECT 51.285 52.535 51.575 52.580 ;
        RECT 55.960 52.440 56.100 52.580 ;
        RECT 63.245 52.580 73.655 52.720 ;
        RECT 63.245 52.535 63.535 52.580 ;
        RECT 65.070 52.520 65.390 52.580 ;
        RECT 73.365 52.535 73.655 52.580 ;
        RECT 73.825 52.535 74.115 52.765 ;
        RECT 74.270 52.520 74.590 52.780 ;
        RECT 75.650 52.520 75.970 52.780 ;
        RECT 78.040 52.765 78.180 53.260 ;
        RECT 78.870 53.200 79.190 53.260 ;
        RECT 77.965 52.535 78.255 52.765 ;
        RECT 81.170 52.720 81.490 52.780 ;
        RECT 82.105 52.720 82.395 52.765 ;
        RECT 81.170 52.580 82.395 52.720 ;
        RECT 81.170 52.520 81.490 52.580 ;
        RECT 82.105 52.535 82.395 52.580 ;
        RECT 82.550 52.520 82.870 52.780 ;
        RECT 83.025 52.535 83.315 52.765 ;
        RECT 83.470 52.720 83.790 52.780 ;
        RECT 83.945 52.720 84.235 52.765 ;
        RECT 83.470 52.580 84.235 52.720 ;
        RECT 52.510 52.380 52.800 52.425 ;
        RECT 50.440 52.240 52.800 52.380 ;
        RECT 52.510 52.195 52.800 52.240 ;
        RECT 55.870 52.380 56.190 52.440 ;
        RECT 59.105 52.380 59.395 52.425 ;
        RECT 55.870 52.240 59.395 52.380 ;
        RECT 55.870 52.180 56.190 52.240 ;
        RECT 59.105 52.195 59.395 52.240 ;
        RECT 65.545 52.380 65.835 52.425 ;
        RECT 68.750 52.380 69.070 52.440 ;
        RECT 65.545 52.240 69.070 52.380 ;
        RECT 65.545 52.195 65.835 52.240 ;
        RECT 68.750 52.180 69.070 52.240 ;
        RECT 69.210 52.180 69.530 52.440 ;
        RECT 75.740 52.380 75.880 52.520 ;
        RECT 78.885 52.380 79.175 52.425 ;
        RECT 81.630 52.380 81.950 52.440 ;
        RECT 75.740 52.240 81.950 52.380 ;
        RECT 83.100 52.380 83.240 52.535 ;
        RECT 83.470 52.520 83.790 52.580 ;
        RECT 83.945 52.535 84.235 52.580 ;
        RECT 85.310 52.520 85.630 52.780 ;
        RECT 85.770 52.720 86.090 52.780 ;
        RECT 86.705 52.720 86.995 52.765 ;
        RECT 85.770 52.580 86.995 52.720 ;
        RECT 85.770 52.520 86.090 52.580 ;
        RECT 86.705 52.535 86.995 52.580 ;
        RECT 84.405 52.380 84.695 52.425 ;
        RECT 83.100 52.240 84.695 52.380 ;
        RECT 78.885 52.195 79.175 52.240 ;
        RECT 81.630 52.180 81.950 52.240 ;
        RECT 84.405 52.195 84.695 52.240 ;
        RECT 86.230 52.380 86.550 52.440 ;
        RECT 87.150 52.380 87.470 52.440 ;
        RECT 86.230 52.240 87.470 52.380 ;
        RECT 86.230 52.180 86.550 52.240 ;
        RECT 87.150 52.180 87.470 52.240 ;
        RECT 20.310 51.900 27.580 52.040 ;
        RECT 20.910 51.840 21.230 51.900 ;
        RECT 23.210 51.840 23.530 51.900 ;
        RECT 27.825 51.855 28.115 52.085 ;
        RECT 48.050 52.040 48.370 52.100 ;
        RECT 49.525 52.040 49.815 52.085 ;
        RECT 51.730 52.040 52.050 52.100 ;
        RECT 48.050 51.900 52.050 52.040 ;
        RECT 48.050 51.840 48.370 51.900 ;
        RECT 49.525 51.855 49.815 51.900 ;
        RECT 51.730 51.840 52.050 51.900 ;
        RECT 58.185 52.040 58.475 52.085 ;
        RECT 62.310 52.040 62.630 52.100 ;
        RECT 58.185 51.900 62.630 52.040 ;
        RECT 58.185 51.855 58.475 51.900 ;
        RECT 62.310 51.840 62.630 51.900 ;
        RECT 65.990 51.840 66.310 52.100 ;
        RECT 68.290 52.040 68.610 52.100 ;
        RECT 75.665 52.040 75.955 52.085 ;
        RECT 68.290 51.900 75.955 52.040 ;
        RECT 68.290 51.840 68.610 51.900 ;
        RECT 75.665 51.855 75.955 51.900 ;
        RECT 76.110 52.040 76.430 52.100 ;
        RECT 77.045 52.040 77.335 52.085 ;
        RECT 76.110 51.900 77.335 52.040 ;
        RECT 76.110 51.840 76.430 51.900 ;
        RECT 77.045 51.855 77.335 51.900 ;
        RECT 80.710 51.840 81.030 52.100 ;
        RECT 12.100 51.220 89.840 51.700 ;
        RECT 13.565 51.020 13.855 51.065 ;
        RECT 18.150 51.020 18.470 51.080 ;
        RECT 13.565 50.880 18.470 51.020 ;
        RECT 13.565 50.835 13.855 50.880 ;
        RECT 18.150 50.820 18.470 50.880 ;
        RECT 25.970 51.020 26.290 51.080 ;
        RECT 28.285 51.020 28.575 51.065 ;
        RECT 25.970 50.880 28.575 51.020 ;
        RECT 25.970 50.820 26.290 50.880 ;
        RECT 28.285 50.835 28.575 50.880 ;
        RECT 30.110 51.020 30.430 51.080 ;
        RECT 31.585 51.020 31.875 51.065 ;
        RECT 30.110 50.880 31.875 51.020 ;
        RECT 30.110 50.820 30.430 50.880 ;
        RECT 31.585 50.835 31.875 50.880 ;
        RECT 32.885 51.020 33.175 51.065 ;
        RECT 33.330 51.020 33.650 51.080 ;
        RECT 32.885 50.880 33.650 51.020 ;
        RECT 32.885 50.835 33.175 50.880 ;
        RECT 33.330 50.820 33.650 50.880 ;
        RECT 48.065 51.020 48.355 51.065 ;
        RECT 48.970 51.020 49.290 51.080 ;
        RECT 48.065 50.880 49.290 51.020 ;
        RECT 48.065 50.835 48.355 50.880 ;
        RECT 48.970 50.820 49.290 50.880 ;
        RECT 55.410 50.820 55.730 51.080 ;
        RECT 58.630 50.820 58.950 51.080 ;
        RECT 60.470 50.820 60.790 51.080 ;
        RECT 69.225 51.020 69.515 51.065 ;
        RECT 69.670 51.020 69.990 51.080 ;
        RECT 69.225 50.880 69.990 51.020 ;
        RECT 69.225 50.835 69.515 50.880 ;
        RECT 69.670 50.820 69.990 50.880 ;
        RECT 71.050 51.020 71.370 51.080 ;
        RECT 71.525 51.020 71.815 51.065 ;
        RECT 71.050 50.880 71.815 51.020 ;
        RECT 71.050 50.820 71.370 50.880 ;
        RECT 71.525 50.835 71.815 50.880 ;
        RECT 18.610 50.680 18.930 50.740 ;
        RECT 18.610 50.540 20.220 50.680 ;
        RECT 18.610 50.480 18.930 50.540 ;
        RECT 19.070 50.385 19.390 50.400 ;
        RECT 19.070 50.155 19.420 50.385 ;
        RECT 19.070 50.140 19.390 50.155 ;
        RECT 15.875 50.000 16.165 50.045 ;
        RECT 18.395 50.000 18.685 50.045 ;
        RECT 19.585 50.000 19.875 50.045 ;
        RECT 15.875 49.860 19.875 50.000 ;
        RECT 20.080 50.000 20.220 50.540 ;
        RECT 20.910 50.480 21.230 50.740 ;
        RECT 21.925 50.680 22.215 50.725 ;
        RECT 21.460 50.540 22.215 50.680 ;
        RECT 20.450 50.140 20.770 50.400 ;
        RECT 21.460 50.000 21.600 50.540 ;
        RECT 21.925 50.495 22.215 50.540 ;
        RECT 26.430 50.680 26.750 50.740 ;
        RECT 29.205 50.680 29.495 50.725 ;
        RECT 26.430 50.540 29.495 50.680 ;
        RECT 26.430 50.480 26.750 50.540 ;
        RECT 29.205 50.495 29.495 50.540 ;
        RECT 30.585 50.680 30.875 50.725 ;
        RECT 34.250 50.680 34.570 50.740 ;
        RECT 38.405 50.680 38.695 50.725 ;
        RECT 30.585 50.540 34.570 50.680 ;
        RECT 30.585 50.495 30.875 50.540 ;
        RECT 34.250 50.480 34.570 50.540 ;
        RECT 34.800 50.540 38.695 50.680 ;
        RECT 23.225 50.340 23.515 50.385 ;
        RECT 20.080 49.860 21.600 50.000 ;
        RECT 22.840 50.200 23.515 50.340 ;
        RECT 15.875 49.815 16.165 49.860 ;
        RECT 18.395 49.815 18.685 49.860 ;
        RECT 19.585 49.815 19.875 49.860 ;
        RECT 16.310 49.660 16.600 49.705 ;
        RECT 17.880 49.660 18.170 49.705 ;
        RECT 19.980 49.660 20.270 49.705 ;
        RECT 16.310 49.520 20.270 49.660 ;
        RECT 16.310 49.475 16.600 49.520 ;
        RECT 17.880 49.475 18.170 49.520 ;
        RECT 19.980 49.475 20.270 49.520 ;
        RECT 21.370 49.660 21.690 49.720 ;
        RECT 22.840 49.705 22.980 50.200 ;
        RECT 23.225 50.155 23.515 50.200 ;
        RECT 24.130 50.140 24.450 50.400 ;
        RECT 30.125 50.155 30.415 50.385 ;
        RECT 30.200 50.000 30.340 50.155 ;
        RECT 33.790 50.140 34.110 50.400 ;
        RECT 34.800 50.385 34.940 50.540 ;
        RECT 38.405 50.495 38.695 50.540 ;
        RECT 42.500 50.680 42.790 50.725 ;
        RECT 47.130 50.680 47.450 50.740 ;
        RECT 67.385 50.680 67.675 50.725 ;
        RECT 70.590 50.680 70.910 50.740 ;
        RECT 42.500 50.540 47.450 50.680 ;
        RECT 42.500 50.495 42.790 50.540 ;
        RECT 47.130 50.480 47.450 50.540 ;
        RECT 48.600 50.540 56.100 50.680 ;
        RECT 34.725 50.155 35.015 50.385 ;
        RECT 35.170 50.140 35.490 50.400 ;
        RECT 37.930 50.340 38.250 50.400 ;
        RECT 48.600 50.385 48.740 50.540 ;
        RECT 55.960 50.400 56.100 50.540 ;
        RECT 67.385 50.540 70.910 50.680 ;
        RECT 67.385 50.495 67.675 50.540 ;
        RECT 70.590 50.480 70.910 50.540 ;
        RECT 39.325 50.340 39.615 50.385 ;
        RECT 37.930 50.200 39.615 50.340 ;
        RECT 37.930 50.140 38.250 50.200 ;
        RECT 39.325 50.155 39.615 50.200 ;
        RECT 48.525 50.155 48.815 50.385 ;
        RECT 48.970 50.340 49.290 50.400 ;
        RECT 49.805 50.340 50.095 50.385 ;
        RECT 48.970 50.200 50.095 50.340 ;
        RECT 48.970 50.140 49.290 50.200 ;
        RECT 49.805 50.155 50.095 50.200 ;
        RECT 55.870 50.140 56.190 50.400 ;
        RECT 60.945 50.340 61.235 50.385 ;
        RECT 65.990 50.340 66.310 50.400 ;
        RECT 66.925 50.340 67.215 50.385 ;
        RECT 71.065 50.340 71.355 50.385 ;
        RECT 60.945 50.200 71.355 50.340 ;
        RECT 71.600 50.340 71.740 50.835 ;
        RECT 73.350 50.820 73.670 51.080 ;
        RECT 75.190 51.020 75.510 51.080 ;
        RECT 85.310 51.020 85.630 51.080 ;
        RECT 88.085 51.020 88.375 51.065 ;
        RECT 75.190 50.880 80.480 51.020 ;
        RECT 75.190 50.820 75.510 50.880 ;
        RECT 79.790 50.680 80.110 50.740 ;
        RECT 78.500 50.540 80.110 50.680 ;
        RECT 74.745 50.340 75.035 50.385 ;
        RECT 71.600 50.200 75.035 50.340 ;
        RECT 60.945 50.155 61.235 50.200 ;
        RECT 30.570 50.000 30.890 50.060 ;
        RECT 36.090 50.000 36.410 50.060 ;
        RECT 30.200 49.860 30.890 50.000 ;
        RECT 30.570 49.800 30.890 49.860 ;
        RECT 32.500 49.860 36.410 50.000 ;
        RECT 22.765 49.660 23.055 49.705 ;
        RECT 21.370 49.520 23.055 49.660 ;
        RECT 21.370 49.460 21.690 49.520 ;
        RECT 22.765 49.475 23.055 49.520 ;
        RECT 23.225 49.660 23.515 49.705 ;
        RECT 26.890 49.660 27.210 49.720 ;
        RECT 32.500 49.705 32.640 49.860 ;
        RECT 36.090 49.800 36.410 49.860 ;
        RECT 40.230 49.800 40.550 50.060 ;
        RECT 41.165 49.815 41.455 50.045 ;
        RECT 42.045 50.000 42.335 50.045 ;
        RECT 43.235 50.000 43.525 50.045 ;
        RECT 45.755 50.000 46.045 50.045 ;
        RECT 42.045 49.860 46.045 50.000 ;
        RECT 42.045 49.815 42.335 49.860 ;
        RECT 43.235 49.815 43.525 49.860 ;
        RECT 45.755 49.815 46.045 49.860 ;
        RECT 49.405 50.000 49.695 50.045 ;
        RECT 50.595 50.000 50.885 50.045 ;
        RECT 53.115 50.000 53.405 50.045 ;
        RECT 49.405 49.860 53.405 50.000 ;
        RECT 49.405 49.815 49.695 49.860 ;
        RECT 50.595 49.815 50.885 49.860 ;
        RECT 53.115 49.815 53.405 49.860 ;
        RECT 54.490 50.000 54.810 50.060 ;
        RECT 61.020 50.000 61.160 50.155 ;
        RECT 65.990 50.140 66.310 50.200 ;
        RECT 66.925 50.155 67.215 50.200 ;
        RECT 71.065 50.155 71.355 50.200 ;
        RECT 74.745 50.155 75.035 50.200 ;
        RECT 75.190 50.140 75.510 50.400 ;
        RECT 75.665 50.340 75.955 50.385 ;
        RECT 76.110 50.340 76.430 50.400 ;
        RECT 75.665 50.200 76.430 50.340 ;
        RECT 75.665 50.155 75.955 50.200 ;
        RECT 76.110 50.140 76.430 50.200 ;
        RECT 76.570 50.340 76.890 50.400 ;
        RECT 78.500 50.385 78.640 50.540 ;
        RECT 79.790 50.480 80.110 50.540 ;
        RECT 77.505 50.340 77.795 50.385 ;
        RECT 76.570 50.200 77.795 50.340 ;
        RECT 76.570 50.140 76.890 50.200 ;
        RECT 77.505 50.155 77.795 50.200 ;
        RECT 78.425 50.155 78.715 50.385 ;
        RECT 78.885 50.155 79.175 50.385 ;
        RECT 79.345 50.340 79.635 50.385 ;
        RECT 80.340 50.340 80.480 50.880 ;
        RECT 85.310 50.880 88.375 51.020 ;
        RECT 85.310 50.820 85.630 50.880 ;
        RECT 88.085 50.835 88.375 50.880 ;
        RECT 80.710 50.680 81.030 50.740 ;
        RECT 82.410 50.680 82.700 50.725 ;
        RECT 80.710 50.540 82.700 50.680 ;
        RECT 80.710 50.480 81.030 50.540 ;
        RECT 82.410 50.495 82.700 50.540 ;
        RECT 85.310 50.340 85.630 50.400 ;
        RECT 79.345 50.200 85.630 50.340 ;
        RECT 79.345 50.155 79.635 50.200 ;
        RECT 54.490 49.860 61.160 50.000 ;
        RECT 23.225 49.520 27.210 49.660 ;
        RECT 23.225 49.475 23.515 49.520 ;
        RECT 26.890 49.460 27.210 49.520 ;
        RECT 32.425 49.475 32.715 49.705 ;
        RECT 34.250 49.460 34.570 49.720 ;
        RECT 38.390 49.660 38.710 49.720 ;
        RECT 41.240 49.660 41.380 49.815 ;
        RECT 54.490 49.800 54.810 49.860 ;
        RECT 61.390 49.800 61.710 50.060 ;
        RECT 68.290 49.800 68.610 50.060 ;
        RECT 71.970 49.800 72.290 50.060 ;
        RECT 73.350 50.000 73.670 50.060 ;
        RECT 75.280 50.000 75.420 50.140 ;
        RECT 78.960 50.000 79.100 50.155 ;
        RECT 73.350 49.860 75.420 50.000 ;
        RECT 78.500 49.860 79.100 50.000 ;
        RECT 73.350 49.800 73.670 49.860 ;
        RECT 78.500 49.720 78.640 49.860 ;
        RECT 38.390 49.520 41.380 49.660 ;
        RECT 41.650 49.660 41.940 49.705 ;
        RECT 43.750 49.660 44.040 49.705 ;
        RECT 45.320 49.660 45.610 49.705 ;
        RECT 41.650 49.520 45.610 49.660 ;
        RECT 38.390 49.460 38.710 49.520 ;
        RECT 41.650 49.475 41.940 49.520 ;
        RECT 43.750 49.475 44.040 49.520 ;
        RECT 45.320 49.475 45.610 49.520 ;
        RECT 49.010 49.660 49.300 49.705 ;
        RECT 51.110 49.660 51.400 49.705 ;
        RECT 52.680 49.660 52.970 49.705 ;
        RECT 49.010 49.520 52.970 49.660 ;
        RECT 49.010 49.475 49.300 49.520 ;
        RECT 51.110 49.475 51.400 49.520 ;
        RECT 52.680 49.475 52.970 49.520 ;
        RECT 78.410 49.460 78.730 49.720 ;
        RECT 21.845 49.320 22.135 49.365 ;
        RECT 22.290 49.320 22.610 49.380 ;
        RECT 21.845 49.180 22.610 49.320 ;
        RECT 21.845 49.135 22.135 49.180 ;
        RECT 22.290 49.120 22.610 49.180 ;
        RECT 29.650 49.320 29.970 49.380 ;
        RECT 31.505 49.320 31.795 49.365 ;
        RECT 33.330 49.320 33.650 49.380 ;
        RECT 29.650 49.180 33.650 49.320 ;
        RECT 29.650 49.120 29.970 49.180 ;
        RECT 31.505 49.135 31.795 49.180 ;
        RECT 33.330 49.120 33.650 49.180 ;
        RECT 55.410 49.320 55.730 49.380 ;
        RECT 60.010 49.320 60.330 49.380 ;
        RECT 62.770 49.320 63.090 49.380 ;
        RECT 55.410 49.180 63.090 49.320 ;
        RECT 55.410 49.120 55.730 49.180 ;
        RECT 60.010 49.120 60.330 49.180 ;
        RECT 62.770 49.120 63.090 49.180 ;
        RECT 65.085 49.320 65.375 49.365 ;
        RECT 65.530 49.320 65.850 49.380 ;
        RECT 65.085 49.180 65.850 49.320 ;
        RECT 65.085 49.135 65.375 49.180 ;
        RECT 65.530 49.120 65.850 49.180 ;
        RECT 71.510 49.320 71.830 49.380 ;
        RECT 79.420 49.320 79.560 50.155 ;
        RECT 85.310 50.140 85.630 50.200 ;
        RECT 81.170 49.800 81.490 50.060 ;
        RECT 82.065 50.000 82.355 50.045 ;
        RECT 83.255 50.000 83.545 50.045 ;
        RECT 85.775 50.000 86.065 50.045 ;
        RECT 82.065 49.860 86.065 50.000 ;
        RECT 82.065 49.815 82.355 49.860 ;
        RECT 83.255 49.815 83.545 49.860 ;
        RECT 85.775 49.815 86.065 49.860 ;
        RECT 80.725 49.660 81.015 49.705 ;
        RECT 81.670 49.660 81.960 49.705 ;
        RECT 83.770 49.660 84.060 49.705 ;
        RECT 85.340 49.660 85.630 49.705 ;
        RECT 80.725 49.520 81.400 49.660 ;
        RECT 80.725 49.475 81.015 49.520 ;
        RECT 71.510 49.180 79.560 49.320 ;
        RECT 81.260 49.320 81.400 49.520 ;
        RECT 81.670 49.520 85.630 49.660 ;
        RECT 81.670 49.475 81.960 49.520 ;
        RECT 83.770 49.475 84.060 49.520 ;
        RECT 85.340 49.475 85.630 49.520 ;
        RECT 82.550 49.320 82.870 49.380 ;
        RECT 81.260 49.180 82.870 49.320 ;
        RECT 71.510 49.120 71.830 49.180 ;
        RECT 82.550 49.120 82.870 49.180 ;
        RECT 12.100 48.500 89.840 48.980 ;
        RECT 20.450 48.300 20.770 48.360 ;
        RECT 14.560 48.160 20.770 48.300 ;
        RECT 14.560 47.665 14.700 48.160 ;
        RECT 20.450 48.100 20.770 48.160 ;
        RECT 20.910 48.300 21.230 48.360 ;
        RECT 21.385 48.300 21.675 48.345 ;
        RECT 33.345 48.300 33.635 48.345 ;
        RECT 38.865 48.300 39.155 48.345 ;
        RECT 20.910 48.160 24.820 48.300 ;
        RECT 20.910 48.100 21.230 48.160 ;
        RECT 21.385 48.115 21.675 48.160 ;
        RECT 14.970 47.960 15.260 48.005 ;
        RECT 17.070 47.960 17.360 48.005 ;
        RECT 18.640 47.960 18.930 48.005 ;
        RECT 14.970 47.820 18.930 47.960 ;
        RECT 14.970 47.775 15.260 47.820 ;
        RECT 17.070 47.775 17.360 47.820 ;
        RECT 18.640 47.775 18.930 47.820 ;
        RECT 19.530 47.960 19.850 48.020 ;
        RECT 24.680 48.005 24.820 48.160 ;
        RECT 33.345 48.160 39.155 48.300 ;
        RECT 33.345 48.115 33.635 48.160 ;
        RECT 38.865 48.115 39.155 48.160 ;
        RECT 47.145 48.300 47.435 48.345 ;
        RECT 48.510 48.300 48.830 48.360 ;
        RECT 47.145 48.160 48.830 48.300 ;
        RECT 47.145 48.115 47.435 48.160 ;
        RECT 48.510 48.100 48.830 48.160 ;
        RECT 51.270 48.100 51.590 48.360 ;
        RECT 53.125 48.115 53.415 48.345 ;
        RECT 54.045 48.300 54.335 48.345 ;
        RECT 61.850 48.300 62.170 48.360 ;
        RECT 54.045 48.160 62.170 48.300 ;
        RECT 54.045 48.115 54.335 48.160 ;
        RECT 21.845 47.960 22.135 48.005 ;
        RECT 19.530 47.820 22.135 47.960 ;
        RECT 19.530 47.760 19.850 47.820 ;
        RECT 21.845 47.775 22.135 47.820 ;
        RECT 24.605 47.775 24.895 48.005 ;
        RECT 26.905 47.960 27.195 48.005 ;
        RECT 33.790 47.960 34.110 48.020 ;
        RECT 26.905 47.820 34.110 47.960 ;
        RECT 26.905 47.775 27.195 47.820 ;
        RECT 14.485 47.435 14.775 47.665 ;
        RECT 15.365 47.620 15.655 47.665 ;
        RECT 16.555 47.620 16.845 47.665 ;
        RECT 19.075 47.620 19.365 47.665 ;
        RECT 15.365 47.480 19.365 47.620 ;
        RECT 21.920 47.620 22.060 47.775 ;
        RECT 33.790 47.760 34.110 47.820 ;
        RECT 34.710 47.960 35.030 48.020 ;
        RECT 35.185 47.960 35.475 48.005 ;
        RECT 35.645 47.960 35.935 48.005 ;
        RECT 34.710 47.820 35.935 47.960 ;
        RECT 34.710 47.760 35.030 47.820 ;
        RECT 35.185 47.775 35.475 47.820 ;
        RECT 35.645 47.775 35.935 47.820 ;
        RECT 37.930 47.960 38.250 48.020 ;
        RECT 53.200 47.960 53.340 48.115 ;
        RECT 61.850 48.100 62.170 48.160 ;
        RECT 63.245 48.300 63.535 48.345 ;
        RECT 65.070 48.300 65.390 48.360 ;
        RECT 67.370 48.300 67.690 48.360 ;
        RECT 63.245 48.160 67.690 48.300 ;
        RECT 63.245 48.115 63.535 48.160 ;
        RECT 65.070 48.100 65.390 48.160 ;
        RECT 67.370 48.100 67.690 48.160 ;
        RECT 70.130 48.300 70.450 48.360 ;
        RECT 72.905 48.300 73.195 48.345 ;
        RECT 73.810 48.300 74.130 48.360 ;
        RECT 70.130 48.160 74.130 48.300 ;
        RECT 70.130 48.100 70.450 48.160 ;
        RECT 72.905 48.115 73.195 48.160 ;
        RECT 73.810 48.100 74.130 48.160 ;
        RECT 86.690 48.300 87.010 48.360 ;
        RECT 88.085 48.300 88.375 48.345 ;
        RECT 86.690 48.160 88.375 48.300 ;
        RECT 86.690 48.100 87.010 48.160 ;
        RECT 88.085 48.115 88.375 48.160 ;
        RECT 55.410 47.960 55.730 48.020 ;
        RECT 37.930 47.820 44.140 47.960 ;
        RECT 53.200 47.820 55.730 47.960 ;
        RECT 37.930 47.760 38.250 47.820 ;
        RECT 41.165 47.620 41.455 47.665 ;
        RECT 21.920 47.480 28.500 47.620 ;
        RECT 15.365 47.435 15.655 47.480 ;
        RECT 16.555 47.435 16.845 47.480 ;
        RECT 19.075 47.435 19.365 47.480 ;
        RECT 14.560 47.280 14.700 47.435 ;
        RECT 14.930 47.280 15.250 47.340 ;
        RECT 15.850 47.325 16.170 47.340 ;
        RECT 15.820 47.280 16.170 47.325 ;
        RECT 14.560 47.140 15.250 47.280 ;
        RECT 15.655 47.140 16.170 47.280 ;
        RECT 14.930 47.080 15.250 47.140 ;
        RECT 15.820 47.095 16.170 47.140 ;
        RECT 15.850 47.080 16.170 47.095 ;
        RECT 21.830 47.280 22.150 47.340 ;
        RECT 23.685 47.280 23.975 47.325 ;
        RECT 24.130 47.280 24.450 47.340 ;
        RECT 25.600 47.325 25.740 47.480 ;
        RECT 21.830 47.140 24.450 47.280 ;
        RECT 21.830 47.080 22.150 47.140 ;
        RECT 23.685 47.095 23.975 47.140 ;
        RECT 24.130 47.080 24.450 47.140 ;
        RECT 25.525 47.095 25.815 47.325 ;
        RECT 25.985 47.280 26.275 47.325 ;
        RECT 26.430 47.280 26.750 47.340 ;
        RECT 25.985 47.140 26.750 47.280 ;
        RECT 25.985 47.095 26.275 47.140 ;
        RECT 26.430 47.080 26.750 47.140 ;
        RECT 27.350 47.080 27.670 47.340 ;
        RECT 28.360 47.325 28.500 47.480 ;
        RECT 37.560 47.480 41.455 47.620 ;
        RECT 28.285 47.095 28.575 47.325 ;
        RECT 35.170 47.280 35.490 47.340 ;
        RECT 37.010 47.280 37.330 47.340 ;
        RECT 37.560 47.325 37.700 47.480 ;
        RECT 41.165 47.435 41.455 47.480 ;
        RECT 37.485 47.280 37.775 47.325 ;
        RECT 35.170 47.140 37.775 47.280 ;
        RECT 35.170 47.080 35.490 47.140 ;
        RECT 37.010 47.080 37.330 47.140 ;
        RECT 37.485 47.095 37.775 47.140 ;
        RECT 37.930 47.280 38.250 47.340 ;
        RECT 39.785 47.280 40.075 47.325 ;
        RECT 37.930 47.140 40.075 47.280 ;
        RECT 37.930 47.080 38.250 47.140 ;
        RECT 39.785 47.095 40.075 47.140 ;
        RECT 40.230 47.080 40.550 47.340 ;
        RECT 44.000 47.325 44.140 47.820 ;
        RECT 55.410 47.760 55.730 47.820 ;
        RECT 56.790 47.960 57.080 48.005 ;
        RECT 58.360 47.960 58.650 48.005 ;
        RECT 60.460 47.960 60.750 48.005 ;
        RECT 56.790 47.820 60.750 47.960 ;
        RECT 56.790 47.775 57.080 47.820 ;
        RECT 58.360 47.775 58.650 47.820 ;
        RECT 60.460 47.775 60.750 47.820 ;
        RECT 64.650 47.960 64.940 48.005 ;
        RECT 66.750 47.960 67.040 48.005 ;
        RECT 68.320 47.960 68.610 48.005 ;
        RECT 64.650 47.820 68.610 47.960 ;
        RECT 64.650 47.775 64.940 47.820 ;
        RECT 66.750 47.775 67.040 47.820 ;
        RECT 68.320 47.775 68.610 47.820 ;
        RECT 70.590 47.960 70.910 48.020 ;
        RECT 71.065 47.960 71.355 48.005 ;
        RECT 80.710 47.960 81.030 48.020 ;
        RECT 70.590 47.820 81.030 47.960 ;
        RECT 70.590 47.760 70.910 47.820 ;
        RECT 71.065 47.775 71.355 47.820 ;
        RECT 80.710 47.760 81.030 47.820 ;
        RECT 81.670 47.960 81.960 48.005 ;
        RECT 83.770 47.960 84.060 48.005 ;
        RECT 85.340 47.960 85.630 48.005 ;
        RECT 81.670 47.820 85.630 47.960 ;
        RECT 81.670 47.775 81.960 47.820 ;
        RECT 83.770 47.775 84.060 47.820 ;
        RECT 85.340 47.775 85.630 47.820 ;
        RECT 49.430 47.620 49.750 47.680 ;
        RECT 49.905 47.620 50.195 47.665 ;
        RECT 52.665 47.620 52.955 47.665 ;
        RECT 49.430 47.480 52.955 47.620 ;
        RECT 49.430 47.420 49.750 47.480 ;
        RECT 49.905 47.435 50.195 47.480 ;
        RECT 52.665 47.435 52.955 47.480 ;
        RECT 56.355 47.620 56.645 47.665 ;
        RECT 58.875 47.620 59.165 47.665 ;
        RECT 60.065 47.620 60.355 47.665 ;
        RECT 64.165 47.620 64.455 47.665 ;
        RECT 56.355 47.480 60.355 47.620 ;
        RECT 56.355 47.435 56.645 47.480 ;
        RECT 58.875 47.435 59.165 47.480 ;
        RECT 60.065 47.435 60.355 47.480 ;
        RECT 61.020 47.480 64.455 47.620 ;
        RECT 40.705 47.095 40.995 47.325 ;
        RECT 43.925 47.095 44.215 47.325 ;
        RECT 45.765 47.095 46.055 47.325 ;
        RECT 46.685 47.280 46.975 47.325 ;
        RECT 53.125 47.280 53.415 47.325 ;
        RECT 46.685 47.140 53.415 47.280 ;
        RECT 46.685 47.095 46.975 47.140 ;
        RECT 53.125 47.095 53.415 47.140 ;
        RECT 55.870 47.280 56.190 47.340 ;
        RECT 61.020 47.325 61.160 47.480 ;
        RECT 64.165 47.435 64.455 47.480 ;
        RECT 65.045 47.620 65.335 47.665 ;
        RECT 66.235 47.620 66.525 47.665 ;
        RECT 68.755 47.620 69.045 47.665 ;
        RECT 65.045 47.480 69.045 47.620 ;
        RECT 65.045 47.435 65.335 47.480 ;
        RECT 66.235 47.435 66.525 47.480 ;
        RECT 68.755 47.435 69.045 47.480 ;
        RECT 69.210 47.620 69.530 47.680 ;
        RECT 81.170 47.620 81.490 47.680 ;
        RECT 69.210 47.480 81.490 47.620 ;
        RECT 69.210 47.420 69.530 47.480 ;
        RECT 81.170 47.420 81.490 47.480 ;
        RECT 82.065 47.620 82.355 47.665 ;
        RECT 83.255 47.620 83.545 47.665 ;
        RECT 85.775 47.620 86.065 47.665 ;
        RECT 82.065 47.480 86.065 47.620 ;
        RECT 82.065 47.435 82.355 47.480 ;
        RECT 83.255 47.435 83.545 47.480 ;
        RECT 85.775 47.435 86.065 47.480 ;
        RECT 60.945 47.280 61.235 47.325 ;
        RECT 55.870 47.140 61.235 47.280 ;
        RECT 18.610 46.940 18.930 47.000 ;
        RECT 22.765 46.940 23.055 46.985 ;
        RECT 26.905 46.940 27.195 46.985 ;
        RECT 18.610 46.800 23.055 46.940 ;
        RECT 18.610 46.740 18.930 46.800 ;
        RECT 22.765 46.755 23.055 46.800 ;
        RECT 23.760 46.800 27.195 46.940 ;
        RECT 23.760 46.660 23.900 46.800 ;
        RECT 26.905 46.755 27.195 46.800 ;
        RECT 30.570 46.940 30.890 47.000 ;
        RECT 38.405 46.940 38.695 46.985 ;
        RECT 40.780 46.940 40.920 47.095 ;
        RECT 41.150 46.940 41.470 47.000 ;
        RECT 43.005 46.940 43.295 46.985 ;
        RECT 30.570 46.800 43.295 46.940 ;
        RECT 45.840 46.940 45.980 47.095 ;
        RECT 52.190 46.940 52.510 47.000 ;
        RECT 45.840 46.800 52.510 46.940 ;
        RECT 53.200 46.940 53.340 47.095 ;
        RECT 55.870 47.080 56.190 47.140 ;
        RECT 60.945 47.095 61.235 47.140 ;
        RECT 61.405 47.095 61.695 47.325 ;
        RECT 62.325 47.280 62.615 47.325 ;
        RECT 62.770 47.280 63.090 47.340 ;
        RECT 65.530 47.325 65.850 47.340 ;
        RECT 65.500 47.280 65.850 47.325 ;
        RECT 62.325 47.140 63.090 47.280 ;
        RECT 65.335 47.140 65.850 47.280 ;
        RECT 62.325 47.095 62.615 47.140 ;
        RECT 58.630 46.940 58.950 47.000 ;
        RECT 53.200 46.800 58.950 46.940 ;
        RECT 30.570 46.740 30.890 46.800 ;
        RECT 38.405 46.755 38.695 46.800 ;
        RECT 41.150 46.740 41.470 46.800 ;
        RECT 43.005 46.755 43.295 46.800 ;
        RECT 52.190 46.740 52.510 46.800 ;
        RECT 58.630 46.740 58.950 46.800 ;
        RECT 59.550 46.985 59.870 47.000 ;
        RECT 59.550 46.940 59.900 46.985 ;
        RECT 59.550 46.800 60.065 46.940 ;
        RECT 59.550 46.755 59.900 46.800 ;
        RECT 59.550 46.740 59.870 46.755 ;
        RECT 20.910 46.600 21.230 46.660 ;
        RECT 22.290 46.600 22.610 46.660 ;
        RECT 23.225 46.600 23.515 46.645 ;
        RECT 20.910 46.460 23.515 46.600 ;
        RECT 20.910 46.400 21.230 46.460 ;
        RECT 22.290 46.400 22.610 46.460 ;
        RECT 23.225 46.415 23.515 46.460 ;
        RECT 23.670 46.400 23.990 46.660 ;
        RECT 27.810 46.400 28.130 46.660 ;
        RECT 32.425 46.600 32.715 46.645 ;
        RECT 32.870 46.600 33.190 46.660 ;
        RECT 32.425 46.460 33.190 46.600 ;
        RECT 32.425 46.415 32.715 46.460 ;
        RECT 32.870 46.400 33.190 46.460 ;
        RECT 33.330 46.600 33.650 46.660 ;
        RECT 35.170 46.600 35.490 46.660 ;
        RECT 33.330 46.460 35.490 46.600 ;
        RECT 33.330 46.400 33.650 46.460 ;
        RECT 35.170 46.400 35.490 46.460 ;
        RECT 36.550 46.400 36.870 46.660 ;
        RECT 37.010 46.600 37.330 46.660 ;
        RECT 40.230 46.600 40.550 46.660 ;
        RECT 37.010 46.460 40.550 46.600 ;
        RECT 37.010 46.400 37.330 46.460 ;
        RECT 40.230 46.400 40.550 46.460 ;
        RECT 42.070 46.400 42.390 46.660 ;
        RECT 46.685 46.600 46.975 46.645 ;
        RECT 56.330 46.600 56.650 46.660 ;
        RECT 61.480 46.600 61.620 47.095 ;
        RECT 62.770 47.080 63.090 47.140 ;
        RECT 65.500 47.095 65.850 47.140 ;
        RECT 65.530 47.080 65.850 47.095 ;
        RECT 71.050 47.280 71.370 47.340 ;
        RECT 72.905 47.280 73.195 47.325 ;
        RECT 74.270 47.280 74.590 47.340 ;
        RECT 71.050 47.140 74.590 47.280 ;
        RECT 71.050 47.080 71.370 47.140 ;
        RECT 72.905 47.095 73.195 47.140 ;
        RECT 74.270 47.080 74.590 47.140 ;
        RECT 74.730 47.080 75.050 47.340 ;
        RECT 75.190 47.280 75.510 47.340 ;
        RECT 76.570 47.280 76.890 47.340 ;
        RECT 77.045 47.280 77.335 47.325 ;
        RECT 75.190 47.140 77.335 47.280 ;
        RECT 75.190 47.080 75.510 47.140 ;
        RECT 76.570 47.080 76.890 47.140 ;
        RECT 77.045 47.095 77.335 47.140 ;
        RECT 77.950 47.080 78.270 47.340 ;
        RECT 78.410 47.080 78.730 47.340 ;
        RECT 78.870 47.080 79.190 47.340 ;
        RECT 82.550 47.325 82.870 47.340 ;
        RECT 82.520 47.280 82.870 47.325 ;
        RECT 82.355 47.140 82.870 47.280 ;
        RECT 82.520 47.095 82.870 47.140 ;
        RECT 82.550 47.080 82.870 47.095 ;
        RECT 67.370 46.940 67.690 47.000 ;
        RECT 78.500 46.940 78.640 47.080 ;
        RECT 82.090 46.940 82.410 47.000 ;
        RECT 67.370 46.800 72.200 46.940 ;
        RECT 78.500 46.800 82.410 46.940 ;
        RECT 67.370 46.740 67.690 46.800 ;
        RECT 72.060 46.645 72.200 46.800 ;
        RECT 82.090 46.740 82.410 46.800 ;
        RECT 46.685 46.460 61.620 46.600 ;
        RECT 46.685 46.415 46.975 46.460 ;
        RECT 56.330 46.400 56.650 46.460 ;
        RECT 71.985 46.415 72.275 46.645 ;
        RECT 80.250 46.400 80.570 46.660 ;
        RECT 80.710 46.600 81.030 46.660 ;
        RECT 81.630 46.600 81.950 46.660 ;
        RECT 88.070 46.600 88.390 46.660 ;
        RECT 80.710 46.460 88.390 46.600 ;
        RECT 80.710 46.400 81.030 46.460 ;
        RECT 81.630 46.400 81.950 46.460 ;
        RECT 88.070 46.400 88.390 46.460 ;
        RECT 12.100 45.780 89.840 46.260 ;
        RECT 21.370 45.580 21.690 45.640 ;
        RECT 13.640 45.440 21.690 45.580 ;
        RECT 13.640 44.945 13.780 45.440 ;
        RECT 21.370 45.380 21.690 45.440 ;
        RECT 21.830 45.380 22.150 45.640 ;
        RECT 22.305 45.395 22.595 45.625 ;
        RECT 23.145 45.580 23.435 45.625 ;
        RECT 27.810 45.580 28.130 45.640 ;
        RECT 23.145 45.440 28.130 45.580 ;
        RECT 23.145 45.395 23.435 45.440 ;
        RECT 14.010 45.040 14.330 45.300 ;
        RECT 16.280 45.240 16.570 45.285 ;
        RECT 22.380 45.240 22.520 45.395 ;
        RECT 27.810 45.380 28.130 45.440 ;
        RECT 30.110 45.380 30.430 45.640 ;
        RECT 37.010 45.580 37.330 45.640 ;
        RECT 31.120 45.440 37.330 45.580 ;
        RECT 16.280 45.100 22.520 45.240 ;
        RECT 16.280 45.055 16.570 45.100 ;
        RECT 24.145 45.055 24.435 45.285 ;
        RECT 29.665 45.240 29.955 45.285 ;
        RECT 31.120 45.240 31.260 45.440 ;
        RECT 37.010 45.380 37.330 45.440 ;
        RECT 37.470 45.380 37.790 45.640 ;
        RECT 47.145 45.580 47.435 45.625 ;
        RECT 48.970 45.580 49.290 45.640 ;
        RECT 54.490 45.580 54.810 45.640 ;
        RECT 47.145 45.440 49.290 45.580 ;
        RECT 47.145 45.395 47.435 45.440 ;
        RECT 48.970 45.380 49.290 45.440 ;
        RECT 49.520 45.440 54.810 45.580 ;
        RECT 49.520 45.240 49.660 45.440 ;
        RECT 54.490 45.380 54.810 45.440 ;
        RECT 63.230 45.580 63.550 45.640 ;
        RECT 74.730 45.580 75.050 45.640 ;
        RECT 63.230 45.440 75.050 45.580 ;
        RECT 63.230 45.380 63.550 45.440 ;
        RECT 74.730 45.380 75.050 45.440 ;
        RECT 87.610 45.380 87.930 45.640 ;
        RECT 55.870 45.240 56.190 45.300 ;
        RECT 69.210 45.240 69.530 45.300 ;
        RECT 81.170 45.240 81.490 45.300 ;
        RECT 29.665 45.100 31.260 45.240 ;
        RECT 31.580 45.100 34.940 45.240 ;
        RECT 29.665 45.055 29.955 45.100 ;
        RECT 13.565 44.715 13.855 44.945 ;
        RECT 14.470 44.700 14.790 44.960 ;
        RECT 14.930 44.700 15.250 44.960 ;
        RECT 17.690 44.900 18.010 44.960 ;
        RECT 24.220 44.900 24.360 45.055 ;
        RECT 25.065 44.900 25.355 44.945 ;
        RECT 17.690 44.760 25.355 44.900 ;
        RECT 17.690 44.700 18.010 44.760 ;
        RECT 25.065 44.715 25.355 44.760 ;
        RECT 25.985 44.715 26.275 44.945 ;
        RECT 15.825 44.560 16.115 44.605 ;
        RECT 17.015 44.560 17.305 44.605 ;
        RECT 19.535 44.560 19.825 44.605 ;
        RECT 26.060 44.560 26.200 44.715 ;
        RECT 26.430 44.700 26.750 44.960 ;
        RECT 26.890 44.700 27.210 44.960 ;
        RECT 28.745 44.715 29.035 44.945 ;
        RECT 15.825 44.420 19.825 44.560 ;
        RECT 15.825 44.375 16.115 44.420 ;
        RECT 17.015 44.375 17.305 44.420 ;
        RECT 19.535 44.375 19.825 44.420 ;
        RECT 23.300 44.420 26.200 44.560 ;
        RECT 28.820 44.560 28.960 44.715 ;
        RECT 30.110 44.700 30.430 44.960 ;
        RECT 30.585 44.900 30.875 44.945 ;
        RECT 31.580 44.900 31.720 45.100 ;
        RECT 34.800 44.960 34.940 45.100 ;
        RECT 45.840 45.100 49.660 45.240 ;
        RECT 51.820 45.100 56.190 45.240 ;
        RECT 30.585 44.760 31.720 44.900 ;
        RECT 31.920 44.900 32.210 44.945 ;
        RECT 33.330 44.900 33.650 44.960 ;
        RECT 31.920 44.760 33.650 44.900 ;
        RECT 30.585 44.715 30.875 44.760 ;
        RECT 31.920 44.715 32.210 44.760 ;
        RECT 33.330 44.700 33.650 44.760 ;
        RECT 34.710 44.900 35.030 44.960 ;
        RECT 38.390 44.900 38.710 44.960 ;
        RECT 34.710 44.760 38.710 44.900 ;
        RECT 34.710 44.700 35.030 44.760 ;
        RECT 38.390 44.700 38.710 44.760 ;
        RECT 39.740 44.900 40.030 44.945 ;
        RECT 41.610 44.900 41.930 44.960 ;
        RECT 45.840 44.945 45.980 45.100 ;
        RECT 39.740 44.760 41.930 44.900 ;
        RECT 39.740 44.715 40.030 44.760 ;
        RECT 41.610 44.700 41.930 44.760 ;
        RECT 45.765 44.715 46.055 44.945 ;
        RECT 46.225 44.900 46.515 44.945 ;
        RECT 48.050 44.900 48.370 44.960 ;
        RECT 46.225 44.760 48.370 44.900 ;
        RECT 46.225 44.715 46.515 44.760 ;
        RECT 48.050 44.700 48.370 44.760 ;
        RECT 48.525 44.900 48.815 44.945 ;
        RECT 50.350 44.900 50.670 44.960 ;
        RECT 51.820 44.945 51.960 45.100 ;
        RECT 55.870 45.040 56.190 45.100 ;
        RECT 64.240 45.100 72.200 45.240 ;
        RECT 48.525 44.760 50.670 44.900 ;
        RECT 48.525 44.715 48.815 44.760 ;
        RECT 50.350 44.700 50.670 44.760 ;
        RECT 51.745 44.715 52.035 44.945 ;
        RECT 53.025 44.900 53.315 44.945 ;
        RECT 52.280 44.760 53.315 44.900 ;
        RECT 31.465 44.560 31.755 44.605 ;
        RECT 32.655 44.560 32.945 44.605 ;
        RECT 35.175 44.560 35.465 44.605 ;
        RECT 28.820 44.420 30.800 44.560 ;
        RECT 15.430 44.220 15.720 44.265 ;
        RECT 17.530 44.220 17.820 44.265 ;
        RECT 19.100 44.220 19.390 44.265 ;
        RECT 15.430 44.080 19.390 44.220 ;
        RECT 15.430 44.035 15.720 44.080 ;
        RECT 17.530 44.035 17.820 44.080 ;
        RECT 19.100 44.035 19.390 44.080 ;
        RECT 16.310 43.880 16.630 43.940 ;
        RECT 18.150 43.880 18.470 43.940 ;
        RECT 23.300 43.925 23.440 44.420 ;
        RECT 28.285 44.220 28.575 44.265 ;
        RECT 29.650 44.220 29.970 44.280 ;
        RECT 28.285 44.080 29.970 44.220 ;
        RECT 28.285 44.035 28.575 44.080 ;
        RECT 29.650 44.020 29.970 44.080 ;
        RECT 23.225 43.880 23.515 43.925 ;
        RECT 16.310 43.740 23.515 43.880 ;
        RECT 30.660 43.880 30.800 44.420 ;
        RECT 31.465 44.420 35.465 44.560 ;
        RECT 31.465 44.375 31.755 44.420 ;
        RECT 32.655 44.375 32.945 44.420 ;
        RECT 35.175 44.375 35.465 44.420 ;
        RECT 39.285 44.560 39.575 44.605 ;
        RECT 40.475 44.560 40.765 44.605 ;
        RECT 42.995 44.560 43.285 44.605 ;
        RECT 39.285 44.420 43.285 44.560 ;
        RECT 39.285 44.375 39.575 44.420 ;
        RECT 40.475 44.375 40.765 44.420 ;
        RECT 42.995 44.375 43.285 44.420 ;
        RECT 47.145 44.560 47.435 44.605 ;
        RECT 47.590 44.560 47.910 44.620 ;
        RECT 47.145 44.420 47.910 44.560 ;
        RECT 47.145 44.375 47.435 44.420 ;
        RECT 47.590 44.360 47.910 44.420 ;
        RECT 48.985 44.560 49.275 44.605 ;
        RECT 49.890 44.560 50.210 44.620 ;
        RECT 52.280 44.560 52.420 44.760 ;
        RECT 53.025 44.715 53.315 44.760 ;
        RECT 54.950 44.900 55.270 44.960 ;
        RECT 59.105 44.900 59.395 44.945 ;
        RECT 54.950 44.760 59.395 44.900 ;
        RECT 54.950 44.700 55.270 44.760 ;
        RECT 59.105 44.715 59.395 44.760 ;
        RECT 62.310 44.700 62.630 44.960 ;
        RECT 64.240 44.945 64.380 45.100 ;
        RECT 69.210 45.040 69.530 45.100 ;
        RECT 64.165 44.715 64.455 44.945 ;
        RECT 64.610 44.900 64.930 44.960 ;
        RECT 72.060 44.945 72.200 45.100 ;
        RECT 81.170 45.100 86.460 45.240 ;
        RECT 81.170 45.040 81.490 45.100 ;
        RECT 65.445 44.900 65.735 44.945 ;
        RECT 64.610 44.760 65.735 44.900 ;
        RECT 64.610 44.700 64.930 44.760 ;
        RECT 65.445 44.715 65.735 44.760 ;
        RECT 71.985 44.715 72.275 44.945 ;
        RECT 72.430 44.900 72.750 44.960 ;
        RECT 73.265 44.900 73.555 44.945 ;
        RECT 72.430 44.760 73.555 44.900 ;
        RECT 72.430 44.700 72.750 44.760 ;
        RECT 73.265 44.715 73.555 44.760 ;
        RECT 80.250 44.900 80.570 44.960 ;
        RECT 86.320 44.945 86.460 45.100 ;
        RECT 84.910 44.900 85.200 44.945 ;
        RECT 80.250 44.760 85.200 44.900 ;
        RECT 80.250 44.700 80.570 44.760 ;
        RECT 84.910 44.715 85.200 44.760 ;
        RECT 86.245 44.715 86.535 44.945 ;
        RECT 86.690 44.700 87.010 44.960 ;
        RECT 48.985 44.420 50.210 44.560 ;
        RECT 48.985 44.375 49.275 44.420 ;
        RECT 49.890 44.360 50.210 44.420 ;
        RECT 50.440 44.420 52.420 44.560 ;
        RECT 52.625 44.560 52.915 44.605 ;
        RECT 53.815 44.560 54.105 44.605 ;
        RECT 56.335 44.560 56.625 44.605 ;
        RECT 52.625 44.420 56.625 44.560 ;
        RECT 50.440 44.265 50.580 44.420 ;
        RECT 52.625 44.375 52.915 44.420 ;
        RECT 53.815 44.375 54.105 44.420 ;
        RECT 56.335 44.375 56.625 44.420 ;
        RECT 65.045 44.560 65.335 44.605 ;
        RECT 66.235 44.560 66.525 44.605 ;
        RECT 68.755 44.560 69.045 44.605 ;
        RECT 65.045 44.420 69.045 44.560 ;
        RECT 65.045 44.375 65.335 44.420 ;
        RECT 66.235 44.375 66.525 44.420 ;
        RECT 68.755 44.375 69.045 44.420 ;
        RECT 72.865 44.560 73.155 44.605 ;
        RECT 74.055 44.560 74.345 44.605 ;
        RECT 76.575 44.560 76.865 44.605 ;
        RECT 72.865 44.420 76.865 44.560 ;
        RECT 72.865 44.375 73.155 44.420 ;
        RECT 74.055 44.375 74.345 44.420 ;
        RECT 76.575 44.375 76.865 44.420 ;
        RECT 81.655 44.560 81.945 44.605 ;
        RECT 84.175 44.560 84.465 44.605 ;
        RECT 85.365 44.560 85.655 44.605 ;
        RECT 81.655 44.420 85.655 44.560 ;
        RECT 81.655 44.375 81.945 44.420 ;
        RECT 84.175 44.375 84.465 44.420 ;
        RECT 85.365 44.375 85.655 44.420 ;
        RECT 31.070 44.220 31.360 44.265 ;
        RECT 33.170 44.220 33.460 44.265 ;
        RECT 34.740 44.220 35.030 44.265 ;
        RECT 31.070 44.080 35.030 44.220 ;
        RECT 31.070 44.035 31.360 44.080 ;
        RECT 33.170 44.035 33.460 44.080 ;
        RECT 34.740 44.035 35.030 44.080 ;
        RECT 38.890 44.220 39.180 44.265 ;
        RECT 40.990 44.220 41.280 44.265 ;
        RECT 42.560 44.220 42.850 44.265 ;
        RECT 38.890 44.080 42.850 44.220 ;
        RECT 38.890 44.035 39.180 44.080 ;
        RECT 40.990 44.035 41.280 44.080 ;
        RECT 42.560 44.035 42.850 44.080 ;
        RECT 50.365 44.035 50.655 44.265 ;
        RECT 52.230 44.220 52.520 44.265 ;
        RECT 54.330 44.220 54.620 44.265 ;
        RECT 55.900 44.220 56.190 44.265 ;
        RECT 52.230 44.080 56.190 44.220 ;
        RECT 52.230 44.035 52.520 44.080 ;
        RECT 54.330 44.035 54.620 44.080 ;
        RECT 55.900 44.035 56.190 44.080 ;
        RECT 64.650 44.220 64.940 44.265 ;
        RECT 66.750 44.220 67.040 44.265 ;
        RECT 68.320 44.220 68.610 44.265 ;
        RECT 64.650 44.080 68.610 44.220 ;
        RECT 64.650 44.035 64.940 44.080 ;
        RECT 66.750 44.035 67.040 44.080 ;
        RECT 68.320 44.035 68.610 44.080 ;
        RECT 71.065 44.220 71.355 44.265 ;
        RECT 71.510 44.220 71.830 44.280 ;
        RECT 71.065 44.080 71.830 44.220 ;
        RECT 71.065 44.035 71.355 44.080 ;
        RECT 71.510 44.020 71.830 44.080 ;
        RECT 72.470 44.220 72.760 44.265 ;
        RECT 74.570 44.220 74.860 44.265 ;
        RECT 76.140 44.220 76.430 44.265 ;
        RECT 72.470 44.080 76.430 44.220 ;
        RECT 72.470 44.035 72.760 44.080 ;
        RECT 74.570 44.035 74.860 44.080 ;
        RECT 76.140 44.035 76.430 44.080 ;
        RECT 82.090 44.220 82.380 44.265 ;
        RECT 83.660 44.220 83.950 44.265 ;
        RECT 85.760 44.220 86.050 44.265 ;
        RECT 82.090 44.080 86.050 44.220 ;
        RECT 82.090 44.035 82.380 44.080 ;
        RECT 83.660 44.035 83.950 44.080 ;
        RECT 85.760 44.035 86.050 44.080 ;
        RECT 36.550 43.880 36.870 43.940 ;
        RECT 39.770 43.880 40.090 43.940 ;
        RECT 45.305 43.880 45.595 43.925 ;
        RECT 46.670 43.880 46.990 43.940 ;
        RECT 30.660 43.740 46.990 43.880 ;
        RECT 16.310 43.680 16.630 43.740 ;
        RECT 18.150 43.680 18.470 43.740 ;
        RECT 23.225 43.695 23.515 43.740 ;
        RECT 36.550 43.680 36.870 43.740 ;
        RECT 39.770 43.680 40.090 43.740 ;
        RECT 45.305 43.695 45.595 43.740 ;
        RECT 46.670 43.680 46.990 43.740 ;
        RECT 58.630 43.880 58.950 43.940 ;
        RECT 60.470 43.880 60.790 43.940 ;
        RECT 58.630 43.740 60.790 43.880 ;
        RECT 58.630 43.680 58.950 43.740 ;
        RECT 60.470 43.680 60.790 43.740 ;
        RECT 76.570 43.880 76.890 43.940 ;
        RECT 78.885 43.880 79.175 43.925 ;
        RECT 76.570 43.740 79.175 43.880 ;
        RECT 76.570 43.680 76.890 43.740 ;
        RECT 78.885 43.695 79.175 43.740 ;
        RECT 79.330 43.680 79.650 43.940 ;
        RECT 12.100 43.060 89.840 43.540 ;
        RECT 18.150 42.860 18.470 42.920 ;
        RECT 21.385 42.860 21.675 42.905 ;
        RECT 18.150 42.720 21.675 42.860 ;
        RECT 18.150 42.660 18.470 42.720 ;
        RECT 21.385 42.675 21.675 42.720 ;
        RECT 18.610 42.520 18.930 42.580 ;
        RECT 15.480 42.380 18.930 42.520 ;
        RECT 21.460 42.520 21.600 42.675 ;
        RECT 22.290 42.660 22.610 42.920 ;
        RECT 23.670 42.660 23.990 42.920 ;
        RECT 30.570 42.860 30.890 42.920 ;
        RECT 24.220 42.720 30.890 42.860 ;
        RECT 24.220 42.520 24.360 42.720 ;
        RECT 30.570 42.660 30.890 42.720 ;
        RECT 32.410 42.660 32.730 42.920 ;
        RECT 35.170 42.860 35.490 42.920 ;
        RECT 37.470 42.860 37.790 42.920 ;
        RECT 40.230 42.860 40.550 42.920 ;
        RECT 41.165 42.860 41.455 42.905 ;
        RECT 35.170 42.720 40.000 42.860 ;
        RECT 35.170 42.660 35.490 42.720 ;
        RECT 37.470 42.660 37.790 42.720 ;
        RECT 21.460 42.380 24.360 42.520 ;
        RECT 26.010 42.520 26.300 42.565 ;
        RECT 28.110 42.520 28.400 42.565 ;
        RECT 29.680 42.520 29.970 42.565 ;
        RECT 26.010 42.380 29.970 42.520 ;
        RECT 15.480 42.225 15.620 42.380 ;
        RECT 18.610 42.320 18.930 42.380 ;
        RECT 26.010 42.335 26.300 42.380 ;
        RECT 28.110 42.335 28.400 42.380 ;
        RECT 29.680 42.335 29.970 42.380 ;
        RECT 34.750 42.520 35.040 42.565 ;
        RECT 36.850 42.520 37.140 42.565 ;
        RECT 38.420 42.520 38.710 42.565 ;
        RECT 34.750 42.380 38.710 42.520 ;
        RECT 39.860 42.520 40.000 42.720 ;
        RECT 40.230 42.720 41.455 42.860 ;
        RECT 40.230 42.660 40.550 42.720 ;
        RECT 41.165 42.675 41.455 42.720 ;
        RECT 41.610 42.660 41.930 42.920 ;
        RECT 42.545 42.675 42.835 42.905 ;
        RECT 42.620 42.520 42.760 42.675 ;
        RECT 63.230 42.660 63.550 42.920 ;
        RECT 64.165 42.860 64.455 42.905 ;
        RECT 64.610 42.860 64.930 42.920 ;
        RECT 64.165 42.720 64.930 42.860 ;
        RECT 64.165 42.675 64.455 42.720 ;
        RECT 64.610 42.660 64.930 42.720 ;
        RECT 71.525 42.860 71.815 42.905 ;
        RECT 72.430 42.860 72.750 42.920 ;
        RECT 71.525 42.720 72.750 42.860 ;
        RECT 71.525 42.675 71.815 42.720 ;
        RECT 72.430 42.660 72.750 42.720 ;
        RECT 78.870 42.860 79.190 42.920 ;
        RECT 79.805 42.860 80.095 42.905 ;
        RECT 78.870 42.720 80.095 42.860 ;
        RECT 78.870 42.660 79.190 42.720 ;
        RECT 79.805 42.675 80.095 42.720 ;
        RECT 39.860 42.380 42.760 42.520 ;
        RECT 81.670 42.520 81.960 42.565 ;
        RECT 83.770 42.520 84.060 42.565 ;
        RECT 85.340 42.520 85.630 42.565 ;
        RECT 81.670 42.380 85.630 42.520 ;
        RECT 34.750 42.335 35.040 42.380 ;
        RECT 36.850 42.335 37.140 42.380 ;
        RECT 38.420 42.335 38.710 42.380 ;
        RECT 81.670 42.335 81.960 42.380 ;
        RECT 83.770 42.335 84.060 42.380 ;
        RECT 85.340 42.335 85.630 42.380 ;
        RECT 15.405 41.995 15.695 42.225 ;
        RECT 16.785 42.180 17.075 42.225 ;
        RECT 18.150 42.180 18.470 42.240 ;
        RECT 16.785 42.040 18.470 42.180 ;
        RECT 16.785 41.995 17.075 42.040 ;
        RECT 18.150 41.980 18.470 42.040 ;
        RECT 20.450 42.180 20.770 42.240 ;
        RECT 22.750 42.180 23.070 42.240 ;
        RECT 25.525 42.180 25.815 42.225 ;
        RECT 20.450 42.040 25.815 42.180 ;
        RECT 20.450 41.980 20.770 42.040 ;
        RECT 22.750 41.980 23.070 42.040 ;
        RECT 25.525 41.995 25.815 42.040 ;
        RECT 26.405 42.180 26.695 42.225 ;
        RECT 27.595 42.180 27.885 42.225 ;
        RECT 30.115 42.180 30.405 42.225 ;
        RECT 26.405 42.040 30.405 42.180 ;
        RECT 26.405 41.995 26.695 42.040 ;
        RECT 27.595 41.995 27.885 42.040 ;
        RECT 30.115 41.995 30.405 42.040 ;
        RECT 35.145 42.180 35.435 42.225 ;
        RECT 36.335 42.180 36.625 42.225 ;
        RECT 38.855 42.180 39.145 42.225 ;
        RECT 35.145 42.040 39.145 42.180 ;
        RECT 35.145 41.995 35.435 42.040 ;
        RECT 36.335 41.995 36.625 42.040 ;
        RECT 38.855 41.995 39.145 42.040 ;
        RECT 52.190 42.180 52.510 42.240 ;
        RECT 52.665 42.180 52.955 42.225 ;
        RECT 52.190 42.040 52.955 42.180 ;
        RECT 52.190 41.980 52.510 42.040 ;
        RECT 52.665 41.995 52.955 42.040 ;
        RECT 59.565 42.180 59.855 42.225 ;
        RECT 61.850 42.180 62.170 42.240 ;
        RECT 62.450 42.180 62.740 42.225 ;
        RECT 59.565 42.040 62.740 42.180 ;
        RECT 59.565 41.995 59.855 42.040 ;
        RECT 61.850 41.980 62.170 42.040 ;
        RECT 62.450 41.995 62.740 42.040 ;
        RECT 67.370 41.980 67.690 42.240 ;
        RECT 81.170 41.980 81.490 42.240 ;
        RECT 82.065 42.180 82.355 42.225 ;
        RECT 83.255 42.180 83.545 42.225 ;
        RECT 85.775 42.180 86.065 42.225 ;
        RECT 82.065 42.040 86.065 42.180 ;
        RECT 82.065 41.995 82.355 42.040 ;
        RECT 83.255 41.995 83.545 42.040 ;
        RECT 85.775 41.995 86.065 42.040 ;
        RECT 14.945 41.840 15.235 41.885 ;
        RECT 20.910 41.840 21.230 41.900 ;
        RECT 25.970 41.840 26.290 41.900 ;
        RECT 14.945 41.700 21.230 41.840 ;
        RECT 14.945 41.655 15.235 41.700 ;
        RECT 20.910 41.640 21.230 41.700 ;
        RECT 22.970 41.700 26.290 41.840 ;
        RECT 22.970 41.670 23.110 41.700 ;
        RECT 17.245 41.500 17.535 41.545 ;
        RECT 17.690 41.500 18.010 41.560 ;
        RECT 17.245 41.360 18.010 41.500 ;
        RECT 17.245 41.315 17.535 41.360 ;
        RECT 17.690 41.300 18.010 41.360 ;
        RECT 18.150 41.545 18.470 41.560 ;
        RECT 18.150 41.315 18.535 41.545 ;
        RECT 19.990 41.500 20.310 41.560 ;
        RECT 21.370 41.545 21.690 41.560 ;
        RECT 22.840 41.545 23.110 41.670 ;
        RECT 25.970 41.640 26.290 41.700 ;
        RECT 26.860 41.840 27.150 41.885 ;
        RECT 29.650 41.840 29.970 41.900 ;
        RECT 32.885 41.840 33.175 41.885 ;
        RECT 26.860 41.700 29.970 41.840 ;
        RECT 26.860 41.655 27.150 41.700 ;
        RECT 29.650 41.640 29.970 41.700 ;
        RECT 31.120 41.700 33.175 41.840 ;
        RECT 20.465 41.500 20.755 41.545 ;
        RECT 18.700 41.360 20.755 41.500 ;
        RECT 18.150 41.300 18.470 41.315 ;
        RECT 17.780 41.160 17.920 41.300 ;
        RECT 18.700 41.160 18.840 41.360 ;
        RECT 19.990 41.300 20.310 41.360 ;
        RECT 20.465 41.315 20.755 41.360 ;
        RECT 21.370 41.315 21.755 41.545 ;
        RECT 22.765 41.530 23.110 41.545 ;
        RECT 22.765 41.315 23.055 41.530 ;
        RECT 21.370 41.300 21.690 41.315 ;
        RECT 17.780 41.020 18.840 41.160 ;
        RECT 19.070 40.960 19.390 41.220 ;
        RECT 19.530 41.160 19.850 41.220 ;
        RECT 20.910 41.160 21.230 41.220 ;
        RECT 23.765 41.160 24.055 41.205 ;
        RECT 19.530 41.020 24.055 41.160 ;
        RECT 19.530 40.960 19.850 41.020 ;
        RECT 20.910 40.960 21.230 41.020 ;
        RECT 23.765 40.975 24.055 41.020 ;
        RECT 24.605 41.160 24.895 41.205 ;
        RECT 26.430 41.160 26.750 41.220 ;
        RECT 31.120 41.160 31.260 41.700 ;
        RECT 32.885 41.655 33.175 41.700 ;
        RECT 33.790 41.640 34.110 41.900 ;
        RECT 34.265 41.840 34.555 41.885 ;
        RECT 34.710 41.840 35.030 41.900 ;
        RECT 34.265 41.700 35.030 41.840 ;
        RECT 34.265 41.655 34.555 41.700 ;
        RECT 34.710 41.640 35.030 41.700 ;
        RECT 41.150 41.840 41.470 41.900 ;
        RECT 45.765 41.840 46.055 41.885 ;
        RECT 41.150 41.700 46.055 41.840 ;
        RECT 41.150 41.640 41.470 41.700 ;
        RECT 45.765 41.655 46.055 41.700 ;
        RECT 46.670 41.640 46.990 41.900 ;
        RECT 55.885 41.655 56.175 41.885 ;
        RECT 33.330 41.300 33.650 41.560 ;
        RECT 35.600 41.500 35.890 41.545 ;
        RECT 36.090 41.500 36.410 41.560 ;
        RECT 35.600 41.360 36.410 41.500 ;
        RECT 35.600 41.315 35.890 41.360 ;
        RECT 36.090 41.300 36.410 41.360 ;
        RECT 42.070 41.545 42.390 41.560 ;
        RECT 42.070 41.315 42.675 41.545 ;
        RECT 43.465 41.500 43.755 41.545 ;
        RECT 46.225 41.500 46.515 41.545 ;
        RECT 43.465 41.360 46.515 41.500 ;
        RECT 55.960 41.500 56.100 41.655 ;
        RECT 60.010 41.640 60.330 41.900 ;
        RECT 60.470 41.840 60.790 41.900 ;
        RECT 61.405 41.840 61.695 41.885 ;
        RECT 60.470 41.700 61.695 41.840 ;
        RECT 60.470 41.640 60.790 41.700 ;
        RECT 61.405 41.655 61.695 41.700 ;
        RECT 69.670 41.840 69.990 41.900 ;
        RECT 71.065 41.840 71.355 41.885 ;
        RECT 69.670 41.700 71.355 41.840 ;
        RECT 69.670 41.640 69.990 41.700 ;
        RECT 71.065 41.655 71.355 41.700 ;
        RECT 72.890 41.640 73.210 41.900 ;
        RECT 73.350 41.640 73.670 41.900 ;
        RECT 73.825 41.840 74.115 41.885 ;
        RECT 74.270 41.840 74.590 41.900 ;
        RECT 73.825 41.700 74.590 41.840 ;
        RECT 73.825 41.655 74.115 41.700 ;
        RECT 74.270 41.640 74.590 41.700 ;
        RECT 74.745 41.840 75.035 41.885 ;
        RECT 75.190 41.840 75.510 41.900 ;
        RECT 74.745 41.700 75.510 41.840 ;
        RECT 74.745 41.655 75.035 41.700 ;
        RECT 75.190 41.640 75.510 41.700 ;
        RECT 76.570 41.840 76.890 41.900 ;
        RECT 77.045 41.840 77.335 41.885 ;
        RECT 76.570 41.700 77.335 41.840 ;
        RECT 76.570 41.640 76.890 41.700 ;
        RECT 77.045 41.655 77.335 41.700 ;
        RECT 77.490 41.840 77.810 41.900 ;
        RECT 77.965 41.840 78.255 41.885 ;
        RECT 77.490 41.700 78.255 41.840 ;
        RECT 77.490 41.640 77.810 41.700 ;
        RECT 77.965 41.655 78.255 41.700 ;
        RECT 78.885 41.840 79.175 41.885 ;
        RECT 79.790 41.840 80.110 41.900 ;
        RECT 78.885 41.700 80.110 41.840 ;
        RECT 78.885 41.655 79.175 41.700 ;
        RECT 79.790 41.640 80.110 41.700 ;
        RECT 61.865 41.500 62.155 41.545 ;
        RECT 62.310 41.500 62.630 41.560 ;
        RECT 55.960 41.360 62.630 41.500 ;
        RECT 43.465 41.315 43.755 41.360 ;
        RECT 46.225 41.315 46.515 41.360 ;
        RECT 61.865 41.315 62.155 41.360 ;
        RECT 42.070 41.300 42.390 41.315 ;
        RECT 62.310 41.300 62.630 41.360 ;
        RECT 66.465 41.500 66.755 41.545 ;
        RECT 71.510 41.500 71.830 41.560 ;
        RECT 66.465 41.360 71.830 41.500 ;
        RECT 66.465 41.315 66.755 41.360 ;
        RECT 71.510 41.300 71.830 41.360 ;
        RECT 78.410 41.500 78.730 41.560 ;
        RECT 79.330 41.500 79.650 41.560 ;
        RECT 78.410 41.360 79.650 41.500 ;
        RECT 78.410 41.300 78.730 41.360 ;
        RECT 79.330 41.300 79.650 41.360 ;
        RECT 82.520 41.500 82.810 41.545 ;
        RECT 84.390 41.500 84.710 41.560 ;
        RECT 82.520 41.360 84.710 41.500 ;
        RECT 82.520 41.315 82.810 41.360 ;
        RECT 84.390 41.300 84.710 41.360 ;
        RECT 24.605 41.020 31.260 41.160 ;
        RECT 56.345 41.160 56.635 41.205 ;
        RECT 56.790 41.160 57.110 41.220 ;
        RECT 56.345 41.020 57.110 41.160 ;
        RECT 24.605 40.975 24.895 41.020 ;
        RECT 26.430 40.960 26.750 41.020 ;
        RECT 56.345 40.975 56.635 41.020 ;
        RECT 56.790 40.960 57.110 41.020 ;
        RECT 65.990 40.960 66.310 41.220 ;
        RECT 70.145 41.160 70.435 41.205 ;
        RECT 72.430 41.160 72.750 41.220 ;
        RECT 70.145 41.020 72.750 41.160 ;
        RECT 70.145 40.975 70.435 41.020 ;
        RECT 72.430 40.960 72.750 41.020 ;
        RECT 74.730 41.160 75.050 41.220 ;
        RECT 78.870 41.160 79.190 41.220 ;
        RECT 86.230 41.160 86.550 41.220 ;
        RECT 74.730 41.020 86.550 41.160 ;
        RECT 74.730 40.960 75.050 41.020 ;
        RECT 78.870 40.960 79.190 41.020 ;
        RECT 86.230 40.960 86.550 41.020 ;
        RECT 87.610 41.160 87.930 41.220 ;
        RECT 88.085 41.160 88.375 41.205 ;
        RECT 87.610 41.020 88.375 41.160 ;
        RECT 87.610 40.960 87.930 41.020 ;
        RECT 88.085 40.975 88.375 41.020 ;
        RECT 12.100 40.340 89.840 40.820 ;
        RECT 25.970 40.140 26.290 40.200 ;
        RECT 22.000 40.000 26.290 40.140 ;
        RECT 20.465 39.460 20.755 39.505 ;
        RECT 22.000 39.460 22.140 40.000 ;
        RECT 25.970 39.940 26.290 40.000 ;
        RECT 34.250 40.140 34.570 40.200 ;
        RECT 38.405 40.140 38.695 40.185 ;
        RECT 34.250 40.000 38.695 40.140 ;
        RECT 34.250 39.940 34.570 40.000 ;
        RECT 38.405 39.955 38.695 40.000 ;
        RECT 40.245 40.140 40.535 40.185 ;
        RECT 41.150 40.140 41.470 40.200 ;
        RECT 40.245 40.000 41.470 40.140 ;
        RECT 40.245 39.955 40.535 40.000 ;
        RECT 22.290 39.800 22.610 39.860 ;
        RECT 23.990 39.800 24.280 39.845 ;
        RECT 30.885 39.800 31.175 39.845 ;
        RECT 22.290 39.660 24.280 39.800 ;
        RECT 22.290 39.600 22.610 39.660 ;
        RECT 23.990 39.615 24.280 39.660 ;
        RECT 24.680 39.660 31.175 39.800 ;
        RECT 20.465 39.320 22.140 39.460 ;
        RECT 20.465 39.275 20.755 39.320 ;
        RECT 22.750 39.260 23.070 39.520 ;
        RECT 24.680 39.460 24.820 39.660 ;
        RECT 30.885 39.615 31.175 39.660 ;
        RECT 31.965 39.615 32.255 39.845 ;
        RECT 36.105 39.800 36.395 39.845 ;
        RECT 40.320 39.800 40.460 39.955 ;
        RECT 41.150 39.940 41.470 40.000 ;
        RECT 50.810 40.140 51.130 40.200 ;
        RECT 54.045 40.140 54.335 40.185 ;
        RECT 50.810 40.000 54.335 40.140 ;
        RECT 50.810 39.940 51.130 40.000 ;
        RECT 54.045 39.955 54.335 40.000 ;
        RECT 58.185 40.140 58.475 40.185 ;
        RECT 61.390 40.140 61.710 40.200 ;
        RECT 58.185 40.000 61.710 40.140 ;
        RECT 58.185 39.955 58.475 40.000 ;
        RECT 61.390 39.940 61.710 40.000 ;
        RECT 62.325 40.140 62.615 40.185 ;
        RECT 62.770 40.140 63.090 40.200 ;
        RECT 62.325 40.000 63.090 40.140 ;
        RECT 62.325 39.955 62.615 40.000 ;
        RECT 62.770 39.940 63.090 40.000 ;
        RECT 63.245 40.140 63.535 40.185 ;
        RECT 66.450 40.140 66.770 40.200 ;
        RECT 63.245 40.000 66.770 40.140 ;
        RECT 63.245 39.955 63.535 40.000 ;
        RECT 66.450 39.940 66.770 40.000 ;
        RECT 66.925 40.140 67.215 40.185 ;
        RECT 71.970 40.140 72.290 40.200 ;
        RECT 66.925 40.000 72.290 40.140 ;
        RECT 66.925 39.955 67.215 40.000 ;
        RECT 71.970 39.940 72.290 40.000 ;
        RECT 74.270 39.940 74.590 40.200 ;
        RECT 77.045 40.140 77.335 40.185 ;
        RECT 77.950 40.140 78.270 40.200 ;
        RECT 77.045 40.000 78.270 40.140 ;
        RECT 77.045 39.955 77.335 40.000 ;
        RECT 77.950 39.940 78.270 40.000 ;
        RECT 80.265 40.140 80.555 40.185 ;
        RECT 82.550 40.140 82.870 40.200 ;
        RECT 80.265 40.000 82.870 40.140 ;
        RECT 80.265 39.955 80.555 40.000 ;
        RECT 82.550 39.940 82.870 40.000 ;
        RECT 84.390 39.940 84.710 40.200 ;
        RECT 84.850 39.940 85.170 40.200 ;
        RECT 86.690 40.140 87.010 40.200 ;
        RECT 86.320 40.000 87.010 40.140 ;
        RECT 36.105 39.660 40.460 39.800 ;
        RECT 59.025 39.800 59.315 39.845 ;
        RECT 59.025 39.660 59.780 39.800 ;
        RECT 36.105 39.615 36.395 39.660 ;
        RECT 59.025 39.615 59.315 39.660 ;
        RECT 23.300 39.320 24.820 39.460 ;
        RECT 26.890 39.460 27.210 39.520 ;
        RECT 32.040 39.460 32.180 39.615 ;
        RECT 26.890 39.320 32.180 39.460 ;
        RECT 39.325 39.460 39.615 39.505 ;
        RECT 40.230 39.460 40.550 39.520 ;
        RECT 39.325 39.320 40.550 39.460 ;
        RECT 20.910 38.920 21.230 39.180 ;
        RECT 22.305 39.120 22.595 39.165 ;
        RECT 23.300 39.120 23.440 39.320 ;
        RECT 26.890 39.260 27.210 39.320 ;
        RECT 39.325 39.275 39.615 39.320 ;
        RECT 40.230 39.260 40.550 39.320 ;
        RECT 40.705 39.275 40.995 39.505 ;
        RECT 54.045 39.275 54.335 39.505 ;
        RECT 22.305 38.980 23.440 39.120 ;
        RECT 23.645 39.120 23.935 39.165 ;
        RECT 24.835 39.120 25.125 39.165 ;
        RECT 27.355 39.120 27.645 39.165 ;
        RECT 23.645 38.980 27.645 39.120 ;
        RECT 22.305 38.935 22.595 38.980 ;
        RECT 23.645 38.935 23.935 38.980 ;
        RECT 24.835 38.935 25.125 38.980 ;
        RECT 27.355 38.935 27.645 38.980 ;
        RECT 39.770 39.120 40.090 39.180 ;
        RECT 40.780 39.120 40.920 39.275 ;
        RECT 39.770 38.980 40.920 39.120 ;
        RECT 54.120 39.120 54.260 39.275 ;
        RECT 54.950 39.260 55.270 39.520 ;
        RECT 55.410 39.260 55.730 39.520 ;
        RECT 55.885 39.460 56.175 39.505 ;
        RECT 56.330 39.460 56.650 39.520 ;
        RECT 55.885 39.320 56.650 39.460 ;
        RECT 55.885 39.275 56.175 39.320 ;
        RECT 56.330 39.260 56.650 39.320 ;
        RECT 55.500 39.120 55.640 39.260 ;
        RECT 54.120 38.980 55.640 39.120 ;
        RECT 39.770 38.920 40.090 38.980 ;
        RECT 56.790 38.920 57.110 39.180 ;
        RECT 59.640 39.120 59.780 39.660 ;
        RECT 60.025 39.615 60.315 39.845 ;
        RECT 71.050 39.800 71.370 39.860 ;
        RECT 68.610 39.660 71.370 39.800 ;
        RECT 60.100 39.460 60.240 39.615 ;
        RECT 60.485 39.460 60.775 39.505 ;
        RECT 62.310 39.460 62.630 39.520 ;
        RECT 64.165 39.460 64.455 39.505 ;
        RECT 68.610 39.460 68.750 39.660 ;
        RECT 71.050 39.600 71.370 39.660 ;
        RECT 71.600 39.660 78.180 39.800 ;
        RECT 71.600 39.505 71.740 39.660 ;
        RECT 60.100 39.320 68.750 39.460 ;
        RECT 69.685 39.460 69.975 39.505 ;
        RECT 69.685 39.320 71.280 39.460 ;
        RECT 60.485 39.275 60.775 39.320 ;
        RECT 62.310 39.260 62.630 39.320 ;
        RECT 64.165 39.275 64.455 39.320 ;
        RECT 69.685 39.275 69.975 39.320 ;
        RECT 61.850 39.120 62.170 39.180 ;
        RECT 62.770 39.120 63.090 39.180 ;
        RECT 59.640 38.980 63.090 39.120 ;
        RECT 61.850 38.920 62.170 38.980 ;
        RECT 62.770 38.920 63.090 38.980 ;
        RECT 65.545 38.935 65.835 39.165 ;
        RECT 71.140 39.120 71.280 39.320 ;
        RECT 71.525 39.275 71.815 39.505 ;
        RECT 72.905 39.275 73.195 39.505 ;
        RECT 73.825 39.460 74.115 39.505 ;
        RECT 74.270 39.460 74.590 39.520 ;
        RECT 73.825 39.320 74.590 39.460 ;
        RECT 73.825 39.275 74.115 39.320 ;
        RECT 72.980 39.120 73.120 39.275 ;
        RECT 74.270 39.260 74.590 39.320 ;
        RECT 75.205 39.275 75.495 39.505 ;
        RECT 74.730 39.120 75.050 39.180 ;
        RECT 71.140 38.980 75.050 39.120 ;
        RECT 75.280 39.120 75.420 39.275 ;
        RECT 76.110 39.260 76.430 39.520 ;
        RECT 78.040 39.505 78.180 39.660 ;
        RECT 78.870 39.600 79.190 39.860 ;
        RECT 79.790 39.800 80.110 39.860 ;
        RECT 86.320 39.845 86.460 40.000 ;
        RECT 86.690 39.940 87.010 40.000 ;
        RECT 79.790 39.660 86.000 39.800 ;
        RECT 79.790 39.600 80.110 39.660 ;
        RECT 77.965 39.460 78.255 39.505 ;
        RECT 78.410 39.460 78.730 39.520 ;
        RECT 77.965 39.320 78.730 39.460 ;
        RECT 77.965 39.275 78.255 39.320 ;
        RECT 78.410 39.260 78.730 39.320 ;
        RECT 79.330 39.260 79.650 39.520 ;
        RECT 81.185 39.490 81.475 39.505 ;
        RECT 81.630 39.490 81.950 39.510 ;
        RECT 81.185 39.350 81.950 39.490 ;
        RECT 81.185 39.275 81.475 39.350 ;
        RECT 81.630 39.250 81.950 39.350 ;
        RECT 82.105 39.290 82.395 39.520 ;
        RECT 82.595 39.505 82.915 39.520 ;
        RECT 82.580 39.460 82.915 39.505 ;
        RECT 83.255 39.460 83.545 39.505 ;
        RECT 85.310 39.460 85.630 39.520 ;
        RECT 85.860 39.505 86.000 39.660 ;
        RECT 86.245 39.615 86.535 39.845 ;
        RECT 82.580 39.320 83.080 39.460 ;
        RECT 83.255 39.320 85.630 39.460 ;
        RECT 76.570 39.120 76.890 39.180 ;
        RECT 75.280 38.980 76.890 39.120 ;
        RECT 23.250 38.780 23.540 38.825 ;
        RECT 25.350 38.780 25.640 38.825 ;
        RECT 26.920 38.780 27.210 38.825 ;
        RECT 23.250 38.640 27.210 38.780 ;
        RECT 23.250 38.595 23.540 38.640 ;
        RECT 25.350 38.595 25.640 38.640 ;
        RECT 26.920 38.595 27.210 38.640 ;
        RECT 34.725 38.780 35.015 38.825 ;
        RECT 37.470 38.780 37.790 38.840 ;
        RECT 65.620 38.780 65.760 38.935 ;
        RECT 74.730 38.920 75.050 38.980 ;
        RECT 76.570 38.920 76.890 38.980 ;
        RECT 77.030 39.120 77.350 39.180 ;
        RECT 77.030 39.080 80.480 39.120 ;
        RECT 82.180 39.080 82.320 39.290 ;
        RECT 82.580 39.275 82.915 39.320 ;
        RECT 83.255 39.275 83.545 39.320 ;
        RECT 82.595 39.260 82.915 39.275 ;
        RECT 85.310 39.260 85.630 39.320 ;
        RECT 85.785 39.275 86.075 39.505 ;
        RECT 86.690 39.260 87.010 39.520 ;
        RECT 87.610 39.260 87.930 39.520 ;
        RECT 77.030 38.980 82.320 39.080 ;
        RECT 77.030 38.920 77.350 38.980 ;
        RECT 80.340 38.940 82.320 38.980 ;
        RECT 34.725 38.640 37.790 38.780 ;
        RECT 34.725 38.595 35.015 38.640 ;
        RECT 37.470 38.580 37.790 38.640 ;
        RECT 62.400 38.640 65.760 38.780 ;
        RECT 23.670 38.440 23.990 38.500 ;
        RECT 29.665 38.440 29.955 38.485 ;
        RECT 23.670 38.300 29.955 38.440 ;
        RECT 23.670 38.240 23.990 38.300 ;
        RECT 29.665 38.255 29.955 38.300 ;
        RECT 30.110 38.240 30.430 38.500 ;
        RECT 30.570 38.440 30.890 38.500 ;
        RECT 31.045 38.440 31.335 38.485 ;
        RECT 30.570 38.300 31.335 38.440 ;
        RECT 30.570 38.240 30.890 38.300 ;
        RECT 31.045 38.255 31.335 38.300 ;
        RECT 33.790 38.240 34.110 38.500 ;
        RECT 56.330 38.240 56.650 38.500 ;
        RECT 59.105 38.440 59.395 38.485 ;
        RECT 60.930 38.440 61.250 38.500 ;
        RECT 62.400 38.485 62.540 38.640 ;
        RECT 62.325 38.440 62.615 38.485 ;
        RECT 59.105 38.300 62.615 38.440 ;
        RECT 59.105 38.255 59.395 38.300 ;
        RECT 60.930 38.240 61.250 38.300 ;
        RECT 62.325 38.255 62.615 38.300 ;
        RECT 65.070 38.240 65.390 38.500 ;
        RECT 65.620 38.440 65.760 38.640 ;
        RECT 68.765 38.780 69.055 38.825 ;
        RECT 82.550 38.780 82.870 38.840 ;
        RECT 68.765 38.640 82.870 38.780 ;
        RECT 68.765 38.595 69.055 38.640 ;
        RECT 82.550 38.580 82.870 38.640 ;
        RECT 70.130 38.440 70.450 38.500 ;
        RECT 65.620 38.300 70.450 38.440 ;
        RECT 70.130 38.240 70.450 38.300 ;
        RECT 70.590 38.240 70.910 38.500 ;
        RECT 71.985 38.440 72.275 38.485 ;
        RECT 75.190 38.440 75.510 38.500 ;
        RECT 71.985 38.300 75.510 38.440 ;
        RECT 71.985 38.255 72.275 38.300 ;
        RECT 75.190 38.240 75.510 38.300 ;
        RECT 75.650 38.440 75.970 38.500 ;
        RECT 81.630 38.440 81.950 38.500 ;
        RECT 75.650 38.300 81.950 38.440 ;
        RECT 75.650 38.240 75.970 38.300 ;
        RECT 81.630 38.240 81.950 38.300 ;
        RECT 12.100 37.620 89.840 38.100 ;
        RECT 25.525 37.420 25.815 37.465 ;
        RECT 25.970 37.420 26.290 37.480 ;
        RECT 25.525 37.280 26.290 37.420 ;
        RECT 25.525 37.235 25.815 37.280 ;
        RECT 25.970 37.220 26.290 37.280 ;
        RECT 39.785 37.420 40.075 37.465 ;
        RECT 41.150 37.420 41.470 37.480 ;
        RECT 39.785 37.280 41.470 37.420 ;
        RECT 39.785 37.235 40.075 37.280 ;
        RECT 41.150 37.220 41.470 37.280 ;
        RECT 59.550 37.220 59.870 37.480 ;
        RECT 66.465 37.420 66.755 37.465 ;
        RECT 66.910 37.420 67.230 37.480 ;
        RECT 66.465 37.280 67.230 37.420 ;
        RECT 66.465 37.235 66.755 37.280 ;
        RECT 66.910 37.220 67.230 37.280 ;
        RECT 69.685 37.420 69.975 37.465 ;
        RECT 77.030 37.420 77.350 37.480 ;
        RECT 86.690 37.420 87.010 37.480 ;
        RECT 69.685 37.280 77.350 37.420 ;
        RECT 69.685 37.235 69.975 37.280 ;
        RECT 77.030 37.220 77.350 37.280 ;
        RECT 82.180 37.280 87.010 37.420 ;
        RECT 19.990 37.080 20.310 37.140 ;
        RECT 26.890 37.080 27.210 37.140 ;
        RECT 19.990 36.940 27.210 37.080 ;
        RECT 19.990 36.880 20.310 36.940 ;
        RECT 26.890 36.880 27.210 36.940 ;
        RECT 28.270 37.080 28.560 37.125 ;
        RECT 29.840 37.080 30.130 37.125 ;
        RECT 31.940 37.080 32.230 37.125 ;
        RECT 28.270 36.940 32.230 37.080 ;
        RECT 28.270 36.895 28.560 36.940 ;
        RECT 29.840 36.895 30.130 36.940 ;
        RECT 31.940 36.895 32.230 36.940 ;
        RECT 33.370 37.080 33.660 37.125 ;
        RECT 35.470 37.080 35.760 37.125 ;
        RECT 37.040 37.080 37.330 37.125 ;
        RECT 33.370 36.940 37.330 37.080 ;
        RECT 33.370 36.895 33.660 36.940 ;
        RECT 35.470 36.895 35.760 36.940 ;
        RECT 37.040 36.895 37.330 36.940 ;
        RECT 77.490 36.880 77.810 37.140 ;
        RECT 80.250 36.880 80.570 37.140 ;
        RECT 27.835 36.740 28.125 36.785 ;
        RECT 30.355 36.740 30.645 36.785 ;
        RECT 31.545 36.740 31.835 36.785 ;
        RECT 27.835 36.600 31.835 36.740 ;
        RECT 27.835 36.555 28.125 36.600 ;
        RECT 30.355 36.555 30.645 36.600 ;
        RECT 31.545 36.555 31.835 36.600 ;
        RECT 33.765 36.740 34.055 36.785 ;
        RECT 34.955 36.740 35.245 36.785 ;
        RECT 37.475 36.740 37.765 36.785 ;
        RECT 76.110 36.740 76.430 36.800 ;
        RECT 33.765 36.600 37.765 36.740 ;
        RECT 33.765 36.555 34.055 36.600 ;
        RECT 34.955 36.555 35.245 36.600 ;
        RECT 37.475 36.555 37.765 36.600 ;
        RECT 60.100 36.600 63.460 36.740 ;
        RECT 32.425 36.400 32.715 36.445 ;
        RECT 32.885 36.400 33.175 36.445 ;
        RECT 32.425 36.260 33.560 36.400 ;
        RECT 32.425 36.215 32.715 36.260 ;
        RECT 32.885 36.215 33.175 36.260 ;
        RECT 30.110 36.060 30.430 36.120 ;
        RECT 31.090 36.060 31.380 36.105 ;
        RECT 30.110 35.920 31.380 36.060 ;
        RECT 30.110 35.860 30.430 35.920 ;
        RECT 31.090 35.875 31.380 35.920 ;
        RECT 33.420 35.720 33.560 36.260 ;
        RECT 34.220 36.215 34.510 36.445 ;
        RECT 56.330 36.400 56.650 36.460 ;
        RECT 60.100 36.445 60.240 36.600 ;
        RECT 59.105 36.400 59.395 36.445 ;
        RECT 56.330 36.260 59.395 36.400 ;
        RECT 33.790 36.060 34.110 36.120 ;
        RECT 34.340 36.060 34.480 36.215 ;
        RECT 56.330 36.200 56.650 36.260 ;
        RECT 59.105 36.215 59.395 36.260 ;
        RECT 60.025 36.215 60.315 36.445 ;
        RECT 60.470 36.200 60.790 36.460 ;
        RECT 60.930 36.400 61.250 36.460 ;
        RECT 63.320 36.445 63.460 36.600 ;
        RECT 72.060 36.600 76.430 36.740 ;
        RECT 77.580 36.740 77.720 36.880 ;
        RECT 82.180 36.740 82.320 37.280 ;
        RECT 86.690 37.220 87.010 37.280 ;
        RECT 83.010 36.880 83.330 37.140 ;
        RECT 77.580 36.600 82.320 36.740 ;
        RECT 83.100 36.740 83.240 36.880 ;
        RECT 83.100 36.600 86.000 36.740 ;
        RECT 61.405 36.400 61.695 36.445 ;
        RECT 60.930 36.260 61.695 36.400 ;
        RECT 60.930 36.200 61.250 36.260 ;
        RECT 61.405 36.215 61.695 36.260 ;
        RECT 63.245 36.400 63.535 36.445 ;
        RECT 65.070 36.400 65.390 36.460 ;
        RECT 63.245 36.260 65.390 36.400 ;
        RECT 63.245 36.215 63.535 36.260 ;
        RECT 65.070 36.200 65.390 36.260 ;
        RECT 67.385 36.400 67.675 36.445 ;
        RECT 67.830 36.400 68.150 36.460 ;
        RECT 67.385 36.260 68.150 36.400 ;
        RECT 67.385 36.215 67.675 36.260 ;
        RECT 67.830 36.200 68.150 36.260 ;
        RECT 69.225 36.400 69.515 36.445 ;
        RECT 70.590 36.400 70.910 36.460 ;
        RECT 69.225 36.260 70.910 36.400 ;
        RECT 69.225 36.215 69.515 36.260 ;
        RECT 70.590 36.200 70.910 36.260 ;
        RECT 72.060 36.120 72.200 36.600 ;
        RECT 76.110 36.540 76.430 36.600 ;
        RECT 72.905 36.400 73.195 36.445 ;
        RECT 77.045 36.400 77.335 36.445 ;
        RECT 77.490 36.400 77.810 36.460 ;
        RECT 78.040 36.445 78.180 36.600 ;
        RECT 72.905 36.260 77.810 36.400 ;
        RECT 72.905 36.215 73.195 36.260 ;
        RECT 77.045 36.215 77.335 36.260 ;
        RECT 77.490 36.200 77.810 36.260 ;
        RECT 77.965 36.215 78.255 36.445 ;
        RECT 78.425 36.215 78.715 36.445 ;
        RECT 78.885 36.400 79.175 36.445 ;
        RECT 79.790 36.400 80.110 36.460 ;
        RECT 82.180 36.445 82.320 36.600 ;
        RECT 85.860 36.460 86.000 36.600 ;
        RECT 81.185 36.400 81.475 36.445 ;
        RECT 78.885 36.260 81.475 36.400 ;
        RECT 78.885 36.215 79.175 36.260 ;
        RECT 33.790 35.920 34.480 36.060 ;
        RECT 71.525 36.060 71.815 36.105 ;
        RECT 71.970 36.060 72.290 36.120 ;
        RECT 71.525 35.920 72.290 36.060 ;
        RECT 33.790 35.860 34.110 35.920 ;
        RECT 71.525 35.875 71.815 35.920 ;
        RECT 71.970 35.860 72.290 35.920 ;
        RECT 74.270 35.860 74.590 36.120 ;
        RECT 75.205 35.875 75.495 36.105 ;
        RECT 75.650 36.060 75.970 36.120 ;
        RECT 76.125 36.060 76.415 36.105 ;
        RECT 75.650 35.920 76.415 36.060 ;
        RECT 78.500 36.060 78.640 36.215 ;
        RECT 79.790 36.200 80.110 36.260 ;
        RECT 81.185 36.215 81.475 36.260 ;
        RECT 82.105 36.215 82.395 36.445 ;
        RECT 83.025 36.215 83.315 36.445 ;
        RECT 84.850 36.400 85.170 36.460 ;
        RECT 85.325 36.400 85.615 36.445 ;
        RECT 84.850 36.260 85.615 36.400 ;
        RECT 79.330 36.060 79.650 36.120 ;
        RECT 80.250 36.060 80.570 36.120 ;
        RECT 78.500 35.920 79.650 36.060 ;
        RECT 34.250 35.720 34.570 35.780 ;
        RECT 33.420 35.580 34.570 35.720 ;
        RECT 34.250 35.520 34.570 35.580 ;
        RECT 60.945 35.720 61.235 35.765 ;
        RECT 61.390 35.720 61.710 35.780 ;
        RECT 60.945 35.580 61.710 35.720 ;
        RECT 60.945 35.535 61.235 35.580 ;
        RECT 61.390 35.520 61.710 35.580 ;
        RECT 63.705 35.720 63.995 35.765 ;
        RECT 64.150 35.720 64.470 35.780 ;
        RECT 63.705 35.580 64.470 35.720 ;
        RECT 63.705 35.535 63.995 35.580 ;
        RECT 64.150 35.520 64.470 35.580 ;
        RECT 68.290 35.520 68.610 35.780 ;
        RECT 73.825 35.720 74.115 35.765 ;
        RECT 74.730 35.720 75.050 35.780 ;
        RECT 73.825 35.580 75.050 35.720 ;
        RECT 75.280 35.720 75.420 35.875 ;
        RECT 75.650 35.860 75.970 35.920 ;
        RECT 76.125 35.875 76.415 35.920 ;
        RECT 77.490 35.720 77.810 35.780 ;
        RECT 75.280 35.580 77.810 35.720 ;
        RECT 73.825 35.535 74.115 35.580 ;
        RECT 74.730 35.520 75.050 35.580 ;
        RECT 77.490 35.520 77.810 35.580 ;
        RECT 78.410 35.720 78.730 35.780 ;
        RECT 78.960 35.720 79.100 35.920 ;
        RECT 79.330 35.860 79.650 35.920 ;
        RECT 79.880 35.920 80.570 36.060 ;
        RECT 79.880 35.765 80.020 35.920 ;
        RECT 80.250 35.860 80.570 35.920 ;
        RECT 81.630 35.860 81.950 36.120 ;
        RECT 83.100 36.060 83.240 36.215 ;
        RECT 84.850 36.200 85.170 36.260 ;
        RECT 85.325 36.215 85.615 36.260 ;
        RECT 85.770 36.200 86.090 36.460 ;
        RECT 86.230 36.200 86.550 36.460 ;
        RECT 87.150 36.200 87.470 36.460 ;
        RECT 82.180 35.920 83.240 36.060 ;
        RECT 78.410 35.580 79.100 35.720 ;
        RECT 78.410 35.520 78.730 35.580 ;
        RECT 79.805 35.535 80.095 35.765 ;
        RECT 80.710 35.720 81.030 35.780 ;
        RECT 82.180 35.720 82.320 35.920 ;
        RECT 80.710 35.580 82.320 35.720 ;
        RECT 83.010 35.720 83.330 35.780 ;
        RECT 83.945 35.720 84.235 35.765 ;
        RECT 83.010 35.580 84.235 35.720 ;
        RECT 80.710 35.520 81.030 35.580 ;
        RECT 83.010 35.520 83.330 35.580 ;
        RECT 83.945 35.535 84.235 35.580 ;
        RECT 12.100 34.900 89.840 35.380 ;
        RECT 53.570 34.700 53.890 34.760 ;
        RECT 56.805 34.700 57.095 34.745 ;
        RECT 60.470 34.700 60.790 34.760 ;
        RECT 53.570 34.560 60.790 34.700 ;
        RECT 53.570 34.500 53.890 34.560 ;
        RECT 56.805 34.515 57.095 34.560 ;
        RECT 60.470 34.500 60.790 34.560 ;
        RECT 66.450 34.700 66.770 34.760 ;
        RECT 70.130 34.700 70.450 34.760 ;
        RECT 66.450 34.560 70.450 34.700 ;
        RECT 66.450 34.500 66.770 34.560 ;
        RECT 70.130 34.500 70.450 34.560 ;
        RECT 70.605 34.700 70.895 34.745 ;
        RECT 76.585 34.700 76.875 34.745 ;
        RECT 70.605 34.560 76.875 34.700 ;
        RECT 70.605 34.515 70.895 34.560 ;
        RECT 76.585 34.515 76.875 34.560 ;
        RECT 83.470 34.700 83.790 34.760 ;
        RECT 83.470 34.560 86.920 34.700 ;
        RECT 83.470 34.500 83.790 34.560 ;
        RECT 52.650 34.360 52.970 34.420 ;
        RECT 54.030 34.360 54.350 34.420 ;
        RECT 59.565 34.360 59.855 34.405 ;
        RECT 61.850 34.360 62.170 34.420 ;
        RECT 52.650 34.220 54.350 34.360 ;
        RECT 52.650 34.160 52.970 34.220 ;
        RECT 54.030 34.160 54.350 34.220 ;
        RECT 57.340 34.220 62.170 34.360 ;
        RECT 70.220 34.360 70.360 34.500 ;
        RECT 73.350 34.360 73.670 34.420 ;
        RECT 75.650 34.360 75.970 34.420 ;
        RECT 70.220 34.220 72.200 34.360 ;
        RECT 57.340 34.065 57.480 34.220 ;
        RECT 59.565 34.175 59.855 34.220 ;
        RECT 61.850 34.160 62.170 34.220 ;
        RECT 56.345 33.835 56.635 34.065 ;
        RECT 57.265 33.835 57.555 34.065 ;
        RECT 58.645 33.835 58.935 34.065 ;
        RECT 60.485 34.020 60.775 34.065 ;
        RECT 60.930 34.020 61.250 34.080 ;
        RECT 60.485 33.880 61.250 34.020 ;
        RECT 60.485 33.835 60.775 33.880 ;
        RECT 56.420 33.680 56.560 33.835 ;
        RECT 58.720 33.680 58.860 33.835 ;
        RECT 60.930 33.820 61.250 33.880 ;
        RECT 62.325 34.020 62.615 34.065 ;
        RECT 65.070 34.020 65.390 34.080 ;
        RECT 62.325 33.880 65.390 34.020 ;
        RECT 62.325 33.835 62.615 33.880 ;
        RECT 65.070 33.820 65.390 33.880 ;
        RECT 71.050 33.820 71.370 34.080 ;
        RECT 72.060 34.020 72.200 34.220 ;
        RECT 73.350 34.220 74.960 34.360 ;
        RECT 73.350 34.160 73.670 34.220 ;
        RECT 74.820 34.065 74.960 34.220 ;
        RECT 75.650 34.220 86.460 34.360 ;
        RECT 75.650 34.160 75.970 34.220 ;
        RECT 74.285 34.020 74.575 34.065 ;
        RECT 72.060 33.880 74.575 34.020 ;
        RECT 74.285 33.835 74.575 33.880 ;
        RECT 74.745 33.835 75.035 34.065 ;
        RECT 75.205 34.020 75.495 34.065 ;
        RECT 75.205 33.880 75.880 34.020 ;
        RECT 75.205 33.835 75.495 33.880 ;
        RECT 56.420 33.540 62.540 33.680 ;
        RECT 54.030 33.340 54.350 33.400 ;
        RECT 57.725 33.340 58.015 33.385 ;
        RECT 54.030 33.200 58.015 33.340 ;
        RECT 54.030 33.140 54.350 33.200 ;
        RECT 57.725 33.155 58.015 33.200 ;
        RECT 62.400 33.060 62.540 33.540 ;
        RECT 66.910 33.480 67.230 33.740 ;
        RECT 67.370 33.480 67.690 33.740 ;
        RECT 71.510 33.480 71.830 33.740 ;
        RECT 63.245 33.340 63.535 33.385 ;
        RECT 71.050 33.340 71.370 33.400 ;
        RECT 63.245 33.200 71.370 33.340 ;
        RECT 63.245 33.155 63.535 33.200 ;
        RECT 71.050 33.140 71.370 33.200 ;
        RECT 62.310 32.800 62.630 33.060 ;
        RECT 64.625 33.000 64.915 33.045 ;
        RECT 65.070 33.000 65.390 33.060 ;
        RECT 64.625 32.860 65.390 33.000 ;
        RECT 64.625 32.815 64.915 32.860 ;
        RECT 65.070 32.800 65.390 32.860 ;
        RECT 68.750 32.800 69.070 33.060 ;
        RECT 72.905 33.000 73.195 33.045 ;
        RECT 73.350 33.000 73.670 33.060 ;
        RECT 72.905 32.860 73.670 33.000 ;
        RECT 74.360 33.000 74.500 33.835 ;
        RECT 74.730 33.340 75.050 33.400 ;
        RECT 75.740 33.340 75.880 33.880 ;
        RECT 76.110 33.820 76.430 34.080 ;
        RECT 78.410 34.020 78.730 34.080 ;
        RECT 81.645 34.020 81.935 34.065 ;
        RECT 78.410 33.880 81.935 34.020 ;
        RECT 78.410 33.820 78.730 33.880 ;
        RECT 81.645 33.835 81.935 33.880 ;
        RECT 82.090 33.820 82.410 34.080 ;
        RECT 82.550 33.820 82.870 34.080 ;
        RECT 83.470 33.820 83.790 34.080 ;
        RECT 86.320 34.065 86.460 34.220 ;
        RECT 85.325 33.835 85.615 34.065 ;
        RECT 85.785 33.835 86.075 34.065 ;
        RECT 86.245 33.835 86.535 34.065 ;
        RECT 86.780 34.020 86.920 34.560 ;
        RECT 87.150 34.020 87.470 34.080 ;
        RECT 86.780 33.880 87.470 34.020 ;
        RECT 77.490 33.680 77.810 33.740 ;
        RECT 79.345 33.680 79.635 33.725 ;
        RECT 77.490 33.540 79.635 33.680 ;
        RECT 77.490 33.480 77.810 33.540 ;
        RECT 79.345 33.495 79.635 33.540 ;
        RECT 79.790 33.680 80.110 33.740 ;
        RECT 85.400 33.680 85.540 33.835 ;
        RECT 79.790 33.540 85.540 33.680 ;
        RECT 79.790 33.480 80.110 33.540 ;
        RECT 74.730 33.200 75.880 33.340 ;
        RECT 76.110 33.340 76.430 33.400 ;
        RECT 82.090 33.340 82.410 33.400 ;
        RECT 85.860 33.340 86.000 33.835 ;
        RECT 87.150 33.820 87.470 33.880 ;
        RECT 76.110 33.200 81.860 33.340 ;
        RECT 74.730 33.140 75.050 33.200 ;
        RECT 76.110 33.140 76.430 33.200 ;
        RECT 78.410 33.000 78.730 33.060 ;
        RECT 74.360 32.860 78.730 33.000 ;
        RECT 72.905 32.815 73.195 32.860 ;
        RECT 73.350 32.800 73.670 32.860 ;
        RECT 78.410 32.800 78.730 32.860 ;
        RECT 80.250 32.800 80.570 33.060 ;
        RECT 81.720 33.000 81.860 33.200 ;
        RECT 82.090 33.200 86.000 33.340 ;
        RECT 82.090 33.140 82.410 33.200 ;
        RECT 83.470 33.000 83.790 33.060 ;
        RECT 81.720 32.860 83.790 33.000 ;
        RECT 83.470 32.800 83.790 32.860 ;
        RECT 83.930 32.800 84.250 33.060 ;
        RECT 12.100 32.180 89.840 32.660 ;
        RECT 51.270 31.980 51.590 32.040 ;
        RECT 51.745 31.980 52.035 32.025 ;
        RECT 51.270 31.840 52.035 31.980 ;
        RECT 51.270 31.780 51.590 31.840 ;
        RECT 51.745 31.795 52.035 31.840 ;
        RECT 62.310 31.780 62.630 32.040 ;
        RECT 70.130 31.980 70.450 32.040 ;
        RECT 70.605 31.980 70.895 32.025 ;
        RECT 70.130 31.840 70.895 31.980 ;
        RECT 70.130 31.780 70.450 31.840 ;
        RECT 70.605 31.795 70.895 31.840 ;
        RECT 77.045 31.980 77.335 32.025 ;
        RECT 77.950 31.980 78.270 32.040 ;
        RECT 77.045 31.840 78.270 31.980 ;
        RECT 77.045 31.795 77.335 31.840 ;
        RECT 77.950 31.780 78.270 31.840 ;
        RECT 55.910 31.640 56.200 31.685 ;
        RECT 58.010 31.640 58.300 31.685 ;
        RECT 59.580 31.640 59.870 31.685 ;
        RECT 55.910 31.500 59.870 31.640 ;
        RECT 55.910 31.455 56.200 31.500 ;
        RECT 58.010 31.455 58.300 31.500 ;
        RECT 59.580 31.455 59.870 31.500 ;
        RECT 64.190 31.640 64.480 31.685 ;
        RECT 66.290 31.640 66.580 31.685 ;
        RECT 67.860 31.640 68.150 31.685 ;
        RECT 64.190 31.500 68.150 31.640 ;
        RECT 64.190 31.455 64.480 31.500 ;
        RECT 66.290 31.455 66.580 31.500 ;
        RECT 67.860 31.455 68.150 31.500 ;
        RECT 79.790 31.640 80.080 31.685 ;
        RECT 81.360 31.640 81.650 31.685 ;
        RECT 83.460 31.640 83.750 31.685 ;
        RECT 79.790 31.500 83.750 31.640 ;
        RECT 79.790 31.455 80.080 31.500 ;
        RECT 81.360 31.455 81.650 31.500 ;
        RECT 83.460 31.455 83.750 31.500 ;
        RECT 85.770 31.440 86.090 31.700 ;
        RECT 52.190 31.300 52.510 31.360 ;
        RECT 52.665 31.300 52.955 31.345 ;
        RECT 52.190 31.160 52.955 31.300 ;
        RECT 52.190 31.100 52.510 31.160 ;
        RECT 52.665 31.115 52.955 31.160 ;
        RECT 56.305 31.300 56.595 31.345 ;
        RECT 57.495 31.300 57.785 31.345 ;
        RECT 60.015 31.300 60.305 31.345 ;
        RECT 56.305 31.160 60.305 31.300 ;
        RECT 56.305 31.115 56.595 31.160 ;
        RECT 57.495 31.115 57.785 31.160 ;
        RECT 60.015 31.115 60.305 31.160 ;
        RECT 64.585 31.300 64.875 31.345 ;
        RECT 65.775 31.300 66.065 31.345 ;
        RECT 68.295 31.300 68.585 31.345 ;
        RECT 64.585 31.160 68.585 31.300 ;
        RECT 64.585 31.115 64.875 31.160 ;
        RECT 65.775 31.115 66.065 31.160 ;
        RECT 68.295 31.115 68.585 31.160 ;
        RECT 71.050 31.300 71.370 31.360 ;
        RECT 74.285 31.300 74.575 31.345 ;
        RECT 71.050 31.160 74.575 31.300 ;
        RECT 71.050 31.100 71.370 31.160 ;
        RECT 74.285 31.115 74.575 31.160 ;
        RECT 79.355 31.300 79.645 31.345 ;
        RECT 81.875 31.300 82.165 31.345 ;
        RECT 83.065 31.300 83.355 31.345 ;
        RECT 79.355 31.160 83.355 31.300 ;
        RECT 85.860 31.300 86.000 31.440 ;
        RECT 85.860 31.160 86.460 31.300 ;
        RECT 79.355 31.115 79.645 31.160 ;
        RECT 81.875 31.115 82.165 31.160 ;
        RECT 83.065 31.115 83.355 31.160 ;
        RECT 50.810 30.960 51.130 31.020 ;
        RECT 51.285 30.960 51.575 31.005 ;
        RECT 53.110 30.960 53.430 31.020 ;
        RECT 50.810 30.820 53.430 30.960 ;
        RECT 50.810 30.760 51.130 30.820 ;
        RECT 51.285 30.775 51.575 30.820 ;
        RECT 53.110 30.760 53.430 30.820 ;
        RECT 53.570 30.760 53.890 31.020 ;
        RECT 54.030 30.760 54.350 31.020 ;
        RECT 55.425 30.960 55.715 31.005 ;
        RECT 55.870 30.960 56.190 31.020 ;
        RECT 55.425 30.820 56.190 30.960 ;
        RECT 55.425 30.775 55.715 30.820 ;
        RECT 55.870 30.760 56.190 30.820 ;
        RECT 63.690 30.760 64.010 31.020 ;
        RECT 65.070 31.005 65.390 31.020 ;
        RECT 65.040 30.960 65.390 31.005 ;
        RECT 73.825 30.960 74.115 31.005 ;
        RECT 78.410 30.960 78.730 31.020 ;
        RECT 79.790 30.960 80.110 31.020 ;
        RECT 64.875 30.820 65.390 30.960 ;
        RECT 65.040 30.775 65.390 30.820 ;
        RECT 65.070 30.760 65.390 30.775 ;
        RECT 65.620 30.820 80.110 30.960 ;
        RECT 54.965 30.620 55.255 30.665 ;
        RECT 56.650 30.620 56.940 30.665 ;
        RECT 54.965 30.480 56.940 30.620 ;
        RECT 54.965 30.435 55.255 30.480 ;
        RECT 56.650 30.435 56.940 30.480 ;
        RECT 64.610 30.620 64.930 30.680 ;
        RECT 65.620 30.620 65.760 30.820 ;
        RECT 73.825 30.775 74.115 30.820 ;
        RECT 78.410 30.760 78.730 30.820 ;
        RECT 79.790 30.760 80.110 30.820 ;
        RECT 81.170 30.960 81.490 31.020 ;
        RECT 86.320 31.005 86.460 31.160 ;
        RECT 83.945 30.960 84.235 31.005 ;
        RECT 81.170 30.820 84.235 30.960 ;
        RECT 81.170 30.760 81.490 30.820 ;
        RECT 83.945 30.775 84.235 30.820 ;
        RECT 85.785 30.775 86.075 31.005 ;
        RECT 86.245 30.775 86.535 31.005 ;
        RECT 73.365 30.620 73.655 30.665 ;
        RECT 64.610 30.480 65.760 30.620 ;
        RECT 68.610 30.480 73.655 30.620 ;
        RECT 64.610 30.420 64.930 30.480 ;
        RECT 52.665 30.280 52.955 30.325 ;
        RECT 54.490 30.280 54.810 30.340 ;
        RECT 52.665 30.140 54.810 30.280 ;
        RECT 52.665 30.095 52.955 30.140 ;
        RECT 54.490 30.080 54.810 30.140 ;
        RECT 60.470 30.280 60.790 30.340 ;
        RECT 66.910 30.280 67.230 30.340 ;
        RECT 68.610 30.280 68.750 30.480 ;
        RECT 73.365 30.435 73.655 30.480 ;
        RECT 80.250 30.620 80.570 30.680 ;
        RECT 82.610 30.620 82.900 30.665 ;
        RECT 80.250 30.480 82.900 30.620 ;
        RECT 85.860 30.620 86.000 30.775 ;
        RECT 86.690 30.760 87.010 31.020 ;
        RECT 87.150 30.960 87.470 31.020 ;
        RECT 87.625 30.960 87.915 31.005 ;
        RECT 87.150 30.820 87.915 30.960 ;
        RECT 87.150 30.760 87.470 30.820 ;
        RECT 87.625 30.775 87.915 30.820 ;
        RECT 88.070 30.620 88.390 30.680 ;
        RECT 85.860 30.480 88.390 30.620 ;
        RECT 80.250 30.420 80.570 30.480 ;
        RECT 82.610 30.435 82.900 30.480 ;
        RECT 88.070 30.420 88.390 30.480 ;
        RECT 60.470 30.140 68.750 30.280 ;
        RECT 71.050 30.280 71.370 30.340 ;
        RECT 71.525 30.280 71.815 30.325 ;
        RECT 71.050 30.140 71.815 30.280 ;
        RECT 60.470 30.080 60.790 30.140 ;
        RECT 66.910 30.080 67.230 30.140 ;
        RECT 71.050 30.080 71.370 30.140 ;
        RECT 71.525 30.095 71.815 30.140 ;
        RECT 84.390 30.080 84.710 30.340 ;
        RECT 12.100 29.460 89.840 29.940 ;
        RECT 61.390 29.260 61.710 29.320 ;
        RECT 47.680 29.120 61.710 29.260 ;
        RECT 47.680 28.965 47.820 29.120 ;
        RECT 61.390 29.060 61.710 29.120 ;
        RECT 64.610 29.060 64.930 29.320 ;
        RECT 47.605 28.735 47.895 28.965 ;
        RECT 50.810 28.920 51.130 28.980 ;
        RECT 52.665 28.920 52.955 28.965 ;
        RECT 50.810 28.780 52.955 28.920 ;
        RECT 50.810 28.720 51.130 28.780 ;
        RECT 52.665 28.735 52.955 28.780 ;
        RECT 53.110 28.720 53.430 28.980 ;
        RECT 53.815 28.920 54.105 28.965 ;
        RECT 55.410 28.920 55.730 28.980 ;
        RECT 53.815 28.780 55.730 28.920 ;
        RECT 53.815 28.735 54.105 28.780 ;
        RECT 55.410 28.720 55.730 28.780 ;
        RECT 70.300 28.920 70.590 28.965 ;
        RECT 71.050 28.920 71.370 28.980 ;
        RECT 75.650 28.920 75.970 28.980 ;
        RECT 81.170 28.920 81.490 28.980 ;
        RECT 70.300 28.780 71.370 28.920 ;
        RECT 70.300 28.735 70.590 28.780 ;
        RECT 71.050 28.720 71.370 28.780 ;
        RECT 72.980 28.780 86.920 28.920 ;
        RECT 48.525 28.580 48.815 28.625 ;
        RECT 48.985 28.580 49.275 28.625 ;
        RECT 48.525 28.440 49.275 28.580 ;
        RECT 48.525 28.395 48.815 28.440 ;
        RECT 48.985 28.395 49.275 28.440 ;
        RECT 49.905 28.580 50.195 28.625 ;
        RECT 49.905 28.440 51.960 28.580 ;
        RECT 49.905 28.395 50.195 28.440 ;
        RECT 50.825 28.055 51.115 28.285 ;
        RECT 51.820 28.240 51.960 28.440 ;
        RECT 52.190 28.380 52.510 28.640 ;
        RECT 54.490 28.380 54.810 28.640 ;
        RECT 57.220 28.580 57.510 28.625 ;
        RECT 58.630 28.580 58.950 28.640 ;
        RECT 57.220 28.440 58.950 28.580 ;
        RECT 57.220 28.395 57.510 28.440 ;
        RECT 58.630 28.380 58.950 28.440 ;
        RECT 71.525 28.580 71.815 28.625 ;
        RECT 71.985 28.580 72.275 28.625 ;
        RECT 72.980 28.580 73.120 28.780 ;
        RECT 75.650 28.720 75.970 28.780 ;
        RECT 81.170 28.720 81.490 28.780 ;
        RECT 73.350 28.625 73.670 28.640 ;
        RECT 71.525 28.440 73.120 28.580 ;
        RECT 73.320 28.580 73.670 28.625 ;
        RECT 83.930 28.580 84.250 28.640 ;
        RECT 86.780 28.625 86.920 28.780 ;
        RECT 85.370 28.580 85.660 28.625 ;
        RECT 73.320 28.440 73.820 28.580 ;
        RECT 83.930 28.440 85.660 28.580 ;
        RECT 71.525 28.395 71.815 28.440 ;
        RECT 71.985 28.395 72.275 28.440 ;
        RECT 73.320 28.395 73.670 28.440 ;
        RECT 73.350 28.380 73.670 28.395 ;
        RECT 83.930 28.380 84.250 28.440 ;
        RECT 85.370 28.395 85.660 28.440 ;
        RECT 86.705 28.395 86.995 28.625 ;
        RECT 53.570 28.240 53.890 28.300 ;
        RECT 51.820 28.100 53.890 28.240 ;
        RECT 50.900 27.900 51.040 28.055 ;
        RECT 53.570 28.040 53.890 28.100 ;
        RECT 55.870 28.040 56.190 28.300 ;
        RECT 56.765 28.240 57.055 28.285 ;
        RECT 57.955 28.240 58.245 28.285 ;
        RECT 60.475 28.240 60.765 28.285 ;
        RECT 56.765 28.100 60.765 28.240 ;
        RECT 56.765 28.055 57.055 28.100 ;
        RECT 57.955 28.055 58.245 28.100 ;
        RECT 60.475 28.055 60.765 28.100 ;
        RECT 66.935 28.240 67.225 28.285 ;
        RECT 69.455 28.240 69.745 28.285 ;
        RECT 70.645 28.240 70.935 28.285 ;
        RECT 66.935 28.100 70.935 28.240 ;
        RECT 66.935 28.055 67.225 28.100 ;
        RECT 69.455 28.055 69.745 28.100 ;
        RECT 70.645 28.055 70.935 28.100 ;
        RECT 72.865 28.240 73.155 28.285 ;
        RECT 74.055 28.240 74.345 28.285 ;
        RECT 76.575 28.240 76.865 28.285 ;
        RECT 72.865 28.100 76.865 28.240 ;
        RECT 72.865 28.055 73.155 28.100 ;
        RECT 74.055 28.055 74.345 28.100 ;
        RECT 76.575 28.055 76.865 28.100 ;
        RECT 82.115 28.240 82.405 28.285 ;
        RECT 84.635 28.240 84.925 28.285 ;
        RECT 85.825 28.240 86.115 28.285 ;
        RECT 82.115 28.100 86.115 28.240 ;
        RECT 82.115 28.055 82.405 28.100 ;
        RECT 84.635 28.055 84.925 28.100 ;
        RECT 85.825 28.055 86.115 28.100 ;
        RECT 56.370 27.900 56.660 27.945 ;
        RECT 58.470 27.900 58.760 27.945 ;
        RECT 60.040 27.900 60.330 27.945 ;
        RECT 50.900 27.760 56.100 27.900 ;
        RECT 46.670 27.360 46.990 27.620 ;
        RECT 51.270 27.360 51.590 27.620 ;
        RECT 55.960 27.560 56.100 27.760 ;
        RECT 56.370 27.760 60.330 27.900 ;
        RECT 56.370 27.715 56.660 27.760 ;
        RECT 58.470 27.715 58.760 27.760 ;
        RECT 60.040 27.715 60.330 27.760 ;
        RECT 62.770 27.700 63.090 27.960 ;
        RECT 67.370 27.900 67.660 27.945 ;
        RECT 68.940 27.900 69.230 27.945 ;
        RECT 71.040 27.900 71.330 27.945 ;
        RECT 67.370 27.760 71.330 27.900 ;
        RECT 67.370 27.715 67.660 27.760 ;
        RECT 68.940 27.715 69.230 27.760 ;
        RECT 71.040 27.715 71.330 27.760 ;
        RECT 72.470 27.900 72.760 27.945 ;
        RECT 74.570 27.900 74.860 27.945 ;
        RECT 76.140 27.900 76.430 27.945 ;
        RECT 72.470 27.760 76.430 27.900 ;
        RECT 72.470 27.715 72.760 27.760 ;
        RECT 74.570 27.715 74.860 27.760 ;
        RECT 76.140 27.715 76.430 27.760 ;
        RECT 79.805 27.900 80.095 27.945 ;
        RECT 81.630 27.900 81.950 27.960 ;
        RECT 79.805 27.760 81.950 27.900 ;
        RECT 79.805 27.715 80.095 27.760 ;
        RECT 81.630 27.700 81.950 27.760 ;
        RECT 82.550 27.900 82.840 27.945 ;
        RECT 84.120 27.900 84.410 27.945 ;
        RECT 86.220 27.900 86.510 27.945 ;
        RECT 82.550 27.760 86.510 27.900 ;
        RECT 82.550 27.715 82.840 27.760 ;
        RECT 84.120 27.715 84.410 27.760 ;
        RECT 86.220 27.715 86.510 27.760 ;
        RECT 60.930 27.560 61.250 27.620 ;
        RECT 55.960 27.420 61.250 27.560 ;
        RECT 60.930 27.360 61.250 27.420 ;
        RECT 78.870 27.360 79.190 27.620 ;
        RECT 12.100 26.740 89.840 27.220 ;
        RECT 55.410 26.340 55.730 26.600 ;
        RECT 60.930 26.540 61.250 26.600 ;
        RECT 62.785 26.540 63.075 26.585 ;
        RECT 64.165 26.540 64.455 26.585 ;
        RECT 60.930 26.400 64.455 26.540 ;
        RECT 60.930 26.340 61.250 26.400 ;
        RECT 62.785 26.355 63.075 26.400 ;
        RECT 64.165 26.355 64.455 26.400 ;
        RECT 65.085 26.540 65.375 26.585 ;
        RECT 67.370 26.540 67.690 26.600 ;
        RECT 65.085 26.400 67.690 26.540 ;
        RECT 65.085 26.355 65.375 26.400 ;
        RECT 67.370 26.340 67.690 26.400 ;
        RECT 73.365 26.540 73.655 26.585 ;
        RECT 77.490 26.540 77.810 26.600 ;
        RECT 84.850 26.540 85.170 26.600 ;
        RECT 88.085 26.540 88.375 26.585 ;
        RECT 73.365 26.400 77.810 26.540 ;
        RECT 73.365 26.355 73.655 26.400 ;
        RECT 77.490 26.340 77.810 26.400 ;
        RECT 78.040 26.400 80.020 26.540 ;
        RECT 56.370 26.200 56.660 26.245 ;
        RECT 58.470 26.200 58.760 26.245 ;
        RECT 60.040 26.200 60.330 26.245 ;
        RECT 56.370 26.060 60.330 26.200 ;
        RECT 56.370 26.015 56.660 26.060 ;
        RECT 58.470 26.015 58.760 26.060 ;
        RECT 60.040 26.015 60.330 26.060 ;
        RECT 66.950 26.200 67.240 26.245 ;
        RECT 69.050 26.200 69.340 26.245 ;
        RECT 70.620 26.200 70.910 26.245 ;
        RECT 76.110 26.200 76.430 26.260 ;
        RECT 78.040 26.200 78.180 26.400 ;
        RECT 66.950 26.060 70.910 26.200 ;
        RECT 66.950 26.015 67.240 26.060 ;
        RECT 69.050 26.015 69.340 26.060 ;
        RECT 70.620 26.015 70.910 26.060 ;
        RECT 71.600 26.060 78.180 26.200 ;
        RECT 78.500 26.060 79.560 26.200 ;
        RECT 46.670 25.860 46.990 25.920 ;
        RECT 46.670 25.720 53.340 25.860 ;
        RECT 46.670 25.660 46.990 25.720 ;
        RECT 50.350 25.320 50.670 25.580 ;
        RECT 52.650 25.320 52.970 25.580 ;
        RECT 53.200 25.520 53.340 25.720 ;
        RECT 55.870 25.660 56.190 25.920 ;
        RECT 56.765 25.860 57.055 25.905 ;
        RECT 57.955 25.860 58.245 25.905 ;
        RECT 60.475 25.860 60.765 25.905 ;
        RECT 56.765 25.720 60.765 25.860 ;
        RECT 56.765 25.675 57.055 25.720 ;
        RECT 57.955 25.675 58.245 25.720 ;
        RECT 60.475 25.675 60.765 25.720 ;
        RECT 63.690 25.860 64.010 25.920 ;
        RECT 66.450 25.860 66.770 25.920 ;
        RECT 63.690 25.720 66.770 25.860 ;
        RECT 63.690 25.660 64.010 25.720 ;
        RECT 66.450 25.660 66.770 25.720 ;
        RECT 67.345 25.860 67.635 25.905 ;
        RECT 68.535 25.860 68.825 25.905 ;
        RECT 71.055 25.860 71.345 25.905 ;
        RECT 67.345 25.720 71.345 25.860 ;
        RECT 67.345 25.675 67.635 25.720 ;
        RECT 68.535 25.675 68.825 25.720 ;
        RECT 71.055 25.675 71.345 25.720 ;
        RECT 57.165 25.520 57.455 25.565 ;
        RECT 71.600 25.520 71.740 26.060 ;
        RECT 76.110 26.000 76.430 26.060 ;
        RECT 75.665 25.860 75.955 25.905 ;
        RECT 78.500 25.860 78.640 26.060 ;
        RECT 75.665 25.720 78.640 25.860 ;
        RECT 75.665 25.675 75.955 25.720 ;
        RECT 53.200 25.380 57.455 25.520 ;
        RECT 57.165 25.335 57.455 25.380 ;
        RECT 61.940 25.380 71.740 25.520 ;
        RECT 71.970 25.520 72.290 25.580 ;
        RECT 73.825 25.520 74.115 25.565 ;
        RECT 77.950 25.520 78.270 25.580 ;
        RECT 71.970 25.380 78.270 25.520 ;
        RECT 52.190 25.180 52.510 25.240 ;
        RECT 61.940 25.180 62.080 25.380 ;
        RECT 71.970 25.320 72.290 25.380 ;
        RECT 73.825 25.335 74.115 25.380 ;
        RECT 77.950 25.320 78.270 25.380 ;
        RECT 78.410 25.320 78.730 25.580 ;
        RECT 79.420 25.565 79.560 26.060 ;
        RECT 78.885 25.335 79.175 25.565 ;
        RECT 79.345 25.335 79.635 25.565 ;
        RECT 79.880 25.520 80.020 26.400 ;
        RECT 84.850 26.400 88.375 26.540 ;
        RECT 84.850 26.340 85.170 26.400 ;
        RECT 88.085 26.355 88.375 26.400 ;
        RECT 81.670 26.200 81.960 26.245 ;
        RECT 83.770 26.200 84.060 26.245 ;
        RECT 85.340 26.200 85.630 26.245 ;
        RECT 81.670 26.060 85.630 26.200 ;
        RECT 81.670 26.015 81.960 26.060 ;
        RECT 83.770 26.015 84.060 26.060 ;
        RECT 85.340 26.015 85.630 26.060 ;
        RECT 81.170 25.660 81.490 25.920 ;
        RECT 82.065 25.860 82.355 25.905 ;
        RECT 83.255 25.860 83.545 25.905 ;
        RECT 85.775 25.860 86.065 25.905 ;
        RECT 82.065 25.720 86.065 25.860 ;
        RECT 82.065 25.675 82.355 25.720 ;
        RECT 83.255 25.675 83.545 25.720 ;
        RECT 85.775 25.675 86.065 25.720 ;
        RECT 80.265 25.520 80.555 25.565 ;
        RECT 79.880 25.380 80.555 25.520 ;
        RECT 80.265 25.335 80.555 25.380 ;
        RECT 82.520 25.520 82.810 25.565 ;
        RECT 84.390 25.520 84.710 25.580 ;
        RECT 82.520 25.380 84.710 25.520 ;
        RECT 82.520 25.335 82.810 25.380 ;
        RECT 52.190 25.040 62.080 25.180 ;
        RECT 62.310 25.180 62.630 25.240 ;
        RECT 64.150 25.225 64.470 25.240 ;
        RECT 63.245 25.180 63.535 25.225 ;
        RECT 62.310 25.040 63.535 25.180 ;
        RECT 52.190 24.980 52.510 25.040 ;
        RECT 62.310 24.980 62.630 25.040 ;
        RECT 63.245 24.995 63.535 25.040 ;
        RECT 64.150 24.995 64.535 25.225 ;
        RECT 67.800 25.180 68.090 25.225 ;
        RECT 68.750 25.180 69.070 25.240 ;
        RECT 67.800 25.040 69.070 25.180 ;
        RECT 67.800 24.995 68.090 25.040 ;
        RECT 64.150 24.980 64.470 24.995 ;
        RECT 68.750 24.980 69.070 25.040 ;
        RECT 74.745 25.180 75.035 25.225 ;
        RECT 76.110 25.180 76.430 25.240 ;
        RECT 74.745 25.040 76.430 25.180 ;
        RECT 78.960 25.180 79.100 25.335 ;
        RECT 84.390 25.320 84.710 25.380 ;
        RECT 85.770 25.180 86.090 25.240 ;
        RECT 78.960 25.040 86.090 25.180 ;
        RECT 74.745 24.995 75.035 25.040 ;
        RECT 76.110 24.980 76.430 25.040 ;
        RECT 85.770 24.980 86.090 25.040 ;
        RECT 49.445 24.840 49.735 24.885 ;
        RECT 50.350 24.840 50.670 24.900 ;
        RECT 49.445 24.700 50.670 24.840 ;
        RECT 49.445 24.655 49.735 24.700 ;
        RECT 50.350 24.640 50.670 24.700 ;
        RECT 77.030 24.640 77.350 24.900 ;
        RECT 12.100 24.020 89.840 24.500 ;
        RECT 52.650 23.820 52.970 23.880 ;
        RECT 53.585 23.820 53.875 23.865 ;
        RECT 52.650 23.680 53.875 23.820 ;
        RECT 52.650 23.620 52.970 23.680 ;
        RECT 53.585 23.635 53.875 23.680 ;
        RECT 58.630 23.620 58.950 23.880 ;
        RECT 60.485 23.820 60.775 23.865 ;
        RECT 62.770 23.820 63.090 23.880 ;
        RECT 60.485 23.680 63.090 23.820 ;
        RECT 60.485 23.635 60.775 23.680 ;
        RECT 62.770 23.620 63.090 23.680 ;
        RECT 76.110 23.820 76.430 23.880 ;
        RECT 77.045 23.820 77.335 23.865 ;
        RECT 79.330 23.820 79.650 23.880 ;
        RECT 76.110 23.680 79.650 23.820 ;
        RECT 76.110 23.620 76.430 23.680 ;
        RECT 77.045 23.635 77.335 23.680 ;
        RECT 79.330 23.620 79.650 23.680 ;
        RECT 80.725 23.820 81.015 23.865 ;
        RECT 86.230 23.820 86.550 23.880 ;
        RECT 80.725 23.680 86.550 23.820 ;
        RECT 80.725 23.635 81.015 23.680 ;
        RECT 86.230 23.620 86.550 23.680 ;
        RECT 48.020 23.480 48.310 23.525 ;
        RECT 51.270 23.480 51.590 23.540 ;
        RECT 48.020 23.340 51.590 23.480 ;
        RECT 48.020 23.295 48.310 23.340 ;
        RECT 51.270 23.280 51.590 23.340 ;
        RECT 66.450 23.480 66.770 23.540 ;
        RECT 75.650 23.480 75.970 23.540 ;
        RECT 66.450 23.340 75.970 23.480 ;
        RECT 66.450 23.280 66.770 23.340 ;
        RECT 34.250 23.140 34.570 23.200 ;
        RECT 70.220 23.185 70.360 23.340 ;
        RECT 75.650 23.280 75.970 23.340 ;
        RECT 79.805 23.480 80.095 23.525 ;
        RECT 80.250 23.480 80.570 23.540 ;
        RECT 79.805 23.340 80.570 23.480 ;
        RECT 79.805 23.295 80.095 23.340 ;
        RECT 80.250 23.280 80.570 23.340 ;
        RECT 82.520 23.480 82.810 23.525 ;
        RECT 83.010 23.480 83.330 23.540 ;
        RECT 82.520 23.340 83.330 23.480 ;
        RECT 82.520 23.295 82.810 23.340 ;
        RECT 83.010 23.280 83.330 23.340 ;
        RECT 46.685 23.140 46.975 23.185 ;
        RECT 34.250 23.000 46.975 23.140 ;
        RECT 34.250 22.940 34.570 23.000 ;
        RECT 46.685 22.955 46.975 23.000 ;
        RECT 70.145 23.140 70.435 23.185 ;
        RECT 71.480 23.140 71.770 23.185 ;
        RECT 77.030 23.140 77.350 23.200 ;
        RECT 70.145 23.000 70.545 23.140 ;
        RECT 71.480 23.000 77.350 23.140 ;
        RECT 70.145 22.955 70.435 23.000 ;
        RECT 71.480 22.955 71.770 23.000 ;
        RECT 77.030 22.940 77.350 23.000 ;
        RECT 77.490 22.940 77.810 23.200 ;
        RECT 77.950 23.140 78.270 23.200 ;
        RECT 78.885 23.140 79.175 23.185 ;
        RECT 79.330 23.140 79.650 23.200 ;
        RECT 77.950 23.000 79.650 23.140 ;
        RECT 77.950 22.940 78.270 23.000 ;
        RECT 78.885 22.955 79.175 23.000 ;
        RECT 79.330 22.940 79.650 23.000 ;
        RECT 81.170 22.940 81.490 23.200 ;
        RECT 47.565 22.800 47.855 22.845 ;
        RECT 48.755 22.800 49.045 22.845 ;
        RECT 51.275 22.800 51.565 22.845 ;
        RECT 47.565 22.660 51.565 22.800 ;
        RECT 47.565 22.615 47.855 22.660 ;
        RECT 48.755 22.615 49.045 22.660 ;
        RECT 51.275 22.615 51.565 22.660 ;
        RECT 60.930 22.600 61.250 22.860 ;
        RECT 61.390 22.600 61.710 22.860 ;
        RECT 71.025 22.800 71.315 22.845 ;
        RECT 72.215 22.800 72.505 22.845 ;
        RECT 74.735 22.800 75.025 22.845 ;
        RECT 71.025 22.660 75.025 22.800 ;
        RECT 71.025 22.615 71.315 22.660 ;
        RECT 72.215 22.615 72.505 22.660 ;
        RECT 74.735 22.615 75.025 22.660 ;
        RECT 82.065 22.800 82.355 22.845 ;
        RECT 83.255 22.800 83.545 22.845 ;
        RECT 85.775 22.800 86.065 22.845 ;
        RECT 82.065 22.660 86.065 22.800 ;
        RECT 82.065 22.615 82.355 22.660 ;
        RECT 83.255 22.615 83.545 22.660 ;
        RECT 85.775 22.615 86.065 22.660 ;
        RECT 47.170 22.460 47.460 22.505 ;
        RECT 49.270 22.460 49.560 22.505 ;
        RECT 50.840 22.460 51.130 22.505 ;
        RECT 47.170 22.320 51.130 22.460 ;
        RECT 47.170 22.275 47.460 22.320 ;
        RECT 49.270 22.275 49.560 22.320 ;
        RECT 50.840 22.275 51.130 22.320 ;
        RECT 70.630 22.460 70.920 22.505 ;
        RECT 72.730 22.460 73.020 22.505 ;
        RECT 74.300 22.460 74.590 22.505 ;
        RECT 70.630 22.320 74.590 22.460 ;
        RECT 70.630 22.275 70.920 22.320 ;
        RECT 72.730 22.275 73.020 22.320 ;
        RECT 74.300 22.275 74.590 22.320 ;
        RECT 75.650 22.460 75.970 22.520 ;
        RECT 78.870 22.460 79.190 22.520 ;
        RECT 75.650 22.320 79.190 22.460 ;
        RECT 75.650 22.260 75.970 22.320 ;
        RECT 78.870 22.260 79.190 22.320 ;
        RECT 81.670 22.460 81.960 22.505 ;
        RECT 83.770 22.460 84.060 22.505 ;
        RECT 85.340 22.460 85.630 22.505 ;
        RECT 81.670 22.320 85.630 22.460 ;
        RECT 81.670 22.275 81.960 22.320 ;
        RECT 83.770 22.275 84.060 22.320 ;
        RECT 85.340 22.275 85.630 22.320 ;
        RECT 78.425 22.120 78.715 22.165 ;
        RECT 79.790 22.120 80.110 22.180 ;
        RECT 78.425 21.980 80.110 22.120 ;
        RECT 78.425 21.935 78.715 21.980 ;
        RECT 79.790 21.920 80.110 21.980 ;
        RECT 80.250 22.120 80.570 22.180 ;
        RECT 88.085 22.120 88.375 22.165 ;
        RECT 80.250 21.980 88.375 22.120 ;
        RECT 80.250 21.920 80.570 21.980 ;
        RECT 88.085 21.935 88.375 21.980 ;
        RECT 12.100 21.300 89.840 21.780 ;
        RECT 80.710 20.900 81.030 21.160 ;
        RECT 82.550 20.900 82.870 21.160 ;
        RECT 85.325 21.100 85.615 21.145 ;
        RECT 86.690 21.100 87.010 21.160 ;
        RECT 85.325 20.960 87.010 21.100 ;
        RECT 85.325 20.915 85.615 20.960 ;
        RECT 86.690 20.900 87.010 20.960 ;
        RECT 87.610 20.900 87.930 21.160 ;
        RECT 48.525 20.760 48.815 20.805 ;
        RECT 50.810 20.760 51.130 20.820 ;
        RECT 48.525 20.620 51.130 20.760 ;
        RECT 48.525 20.575 48.815 20.620 ;
        RECT 50.810 20.560 51.130 20.620 ;
        RECT 56.805 20.760 57.095 20.805 ;
        RECT 60.930 20.760 61.250 20.820 ;
        RECT 56.805 20.620 61.250 20.760 ;
        RECT 56.805 20.575 57.095 20.620 ;
        RECT 60.930 20.560 61.250 20.620 ;
        RECT 79.330 20.760 79.650 20.820 ;
        RECT 79.330 20.620 83.700 20.760 ;
        RECT 79.330 20.560 79.650 20.620 ;
        RECT 43.925 20.420 44.215 20.465 ;
        RECT 53.110 20.420 53.430 20.480 ;
        RECT 43.925 20.280 53.430 20.420 ;
        RECT 43.925 20.235 44.215 20.280 ;
        RECT 53.110 20.220 53.430 20.280 ;
        RECT 42.070 20.080 42.390 20.140 ;
        RECT 42.545 20.080 42.835 20.125 ;
        RECT 42.070 19.940 42.835 20.080 ;
        RECT 42.070 19.880 42.390 19.940 ;
        RECT 42.545 19.895 42.835 19.940 ;
        RECT 50.350 19.880 50.670 20.140 ;
        RECT 52.650 20.080 52.970 20.140 ;
        RECT 53.585 20.080 53.875 20.125 ;
        RECT 52.650 19.940 53.875 20.080 ;
        RECT 52.650 19.880 52.970 19.940 ;
        RECT 53.585 19.895 53.875 19.940 ;
        RECT 72.905 20.080 73.195 20.125 ;
        RECT 75.650 20.080 75.970 20.140 ;
        RECT 72.905 19.940 75.970 20.080 ;
        RECT 72.905 19.895 73.195 19.940 ;
        RECT 75.650 19.880 75.970 19.940 ;
        RECT 76.110 19.880 76.430 20.140 ;
        RECT 76.570 20.080 76.890 20.140 ;
        RECT 79.345 20.080 79.635 20.125 ;
        RECT 76.570 19.940 79.635 20.080 ;
        RECT 76.570 19.880 76.890 19.940 ;
        RECT 79.345 19.895 79.635 19.940 ;
        RECT 79.790 19.880 80.110 20.140 ;
        RECT 80.250 20.080 80.570 20.140 ;
        RECT 83.560 20.125 83.700 20.620 ;
        RECT 81.645 20.080 81.935 20.125 ;
        RECT 80.250 19.940 81.935 20.080 ;
        RECT 80.250 19.880 80.570 19.940 ;
        RECT 81.645 19.895 81.935 19.940 ;
        RECT 83.485 19.895 83.775 20.125 ;
        RECT 84.405 20.080 84.695 20.125 ;
        RECT 84.850 20.080 85.170 20.140 ;
        RECT 86.705 20.080 86.995 20.125 ;
        RECT 84.405 19.940 86.995 20.080 ;
        RECT 84.405 19.895 84.695 19.940 ;
        RECT 84.850 19.880 85.170 19.940 ;
        RECT 86.705 19.895 86.995 19.940 ;
        RECT 45.290 19.740 45.610 19.800 ;
        RECT 47.605 19.740 47.895 19.785 ;
        RECT 45.290 19.600 47.895 19.740 ;
        RECT 45.290 19.540 45.610 19.600 ;
        RECT 47.605 19.555 47.895 19.600 ;
        RECT 54.950 19.740 55.270 19.800 ;
        RECT 55.885 19.740 56.175 19.785 ;
        RECT 54.950 19.600 56.175 19.740 ;
        RECT 54.950 19.540 55.270 19.600 ;
        RECT 55.885 19.555 56.175 19.600 ;
        RECT 48.510 19.400 48.830 19.460 ;
        RECT 49.445 19.400 49.735 19.445 ;
        RECT 48.510 19.260 49.735 19.400 ;
        RECT 48.510 19.200 48.830 19.260 ;
        RECT 49.445 19.215 49.735 19.260 ;
        RECT 51.730 19.400 52.050 19.460 ;
        RECT 52.665 19.400 52.955 19.445 ;
        RECT 51.730 19.260 52.955 19.400 ;
        RECT 51.730 19.200 52.050 19.260 ;
        RECT 52.665 19.215 52.955 19.260 ;
        RECT 71.050 19.400 71.370 19.460 ;
        RECT 71.985 19.400 72.275 19.445 ;
        RECT 71.050 19.260 72.275 19.400 ;
        RECT 71.050 19.200 71.370 19.260 ;
        RECT 71.985 19.215 72.275 19.260 ;
        RECT 74.270 19.400 74.590 19.460 ;
        RECT 75.205 19.400 75.495 19.445 ;
        RECT 74.270 19.260 75.495 19.400 ;
        RECT 74.270 19.200 74.590 19.260 ;
        RECT 75.205 19.215 75.495 19.260 ;
        RECT 77.490 19.400 77.810 19.460 ;
        RECT 78.425 19.400 78.715 19.445 ;
        RECT 77.490 19.260 78.715 19.400 ;
        RECT 77.490 19.200 77.810 19.260 ;
        RECT 78.425 19.215 78.715 19.260 ;
        RECT 12.100 18.580 89.840 19.060 ;
      LAYER met2 ;
        RECT 118.795 224.565 119.455 225.215 ;
        RECT 121.530 224.805 122.190 225.455 ;
        RECT 124.275 224.945 124.935 225.595 ;
        RECT 127.145 224.965 127.805 225.615 ;
        RECT 129.605 224.960 130.265 225.610 ;
        RECT 132.985 224.945 133.645 225.595 ;
        RECT 134.915 225.075 135.575 225.725 ;
        RECT 137.630 224.895 138.410 225.575 ;
        RECT 69.205 222.560 69.595 222.640 ;
        RECT 69.205 222.420 127.660 222.560 ;
        RECT 69.205 222.340 69.595 222.420 ;
        RECT 72.120 222.090 72.420 222.215 ;
        RECT 72.120 221.950 126.920 222.090 ;
        RECT 72.120 221.825 72.420 221.950 ;
        RECT 74.770 221.725 75.160 221.785 ;
        RECT 125.240 221.770 125.770 221.780 ;
        RECT 125.240 221.725 125.805 221.770 ;
        RECT 74.770 221.540 125.805 221.725 ;
        RECT 74.770 221.485 75.160 221.540 ;
        RECT 125.240 221.490 125.805 221.540 ;
        RECT 126.780 221.620 126.920 221.950 ;
        RECT 127.520 222.060 127.660 222.420 ;
        RECT 149.680 222.060 150.000 222.120 ;
        RECT 127.520 221.920 150.000 222.060 ;
        RECT 149.680 221.860 150.000 221.920 ;
        RECT 125.240 221.480 125.770 221.490 ;
        RECT 126.780 221.480 140.200 221.620 ;
        RECT 138.880 221.310 139.370 221.320 ;
        RECT 80.275 221.240 80.665 221.305 ;
        RECT 82.770 221.240 83.840 221.280 ;
        RECT 80.275 221.160 117.550 221.240 ;
        RECT 138.880 221.160 139.405 221.310 ;
        RECT 80.275 221.120 139.405 221.160 ;
        RECT 80.275 221.070 82.940 221.120 ;
        RECT 83.620 221.070 139.405 221.120 ;
        RECT 80.275 221.005 80.665 221.070 ;
        RECT 117.055 221.030 139.405 221.070 ;
        RECT 117.055 221.020 139.370 221.030 ;
        RECT 83.085 220.900 83.475 220.980 ;
        RECT 117.055 220.965 139.130 221.020 ;
        RECT 140.060 221.000 140.200 221.480 ;
        RECT 149.120 221.000 149.440 221.060 ;
        RECT 83.085 220.800 116.760 220.900 ;
        RECT 140.060 220.860 149.440 221.000 ;
        RECT 149.120 220.800 149.440 220.860 ;
        RECT 83.085 220.760 133.370 220.800 ;
        RECT 83.085 220.680 83.475 220.760 ;
        RECT 116.620 220.660 133.370 220.760 ;
        RECT 85.785 220.525 86.175 220.595 ;
        RECT 115.915 220.580 116.285 220.585 ;
        RECT 115.570 220.525 116.285 220.580 ;
        RECT 85.785 220.365 116.285 220.525 ;
        RECT 85.785 220.295 86.175 220.365 ;
        RECT 115.570 220.310 116.285 220.365 ;
        RECT 115.915 220.305 116.285 220.310 ;
        RECT 91.280 220.140 91.670 220.220 ;
        RECT 132.220 220.210 132.610 220.480 ;
        RECT 93.670 220.140 94.650 220.160 ;
        RECT 116.845 220.140 132.610 220.210 ;
        RECT 91.280 220.040 132.610 220.140 ;
        RECT 133.230 220.250 133.370 220.660 ;
        RECT 148.660 220.250 148.920 220.340 ;
        RECT 133.230 220.110 148.920 220.250 ;
        RECT 91.280 220.035 132.510 220.040 ;
        RECT 91.280 220.020 117.005 220.035 ;
        RECT 148.660 220.020 148.920 220.110 ;
        RECT 91.280 219.995 93.810 220.020 ;
        RECT 94.490 220.000 117.005 220.020 ;
        RECT 94.490 219.995 116.860 220.000 ;
        RECT 91.280 219.920 91.670 219.995 ;
        RECT 93.955 219.800 94.345 219.880 ;
        RECT 148.110 219.800 148.430 219.860 ;
        RECT 93.955 219.660 148.430 219.800 ;
        RECT 88.600 219.490 88.900 219.615 ;
        RECT 93.955 219.580 94.345 219.660 ;
        RECT 148.110 219.600 148.430 219.660 ;
        RECT 88.600 219.440 93.810 219.490 ;
        RECT 94.490 219.440 111.950 219.490 ;
        RECT 88.600 219.350 111.950 219.440 ;
        RECT 88.600 219.225 88.900 219.350 ;
        RECT 93.560 219.310 94.730 219.350 ;
        RECT 93.670 219.290 94.610 219.310 ;
        RECT 77.535 219.090 77.925 219.170 ;
        RECT 96.090 219.090 111.560 219.180 ;
        RECT 77.535 219.080 88.440 219.090 ;
        RECT 89.070 219.080 111.560 219.090 ;
        RECT 77.535 219.040 111.560 219.080 ;
        RECT 77.535 218.950 96.230 219.040 ;
        RECT 77.535 218.870 77.925 218.950 ;
        RECT 88.330 218.940 89.190 218.950 ;
        RECT 66.485 218.730 66.875 218.810 ;
        RECT 96.750 218.730 111.150 218.830 ;
        RECT 66.485 218.690 111.150 218.730 ;
        RECT 66.485 218.590 96.890 218.690 ;
        RECT 66.485 218.510 66.875 218.590 ;
        RECT 63.655 218.200 64.045 218.280 ;
        RECT 63.655 218.060 110.150 218.200 ;
        RECT 63.655 217.980 64.045 218.060 ;
        RECT 95.395 217.375 95.655 217.695 ;
        RECT 45.310 181.510 45.590 185.510 ;
        RECT 71.070 181.510 71.350 185.510 ;
        RECT 74.290 181.510 74.570 185.510 ;
        RECT 80.730 181.510 81.010 185.510 ;
        RECT 83.950 181.510 84.230 185.510 ;
        RECT 27.650 173.675 29.190 174.045 ;
        RECT 45.380 173.510 45.520 181.510 ;
        RECT 71.140 173.510 71.280 181.510 ;
        RECT 45.320 173.190 45.580 173.510 ;
        RECT 71.080 173.190 71.340 173.510 ;
        RECT 71.540 173.190 71.800 173.510 ;
        RECT 47.160 172.170 47.420 172.490 ;
        RECT 59.580 172.170 59.840 172.490 ;
        RECT 60.960 172.170 61.220 172.490 ;
        RECT 63.260 172.170 63.520 172.490 ;
        RECT 64.180 172.170 64.440 172.490 ;
        RECT 30.950 170.955 32.490 171.325 ;
        RECT 42.560 169.790 42.820 170.110 ;
        RECT 43.480 169.790 43.740 170.110 ;
        RECT 43.940 169.790 44.200 170.110 ;
        RECT 41.640 169.110 41.900 169.430 ;
        RECT 42.100 169.110 42.360 169.430 ;
        RECT 40.260 168.770 40.520 169.090 ;
        RECT 27.650 168.235 29.190 168.605 ;
        RECT 40.320 166.710 40.460 168.770 ;
        RECT 41.700 167.585 41.840 169.110 ;
        RECT 41.630 167.215 41.910 167.585 ;
        RECT 40.260 166.390 40.520 166.710 ;
        RECT 41.180 166.390 41.440 166.710 ;
        RECT 30.950 165.515 32.490 165.885 ;
        RECT 37.040 164.010 37.300 164.330 ;
        RECT 27.650 162.795 29.190 163.165 ;
        RECT 37.100 162.630 37.240 164.010 ;
        RECT 41.240 163.990 41.380 166.390 ;
        RECT 42.160 164.670 42.300 169.110 ;
        RECT 42.620 166.905 42.760 169.790 ;
        RECT 42.550 166.535 42.830 166.905 ;
        RECT 43.540 165.350 43.680 169.790 ;
        RECT 43.480 165.030 43.740 165.350 ;
        RECT 42.100 164.350 42.360 164.670 ;
        RECT 41.180 163.670 41.440 163.990 ;
        RECT 40.260 163.330 40.520 163.650 ;
        RECT 37.040 162.310 37.300 162.630 ;
        RECT 30.950 160.075 32.490 160.445 ;
        RECT 36.120 158.910 36.380 159.230 ;
        RECT 7.130 158.375 7.410 158.745 ;
        RECT 7.200 96.670 7.340 158.375 ;
        RECT 34.280 157.890 34.540 158.210 ;
        RECT 27.650 157.355 29.190 157.725 ;
        RECT 30.950 154.635 32.490 155.005 ;
        RECT 34.340 153.790 34.480 157.890 ;
        RECT 35.200 155.170 35.460 155.490 ;
        RECT 34.280 153.470 34.540 153.790 ;
        RECT 27.650 151.915 29.190 152.285 ;
        RECT 35.260 150.730 35.400 155.170 ;
        RECT 36.180 154.130 36.320 158.910 ;
        RECT 37.100 158.890 37.240 162.310 ;
        RECT 38.880 161.290 39.140 161.610 ;
        RECT 38.940 159.570 39.080 161.290 ;
        RECT 40.320 159.910 40.460 163.330 ;
        RECT 41.240 161.610 41.380 163.670 ;
        RECT 44.000 162.030 44.140 169.790 ;
        RECT 44.860 169.450 45.120 169.770 ;
        RECT 44.400 164.350 44.660 164.670 ;
        RECT 43.540 161.890 44.140 162.030 ;
        RECT 41.180 161.290 41.440 161.610 ;
        RECT 41.640 160.950 41.900 161.270 ;
        RECT 40.260 159.590 40.520 159.910 ;
        RECT 40.720 159.590 40.980 159.910 ;
        RECT 38.880 159.250 39.140 159.570 ;
        RECT 37.500 158.910 37.760 159.230 ;
        RECT 37.040 158.570 37.300 158.890 ;
        RECT 37.100 157.190 37.240 158.570 ;
        RECT 37.040 156.870 37.300 157.190 ;
        RECT 37.100 155.490 37.240 156.870 ;
        RECT 37.560 156.170 37.700 158.910 ;
        RECT 37.500 155.850 37.760 156.170 ;
        RECT 40.780 155.910 40.920 159.590 ;
        RECT 41.700 158.210 41.840 160.950 ;
        RECT 41.640 157.890 41.900 158.210 ;
        RECT 43.540 157.190 43.680 161.890 ;
        RECT 43.940 161.290 44.200 161.610 ;
        RECT 44.000 159.230 44.140 161.290 ;
        RECT 43.940 158.910 44.200 159.230 ;
        RECT 44.460 158.630 44.600 164.350 ;
        RECT 44.920 164.330 45.060 169.450 ;
        RECT 47.220 168.070 47.360 172.170 ;
        RECT 58.660 171.490 58.920 171.810 ;
        RECT 52.220 169.790 52.480 170.110 ;
        RECT 48.540 168.770 48.800 169.090 ;
        RECT 47.160 167.750 47.420 168.070 ;
        RECT 47.220 167.050 47.360 167.750 ;
        RECT 48.600 167.390 48.740 168.770 ;
        RECT 52.280 168.070 52.420 169.790 ;
        RECT 52.220 167.750 52.480 168.070 ;
        RECT 48.540 167.070 48.800 167.390 ;
        RECT 47.160 166.730 47.420 167.050 ;
        RECT 49.000 166.790 49.260 167.050 ;
        RECT 48.600 166.730 49.260 166.790 ;
        RECT 53.600 166.730 53.860 167.050 ;
        RECT 54.980 166.730 55.240 167.050 ;
        RECT 48.600 166.650 49.200 166.730 ;
        RECT 46.240 166.050 46.500 166.370 ;
        RECT 46.300 165.010 46.440 166.050 ;
        RECT 46.240 164.690 46.500 165.010 ;
        RECT 44.860 164.010 45.120 164.330 ;
        RECT 46.700 164.010 46.960 164.330 ;
        RECT 44.000 158.490 44.600 158.630 ;
        RECT 42.100 156.870 42.360 157.190 ;
        RECT 43.480 156.870 43.740 157.190 ;
        RECT 41.170 156.335 41.450 156.705 ;
        RECT 41.240 156.170 41.380 156.335 ;
        RECT 39.860 155.770 40.920 155.910 ;
        RECT 41.180 155.850 41.440 156.170 ;
        RECT 42.160 155.830 42.300 156.870 ;
        RECT 42.560 156.530 42.820 156.850 ;
        RECT 37.040 155.170 37.300 155.490 ;
        RECT 39.860 154.470 40.000 155.770 ;
        RECT 42.100 155.510 42.360 155.830 ;
        RECT 40.260 155.170 40.520 155.490 ;
        RECT 41.180 155.170 41.440 155.490 ;
        RECT 40.320 154.470 40.460 155.170 ;
        RECT 39.800 154.150 40.060 154.470 ;
        RECT 40.260 154.150 40.520 154.470 ;
        RECT 36.120 153.810 36.380 154.130 ;
        RECT 40.720 153.810 40.980 154.130 ;
        RECT 39.800 153.470 40.060 153.790 ;
        RECT 39.860 151.150 40.000 153.470 ;
        RECT 40.780 151.750 40.920 153.810 ;
        RECT 41.240 153.790 41.380 155.170 ;
        RECT 41.180 153.470 41.440 153.790 ;
        RECT 42.620 153.110 42.760 156.530 ;
        RECT 43.010 156.335 43.290 156.705 ;
        RECT 43.080 153.110 43.220 156.335 ;
        RECT 42.560 152.790 42.820 153.110 ;
        RECT 43.020 152.790 43.280 153.110 ;
        RECT 40.720 151.430 40.980 151.750 ;
        RECT 39.860 151.010 40.920 151.150 ;
        RECT 40.780 150.730 40.920 151.010 ;
        RECT 42.620 150.730 42.760 152.790 ;
        RECT 35.200 150.410 35.460 150.730 ;
        RECT 40.720 150.410 40.980 150.730 ;
        RECT 42.560 150.410 42.820 150.730 ;
        RECT 21.400 150.070 21.660 150.390 ;
        RECT 19.560 148.030 19.820 148.350 ;
        RECT 18.640 144.630 18.900 144.950 ;
        RECT 17.260 143.270 17.520 143.590 ;
        RECT 14.960 142.590 15.220 142.910 ;
        RECT 15.020 140.530 15.160 142.590 ;
        RECT 16.800 142.250 17.060 142.570 ;
        RECT 14.960 140.210 15.220 140.530 ;
        RECT 10.810 134.575 11.090 134.945 ;
        RECT 10.880 134.410 11.020 134.575 ;
        RECT 10.820 134.090 11.080 134.410 ;
        RECT 16.860 132.710 17.000 142.250 ;
        RECT 16.800 132.390 17.060 132.710 ;
        RECT 15.880 131.370 16.140 131.690 ;
        RECT 15.420 130.690 15.680 131.010 ;
        RECT 15.480 128.970 15.620 130.690 ;
        RECT 15.940 129.990 16.080 131.370 ;
        RECT 15.880 129.670 16.140 129.990 ;
        RECT 13.580 128.650 13.840 128.970 ;
        RECT 15.420 128.650 15.680 128.970 ;
        RECT 16.800 128.650 17.060 128.970 ;
        RECT 13.640 126.590 13.780 128.650 ;
        RECT 13.580 126.270 13.840 126.590 ;
        RECT 14.960 126.270 15.220 126.590 ;
        RECT 15.020 124.550 15.160 126.270 ;
        RECT 14.960 124.230 15.220 124.550 ;
        RECT 16.860 123.870 17.000 128.650 ;
        RECT 16.800 123.550 17.060 123.870 ;
        RECT 10.820 115.390 11.080 115.710 ;
        RECT 10.880 114.545 11.020 115.390 ;
        RECT 10.810 114.175 11.090 114.545 ;
        RECT 16.860 113.330 17.000 123.550 ;
        RECT 17.320 123.530 17.460 143.270 ;
        RECT 18.180 142.930 18.440 143.250 ;
        RECT 17.720 142.250 17.980 142.570 ;
        RECT 17.780 140.870 17.920 142.250 ;
        RECT 17.720 140.550 17.980 140.870 ;
        RECT 18.240 140.780 18.380 142.930 ;
        RECT 18.700 142.230 18.840 144.630 ;
        RECT 18.640 141.910 18.900 142.230 ;
        RECT 19.620 140.870 19.760 148.030 ;
        RECT 20.480 147.690 20.740 148.010 ;
        RECT 20.540 145.290 20.680 147.690 ;
        RECT 20.480 144.970 20.740 145.290 ;
        RECT 20.940 143.270 21.200 143.590 ;
        RECT 20.480 143.105 20.740 143.250 ;
        RECT 20.470 142.990 20.750 143.105 ;
        RECT 20.080 142.850 20.750 142.990 ;
        RECT 18.240 140.640 19.300 140.780 ;
        RECT 19.160 140.190 19.300 140.640 ;
        RECT 19.560 140.550 19.820 140.870 ;
        RECT 18.640 139.870 18.900 140.190 ;
        RECT 19.100 139.870 19.360 140.190 ;
        RECT 19.550 140.015 19.830 140.385 ;
        RECT 18.700 137.810 18.840 139.870 ;
        RECT 18.640 137.490 18.900 137.810 ;
        RECT 19.620 131.690 19.760 140.015 ;
        RECT 19.560 131.370 19.820 131.690 ;
        RECT 19.560 128.310 19.820 128.630 ;
        RECT 19.620 124.550 19.760 128.310 ;
        RECT 19.560 124.230 19.820 124.550 ;
        RECT 20.080 124.210 20.220 142.850 ;
        RECT 20.470 142.735 20.750 142.850 ;
        RECT 21.000 142.425 21.140 143.270 ;
        RECT 21.460 142.570 21.600 150.070 ;
        RECT 30.950 149.195 32.490 149.565 ;
        RECT 23.700 148.030 23.960 148.350 ;
        RECT 30.140 148.030 30.400 148.350 ;
        RECT 40.260 148.030 40.520 148.350 ;
        RECT 23.240 144.290 23.500 144.610 ;
        RECT 20.930 142.055 21.210 142.425 ;
        RECT 21.400 142.250 21.660 142.570 ;
        RECT 23.300 142.480 23.440 144.290 ;
        RECT 22.840 142.340 23.440 142.480 ;
        RECT 20.480 140.550 20.740 140.870 ;
        RECT 20.540 140.385 20.680 140.550 ;
        RECT 20.470 140.015 20.750 140.385 ;
        RECT 21.460 139.760 21.600 142.250 ;
        RECT 21.860 141.910 22.120 142.230 ;
        RECT 21.920 141.745 22.060 141.910 ;
        RECT 21.850 141.375 22.130 141.745 ;
        RECT 22.320 139.760 22.580 139.850 ;
        RECT 21.460 139.620 22.580 139.760 ;
        RECT 20.940 138.850 21.200 139.170 ;
        RECT 21.000 132.030 21.140 138.850 ;
        RECT 20.940 131.710 21.200 132.030 ;
        RECT 21.920 129.310 22.060 139.620 ;
        RECT 22.320 139.530 22.580 139.620 ;
        RECT 22.840 139.170 22.980 142.340 ;
        RECT 23.760 141.890 23.900 148.030 ;
        RECT 25.540 147.350 25.800 147.670 ;
        RECT 25.600 145.290 25.740 147.350 ;
        RECT 26.460 147.010 26.720 147.330 ;
        RECT 25.540 144.970 25.800 145.290 ;
        RECT 26.000 144.290 26.260 144.610 ;
        RECT 26.060 143.590 26.200 144.290 ;
        RECT 26.000 143.270 26.260 143.590 ;
        RECT 24.160 142.590 24.420 142.910 ;
        RECT 23.700 141.570 23.960 141.890 ;
        RECT 24.220 141.745 24.360 142.590 ;
        RECT 23.240 139.530 23.500 139.850 ;
        RECT 22.780 138.850 23.040 139.170 ;
        RECT 22.320 137.490 22.580 137.810 ;
        RECT 21.860 128.990 22.120 129.310 ;
        RECT 22.380 128.970 22.520 137.490 ;
        RECT 22.840 136.450 22.980 138.850 ;
        RECT 23.300 137.810 23.440 139.530 ;
        RECT 23.240 137.490 23.500 137.810 ;
        RECT 23.760 136.790 23.900 141.570 ;
        RECT 24.150 141.375 24.430 141.745 ;
        RECT 25.540 140.550 25.800 140.870 ;
        RECT 25.600 139.510 25.740 140.550 ;
        RECT 26.000 139.760 26.260 139.850 ;
        RECT 26.520 139.760 26.660 147.010 ;
        RECT 27.650 146.475 29.190 146.845 ;
        RECT 27.380 144.970 27.640 145.290 ;
        RECT 26.920 144.630 27.180 144.950 ;
        RECT 26.000 139.620 26.660 139.760 ;
        RECT 26.000 139.530 26.260 139.620 ;
        RECT 24.160 139.190 24.420 139.510 ;
        RECT 25.540 139.190 25.800 139.510 ;
        RECT 23.700 136.470 23.960 136.790 ;
        RECT 22.780 136.130 23.040 136.450 ;
        RECT 24.220 136.190 24.360 139.190 ;
        RECT 26.520 138.150 26.660 139.620 ;
        RECT 26.460 137.830 26.720 138.150 ;
        RECT 21.400 128.650 21.660 128.970 ;
        RECT 22.320 128.650 22.580 128.970 ;
        RECT 21.460 127.270 21.600 128.650 ;
        RECT 21.860 127.970 22.120 128.290 ;
        RECT 22.320 128.200 22.580 128.290 ;
        RECT 22.840 128.200 22.980 136.130 ;
        RECT 23.760 136.050 24.360 136.190 ;
        RECT 23.760 132.030 23.900 136.050 ;
        RECT 24.160 133.410 24.420 133.730 ;
        RECT 24.220 132.030 24.360 133.410 ;
        RECT 24.620 132.050 24.880 132.370 ;
        RECT 23.700 131.710 23.960 132.030 ;
        RECT 24.160 131.710 24.420 132.030 ;
        RECT 23.760 131.430 23.900 131.710 ;
        RECT 23.760 131.290 24.360 131.430 ;
        RECT 23.700 130.690 23.960 131.010 ;
        RECT 23.760 128.970 23.900 130.690 ;
        RECT 23.700 128.825 23.960 128.970 ;
        RECT 23.240 128.310 23.500 128.630 ;
        RECT 23.690 128.455 23.970 128.825 ;
        RECT 22.320 128.060 22.980 128.200 ;
        RECT 22.320 127.970 22.580 128.060 ;
        RECT 21.400 126.950 21.660 127.270 ;
        RECT 21.920 126.590 22.060 127.970 ;
        RECT 22.380 126.590 22.520 127.970 ;
        RECT 23.300 126.590 23.440 128.310 ;
        RECT 20.940 126.270 21.200 126.590 ;
        RECT 21.860 126.270 22.120 126.590 ;
        RECT 22.320 126.270 22.580 126.590 ;
        RECT 23.240 126.270 23.500 126.590 ;
        RECT 23.700 126.270 23.960 126.590 ;
        RECT 20.020 124.120 20.280 124.210 ;
        RECT 20.020 123.980 20.680 124.120 ;
        RECT 20.020 123.890 20.280 123.980 ;
        RECT 17.260 123.210 17.520 123.530 ;
        RECT 18.180 123.210 18.440 123.530 ;
        RECT 16.800 113.010 17.060 113.330 ;
        RECT 17.320 112.990 17.460 123.210 ;
        RECT 17.720 121.510 17.980 121.830 ;
        RECT 17.260 112.670 17.520 112.990 ;
        RECT 17.780 112.505 17.920 121.510 ;
        RECT 18.240 120.470 18.380 123.210 ;
        RECT 19.100 122.530 19.360 122.850 ;
        RECT 19.160 121.830 19.300 122.530 ;
        RECT 19.100 121.510 19.360 121.830 ;
        RECT 18.640 120.490 18.900 120.810 ;
        RECT 18.180 120.150 18.440 120.470 ;
        RECT 18.700 118.410 18.840 120.490 ;
        RECT 18.240 118.270 18.840 118.410 ;
        RECT 17.710 112.135 17.990 112.505 ;
        RECT 17.720 111.990 17.980 112.135 ;
        RECT 14.040 111.650 14.300 111.970 ;
        RECT 13.580 109.610 13.840 109.930 ;
        RECT 13.640 108.230 13.780 109.610 ;
        RECT 13.580 107.910 13.840 108.230 ;
        RECT 13.640 107.550 13.780 107.910 ;
        RECT 13.580 107.230 13.840 107.550 ;
        RECT 14.100 107.210 14.240 111.650 ;
        RECT 14.040 106.890 14.300 107.210 ;
        RECT 18.240 103.810 18.380 118.270 ;
        RECT 20.540 112.990 20.680 123.980 ;
        RECT 21.000 123.530 21.140 126.270 ;
        RECT 21.400 125.250 21.660 125.570 ;
        RECT 21.460 124.550 21.600 125.250 ;
        RECT 21.400 124.230 21.660 124.550 ;
        RECT 21.460 123.530 21.600 124.230 ;
        RECT 21.920 124.210 22.060 126.270 ;
        RECT 21.860 123.890 22.120 124.210 ;
        RECT 23.240 123.550 23.500 123.870 ;
        RECT 20.940 123.210 21.200 123.530 ;
        RECT 21.400 123.210 21.660 123.530 ;
        RECT 22.780 123.210 23.040 123.530 ;
        RECT 21.000 121.830 21.140 123.210 ;
        RECT 21.460 122.590 21.600 123.210 ;
        RECT 21.860 123.100 22.120 123.190 ;
        RECT 21.860 122.960 22.520 123.100 ;
        RECT 21.860 122.870 22.120 122.960 ;
        RECT 21.460 122.450 22.060 122.590 ;
        RECT 20.940 121.510 21.200 121.830 ;
        RECT 21.920 121.150 22.060 122.450 ;
        RECT 21.860 120.830 22.120 121.150 ;
        RECT 22.380 120.130 22.520 122.960 ;
        RECT 22.840 120.810 22.980 123.210 ;
        RECT 22.780 120.490 23.040 120.810 ;
        RECT 22.320 119.810 22.580 120.130 ;
        RECT 22.380 115.710 22.520 119.810 ;
        RECT 23.300 119.110 23.440 123.550 ;
        RECT 23.240 118.790 23.500 119.110 ;
        RECT 23.240 118.410 23.500 118.430 ;
        RECT 23.760 118.410 23.900 126.270 ;
        RECT 24.220 121.830 24.360 131.290 ;
        RECT 24.680 128.970 24.820 132.050 ;
        RECT 26.520 132.030 26.660 137.830 ;
        RECT 26.980 136.790 27.120 144.630 ;
        RECT 27.440 143.250 27.580 144.970 ;
        RECT 29.680 144.630 29.940 144.950 ;
        RECT 27.380 142.930 27.640 143.250 ;
        RECT 27.440 141.890 27.580 142.930 ;
        RECT 27.380 141.570 27.640 141.890 ;
        RECT 27.650 141.035 29.190 141.405 ;
        RECT 29.740 140.530 29.880 144.630 ;
        RECT 30.200 143.590 30.340 148.030 ;
        RECT 35.660 147.350 35.920 147.670 ;
        RECT 34.740 144.970 35.000 145.290 ;
        RECT 32.900 144.290 33.160 144.610 ;
        RECT 30.950 143.755 32.490 144.125 ;
        RECT 30.140 143.270 30.400 143.590 ;
        RECT 29.680 140.210 29.940 140.530 ;
        RECT 27.840 139.870 28.100 140.190 ;
        RECT 27.900 139.170 28.040 139.870 ;
        RECT 28.760 139.190 29.020 139.510 ;
        RECT 27.840 138.850 28.100 139.170 ;
        RECT 28.820 137.130 28.960 139.190 ;
        RECT 29.680 138.850 29.940 139.170 ;
        RECT 28.760 136.810 29.020 137.130 ;
        RECT 26.920 136.470 27.180 136.790 ;
        RECT 27.650 135.595 29.190 135.965 ;
        RECT 29.740 134.750 29.880 138.850 ;
        RECT 30.200 137.810 30.340 143.270 ;
        RECT 30.590 142.735 30.870 143.105 ;
        RECT 30.660 140.190 30.800 142.735 ;
        RECT 31.520 142.590 31.780 142.910 ;
        RECT 30.600 139.870 30.860 140.190 ;
        RECT 30.600 139.190 30.860 139.510 ;
        RECT 30.140 137.490 30.400 137.810 ;
        RECT 29.680 134.430 29.940 134.750 ;
        RECT 29.740 132.710 29.880 134.430 ;
        RECT 29.680 132.390 29.940 132.710 ;
        RECT 30.200 132.370 30.340 137.490 ;
        RECT 30.660 137.470 30.800 139.190 ;
        RECT 31.580 139.170 31.720 142.590 ;
        RECT 31.970 142.055 32.250 142.425 ;
        RECT 32.040 140.190 32.180 142.055 ;
        RECT 31.980 139.870 32.240 140.190 ;
        RECT 31.520 138.850 31.780 139.170 ;
        RECT 32.040 139.080 32.180 139.870 ;
        RECT 32.960 139.510 33.100 144.290 ;
        RECT 34.800 141.890 34.940 144.970 ;
        RECT 34.740 141.570 35.000 141.890 ;
        RECT 34.280 139.870 34.540 140.190 ;
        RECT 33.360 139.530 33.620 139.850 ;
        RECT 32.900 139.190 33.160 139.510 ;
        RECT 32.040 138.940 32.765 139.080 ;
        RECT 32.625 138.910 32.765 138.940 ;
        RECT 32.625 138.770 33.100 138.910 ;
        RECT 30.950 138.315 32.490 138.685 ;
        RECT 30.600 137.150 30.860 137.470 ;
        RECT 30.660 136.450 30.800 137.150 ;
        RECT 30.600 136.130 30.860 136.450 ;
        RECT 30.660 132.620 30.800 136.130 ;
        RECT 30.950 132.875 32.490 133.245 ;
        RECT 30.660 132.480 31.260 132.620 ;
        RECT 30.140 132.050 30.400 132.370 ;
        RECT 26.460 131.710 26.720 132.030 ;
        RECT 26.000 131.370 26.260 131.690 ;
        RECT 30.200 131.430 30.340 132.050 ;
        RECT 31.120 131.690 31.260 132.480 ;
        RECT 25.540 131.030 25.800 131.350 ;
        RECT 24.620 128.650 24.880 128.970 ;
        RECT 25.080 126.500 25.340 126.590 ;
        RECT 25.600 126.500 25.740 131.030 ;
        RECT 26.060 128.710 26.200 131.370 ;
        RECT 29.680 131.030 29.940 131.350 ;
        RECT 30.200 131.290 30.800 131.430 ;
        RECT 31.060 131.370 31.320 131.690 ;
        RECT 26.920 130.690 27.180 131.010 ;
        RECT 26.460 129.505 26.720 129.650 ;
        RECT 26.450 129.135 26.730 129.505 ;
        RECT 26.980 128.970 27.120 130.690 ;
        RECT 27.650 130.155 29.190 130.525 ;
        RECT 27.840 129.670 28.100 129.990 ;
        RECT 26.060 128.570 26.660 128.710 ;
        RECT 26.920 128.650 27.180 128.970 ;
        RECT 26.520 128.030 26.660 128.570 ;
        RECT 26.920 128.030 27.180 128.290 ;
        RECT 26.520 127.970 27.180 128.030 ;
        RECT 26.520 127.890 27.120 127.970 ;
        RECT 25.080 126.360 25.740 126.500 ;
        RECT 25.080 126.270 25.340 126.360 ;
        RECT 24.620 125.930 24.880 126.250 ;
        RECT 24.160 121.510 24.420 121.830 ;
        RECT 23.240 118.340 23.900 118.410 ;
        RECT 22.840 118.270 23.900 118.340 ;
        RECT 22.840 118.200 23.500 118.270 ;
        RECT 22.320 115.390 22.580 115.710 ;
        RECT 20.480 112.900 20.740 112.990 ;
        RECT 19.620 112.760 20.740 112.900 ;
        RECT 18.640 112.560 18.900 112.650 ;
        RECT 19.620 112.560 19.760 112.760 ;
        RECT 20.480 112.670 20.740 112.760 ;
        RECT 18.640 112.420 19.760 112.560 ;
        RECT 20.940 112.505 21.200 112.650 ;
        RECT 18.640 112.330 18.900 112.420 ;
        RECT 20.930 112.135 21.210 112.505 ;
        RECT 18.640 111.650 18.900 111.970 ;
        RECT 18.700 110.610 18.840 111.650 ;
        RECT 18.640 110.290 18.900 110.610 ;
        RECT 21.000 110.270 21.140 112.135 ;
        RECT 21.400 111.990 21.660 112.310 ;
        RECT 20.940 109.950 21.200 110.270 ;
        RECT 21.000 107.890 21.140 109.950 ;
        RECT 21.460 109.930 21.600 111.990 ;
        RECT 22.380 110.950 22.520 115.390 ;
        RECT 22.320 110.630 22.580 110.950 ;
        RECT 22.380 110.270 22.520 110.630 ;
        RECT 22.320 109.950 22.580 110.270 ;
        RECT 21.400 109.610 21.660 109.930 ;
        RECT 20.940 107.570 21.200 107.890 ;
        RECT 18.180 103.490 18.440 103.810 ;
        RECT 20.020 103.490 20.280 103.810 ;
        RECT 22.320 103.720 22.580 103.810 ;
        RECT 22.840 103.720 22.980 118.200 ;
        RECT 23.240 118.110 23.500 118.200 ;
        RECT 24.680 116.390 24.820 125.930 ;
        RECT 24.620 116.070 24.880 116.390 ;
        RECT 23.240 115.390 23.500 115.710 ;
        RECT 23.300 113.670 23.440 115.390 ;
        RECT 23.700 114.370 23.960 114.690 ;
        RECT 23.240 113.350 23.500 113.670 ;
        RECT 23.760 112.650 23.900 114.370 ;
        RECT 23.700 112.330 23.960 112.650 ;
        RECT 23.760 106.530 23.900 112.330 ;
        RECT 24.680 111.030 24.820 116.070 ;
        RECT 25.140 111.710 25.280 126.270 ;
        RECT 26.980 126.250 27.120 127.890 ;
        RECT 27.900 126.590 28.040 129.670 ;
        RECT 27.840 126.270 28.100 126.590 ;
        RECT 26.920 125.930 27.180 126.250 ;
        RECT 25.540 125.250 25.800 125.570 ;
        RECT 26.920 125.250 27.180 125.570 ;
        RECT 25.600 123.530 25.740 125.250 ;
        RECT 25.540 123.210 25.800 123.530 ;
        RECT 26.980 123.440 27.120 125.250 ;
        RECT 27.650 124.715 29.190 125.085 ;
        RECT 27.380 123.440 27.640 123.530 ;
        RECT 26.980 123.300 27.640 123.440 ;
        RECT 25.540 121.510 25.800 121.830 ;
        RECT 25.600 113.670 25.740 121.510 ;
        RECT 26.980 121.150 27.120 123.300 ;
        RECT 27.380 123.210 27.640 123.300 ;
        RECT 29.740 123.270 29.880 131.030 ;
        RECT 30.140 130.690 30.400 131.010 ;
        RECT 27.840 122.870 28.100 123.190 ;
        RECT 28.820 123.130 29.880 123.270 ;
        RECT 26.920 120.830 27.180 121.150 ;
        RECT 27.900 120.470 28.040 122.870 ;
        RECT 28.820 121.150 28.960 123.130 ;
        RECT 30.200 122.850 30.340 130.690 ;
        RECT 30.660 125.910 30.800 131.290 ;
        RECT 31.120 129.990 31.260 131.370 ;
        RECT 31.060 129.670 31.320 129.990 ;
        RECT 31.520 129.220 31.780 129.310 ;
        RECT 32.960 129.220 33.100 138.770 ;
        RECT 33.420 138.150 33.560 139.530 ;
        RECT 34.340 138.150 34.480 139.870 ;
        RECT 33.360 137.830 33.620 138.150 ;
        RECT 34.280 137.830 34.540 138.150 ;
        RECT 33.420 137.130 33.560 137.830 ;
        RECT 33.360 136.810 33.620 137.130 ;
        RECT 33.420 129.990 33.560 136.810 ;
        RECT 34.800 134.070 34.940 141.570 ;
        RECT 35.720 139.510 35.860 147.350 ;
        RECT 36.580 144.630 36.840 144.950 ;
        RECT 36.110 142.735 36.390 143.105 ;
        RECT 35.660 139.190 35.920 139.510 ;
        RECT 36.180 139.170 36.320 142.735 ;
        RECT 36.640 140.530 36.780 144.630 ;
        RECT 40.320 144.610 40.460 148.030 ;
        RECT 37.960 144.290 38.220 144.610 ;
        RECT 40.260 144.290 40.520 144.610 ;
        RECT 37.040 141.570 37.300 141.890 ;
        RECT 36.580 140.210 36.840 140.530 ;
        RECT 36.580 139.760 36.840 139.850 ;
        RECT 37.100 139.760 37.240 141.570 ;
        RECT 38.020 139.850 38.160 144.290 ;
        RECT 36.580 139.620 37.240 139.760 ;
        RECT 36.580 139.530 36.840 139.620 ;
        RECT 35.200 138.850 35.460 139.170 ;
        RECT 36.120 138.850 36.380 139.170 ;
        RECT 35.260 137.470 35.400 138.850 ;
        RECT 35.200 137.150 35.460 137.470 ;
        RECT 35.660 137.150 35.920 137.470 ;
        RECT 35.720 136.450 35.860 137.150 ;
        RECT 35.660 136.130 35.920 136.450 ;
        RECT 34.740 133.750 35.000 134.070 ;
        RECT 34.800 132.030 34.940 133.750 ;
        RECT 35.720 132.030 35.860 136.130 ;
        RECT 34.740 131.710 35.000 132.030 ;
        RECT 35.660 131.710 35.920 132.030 ;
        RECT 33.820 130.690 34.080 131.010 ;
        RECT 33.360 129.670 33.620 129.990 ;
        RECT 33.880 129.310 34.020 130.690 ;
        RECT 31.520 129.080 33.560 129.220 ;
        RECT 31.520 128.990 31.780 129.080 ;
        RECT 33.420 128.710 33.560 129.080 ;
        RECT 33.820 128.990 34.080 129.310 ;
        RECT 32.440 128.540 32.700 128.630 ;
        RECT 33.420 128.570 34.020 128.710 ;
        RECT 32.440 128.400 33.100 128.540 ;
        RECT 32.440 128.310 32.700 128.400 ;
        RECT 30.950 127.435 32.490 127.805 ;
        RECT 30.600 125.590 30.860 125.910 ;
        RECT 29.680 122.530 29.940 122.850 ;
        RECT 30.140 122.530 30.400 122.850 ;
        RECT 30.600 122.530 30.860 122.850 ;
        RECT 28.760 120.830 29.020 121.150 ;
        RECT 27.840 120.150 28.100 120.470 ;
        RECT 27.650 119.275 29.190 119.645 ;
        RECT 28.760 118.790 29.020 119.110 ;
        RECT 28.300 118.450 28.560 118.770 ;
        RECT 26.460 117.770 26.720 118.090 ;
        RECT 26.000 117.430 26.260 117.750 ;
        RECT 26.060 116.390 26.200 117.430 ;
        RECT 26.000 116.070 26.260 116.390 ;
        RECT 26.000 115.390 26.260 115.710 ;
        RECT 26.060 114.690 26.200 115.390 ;
        RECT 26.000 114.370 26.260 114.690 ;
        RECT 25.540 113.350 25.800 113.670 ;
        RECT 25.140 111.570 25.740 111.710 ;
        RECT 24.680 110.890 25.280 111.030 ;
        RECT 24.620 109.950 24.880 110.270 ;
        RECT 24.680 108.230 24.820 109.950 ;
        RECT 24.620 107.910 24.880 108.230 ;
        RECT 23.700 106.210 23.960 106.530 ;
        RECT 23.760 105.510 23.900 106.210 ;
        RECT 23.700 105.190 23.960 105.510 ;
        RECT 25.140 105.170 25.280 110.890 ;
        RECT 25.080 104.850 25.340 105.170 ;
        RECT 22.320 103.580 22.980 103.720 ;
        RECT 22.320 103.490 22.580 103.580 ;
        RECT 18.640 99.300 18.900 99.390 ;
        RECT 18.640 99.160 19.300 99.300 ;
        RECT 18.640 99.070 18.900 99.160 ;
        RECT 17.260 98.050 17.520 98.370 ;
        RECT 16.340 97.030 16.600 97.350 ;
        RECT 7.140 96.350 7.400 96.670 ;
        RECT 15.420 95.670 15.680 95.990 ;
        RECT 13.580 95.560 13.840 95.650 ;
        RECT 13.580 95.420 14.240 95.560 ;
        RECT 13.580 95.330 13.840 95.420 ;
        RECT 13.580 93.630 13.840 93.950 ;
        RECT 13.640 91.230 13.780 93.630 ;
        RECT 13.580 90.910 13.840 91.230 ;
        RECT 13.640 88.510 13.780 90.910 ;
        RECT 14.100 90.890 14.240 95.420 ;
        RECT 14.500 95.330 14.760 95.650 ;
        RECT 14.040 90.570 14.300 90.890 ;
        RECT 13.580 88.190 13.840 88.510 ;
        RECT 14.560 83.750 14.700 95.330 ;
        RECT 14.960 88.190 15.220 88.510 ;
        RECT 15.020 86.470 15.160 88.190 ;
        RECT 15.480 86.470 15.620 95.670 ;
        RECT 15.880 95.330 16.140 95.650 ;
        RECT 15.940 93.950 16.080 95.330 ;
        RECT 15.880 93.630 16.140 93.950 ;
        RECT 14.960 86.150 15.220 86.470 ;
        RECT 15.420 86.150 15.680 86.470 ;
        RECT 16.400 85.110 16.540 97.030 ;
        RECT 16.800 88.190 17.060 88.510 ;
        RECT 16.340 85.020 16.600 85.110 ;
        RECT 15.940 84.880 16.600 85.020 ;
        RECT 14.500 83.430 14.760 83.750 ;
        RECT 14.960 73.910 15.220 74.230 ;
        RECT 15.020 72.870 15.160 73.910 ;
        RECT 14.960 72.550 15.220 72.870 ;
        RECT 15.940 72.190 16.080 84.880 ;
        RECT 16.340 84.790 16.600 84.880 ;
        RECT 16.860 83.070 17.000 88.190 ;
        RECT 17.320 83.070 17.460 98.050 ;
        RECT 18.640 96.185 18.900 96.330 ;
        RECT 18.180 95.670 18.440 95.990 ;
        RECT 18.630 95.815 18.910 96.185 ;
        RECT 18.240 91.910 18.380 95.670 ;
        RECT 19.160 95.650 19.300 99.160 ;
        RECT 20.080 96.330 20.220 103.490 ;
        RECT 21.860 99.070 22.120 99.390 ;
        RECT 20.540 97.350 21.140 97.430 ;
        RECT 20.540 97.290 21.200 97.350 ;
        RECT 20.020 96.010 20.280 96.330 ;
        RECT 18.640 95.330 18.900 95.650 ;
        RECT 19.100 95.330 19.360 95.650 ;
        RECT 18.180 91.590 18.440 91.910 ;
        RECT 16.800 82.750 17.060 83.070 ;
        RECT 17.260 82.750 17.520 83.070 ;
        RECT 16.860 77.630 17.000 82.750 ;
        RECT 16.800 77.310 17.060 77.630 ;
        RECT 16.340 76.290 16.600 76.610 ;
        RECT 16.400 72.870 16.540 76.290 ;
        RECT 16.340 72.550 16.600 72.870 ;
        RECT 16.860 72.190 17.000 77.310 ;
        RECT 15.880 71.870 16.140 72.190 ;
        RECT 16.800 71.870 17.060 72.190 ;
        RECT 14.040 68.470 14.300 68.790 ;
        RECT 14.100 67.430 14.240 68.470 ;
        RECT 15.420 68.130 15.680 68.450 ;
        RECT 14.040 67.110 14.300 67.430 ;
        RECT 15.480 64.710 15.620 68.130 ;
        RECT 15.940 67.090 16.080 71.870 ;
        RECT 18.240 71.850 18.380 91.590 ;
        RECT 18.700 83.750 18.840 95.330 ;
        RECT 18.640 83.430 18.900 83.750 ;
        RECT 19.160 83.070 19.300 95.330 ;
        RECT 20.540 93.350 20.680 97.290 ;
        RECT 20.940 97.030 21.200 97.290 ;
        RECT 21.400 96.690 21.660 97.010 ;
        RECT 21.460 94.630 21.600 96.690 ;
        RECT 21.920 96.330 22.060 99.070 ;
        RECT 21.860 96.010 22.120 96.330 ;
        RECT 21.400 94.310 21.660 94.630 ;
        RECT 20.540 93.210 21.140 93.350 ;
        RECT 21.000 90.550 21.140 93.210 ;
        RECT 20.940 90.230 21.200 90.550 ;
        RECT 21.000 88.590 21.140 90.230 ;
        RECT 21.460 89.190 21.600 94.310 ;
        RECT 21.920 90.210 22.060 96.010 ;
        RECT 22.380 95.650 22.520 103.490 ;
        RECT 25.600 99.730 25.740 111.570 ;
        RECT 26.060 109.250 26.200 114.370 ;
        RECT 26.520 110.610 26.660 117.770 ;
        RECT 28.360 115.710 28.500 118.450 ;
        RECT 28.820 115.710 28.960 118.790 ;
        RECT 29.740 118.430 29.880 122.530 ;
        RECT 30.140 120.830 30.400 121.150 ;
        RECT 30.200 120.470 30.340 120.830 ;
        RECT 30.140 120.150 30.400 120.470 ;
        RECT 29.680 118.110 29.940 118.430 ;
        RECT 30.200 117.750 30.340 120.150 ;
        RECT 30.660 118.090 30.800 122.530 ;
        RECT 30.950 121.995 32.490 122.365 ;
        RECT 31.520 120.490 31.780 120.810 ;
        RECT 31.060 119.810 31.320 120.130 ;
        RECT 30.600 117.770 30.860 118.090 ;
        RECT 30.140 117.430 30.400 117.750 ;
        RECT 29.680 117.090 29.940 117.410 ;
        RECT 31.120 117.320 31.260 119.810 ;
        RECT 31.580 119.110 31.720 120.490 ;
        RECT 31.980 120.150 32.240 120.470 ;
        RECT 31.520 118.790 31.780 119.110 ;
        RECT 32.040 118.770 32.180 120.150 ;
        RECT 31.980 118.450 32.240 118.770 ;
        RECT 30.660 117.180 31.260 117.320 ;
        RECT 28.300 115.390 28.560 115.710 ;
        RECT 28.760 115.390 29.020 115.710 ;
        RECT 27.650 113.835 29.190 114.205 ;
        RECT 28.300 112.330 28.560 112.650 ;
        RECT 29.220 112.330 29.480 112.650 ;
        RECT 27.370 110.775 27.650 111.145 ;
        RECT 28.360 110.950 28.500 112.330 ;
        RECT 26.460 110.290 26.720 110.610 ;
        RECT 26.000 108.930 26.260 109.250 ;
        RECT 26.520 105.170 26.660 110.290 ;
        RECT 27.440 110.270 27.580 110.775 ;
        RECT 28.300 110.630 28.560 110.950 ;
        RECT 27.380 109.950 27.640 110.270 ;
        RECT 26.920 109.610 27.180 109.930 ;
        RECT 29.280 109.670 29.420 112.330 ;
        RECT 29.740 110.270 29.880 117.090 ;
        RECT 30.140 114.370 30.400 114.690 ;
        RECT 29.680 109.950 29.940 110.270 ;
        RECT 26.980 108.140 27.120 109.610 ;
        RECT 29.280 109.530 29.880 109.670 ;
        RECT 27.650 108.395 29.190 108.765 ;
        RECT 27.380 108.140 27.640 108.230 ;
        RECT 26.980 108.000 27.640 108.140 ;
        RECT 27.380 107.910 27.640 108.000 ;
        RECT 28.300 107.910 28.560 108.230 ;
        RECT 29.220 107.910 29.480 108.230 ;
        RECT 27.840 106.890 28.100 107.210 ;
        RECT 27.380 106.550 27.640 106.870 ;
        RECT 27.440 105.510 27.580 106.550 ;
        RECT 27.380 105.190 27.640 105.510 ;
        RECT 26.460 104.850 26.720 105.170 ;
        RECT 27.900 104.830 28.040 106.890 ;
        RECT 28.360 106.530 28.500 107.910 ;
        RECT 28.760 106.890 29.020 107.210 ;
        RECT 28.300 106.210 28.560 106.530 ;
        RECT 26.920 104.510 27.180 104.830 ;
        RECT 27.840 104.510 28.100 104.830 ;
        RECT 26.460 103.830 26.720 104.150 ;
        RECT 26.520 100.070 26.660 103.830 ;
        RECT 26.980 102.700 27.120 104.510 ;
        RECT 27.900 104.345 28.040 104.510 ;
        RECT 27.830 103.975 28.110 104.345 ;
        RECT 28.360 103.810 28.500 106.210 ;
        RECT 28.820 104.490 28.960 106.890 ;
        RECT 28.760 104.170 29.020 104.490 ;
        RECT 29.280 104.150 29.420 107.910 ;
        RECT 29.220 103.830 29.480 104.150 ;
        RECT 28.300 103.490 28.560 103.810 ;
        RECT 27.650 102.955 29.190 103.325 ;
        RECT 26.980 102.560 27.580 102.700 ;
        RECT 26.460 99.750 26.720 100.070 ;
        RECT 27.440 99.730 27.580 102.560 ;
        RECT 22.780 99.410 23.040 99.730 ;
        RECT 25.540 99.410 25.800 99.730 ;
        RECT 27.380 99.410 27.640 99.730 ;
        RECT 22.320 95.330 22.580 95.650 ;
        RECT 22.310 93.775 22.590 94.145 ;
        RECT 22.320 93.630 22.580 93.775 ;
        RECT 21.860 89.890 22.120 90.210 ;
        RECT 21.400 88.870 21.660 89.190 ;
        RECT 21.000 88.450 21.600 88.590 ;
        RECT 20.480 87.510 20.740 87.830 ;
        RECT 20.020 86.150 20.280 86.470 ;
        RECT 20.080 85.985 20.220 86.150 ;
        RECT 20.010 85.615 20.290 85.985 ;
        RECT 20.540 85.790 20.680 87.510 ;
        RECT 21.460 87.490 21.600 88.450 ;
        RECT 21.920 88.420 22.060 89.890 ;
        RECT 22.320 88.420 22.580 88.510 ;
        RECT 21.920 88.280 22.580 88.420 ;
        RECT 21.400 87.170 21.660 87.490 ;
        RECT 20.930 86.295 21.210 86.665 ;
        RECT 20.480 85.470 20.740 85.790 ;
        RECT 21.000 85.450 21.140 86.295 ;
        RECT 20.940 85.130 21.200 85.450 ;
        RECT 19.100 82.750 19.360 83.070 ;
        RECT 20.940 77.990 21.200 78.310 ;
        RECT 18.640 76.970 18.900 77.290 ;
        RECT 18.700 75.250 18.840 76.970 ;
        RECT 18.640 74.930 18.900 75.250 ;
        RECT 18.700 72.530 18.840 74.930 ;
        RECT 21.000 74.570 21.140 77.990 ;
        RECT 20.940 74.480 21.200 74.570 ;
        RECT 20.540 74.340 21.200 74.480 ;
        RECT 18.640 72.270 18.900 72.530 ;
        RECT 18.640 72.210 20.220 72.270 ;
        RECT 18.700 72.130 20.220 72.210 ;
        RECT 18.180 71.530 18.440 71.850 ;
        RECT 19.100 71.530 19.360 71.850 ;
        RECT 19.160 69.130 19.300 71.530 ;
        RECT 19.560 71.190 19.820 71.510 ;
        RECT 19.100 68.810 19.360 69.130 ;
        RECT 17.720 68.130 17.980 68.450 ;
        RECT 18.180 68.130 18.440 68.450 ;
        RECT 17.780 67.430 17.920 68.130 ;
        RECT 17.720 67.110 17.980 67.430 ;
        RECT 15.880 66.770 16.140 67.090 ;
        RECT 15.420 64.390 15.680 64.710 ;
        RECT 14.960 63.030 15.220 63.350 ;
        RECT 15.020 61.990 15.160 63.030 ;
        RECT 14.960 61.670 15.220 61.990 ;
        RECT 15.940 60.290 16.080 66.770 ;
        RECT 17.780 63.350 17.920 67.110 ;
        RECT 17.720 63.030 17.980 63.350 ;
        RECT 16.800 62.690 17.060 63.010 ;
        RECT 16.860 61.650 17.000 62.690 ;
        RECT 16.800 61.330 17.060 61.650 ;
        RECT 15.880 59.970 16.140 60.290 ;
        RECT 15.940 53.830 16.080 59.970 ;
        RECT 15.880 53.510 16.140 53.830 ;
        RECT 14.500 53.170 14.760 53.490 ;
        RECT 14.040 52.150 14.300 52.470 ;
        RECT 14.100 45.330 14.240 52.150 ;
        RECT 14.040 45.010 14.300 45.330 ;
        RECT 14.560 44.990 14.700 53.170 ;
        RECT 15.420 51.810 15.680 52.130 ;
        RECT 14.960 47.050 15.220 47.370 ;
        RECT 15.480 47.280 15.620 51.810 ;
        RECT 15.940 47.790 16.080 53.510 ;
        RECT 16.860 52.470 17.000 61.330 ;
        RECT 18.240 61.310 18.380 68.130 ;
        RECT 19.620 63.010 19.760 71.190 ;
        RECT 20.080 69.470 20.220 72.130 ;
        RECT 20.540 71.850 20.680 74.340 ;
        RECT 20.940 74.250 21.200 74.340 ;
        RECT 20.940 73.570 21.200 73.890 ;
        RECT 21.000 72.530 21.140 73.570 ;
        RECT 20.940 72.210 21.200 72.530 ;
        RECT 20.480 71.760 20.740 71.850 ;
        RECT 20.480 71.620 21.140 71.760 ;
        RECT 20.480 71.530 20.740 71.620 ;
        RECT 20.020 69.150 20.280 69.470 ;
        RECT 20.480 68.470 20.740 68.790 ;
        RECT 20.540 64.710 20.680 68.470 ;
        RECT 21.000 68.305 21.140 71.620 ;
        RECT 20.930 67.935 21.210 68.305 ;
        RECT 20.940 67.110 21.200 67.430 ;
        RECT 21.000 65.470 21.140 67.110 ;
        RECT 21.460 66.150 21.600 87.170 ;
        RECT 21.920 86.130 22.060 88.280 ;
        RECT 22.320 88.190 22.580 88.280 ;
        RECT 22.840 86.380 22.980 99.410 ;
        RECT 27.650 97.515 29.190 97.885 ;
        RECT 29.740 97.350 29.880 109.530 ;
        RECT 30.200 107.550 30.340 114.370 ;
        RECT 30.660 113.330 30.800 117.180 ;
        RECT 30.950 116.555 32.490 116.925 ;
        RECT 32.960 116.390 33.100 128.400 ;
        RECT 33.880 128.290 34.020 128.570 ;
        RECT 34.280 128.310 34.540 128.630 ;
        RECT 33.360 127.970 33.620 128.290 ;
        RECT 33.820 127.970 34.080 128.290 ;
        RECT 33.420 126.590 33.560 127.970 ;
        RECT 33.360 126.270 33.620 126.590 ;
        RECT 33.360 122.530 33.620 122.850 ;
        RECT 33.420 120.470 33.560 122.530 ;
        RECT 33.880 121.490 34.020 127.970 ;
        RECT 33.820 121.170 34.080 121.490 ;
        RECT 33.360 120.150 33.620 120.470 ;
        RECT 33.880 119.870 34.020 121.170 ;
        RECT 34.340 120.810 34.480 128.310 ;
        RECT 34.800 126.930 34.940 131.710 ;
        RECT 35.660 131.030 35.920 131.350 ;
        RECT 34.740 126.610 35.000 126.930 ;
        RECT 35.720 121.150 35.860 131.030 ;
        RECT 36.180 129.310 36.320 138.850 ;
        RECT 37.100 137.810 37.240 139.620 ;
        RECT 37.960 139.530 38.220 139.850 ;
        RECT 37.040 137.490 37.300 137.810 ;
        RECT 36.120 128.990 36.380 129.310 ;
        RECT 37.100 128.630 37.240 137.490 ;
        RECT 39.340 136.810 39.600 137.130 ;
        RECT 39.400 135.430 39.540 136.810 ;
        RECT 39.340 135.110 39.600 135.430 ;
        RECT 40.780 135.090 40.920 150.410 ;
        RECT 41.640 148.370 41.900 148.690 ;
        RECT 44.000 148.430 44.140 158.490 ;
        RECT 44.920 151.070 45.060 164.010 ;
        RECT 46.760 162.630 46.900 164.010 ;
        RECT 46.700 162.310 46.960 162.630 ;
        RECT 48.600 161.610 48.740 166.650 ;
        RECT 50.840 166.390 51.100 166.710 ;
        RECT 49.000 166.050 49.260 166.370 ;
        RECT 49.060 164.670 49.200 166.050 ;
        RECT 49.000 164.350 49.260 164.670 ;
        RECT 49.000 161.970 49.260 162.290 ;
        RECT 49.060 161.610 49.200 161.970 ;
        RECT 50.900 161.610 51.040 166.390 ;
        RECT 53.660 163.650 53.800 166.730 ;
        RECT 55.040 164.670 55.180 166.730 ;
        RECT 58.720 166.710 58.860 171.490 ;
        RECT 58.720 166.570 59.320 166.710 ;
        RECT 54.980 164.350 55.240 164.670 ;
        RECT 56.360 164.350 56.620 164.670 ;
        RECT 53.600 163.330 53.860 163.650 ;
        RECT 48.540 161.290 48.800 161.610 ;
        RECT 49.000 161.290 49.260 161.610 ;
        RECT 50.840 161.290 51.100 161.610 ;
        RECT 52.220 161.290 52.480 161.610 ;
        RECT 52.680 161.290 52.940 161.610 ;
        RECT 46.700 160.610 46.960 160.930 ;
        RECT 46.760 159.570 46.900 160.610 ;
        RECT 46.700 159.250 46.960 159.570 ;
        RECT 46.240 158.910 46.500 159.230 ;
        RECT 45.320 157.890 45.580 158.210 ;
        RECT 45.380 156.510 45.520 157.890 ;
        RECT 45.780 156.870 46.040 157.190 ;
        RECT 45.320 156.190 45.580 156.510 ;
        RECT 44.860 150.750 45.120 151.070 ;
        RECT 44.400 149.730 44.660 150.050 ;
        RECT 41.180 147.010 41.440 147.330 ;
        RECT 41.240 142.910 41.380 147.010 ;
        RECT 41.700 146.310 41.840 148.370 ;
        RECT 42.100 148.030 42.360 148.350 ;
        RECT 43.020 148.030 43.280 148.350 ;
        RECT 43.540 148.290 44.140 148.430 ;
        RECT 41.640 145.990 41.900 146.310 ;
        RECT 42.160 145.970 42.300 148.030 ;
        RECT 42.560 147.690 42.820 148.010 ;
        RECT 42.100 145.650 42.360 145.970 ;
        RECT 41.640 144.290 41.900 144.610 ;
        RECT 41.180 142.590 41.440 142.910 ;
        RECT 41.180 139.190 41.440 139.510 ;
        RECT 41.240 138.150 41.380 139.190 ;
        RECT 41.180 137.830 41.440 138.150 ;
        RECT 41.700 135.430 41.840 144.290 ;
        RECT 42.100 142.930 42.360 143.250 ;
        RECT 42.160 139.850 42.300 142.930 ;
        RECT 42.100 139.530 42.360 139.850 ;
        RECT 42.620 136.790 42.760 147.690 ;
        RECT 43.080 144.950 43.220 148.030 ;
        RECT 43.540 146.310 43.680 148.290 ;
        RECT 43.480 145.990 43.740 146.310 ;
        RECT 43.020 144.630 43.280 144.950 ;
        RECT 43.080 140.870 43.220 144.630 ;
        RECT 43.020 140.550 43.280 140.870 ;
        RECT 42.560 136.470 42.820 136.790 ;
        RECT 41.640 135.110 41.900 135.430 ;
        RECT 40.720 134.770 40.980 135.090 ;
        RECT 39.800 134.430 40.060 134.750 ;
        RECT 37.500 131.030 37.760 131.350 ;
        RECT 37.960 131.030 38.220 131.350 ;
        RECT 37.560 129.990 37.700 131.030 ;
        RECT 37.500 129.670 37.760 129.990 ;
        RECT 37.040 128.310 37.300 128.630 ;
        RECT 36.120 125.250 36.380 125.570 ;
        RECT 35.660 120.830 35.920 121.150 ;
        RECT 34.280 120.490 34.540 120.810 ;
        RECT 33.420 119.730 34.020 119.870 ;
        RECT 34.740 119.810 35.000 120.130 ;
        RECT 33.420 116.390 33.560 119.730 ;
        RECT 33.820 117.770 34.080 118.090 ;
        RECT 32.900 116.070 33.160 116.390 ;
        RECT 33.360 116.070 33.620 116.390 ;
        RECT 31.520 115.730 31.780 116.050 ;
        RECT 31.060 115.390 31.320 115.710 ;
        RECT 30.600 113.010 30.860 113.330 ;
        RECT 31.120 112.650 31.260 115.390 ;
        RECT 31.580 113.330 31.720 115.730 ;
        RECT 31.980 115.050 32.240 115.370 ;
        RECT 31.520 113.010 31.780 113.330 ;
        RECT 32.040 112.990 32.180 115.050 ;
        RECT 32.960 115.030 33.100 116.070 ;
        RECT 32.900 114.710 33.160 115.030 ;
        RECT 31.980 112.670 32.240 112.990 ;
        RECT 32.960 112.650 33.100 114.710 ;
        RECT 31.060 112.330 31.320 112.650 ;
        RECT 32.900 112.330 33.160 112.650 ;
        RECT 33.420 112.310 33.560 116.070 ;
        RECT 33.360 111.990 33.620 112.310 ;
        RECT 30.600 111.650 30.860 111.970 ;
        RECT 30.660 108.230 30.800 111.650 ;
        RECT 30.950 111.115 32.490 111.485 ;
        RECT 32.900 109.610 33.160 109.930 ;
        RECT 31.060 109.270 31.320 109.590 ;
        RECT 30.600 107.910 30.860 108.230 ;
        RECT 30.140 107.230 30.400 107.550 ;
        RECT 30.200 104.830 30.340 107.230 ;
        RECT 31.120 107.210 31.260 109.270 ;
        RECT 32.440 107.230 32.700 107.550 ;
        RECT 31.060 106.890 31.320 107.210 ;
        RECT 32.500 107.065 32.640 107.230 ;
        RECT 32.430 106.695 32.710 107.065 ;
        RECT 30.950 105.675 32.490 106.045 ;
        RECT 32.960 105.510 33.100 109.610 ;
        RECT 33.880 107.210 34.020 117.770 ;
        RECT 34.800 116.050 34.940 119.810 ;
        RECT 35.720 118.430 35.860 120.830 ;
        RECT 35.660 118.110 35.920 118.430 ;
        RECT 34.740 115.730 35.000 116.050 ;
        RECT 35.660 115.730 35.920 116.050 ;
        RECT 35.720 115.110 35.860 115.730 ;
        RECT 36.180 115.710 36.320 125.250 ;
        RECT 36.120 115.390 36.380 115.710 ;
        RECT 35.720 114.970 36.320 115.110 ;
        RECT 34.740 114.370 35.000 114.690 ;
        RECT 35.660 114.370 35.920 114.690 ;
        RECT 34.800 107.210 34.940 114.370 ;
        RECT 33.350 106.695 33.630 107.065 ;
        RECT 33.820 106.890 34.080 107.210 ;
        RECT 34.740 106.890 35.000 107.210 ;
        RECT 35.720 106.870 35.860 114.370 ;
        RECT 36.180 113.750 36.320 114.970 ;
        RECT 36.180 113.610 36.780 113.750 ;
        RECT 30.600 105.190 30.860 105.510 ;
        RECT 32.900 105.190 33.160 105.510 ;
        RECT 30.140 104.510 30.400 104.830 ;
        RECT 30.140 103.490 30.400 103.810 ;
        RECT 23.240 97.030 23.500 97.350 ;
        RECT 29.680 97.030 29.940 97.350 ;
        RECT 23.300 96.330 23.440 97.030 ;
        RECT 23.760 96.610 24.820 96.750 ;
        RECT 25.540 96.690 25.800 97.010 ;
        RECT 23.760 96.330 23.900 96.610 ;
        RECT 23.240 96.010 23.500 96.330 ;
        RECT 23.700 96.010 23.960 96.330 ;
        RECT 23.300 90.210 23.440 96.010 ;
        RECT 24.160 95.670 24.420 95.990 ;
        RECT 23.700 95.330 23.960 95.650 ;
        RECT 23.240 89.890 23.500 90.210 ;
        RECT 23.300 88.850 23.440 89.890 ;
        RECT 23.240 88.530 23.500 88.850 ;
        RECT 22.380 86.240 22.980 86.380 ;
        RECT 21.860 85.810 22.120 86.130 ;
        RECT 22.380 85.305 22.520 86.240 ;
        RECT 22.770 85.615 23.050 85.985 ;
        RECT 22.310 84.935 22.590 85.305 ;
        RECT 22.380 84.770 22.520 84.935 ;
        RECT 22.320 84.450 22.580 84.770 ;
        RECT 22.380 78.310 22.520 84.450 ;
        RECT 22.840 79.240 22.980 85.615 ;
        RECT 23.240 85.470 23.500 85.790 ;
        RECT 23.300 80.010 23.440 85.470 ;
        RECT 23.760 85.450 23.900 95.330 ;
        RECT 24.220 93.950 24.360 95.670 ;
        RECT 24.160 93.630 24.420 93.950 ;
        RECT 24.160 89.890 24.420 90.210 ;
        RECT 24.220 89.190 24.360 89.890 ;
        RECT 24.160 88.870 24.420 89.190 ;
        RECT 24.680 88.510 24.820 96.610 ;
        RECT 25.600 96.330 25.740 96.690 ;
        RECT 25.540 96.010 25.800 96.330 ;
        RECT 26.000 96.185 26.260 96.330 ;
        RECT 25.990 95.815 26.270 96.185 ;
        RECT 25.080 93.630 25.340 93.950 ;
        RECT 25.140 91.910 25.280 93.630 ;
        RECT 25.540 92.610 25.800 92.930 ;
        RECT 25.080 91.590 25.340 91.910 ;
        RECT 25.600 90.890 25.740 92.610 ;
        RECT 25.540 90.570 25.800 90.890 ;
        RECT 24.620 88.190 24.880 88.510 ;
        RECT 24.680 87.830 24.820 88.190 ;
        RECT 26.060 88.080 26.200 95.815 ;
        RECT 26.920 95.670 27.180 95.990 ;
        RECT 26.980 92.930 27.120 95.670 ;
        RECT 26.920 92.610 27.180 92.930 ;
        RECT 26.980 90.890 27.120 92.610 ;
        RECT 27.650 92.075 29.190 92.445 ;
        RECT 29.740 90.890 29.880 97.030 ;
        RECT 30.200 91.230 30.340 103.490 ;
        RECT 30.140 90.910 30.400 91.230 ;
        RECT 26.920 90.570 27.180 90.890 ;
        RECT 27.840 90.570 28.100 90.890 ;
        RECT 29.680 90.570 29.940 90.890 ;
        RECT 26.460 90.230 26.720 90.550 ;
        RECT 26.520 89.190 26.660 90.230 ;
        RECT 26.460 88.870 26.720 89.190 ;
        RECT 26.980 88.510 27.120 90.570 ;
        RECT 27.380 89.890 27.640 90.210 ;
        RECT 26.920 88.190 27.180 88.510 ;
        RECT 26.460 88.080 26.720 88.170 ;
        RECT 26.060 87.940 26.720 88.080 ;
        RECT 24.620 87.510 24.880 87.830 ;
        RECT 24.680 86.130 24.820 87.510 ;
        RECT 26.060 86.470 26.200 87.940 ;
        RECT 26.460 87.850 26.720 87.940 ;
        RECT 27.440 87.910 27.580 89.890 ;
        RECT 27.900 88.510 28.040 90.570 ;
        RECT 30.140 90.230 30.400 90.550 ;
        RECT 29.220 89.890 29.480 90.210 ;
        RECT 27.840 88.190 28.100 88.510 ;
        RECT 28.300 88.190 28.560 88.510 ;
        RECT 26.980 87.770 27.580 87.910 ;
        RECT 28.360 87.830 28.500 88.190 ;
        RECT 26.000 86.150 26.260 86.470 ;
        RECT 26.980 86.380 27.120 87.770 ;
        RECT 28.300 87.510 28.560 87.830 ;
        RECT 29.280 87.490 29.420 89.890 ;
        RECT 29.680 88.870 29.940 89.190 ;
        RECT 29.220 87.170 29.480 87.490 ;
        RECT 29.740 87.230 29.880 88.870 ;
        RECT 30.200 88.510 30.340 90.230 ;
        RECT 30.140 88.190 30.400 88.510 ;
        RECT 29.740 87.090 30.340 87.230 ;
        RECT 27.650 86.635 29.190 87.005 ;
        RECT 26.980 86.240 27.580 86.380 ;
        RECT 24.620 85.810 24.880 86.130 ;
        RECT 26.060 85.450 26.200 86.150 ;
        RECT 23.700 85.130 23.960 85.450 ;
        RECT 26.000 85.130 26.260 85.450 ;
        RECT 26.920 85.305 27.180 85.450 ;
        RECT 25.080 84.790 25.340 85.110 ;
        RECT 26.910 84.935 27.190 85.305 ;
        RECT 25.140 83.750 25.280 84.790 ;
        RECT 26.000 84.450 26.260 84.770 ;
        RECT 26.460 84.450 26.720 84.770 ;
        RECT 25.080 83.430 25.340 83.750 ;
        RECT 23.240 79.690 23.500 80.010 ;
        RECT 22.840 79.100 23.440 79.240 ;
        RECT 22.320 77.990 22.580 78.310 ;
        RECT 22.320 74.930 22.580 75.250 ;
        RECT 21.860 74.250 22.120 74.570 ;
        RECT 21.920 69.810 22.060 74.250 ;
        RECT 22.380 72.190 22.520 74.930 ;
        RECT 22.780 73.910 23.040 74.230 ;
        RECT 22.320 71.870 22.580 72.190 ;
        RECT 22.320 70.850 22.580 71.170 ;
        RECT 21.860 69.490 22.120 69.810 ;
        RECT 22.380 68.450 22.520 70.850 ;
        RECT 22.840 70.150 22.980 73.910 ;
        RECT 22.780 69.830 23.040 70.150 ;
        RECT 22.320 68.130 22.580 68.450 ;
        RECT 23.300 67.510 23.440 79.100 ;
        RECT 23.700 79.010 23.960 79.330 ;
        RECT 23.760 75.105 23.900 79.010 ;
        RECT 24.610 77.455 24.890 77.825 ;
        RECT 25.540 77.650 25.800 77.970 ;
        RECT 24.620 77.310 24.880 77.455 ;
        RECT 24.620 76.860 24.880 76.950 ;
        RECT 24.220 76.720 24.880 76.860 ;
        RECT 23.690 74.735 23.970 75.105 ;
        RECT 24.220 74.310 24.360 76.720 ;
        RECT 24.620 76.630 24.880 76.720 ;
        RECT 24.610 76.095 24.890 76.465 ;
        RECT 25.080 76.290 25.340 76.610 ;
        RECT 24.680 74.570 24.820 76.095 ;
        RECT 23.760 74.230 24.360 74.310 ;
        RECT 24.620 74.250 24.880 74.570 ;
        RECT 23.700 74.170 24.360 74.230 ;
        RECT 23.700 73.910 23.960 74.170 ;
        RECT 24.160 73.570 24.420 73.890 ;
        RECT 23.700 71.080 23.960 71.170 ;
        RECT 24.220 71.080 24.360 73.570 ;
        RECT 24.680 71.590 24.820 74.250 ;
        RECT 25.140 72.190 25.280 76.290 ;
        RECT 25.600 72.870 25.740 77.650 ;
        RECT 26.060 75.105 26.200 84.450 ;
        RECT 26.520 76.610 26.660 84.450 ;
        RECT 27.440 82.300 27.580 86.240 ;
        RECT 29.680 86.150 29.940 86.470 ;
        RECT 26.980 82.160 27.580 82.300 ;
        RECT 26.980 80.350 27.120 82.160 ;
        RECT 27.650 81.195 29.190 81.565 ;
        RECT 26.920 80.030 27.180 80.350 ;
        RECT 26.980 77.290 27.120 80.030 ;
        RECT 29.740 80.010 29.880 86.150 ;
        RECT 30.200 83.070 30.340 87.090 ;
        RECT 30.660 86.470 30.800 105.190 ;
        RECT 32.430 104.655 32.710 105.025 ;
        RECT 32.440 104.510 32.700 104.655 ;
        RECT 30.950 100.235 32.490 100.605 ;
        RECT 31.520 99.070 31.780 99.390 ;
        RECT 32.440 99.070 32.700 99.390 ;
        RECT 31.580 96.330 31.720 99.070 ;
        RECT 32.500 96.330 32.640 99.070 ;
        RECT 33.420 97.350 33.560 106.695 ;
        RECT 35.660 106.550 35.920 106.870 ;
        RECT 35.720 104.830 35.860 106.550 ;
        RECT 36.120 106.210 36.380 106.530 ;
        RECT 36.180 105.170 36.320 106.210 ;
        RECT 36.120 104.850 36.380 105.170 ;
        RECT 36.640 105.025 36.780 113.610 ;
        RECT 37.100 109.930 37.240 128.310 ;
        RECT 38.020 128.290 38.160 131.030 ;
        RECT 37.500 127.970 37.760 128.290 ;
        RECT 37.960 127.970 38.220 128.290 ;
        RECT 37.560 123.530 37.700 127.970 ;
        RECT 38.020 125.570 38.160 127.970 ;
        RECT 37.960 125.250 38.220 125.570 ;
        RECT 37.500 123.210 37.760 123.530 ;
        RECT 38.420 123.210 38.680 123.530 ;
        RECT 37.960 120.490 38.220 120.810 ;
        RECT 37.500 120.150 37.760 120.470 ;
        RECT 37.560 116.050 37.700 120.150 ;
        RECT 37.500 115.730 37.760 116.050 ;
        RECT 38.020 113.330 38.160 120.490 ;
        RECT 38.480 118.770 38.620 123.210 ;
        RECT 38.880 120.830 39.140 121.150 ;
        RECT 38.420 118.450 38.680 118.770 ;
        RECT 38.480 118.090 38.620 118.450 ;
        RECT 38.420 117.770 38.680 118.090 ;
        RECT 38.480 113.330 38.620 117.770 ;
        RECT 37.960 113.010 38.220 113.330 ;
        RECT 38.420 113.010 38.680 113.330 ;
        RECT 37.040 109.610 37.300 109.930 ;
        RECT 38.020 108.230 38.160 113.010 ;
        RECT 38.940 112.650 39.080 120.830 ;
        RECT 39.860 115.710 40.000 134.430 ;
        RECT 42.620 134.410 42.760 136.470 ;
        RECT 42.560 134.090 42.820 134.410 ;
        RECT 42.100 131.710 42.360 132.030 ;
        RECT 42.160 129.990 42.300 131.710 ;
        RECT 42.100 129.670 42.360 129.990 ;
        RECT 43.540 129.310 43.680 145.990 ;
        RECT 43.940 141.570 44.200 141.890 ;
        RECT 43.480 128.990 43.740 129.310 ;
        RECT 41.180 122.530 41.440 122.850 ;
        RECT 40.720 117.770 40.980 118.090 ;
        RECT 40.260 117.090 40.520 117.410 ;
        RECT 39.800 115.390 40.060 115.710 ;
        RECT 39.340 114.370 39.600 114.690 ;
        RECT 38.880 112.330 39.140 112.650 ;
        RECT 38.940 110.950 39.080 112.330 ;
        RECT 38.880 110.630 39.140 110.950 ;
        RECT 37.960 107.910 38.220 108.230 ;
        RECT 38.940 105.510 39.080 110.630 ;
        RECT 38.880 105.190 39.140 105.510 ;
        RECT 35.660 104.510 35.920 104.830 ;
        RECT 36.570 104.655 36.850 105.025 ;
        RECT 39.400 103.810 39.540 114.370 ;
        RECT 39.860 109.590 40.000 115.390 ;
        RECT 40.320 112.990 40.460 117.090 ;
        RECT 40.780 116.050 40.920 117.770 ;
        RECT 40.720 115.730 40.980 116.050 ;
        RECT 41.240 115.710 41.380 122.530 ;
        RECT 41.640 117.430 41.900 117.750 ;
        RECT 41.700 116.050 41.840 117.430 ;
        RECT 41.640 115.730 41.900 116.050 ;
        RECT 41.180 115.390 41.440 115.710 ;
        RECT 43.020 113.350 43.280 113.670 ;
        RECT 40.260 112.670 40.520 112.990 ;
        RECT 43.080 110.610 43.220 113.350 ;
        RECT 43.020 110.290 43.280 110.610 ;
        RECT 39.800 109.270 40.060 109.590 ;
        RECT 41.180 104.170 41.440 104.490 ;
        RECT 39.340 103.490 39.600 103.810 ;
        RECT 39.800 103.490 40.060 103.810 ;
        RECT 36.580 100.770 36.840 101.090 ;
        RECT 36.640 99.390 36.780 100.770 ;
        RECT 39.860 99.390 40.000 103.490 ;
        RECT 41.240 101.770 41.380 104.170 ;
        RECT 41.180 101.450 41.440 101.770 ;
        RECT 41.240 99.390 41.380 101.450 ;
        RECT 41.640 101.110 41.900 101.430 ;
        RECT 41.700 99.730 41.840 101.110 ;
        RECT 42.100 100.770 42.360 101.090 ;
        RECT 41.640 99.410 41.900 99.730 ;
        RECT 36.580 99.070 36.840 99.390 ;
        RECT 39.800 99.070 40.060 99.390 ;
        RECT 41.180 99.070 41.440 99.390 ;
        RECT 33.360 97.030 33.620 97.350 ;
        RECT 31.520 96.010 31.780 96.330 ;
        RECT 32.440 96.010 32.700 96.330 ;
        RECT 32.500 95.650 32.640 96.010 ;
        RECT 32.440 95.330 32.700 95.650 ;
        RECT 30.950 94.795 32.490 95.165 ;
        RECT 33.420 94.710 33.560 97.030 ;
        RECT 37.040 95.330 37.300 95.650 ;
        RECT 33.420 94.570 34.020 94.710 ;
        RECT 31.980 93.970 32.240 94.290 ;
        RECT 33.360 93.970 33.620 94.290 ;
        RECT 32.040 91.230 32.180 93.970 ;
        RECT 32.900 92.610 33.160 92.930 ;
        RECT 32.960 91.910 33.100 92.610 ;
        RECT 32.900 91.590 33.160 91.910 ;
        RECT 31.980 90.910 32.240 91.230 ;
        RECT 32.900 90.910 33.160 91.230 ;
        RECT 30.950 89.355 32.490 89.725 ;
        RECT 31.980 88.530 32.240 88.850 ;
        RECT 31.520 87.510 31.780 87.830 ;
        RECT 31.060 87.170 31.320 87.490 ;
        RECT 30.600 86.150 30.860 86.470 ;
        RECT 31.120 85.870 31.260 87.170 ;
        RECT 30.660 85.790 31.260 85.870 ;
        RECT 30.600 85.730 31.260 85.790 ;
        RECT 30.600 85.470 30.860 85.730 ;
        RECT 30.140 82.750 30.400 83.070 ;
        RECT 30.140 81.730 30.400 82.050 ;
        RECT 28.300 79.690 28.560 80.010 ;
        RECT 29.680 79.690 29.940 80.010 ;
        RECT 27.840 79.010 28.100 79.330 ;
        RECT 27.900 77.630 28.040 79.010 ;
        RECT 27.840 77.310 28.100 77.630 ;
        RECT 26.920 76.970 27.180 77.290 ;
        RECT 28.360 76.950 28.500 79.690 ;
        RECT 29.680 79.010 29.940 79.330 ;
        RECT 28.760 77.310 29.020 77.630 ;
        RECT 28.300 76.630 28.560 76.950 ;
        RECT 28.820 76.610 28.960 77.310 ;
        RECT 26.460 76.290 26.720 76.610 ;
        RECT 26.920 76.290 27.180 76.610 ;
        RECT 28.760 76.290 29.020 76.610 ;
        RECT 25.990 74.735 26.270 75.105 ;
        RECT 25.540 72.550 25.800 72.870 ;
        RECT 26.520 72.190 26.660 76.290 ;
        RECT 25.080 71.870 25.340 72.190 ;
        RECT 26.460 71.870 26.720 72.190 ;
        RECT 24.680 71.450 25.280 71.590 ;
        RECT 26.000 71.530 26.260 71.850 ;
        RECT 23.700 70.940 24.360 71.080 ;
        RECT 23.700 70.850 23.960 70.940 ;
        RECT 24.620 70.850 24.880 71.170 ;
        RECT 23.690 69.380 23.970 69.665 ;
        RECT 23.690 69.295 24.360 69.380 ;
        RECT 23.700 69.240 24.360 69.295 ;
        RECT 23.700 69.150 23.960 69.240 ;
        RECT 22.840 67.370 23.440 67.510 ;
        RECT 22.840 67.090 22.980 67.370 ;
        RECT 22.320 66.770 22.580 67.090 ;
        RECT 22.780 66.770 23.040 67.090 ;
        RECT 21.460 66.010 22.060 66.150 ;
        RECT 21.920 65.730 22.060 66.010 ;
        RECT 21.400 65.470 21.660 65.730 ;
        RECT 21.000 65.410 21.660 65.470 ;
        RECT 21.860 65.410 22.120 65.730 ;
        RECT 21.000 65.330 21.600 65.410 ;
        RECT 22.380 64.710 22.520 66.770 ;
        RECT 20.480 64.390 20.740 64.710 ;
        RECT 22.320 64.390 22.580 64.710 ;
        RECT 20.480 63.370 20.740 63.690 ;
        RECT 19.560 62.690 19.820 63.010 ;
        RECT 19.620 61.650 19.760 62.690 ;
        RECT 19.560 61.330 19.820 61.650 ;
        RECT 18.180 60.990 18.440 61.310 ;
        RECT 18.240 53.150 18.380 60.990 ;
        RECT 20.540 58.590 20.680 63.370 ;
        RECT 22.320 63.030 22.580 63.350 ;
        RECT 20.480 58.270 20.740 58.590 ;
        RECT 18.180 52.830 18.440 53.150 ;
        RECT 18.240 52.550 18.380 52.830 ;
        RECT 16.800 52.380 17.060 52.470 ;
        RECT 18.240 52.410 18.840 52.550 ;
        RECT 16.800 52.240 17.920 52.380 ;
        RECT 16.800 52.150 17.060 52.240 ;
        RECT 15.940 47.650 16.540 47.790 ;
        RECT 15.880 47.280 16.140 47.370 ;
        RECT 15.480 47.140 16.140 47.280 ;
        RECT 15.880 47.050 16.140 47.140 ;
        RECT 15.020 44.990 15.160 47.050 ;
        RECT 14.500 44.670 14.760 44.990 ;
        RECT 14.960 44.670 15.220 44.990 ;
        RECT 16.400 43.970 16.540 47.650 ;
        RECT 17.780 44.990 17.920 52.240 ;
        RECT 18.180 51.810 18.440 52.130 ;
        RECT 18.240 51.110 18.380 51.810 ;
        RECT 18.180 50.790 18.440 51.110 ;
        RECT 18.700 50.770 18.840 52.410 ;
        RECT 18.640 50.450 18.900 50.770 ;
        RECT 18.700 47.030 18.840 50.450 ;
        RECT 20.540 50.430 20.680 58.270 ;
        RECT 21.400 55.210 21.660 55.530 ;
        RECT 21.460 52.470 21.600 55.210 ;
        RECT 22.380 52.810 22.520 63.030 ;
        RECT 22.840 61.990 22.980 66.770 ;
        RECT 24.220 66.750 24.360 69.240 ;
        RECT 23.700 66.430 23.960 66.750 ;
        RECT 24.160 66.430 24.420 66.750 ;
        RECT 23.760 65.730 23.900 66.430 ;
        RECT 23.700 65.410 23.960 65.730 ;
        RECT 24.160 65.410 24.420 65.730 ;
        RECT 22.780 61.670 23.040 61.990 ;
        RECT 22.840 59.270 22.980 61.670 ;
        RECT 23.760 60.630 23.900 65.410 ;
        RECT 24.220 61.310 24.360 65.410 ;
        RECT 24.160 60.990 24.420 61.310 ;
        RECT 23.700 60.310 23.960 60.630 ;
        RECT 22.780 58.950 23.040 59.270 ;
        RECT 24.680 58.250 24.820 70.850 ;
        RECT 23.240 57.930 23.500 58.250 ;
        RECT 24.620 57.930 24.880 58.250 ;
        RECT 23.300 56.550 23.440 57.930 ;
        RECT 23.240 56.230 23.500 56.550 ;
        RECT 23.240 55.550 23.500 55.870 ;
        RECT 22.320 52.490 22.580 52.810 ;
        RECT 21.400 52.150 21.660 52.470 ;
        RECT 20.940 51.810 21.200 52.130 ;
        RECT 21.000 50.770 21.140 51.810 ;
        RECT 20.940 50.450 21.200 50.770 ;
        RECT 19.100 50.110 19.360 50.430 ;
        RECT 20.480 50.110 20.740 50.430 ;
        RECT 18.640 46.710 18.900 47.030 ;
        RECT 17.720 44.670 17.980 44.990 ;
        RECT 16.340 43.650 16.600 43.970 ;
        RECT 17.780 41.590 17.920 44.670 ;
        RECT 18.180 43.650 18.440 43.970 ;
        RECT 18.240 42.950 18.380 43.650 ;
        RECT 18.180 42.630 18.440 42.950 ;
        RECT 18.700 42.610 18.840 46.710 ;
        RECT 18.640 42.290 18.900 42.610 ;
        RECT 18.180 41.950 18.440 42.270 ;
        RECT 18.240 41.590 18.380 41.950 ;
        RECT 17.720 41.270 17.980 41.590 ;
        RECT 18.180 41.270 18.440 41.590 ;
        RECT 19.160 41.250 19.300 50.110 ;
        RECT 20.540 48.390 20.680 50.110 ;
        RECT 21.000 48.390 21.140 50.450 ;
        RECT 21.400 49.430 21.660 49.750 ;
        RECT 20.480 48.070 20.740 48.390 ;
        RECT 20.940 48.070 21.200 48.390 ;
        RECT 19.560 47.730 19.820 48.050 ;
        RECT 19.620 41.250 19.760 47.730 ;
        RECT 20.540 42.270 20.680 48.070 ;
        RECT 20.940 46.370 21.200 46.690 ;
        RECT 20.480 41.950 20.740 42.270 ;
        RECT 21.000 41.930 21.140 46.370 ;
        RECT 21.460 45.670 21.600 49.430 ;
        RECT 22.380 49.410 22.520 52.490 ;
        RECT 23.300 52.130 23.440 55.550 ;
        RECT 24.620 55.210 24.880 55.530 ;
        RECT 24.680 53.830 24.820 55.210 ;
        RECT 24.620 53.510 24.880 53.830 ;
        RECT 25.140 53.150 25.280 71.450 ;
        RECT 26.060 70.110 26.200 71.530 ;
        RECT 25.600 69.970 26.200 70.110 ;
        RECT 25.600 65.470 25.740 69.970 ;
        RECT 26.000 68.470 26.260 68.790 ;
        RECT 26.060 66.070 26.200 68.470 ;
        RECT 26.460 68.130 26.720 68.450 ;
        RECT 26.520 67.430 26.660 68.130 ;
        RECT 26.460 67.110 26.720 67.430 ;
        RECT 26.460 66.430 26.720 66.750 ;
        RECT 26.000 65.750 26.260 66.070 ;
        RECT 26.520 65.470 26.660 66.430 ;
        RECT 25.600 65.330 26.660 65.470 ;
        RECT 25.600 63.350 25.740 65.330 ;
        RECT 25.540 63.030 25.800 63.350 ;
        RECT 26.980 61.310 27.120 76.290 ;
        RECT 27.650 75.755 29.190 76.125 ;
        RECT 27.840 75.105 28.100 75.250 ;
        RECT 27.830 74.735 28.110 75.105 ;
        RECT 27.840 74.425 28.100 74.570 ;
        RECT 27.830 74.055 28.110 74.425 ;
        RECT 27.380 73.570 27.640 73.890 ;
        RECT 27.440 72.190 27.580 73.570 ;
        RECT 27.380 71.870 27.640 72.190 ;
        RECT 27.650 70.315 29.190 70.685 ;
        RECT 29.740 70.110 29.880 79.010 ;
        RECT 30.200 71.170 30.340 81.730 ;
        RECT 30.660 79.670 30.800 85.470 ;
        RECT 31.580 85.450 31.720 87.510 ;
        RECT 31.060 85.305 31.320 85.450 ;
        RECT 31.050 84.935 31.330 85.305 ;
        RECT 31.520 85.130 31.780 85.450 ;
        RECT 32.040 85.305 32.180 88.530 ;
        RECT 32.430 85.615 32.710 85.985 ;
        RECT 32.500 85.450 32.640 85.615 ;
        RECT 31.970 84.935 32.250 85.305 ;
        RECT 32.440 85.130 32.700 85.450 ;
        RECT 30.950 83.915 32.490 84.285 ;
        RECT 31.060 83.430 31.320 83.750 ;
        RECT 31.120 80.350 31.260 83.430 ;
        RECT 32.440 82.750 32.700 83.070 ;
        RECT 31.060 80.030 31.320 80.350 ;
        RECT 30.600 79.350 30.860 79.670 ;
        RECT 30.660 77.825 30.800 79.350 ;
        RECT 32.500 79.330 32.640 82.750 ;
        RECT 32.960 80.010 33.100 90.910 ;
        RECT 33.420 86.470 33.560 93.970 ;
        RECT 33.360 86.150 33.620 86.470 ;
        RECT 33.880 85.790 34.020 94.570 ;
        RECT 34.740 93.630 35.000 93.950 ;
        RECT 36.120 93.630 36.380 93.950 ;
        RECT 34.280 92.610 34.540 92.930 ;
        RECT 34.340 90.890 34.480 92.610 ;
        RECT 34.280 90.570 34.540 90.890 ;
        RECT 34.800 88.850 34.940 93.630 ;
        RECT 35.200 93.290 35.460 93.610 ;
        RECT 35.260 88.850 35.400 93.290 ;
        RECT 35.660 92.610 35.920 92.930 ;
        RECT 34.740 88.530 35.000 88.850 ;
        RECT 35.200 88.530 35.460 88.850 ;
        RECT 34.280 87.510 34.540 87.830 ;
        RECT 35.200 87.510 35.460 87.830 ;
        RECT 33.820 85.470 34.080 85.790 ;
        RECT 33.820 83.090 34.080 83.410 ;
        RECT 33.880 80.010 34.020 83.090 ;
        RECT 34.340 83.070 34.480 87.510 ;
        RECT 34.740 87.170 35.000 87.490 ;
        RECT 34.800 86.470 34.940 87.170 ;
        RECT 34.740 86.150 35.000 86.470 ;
        RECT 34.800 85.450 34.940 86.150 ;
        RECT 34.740 85.130 35.000 85.450 ;
        RECT 34.280 82.750 34.540 83.070 ;
        RECT 34.800 81.030 34.940 85.130 ;
        RECT 35.260 83.750 35.400 87.510 ;
        RECT 35.720 87.490 35.860 92.610 ;
        RECT 36.180 91.910 36.320 93.630 ;
        RECT 36.120 91.590 36.380 91.910 ;
        RECT 36.180 89.190 36.320 91.590 ;
        RECT 36.580 90.230 36.840 90.550 ;
        RECT 36.640 89.190 36.780 90.230 ;
        RECT 36.120 88.870 36.380 89.190 ;
        RECT 36.580 88.870 36.840 89.190 ;
        RECT 35.660 87.170 35.920 87.490 ;
        RECT 36.180 85.450 36.320 88.870 ;
        RECT 36.120 85.130 36.380 85.450 ;
        RECT 35.660 84.790 35.920 85.110 ;
        RECT 35.720 84.625 35.860 84.790 ;
        RECT 35.650 84.255 35.930 84.625 ;
        RECT 35.200 83.660 35.460 83.750 ;
        RECT 35.200 83.520 36.320 83.660 ;
        RECT 35.200 83.430 35.460 83.520 ;
        RECT 34.740 80.710 35.000 81.030 ;
        RECT 32.900 79.690 33.160 80.010 ;
        RECT 33.820 79.690 34.080 80.010 ;
        RECT 32.440 79.010 32.700 79.330 ;
        RECT 30.950 78.475 32.490 78.845 ;
        RECT 32.440 77.990 32.700 78.310 ;
        RECT 30.590 77.455 30.870 77.825 ;
        RECT 32.500 77.630 32.640 77.990 ;
        RECT 32.440 77.310 32.700 77.630 ;
        RECT 31.060 76.630 31.320 76.950 ;
        RECT 30.600 75.270 30.860 75.590 ;
        RECT 30.140 70.850 30.400 71.170 ;
        RECT 29.740 69.970 30.340 70.110 ;
        RECT 29.680 68.810 29.940 69.130 ;
        RECT 27.370 67.935 27.650 68.305 ;
        RECT 28.760 68.130 29.020 68.450 ;
        RECT 27.440 66.750 27.580 67.935 ;
        RECT 28.820 67.430 28.960 68.130 ;
        RECT 28.760 67.110 29.020 67.430 ;
        RECT 27.380 66.430 27.640 66.750 ;
        RECT 29.740 66.150 29.880 68.810 ;
        RECT 30.200 66.750 30.340 69.970 ;
        RECT 30.660 69.130 30.800 75.270 ;
        RECT 31.120 74.910 31.260 76.630 ;
        RECT 31.060 74.590 31.320 74.910 ;
        RECT 32.500 74.310 32.640 77.310 ;
        RECT 32.960 75.590 33.100 79.690 ;
        RECT 33.880 78.310 34.020 79.690 ;
        RECT 34.280 79.010 34.540 79.330 ;
        RECT 34.740 79.010 35.000 79.330 ;
        RECT 33.820 77.990 34.080 78.310 ;
        RECT 33.360 76.290 33.620 76.610 ;
        RECT 32.900 75.270 33.160 75.590 ;
        RECT 32.960 74.910 33.100 75.270 ;
        RECT 32.900 74.590 33.160 74.910 ;
        RECT 32.500 74.170 33.100 74.310 ;
        RECT 30.950 73.035 32.490 73.405 ;
        RECT 31.050 72.015 31.330 72.385 ;
        RECT 31.120 71.510 31.260 72.015 ;
        RECT 31.520 71.870 31.780 72.190 ;
        RECT 31.060 71.190 31.320 71.510 ;
        RECT 30.600 68.810 30.860 69.130 ;
        RECT 30.660 67.090 30.800 68.810 ;
        RECT 31.120 68.790 31.260 71.190 ;
        RECT 31.580 70.345 31.720 71.870 ;
        RECT 31.510 69.975 31.790 70.345 ;
        RECT 32.440 70.060 32.700 70.150 ;
        RECT 32.960 70.060 33.100 74.170 ;
        RECT 33.420 71.850 33.560 76.290 ;
        RECT 34.340 72.190 34.480 79.010 ;
        RECT 34.800 72.190 34.940 79.010 ;
        RECT 35.200 77.310 35.460 77.630 ;
        RECT 35.260 72.870 35.400 77.310 ;
        RECT 35.660 76.290 35.920 76.610 ;
        RECT 35.720 72.870 35.860 76.290 ;
        RECT 35.200 72.550 35.460 72.870 ;
        RECT 35.660 72.550 35.920 72.870 ;
        RECT 36.180 72.190 36.320 83.520 ;
        RECT 37.100 83.150 37.240 95.330 ;
        RECT 37.960 93.970 38.220 94.290 ;
        RECT 38.020 90.210 38.160 93.970 ;
        RECT 42.160 92.930 42.300 100.770 ;
        RECT 43.480 99.410 43.740 99.730 ;
        RECT 43.540 97.350 43.680 99.410 ;
        RECT 43.480 97.030 43.740 97.350 ;
        RECT 42.100 92.610 42.360 92.930 ;
        RECT 37.960 89.890 38.220 90.210 ;
        RECT 38.020 86.470 38.160 89.890 ;
        RECT 38.880 88.530 39.140 88.850 ;
        RECT 37.960 86.150 38.220 86.470 ;
        RECT 38.020 85.450 38.160 86.150 ;
        RECT 37.960 85.130 38.220 85.450 ;
        RECT 37.500 84.790 37.760 85.110 ;
        RECT 37.560 83.750 37.700 84.790 ;
        RECT 38.420 84.450 38.680 84.770 ;
        RECT 37.500 83.430 37.760 83.750 ;
        RECT 36.580 82.750 36.840 83.070 ;
        RECT 37.100 83.010 38.160 83.150 ;
        RECT 36.640 79.330 36.780 82.750 ;
        RECT 38.020 80.690 38.160 83.010 ;
        RECT 38.480 82.730 38.620 84.450 ;
        RECT 38.420 82.410 38.680 82.730 ;
        RECT 37.960 80.370 38.220 80.690 ;
        RECT 37.040 79.690 37.300 80.010 ;
        RECT 37.500 79.690 37.760 80.010 ;
        RECT 36.580 79.010 36.840 79.330 ;
        RECT 36.640 74.910 36.780 79.010 ;
        RECT 36.580 74.590 36.840 74.910 ;
        RECT 34.280 71.870 34.540 72.190 ;
        RECT 34.740 71.870 35.000 72.190 ;
        RECT 35.200 71.870 35.460 72.190 ;
        RECT 36.120 71.870 36.380 72.190 ;
        RECT 33.360 71.530 33.620 71.850 ;
        RECT 33.360 70.850 33.620 71.170 ;
        RECT 34.280 70.910 34.540 71.170 ;
        RECT 33.880 70.850 34.540 70.910 ;
        RECT 32.440 69.920 33.100 70.060 ;
        RECT 32.440 69.830 32.700 69.920 ;
        RECT 31.060 68.470 31.320 68.790 ;
        RECT 32.900 68.470 33.160 68.790 ;
        RECT 30.950 67.595 32.490 67.965 ;
        RECT 32.960 67.430 33.100 68.470 ;
        RECT 31.060 67.110 31.320 67.430 ;
        RECT 32.900 67.110 33.160 67.430 ;
        RECT 30.600 66.770 30.860 67.090 ;
        RECT 30.140 66.430 30.400 66.750 ;
        RECT 29.740 66.010 30.340 66.150 ;
        RECT 27.650 64.875 29.190 65.245 ;
        RECT 29.210 63.855 29.490 64.225 ;
        RECT 29.680 64.050 29.940 64.370 ;
        RECT 29.280 63.690 29.420 63.855 ;
        RECT 27.380 63.370 27.640 63.690 ;
        RECT 29.220 63.370 29.480 63.690 ;
        RECT 26.920 60.990 27.180 61.310 ;
        RECT 27.440 60.710 27.580 63.370 ;
        RECT 26.980 60.570 27.580 60.710 ;
        RECT 29.280 60.630 29.420 63.370 ;
        RECT 26.460 58.270 26.720 58.590 ;
        RECT 26.000 55.890 26.260 56.210 ;
        RECT 25.080 52.830 25.340 53.150 ;
        RECT 24.160 52.490 24.420 52.810 ;
        RECT 23.700 52.150 23.960 52.470 ;
        RECT 23.240 51.810 23.500 52.130 ;
        RECT 22.320 49.090 22.580 49.410 ;
        RECT 21.860 47.050 22.120 47.370 ;
        RECT 21.920 45.670 22.060 47.050 ;
        RECT 22.380 46.690 22.520 49.090 ;
        RECT 23.760 46.690 23.900 52.150 ;
        RECT 24.220 50.430 24.360 52.490 ;
        RECT 26.060 51.110 26.200 55.890 ;
        RECT 26.520 55.870 26.660 58.270 ;
        RECT 26.460 55.550 26.720 55.870 ;
        RECT 26.980 55.270 27.120 60.570 ;
        RECT 29.220 60.310 29.480 60.630 ;
        RECT 27.650 59.435 29.190 59.805 ;
        RECT 29.220 57.250 29.480 57.570 ;
        RECT 26.520 55.130 27.120 55.270 ;
        RECT 29.280 55.270 29.420 57.250 ;
        RECT 29.740 56.210 29.880 64.050 ;
        RECT 30.200 63.350 30.340 66.010 ;
        RECT 31.120 63.690 31.260 67.110 ;
        RECT 31.980 66.770 32.240 67.090 ;
        RECT 31.060 63.370 31.320 63.690 ;
        RECT 30.140 63.030 30.400 63.350 ;
        RECT 32.040 63.010 32.180 66.770 ;
        RECT 32.900 65.750 33.160 66.070 ;
        RECT 32.960 64.710 33.100 65.750 ;
        RECT 32.900 64.390 33.160 64.710 ;
        RECT 30.600 62.690 30.860 63.010 ;
        RECT 31.980 62.690 32.240 63.010 ;
        RECT 30.660 61.390 30.800 62.690 ;
        RECT 30.950 62.155 32.490 62.525 ;
        RECT 30.140 60.990 30.400 61.310 ;
        RECT 30.660 61.250 31.260 61.390 ;
        RECT 30.200 58.250 30.340 60.990 ;
        RECT 30.600 60.310 30.860 60.630 ;
        RECT 30.140 57.930 30.400 58.250 ;
        RECT 30.200 56.550 30.340 57.930 ;
        RECT 30.140 56.230 30.400 56.550 ;
        RECT 29.680 55.890 29.940 56.210 ;
        RECT 29.280 55.130 29.880 55.270 ;
        RECT 26.520 53.150 26.660 55.130 ;
        RECT 26.920 54.530 27.180 54.850 ;
        RECT 26.980 53.830 27.120 54.530 ;
        RECT 27.650 53.995 29.190 54.365 ;
        RECT 26.920 53.510 27.180 53.830 ;
        RECT 26.460 52.830 26.720 53.150 ;
        RECT 26.000 50.790 26.260 51.110 ;
        RECT 26.520 50.770 26.660 52.830 ;
        RECT 26.460 50.450 26.720 50.770 ;
        RECT 24.160 50.110 24.420 50.430 ;
        RECT 24.220 47.370 24.360 50.110 ;
        RECT 26.520 47.370 26.660 50.450 ;
        RECT 26.920 49.430 27.180 49.750 ;
        RECT 26.980 48.300 27.120 49.430 ;
        RECT 29.740 49.410 29.880 55.130 ;
        RECT 30.660 53.830 30.800 60.310 ;
        RECT 31.120 57.910 31.260 61.250 ;
        RECT 31.510 61.135 31.790 61.505 ;
        RECT 31.520 60.990 31.780 61.135 ;
        RECT 32.900 60.650 33.160 60.970 ;
        RECT 31.060 57.590 31.320 57.910 ;
        RECT 30.950 56.715 32.490 57.085 ;
        RECT 30.600 53.510 30.860 53.830 ;
        RECT 30.140 50.790 30.400 51.110 ;
        RECT 29.680 49.090 29.940 49.410 ;
        RECT 27.650 48.555 29.190 48.925 ;
        RECT 26.980 48.160 27.580 48.300 ;
        RECT 27.440 47.370 27.580 48.160 ;
        RECT 24.160 47.050 24.420 47.370 ;
        RECT 26.460 47.280 26.720 47.370 ;
        RECT 26.060 47.140 26.720 47.280 ;
        RECT 22.320 46.370 22.580 46.690 ;
        RECT 23.700 46.370 23.960 46.690 ;
        RECT 21.400 45.350 21.660 45.670 ;
        RECT 21.860 45.350 22.120 45.670 ;
        RECT 23.760 42.950 23.900 46.370 ;
        RECT 22.320 42.630 22.580 42.950 ;
        RECT 23.700 42.630 23.960 42.950 ;
        RECT 20.940 41.610 21.200 41.930 ;
        RECT 20.020 41.270 20.280 41.590 ;
        RECT 21.390 41.415 21.670 41.785 ;
        RECT 21.400 41.270 21.660 41.415 ;
        RECT 19.100 40.930 19.360 41.250 ;
        RECT 19.560 40.930 19.820 41.250 ;
        RECT 20.080 37.170 20.220 41.270 ;
        RECT 20.940 40.930 21.200 41.250 ;
        RECT 21.000 39.210 21.140 40.930 ;
        RECT 22.380 39.890 22.520 42.630 ;
        RECT 22.780 41.950 23.040 42.270 ;
        RECT 22.320 39.570 22.580 39.890 ;
        RECT 22.840 39.550 22.980 41.950 ;
        RECT 22.780 39.230 23.040 39.550 ;
        RECT 20.940 38.890 21.200 39.210 ;
        RECT 23.760 38.530 23.900 42.630 ;
        RECT 26.060 41.930 26.200 47.140 ;
        RECT 26.460 47.050 26.720 47.140 ;
        RECT 27.380 47.050 27.640 47.370 ;
        RECT 27.840 46.370 28.100 46.690 ;
        RECT 27.900 45.670 28.040 46.370 ;
        RECT 30.200 45.670 30.340 50.790 ;
        RECT 30.660 50.090 30.800 53.510 ;
        RECT 32.960 52.810 33.100 60.650 ;
        RECT 32.900 52.490 33.160 52.810 ;
        RECT 30.950 51.275 32.490 51.645 ;
        RECT 30.600 49.770 30.860 50.090 ;
        RECT 32.960 47.225 33.100 52.490 ;
        RECT 33.420 51.110 33.560 70.850 ;
        RECT 33.880 70.770 34.480 70.850 ;
        RECT 33.880 58.250 34.020 70.770 ;
        RECT 35.260 70.150 35.400 71.870 ;
        RECT 36.180 70.910 36.320 71.870 ;
        RECT 36.640 71.510 36.780 74.590 ;
        RECT 36.580 71.190 36.840 71.510 ;
        RECT 36.180 70.770 36.780 70.910 ;
        RECT 35.200 69.830 35.460 70.150 ;
        RECT 36.640 68.790 36.780 70.770 ;
        RECT 37.100 69.130 37.240 79.690 ;
        RECT 37.560 69.470 37.700 79.690 ;
        RECT 37.500 69.150 37.760 69.470 ;
        RECT 37.040 68.810 37.300 69.130 ;
        RECT 36.580 68.470 36.840 68.790 ;
        RECT 35.660 68.130 35.920 68.450 ;
        RECT 35.720 66.750 35.860 68.130 ;
        RECT 37.560 67.430 37.700 69.150 ;
        RECT 37.500 67.110 37.760 67.430 ;
        RECT 35.660 66.430 35.920 66.750 ;
        RECT 34.740 66.090 35.000 66.410 ;
        RECT 34.280 63.260 34.540 63.350 ;
        RECT 34.800 63.260 34.940 66.090 ;
        RECT 35.200 64.390 35.460 64.710 ;
        RECT 35.260 63.690 35.400 64.390 ;
        RECT 35.200 63.370 35.460 63.690 ;
        RECT 34.280 63.120 34.940 63.260 ;
        RECT 34.280 63.030 34.540 63.120 ;
        RECT 34.800 61.310 34.940 63.120 ;
        RECT 35.260 61.650 35.400 63.370 ;
        RECT 35.720 63.350 35.860 66.430 ;
        RECT 37.560 64.710 37.700 67.110 ;
        RECT 37.500 64.390 37.760 64.710 ;
        RECT 35.660 63.030 35.920 63.350 ;
        RECT 35.200 61.330 35.460 61.650 ;
        RECT 34.740 60.990 35.000 61.310 ;
        RECT 33.820 57.930 34.080 58.250 ;
        RECT 33.880 56.630 34.020 57.930 ;
        RECT 33.880 56.490 34.480 56.630 ;
        RECT 33.820 55.210 34.080 55.530 ;
        RECT 33.360 50.790 33.620 51.110 ;
        RECT 33.880 50.430 34.020 55.210 ;
        RECT 34.340 52.810 34.480 56.490 ;
        RECT 34.280 52.490 34.540 52.810 ;
        RECT 34.280 50.450 34.540 50.770 ;
        RECT 33.820 50.110 34.080 50.430 ;
        RECT 34.340 49.750 34.480 50.450 ;
        RECT 34.280 49.430 34.540 49.750 ;
        RECT 33.360 49.090 33.620 49.410 ;
        RECT 30.600 46.710 30.860 47.030 ;
        RECT 32.890 46.855 33.170 47.225 ;
        RECT 27.840 45.350 28.100 45.670 ;
        RECT 30.140 45.350 30.400 45.670 ;
        RECT 26.460 44.670 26.720 44.990 ;
        RECT 26.910 44.815 27.190 45.185 ;
        RECT 30.660 45.070 30.800 46.710 ;
        RECT 33.420 46.690 33.560 49.090 ;
        RECT 33.820 47.730 34.080 48.050 ;
        RECT 32.900 46.370 33.160 46.690 ;
        RECT 33.360 46.370 33.620 46.690 ;
        RECT 30.950 45.835 32.490 46.205 ;
        RECT 30.200 44.990 30.800 45.070 ;
        RECT 30.140 44.930 30.800 44.990 ;
        RECT 26.920 44.670 27.180 44.815 ;
        RECT 30.140 44.670 30.400 44.930 ;
        RECT 32.430 44.815 32.710 45.185 ;
        RECT 32.960 45.070 33.100 46.370 ;
        RECT 32.960 44.990 33.560 45.070 ;
        RECT 32.960 44.930 33.620 44.990 ;
        RECT 26.000 41.610 26.260 41.930 ;
        RECT 26.060 40.230 26.200 41.610 ;
        RECT 26.520 41.250 26.660 44.670 ;
        RECT 29.680 43.990 29.940 44.310 ;
        RECT 27.650 43.115 29.190 43.485 ;
        RECT 29.740 41.930 29.880 43.990 ;
        RECT 32.500 42.950 32.640 44.815 ;
        RECT 33.360 44.670 33.620 44.930 ;
        RECT 30.600 42.630 30.860 42.950 ;
        RECT 32.440 42.630 32.700 42.950 ;
        RECT 29.680 41.610 29.940 41.930 ;
        RECT 26.460 40.930 26.720 41.250 ;
        RECT 26.000 39.910 26.260 40.230 ;
        RECT 23.700 38.210 23.960 38.530 ;
        RECT 26.060 37.510 26.200 39.910 ;
        RECT 26.920 39.230 27.180 39.550 ;
        RECT 26.000 37.190 26.260 37.510 ;
        RECT 26.980 37.170 27.120 39.230 ;
        RECT 30.660 38.530 30.800 42.630 ;
        RECT 33.880 41.930 34.020 47.730 ;
        RECT 33.350 41.415 33.630 41.785 ;
        RECT 33.820 41.610 34.080 41.930 ;
        RECT 33.360 41.270 33.620 41.415 ;
        RECT 30.950 40.395 32.490 40.765 ;
        RECT 34.340 40.230 34.480 49.430 ;
        RECT 34.800 48.050 34.940 60.990 ;
        RECT 35.260 59.270 35.400 61.330 ;
        RECT 36.120 59.970 36.380 60.290 ;
        RECT 35.200 58.950 35.460 59.270 ;
        RECT 36.180 56.210 36.320 59.970 ;
        RECT 36.120 55.890 36.380 56.210 ;
        RECT 38.020 55.870 38.160 80.370 ;
        RECT 38.420 79.865 38.680 80.010 ;
        RECT 38.410 79.495 38.690 79.865 ;
        RECT 38.940 70.345 39.080 88.530 ;
        RECT 43.480 88.190 43.740 88.510 ;
        RECT 42.560 87.170 42.820 87.490 ;
        RECT 41.180 86.150 41.440 86.470 ;
        RECT 39.340 84.450 39.600 84.770 ;
        RECT 39.400 77.030 39.540 84.450 ;
        RECT 41.240 83.750 41.380 86.150 ;
        RECT 42.620 85.450 42.760 87.170 ;
        RECT 43.540 86.470 43.680 88.190 ;
        RECT 43.480 86.150 43.740 86.470 ;
        RECT 42.560 85.130 42.820 85.450 ;
        RECT 41.180 83.430 41.440 83.750 ;
        RECT 41.240 80.350 41.380 83.430 ;
        RECT 41.180 80.030 41.440 80.350 ;
        RECT 42.560 80.030 42.820 80.350 ;
        RECT 40.250 79.495 40.530 79.865 ;
        RECT 39.400 76.950 40.000 77.030 ;
        RECT 39.400 76.890 40.060 76.950 ;
        RECT 39.800 76.630 40.060 76.890 ;
        RECT 39.340 73.570 39.600 73.890 ;
        RECT 39.400 72.190 39.540 73.570 ;
        RECT 39.340 71.870 39.600 72.190 ;
        RECT 38.870 69.975 39.150 70.345 ;
        RECT 38.940 67.090 39.080 69.975 ;
        RECT 39.800 68.360 40.060 68.450 ;
        RECT 40.320 68.360 40.460 79.495 ;
        RECT 41.180 79.010 41.440 79.330 ;
        RECT 41.240 77.630 41.380 79.010 ;
        RECT 42.100 77.990 42.360 78.310 ;
        RECT 40.720 77.310 40.980 77.630 ;
        RECT 41.180 77.310 41.440 77.630 ;
        RECT 41.640 77.310 41.900 77.630 ;
        RECT 40.780 74.230 40.920 77.310 ;
        RECT 41.700 74.570 41.840 77.310 ;
        RECT 41.640 74.250 41.900 74.570 ;
        RECT 40.720 73.910 40.980 74.230 ;
        RECT 40.780 72.530 40.920 73.910 ;
        RECT 40.720 72.210 40.980 72.530 ;
        RECT 40.780 70.150 40.920 72.210 ;
        RECT 41.180 71.530 41.440 71.850 ;
        RECT 40.720 69.830 40.980 70.150 ;
        RECT 39.800 68.220 40.460 68.360 ;
        RECT 39.800 68.130 40.060 68.220 ;
        RECT 38.880 66.770 39.140 67.090 ;
        RECT 38.420 57.590 38.680 57.910 ;
        RECT 38.480 56.550 38.620 57.590 ;
        RECT 38.940 57.570 39.080 66.770 ;
        RECT 39.340 63.710 39.600 64.030 ;
        RECT 38.880 57.250 39.140 57.570 ;
        RECT 38.420 56.230 38.680 56.550 ;
        RECT 37.960 55.550 38.220 55.870 ;
        RECT 38.020 53.490 38.160 55.550 ;
        RECT 38.940 55.530 39.080 57.250 ;
        RECT 38.880 55.210 39.140 55.530 ;
        RECT 39.400 54.850 39.540 63.710 ;
        RECT 39.800 57.930 40.060 58.250 ;
        RECT 39.340 54.530 39.600 54.850 ;
        RECT 37.960 53.170 38.220 53.490 ;
        RECT 39.860 52.470 40.000 57.930 ;
        RECT 40.320 55.190 40.460 68.220 ;
        RECT 41.240 65.730 41.380 71.530 ;
        RECT 41.700 71.170 41.840 74.250 ;
        RECT 41.640 70.850 41.900 71.170 ;
        RECT 42.160 66.750 42.300 77.990 ;
        RECT 42.620 75.590 42.760 80.030 ;
        RECT 43.020 79.350 43.280 79.670 ;
        RECT 42.560 75.270 42.820 75.590 ;
        RECT 43.080 75.250 43.220 79.350 ;
        RECT 43.020 74.930 43.280 75.250 ;
        RECT 44.000 74.570 44.140 141.570 ;
        RECT 44.460 128.970 44.600 149.730 ;
        RECT 44.920 139.170 45.060 150.750 ;
        RECT 45.840 149.030 45.980 156.870 ;
        RECT 46.300 154.130 46.440 158.910 ;
        RECT 47.150 156.335 47.430 156.705 ;
        RECT 47.160 156.190 47.420 156.335 ;
        RECT 48.600 154.470 48.740 161.290 ;
        RECT 49.060 159.910 49.200 161.290 ;
        RECT 49.000 159.590 49.260 159.910 ;
        RECT 50.900 158.210 51.040 161.290 ;
        RECT 50.840 157.890 51.100 158.210 ;
        RECT 50.900 156.170 51.040 157.890 ;
        RECT 50.840 155.850 51.100 156.170 ;
        RECT 49.920 155.170 50.180 155.490 ;
        RECT 49.980 154.470 50.120 155.170 ;
        RECT 48.540 154.150 48.800 154.470 ;
        RECT 49.920 154.150 50.180 154.470 ;
        RECT 46.240 153.810 46.500 154.130 ;
        RECT 45.780 148.710 46.040 149.030 ;
        RECT 45.780 148.030 46.040 148.350 ;
        RECT 45.840 145.970 45.980 148.030 ;
        RECT 45.780 145.650 46.040 145.970 ;
        RECT 45.840 139.170 45.980 145.650 ;
        RECT 46.300 143.250 46.440 153.810 ;
        RECT 50.900 151.150 51.040 155.850 ;
        RECT 51.760 155.170 52.020 155.490 ;
        RECT 51.820 154.130 51.960 155.170 ;
        RECT 51.760 153.810 52.020 154.130 ;
        RECT 51.300 153.470 51.560 153.790 ;
        RECT 51.360 151.750 51.500 153.470 ;
        RECT 51.760 152.450 52.020 152.770 ;
        RECT 51.820 151.750 51.960 152.450 ;
        RECT 51.300 151.430 51.560 151.750 ;
        RECT 51.760 151.430 52.020 151.750 ;
        RECT 50.900 151.010 51.500 151.150 ;
        RECT 47.620 150.070 47.880 150.390 ;
        RECT 47.680 148.350 47.820 150.070 ;
        RECT 50.840 149.730 51.100 150.050 ;
        RECT 47.620 148.030 47.880 148.350 ;
        RECT 50.380 148.030 50.640 148.350 ;
        RECT 47.680 143.590 47.820 148.030 ;
        RECT 50.440 145.290 50.580 148.030 ;
        RECT 50.380 144.970 50.640 145.290 ;
        RECT 49.000 144.290 49.260 144.610 ;
        RECT 47.620 143.270 47.880 143.590 ;
        RECT 46.240 142.930 46.500 143.250 ;
        RECT 47.160 142.590 47.420 142.910 ;
        RECT 47.220 140.870 47.360 142.590 ;
        RECT 47.160 140.550 47.420 140.870 ;
        RECT 49.060 140.190 49.200 144.290 ;
        RECT 50.440 143.590 50.580 144.970 ;
        RECT 50.380 143.270 50.640 143.590 ;
        RECT 49.000 139.870 49.260 140.190 ;
        RECT 46.240 139.530 46.500 139.850 ;
        RECT 44.860 138.850 45.120 139.170 ;
        RECT 45.780 138.850 46.040 139.170 ;
        RECT 44.920 136.190 45.060 138.850 ;
        RECT 45.840 137.470 45.980 138.850 ;
        RECT 46.300 137.470 46.440 139.530 ;
        RECT 47.620 137.490 47.880 137.810 ;
        RECT 45.780 137.150 46.040 137.470 ;
        RECT 46.240 137.150 46.500 137.470 ;
        RECT 44.920 136.050 45.520 136.190 ;
        RECT 44.850 135.255 45.130 135.625 ;
        RECT 44.860 135.110 45.120 135.255 ;
        RECT 44.920 132.710 45.060 135.110 ;
        RECT 45.380 134.750 45.520 136.050 ;
        RECT 45.840 135.430 45.980 137.150 ;
        RECT 45.780 135.110 46.040 135.430 ;
        RECT 46.300 134.830 46.440 137.150 ;
        RECT 47.150 135.255 47.430 135.625 ;
        RECT 47.160 135.110 47.420 135.255 ;
        RECT 45.320 134.430 45.580 134.750 ;
        RECT 45.840 134.690 46.440 134.830 ;
        RECT 44.860 132.390 45.120 132.710 ;
        RECT 45.380 131.010 45.520 134.430 ;
        RECT 45.840 134.410 45.980 134.690 ;
        RECT 45.780 134.090 46.040 134.410 ;
        RECT 46.700 134.090 46.960 134.410 ;
        RECT 45.840 132.370 45.980 134.090 ;
        RECT 46.240 133.410 46.500 133.730 ;
        RECT 45.780 132.050 46.040 132.370 ;
        RECT 45.320 130.690 45.580 131.010 ;
        RECT 44.400 128.650 44.660 128.970 ;
        RECT 46.300 118.410 46.440 133.410 ;
        RECT 46.760 124.550 46.900 134.090 ;
        RECT 47.220 132.710 47.360 135.110 ;
        RECT 47.680 134.070 47.820 137.490 ;
        RECT 48.080 134.770 48.340 135.090 ;
        RECT 47.620 133.750 47.880 134.070 ;
        RECT 47.160 132.390 47.420 132.710 ;
        RECT 46.700 124.230 46.960 124.550 ;
        RECT 44.920 118.270 46.440 118.410 ;
        RECT 44.400 117.430 44.660 117.750 ;
        RECT 44.460 116.390 44.600 117.430 ;
        RECT 44.400 116.070 44.660 116.390 ;
        RECT 44.400 104.510 44.660 104.830 ;
        RECT 44.460 97.350 44.600 104.510 ;
        RECT 44.400 97.030 44.660 97.350 ;
        RECT 43.020 74.250 43.280 74.570 ;
        RECT 43.940 74.250 44.200 74.570 ;
        RECT 43.080 72.870 43.220 74.250 ;
        RECT 43.480 73.570 43.740 73.890 ;
        RECT 43.020 72.550 43.280 72.870 ;
        RECT 43.020 68.470 43.280 68.790 ;
        RECT 42.100 66.430 42.360 66.750 ;
        RECT 43.080 66.070 43.220 68.470 ;
        RECT 42.560 65.750 42.820 66.070 ;
        RECT 43.020 65.750 43.280 66.070 ;
        RECT 41.180 65.410 41.440 65.730 ;
        RECT 42.620 61.990 42.760 65.750 ;
        RECT 42.560 61.670 42.820 61.990 ;
        RECT 42.620 59.270 42.760 61.670 ;
        RECT 43.540 61.310 43.680 73.570 ;
        RECT 44.920 70.110 45.060 118.270 ;
        RECT 45.780 117.430 46.040 117.750 ;
        RECT 45.840 115.710 45.980 117.430 ;
        RECT 47.680 116.050 47.820 133.750 ;
        RECT 48.140 131.690 48.280 134.770 ;
        RECT 50.900 134.750 51.040 149.730 ;
        RECT 51.360 145.970 51.500 151.010 ;
        RECT 51.820 150.730 51.960 151.430 ;
        RECT 51.760 150.410 52.020 150.730 ;
        RECT 52.280 149.030 52.420 161.290 ;
        RECT 52.740 156.170 52.880 161.290 ;
        RECT 53.660 160.930 53.800 163.330 ;
        RECT 55.040 162.290 55.180 164.350 ;
        RECT 56.420 162.630 56.560 164.350 ;
        RECT 55.900 162.310 56.160 162.630 ;
        RECT 56.360 162.310 56.620 162.630 ;
        RECT 54.980 161.970 55.240 162.290 ;
        RECT 54.060 161.290 54.320 161.610 ;
        RECT 53.600 160.610 53.860 160.930 ;
        RECT 53.660 156.170 53.800 160.610 ;
        RECT 54.120 157.190 54.260 161.290 ;
        RECT 54.520 159.590 54.780 159.910 ;
        RECT 54.060 156.870 54.320 157.190 ;
        RECT 54.580 156.850 54.720 159.590 ;
        RECT 54.520 156.530 54.780 156.850 ;
        RECT 54.580 156.170 54.720 156.530 ;
        RECT 52.680 155.850 52.940 156.170 ;
        RECT 53.600 155.850 53.860 156.170 ;
        RECT 54.520 155.850 54.780 156.170 ;
        RECT 52.740 151.410 52.880 155.850 ;
        RECT 52.680 151.090 52.940 151.410 ;
        RECT 53.660 150.390 53.800 155.850 ;
        RECT 54.580 154.550 54.720 155.850 ;
        RECT 54.120 154.410 54.720 154.550 ;
        RECT 54.120 152.770 54.260 154.410 ;
        RECT 55.040 153.870 55.180 161.970 ;
        RECT 55.440 160.610 55.700 160.930 ;
        RECT 55.500 156.170 55.640 160.610 ;
        RECT 55.960 159.910 56.100 162.310 ;
        RECT 56.360 161.630 56.620 161.950 ;
        RECT 57.740 161.630 58.000 161.950 ;
        RECT 55.900 159.590 56.160 159.910 ;
        RECT 55.900 157.890 56.160 158.210 ;
        RECT 55.960 156.170 56.100 157.890 ;
        RECT 56.420 157.190 56.560 161.630 ;
        RECT 57.280 161.290 57.540 161.610 ;
        RECT 57.340 159.570 57.480 161.290 ;
        RECT 57.280 159.250 57.540 159.570 ;
        RECT 56.820 158.910 57.080 159.230 ;
        RECT 56.360 156.870 56.620 157.190 ;
        RECT 56.360 156.190 56.620 156.510 ;
        RECT 55.440 155.850 55.700 156.170 ;
        RECT 55.900 155.850 56.160 156.170 ;
        RECT 54.580 153.790 55.180 153.870 ;
        RECT 54.520 153.730 55.180 153.790 ;
        RECT 54.520 153.470 54.780 153.730 ;
        RECT 54.060 152.450 54.320 152.770 ;
        RECT 55.040 150.390 55.180 153.730 ;
        RECT 53.600 150.070 53.860 150.390 ;
        RECT 54.980 150.070 55.240 150.390 ;
        RECT 52.220 148.710 52.480 149.030 ;
        RECT 52.680 147.690 52.940 148.010 ;
        RECT 51.300 145.650 51.560 145.970 ;
        RECT 52.740 138.150 52.880 147.690 ;
        RECT 55.040 145.290 55.180 150.070 ;
        RECT 56.420 148.010 56.560 156.190 ;
        RECT 56.880 151.750 57.020 158.910 ;
        RECT 57.340 156.510 57.480 159.250 ;
        RECT 57.280 156.190 57.540 156.510 ;
        RECT 57.280 153.470 57.540 153.790 ;
        RECT 57.340 151.750 57.480 153.470 ;
        RECT 56.820 151.430 57.080 151.750 ;
        RECT 57.280 151.430 57.540 151.750 ;
        RECT 57.800 151.070 57.940 161.630 ;
        RECT 59.180 161.465 59.320 166.570 ;
        RECT 58.660 160.950 58.920 161.270 ;
        RECT 59.110 161.095 59.390 161.465 ;
        RECT 58.200 157.890 58.460 158.210 ;
        RECT 58.260 157.190 58.400 157.890 ;
        RECT 58.720 157.190 58.860 160.950 ;
        RECT 59.640 159.230 59.780 172.170 ;
        RECT 60.500 171.490 60.760 171.810 ;
        RECT 60.560 170.450 60.700 171.490 ;
        RECT 60.500 170.130 60.760 170.450 ;
        RECT 60.500 169.450 60.760 169.770 ;
        RECT 60.560 167.730 60.700 169.450 ;
        RECT 60.500 167.410 60.760 167.730 ;
        RECT 61.020 166.710 61.160 172.170 ;
        RECT 63.320 170.790 63.460 172.170 ;
        RECT 63.260 170.470 63.520 170.790 ;
        RECT 61.880 169.110 62.140 169.430 ;
        RECT 61.420 167.410 61.680 167.730 ;
        RECT 60.040 166.390 60.300 166.710 ;
        RECT 60.560 166.570 61.160 166.710 ;
        RECT 60.100 161.950 60.240 166.390 ;
        RECT 60.040 161.630 60.300 161.950 ;
        RECT 60.560 160.105 60.700 166.570 ;
        RECT 60.490 159.735 60.770 160.105 ;
        RECT 60.960 159.590 61.220 159.910 ;
        RECT 60.500 159.250 60.760 159.570 ;
        RECT 59.580 158.910 59.840 159.230 ;
        RECT 60.040 158.230 60.300 158.550 ;
        RECT 58.200 156.870 58.460 157.190 ;
        RECT 58.660 156.870 58.920 157.190 ;
        RECT 60.100 156.170 60.240 158.230 ;
        RECT 60.040 155.850 60.300 156.170 ;
        RECT 58.200 155.170 58.460 155.490 ;
        RECT 59.120 155.170 59.380 155.490 ;
        RECT 57.740 150.750 58.000 151.070 ;
        RECT 56.360 147.690 56.620 148.010 ;
        RECT 57.800 147.330 57.940 150.750 ;
        RECT 57.740 147.010 58.000 147.330 ;
        RECT 54.980 144.970 55.240 145.290 ;
        RECT 55.040 143.250 55.180 144.970 ;
        RECT 57.800 143.590 57.940 147.010 ;
        RECT 57.740 143.270 58.000 143.590 ;
        RECT 54.980 142.930 55.240 143.250 ;
        RECT 54.520 141.570 54.780 141.890 ;
        RECT 53.140 140.550 53.400 140.870 ;
        RECT 52.680 137.830 52.940 138.150 ;
        RECT 51.760 137.150 52.020 137.470 ;
        RECT 51.820 135.430 51.960 137.150 ;
        RECT 51.760 135.110 52.020 135.430 ;
        RECT 50.840 134.430 51.100 134.750 ;
        RECT 49.920 132.050 50.180 132.370 ;
        RECT 48.080 131.370 48.340 131.690 ;
        RECT 49.000 130.690 49.260 131.010 ;
        RECT 49.060 128.970 49.200 130.690 ;
        RECT 49.000 128.650 49.260 128.970 ;
        RECT 49.980 124.550 50.120 132.050 ;
        RECT 50.900 129.990 51.040 134.430 ;
        RECT 52.740 134.410 52.880 137.830 ;
        RECT 53.200 134.750 53.340 140.550 ;
        RECT 54.580 139.850 54.720 141.570 ;
        RECT 55.040 139.850 55.180 142.930 ;
        RECT 57.800 142.570 57.940 143.270 ;
        RECT 58.260 142.570 58.400 155.170 ;
        RECT 59.180 150.730 59.320 155.170 ;
        RECT 60.100 154.130 60.240 155.850 ;
        RECT 60.040 153.810 60.300 154.130 ;
        RECT 60.560 153.110 60.700 159.250 ;
        RECT 61.020 154.470 61.160 159.590 ;
        RECT 61.480 158.550 61.620 167.410 ;
        RECT 61.940 161.270 62.080 169.110 ;
        RECT 63.260 168.770 63.520 169.090 ;
        RECT 63.320 167.390 63.460 168.770 ;
        RECT 64.240 168.070 64.380 172.170 ;
        RECT 69.240 171.830 69.500 172.150 ;
        RECT 70.610 171.975 70.890 172.345 ;
        RECT 71.600 172.150 71.740 173.190 ;
        RECT 74.360 173.170 74.500 181.510 ;
        RECT 80.800 173.510 80.940 181.510 ;
        RECT 80.740 173.190 81.000 173.510 ;
        RECT 83.040 173.190 83.300 173.510 ;
        RECT 74.300 172.850 74.560 173.170 ;
        RECT 76.200 172.770 78.180 172.910 ;
        RECT 76.200 172.490 76.340 172.770 ;
        RECT 76.140 172.170 76.400 172.490 ;
        RECT 78.040 172.150 78.180 172.770 ;
        RECT 83.100 172.490 83.240 173.190 ;
        RECT 84.020 172.830 84.160 181.510 ;
        RECT 89.020 173.190 89.280 173.510 ;
        RECT 83.960 172.510 84.220 172.830 ;
        RECT 81.200 172.170 81.460 172.490 ;
        RECT 83.040 172.345 83.300 172.490 ;
        RECT 70.620 171.830 70.880 171.975 ;
        RECT 71.540 171.830 71.800 172.150 ;
        RECT 73.380 171.830 73.640 172.150 ;
        RECT 73.840 171.830 74.100 172.150 ;
        RECT 77.520 171.830 77.780 172.150 ;
        RECT 77.980 171.830 78.240 172.150 ;
        RECT 78.440 171.830 78.700 172.150 ;
        RECT 79.820 171.830 80.080 172.150 ;
        RECT 67.860 171.490 68.120 171.810 ;
        RECT 69.300 171.665 69.440 171.830 ;
        RECT 66.940 169.450 67.200 169.770 ;
        RECT 66.470 168.575 66.750 168.945 ;
        RECT 64.180 167.750 64.440 168.070 ;
        RECT 63.260 167.070 63.520 167.390 ;
        RECT 64.240 166.790 64.380 167.750 ;
        RECT 65.090 167.215 65.370 167.585 ;
        RECT 63.780 166.650 64.380 166.790 ;
        RECT 62.800 165.030 63.060 165.350 ;
        RECT 61.880 160.950 62.140 161.270 ;
        RECT 61.420 158.230 61.680 158.550 ;
        RECT 61.880 158.230 62.140 158.550 ;
        RECT 60.960 154.150 61.220 154.470 ;
        RECT 60.500 152.790 60.760 153.110 ;
        RECT 61.940 151.830 62.080 158.230 ;
        RECT 62.860 156.850 63.000 165.030 ;
        RECT 63.260 158.570 63.520 158.890 ;
        RECT 62.800 156.530 63.060 156.850 ;
        RECT 62.340 156.190 62.600 156.510 ;
        RECT 62.400 152.770 62.540 156.190 ;
        RECT 62.340 152.450 62.600 152.770 ;
        RECT 61.940 151.690 62.540 151.830 ;
        RECT 59.120 150.410 59.380 150.730 ;
        RECT 59.120 149.730 59.380 150.050 ;
        RECT 59.180 149.030 59.320 149.730 ;
        RECT 59.120 148.710 59.380 149.030 ;
        RECT 62.400 148.010 62.540 151.690 ;
        RECT 62.790 150.895 63.070 151.265 ;
        RECT 60.960 147.690 61.220 148.010 ;
        RECT 62.340 147.690 62.600 148.010 ;
        RECT 59.580 144.630 59.840 144.950 ;
        RECT 57.740 142.250 58.000 142.570 ;
        RECT 58.200 142.250 58.460 142.570 ;
        RECT 57.800 140.870 57.940 142.250 ;
        RECT 58.260 140.870 58.400 142.250 ;
        RECT 57.740 140.550 58.000 140.870 ;
        RECT 58.200 140.550 58.460 140.870 ;
        RECT 54.520 139.530 54.780 139.850 ;
        RECT 54.980 139.530 55.240 139.850 ;
        RECT 53.140 134.430 53.400 134.750 ;
        RECT 52.680 134.090 52.940 134.410 ;
        RECT 53.200 132.710 53.340 134.430 ;
        RECT 53.140 132.390 53.400 132.710 ;
        RECT 53.200 131.690 53.340 132.390 ;
        RECT 55.040 132.030 55.180 139.530 ;
        RECT 55.440 139.190 55.700 139.510 ;
        RECT 55.500 138.150 55.640 139.190 ;
        RECT 55.440 137.830 55.700 138.150 ;
        RECT 58.660 137.150 58.920 137.470 ;
        RECT 57.740 136.810 58.000 137.130 ;
        RECT 57.280 133.750 57.540 134.070 ;
        RECT 54.980 131.710 55.240 132.030 ;
        RECT 53.140 131.370 53.400 131.690 ;
        RECT 57.340 129.990 57.480 133.750 ;
        RECT 57.800 129.990 57.940 136.810 ;
        RECT 50.840 129.670 51.100 129.990 ;
        RECT 57.280 129.670 57.540 129.990 ;
        RECT 57.740 129.670 58.000 129.990 ;
        RECT 52.680 128.650 52.940 128.970 ;
        RECT 55.900 128.650 56.160 128.970 ;
        RECT 52.740 126.930 52.880 128.650 ;
        RECT 54.980 127.970 55.240 128.290 ;
        RECT 52.680 126.610 52.940 126.930 ;
        RECT 52.740 126.250 52.880 126.610 ;
        RECT 52.680 125.930 52.940 126.250 ;
        RECT 49.920 124.230 50.180 124.550 ;
        RECT 48.080 123.550 48.340 123.870 ;
        RECT 48.140 121.490 48.280 123.550 ;
        RECT 49.460 123.210 49.720 123.530 ;
        RECT 48.540 122.870 48.800 123.190 ;
        RECT 48.080 121.170 48.340 121.490 ;
        RECT 48.140 120.810 48.280 121.170 ;
        RECT 48.080 120.490 48.340 120.810 ;
        RECT 47.620 115.730 47.880 116.050 ;
        RECT 45.780 115.390 46.040 115.710 ;
        RECT 48.140 112.650 48.280 120.490 ;
        RECT 48.600 119.110 48.740 122.870 ;
        RECT 49.000 120.830 49.260 121.150 ;
        RECT 49.060 119.110 49.200 120.830 ;
        RECT 48.540 118.790 48.800 119.110 ;
        RECT 49.000 118.790 49.260 119.110 ;
        RECT 49.520 118.410 49.660 123.210 ;
        RECT 49.060 118.270 49.660 118.410 ;
        RECT 49.060 113.670 49.200 118.270 ;
        RECT 52.220 117.090 52.480 117.410 ;
        RECT 51.300 115.050 51.560 115.370 ;
        RECT 49.920 114.370 50.180 114.690 ;
        RECT 49.000 113.350 49.260 113.670 ;
        RECT 48.080 112.330 48.340 112.650 ;
        RECT 48.140 109.930 48.280 112.330 ;
        RECT 49.060 110.270 49.200 113.350 ;
        RECT 49.000 109.950 49.260 110.270 ;
        RECT 48.080 109.610 48.340 109.930 ;
        RECT 48.540 109.610 48.800 109.930 ;
        RECT 46.240 108.930 46.500 109.250 ;
        RECT 46.300 107.210 46.440 108.930 ;
        RECT 47.620 107.910 47.880 108.230 ;
        RECT 45.780 106.890 46.040 107.210 ;
        RECT 46.240 106.890 46.500 107.210 ;
        RECT 45.840 101.510 45.980 106.890 ;
        RECT 47.160 106.550 47.420 106.870 ;
        RECT 47.220 103.810 47.360 106.550 ;
        RECT 47.160 103.490 47.420 103.810 ;
        RECT 45.380 101.370 45.980 101.510 ;
        RECT 45.380 99.390 45.520 101.370 ;
        RECT 45.780 100.770 46.040 101.090 ;
        RECT 47.220 100.830 47.360 103.490 ;
        RECT 47.680 101.430 47.820 107.910 ;
        RECT 48.140 104.490 48.280 109.610 ;
        RECT 48.600 107.550 48.740 109.610 ;
        RECT 48.540 107.230 48.800 107.550 ;
        RECT 49.980 107.210 50.120 114.370 ;
        RECT 51.360 112.650 51.500 115.050 ;
        RECT 51.300 112.330 51.560 112.650 ;
        RECT 50.840 111.990 51.100 112.310 ;
        RECT 50.900 110.950 51.040 111.990 ;
        RECT 50.840 110.630 51.100 110.950 ;
        RECT 50.380 107.570 50.640 107.890 ;
        RECT 49.920 106.890 50.180 107.210 ;
        RECT 48.540 106.210 48.800 106.530 ;
        RECT 48.600 105.510 48.740 106.210 ;
        RECT 49.980 105.590 50.120 106.890 ;
        RECT 48.540 105.190 48.800 105.510 ;
        RECT 49.520 105.450 50.120 105.590 ;
        RECT 48.080 104.170 48.340 104.490 ;
        RECT 48.140 101.770 48.280 104.170 ;
        RECT 48.080 101.450 48.340 101.770 ;
        RECT 47.620 101.110 47.880 101.430 ;
        RECT 48.080 100.830 48.340 101.090 ;
        RECT 47.220 100.770 48.340 100.830 ;
        RECT 45.320 99.070 45.580 99.390 ;
        RECT 45.840 96.330 45.980 100.770 ;
        RECT 47.220 100.690 48.280 100.770 ;
        RECT 46.240 99.750 46.500 100.070 ;
        RECT 46.300 96.330 46.440 99.750 ;
        RECT 45.780 96.010 46.040 96.330 ;
        RECT 46.240 96.010 46.500 96.330 ;
        RECT 47.160 90.570 47.420 90.890 ;
        RECT 47.220 85.790 47.360 90.570 ;
        RECT 47.680 86.470 47.820 100.690 ;
        RECT 48.600 99.730 48.740 105.190 ;
        RECT 49.520 102.450 49.660 105.450 ;
        RECT 49.920 104.850 50.180 105.170 ;
        RECT 49.460 102.130 49.720 102.450 ;
        RECT 49.000 101.450 49.260 101.770 ;
        RECT 49.060 100.070 49.200 101.450 ;
        RECT 49.980 101.090 50.120 104.850 ;
        RECT 50.440 103.810 50.580 107.570 ;
        RECT 51.300 106.890 51.560 107.210 ;
        RECT 50.840 106.550 51.100 106.870 ;
        RECT 50.380 103.490 50.640 103.810 ;
        RECT 49.920 100.770 50.180 101.090 ;
        RECT 49.000 99.750 49.260 100.070 ;
        RECT 48.540 99.410 48.800 99.730 ;
        RECT 48.600 96.750 48.740 99.410 ;
        RECT 50.440 98.710 50.580 103.490 ;
        RECT 50.900 102.790 51.040 106.550 ;
        RECT 50.840 102.470 51.100 102.790 ;
        RECT 50.380 98.390 50.640 98.710 ;
        RECT 48.140 96.610 50.120 96.750 ;
        RECT 50.380 96.690 50.640 97.010 ;
        RECT 48.140 96.330 48.280 96.610 ;
        RECT 49.980 96.330 50.120 96.610 ;
        RECT 48.080 96.010 48.340 96.330 ;
        RECT 48.540 96.010 48.800 96.330 ;
        RECT 49.920 96.010 50.180 96.330 ;
        RECT 48.600 94.630 48.740 96.010 ;
        RECT 48.540 94.310 48.800 94.630 ;
        RECT 49.980 93.610 50.120 96.010 ;
        RECT 50.440 94.290 50.580 96.690 ;
        RECT 50.900 95.990 51.040 102.470 ;
        RECT 50.840 95.670 51.100 95.990 ;
        RECT 51.360 94.630 51.500 106.890 ;
        RECT 51.760 102.470 52.020 102.790 ;
        RECT 51.300 94.310 51.560 94.630 ;
        RECT 50.380 93.970 50.640 94.290 ;
        RECT 49.920 93.290 50.180 93.610 ;
        RECT 50.440 88.510 50.580 93.970 ;
        RECT 51.820 93.350 51.960 102.470 ;
        RECT 52.280 101.430 52.420 117.090 ;
        RECT 52.740 115.710 52.880 125.930 ;
        RECT 54.060 123.550 54.320 123.870 ;
        RECT 54.120 123.385 54.260 123.550 ;
        RECT 54.050 123.015 54.330 123.385 ;
        RECT 54.060 122.530 54.320 122.850 ;
        RECT 54.120 120.470 54.260 122.530 ;
        RECT 54.060 120.150 54.320 120.470 ;
        RECT 55.040 119.305 55.180 127.970 ;
        RECT 55.960 125.570 56.100 128.650 ;
        RECT 55.900 125.250 56.160 125.570 ;
        RECT 57.800 124.550 57.940 129.670 ;
        RECT 57.740 124.230 58.000 124.550 ;
        RECT 58.190 124.375 58.470 124.745 ;
        RECT 57.280 123.550 57.540 123.870 ;
        RECT 55.440 123.210 55.700 123.530 ;
        RECT 55.500 121.830 55.640 123.210 ;
        RECT 55.440 121.510 55.700 121.830 ;
        RECT 55.900 119.810 56.160 120.130 ;
        RECT 56.820 119.810 57.080 120.130 ;
        RECT 54.970 118.935 55.250 119.305 ;
        RECT 53.600 118.110 53.860 118.430 ;
        RECT 53.140 117.770 53.400 118.090 ;
        RECT 52.680 115.390 52.940 115.710 ;
        RECT 53.200 112.990 53.340 117.770 ;
        RECT 53.140 112.670 53.400 112.990 ;
        RECT 53.200 107.890 53.340 112.670 ;
        RECT 53.660 111.825 53.800 118.110 ;
        RECT 54.060 117.430 54.320 117.750 ;
        RECT 54.120 114.690 54.260 117.430 ;
        RECT 55.960 117.410 56.100 119.810 ;
        RECT 56.360 117.770 56.620 118.090 ;
        RECT 55.900 117.090 56.160 117.410 ;
        RECT 55.440 115.390 55.700 115.710 ;
        RECT 54.060 114.370 54.320 114.690 ;
        RECT 55.500 113.670 55.640 115.390 ;
        RECT 55.440 113.350 55.700 113.670 ;
        RECT 56.420 112.650 56.560 117.770 ;
        RECT 56.360 112.330 56.620 112.650 ;
        RECT 53.590 111.455 53.870 111.825 ;
        RECT 56.420 110.610 56.560 112.330 ;
        RECT 56.360 110.290 56.620 110.610 ;
        RECT 53.140 107.570 53.400 107.890 ;
        RECT 52.680 106.550 52.940 106.870 ;
        RECT 52.220 101.110 52.480 101.430 ;
        RECT 52.220 99.750 52.480 100.070 ;
        RECT 52.280 93.950 52.420 99.750 ;
        RECT 52.220 93.630 52.480 93.950 ;
        RECT 51.820 93.210 52.420 93.350 ;
        RECT 51.300 91.590 51.560 91.910 ;
        RECT 51.360 88.510 51.500 91.590 ;
        RECT 51.760 90.230 52.020 90.550 ;
        RECT 51.820 89.190 51.960 90.230 ;
        RECT 51.760 88.870 52.020 89.190 ;
        RECT 50.380 88.190 50.640 88.510 ;
        RECT 51.300 88.190 51.560 88.510 ;
        RECT 47.620 86.150 47.880 86.470 ;
        RECT 49.460 86.150 49.720 86.470 ;
        RECT 47.160 85.470 47.420 85.790 ;
        RECT 47.220 83.070 47.360 85.470 ;
        RECT 48.540 85.130 48.800 85.450 ;
        RECT 48.080 84.450 48.340 84.770 ;
        RECT 48.140 83.750 48.280 84.450 ;
        RECT 48.080 83.430 48.340 83.750 ;
        RECT 47.160 82.750 47.420 83.070 ;
        RECT 46.700 79.920 46.960 80.010 ;
        RECT 47.220 79.920 47.360 82.750 ;
        RECT 48.140 80.010 48.280 83.430 ;
        RECT 46.700 79.780 47.360 79.920 ;
        RECT 46.700 79.690 46.960 79.780 ;
        RECT 48.080 79.690 48.340 80.010 ;
        RECT 46.760 77.630 46.900 79.690 ;
        RECT 48.600 79.670 48.740 85.130 ;
        RECT 49.520 80.010 49.660 86.150 ;
        RECT 50.440 84.625 50.580 88.190 ;
        RECT 51.300 87.170 51.560 87.490 ;
        RECT 50.830 85.615 51.110 85.985 ;
        RECT 50.840 85.470 51.100 85.615 ;
        RECT 50.370 84.255 50.650 84.625 ;
        RECT 50.440 80.690 50.580 84.255 ;
        RECT 51.360 83.410 51.500 87.170 ;
        RECT 51.300 83.090 51.560 83.410 ;
        RECT 50.380 80.370 50.640 80.690 ;
        RECT 51.360 80.010 51.500 83.090 ;
        RECT 51.820 80.690 51.960 88.870 ;
        RECT 52.280 88.510 52.420 93.210 ;
        RECT 52.220 88.190 52.480 88.510 ;
        RECT 51.760 80.370 52.020 80.690 ;
        RECT 49.460 79.690 49.720 80.010 ;
        RECT 51.300 79.690 51.560 80.010 ;
        RECT 48.540 79.350 48.800 79.670 ;
        RECT 48.080 79.010 48.340 79.330 ;
        RECT 47.160 77.650 47.420 77.970 ;
        RECT 46.700 77.310 46.960 77.630 ;
        RECT 45.320 73.570 45.580 73.890 ;
        RECT 45.380 72.190 45.520 73.570 ;
        RECT 46.760 72.190 46.900 77.310 ;
        RECT 45.320 71.870 45.580 72.190 ;
        RECT 46.700 71.870 46.960 72.190 ;
        RECT 44.920 69.970 45.520 70.110 ;
        RECT 43.480 60.990 43.740 61.310 ;
        RECT 42.560 58.950 42.820 59.270 ;
        RECT 41.180 57.930 41.440 58.250 ;
        RECT 41.240 56.550 41.380 57.930 ;
        RECT 43.540 57.570 43.680 60.990 ;
        RECT 44.860 59.970 45.120 60.290 ;
        RECT 43.480 57.250 43.740 57.570 ;
        RECT 41.180 56.230 41.440 56.550 ;
        RECT 40.260 54.870 40.520 55.190 ;
        RECT 38.420 52.150 38.680 52.470 ;
        RECT 39.800 52.150 40.060 52.470 ;
        RECT 35.200 50.110 35.460 50.430 ;
        RECT 37.960 50.110 38.220 50.430 ;
        RECT 34.740 47.730 35.000 48.050 ;
        RECT 35.260 47.370 35.400 50.110 ;
        RECT 36.120 49.770 36.380 50.090 ;
        RECT 35.200 47.050 35.460 47.370 ;
        RECT 35.200 46.370 35.460 46.690 ;
        RECT 34.740 44.670 35.000 44.990 ;
        RECT 34.800 41.930 34.940 44.670 ;
        RECT 35.260 42.950 35.400 46.370 ;
        RECT 35.200 42.630 35.460 42.950 ;
        RECT 34.740 41.610 35.000 41.930 ;
        RECT 34.280 39.910 34.540 40.230 ;
        RECT 34.800 39.630 34.940 41.610 ;
        RECT 36.180 41.590 36.320 49.770 ;
        RECT 38.020 48.050 38.160 50.110 ;
        RECT 38.480 49.750 38.620 52.150 ;
        RECT 40.320 50.090 40.460 54.870 ;
        RECT 44.920 52.810 45.060 59.970 ;
        RECT 44.860 52.490 45.120 52.810 ;
        RECT 40.260 49.770 40.520 50.090 ;
        RECT 38.420 49.430 38.680 49.750 ;
        RECT 37.960 47.730 38.220 48.050 ;
        RECT 38.020 47.370 38.160 47.730 ;
        RECT 37.040 47.280 37.300 47.370 ;
        RECT 37.040 47.140 37.700 47.280 ;
        RECT 37.040 47.050 37.300 47.140 ;
        RECT 36.580 46.370 36.840 46.690 ;
        RECT 37.040 46.370 37.300 46.690 ;
        RECT 36.640 45.070 36.780 46.370 ;
        RECT 37.100 45.670 37.240 46.370 ;
        RECT 37.560 45.670 37.700 47.140 ;
        RECT 37.960 47.050 38.220 47.370 ;
        RECT 37.040 45.350 37.300 45.670 ;
        RECT 37.500 45.350 37.760 45.670 ;
        RECT 38.020 45.070 38.160 47.050 ;
        RECT 36.640 44.930 38.160 45.070 ;
        RECT 38.480 44.990 38.620 49.430 ;
        RECT 40.260 47.050 40.520 47.370 ;
        RECT 40.320 46.690 40.460 47.050 ;
        RECT 41.180 46.710 41.440 47.030 ;
        RECT 40.260 46.370 40.520 46.690 ;
        RECT 36.640 43.970 36.780 44.930 ;
        RECT 38.420 44.670 38.680 44.990 ;
        RECT 36.580 43.650 36.840 43.970 ;
        RECT 39.800 43.650 40.060 43.970 ;
        RECT 37.500 42.630 37.760 42.950 ;
        RECT 36.120 41.270 36.380 41.590 ;
        RECT 34.340 39.490 34.940 39.630 ;
        RECT 30.140 38.210 30.400 38.530 ;
        RECT 30.600 38.210 30.860 38.530 ;
        RECT 33.820 38.210 34.080 38.530 ;
        RECT 27.650 37.675 29.190 38.045 ;
        RECT 20.020 36.850 20.280 37.170 ;
        RECT 26.920 36.850 27.180 37.170 ;
        RECT 30.200 36.150 30.340 38.210 ;
        RECT 33.880 36.150 34.020 38.210 ;
        RECT 30.140 35.830 30.400 36.150 ;
        RECT 33.820 35.830 34.080 36.150 ;
        RECT 34.340 35.810 34.480 39.490 ;
        RECT 37.560 38.870 37.700 42.630 ;
        RECT 39.860 39.210 40.000 43.650 ;
        RECT 40.320 42.950 40.460 46.370 ;
        RECT 40.260 42.630 40.520 42.950 ;
        RECT 40.320 39.550 40.460 42.630 ;
        RECT 41.240 41.930 41.380 46.710 ;
        RECT 42.100 46.370 42.360 46.690 ;
        RECT 41.640 44.670 41.900 44.990 ;
        RECT 41.700 42.950 41.840 44.670 ;
        RECT 41.640 42.630 41.900 42.950 ;
        RECT 41.180 41.610 41.440 41.930 ;
        RECT 41.240 40.230 41.380 41.610 ;
        RECT 42.160 41.590 42.300 46.370 ;
        RECT 42.100 41.270 42.360 41.590 ;
        RECT 41.180 39.910 41.440 40.230 ;
        RECT 40.260 39.230 40.520 39.550 ;
        RECT 39.800 38.890 40.060 39.210 ;
        RECT 37.500 38.550 37.760 38.870 ;
        RECT 41.240 37.510 41.380 39.910 ;
        RECT 45.380 38.385 45.520 69.970 ;
        RECT 46.760 69.130 46.900 71.870 ;
        RECT 47.220 71.170 47.360 77.650 ;
        RECT 48.140 77.630 48.280 79.010 ;
        RECT 48.080 77.310 48.340 77.630 ;
        RECT 47.620 74.250 47.880 74.570 ;
        RECT 48.080 74.250 48.340 74.570 ;
        RECT 47.680 72.190 47.820 74.250 ;
        RECT 48.140 72.870 48.280 74.250 ;
        RECT 48.080 72.550 48.340 72.870 ;
        RECT 47.620 71.870 47.880 72.190 ;
        RECT 47.620 71.190 47.880 71.510 ;
        RECT 47.160 70.850 47.420 71.170 ;
        RECT 47.680 70.110 47.820 71.190 ;
        RECT 48.080 70.850 48.340 71.170 ;
        RECT 47.220 69.970 47.820 70.110 ;
        RECT 46.700 68.810 46.960 69.130 ;
        RECT 46.240 66.660 46.500 66.750 ;
        RECT 46.760 66.660 46.900 68.810 ;
        RECT 46.240 66.520 46.900 66.660 ;
        RECT 46.240 66.430 46.500 66.520 ;
        RECT 47.220 63.010 47.360 69.970 ;
        RECT 48.140 67.090 48.280 70.850 ;
        RECT 48.080 66.770 48.340 67.090 ;
        RECT 48.600 66.750 48.740 79.350 ;
        RECT 48.540 66.430 48.800 66.750 ;
        RECT 49.520 64.710 49.660 79.690 ;
        RECT 52.280 78.310 52.420 88.190 ;
        RECT 52.740 82.730 52.880 106.550 ;
        RECT 53.200 102.870 53.340 107.570 ;
        RECT 53.600 107.230 53.860 107.550 ;
        RECT 53.660 103.810 53.800 107.230 ;
        RECT 56.880 107.210 57.020 119.810 ;
        RECT 57.340 113.330 57.480 123.550 ;
        RECT 58.260 118.410 58.400 124.375 ;
        RECT 58.720 121.150 58.860 137.150 ;
        RECT 59.640 137.130 59.780 144.630 ;
        RECT 60.500 140.550 60.760 140.870 ;
        RECT 60.040 139.190 60.300 139.510 ;
        RECT 60.100 138.150 60.240 139.190 ;
        RECT 60.560 138.150 60.700 140.550 ;
        RECT 60.040 137.830 60.300 138.150 ;
        RECT 60.500 137.830 60.760 138.150 ;
        RECT 59.580 136.810 59.840 137.130 ;
        RECT 60.040 129.670 60.300 129.990 ;
        RECT 60.100 129.310 60.240 129.670 ;
        RECT 59.580 128.990 59.840 129.310 ;
        RECT 60.040 128.990 60.300 129.310 ;
        RECT 59.640 127.270 59.780 128.990 ;
        RECT 59.580 126.950 59.840 127.270 ;
        RECT 59.640 126.590 59.780 126.950 ;
        RECT 59.120 126.270 59.380 126.590 ;
        RECT 59.580 126.270 59.840 126.590 ;
        RECT 59.180 124.550 59.320 126.270 ;
        RECT 59.120 124.230 59.380 124.550 ;
        RECT 60.040 123.210 60.300 123.530 ;
        RECT 59.580 122.530 59.840 122.850 ;
        RECT 59.640 121.150 59.780 122.530 ;
        RECT 58.660 120.830 58.920 121.150 ;
        RECT 59.580 120.830 59.840 121.150 ;
        RECT 59.120 120.490 59.380 120.810 ;
        RECT 59.180 118.680 59.320 120.490 ;
        RECT 59.580 118.680 59.840 118.770 ;
        RECT 59.180 118.540 59.840 118.680 ;
        RECT 58.660 118.410 58.920 118.430 ;
        RECT 58.260 118.270 58.920 118.410 ;
        RECT 58.660 118.110 58.920 118.270 ;
        RECT 58.200 117.770 58.460 118.090 ;
        RECT 57.740 117.430 58.000 117.750 ;
        RECT 57.800 116.050 57.940 117.430 ;
        RECT 57.740 115.730 58.000 116.050 ;
        RECT 57.280 113.010 57.540 113.330 ;
        RECT 55.900 106.890 56.160 107.210 ;
        RECT 56.820 106.890 57.080 107.210 ;
        RECT 54.060 106.210 54.320 106.530 ;
        RECT 54.120 105.170 54.260 106.210 ;
        RECT 54.060 104.850 54.320 105.170 ;
        RECT 55.960 104.610 56.100 106.890 ;
        RECT 56.880 104.610 57.020 106.890 ;
        RECT 55.960 104.470 56.560 104.610 ;
        RECT 56.880 104.470 57.480 104.610 ;
        RECT 56.420 103.810 56.560 104.470 ;
        RECT 56.820 103.830 57.080 104.150 ;
        RECT 53.600 103.720 53.860 103.810 ;
        RECT 53.600 103.580 54.260 103.720 ;
        RECT 53.600 103.490 53.860 103.580 ;
        RECT 53.200 102.730 53.800 102.870 ;
        RECT 53.140 101.110 53.400 101.430 ;
        RECT 53.200 94.630 53.340 101.110 ;
        RECT 53.660 98.370 53.800 102.730 ;
        RECT 54.120 101.770 54.260 103.580 ;
        RECT 56.360 103.490 56.620 103.810 ;
        RECT 56.420 102.450 56.560 103.490 ;
        RECT 56.880 102.790 57.020 103.830 ;
        RECT 56.820 102.470 57.080 102.790 ;
        RECT 55.440 102.130 55.700 102.450 ;
        RECT 56.360 102.130 56.620 102.450 ;
        RECT 54.980 101.790 55.240 102.110 ;
        RECT 54.060 101.450 54.320 101.770 ;
        RECT 54.520 101.450 54.780 101.770 ;
        RECT 54.120 98.790 54.260 101.450 ;
        RECT 54.580 99.730 54.720 101.450 ;
        RECT 54.520 99.410 54.780 99.730 ;
        RECT 55.040 99.390 55.180 101.790 ;
        RECT 55.500 101.090 55.640 102.130 ;
        RECT 56.420 101.430 56.560 102.130 ;
        RECT 56.360 101.110 56.620 101.430 ;
        RECT 55.440 100.770 55.700 101.090 ;
        RECT 54.980 99.300 55.240 99.390 ;
        RECT 55.900 99.300 56.160 99.390 ;
        RECT 56.420 99.300 56.560 101.110 ;
        RECT 57.340 100.070 57.480 104.470 ;
        RECT 57.280 99.750 57.540 100.070 ;
        RECT 54.980 99.160 55.640 99.300 ;
        RECT 54.980 99.070 55.240 99.160 ;
        RECT 54.120 98.650 54.720 98.790 ;
        RECT 54.580 98.370 54.720 98.650 ;
        RECT 53.600 98.050 53.860 98.370 ;
        RECT 54.520 98.050 54.780 98.370 ;
        RECT 53.140 94.310 53.400 94.630 ;
        RECT 53.200 91.910 53.340 94.310 ;
        RECT 53.660 93.950 53.800 98.050 ;
        RECT 53.600 93.630 53.860 93.950 ;
        RECT 53.140 91.590 53.400 91.910 ;
        RECT 53.130 90.375 53.410 90.745 ;
        RECT 53.600 90.570 53.860 90.890 ;
        RECT 53.200 90.210 53.340 90.375 ;
        RECT 53.140 89.890 53.400 90.210 ;
        RECT 53.660 89.190 53.800 90.570 ;
        RECT 54.060 89.890 54.320 90.210 ;
        RECT 53.600 88.870 53.860 89.190 ;
        RECT 53.660 85.360 53.800 88.870 ;
        RECT 54.120 87.910 54.260 89.890 ;
        RECT 54.580 89.190 54.720 98.050 ;
        RECT 54.980 93.290 55.240 93.610 ;
        RECT 54.520 88.870 54.780 89.190 ;
        RECT 54.510 88.335 54.790 88.705 ;
        RECT 55.040 88.510 55.180 93.290 ;
        RECT 55.500 91.910 55.640 99.160 ;
        RECT 55.900 99.160 56.560 99.300 ;
        RECT 55.900 99.070 56.160 99.160 ;
        RECT 55.900 98.390 56.160 98.710 ;
        RECT 55.960 94.290 56.100 98.390 ;
        RECT 55.900 93.970 56.160 94.290 ;
        RECT 55.440 91.820 55.700 91.910 ;
        RECT 55.440 91.680 56.100 91.820 ;
        RECT 55.440 91.590 55.700 91.680 ;
        RECT 55.440 90.910 55.700 91.230 ;
        RECT 55.500 89.190 55.640 90.910 ;
        RECT 55.440 88.870 55.700 89.190 ;
        RECT 54.520 88.190 54.780 88.335 ;
        RECT 54.980 88.190 55.240 88.510 ;
        RECT 54.120 87.770 55.180 87.910 ;
        RECT 55.040 86.470 55.180 87.770 ;
        RECT 55.500 86.470 55.640 88.870 ;
        RECT 54.980 86.150 55.240 86.470 ;
        RECT 55.440 86.150 55.700 86.470 ;
        RECT 54.060 85.360 54.320 85.450 ;
        RECT 53.660 85.220 54.320 85.360 ;
        RECT 54.060 85.130 54.320 85.220 ;
        RECT 53.140 84.450 53.400 84.770 ;
        RECT 52.680 82.410 52.940 82.730 ;
        RECT 52.740 80.350 52.880 82.410 ;
        RECT 52.680 80.030 52.940 80.350 ;
        RECT 52.220 77.990 52.480 78.310 ;
        RECT 53.200 71.850 53.340 84.450 ;
        RECT 54.060 81.730 54.320 82.050 ;
        RECT 54.120 80.690 54.260 81.730 ;
        RECT 55.040 80.690 55.180 86.150 ;
        RECT 55.440 85.305 55.700 85.450 ;
        RECT 55.430 84.935 55.710 85.305 ;
        RECT 55.440 84.450 55.700 84.770 ;
        RECT 54.060 80.370 54.320 80.690 ;
        RECT 54.980 80.370 55.240 80.690 ;
        RECT 54.120 77.630 54.260 80.370 ;
        RECT 55.500 79.865 55.640 84.450 ;
        RECT 55.960 83.750 56.100 91.680 ;
        RECT 56.420 90.890 56.560 99.160 ;
        RECT 57.800 97.350 57.940 115.730 ;
        RECT 58.260 113.330 58.400 117.770 ;
        RECT 58.720 116.050 58.860 118.110 ;
        RECT 58.660 115.730 58.920 116.050 ;
        RECT 59.180 115.280 59.320 118.540 ;
        RECT 59.580 118.450 59.840 118.540 ;
        RECT 58.720 115.140 59.320 115.280 ;
        RECT 58.200 113.010 58.460 113.330 ;
        RECT 58.200 112.330 58.460 112.650 ;
        RECT 58.260 110.950 58.400 112.330 ;
        RECT 58.200 110.630 58.460 110.950 ;
        RECT 58.720 110.270 58.860 115.140 ;
        RECT 59.580 112.330 59.840 112.650 ;
        RECT 59.120 110.290 59.380 110.610 ;
        RECT 58.660 109.950 58.920 110.270 ;
        RECT 59.180 106.530 59.320 110.290 ;
        RECT 59.120 106.210 59.380 106.530 ;
        RECT 58.200 104.170 58.460 104.490 ;
        RECT 58.260 102.790 58.400 104.170 ;
        RECT 58.200 102.470 58.460 102.790 ;
        RECT 58.260 99.730 58.400 102.470 ;
        RECT 58.660 101.450 58.920 101.770 ;
        RECT 58.200 99.410 58.460 99.730 ;
        RECT 57.740 97.030 58.000 97.350 ;
        RECT 57.280 90.910 57.540 91.230 ;
        RECT 56.360 90.570 56.620 90.890 ;
        RECT 56.820 90.230 57.080 90.550 ;
        RECT 56.360 89.890 56.620 90.210 ;
        RECT 56.420 88.170 56.560 89.890 ;
        RECT 56.880 88.705 57.020 90.230 ;
        RECT 57.340 88.850 57.480 90.910 ;
        RECT 56.810 88.335 57.090 88.705 ;
        RECT 57.280 88.530 57.540 88.850 ;
        RECT 56.360 87.850 56.620 88.170 ;
        RECT 57.280 87.850 57.540 88.170 ;
        RECT 56.360 87.170 56.620 87.490 ;
        RECT 56.820 87.170 57.080 87.490 ;
        RECT 56.420 86.470 56.560 87.170 ;
        RECT 56.360 86.150 56.620 86.470 ;
        RECT 56.350 85.615 56.630 85.985 ;
        RECT 56.420 85.450 56.560 85.615 ;
        RECT 56.360 85.130 56.620 85.450 ;
        RECT 55.900 83.430 56.160 83.750 ;
        RECT 55.960 82.390 56.100 83.430 ;
        RECT 55.900 82.070 56.160 82.390 ;
        RECT 56.420 80.350 56.560 85.130 ;
        RECT 56.360 80.030 56.620 80.350 ;
        RECT 55.430 79.495 55.710 79.865 ;
        RECT 54.060 77.310 54.320 77.630 ;
        RECT 54.980 74.250 55.240 74.570 ;
        RECT 52.220 71.530 52.480 71.850 ;
        RECT 53.140 71.530 53.400 71.850 ;
        RECT 52.280 70.150 52.420 71.530 ;
        RECT 52.220 69.830 52.480 70.150 ;
        RECT 52.210 69.295 52.490 69.665 ;
        RECT 52.280 69.130 52.420 69.295 ;
        RECT 52.220 68.810 52.480 69.130 ;
        RECT 49.920 68.130 50.180 68.450 ;
        RECT 51.760 68.130 52.020 68.450 ;
        RECT 49.980 67.430 50.120 68.130 ;
        RECT 49.920 67.110 50.180 67.430 ;
        RECT 50.840 66.090 51.100 66.410 ;
        RECT 49.460 64.390 49.720 64.710 ;
        RECT 50.900 63.350 51.040 66.090 ;
        RECT 51.300 64.390 51.560 64.710 ;
        RECT 50.840 63.030 51.100 63.350 ;
        RECT 47.160 62.690 47.420 63.010 ;
        RECT 50.380 62.690 50.640 63.010 ;
        RECT 47.220 60.030 47.360 62.690 ;
        RECT 49.920 61.330 50.180 61.650 ;
        RECT 49.460 60.650 49.720 60.970 ;
        RECT 47.620 60.310 47.880 60.630 ;
        RECT 46.300 59.890 47.360 60.030 ;
        RECT 46.300 59.270 46.440 59.890 ;
        RECT 46.240 58.950 46.500 59.270 ;
        RECT 47.160 58.610 47.420 58.930 ;
        RECT 47.220 50.770 47.360 58.610 ;
        RECT 47.160 50.450 47.420 50.770 ;
        RECT 47.680 44.650 47.820 60.310 ;
        RECT 49.000 59.970 49.260 60.290 ;
        RECT 49.060 58.590 49.200 59.970 ;
        RECT 49.000 58.270 49.260 58.590 ;
        RECT 49.520 58.250 49.660 60.650 ;
        RECT 49.980 59.270 50.120 61.330 ;
        RECT 50.440 59.270 50.580 62.690 ;
        RECT 50.840 60.650 51.100 60.970 ;
        RECT 49.920 58.950 50.180 59.270 ;
        RECT 50.380 58.950 50.640 59.270 ;
        RECT 48.080 57.930 48.340 58.250 ;
        RECT 49.460 57.930 49.720 58.250 ;
        RECT 48.140 53.150 48.280 57.930 ;
        RECT 49.520 57.310 49.660 57.930 ;
        RECT 49.060 57.170 49.660 57.310 ;
        RECT 48.540 55.210 48.800 55.530 ;
        RECT 48.600 53.830 48.740 55.210 ;
        RECT 48.540 53.510 48.800 53.830 ;
        RECT 48.080 52.830 48.340 53.150 ;
        RECT 48.540 52.150 48.800 52.470 ;
        RECT 48.080 51.810 48.340 52.130 ;
        RECT 48.140 44.990 48.280 51.810 ;
        RECT 48.600 48.390 48.740 52.150 ;
        RECT 49.060 51.110 49.200 57.170 ;
        RECT 49.460 56.230 49.720 56.550 ;
        RECT 49.520 53.830 49.660 56.230 ;
        RECT 49.980 55.870 50.120 58.950 ;
        RECT 50.380 57.250 50.640 57.570 ;
        RECT 49.920 55.550 50.180 55.870 ;
        RECT 49.460 53.510 49.720 53.830 ;
        RECT 49.000 51.020 49.260 51.110 ;
        RECT 49.000 50.880 49.660 51.020 ;
        RECT 49.000 50.790 49.260 50.880 ;
        RECT 49.000 50.110 49.260 50.430 ;
        RECT 48.540 48.070 48.800 48.390 ;
        RECT 49.060 45.670 49.200 50.110 ;
        RECT 49.520 47.710 49.660 50.880 ;
        RECT 49.460 47.390 49.720 47.710 ;
        RECT 49.000 45.350 49.260 45.670 ;
        RECT 50.440 44.990 50.580 57.250 ;
        RECT 48.080 44.670 48.340 44.990 ;
        RECT 50.380 44.670 50.640 44.990 ;
        RECT 47.620 44.330 47.880 44.650 ;
        RECT 49.920 44.390 50.180 44.650 ;
        RECT 50.900 44.390 51.040 60.650 ;
        RECT 51.360 48.390 51.500 64.390 ;
        RECT 51.820 63.350 51.960 68.130 ;
        RECT 53.140 66.430 53.400 66.750 ;
        RECT 54.060 66.430 54.320 66.750 ;
        RECT 52.680 65.585 52.940 65.730 ;
        RECT 52.670 65.215 52.950 65.585 ;
        RECT 52.220 64.390 52.480 64.710 ;
        RECT 51.760 63.030 52.020 63.350 ;
        RECT 52.280 63.010 52.420 64.390 ;
        RECT 52.680 63.430 52.940 63.690 ;
        RECT 53.200 63.430 53.340 66.430 ;
        RECT 54.120 63.690 54.260 66.430 ;
        RECT 55.040 64.370 55.180 74.250 ;
        RECT 55.500 73.890 55.640 79.495 ;
        RECT 55.890 74.735 56.170 75.105 ;
        RECT 55.960 74.570 56.100 74.735 ;
        RECT 56.420 74.570 56.560 80.030 ;
        RECT 55.900 74.250 56.160 74.570 ;
        RECT 56.360 74.250 56.620 74.570 ;
        RECT 55.440 73.570 55.700 73.890 ;
        RECT 55.500 69.470 55.640 73.570 ;
        RECT 56.360 71.530 56.620 71.850 ;
        RECT 55.900 71.190 56.160 71.510 ;
        RECT 55.960 69.665 56.100 71.190 ;
        RECT 55.440 69.150 55.700 69.470 ;
        RECT 55.890 69.295 56.170 69.665 ;
        RECT 55.960 67.090 56.100 69.295 ;
        RECT 55.900 66.770 56.160 67.090 ;
        RECT 56.420 65.730 56.560 71.530 ;
        RECT 56.880 69.130 57.020 87.170 ;
        RECT 57.340 85.450 57.480 87.850 ;
        RECT 57.280 85.130 57.540 85.450 ;
        RECT 57.280 82.070 57.540 82.390 ;
        RECT 57.340 77.630 57.480 82.070 ;
        RECT 57.800 77.970 57.940 97.030 ;
        RECT 58.200 93.970 58.460 94.290 ;
        RECT 58.260 87.490 58.400 93.970 ;
        RECT 58.720 90.890 58.860 101.450 ;
        RECT 59.180 100.070 59.320 106.210 ;
        RECT 59.640 104.150 59.780 112.330 ;
        RECT 60.100 106.870 60.240 123.210 ;
        RECT 60.500 120.830 60.760 121.150 ;
        RECT 60.560 119.110 60.700 120.830 ;
        RECT 60.500 118.790 60.760 119.110 ;
        RECT 60.500 117.090 60.760 117.410 ;
        RECT 60.560 115.710 60.700 117.090 ;
        RECT 61.020 116.390 61.160 147.690 ;
        RECT 62.400 145.630 62.540 147.690 ;
        RECT 62.340 145.310 62.600 145.630 ;
        RECT 62.860 144.610 63.000 150.895 ;
        RECT 62.800 144.290 63.060 144.610 ;
        RECT 62.800 141.910 63.060 142.230 ;
        RECT 61.870 140.695 62.150 141.065 ;
        RECT 61.420 136.470 61.680 136.790 ;
        RECT 61.480 132.905 61.620 136.470 ;
        RECT 61.940 135.430 62.080 140.695 ;
        RECT 61.880 135.110 62.140 135.430 ;
        RECT 62.860 134.410 63.000 141.910 ;
        RECT 63.320 134.750 63.460 158.570 ;
        RECT 63.780 156.170 63.920 166.650 ;
        RECT 64.180 166.050 64.440 166.370 ;
        RECT 64.240 159.910 64.380 166.050 ;
        RECT 64.180 159.590 64.440 159.910 ;
        RECT 65.160 156.170 65.300 167.215 ;
        RECT 66.540 164.070 66.680 168.575 ;
        RECT 67.000 165.350 67.140 169.450 ;
        RECT 66.940 165.030 67.200 165.350 ;
        RECT 66.540 163.930 67.140 164.070 ;
        RECT 66.020 163.330 66.280 163.650 ;
        RECT 66.480 163.330 66.740 163.650 ;
        RECT 66.080 162.630 66.220 163.330 ;
        RECT 66.020 162.310 66.280 162.630 ;
        RECT 65.560 160.950 65.820 161.270 ;
        RECT 65.620 156.850 65.760 160.950 ;
        RECT 66.080 159.910 66.220 162.310 ;
        RECT 66.020 159.590 66.280 159.910 ;
        RECT 66.540 159.310 66.680 163.330 ;
        RECT 66.080 159.170 66.680 159.310 ;
        RECT 65.560 156.530 65.820 156.850 ;
        RECT 63.720 155.850 63.980 156.170 ;
        RECT 64.640 155.850 64.900 156.170 ;
        RECT 65.100 155.850 65.360 156.170 ;
        RECT 64.700 155.345 64.840 155.850 ;
        RECT 64.630 154.975 64.910 155.345 ;
        RECT 64.640 154.150 64.900 154.470 ;
        RECT 64.180 152.450 64.440 152.770 ;
        RECT 64.240 150.730 64.380 152.450 ;
        RECT 64.700 150.730 64.840 154.150 ;
        RECT 64.180 150.410 64.440 150.730 ;
        RECT 64.640 150.410 64.900 150.730 ;
        RECT 64.700 146.310 64.840 150.410 ;
        RECT 64.640 145.990 64.900 146.310 ;
        RECT 66.080 145.630 66.220 159.170 ;
        RECT 67.000 155.230 67.140 163.930 ;
        RECT 67.400 157.890 67.660 158.210 ;
        RECT 67.460 156.170 67.600 157.890 ;
        RECT 67.920 156.850 68.060 171.490 ;
        RECT 69.230 171.295 69.510 171.665 ;
        RECT 72.460 171.490 72.720 171.810 ;
        RECT 68.320 164.350 68.580 164.670 ;
        RECT 68.380 159.910 68.520 164.350 ;
        RECT 68.780 160.610 69.040 160.930 ;
        RECT 68.320 159.590 68.580 159.910 ;
        RECT 68.320 158.230 68.580 158.550 ;
        RECT 67.860 156.530 68.120 156.850 ;
        RECT 68.380 156.510 68.520 158.230 ;
        RECT 68.320 156.190 68.580 156.510 ;
        RECT 67.400 155.850 67.660 156.170 ;
        RECT 67.000 155.090 68.520 155.230 ;
        RECT 67.860 153.130 68.120 153.450 ;
        RECT 67.920 150.730 68.060 153.130 ;
        RECT 67.860 150.410 68.120 150.730 ;
        RECT 66.480 148.710 66.740 149.030 ;
        RECT 66.020 145.310 66.280 145.630 ;
        RECT 66.020 144.290 66.280 144.610 ;
        RECT 65.550 139.335 65.830 139.705 ;
        RECT 65.620 139.170 65.760 139.335 ;
        RECT 65.560 138.850 65.820 139.170 ;
        RECT 65.100 137.150 65.360 137.470 ;
        RECT 63.260 134.430 63.520 134.750 ;
        RECT 62.800 134.090 63.060 134.410 ;
        RECT 61.410 132.535 61.690 132.905 ;
        RECT 63.320 132.710 63.460 134.430 ;
        RECT 63.260 132.390 63.520 132.710 ;
        RECT 62.800 131.710 63.060 132.030 ;
        RECT 64.640 131.710 64.900 132.030 ;
        RECT 61.880 129.330 62.140 129.650 ;
        RECT 61.420 128.030 61.680 128.290 ;
        RECT 61.940 128.030 62.080 129.330 ;
        RECT 61.420 127.970 62.080 128.030 ;
        RECT 62.340 127.970 62.600 128.290 ;
        RECT 61.480 127.890 62.080 127.970 ;
        RECT 61.420 125.930 61.680 126.250 ;
        RECT 61.480 123.530 61.620 125.930 ;
        RECT 61.880 125.250 62.140 125.570 ;
        RECT 61.940 124.550 62.080 125.250 ;
        RECT 61.880 124.230 62.140 124.550 ;
        RECT 61.420 123.210 61.680 123.530 ;
        RECT 61.940 121.490 62.080 124.230 ;
        RECT 62.400 122.850 62.540 127.970 ;
        RECT 62.860 125.910 63.000 131.710 ;
        RECT 64.180 131.370 64.440 131.690 ;
        RECT 63.720 130.690 63.980 131.010 ;
        RECT 63.780 129.310 63.920 130.690 ;
        RECT 63.720 128.990 63.980 129.310 ;
        RECT 63.260 128.650 63.520 128.970 ;
        RECT 63.320 128.290 63.460 128.650 ;
        RECT 63.260 127.970 63.520 128.290 ;
        RECT 63.720 127.970 63.980 128.290 ;
        RECT 63.780 127.180 63.920 127.970 ;
        RECT 63.320 127.040 63.920 127.180 ;
        RECT 62.800 125.590 63.060 125.910 ;
        RECT 62.790 125.055 63.070 125.425 ;
        RECT 62.860 124.550 63.000 125.055 ;
        RECT 62.800 124.230 63.060 124.550 ;
        RECT 63.320 123.950 63.460 127.040 ;
        RECT 64.240 126.930 64.380 131.370 ;
        RECT 64.180 126.610 64.440 126.930 ;
        RECT 63.720 126.270 63.980 126.590 ;
        RECT 62.860 123.810 63.460 123.950 ;
        RECT 62.860 123.530 63.000 123.810 ;
        RECT 62.800 123.210 63.060 123.530 ;
        RECT 63.260 123.210 63.520 123.530 ;
        RECT 62.340 122.530 62.600 122.850 ;
        RECT 61.880 121.170 62.140 121.490 ;
        RECT 61.420 120.830 61.680 121.150 ;
        RECT 60.960 116.070 61.220 116.390 ;
        RECT 60.500 115.390 60.760 115.710 ;
        RECT 61.020 113.330 61.160 116.070 ;
        RECT 60.960 113.010 61.220 113.330 ;
        RECT 60.500 112.330 60.760 112.650 ;
        RECT 60.560 108.230 60.700 112.330 ;
        RECT 61.480 112.310 61.620 120.830 ;
        RECT 62.400 115.370 62.540 122.530 ;
        RECT 62.800 115.730 63.060 116.050 ;
        RECT 62.340 115.050 62.600 115.370 ;
        RECT 61.420 111.990 61.680 112.310 ;
        RECT 61.880 111.650 62.140 111.970 ;
        RECT 61.940 110.270 62.080 111.650 ;
        RECT 61.880 109.950 62.140 110.270 ;
        RECT 60.960 109.610 61.220 109.930 ;
        RECT 60.500 107.910 60.760 108.230 ;
        RECT 60.500 106.890 60.760 107.210 ;
        RECT 60.040 106.550 60.300 106.870 ;
        RECT 60.100 105.510 60.240 106.550 ;
        RECT 60.040 105.190 60.300 105.510 ;
        RECT 60.040 104.510 60.300 104.830 ;
        RECT 59.580 103.830 59.840 104.150 ;
        RECT 59.580 101.110 59.840 101.430 ;
        RECT 59.120 99.750 59.380 100.070 ;
        RECT 59.180 91.570 59.320 99.750 ;
        RECT 59.640 99.390 59.780 101.110 ;
        RECT 60.100 101.090 60.240 104.510 ;
        RECT 60.040 100.770 60.300 101.090 ;
        RECT 59.580 99.070 59.840 99.390 ;
        RECT 59.640 98.370 59.780 99.070 ;
        RECT 60.040 98.730 60.300 99.050 ;
        RECT 59.580 98.050 59.840 98.370 ;
        RECT 60.100 93.610 60.240 98.730 ;
        RECT 60.560 94.630 60.700 106.890 ;
        RECT 61.020 105.510 61.160 109.610 ;
        RECT 61.880 109.270 62.140 109.590 ;
        RECT 61.420 108.930 61.680 109.250 ;
        RECT 60.960 105.190 61.220 105.510 ;
        RECT 61.020 102.110 61.160 105.190 ;
        RECT 60.960 101.790 61.220 102.110 ;
        RECT 61.480 101.680 61.620 108.930 ;
        RECT 61.940 107.210 62.080 109.270 ;
        RECT 61.880 106.890 62.140 107.210 ;
        RECT 61.880 106.210 62.140 106.530 ;
        RECT 61.940 105.510 62.080 106.210 ;
        RECT 61.880 105.190 62.140 105.510 ;
        RECT 62.400 104.830 62.540 115.050 ;
        RECT 62.860 110.950 63.000 115.730 ;
        RECT 63.320 115.370 63.460 123.210 ;
        RECT 63.780 115.710 63.920 126.270 ;
        RECT 64.240 121.150 64.380 126.610 ;
        RECT 64.700 124.550 64.840 131.710 ;
        RECT 65.160 128.970 65.300 137.150 ;
        RECT 66.080 136.450 66.220 144.290 ;
        RECT 66.540 140.530 66.680 148.710 ;
        RECT 67.920 148.690 68.060 150.410 ;
        RECT 67.860 148.370 68.120 148.690 ;
        RECT 67.860 145.990 68.120 146.310 ;
        RECT 67.920 143.590 68.060 145.990 ;
        RECT 67.860 143.270 68.120 143.590 ;
        RECT 66.480 140.270 66.740 140.530 ;
        RECT 66.480 140.210 67.140 140.270 ;
        RECT 66.540 140.130 67.140 140.210 ;
        RECT 67.000 137.810 67.140 140.130 ;
        RECT 66.940 137.490 67.200 137.810 ;
        RECT 66.020 136.130 66.280 136.450 ;
        RECT 66.480 134.430 66.740 134.750 ;
        RECT 66.540 129.650 66.680 134.430 ;
        RECT 66.940 133.410 67.200 133.730 ;
        RECT 67.400 133.410 67.660 133.730 ;
        RECT 67.860 133.410 68.120 133.730 ;
        RECT 66.480 129.330 66.740 129.650 ;
        RECT 65.100 128.880 65.360 128.970 ;
        RECT 65.100 128.740 65.760 128.880 ;
        RECT 65.100 128.650 65.360 128.740 ;
        RECT 65.100 127.970 65.360 128.290 ;
        RECT 65.160 125.425 65.300 127.970 ;
        RECT 65.090 125.055 65.370 125.425 ;
        RECT 64.640 124.230 64.900 124.550 ;
        RECT 64.640 123.590 64.900 123.910 ;
        RECT 64.180 120.830 64.440 121.150 ;
        RECT 64.240 117.750 64.380 120.830 ;
        RECT 64.700 119.110 64.840 123.590 ;
        RECT 64.640 118.790 64.900 119.110 ;
        RECT 65.160 118.410 65.300 125.055 ;
        RECT 65.620 124.745 65.760 128.740 ;
        RECT 66.470 128.455 66.750 128.825 ;
        RECT 66.540 126.930 66.680 128.455 ;
        RECT 66.480 126.610 66.740 126.930 ;
        RECT 66.020 126.270 66.280 126.590 ;
        RECT 65.550 124.375 65.830 124.745 ;
        RECT 66.080 124.550 66.220 126.270 ;
        RECT 66.020 124.230 66.280 124.550 ;
        RECT 66.540 123.950 66.680 126.610 ;
        RECT 67.000 126.590 67.140 133.410 ;
        RECT 67.460 130.865 67.600 133.410 ;
        RECT 67.390 130.495 67.670 130.865 ;
        RECT 67.920 129.990 68.060 133.410 ;
        RECT 68.380 132.030 68.520 155.090 ;
        RECT 68.840 139.705 68.980 160.610 ;
        RECT 69.300 155.490 69.440 171.295 ;
        RECT 69.700 169.110 69.960 169.430 ;
        RECT 69.760 161.610 69.900 169.110 ;
        RECT 72.000 166.390 72.260 166.710 ;
        RECT 71.540 164.350 71.800 164.670 ;
        RECT 70.160 161.630 70.420 161.950 ;
        RECT 69.700 161.290 69.960 161.610 ;
        RECT 70.220 158.890 70.360 161.630 ;
        RECT 70.620 160.950 70.880 161.270 ;
        RECT 70.680 159.570 70.820 160.950 ;
        RECT 70.620 159.250 70.880 159.570 ;
        RECT 70.160 158.570 70.420 158.890 ;
        RECT 71.600 157.190 71.740 164.350 ;
        RECT 72.060 161.270 72.200 166.390 ;
        RECT 72.000 160.950 72.260 161.270 ;
        RECT 72.520 158.890 72.660 171.490 ;
        RECT 73.440 170.790 73.580 171.830 ;
        RECT 73.900 170.790 74.040 171.830 ;
        RECT 73.380 170.470 73.640 170.790 ;
        RECT 73.840 170.470 74.100 170.790 ;
        RECT 72.920 160.610 73.180 160.930 ;
        RECT 72.980 159.910 73.120 160.610 ;
        RECT 72.920 159.590 73.180 159.910 ;
        RECT 72.000 158.570 72.260 158.890 ;
        RECT 72.460 158.570 72.720 158.890 ;
        RECT 71.540 156.870 71.800 157.190 ;
        RECT 72.060 156.510 72.200 158.570 ;
        RECT 70.160 156.190 70.420 156.510 ;
        RECT 72.000 156.190 72.260 156.510 ;
        RECT 72.920 156.190 73.180 156.510 ;
        RECT 69.240 155.170 69.500 155.490 ;
        RECT 69.700 155.170 69.960 155.490 ;
        RECT 69.760 154.130 69.900 155.170 ;
        RECT 69.700 153.810 69.960 154.130 ;
        RECT 69.700 148.030 69.960 148.350 ;
        RECT 69.760 143.590 69.900 148.030 ;
        RECT 69.700 143.270 69.960 143.590 ;
        RECT 70.220 142.990 70.360 156.190 ;
        RECT 72.980 155.490 73.120 156.190 ;
        RECT 71.080 155.170 71.340 155.490 ;
        RECT 72.920 155.170 73.180 155.490 ;
        RECT 70.620 149.730 70.880 150.050 ;
        RECT 70.680 145.630 70.820 149.730 ;
        RECT 70.620 145.310 70.880 145.630 ;
        RECT 69.760 142.850 70.360 142.990 ;
        RECT 69.760 142.570 69.900 142.850 ;
        RECT 69.700 142.250 69.960 142.570 ;
        RECT 68.770 139.335 69.050 139.705 ;
        RECT 69.760 135.430 69.900 142.250 ;
        RECT 70.610 140.015 70.890 140.385 ;
        RECT 69.700 135.110 69.960 135.430 ;
        RECT 68.320 131.710 68.580 132.030 ;
        RECT 69.760 131.690 69.900 135.110 ;
        RECT 69.700 131.370 69.960 131.690 ;
        RECT 67.860 129.670 68.120 129.990 ;
        RECT 67.400 128.990 67.660 129.310 ;
        RECT 67.460 128.825 67.600 128.990 ;
        RECT 67.390 128.455 67.670 128.825 ;
        RECT 67.860 128.650 68.120 128.970 ;
        RECT 66.940 126.270 67.200 126.590 ;
        RECT 66.940 125.590 67.200 125.910 ;
        RECT 67.000 124.550 67.140 125.590 ;
        RECT 66.940 124.230 67.200 124.550 ;
        RECT 65.560 123.550 65.820 123.870 ;
        RECT 66.080 123.810 66.680 123.950 ;
        RECT 67.920 123.950 68.060 128.650 ;
        RECT 69.240 128.310 69.500 128.630 ;
        RECT 69.300 126.590 69.440 128.310 ;
        RECT 69.240 126.270 69.500 126.590 ;
        RECT 65.620 120.130 65.760 123.550 ;
        RECT 65.560 119.810 65.820 120.130 ;
        RECT 66.080 118.770 66.220 123.810 ;
        RECT 66.940 123.550 67.200 123.870 ;
        RECT 67.920 123.810 68.520 123.950 ;
        RECT 66.480 123.210 66.740 123.530 ;
        RECT 66.540 122.850 66.680 123.210 ;
        RECT 66.480 122.530 66.740 122.850 ;
        RECT 67.000 122.025 67.140 123.550 ;
        RECT 67.860 123.385 68.120 123.530 ;
        RECT 67.400 122.870 67.660 123.190 ;
        RECT 67.850 123.015 68.130 123.385 ;
        RECT 67.460 122.705 67.600 122.870 ;
        RECT 67.390 122.335 67.670 122.705 ;
        RECT 66.930 121.655 67.210 122.025 ;
        RECT 67.400 121.510 67.660 121.830 ;
        RECT 66.020 118.450 66.280 118.770 ;
        RECT 64.700 118.270 65.300 118.410 ;
        RECT 66.940 118.340 67.200 118.430 ;
        RECT 67.460 118.340 67.600 121.510 ;
        RECT 64.180 117.430 64.440 117.750 ;
        RECT 63.720 115.390 63.980 115.710 ;
        RECT 64.180 115.390 64.440 115.710 ;
        RECT 63.260 115.050 63.520 115.370 ;
        RECT 62.800 110.630 63.060 110.950 ;
        RECT 63.260 110.290 63.520 110.610 ;
        RECT 62.800 107.230 63.060 107.550 ;
        RECT 62.340 104.510 62.600 104.830 ;
        RECT 62.400 102.450 62.540 104.510 ;
        RECT 62.340 102.130 62.600 102.450 ;
        RECT 62.860 101.770 63.000 107.230 ;
        RECT 63.320 104.830 63.460 110.290 ;
        RECT 63.780 107.210 63.920 115.390 ;
        RECT 64.240 112.560 64.380 115.390 ;
        RECT 64.700 113.330 64.840 118.270 ;
        RECT 66.940 118.200 67.600 118.340 ;
        RECT 66.940 118.110 67.200 118.200 ;
        RECT 65.100 117.770 65.360 118.090 ;
        RECT 65.160 115.710 65.300 117.770 ;
        RECT 66.480 117.430 66.740 117.750 ;
        RECT 65.100 115.390 65.360 115.710 ;
        RECT 65.160 113.670 65.300 115.390 ;
        RECT 66.540 115.370 66.680 117.430 ;
        RECT 66.940 116.070 67.200 116.390 ;
        RECT 66.020 115.110 66.280 115.370 ;
        RECT 65.620 115.050 66.280 115.110 ;
        RECT 66.480 115.050 66.740 115.370 ;
        RECT 65.620 114.970 66.220 115.050 ;
        RECT 65.100 113.350 65.360 113.670 ;
        RECT 64.640 113.010 64.900 113.330 ;
        RECT 65.100 112.560 65.360 112.650 ;
        RECT 64.240 112.420 65.360 112.560 ;
        RECT 65.100 112.330 65.360 112.420 ;
        RECT 64.180 107.910 64.440 108.230 ;
        RECT 63.720 106.890 63.980 107.210 ;
        RECT 63.720 106.210 63.980 106.530 ;
        RECT 63.260 104.510 63.520 104.830 ;
        RECT 61.880 101.680 62.140 101.770 ;
        RECT 62.800 101.680 63.060 101.770 ;
        RECT 61.480 101.540 62.140 101.680 ;
        RECT 61.880 101.450 62.140 101.540 ;
        RECT 62.400 101.540 63.060 101.680 ;
        RECT 60.960 100.770 61.220 101.090 ;
        RECT 60.500 94.310 60.760 94.630 ;
        RECT 60.040 93.290 60.300 93.610 ;
        RECT 61.020 91.910 61.160 100.770 ;
        RECT 61.420 98.050 61.680 98.370 ;
        RECT 60.960 91.590 61.220 91.910 ;
        RECT 59.120 91.250 59.380 91.570 ;
        RECT 58.660 90.570 58.920 90.890 ;
        RECT 60.500 90.570 60.760 90.890 ;
        RECT 58.660 89.890 58.920 90.210 ;
        RECT 59.580 89.890 59.840 90.210 ;
        RECT 58.200 87.170 58.460 87.490 ;
        RECT 58.720 85.450 58.860 89.890 ;
        RECT 59.640 88.170 59.780 89.890 ;
        RECT 60.040 88.190 60.300 88.510 ;
        RECT 59.580 87.850 59.840 88.170 ;
        RECT 59.120 86.150 59.380 86.470 ;
        RECT 59.180 85.450 59.320 86.150 ;
        RECT 59.640 86.130 59.780 87.850 ;
        RECT 59.580 85.810 59.840 86.130 ;
        RECT 58.200 85.130 58.460 85.450 ;
        RECT 58.660 85.130 58.920 85.450 ;
        RECT 59.120 85.130 59.380 85.450 ;
        RECT 59.580 85.130 59.840 85.450 ;
        RECT 58.260 84.770 58.400 85.130 ;
        RECT 58.200 84.450 58.460 84.770 ;
        RECT 59.640 84.625 59.780 85.130 ;
        RECT 58.260 82.300 58.400 84.450 ;
        RECT 59.570 84.255 59.850 84.625 ;
        RECT 60.100 83.750 60.240 88.190 ;
        RECT 60.560 87.490 60.700 90.570 ;
        RECT 61.020 88.170 61.160 91.590 ;
        RECT 60.960 87.850 61.220 88.170 ;
        RECT 60.500 87.170 60.760 87.490 ;
        RECT 60.560 85.790 60.700 87.170 ;
        RECT 60.960 85.810 61.220 86.130 ;
        RECT 60.500 85.470 60.760 85.790 ;
        RECT 60.560 83.750 60.700 85.470 ;
        RECT 61.020 83.750 61.160 85.810 ;
        RECT 61.480 85.450 61.620 98.050 ;
        RECT 61.940 89.190 62.080 101.450 ;
        RECT 62.400 93.270 62.540 101.540 ;
        RECT 62.800 101.450 63.060 101.540 ;
        RECT 63.780 101.430 63.920 106.210 ;
        RECT 63.720 101.110 63.980 101.430 ;
        RECT 64.240 99.390 64.380 107.910 ;
        RECT 65.160 106.870 65.300 112.330 ;
        RECT 65.100 106.550 65.360 106.870 ;
        RECT 64.640 106.210 64.900 106.530 ;
        RECT 64.700 105.510 64.840 106.210 ;
        RECT 64.640 105.190 64.900 105.510 ;
        RECT 64.700 101.770 64.840 105.190 ;
        RECT 65.100 104.740 65.360 104.830 ;
        RECT 65.620 104.740 65.760 114.970 ;
        RECT 66.020 114.370 66.280 114.690 ;
        RECT 66.080 112.650 66.220 114.370 ;
        RECT 66.020 112.330 66.280 112.650 ;
        RECT 65.100 104.600 65.760 104.740 ;
        RECT 65.100 104.510 65.360 104.600 ;
        RECT 66.020 104.510 66.280 104.830 ;
        RECT 65.160 102.790 65.300 104.510 ;
        RECT 66.080 102.790 66.220 104.510 ;
        RECT 65.100 102.470 65.360 102.790 ;
        RECT 66.020 102.470 66.280 102.790 ;
        RECT 64.640 101.450 64.900 101.770 ;
        RECT 65.100 100.770 65.360 101.090 ;
        RECT 64.180 99.300 64.440 99.390 ;
        RECT 63.780 99.160 64.440 99.300 ;
        RECT 62.790 97.175 63.070 97.545 ;
        RECT 62.340 92.950 62.600 93.270 ;
        RECT 62.340 90.230 62.600 90.550 ;
        RECT 61.880 88.870 62.140 89.190 ;
        RECT 61.420 85.130 61.680 85.450 ;
        RECT 61.870 84.935 62.150 85.305 ;
        RECT 61.420 84.450 61.680 84.770 ;
        RECT 60.040 83.430 60.300 83.750 ;
        RECT 60.500 83.430 60.760 83.750 ;
        RECT 60.960 83.430 61.220 83.750 ;
        RECT 59.120 83.090 59.380 83.410 ;
        RECT 58.660 82.300 58.920 82.390 ;
        RECT 58.260 82.160 58.920 82.300 ;
        RECT 58.660 82.070 58.920 82.160 ;
        RECT 59.180 81.030 59.320 83.090 ;
        RECT 59.580 82.750 59.840 83.070 ;
        RECT 59.640 82.050 59.780 82.750 ;
        RECT 59.580 81.730 59.840 82.050 ;
        RECT 59.120 80.710 59.380 81.030 ;
        RECT 59.180 78.310 59.320 80.710 ;
        RECT 59.580 80.370 59.840 80.690 ;
        RECT 59.640 78.390 59.780 80.370 ;
        RECT 60.100 79.330 60.240 83.430 ;
        RECT 60.500 82.750 60.760 83.070 ;
        RECT 60.560 81.030 60.700 82.750 ;
        RECT 60.960 82.070 61.220 82.390 ;
        RECT 60.500 80.710 60.760 81.030 ;
        RECT 60.040 79.010 60.300 79.330 ;
        RECT 61.020 78.390 61.160 82.070 ;
        RECT 59.120 77.990 59.380 78.310 ;
        RECT 59.640 78.250 61.160 78.390 ;
        RECT 57.740 77.650 58.000 77.970 ;
        RECT 57.280 77.310 57.540 77.630 ;
        RECT 56.820 68.810 57.080 69.130 ;
        RECT 56.360 65.410 56.620 65.730 ;
        RECT 54.980 64.050 55.240 64.370 ;
        RECT 57.800 63.690 57.940 77.650 ;
        RECT 59.640 77.630 59.780 78.250 ;
        RECT 59.580 77.310 59.840 77.630 ;
        RECT 59.120 76.970 59.380 77.290 ;
        RECT 59.180 64.710 59.320 76.970 ;
        RECT 59.640 74.570 59.780 77.310 ;
        RECT 60.500 76.970 60.760 77.290 ;
        RECT 59.580 74.250 59.840 74.570 ;
        RECT 60.040 74.250 60.300 74.570 ;
        RECT 60.100 72.870 60.240 74.250 ;
        RECT 60.040 72.550 60.300 72.870 ;
        RECT 60.100 70.150 60.240 72.550 ;
        RECT 60.560 72.530 60.700 76.970 ;
        RECT 60.500 72.210 60.760 72.530 ;
        RECT 60.040 69.830 60.300 70.150 ;
        RECT 60.040 68.130 60.300 68.450 ;
        RECT 60.100 66.830 60.240 68.130 ;
        RECT 60.560 67.430 60.700 72.210 ;
        RECT 60.500 67.110 60.760 67.430 ;
        RECT 60.100 66.690 60.700 66.830 ;
        RECT 59.120 64.390 59.380 64.710 ;
        RECT 52.680 63.370 53.340 63.430 ;
        RECT 54.060 63.370 54.320 63.690 ;
        RECT 57.740 63.370 58.000 63.690 ;
        RECT 52.740 63.290 53.340 63.370 ;
        RECT 52.220 62.690 52.480 63.010 ;
        RECT 51.760 60.990 52.020 61.310 ;
        RECT 51.820 56.550 51.960 60.990 ;
        RECT 52.220 59.970 52.480 60.290 ;
        RECT 52.280 58.250 52.420 59.970 ;
        RECT 52.220 57.930 52.480 58.250 ;
        RECT 51.760 56.230 52.020 56.550 ;
        RECT 52.280 54.590 52.420 57.930 ;
        RECT 52.680 54.590 52.940 54.850 ;
        RECT 52.280 54.530 52.940 54.590 ;
        RECT 52.280 54.450 52.880 54.530 ;
        RECT 51.760 52.040 52.020 52.130 ;
        RECT 52.280 52.040 52.420 54.450 ;
        RECT 51.760 51.900 52.420 52.040 ;
        RECT 51.760 51.810 52.020 51.900 ;
        RECT 51.300 48.070 51.560 48.390 ;
        RECT 49.920 44.330 51.040 44.390 ;
        RECT 49.980 44.250 51.040 44.330 ;
        RECT 46.700 43.650 46.960 43.970 ;
        RECT 46.760 41.930 46.900 43.650 ;
        RECT 46.700 41.610 46.960 41.930 ;
        RECT 50.900 40.230 51.040 44.250 ;
        RECT 50.840 39.910 51.100 40.230 ;
        RECT 45.310 38.015 45.590 38.385 ;
        RECT 41.180 37.190 41.440 37.510 ;
        RECT 34.280 35.490 34.540 35.810 ;
        RECT 30.950 34.955 32.490 35.325 ;
        RECT 27.650 32.235 29.190 32.605 ;
        RECT 30.950 29.515 32.490 29.885 ;
        RECT 27.650 26.795 29.190 27.165 ;
        RECT 30.950 24.075 32.490 24.445 ;
        RECT 34.340 23.230 34.480 35.490 ;
        RECT 51.360 32.070 51.500 48.070 ;
        RECT 52.220 46.710 52.480 47.030 ;
        RECT 52.280 42.270 52.420 46.710 ;
        RECT 52.220 41.950 52.480 42.270 ;
        RECT 52.680 34.130 52.940 34.450 ;
        RECT 51.300 31.750 51.560 32.070 ;
        RECT 52.220 31.070 52.480 31.390 ;
        RECT 50.840 30.730 51.100 31.050 ;
        RECT 50.900 29.010 51.040 30.730 ;
        RECT 50.840 28.690 51.100 29.010 ;
        RECT 50.370 27.815 50.650 28.185 ;
        RECT 46.700 27.330 46.960 27.650 ;
        RECT 46.760 25.950 46.900 27.330 ;
        RECT 46.700 25.630 46.960 25.950 ;
        RECT 50.440 25.610 50.580 27.815 ;
        RECT 50.380 25.290 50.640 25.610 ;
        RECT 50.380 24.610 50.640 24.930 ;
        RECT 34.280 22.910 34.540 23.230 ;
        RECT 27.650 21.355 29.190 21.725 ;
        RECT 50.440 20.170 50.580 24.610 ;
        RECT 50.900 20.850 51.040 28.690 ;
        RECT 52.280 28.670 52.420 31.070 ;
        RECT 52.740 30.110 52.880 34.130 ;
        RECT 53.200 31.050 53.340 63.290 ;
        RECT 53.600 34.470 53.860 34.790 ;
        RECT 53.660 31.050 53.800 34.470 ;
        RECT 54.120 34.450 54.260 63.370 ;
        RECT 55.440 60.990 55.700 61.310 ;
        RECT 54.520 55.210 54.780 55.530 ;
        RECT 54.580 50.090 54.720 55.210 ;
        RECT 55.500 51.110 55.640 60.990 ;
        RECT 59.120 60.650 59.380 60.970 ;
        RECT 59.180 58.250 59.320 60.650 ;
        RECT 59.120 57.930 59.380 58.250 ;
        RECT 55.900 55.550 56.160 55.870 ;
        RECT 58.660 55.550 58.920 55.870 ;
        RECT 55.960 52.470 56.100 55.550 ;
        RECT 55.900 52.150 56.160 52.470 ;
        RECT 55.440 50.790 55.700 51.110 ;
        RECT 54.520 49.770 54.780 50.090 ;
        RECT 54.580 45.670 54.720 49.770 ;
        RECT 55.500 49.410 55.640 50.790 ;
        RECT 55.960 50.430 56.100 52.150 ;
        RECT 58.720 51.110 58.860 55.550 ;
        RECT 58.660 50.790 58.920 51.110 ;
        RECT 55.900 50.110 56.160 50.430 ;
        RECT 55.440 49.090 55.700 49.410 ;
        RECT 55.500 48.050 55.640 49.090 ;
        RECT 55.440 47.730 55.700 48.050 ;
        RECT 54.520 45.350 54.780 45.670 ;
        RECT 54.980 44.670 55.240 44.990 ;
        RECT 55.040 39.550 55.180 44.670 ;
        RECT 55.500 39.550 55.640 47.730 ;
        RECT 55.960 47.370 56.100 50.110 ;
        RECT 55.900 47.050 56.160 47.370 ;
        RECT 55.960 45.330 56.100 47.050 ;
        RECT 58.660 46.940 58.920 47.030 ;
        RECT 59.180 46.940 59.320 57.930 ;
        RECT 60.560 54.850 60.700 66.690 ;
        RECT 61.480 62.865 61.620 84.450 ;
        RECT 61.940 83.750 62.080 84.935 ;
        RECT 61.880 83.430 62.140 83.750 ;
        RECT 61.940 83.070 62.080 83.430 ;
        RECT 61.880 82.750 62.140 83.070 ;
        RECT 62.400 80.430 62.540 90.230 ;
        RECT 61.940 80.350 62.540 80.430 ;
        RECT 61.880 80.290 62.540 80.350 ;
        RECT 61.880 80.030 62.140 80.290 ;
        RECT 61.940 79.330 62.080 80.030 ;
        RECT 61.880 79.010 62.140 79.330 ;
        RECT 61.940 78.310 62.080 79.010 ;
        RECT 61.880 77.990 62.140 78.310 ;
        RECT 61.940 74.910 62.080 77.990 ;
        RECT 62.860 77.630 63.000 97.175 ;
        RECT 63.780 95.390 63.920 99.160 ;
        RECT 64.180 99.070 64.440 99.160 ;
        RECT 65.160 96.670 65.300 100.770 ;
        RECT 65.100 96.350 65.360 96.670 ;
        RECT 63.320 95.250 63.920 95.390 ;
        RECT 63.320 91.230 63.460 95.250 ;
        RECT 63.720 94.310 63.980 94.630 ;
        RECT 63.260 90.910 63.520 91.230 ;
        RECT 63.320 87.830 63.460 90.910 ;
        RECT 63.780 88.850 63.920 94.310 ;
        RECT 64.640 93.290 64.900 93.610 ;
        RECT 64.170 91.055 64.450 91.425 ;
        RECT 64.240 89.190 64.380 91.055 ;
        RECT 64.180 88.870 64.440 89.190 ;
        RECT 63.720 88.530 63.980 88.850 ;
        RECT 63.260 87.510 63.520 87.830 ;
        RECT 63.260 84.450 63.520 84.770 ;
        RECT 63.320 80.690 63.460 84.450 ;
        RECT 63.780 83.830 63.920 88.530 ;
        RECT 64.180 87.850 64.440 88.170 ;
        RECT 64.240 84.770 64.380 87.850 ;
        RECT 64.700 85.110 64.840 93.290 ;
        RECT 65.560 92.950 65.820 93.270 ;
        RECT 65.100 91.250 65.360 91.570 ;
        RECT 65.160 87.490 65.300 91.250 ;
        RECT 65.100 87.170 65.360 87.490 ;
        RECT 65.160 86.130 65.300 87.170 ;
        RECT 65.100 85.810 65.360 86.130 ;
        RECT 65.620 85.450 65.760 92.950 ;
        RECT 66.020 89.890 66.280 90.210 ;
        RECT 66.080 88.850 66.220 89.890 ;
        RECT 66.020 88.530 66.280 88.850 ;
        RECT 66.080 85.790 66.220 88.530 ;
        RECT 66.020 85.470 66.280 85.790 ;
        RECT 65.560 85.130 65.820 85.450 ;
        RECT 67.000 85.190 67.140 116.070 ;
        RECT 67.460 112.990 67.600 118.200 ;
        RECT 67.860 117.830 68.120 118.090 ;
        RECT 68.380 117.830 68.520 123.810 ;
        RECT 68.780 123.550 69.040 123.870 ;
        RECT 68.840 120.470 68.980 123.550 ;
        RECT 69.230 122.590 69.510 122.705 ;
        RECT 69.760 122.590 69.900 131.370 ;
        RECT 70.680 131.010 70.820 140.015 ;
        RECT 70.620 130.690 70.880 131.010 ;
        RECT 70.680 127.270 70.820 130.690 ;
        RECT 70.620 126.950 70.880 127.270 ;
        RECT 70.160 126.270 70.420 126.590 ;
        RECT 70.620 126.500 70.880 126.590 ;
        RECT 71.140 126.500 71.280 155.170 ;
        RECT 73.440 154.130 73.580 170.470 ;
        RECT 73.900 156.590 74.040 170.470 ;
        RECT 76.600 170.130 76.860 170.450 ;
        RECT 74.300 169.790 74.560 170.110 ;
        RECT 75.220 169.790 75.480 170.110 ;
        RECT 74.360 159.570 74.500 169.790 ;
        RECT 75.280 168.070 75.420 169.790 ;
        RECT 76.140 169.450 76.400 169.770 ;
        RECT 75.220 167.750 75.480 168.070 ;
        RECT 75.680 167.750 75.940 168.070 ;
        RECT 75.740 167.585 75.880 167.750 ;
        RECT 75.670 167.215 75.950 167.585 ;
        RECT 76.200 167.050 76.340 169.450 ;
        RECT 75.220 166.730 75.480 167.050 ;
        RECT 76.140 166.730 76.400 167.050 ;
        RECT 74.760 166.050 75.020 166.370 ;
        RECT 74.820 165.545 74.960 166.050 ;
        RECT 74.750 165.175 75.030 165.545 ;
        RECT 75.280 165.010 75.420 166.730 ;
        RECT 75.220 164.690 75.480 165.010 ;
        RECT 74.760 164.350 75.020 164.670 ;
        RECT 74.300 159.250 74.560 159.570 ;
        RECT 73.900 156.450 74.500 156.590 ;
        RECT 74.360 155.830 74.500 156.450 ;
        RECT 73.840 155.510 74.100 155.830 ;
        RECT 74.300 155.510 74.560 155.830 ;
        RECT 73.380 153.810 73.640 154.130 ;
        RECT 73.900 153.110 74.040 155.510 ;
        RECT 73.840 152.790 74.100 153.110 ;
        RECT 74.360 152.910 74.500 155.510 ;
        RECT 74.820 155.490 74.960 164.350 ;
        RECT 76.660 161.610 76.800 170.130 ;
        RECT 77.060 168.770 77.320 169.090 ;
        RECT 77.120 164.670 77.260 168.770 ;
        RECT 77.580 165.010 77.720 171.830 ;
        RECT 78.040 170.190 78.180 171.830 ;
        RECT 78.500 170.790 78.640 171.830 ;
        RECT 78.900 171.490 79.160 171.810 ;
        RECT 78.960 170.790 79.100 171.490 ;
        RECT 78.440 170.470 78.700 170.790 ;
        RECT 78.900 170.470 79.160 170.790 ;
        RECT 78.040 170.050 78.640 170.190 ;
        RECT 78.500 169.625 78.640 170.050 ;
        RECT 78.900 169.790 79.160 170.110 ;
        RECT 78.430 169.255 78.710 169.625 ;
        RECT 78.440 168.770 78.700 169.090 ;
        RECT 77.970 167.215 78.250 167.585 ;
        RECT 78.040 165.350 78.180 167.215 ;
        RECT 78.500 166.710 78.640 168.770 ;
        RECT 78.960 166.710 79.100 169.790 ;
        RECT 79.880 169.770 80.020 171.830 ;
        RECT 80.740 171.720 81.000 171.810 ;
        RECT 80.340 171.580 81.000 171.720 ;
        RECT 79.350 169.255 79.630 169.625 ;
        RECT 79.820 169.450 80.080 169.770 ;
        RECT 79.420 167.585 79.560 169.255 ;
        RECT 79.350 167.215 79.630 167.585 ;
        RECT 80.340 166.710 80.480 171.580 ;
        RECT 80.740 171.490 81.000 171.580 ;
        RECT 81.260 170.450 81.400 172.170 ;
        RECT 83.030 171.975 83.310 172.345 ;
        RECT 83.500 172.170 83.760 172.490 ;
        RECT 87.180 172.170 87.440 172.490 ;
        RECT 83.040 171.490 83.300 171.810 ;
        RECT 81.200 170.130 81.460 170.450 ;
        RECT 81.660 169.790 81.920 170.110 ;
        RECT 80.740 169.450 81.000 169.770 ;
        RECT 78.440 166.390 78.700 166.710 ;
        RECT 78.900 166.390 79.160 166.710 ;
        RECT 79.880 166.570 80.480 166.710 ;
        RECT 77.980 165.030 78.240 165.350 ;
        RECT 77.520 164.690 77.780 165.010 ;
        RECT 77.060 164.350 77.320 164.670 ;
        RECT 76.600 161.290 76.860 161.610 ;
        RECT 77.060 158.910 77.320 159.230 ;
        RECT 77.120 158.745 77.260 158.910 ;
        RECT 77.050 158.375 77.330 158.745 ;
        RECT 77.120 158.210 77.260 158.375 ;
        RECT 77.060 157.890 77.320 158.210 ;
        RECT 77.060 156.870 77.320 157.190 ;
        RECT 75.220 155.510 75.480 155.830 ;
        RECT 74.760 155.170 75.020 155.490 ;
        RECT 74.820 154.470 74.960 155.170 ;
        RECT 74.760 154.150 75.020 154.470 ;
        RECT 75.280 153.450 75.420 155.510 ;
        RECT 77.120 154.470 77.260 156.870 ;
        RECT 77.060 154.150 77.320 154.470 ;
        RECT 75.220 153.130 75.480 153.450 ;
        RECT 74.360 152.770 74.960 152.910 ;
        RECT 73.380 151.090 73.640 151.410 ;
        RECT 71.540 150.070 71.800 150.390 ;
        RECT 71.600 149.030 71.740 150.070 ;
        RECT 71.540 148.710 71.800 149.030 ;
        RECT 71.540 148.030 71.800 148.350 ;
        RECT 71.600 146.505 71.740 148.030 ;
        RECT 72.000 147.690 72.260 148.010 ;
        RECT 71.530 146.135 71.810 146.505 ;
        RECT 71.540 144.970 71.800 145.290 ;
        RECT 71.600 134.410 71.740 144.970 ;
        RECT 71.540 134.090 71.800 134.410 ;
        RECT 71.600 132.710 71.740 134.090 ;
        RECT 71.540 132.390 71.800 132.710 ;
        RECT 71.540 130.690 71.800 131.010 ;
        RECT 71.600 128.630 71.740 130.690 ;
        RECT 71.540 128.310 71.800 128.630 ;
        RECT 72.060 127.270 72.200 147.690 ;
        RECT 72.460 144.290 72.720 144.610 ;
        RECT 72.520 139.850 72.660 144.290 ;
        RECT 72.920 142.930 73.180 143.250 ;
        RECT 72.460 139.530 72.720 139.850 ;
        RECT 72.980 137.470 73.120 142.930 ;
        RECT 73.440 142.910 73.580 151.090 ;
        RECT 74.300 147.010 74.560 147.330 ;
        RECT 73.840 145.310 74.100 145.630 ;
        RECT 73.380 142.590 73.640 142.910 ;
        RECT 73.900 142.820 74.040 145.310 ;
        RECT 74.360 145.290 74.500 147.010 ;
        RECT 74.300 144.970 74.560 145.290 ;
        RECT 73.900 142.680 74.500 142.820 ;
        RECT 73.830 142.055 74.110 142.425 ;
        RECT 73.900 141.890 74.040 142.055 ;
        RECT 73.840 141.570 74.100 141.890 ;
        RECT 73.900 139.170 74.040 141.570 ;
        RECT 73.380 138.850 73.640 139.170 ;
        RECT 73.840 138.850 74.100 139.170 ;
        RECT 73.440 137.810 73.580 138.850 ;
        RECT 73.380 137.490 73.640 137.810 ;
        RECT 73.900 137.470 74.040 138.850 ;
        RECT 72.920 137.150 73.180 137.470 ;
        RECT 73.840 137.150 74.100 137.470 ;
        RECT 72.460 129.670 72.720 129.990 ;
        RECT 71.540 126.950 71.800 127.270 ;
        RECT 72.000 126.950 72.260 127.270 ;
        RECT 70.620 126.360 71.280 126.500 ;
        RECT 70.620 126.270 70.880 126.360 ;
        RECT 70.220 123.190 70.360 126.270 ;
        RECT 70.680 126.105 70.820 126.270 ;
        RECT 70.610 125.735 70.890 126.105 ;
        RECT 71.600 125.310 71.740 126.950 ;
        RECT 72.000 126.270 72.260 126.590 ;
        RECT 71.140 125.170 71.740 125.310 ;
        RECT 70.620 123.210 70.880 123.530 ;
        RECT 70.160 122.870 70.420 123.190 ;
        RECT 69.230 122.450 69.900 122.590 ;
        RECT 69.230 122.335 69.510 122.450 ;
        RECT 68.780 120.150 69.040 120.470 ;
        RECT 68.770 118.935 69.050 119.305 ;
        RECT 68.840 118.430 68.980 118.935 ;
        RECT 68.780 118.110 69.040 118.430 ;
        RECT 67.860 117.770 68.520 117.830 ;
        RECT 67.920 117.690 68.520 117.770 ;
        RECT 67.920 116.050 68.060 117.690 ;
        RECT 69.300 117.320 69.440 122.335 ;
        RECT 68.380 117.180 69.440 117.320 ;
        RECT 68.380 116.390 68.520 117.180 ;
        RECT 68.320 116.070 68.580 116.390 ;
        RECT 67.860 115.730 68.120 116.050 ;
        RECT 68.320 115.440 68.580 115.760 ;
        RECT 68.380 114.430 68.520 115.440 ;
        RECT 69.700 115.390 69.960 115.710 ;
        RECT 67.920 114.290 68.520 114.430 ;
        RECT 67.400 112.670 67.660 112.990 ;
        RECT 67.460 110.610 67.600 112.670 ;
        RECT 67.920 112.650 68.060 114.290 ;
        RECT 68.310 113.495 68.590 113.865 ;
        RECT 69.760 113.670 69.900 115.390 ;
        RECT 68.320 113.350 68.580 113.495 ;
        RECT 69.700 113.350 69.960 113.670 ;
        RECT 67.860 112.560 68.120 112.650 ;
        RECT 67.860 112.420 68.520 112.560 ;
        RECT 67.860 112.330 68.120 112.420 ;
        RECT 67.400 110.290 67.660 110.610 ;
        RECT 67.400 109.610 67.660 109.930 ;
        RECT 67.460 105.025 67.600 109.610 ;
        RECT 68.380 108.230 68.520 112.420 ;
        RECT 69.700 112.330 69.960 112.650 ;
        RECT 68.780 111.650 69.040 111.970 ;
        RECT 68.320 107.910 68.580 108.230 ;
        RECT 67.860 107.570 68.120 107.890 ;
        RECT 67.390 104.655 67.670 105.025 ;
        RECT 67.920 104.830 68.060 107.570 ;
        RECT 68.320 104.850 68.580 105.170 ;
        RECT 67.400 104.510 67.660 104.655 ;
        RECT 67.860 104.510 68.120 104.830 ;
        RECT 67.860 101.450 68.120 101.770 ;
        RECT 67.920 99.730 68.060 101.450 ;
        RECT 67.860 99.410 68.120 99.730 ;
        RECT 67.400 99.070 67.660 99.390 ;
        RECT 67.460 97.350 67.600 99.070 ;
        RECT 68.380 97.350 68.520 104.850 ;
        RECT 67.400 97.030 67.660 97.350 ;
        RECT 68.320 97.030 68.580 97.350 ;
        RECT 67.860 93.630 68.120 93.950 ;
        RECT 67.920 92.840 68.060 93.630 ;
        RECT 68.380 93.610 68.520 97.030 ;
        RECT 68.320 93.290 68.580 93.610 ;
        RECT 67.920 92.700 68.520 92.840 ;
        RECT 67.860 88.190 68.120 88.510 ;
        RECT 67.920 85.985 68.060 88.190 ;
        RECT 67.850 85.615 68.130 85.985 ;
        RECT 68.380 85.450 68.520 92.700 ;
        RECT 68.840 90.890 68.980 111.650 ;
        RECT 69.240 103.490 69.500 103.810 ;
        RECT 69.300 101.770 69.440 103.490 ;
        RECT 69.760 102.790 69.900 112.330 ;
        RECT 70.220 104.830 70.360 122.870 ;
        RECT 70.680 113.330 70.820 123.210 ;
        RECT 70.620 113.010 70.880 113.330 ;
        RECT 71.140 112.650 71.280 125.170 ;
        RECT 71.540 123.550 71.800 123.870 ;
        RECT 71.600 121.150 71.740 123.550 ;
        RECT 71.540 120.830 71.800 121.150 ;
        RECT 71.540 118.450 71.800 118.770 ;
        RECT 71.600 117.945 71.740 118.450 ;
        RECT 71.530 117.575 71.810 117.945 ;
        RECT 71.540 113.010 71.800 113.330 ;
        RECT 71.080 112.330 71.340 112.650 ;
        RECT 71.080 111.650 71.340 111.970 ;
        RECT 71.140 110.270 71.280 111.650 ;
        RECT 71.080 109.950 71.340 110.270 ;
        RECT 71.080 107.570 71.340 107.890 ;
        RECT 70.160 104.510 70.420 104.830 ;
        RECT 69.700 102.470 69.960 102.790 ;
        RECT 69.240 101.450 69.500 101.770 ;
        RECT 71.140 95.990 71.280 107.570 ;
        RECT 71.080 95.670 71.340 95.990 ;
        RECT 71.140 93.950 71.280 95.670 ;
        RECT 71.080 93.630 71.340 93.950 ;
        RECT 71.600 93.350 71.740 113.010 ;
        RECT 72.060 107.890 72.200 126.270 ;
        RECT 72.520 126.250 72.660 129.670 ;
        RECT 72.460 125.930 72.720 126.250 ;
        RECT 72.460 122.530 72.720 122.850 ;
        RECT 72.520 112.990 72.660 122.530 ;
        RECT 72.980 117.750 73.120 137.150 ;
        RECT 73.380 133.410 73.640 133.730 ;
        RECT 74.360 133.470 74.500 142.680 ;
        RECT 74.820 140.190 74.960 152.770 ;
        RECT 75.220 152.450 75.480 152.770 ;
        RECT 75.280 149.030 75.420 152.450 ;
        RECT 75.220 148.710 75.480 149.030 ;
        RECT 74.760 139.870 75.020 140.190 ;
        RECT 73.440 132.710 73.580 133.410 ;
        RECT 73.900 133.330 74.500 133.470 ;
        RECT 73.380 132.390 73.640 132.710 ;
        RECT 73.900 124.550 74.040 133.330 ;
        RECT 74.300 132.390 74.560 132.710 ;
        RECT 73.840 124.230 74.100 124.550 ;
        RECT 73.840 123.550 74.100 123.870 ;
        RECT 73.380 122.530 73.640 122.850 ;
        RECT 73.440 118.090 73.580 122.530 ;
        RECT 73.900 119.110 74.040 123.550 ;
        RECT 73.840 118.790 74.100 119.110 ;
        RECT 74.360 118.410 74.500 132.390 ;
        RECT 74.820 129.650 74.960 139.870 ;
        RECT 75.680 139.705 75.940 139.850 ;
        RECT 75.670 139.335 75.950 139.705 ;
        RECT 76.140 139.190 76.400 139.510 ;
        RECT 76.200 136.450 76.340 139.190 ;
        RECT 76.140 136.130 76.400 136.450 ;
        RECT 75.680 134.430 75.940 134.750 ;
        RECT 75.220 131.710 75.480 132.030 ;
        RECT 74.760 129.330 75.020 129.650 ;
        RECT 74.820 128.970 74.960 129.330 ;
        RECT 74.760 128.650 75.020 128.970 ;
        RECT 74.760 124.230 75.020 124.550 ;
        RECT 74.820 119.110 74.960 124.230 ;
        RECT 74.760 118.790 75.020 119.110 ;
        RECT 74.360 118.270 74.960 118.410 ;
        RECT 73.380 117.770 73.640 118.090 ;
        RECT 72.920 117.430 73.180 117.750 ;
        RECT 72.920 114.370 73.180 114.690 ;
        RECT 72.980 112.990 73.120 114.370 ;
        RECT 72.460 112.670 72.720 112.990 ;
        RECT 72.920 112.670 73.180 112.990 ;
        RECT 72.460 110.290 72.720 110.610 ;
        RECT 72.000 107.570 72.260 107.890 ;
        RECT 72.000 106.210 72.260 106.530 ;
        RECT 72.060 104.490 72.200 106.210 ;
        RECT 72.520 105.170 72.660 110.290 ;
        RECT 74.300 106.550 74.560 106.870 ;
        RECT 72.460 104.850 72.720 105.170 ;
        RECT 72.000 104.170 72.260 104.490 ;
        RECT 72.920 100.770 73.180 101.090 ;
        RECT 71.990 99.895 72.270 100.265 ;
        RECT 72.060 94.630 72.200 99.895 ;
        RECT 72.000 94.310 72.260 94.630 ;
        RECT 72.980 93.950 73.120 100.770 ;
        RECT 73.380 98.050 73.640 98.370 ;
        RECT 73.440 96.330 73.580 98.050 ;
        RECT 73.380 96.010 73.640 96.330 ;
        RECT 72.920 93.630 73.180 93.950 ;
        RECT 70.220 93.210 71.740 93.350 ;
        RECT 69.700 92.610 69.960 92.930 ;
        RECT 68.780 90.570 69.040 90.890 ;
        RECT 64.640 84.790 64.900 85.110 ;
        RECT 64.180 84.450 64.440 84.770 ;
        RECT 63.780 83.690 64.380 83.830 ;
        RECT 63.720 83.090 63.980 83.410 ;
        RECT 63.260 80.370 63.520 80.690 ;
        RECT 63.780 80.010 63.920 83.090 ;
        RECT 63.720 79.690 63.980 80.010 ;
        RECT 62.800 77.310 63.060 77.630 ;
        RECT 64.240 75.250 64.380 83.690 ;
        RECT 64.700 83.150 64.840 84.790 ;
        RECT 65.620 83.750 65.760 85.130 ;
        RECT 66.540 85.050 67.140 85.190 ;
        RECT 68.320 85.130 68.580 85.450 ;
        RECT 68.840 85.360 68.980 90.570 ;
        RECT 69.240 89.890 69.500 90.210 ;
        RECT 69.300 88.170 69.440 89.890 ;
        RECT 69.240 87.850 69.500 88.170 ;
        RECT 69.240 85.360 69.500 85.450 ;
        RECT 68.840 85.220 69.500 85.360 ;
        RECT 69.240 85.130 69.500 85.220 ;
        RECT 65.560 83.430 65.820 83.750 ;
        RECT 64.700 83.070 65.300 83.150 ;
        RECT 64.700 83.010 65.360 83.070 ;
        RECT 65.100 82.750 65.360 83.010 ;
        RECT 65.550 82.895 65.830 83.265 ;
        RECT 65.560 82.750 65.820 82.895 ;
        RECT 64.640 82.410 64.900 82.730 ;
        RECT 64.700 80.010 64.840 82.410 ;
        RECT 65.160 80.350 65.300 82.750 ;
        RECT 66.540 80.430 66.680 85.050 ;
        RECT 66.940 84.450 67.200 84.770 ;
        RECT 67.000 82.730 67.140 84.450 ;
        RECT 68.380 83.070 68.520 85.130 ;
        RECT 69.760 84.770 69.900 92.610 ;
        RECT 69.240 84.625 69.500 84.770 ;
        RECT 69.230 84.255 69.510 84.625 ;
        RECT 69.700 84.450 69.960 84.770 ;
        RECT 68.320 82.750 68.580 83.070 ;
        RECT 66.940 82.410 67.200 82.730 ;
        RECT 68.780 82.070 69.040 82.390 ;
        RECT 67.400 81.730 67.660 82.050 ;
        RECT 68.320 81.730 68.580 82.050 ;
        RECT 65.100 80.030 65.360 80.350 ;
        RECT 66.540 80.290 67.140 80.430 ;
        RECT 64.640 79.865 64.900 80.010 ;
        RECT 64.630 79.495 64.910 79.865 ;
        RECT 66.020 79.750 66.280 80.010 ;
        RECT 66.020 79.690 66.680 79.750 ;
        RECT 66.080 79.610 66.680 79.690 ;
        RECT 64.180 74.930 64.440 75.250 ;
        RECT 61.880 74.590 62.140 74.910 ;
        RECT 66.540 74.570 66.680 79.610 ;
        RECT 67.000 77.630 67.140 80.290 ;
        RECT 67.460 79.670 67.600 81.730 ;
        RECT 67.400 79.350 67.660 79.670 ;
        RECT 66.940 77.310 67.200 77.630 ;
        RECT 66.480 74.250 66.740 74.570 ;
        RECT 65.560 73.570 65.820 73.890 ;
        RECT 64.180 70.850 64.440 71.170 ;
        RECT 63.720 68.810 63.980 69.130 ;
        RECT 63.780 66.750 63.920 68.810 ;
        RECT 64.240 67.090 64.380 70.850 ;
        RECT 65.620 69.470 65.760 73.570 ;
        RECT 66.540 69.470 66.680 74.250 ;
        RECT 67.000 72.530 67.140 77.310 ;
        RECT 67.400 76.290 67.660 76.610 ;
        RECT 67.860 76.290 68.120 76.610 ;
        RECT 67.460 72.870 67.600 76.290 ;
        RECT 67.920 74.570 68.060 76.290 ;
        RECT 67.860 74.250 68.120 74.570 ;
        RECT 67.400 72.550 67.660 72.870 ;
        RECT 66.940 72.210 67.200 72.530 ;
        RECT 67.000 71.850 67.140 72.210 ;
        RECT 68.380 72.190 68.520 81.730 ;
        RECT 68.840 77.290 68.980 82.070 ;
        RECT 68.780 76.970 69.040 77.290 ;
        RECT 68.320 71.870 68.580 72.190 ;
        RECT 69.760 71.850 69.900 84.450 ;
        RECT 66.940 71.530 67.200 71.850 ;
        RECT 69.700 71.530 69.960 71.850 ;
        RECT 68.320 71.190 68.580 71.510 ;
        RECT 67.860 70.850 68.120 71.170 ;
        RECT 65.560 69.150 65.820 69.470 ;
        RECT 66.480 69.150 66.740 69.470 ;
        RECT 66.020 68.810 66.280 69.130 ;
        RECT 65.100 68.130 65.360 68.450 ;
        RECT 64.180 66.770 64.440 67.090 ;
        RECT 63.720 66.430 63.980 66.750 ;
        RECT 65.160 63.690 65.300 68.130 ;
        RECT 66.080 67.430 66.220 68.810 ;
        RECT 67.920 68.790 68.060 70.850 ;
        RECT 67.860 68.470 68.120 68.790 ;
        RECT 67.850 67.935 68.130 68.305 ;
        RECT 66.020 67.110 66.280 67.430 ;
        RECT 66.940 66.430 67.200 66.750 ;
        RECT 65.100 63.370 65.360 63.690 ;
        RECT 61.410 62.495 61.690 62.865 ;
        RECT 61.420 59.970 61.680 60.290 ;
        RECT 60.500 54.530 60.760 54.850 ;
        RECT 60.560 51.110 60.700 54.530 ;
        RECT 60.500 50.790 60.760 51.110 ;
        RECT 61.480 50.090 61.620 59.970 ;
        RECT 63.720 57.590 63.980 57.910 ;
        RECT 64.180 57.590 64.440 57.910 ;
        RECT 63.780 53.830 63.920 57.590 ;
        RECT 64.240 55.870 64.380 57.590 ;
        RECT 64.180 55.550 64.440 55.870 ;
        RECT 63.720 53.510 63.980 53.830 ;
        RECT 65.160 52.810 65.300 63.370 ;
        RECT 67.000 63.350 67.140 66.430 ;
        RECT 66.940 63.030 67.200 63.350 ;
        RECT 67.000 61.310 67.140 63.030 ;
        RECT 66.940 60.990 67.200 61.310 ;
        RECT 67.000 57.910 67.140 60.990 ;
        RECT 66.940 57.590 67.200 57.910 ;
        RECT 66.930 55.695 67.210 56.065 ;
        RECT 66.480 52.830 66.740 53.150 ;
        RECT 65.100 52.490 65.360 52.810 ;
        RECT 62.340 51.810 62.600 52.130 ;
        RECT 66.020 51.810 66.280 52.130 ;
        RECT 61.420 49.770 61.680 50.090 ;
        RECT 60.040 49.090 60.300 49.410 ;
        RECT 58.660 46.800 59.320 46.940 ;
        RECT 58.660 46.710 58.920 46.800 ;
        RECT 59.580 46.710 59.840 47.030 ;
        RECT 56.360 46.370 56.620 46.690 ;
        RECT 55.900 45.010 56.160 45.330 ;
        RECT 54.980 39.230 55.240 39.550 ;
        RECT 55.440 39.230 55.700 39.550 ;
        RECT 54.060 34.130 54.320 34.450 ;
        RECT 54.060 33.110 54.320 33.430 ;
        RECT 54.120 31.050 54.260 33.110 ;
        RECT 55.960 31.050 56.100 45.010 ;
        RECT 56.420 39.550 56.560 46.370 ;
        RECT 58.720 43.970 58.860 46.710 ;
        RECT 58.660 43.650 58.920 43.970 ;
        RECT 56.820 40.930 57.080 41.250 ;
        RECT 56.360 39.230 56.620 39.550 ;
        RECT 56.880 39.210 57.020 40.930 ;
        RECT 56.820 38.890 57.080 39.210 ;
        RECT 56.360 38.210 56.620 38.530 ;
        RECT 56.420 36.490 56.560 38.210 ;
        RECT 59.640 37.510 59.780 46.710 ;
        RECT 60.100 41.930 60.240 49.090 ;
        RECT 60.500 43.650 60.760 43.970 ;
        RECT 60.560 41.930 60.700 43.650 ;
        RECT 60.040 41.610 60.300 41.930 ;
        RECT 60.500 41.610 60.760 41.930 ;
        RECT 61.480 40.230 61.620 49.770 ;
        RECT 61.880 48.070 62.140 48.390 ;
        RECT 61.940 42.270 62.080 48.070 ;
        RECT 62.400 44.990 62.540 51.810 ;
        RECT 66.080 50.430 66.220 51.810 ;
        RECT 66.020 50.110 66.280 50.430 ;
        RECT 62.800 49.090 63.060 49.410 ;
        RECT 65.560 49.090 65.820 49.410 ;
        RECT 62.860 47.370 63.000 49.090 ;
        RECT 65.100 48.070 65.360 48.390 ;
        RECT 62.800 47.050 63.060 47.370 ;
        RECT 63.260 45.350 63.520 45.670 ;
        RECT 62.340 44.670 62.600 44.990 ;
        RECT 61.880 41.950 62.140 42.270 ;
        RECT 62.400 41.590 62.540 44.670 ;
        RECT 63.320 42.950 63.460 45.350 ;
        RECT 64.640 44.670 64.900 44.990 ;
        RECT 64.700 42.950 64.840 44.670 ;
        RECT 63.260 42.860 63.520 42.950 ;
        RECT 62.860 42.720 63.520 42.860 ;
        RECT 62.340 41.270 62.600 41.590 ;
        RECT 62.860 40.230 63.000 42.720 ;
        RECT 63.260 42.630 63.520 42.720 ;
        RECT 64.640 42.630 64.900 42.950 ;
        RECT 61.420 39.910 61.680 40.230 ;
        RECT 62.800 39.910 63.060 40.230 ;
        RECT 62.340 39.230 62.600 39.550 ;
        RECT 61.880 38.890 62.140 39.210 ;
        RECT 60.960 38.210 61.220 38.530 ;
        RECT 59.580 37.190 59.840 37.510 ;
        RECT 61.020 36.490 61.160 38.210 ;
        RECT 56.360 36.170 56.620 36.490 ;
        RECT 60.500 36.170 60.760 36.490 ;
        RECT 60.960 36.170 61.220 36.490 ;
        RECT 60.560 34.790 60.700 36.170 ;
        RECT 60.500 34.470 60.760 34.790 ;
        RECT 61.020 34.110 61.160 36.170 ;
        RECT 61.420 35.490 61.680 35.810 ;
        RECT 60.960 33.790 61.220 34.110 ;
        RECT 53.140 30.730 53.400 31.050 ;
        RECT 53.600 30.730 53.860 31.050 ;
        RECT 54.060 30.730 54.320 31.050 ;
        RECT 55.900 30.730 56.160 31.050 ;
        RECT 52.740 29.970 53.340 30.110 ;
        RECT 53.200 29.010 53.340 29.970 ;
        RECT 53.140 28.690 53.400 29.010 ;
        RECT 52.220 28.350 52.480 28.670 ;
        RECT 51.300 27.330 51.560 27.650 ;
        RECT 51.360 23.570 51.500 27.330 ;
        RECT 52.280 25.270 52.420 28.350 ;
        RECT 52.680 25.290 52.940 25.610 ;
        RECT 52.220 24.950 52.480 25.270 ;
        RECT 52.740 23.910 52.880 25.290 ;
        RECT 52.680 23.590 52.940 23.910 ;
        RECT 51.300 23.250 51.560 23.570 ;
        RECT 50.840 20.530 51.100 20.850 ;
        RECT 52.740 20.170 52.880 23.590 ;
        RECT 53.200 20.510 53.340 28.690 ;
        RECT 53.660 28.330 53.800 30.730 ;
        RECT 54.520 30.050 54.780 30.370 ;
        RECT 54.580 28.670 54.720 30.050 ;
        RECT 55.440 28.690 55.700 29.010 ;
        RECT 54.520 28.350 54.780 28.670 ;
        RECT 53.600 28.010 53.860 28.330 ;
        RECT 55.500 26.630 55.640 28.690 ;
        RECT 55.960 28.330 56.100 30.730 ;
        RECT 60.500 30.050 60.760 30.370 ;
        RECT 58.660 28.350 58.920 28.670 ;
        RECT 55.900 28.010 56.160 28.330 ;
        RECT 55.440 26.310 55.700 26.630 ;
        RECT 55.960 25.950 56.100 28.010 ;
        RECT 55.900 25.630 56.160 25.950 ;
        RECT 58.720 23.910 58.860 28.350 ;
        RECT 60.560 26.030 60.700 30.050 ;
        RECT 61.020 27.650 61.160 33.790 ;
        RECT 61.480 29.350 61.620 35.490 ;
        RECT 61.940 34.450 62.080 38.890 ;
        RECT 61.880 34.130 62.140 34.450 ;
        RECT 62.400 33.090 62.540 39.230 ;
        RECT 62.860 39.210 63.000 39.910 ;
        RECT 62.800 38.890 63.060 39.210 ;
        RECT 65.160 38.530 65.300 48.070 ;
        RECT 65.620 47.370 65.760 49.090 ;
        RECT 65.560 47.050 65.820 47.370 ;
        RECT 66.080 41.250 66.220 50.110 ;
        RECT 66.020 40.930 66.280 41.250 ;
        RECT 65.100 38.210 65.360 38.530 ;
        RECT 62.790 36.655 63.070 37.025 ;
        RECT 62.340 32.770 62.600 33.090 ;
        RECT 62.400 32.070 62.540 32.770 ;
        RECT 62.340 31.750 62.600 32.070 ;
        RECT 61.420 29.030 61.680 29.350 ;
        RECT 60.960 27.330 61.220 27.650 ;
        RECT 61.020 26.630 61.160 27.330 ;
        RECT 60.960 26.310 61.220 26.630 ;
        RECT 60.560 25.890 61.160 26.030 ;
        RECT 58.660 23.590 58.920 23.910 ;
        RECT 61.020 22.890 61.160 25.890 ;
        RECT 61.480 22.890 61.620 29.030 ;
        RECT 62.400 25.270 62.540 31.750 ;
        RECT 62.860 27.990 63.000 36.655 ;
        RECT 65.160 36.490 65.300 38.210 ;
        RECT 66.080 36.910 66.220 40.930 ;
        RECT 66.540 40.230 66.680 52.830 ;
        RECT 66.480 39.910 66.740 40.230 ;
        RECT 67.000 37.510 67.140 55.695 ;
        RECT 67.920 54.850 68.060 67.935 ;
        RECT 68.380 67.090 68.520 71.190 ;
        RECT 68.320 66.770 68.580 67.090 ;
        RECT 69.760 64.790 69.900 71.530 ;
        RECT 70.220 68.985 70.360 93.210 ;
        RECT 71.540 91.590 71.800 91.910 ;
        RECT 71.080 89.890 71.340 90.210 ;
        RECT 71.140 85.110 71.280 89.890 ;
        RECT 71.080 84.790 71.340 85.110 ;
        RECT 71.140 79.670 71.280 84.790 ;
        RECT 71.600 84.770 71.740 91.590 ;
        RECT 72.000 90.570 72.260 90.890 ;
        RECT 72.920 90.570 73.180 90.890 ;
        RECT 73.840 90.570 74.100 90.890 ;
        RECT 72.060 87.910 72.200 90.570 ;
        RECT 72.980 89.385 73.120 90.570 ;
        RECT 73.380 89.890 73.640 90.210 ;
        RECT 72.910 89.015 73.190 89.385 ;
        RECT 72.920 88.190 73.180 88.510 ;
        RECT 72.060 87.770 72.660 87.910 ;
        RECT 72.520 87.490 72.660 87.770 ;
        RECT 72.460 87.170 72.720 87.490 ;
        RECT 72.980 85.110 73.120 88.190 ;
        RECT 73.440 85.110 73.580 89.890 ;
        RECT 73.900 88.850 74.040 90.570 ;
        RECT 73.840 88.530 74.100 88.850 ;
        RECT 73.840 87.850 74.100 88.170 ;
        RECT 72.920 84.790 73.180 85.110 ;
        RECT 73.380 84.790 73.640 85.110 ;
        RECT 71.540 84.450 71.800 84.770 ;
        RECT 71.080 79.350 71.340 79.670 ;
        RECT 70.620 79.010 70.880 79.330 ;
        RECT 70.680 78.310 70.820 79.010 ;
        RECT 70.620 77.990 70.880 78.310 ;
        RECT 71.600 75.590 71.740 84.450 ;
        RECT 72.920 82.410 73.180 82.730 ;
        RECT 72.980 79.330 73.120 82.410 ;
        RECT 73.440 80.350 73.580 84.790 ;
        RECT 73.380 80.030 73.640 80.350 ;
        RECT 72.920 79.010 73.180 79.330 ;
        RECT 73.380 79.240 73.640 79.330 ;
        RECT 73.900 79.240 74.040 87.850 ;
        RECT 73.380 79.100 74.040 79.240 ;
        RECT 73.380 79.010 73.640 79.100 ;
        RECT 72.980 77.970 73.120 79.010 ;
        RECT 72.920 77.650 73.180 77.970 ;
        RECT 71.540 75.270 71.800 75.590 ;
        RECT 70.150 68.615 70.430 68.985 ;
        RECT 69.760 64.650 70.820 64.790 ;
        RECT 70.160 62.690 70.420 63.010 ;
        RECT 68.780 57.250 69.040 57.570 ;
        RECT 68.840 56.210 68.980 57.250 ;
        RECT 68.780 55.890 69.040 56.210 ;
        RECT 67.860 54.530 68.120 54.850 ;
        RECT 67.860 53.170 68.120 53.490 ;
        RECT 67.400 52.830 67.660 53.150 ;
        RECT 67.460 48.390 67.600 52.830 ;
        RECT 67.400 48.070 67.660 48.390 ;
        RECT 67.400 46.710 67.660 47.030 ;
        RECT 67.460 42.270 67.600 46.710 ;
        RECT 67.400 41.950 67.660 42.270 ;
        RECT 66.940 37.190 67.200 37.510 ;
        RECT 66.080 36.770 67.140 36.910 ;
        RECT 65.100 36.170 65.360 36.490 ;
        RECT 64.180 35.490 64.440 35.810 ;
        RECT 63.720 30.730 63.980 31.050 ;
        RECT 62.800 27.670 63.060 27.990 ;
        RECT 62.340 24.950 62.600 25.270 ;
        RECT 62.860 23.910 63.000 27.670 ;
        RECT 63.780 25.950 63.920 30.730 ;
        RECT 63.720 25.630 63.980 25.950 ;
        RECT 64.240 25.270 64.380 35.490 ;
        RECT 65.160 34.110 65.300 36.170 ;
        RECT 66.470 34.615 66.750 34.985 ;
        RECT 66.480 34.470 66.740 34.615 ;
        RECT 65.100 33.790 65.360 34.110 ;
        RECT 67.000 33.770 67.140 36.770 ;
        RECT 67.920 36.490 68.060 53.170 ;
        RECT 68.840 52.470 68.980 55.890 ;
        RECT 69.700 55.550 69.960 55.870 ;
        RECT 68.780 52.150 69.040 52.470 ;
        RECT 69.240 52.150 69.500 52.470 ;
        RECT 68.320 51.810 68.580 52.130 ;
        RECT 68.380 50.090 68.520 51.810 ;
        RECT 68.320 49.770 68.580 50.090 ;
        RECT 69.300 47.710 69.440 52.150 ;
        RECT 69.760 51.110 69.900 55.550 ;
        RECT 69.700 50.790 69.960 51.110 ;
        RECT 70.220 50.510 70.360 62.690 ;
        RECT 70.680 50.770 70.820 64.650 ;
        RECT 72.920 64.620 73.180 64.710 ;
        RECT 73.440 64.620 73.580 79.010 ;
        RECT 74.360 71.510 74.500 106.550 ;
        RECT 74.820 96.330 74.960 118.270 ;
        RECT 75.280 113.670 75.420 131.710 ;
        RECT 75.740 129.310 75.880 134.430 ;
        RECT 77.120 134.410 77.260 154.150 ;
        RECT 77.580 136.450 77.720 164.690 ;
        RECT 79.360 161.970 79.620 162.290 ;
        RECT 78.440 161.290 78.700 161.610 ;
        RECT 77.980 160.950 78.240 161.270 ;
        RECT 78.040 159.230 78.180 160.950 ;
        RECT 77.980 158.910 78.240 159.230 ;
        RECT 78.040 155.910 78.180 158.910 ;
        RECT 78.500 156.510 78.640 161.290 ;
        RECT 79.420 159.230 79.560 161.970 ;
        RECT 79.880 161.610 80.020 166.570 ;
        RECT 80.800 162.030 80.940 169.450 ;
        RECT 81.190 169.255 81.470 169.625 ;
        RECT 81.260 169.090 81.400 169.255 ;
        RECT 81.200 168.770 81.460 169.090 ;
        RECT 81.200 166.730 81.460 167.050 ;
        RECT 80.340 161.890 80.940 162.030 ;
        RECT 79.820 161.290 80.080 161.610 ;
        RECT 79.360 158.910 79.620 159.230 ;
        RECT 78.900 158.570 79.160 158.890 ;
        RECT 78.440 156.190 78.700 156.510 ;
        RECT 78.040 155.770 78.640 155.910 ;
        RECT 77.980 155.170 78.240 155.490 ;
        RECT 78.040 150.730 78.180 155.170 ;
        RECT 78.500 150.730 78.640 155.770 ;
        RECT 78.960 153.790 79.100 158.570 ;
        RECT 79.420 155.490 79.560 158.910 ;
        RECT 79.360 155.170 79.620 155.490 ;
        RECT 78.900 153.470 79.160 153.790 ;
        RECT 78.960 151.750 79.100 153.470 ;
        RECT 79.420 153.190 79.560 155.170 ;
        RECT 79.820 154.150 80.080 154.470 ;
        RECT 79.880 153.790 80.020 154.150 ;
        RECT 79.820 153.470 80.080 153.790 ;
        RECT 79.420 153.050 80.020 153.190 ;
        RECT 79.360 152.450 79.620 152.770 ;
        RECT 78.900 151.430 79.160 151.750 ;
        RECT 79.420 151.410 79.560 152.450 ;
        RECT 79.360 151.090 79.620 151.410 ;
        RECT 79.880 151.070 80.020 153.050 ;
        RECT 79.820 150.750 80.080 151.070 ;
        RECT 77.980 150.410 78.240 150.730 ;
        RECT 78.440 150.410 78.700 150.730 ;
        RECT 80.340 150.470 80.480 161.890 ;
        RECT 81.260 161.610 81.400 166.730 ;
        RECT 81.200 161.290 81.460 161.610 ;
        RECT 80.740 160.950 81.000 161.270 ;
        RECT 80.800 157.190 80.940 160.950 ;
        RECT 81.260 159.230 81.400 161.290 ;
        RECT 81.720 159.230 81.860 169.790 ;
        RECT 82.120 169.110 82.380 169.430 ;
        RECT 82.180 167.050 82.320 169.110 ;
        RECT 82.120 166.730 82.380 167.050 ;
        RECT 82.580 166.730 82.840 167.050 ;
        RECT 81.200 158.910 81.460 159.230 ;
        RECT 81.660 158.910 81.920 159.230 ;
        RECT 80.740 156.870 81.000 157.190 ;
        RECT 80.740 155.850 81.000 156.170 ;
        RECT 80.800 153.110 80.940 155.850 ;
        RECT 80.740 152.790 81.000 153.110 ;
        RECT 81.260 151.070 81.400 158.910 ;
        RECT 81.660 153.470 81.920 153.790 ;
        RECT 81.720 153.305 81.860 153.470 ;
        RECT 81.650 152.935 81.930 153.305 ;
        RECT 80.740 150.750 81.000 151.070 ;
        RECT 81.200 150.750 81.460 151.070 ;
        RECT 77.980 145.990 78.240 146.310 ;
        RECT 77.520 136.130 77.780 136.450 ;
        RECT 76.130 133.895 76.410 134.265 ;
        RECT 77.060 134.090 77.320 134.410 ;
        RECT 76.200 131.350 76.340 133.895 ;
        RECT 76.600 133.750 76.860 134.070 ;
        RECT 76.140 131.030 76.400 131.350 ;
        RECT 76.660 130.070 76.800 133.750 ;
        RECT 77.120 131.350 77.260 134.090 ;
        RECT 78.040 132.030 78.180 145.990 ;
        RECT 78.500 140.440 78.640 150.410 ;
        RECT 79.880 150.330 80.480 150.470 ;
        RECT 79.360 147.010 79.620 147.330 ;
        RECT 79.420 143.590 79.560 147.010 ;
        RECT 79.360 143.270 79.620 143.590 ;
        RECT 79.360 140.440 79.620 140.530 ;
        RECT 78.500 140.300 79.620 140.440 ;
        RECT 79.360 140.210 79.620 140.300 ;
        RECT 78.900 136.810 79.160 137.130 ;
        RECT 78.440 136.470 78.700 136.790 ;
        RECT 78.500 132.030 78.640 136.470 ;
        RECT 78.960 134.750 79.100 136.810 ;
        RECT 78.900 134.430 79.160 134.750 ;
        RECT 79.420 134.150 79.560 140.210 ;
        RECT 78.960 134.010 79.560 134.150 ;
        RECT 77.980 131.710 78.240 132.030 ;
        RECT 78.440 131.710 78.700 132.030 ;
        RECT 77.060 131.030 77.320 131.350 ;
        RECT 76.660 129.930 77.720 130.070 ;
        RECT 78.040 129.990 78.180 131.710 ;
        RECT 78.440 131.030 78.700 131.350 ;
        RECT 76.600 129.330 76.860 129.650 ;
        RECT 75.680 128.990 75.940 129.310 ;
        RECT 76.140 128.990 76.400 129.310 ;
        RECT 75.740 127.270 75.880 128.990 ;
        RECT 75.680 126.950 75.940 127.270 ;
        RECT 75.670 124.375 75.950 124.745 ;
        RECT 75.740 120.470 75.880 124.375 ;
        RECT 76.200 124.210 76.340 128.990 ;
        RECT 76.140 123.890 76.400 124.210 ;
        RECT 76.140 122.870 76.400 123.190 ;
        RECT 76.200 120.810 76.340 122.870 ;
        RECT 76.140 120.490 76.400 120.810 ;
        RECT 75.680 120.150 75.940 120.470 ;
        RECT 75.680 114.370 75.940 114.690 ;
        RECT 75.220 113.350 75.480 113.670 ;
        RECT 75.740 112.650 75.880 114.370 ;
        RECT 75.680 112.330 75.940 112.650 ;
        RECT 76.660 112.310 76.800 129.330 ;
        RECT 77.580 128.290 77.720 129.930 ;
        RECT 77.980 129.670 78.240 129.990 ;
        RECT 77.060 127.970 77.320 128.290 ;
        RECT 77.520 127.970 77.780 128.290 ;
        RECT 77.120 126.930 77.260 127.970 ;
        RECT 77.580 126.930 77.720 127.970 ;
        RECT 77.060 126.610 77.320 126.930 ;
        RECT 77.520 126.610 77.780 126.930 ;
        RECT 77.980 125.590 78.240 125.910 ;
        RECT 78.040 123.530 78.180 125.590 ;
        RECT 77.060 123.210 77.320 123.530 ;
        RECT 77.980 123.210 78.240 123.530 ;
        RECT 77.120 122.850 77.260 123.210 ;
        RECT 77.060 122.530 77.320 122.850 ;
        RECT 77.060 119.810 77.320 120.130 ;
        RECT 77.120 116.390 77.260 119.810 ;
        RECT 78.500 119.110 78.640 131.030 ;
        RECT 78.960 128.970 79.100 134.010 ;
        RECT 79.360 131.710 79.620 132.030 ;
        RECT 79.880 131.940 80.020 150.330 ;
        RECT 80.280 149.730 80.540 150.050 ;
        RECT 80.340 144.950 80.480 149.730 ;
        RECT 80.800 146.310 80.940 150.750 ;
        RECT 80.740 145.990 81.000 146.310 ;
        RECT 81.260 145.290 81.400 150.750 ;
        RECT 82.180 148.690 82.320 166.730 ;
        RECT 82.640 164.670 82.780 166.730 ;
        RECT 82.580 164.350 82.840 164.670 ;
        RECT 82.640 155.230 82.780 164.350 ;
        RECT 83.100 156.170 83.240 171.490 ;
        RECT 83.560 168.070 83.700 172.170 ;
        RECT 84.880 171.830 85.140 172.150 ;
        RECT 85.340 171.830 85.600 172.150 ;
        RECT 85.800 171.830 86.060 172.150 ;
        RECT 83.960 171.490 84.220 171.810 ;
        RECT 83.500 167.750 83.760 168.070 ;
        RECT 83.500 164.010 83.760 164.330 ;
        RECT 83.560 160.785 83.700 164.010 ;
        RECT 83.490 160.415 83.770 160.785 ;
        RECT 83.490 157.695 83.770 158.065 ;
        RECT 83.040 155.850 83.300 156.170 ;
        RECT 82.640 155.090 83.240 155.230 ;
        RECT 83.100 153.790 83.240 155.090 ;
        RECT 83.040 153.470 83.300 153.790 ;
        RECT 82.580 152.790 82.840 153.110 ;
        RECT 82.120 148.600 82.380 148.690 ;
        RECT 81.720 148.460 82.380 148.600 ;
        RECT 81.200 144.970 81.460 145.290 ;
        RECT 80.280 144.630 80.540 144.950 ;
        RECT 81.260 142.910 81.400 144.970 ;
        RECT 80.280 142.590 80.540 142.910 ;
        RECT 81.200 142.590 81.460 142.910 ;
        RECT 80.340 140.870 80.480 142.590 ;
        RECT 80.280 140.550 80.540 140.870 ;
        RECT 80.740 138.850 81.000 139.170 ;
        RECT 80.800 138.150 80.940 138.850 ;
        RECT 80.740 137.830 81.000 138.150 ;
        RECT 81.260 137.810 81.400 142.590 ;
        RECT 81.200 137.490 81.460 137.810 ;
        RECT 80.740 136.810 81.000 137.130 ;
        RECT 80.800 135.430 80.940 136.810 ;
        RECT 80.740 135.110 81.000 135.430 ;
        RECT 81.260 134.750 81.400 137.490 ;
        RECT 81.200 134.430 81.460 134.750 ;
        RECT 81.260 132.030 81.400 134.430 ;
        RECT 81.720 132.370 81.860 148.460 ;
        RECT 82.120 148.370 82.380 148.460 ;
        RECT 82.120 144.290 82.380 144.610 ;
        RECT 82.180 138.150 82.320 144.290 ;
        RECT 82.120 137.830 82.380 138.150 ;
        RECT 82.640 137.470 82.780 152.790 ;
        RECT 83.100 151.750 83.240 153.470 ;
        RECT 83.560 153.110 83.700 157.695 ;
        RECT 84.020 154.130 84.160 171.490 ;
        RECT 84.940 170.450 85.080 171.830 ;
        RECT 84.880 170.130 85.140 170.450 ;
        RECT 85.400 170.190 85.540 171.830 ;
        RECT 85.860 171.665 86.000 171.830 ;
        RECT 85.790 171.295 86.070 171.665 ;
        RECT 85.400 170.110 86.460 170.190 ;
        RECT 85.400 170.050 86.520 170.110 ;
        RECT 86.260 169.790 86.520 170.050 ;
        RECT 84.880 169.450 85.140 169.770 ;
        RECT 85.800 169.450 86.060 169.770 ;
        RECT 84.420 168.770 84.680 169.090 ;
        RECT 84.940 168.945 85.080 169.450 ;
        RECT 84.480 168.265 84.620 168.770 ;
        RECT 84.870 168.575 85.150 168.945 ;
        RECT 84.410 167.895 84.690 168.265 ;
        RECT 85.860 163.990 86.000 169.450 ;
        RECT 86.320 167.390 86.460 169.790 ;
        RECT 87.240 168.945 87.380 172.170 ;
        RECT 87.640 171.830 87.900 172.150 ;
        RECT 87.170 168.575 87.450 168.945 ;
        RECT 86.720 167.410 86.980 167.730 ;
        RECT 86.260 167.070 86.520 167.390 ;
        RECT 85.800 163.670 86.060 163.990 ;
        RECT 85.340 163.330 85.600 163.650 ;
        RECT 84.420 158.910 84.680 159.230 ;
        RECT 84.480 157.190 84.620 158.910 ;
        RECT 84.420 156.870 84.680 157.190 ;
        RECT 84.880 156.190 85.140 156.510 ;
        RECT 83.960 153.810 84.220 154.130 ;
        RECT 83.960 153.130 84.220 153.450 ;
        RECT 83.500 152.790 83.760 153.110 ;
        RECT 83.040 151.430 83.300 151.750 ;
        RECT 83.040 150.070 83.300 150.390 ;
        RECT 83.100 149.030 83.240 150.070 ;
        RECT 83.500 149.730 83.760 150.050 ;
        RECT 83.040 148.710 83.300 149.030 ;
        RECT 83.560 147.865 83.700 149.730 ;
        RECT 83.490 147.495 83.770 147.865 ;
        RECT 83.500 144.630 83.760 144.950 ;
        RECT 83.040 144.290 83.300 144.610 ;
        RECT 83.100 141.890 83.240 144.290 ;
        RECT 83.040 141.570 83.300 141.890 ;
        RECT 82.580 137.150 82.840 137.470 ;
        RECT 82.580 133.750 82.840 134.070 ;
        RECT 81.660 132.050 81.920 132.370 ;
        RECT 79.880 131.800 80.940 131.940 ;
        RECT 79.420 129.650 79.560 131.710 ;
        RECT 80.280 131.030 80.540 131.350 ;
        RECT 79.820 130.690 80.080 131.010 ;
        RECT 79.880 130.185 80.020 130.690 ;
        RECT 79.810 129.815 80.090 130.185 ;
        RECT 79.360 129.330 79.620 129.650 ;
        RECT 78.900 128.650 79.160 128.970 ;
        RECT 78.960 127.350 79.100 128.650 ;
        RECT 78.960 127.210 80.020 127.350 ;
        RECT 78.890 123.695 79.170 124.065 ;
        RECT 78.960 123.530 79.100 123.695 ;
        RECT 78.900 123.210 79.160 123.530 ;
        RECT 78.440 118.790 78.700 119.110 ;
        RECT 77.520 118.110 77.780 118.430 ;
        RECT 77.980 118.110 78.240 118.430 ;
        RECT 78.960 118.410 79.100 123.210 ;
        RECT 79.360 120.830 79.620 121.150 ;
        RECT 78.500 118.270 79.100 118.410 ;
        RECT 77.060 116.070 77.320 116.390 ;
        RECT 77.580 113.070 77.720 118.110 ;
        RECT 78.040 114.690 78.180 118.110 ;
        RECT 78.500 116.050 78.640 118.270 ;
        RECT 78.900 117.430 79.160 117.750 ;
        RECT 78.960 116.390 79.100 117.430 ;
        RECT 79.420 116.390 79.560 120.830 ;
        RECT 78.900 116.070 79.160 116.390 ;
        RECT 79.360 116.070 79.620 116.390 ;
        RECT 78.440 115.730 78.700 116.050 ;
        RECT 77.980 114.370 78.240 114.690 ;
        RECT 78.500 113.330 78.640 115.730 ;
        RECT 77.120 112.930 77.720 113.070 ;
        RECT 78.440 113.010 78.700 113.330 ;
        RECT 76.600 111.990 76.860 112.310 ;
        RECT 75.220 104.850 75.480 105.170 ;
        RECT 74.760 96.010 75.020 96.330 ;
        RECT 74.820 71.850 74.960 96.010 ;
        RECT 75.280 90.550 75.420 104.850 ;
        RECT 76.140 104.170 76.400 104.490 ;
        RECT 76.200 102.450 76.340 104.170 ;
        RECT 76.140 102.130 76.400 102.450 ;
        RECT 76.200 101.770 76.340 102.130 ;
        RECT 76.140 101.450 76.400 101.770 ;
        RECT 76.140 99.750 76.400 100.070 ;
        RECT 76.200 96.330 76.340 99.750 ;
        RECT 75.670 95.815 75.950 96.185 ;
        RECT 76.140 96.010 76.400 96.330 ;
        RECT 75.740 94.630 75.880 95.815 ;
        RECT 75.680 94.310 75.940 94.630 ;
        RECT 76.660 94.030 76.800 111.990 ;
        RECT 77.120 102.790 77.260 112.930 ;
        RECT 78.960 112.650 79.100 116.070 ;
        RECT 79.880 115.790 80.020 127.210 ;
        RECT 80.340 118.430 80.480 131.030 ;
        RECT 80.800 122.850 80.940 131.800 ;
        RECT 81.200 131.710 81.460 132.030 ;
        RECT 81.720 131.430 81.860 132.050 ;
        RECT 81.260 131.350 81.860 131.430 ;
        RECT 81.200 131.290 81.860 131.350 ;
        RECT 81.200 131.030 81.460 131.290 ;
        RECT 82.640 131.010 82.780 133.750 ;
        RECT 82.580 130.690 82.840 131.010 ;
        RECT 83.040 130.690 83.300 131.010 ;
        RECT 81.200 129.670 81.460 129.990 ;
        RECT 82.110 129.815 82.390 130.185 ;
        RECT 81.260 128.970 81.400 129.670 ;
        RECT 82.180 129.650 82.320 129.815 ;
        RECT 82.120 129.330 82.380 129.650 ;
        RECT 81.200 128.650 81.460 128.970 ;
        RECT 81.660 128.650 81.920 128.970 ;
        RECT 81.720 127.270 81.860 128.650 ;
        RECT 81.660 126.950 81.920 127.270 ;
        RECT 82.570 127.095 82.850 127.465 ;
        RECT 82.120 126.270 82.380 126.590 ;
        RECT 80.740 122.530 81.000 122.850 ;
        RECT 80.280 118.110 80.540 118.430 ;
        RECT 80.800 117.150 80.940 122.530 ;
        RECT 82.180 121.830 82.320 126.270 ;
        RECT 82.640 126.250 82.780 127.095 ;
        RECT 82.580 125.930 82.840 126.250 ;
        RECT 83.100 125.570 83.240 130.690 ;
        RECT 83.560 128.630 83.700 144.630 ;
        RECT 84.020 144.610 84.160 153.130 ;
        RECT 84.420 150.410 84.680 150.730 ;
        RECT 84.480 148.350 84.620 150.410 ;
        RECT 84.420 148.030 84.680 148.350 ;
        RECT 84.940 144.950 85.080 156.190 ;
        RECT 85.400 148.350 85.540 163.330 ;
        RECT 86.250 159.055 86.530 159.425 ;
        RECT 85.800 157.890 86.060 158.210 ;
        RECT 85.860 156.170 86.000 157.890 ;
        RECT 85.800 155.850 86.060 156.170 ;
        RECT 86.320 154.550 86.460 159.055 ;
        RECT 85.860 154.470 86.460 154.550 ;
        RECT 85.860 154.410 86.520 154.470 ;
        RECT 85.860 148.350 86.000 154.410 ;
        RECT 86.260 154.150 86.520 154.410 ;
        RECT 86.250 153.615 86.530 153.985 ;
        RECT 86.780 153.790 86.920 167.410 ;
        RECT 87.240 167.050 87.380 168.575 ;
        RECT 87.180 166.730 87.440 167.050 ;
        RECT 87.180 166.050 87.440 166.370 ;
        RECT 86.260 153.470 86.520 153.615 ;
        RECT 86.720 153.470 86.980 153.790 ;
        RECT 87.240 148.350 87.380 166.050 ;
        RECT 87.700 159.910 87.840 171.830 ;
        RECT 88.560 167.070 88.820 167.390 ;
        RECT 88.090 164.495 88.370 164.865 ;
        RECT 88.100 164.350 88.360 164.495 ;
        RECT 88.100 163.670 88.360 163.990 ;
        RECT 88.160 162.630 88.300 163.670 ;
        RECT 88.100 162.310 88.360 162.630 ;
        RECT 87.640 159.590 87.900 159.910 ;
        RECT 88.090 154.295 88.370 154.665 ;
        RECT 88.160 153.790 88.300 154.295 ;
        RECT 88.100 153.470 88.360 153.790 ;
        RECT 85.340 148.030 85.600 148.350 ;
        RECT 85.800 148.030 86.060 148.350 ;
        RECT 87.180 148.030 87.440 148.350 ;
        RECT 88.100 148.030 88.360 148.350 ;
        RECT 85.340 147.350 85.600 147.670 ;
        RECT 85.400 145.290 85.540 147.350 ;
        RECT 87.640 147.010 87.900 147.330 ;
        RECT 85.340 144.970 85.600 145.290 ;
        RECT 86.720 144.970 86.980 145.290 ;
        RECT 87.180 144.970 87.440 145.290 ;
        RECT 84.880 144.630 85.140 144.950 ;
        RECT 83.960 144.290 84.220 144.610 ;
        RECT 84.420 144.290 84.680 144.610 ;
        RECT 84.480 143.250 84.620 144.290 ;
        RECT 84.420 142.930 84.680 143.250 ;
        RECT 84.420 137.150 84.680 137.470 ;
        RECT 84.880 137.150 85.140 137.470 ;
        RECT 84.480 134.945 84.620 137.150 ;
        RECT 84.410 134.575 84.690 134.945 ;
        RECT 84.420 133.410 84.680 133.730 ;
        RECT 83.960 131.710 84.220 132.030 ;
        RECT 84.020 129.990 84.160 131.710 ;
        RECT 84.480 129.990 84.620 133.410 ;
        RECT 84.940 131.010 85.080 137.150 ;
        RECT 85.400 132.710 85.540 144.970 ;
        RECT 85.800 139.705 86.060 139.850 ;
        RECT 85.790 139.335 86.070 139.705 ;
        RECT 85.800 136.130 86.060 136.450 ;
        RECT 85.340 132.390 85.600 132.710 ;
        RECT 85.860 132.110 86.000 136.130 ;
        RECT 85.400 131.970 86.000 132.110 ;
        RECT 84.880 130.690 85.140 131.010 ;
        RECT 83.960 129.670 84.220 129.990 ;
        RECT 84.420 129.670 84.680 129.990 ;
        RECT 84.420 128.650 84.680 128.970 ;
        RECT 83.500 128.540 83.760 128.630 ;
        RECT 83.500 128.400 84.160 128.540 ;
        RECT 83.500 128.310 83.760 128.400 ;
        RECT 83.500 126.270 83.760 126.590 ;
        RECT 83.040 125.250 83.300 125.570 ;
        RECT 82.570 123.695 82.850 124.065 ;
        RECT 82.120 121.510 82.380 121.830 ;
        RECT 81.660 120.150 81.920 120.470 ;
        RECT 81.200 118.790 81.460 119.110 ;
        RECT 80.340 117.010 80.940 117.150 ;
        RECT 80.340 116.050 80.480 117.010 ;
        RECT 81.260 116.300 81.400 118.790 ;
        RECT 80.800 116.160 81.400 116.300 ;
        RECT 79.420 115.650 80.020 115.790 ;
        RECT 80.280 115.730 80.540 116.050 ;
        RECT 77.520 112.330 77.780 112.650 ;
        RECT 78.900 112.330 79.160 112.650 ;
        RECT 77.580 109.250 77.720 112.330 ;
        RECT 78.440 111.990 78.700 112.310 ;
        RECT 78.500 110.950 78.640 111.990 ;
        RECT 78.440 110.630 78.700 110.950 ;
        RECT 77.520 108.930 77.780 109.250 ;
        RECT 77.580 107.210 77.720 108.930 ;
        RECT 77.520 107.120 77.780 107.210 ;
        RECT 77.520 106.980 78.180 107.120 ;
        RECT 77.520 106.890 77.780 106.980 ;
        RECT 78.040 104.490 78.180 106.980 ;
        RECT 78.440 106.550 78.700 106.870 ;
        RECT 78.500 105.510 78.640 106.550 ;
        RECT 79.420 105.510 79.560 115.650 ;
        RECT 80.340 112.220 80.480 115.730 ;
        RECT 79.880 112.080 80.480 112.220 ;
        RECT 79.880 110.610 80.020 112.080 ;
        RECT 80.800 111.710 80.940 116.160 ;
        RECT 81.720 115.710 81.860 120.150 ;
        RECT 82.180 118.090 82.320 121.510 ;
        RECT 82.120 117.770 82.380 118.090 ;
        RECT 82.640 117.410 82.780 123.695 ;
        RECT 83.560 122.850 83.700 126.270 ;
        RECT 84.020 124.550 84.160 128.400 ;
        RECT 84.480 126.590 84.620 128.650 ;
        RECT 84.420 126.270 84.680 126.590 ;
        RECT 84.880 125.930 85.140 126.250 ;
        RECT 83.960 124.230 84.220 124.550 ;
        RECT 83.500 122.530 83.760 122.850 ;
        RECT 83.030 120.295 83.310 120.665 ;
        RECT 83.100 117.750 83.240 120.295 ;
        RECT 83.560 118.090 83.700 122.530 ;
        RECT 83.500 117.770 83.760 118.090 ;
        RECT 83.040 117.430 83.300 117.750 ;
        RECT 82.580 117.090 82.840 117.410 ;
        RECT 81.200 115.390 81.460 115.710 ;
        RECT 81.660 115.390 81.920 115.710 ;
        RECT 81.260 114.690 81.400 115.390 ;
        RECT 83.500 114.710 83.760 115.030 ;
        RECT 81.200 114.370 81.460 114.690 ;
        RECT 80.340 111.570 80.940 111.710 ;
        RECT 80.340 110.610 80.480 111.570 ;
        RECT 80.730 110.775 81.010 111.145 ;
        RECT 80.740 110.630 81.000 110.775 ;
        RECT 79.820 110.290 80.080 110.610 ;
        RECT 80.280 110.290 80.540 110.610 ;
        RECT 80.280 108.140 80.540 108.230 ;
        RECT 79.880 108.000 80.540 108.140 ;
        RECT 78.440 105.190 78.700 105.510 ;
        RECT 79.360 105.190 79.620 105.510 ;
        RECT 78.430 104.655 78.710 105.025 ;
        RECT 79.360 104.740 79.620 104.830 ;
        RECT 77.980 104.170 78.240 104.490 ;
        RECT 77.510 103.295 77.790 103.665 ;
        RECT 77.060 102.470 77.320 102.790 ;
        RECT 77.580 100.070 77.720 103.295 ;
        RECT 77.520 99.750 77.780 100.070 ;
        RECT 78.040 99.390 78.180 104.170 ;
        RECT 77.980 99.070 78.240 99.390 ;
        RECT 77.060 98.390 77.320 98.710 ;
        RECT 77.120 96.330 77.260 98.390 ;
        RECT 77.060 96.010 77.320 96.330 ;
        RECT 77.980 96.010 78.240 96.330 ;
        RECT 76.660 93.950 77.260 94.030 ;
        RECT 76.140 93.630 76.400 93.950 ;
        RECT 76.660 93.890 77.320 93.950 ;
        RECT 77.060 93.630 77.320 93.890 ;
        RECT 75.680 91.250 75.940 91.570 ;
        RECT 75.220 90.230 75.480 90.550 ;
        RECT 75.220 85.810 75.480 86.130 ;
        RECT 75.280 82.050 75.420 85.810 ;
        RECT 75.740 84.770 75.880 91.250 ;
        RECT 76.200 89.950 76.340 93.630 ;
        RECT 76.600 90.745 76.860 90.890 ;
        RECT 76.590 90.375 76.870 90.745 ;
        RECT 76.600 89.950 76.860 90.210 ;
        RECT 76.200 89.890 76.860 89.950 ;
        RECT 76.200 89.810 76.800 89.890 ;
        RECT 76.200 88.510 76.340 89.810 ;
        RECT 77.120 88.850 77.260 93.630 ;
        RECT 78.040 92.930 78.180 96.010 ;
        RECT 77.980 92.610 78.240 92.930 ;
        RECT 77.060 88.530 77.320 88.850 ;
        RECT 78.500 88.590 78.640 104.655 ;
        RECT 78.960 104.600 79.620 104.740 ;
        RECT 78.960 94.630 79.100 104.600 ;
        RECT 79.360 104.510 79.620 104.600 ;
        RECT 79.880 101.770 80.020 108.000 ;
        RECT 80.280 107.910 80.540 108.000 ;
        RECT 81.260 105.590 81.400 114.370 ;
        RECT 82.120 113.350 82.380 113.670 ;
        RECT 81.660 111.990 81.920 112.310 ;
        RECT 81.720 110.950 81.860 111.990 ;
        RECT 82.180 110.950 82.320 113.350 ;
        RECT 81.660 110.630 81.920 110.950 ;
        RECT 82.120 110.630 82.380 110.950 ;
        RECT 83.560 110.270 83.700 114.710 ;
        RECT 83.500 109.950 83.760 110.270 ;
        RECT 84.020 109.930 84.160 124.230 ;
        RECT 84.420 115.730 84.680 116.050 ;
        RECT 84.480 110.270 84.620 115.730 ;
        RECT 84.420 109.950 84.680 110.270 ;
        RECT 83.960 109.610 84.220 109.930 ;
        RECT 83.500 109.270 83.760 109.590 ;
        RECT 82.570 106.695 82.850 107.065 ;
        RECT 82.640 106.530 82.780 106.695 ;
        RECT 82.580 106.210 82.840 106.530 ;
        RECT 80.800 105.450 81.400 105.590 ;
        RECT 79.820 101.450 80.080 101.770 ;
        RECT 80.280 101.450 80.540 101.770 ;
        RECT 79.360 99.070 79.620 99.390 ;
        RECT 79.420 97.350 79.560 99.070 ;
        RECT 79.360 97.030 79.620 97.350 ;
        RECT 78.900 94.310 79.160 94.630 ;
        RECT 79.880 94.030 80.020 101.450 ;
        RECT 80.340 94.630 80.480 101.450 ;
        RECT 80.800 97.010 80.940 105.450 ;
        RECT 81.200 104.850 81.460 105.170 ;
        RECT 80.740 96.690 81.000 97.010 ;
        RECT 80.800 95.390 80.940 96.690 ;
        RECT 81.260 96.330 81.400 104.850 ;
        RECT 81.660 104.510 81.920 104.830 ;
        RECT 81.720 102.790 81.860 104.510 ;
        RECT 82.120 103.490 82.380 103.810 ;
        RECT 81.660 102.470 81.920 102.790 ;
        RECT 82.180 101.770 82.320 103.490 ;
        RECT 83.560 102.790 83.700 109.270 ;
        RECT 83.500 102.470 83.760 102.790 ;
        RECT 82.580 102.130 82.840 102.450 ;
        RECT 83.560 102.305 83.700 102.470 ;
        RECT 82.120 101.450 82.380 101.770 ;
        RECT 82.180 97.350 82.320 101.450 ;
        RECT 82.120 97.030 82.380 97.350 ;
        RECT 81.200 96.010 81.460 96.330 ;
        RECT 80.800 95.250 81.400 95.390 ;
        RECT 81.660 95.330 81.920 95.650 ;
        RECT 80.280 94.310 80.540 94.630 ;
        RECT 79.420 93.950 80.020 94.030 ;
        RECT 79.360 93.890 80.020 93.950 ;
        RECT 79.360 93.630 79.620 93.890 ;
        RECT 80.730 93.775 81.010 94.145 ;
        RECT 80.740 93.630 81.000 93.775 ;
        RECT 79.810 93.095 80.090 93.465 ;
        RECT 80.280 93.290 80.540 93.610 ;
        RECT 78.890 90.375 79.170 90.745 ;
        RECT 76.140 88.190 76.400 88.510 ;
        RECT 77.120 87.830 77.260 88.530 ;
        RECT 78.040 88.450 78.640 88.590 ;
        RECT 77.060 87.510 77.320 87.830 ;
        RECT 76.600 86.150 76.860 86.470 ;
        RECT 75.680 84.450 75.940 84.770 ;
        RECT 75.680 82.410 75.940 82.730 ;
        RECT 75.220 81.730 75.480 82.050 ;
        RECT 75.740 79.330 75.880 82.410 ;
        RECT 76.660 80.690 76.800 86.150 ;
        RECT 77.520 85.130 77.780 85.450 ;
        RECT 77.050 82.895 77.330 83.265 ;
        RECT 77.060 82.750 77.320 82.895 ;
        RECT 76.600 80.370 76.860 80.690 ;
        RECT 76.140 80.030 76.400 80.350 ;
        RECT 75.680 79.010 75.940 79.330 ;
        RECT 75.210 77.455 75.490 77.825 ;
        RECT 76.200 77.630 76.340 80.030 ;
        RECT 74.760 71.530 75.020 71.850 ;
        RECT 74.300 71.190 74.560 71.510 ;
        RECT 74.300 69.150 74.560 69.470 ;
        RECT 73.830 68.615 74.110 68.985 ;
        RECT 73.900 64.710 74.040 68.615 ;
        RECT 74.360 67.430 74.500 69.150 ;
        RECT 74.300 67.110 74.560 67.430 ;
        RECT 74.820 66.660 74.960 71.530 ;
        RECT 75.280 67.430 75.420 77.455 ;
        RECT 76.140 77.310 76.400 77.630 ;
        RECT 75.680 76.970 75.940 77.290 ;
        RECT 75.740 75.250 75.880 76.970 ;
        RECT 76.660 76.950 76.800 80.370 ;
        RECT 77.580 78.310 77.720 85.130 ;
        RECT 77.520 77.990 77.780 78.310 ;
        RECT 76.600 76.630 76.860 76.950 ;
        RECT 76.140 75.270 76.400 75.590 ;
        RECT 75.680 74.930 75.940 75.250 ;
        RECT 76.200 74.480 76.340 75.270 ;
        RECT 75.740 74.340 76.340 74.480 ;
        RECT 75.220 67.110 75.480 67.430 ;
        RECT 74.820 66.520 75.420 66.660 ;
        RECT 74.750 65.895 75.030 66.265 ;
        RECT 72.920 64.480 73.580 64.620 ;
        RECT 72.920 64.390 73.180 64.480 ;
        RECT 73.840 64.390 74.100 64.710 ;
        RECT 71.080 58.270 71.340 58.590 ;
        RECT 72.450 58.415 72.730 58.785 ;
        RECT 71.140 56.745 71.280 58.270 ;
        RECT 72.520 58.250 72.660 58.415 ;
        RECT 72.460 57.930 72.720 58.250 ;
        RECT 72.000 57.590 72.260 57.910 ;
        RECT 71.070 56.375 71.350 56.745 ;
        RECT 71.080 56.230 71.340 56.375 ;
        RECT 71.140 51.110 71.280 56.230 ;
        RECT 72.060 55.870 72.200 57.590 ;
        RECT 73.900 56.310 74.040 64.390 ;
        RECT 74.820 61.990 74.960 65.895 ;
        RECT 74.760 61.670 75.020 61.990 ;
        RECT 73.900 56.170 74.960 56.310 ;
        RECT 72.000 55.550 72.260 55.870 ;
        RECT 73.380 55.550 73.640 55.870 ;
        RECT 72.920 54.530 73.180 54.850 ;
        RECT 71.080 50.790 71.340 51.110 ;
        RECT 69.760 50.370 70.360 50.510 ;
        RECT 70.620 50.450 70.880 50.770 ;
        RECT 69.240 47.390 69.500 47.710 ;
        RECT 69.300 45.330 69.440 47.390 ;
        RECT 69.240 45.010 69.500 45.330 ;
        RECT 69.760 41.930 69.900 50.370 ;
        RECT 70.160 48.070 70.420 48.390 ;
        RECT 69.700 41.610 69.960 41.930 ;
        RECT 70.220 38.530 70.360 48.070 ;
        RECT 70.680 48.050 70.820 50.450 ;
        RECT 72.000 49.770 72.260 50.090 ;
        RECT 71.540 49.090 71.800 49.410 ;
        RECT 70.620 47.730 70.880 48.050 ;
        RECT 71.080 47.050 71.340 47.370 ;
        RECT 70.610 45.495 70.890 45.865 ;
        RECT 70.680 38.530 70.820 45.495 ;
        RECT 71.140 39.890 71.280 47.050 ;
        RECT 71.600 44.310 71.740 49.090 ;
        RECT 71.540 43.990 71.800 44.310 ;
        RECT 71.600 41.590 71.740 43.990 ;
        RECT 71.540 41.270 71.800 41.590 ;
        RECT 72.060 40.230 72.200 49.770 ;
        RECT 72.980 47.225 73.120 54.530 ;
        RECT 73.440 51.110 73.580 55.550 ;
        RECT 73.840 53.510 74.100 53.830 ;
        RECT 73.380 50.790 73.640 51.110 ;
        RECT 73.380 49.770 73.640 50.090 ;
        RECT 72.910 46.855 73.190 47.225 ;
        RECT 72.460 44.670 72.720 44.990 ;
        RECT 72.520 42.950 72.660 44.670 ;
        RECT 72.460 42.630 72.720 42.950 ;
        RECT 72.980 41.930 73.120 46.855 ;
        RECT 73.440 41.930 73.580 49.770 ;
        RECT 73.900 48.390 74.040 53.510 ;
        RECT 74.300 52.490 74.560 52.810 ;
        RECT 73.840 48.070 74.100 48.390 ;
        RECT 74.360 47.370 74.500 52.490 ;
        RECT 74.820 50.340 74.960 56.170 ;
        RECT 75.280 51.110 75.420 66.520 ;
        RECT 75.740 63.690 75.880 74.340 ;
        RECT 76.660 69.810 76.800 76.630 ;
        RECT 77.580 75.670 77.720 77.990 ;
        RECT 77.120 75.530 77.720 75.670 ;
        RECT 77.120 74.570 77.260 75.530 ;
        RECT 77.520 74.930 77.780 75.250 ;
        RECT 77.060 74.250 77.320 74.570 ;
        RECT 77.060 73.570 77.320 73.890 ;
        RECT 77.120 72.870 77.260 73.570 ;
        RECT 77.060 72.550 77.320 72.870 ;
        RECT 77.580 72.530 77.720 74.930 ;
        RECT 77.520 72.210 77.780 72.530 ;
        RECT 77.520 70.850 77.780 71.170 ;
        RECT 76.600 69.490 76.860 69.810 ;
        RECT 77.580 69.130 77.720 70.850 ;
        RECT 76.140 68.810 76.400 69.130 ;
        RECT 77.520 68.810 77.780 69.130 ;
        RECT 76.200 68.450 76.340 68.810 ;
        RECT 76.140 68.130 76.400 68.450 ;
        RECT 76.590 67.935 76.870 68.305 ;
        RECT 77.060 68.130 77.320 68.450 ;
        RECT 76.140 66.430 76.400 66.750 ;
        RECT 76.200 64.030 76.340 66.430 ;
        RECT 76.660 66.070 76.800 67.935 ;
        RECT 77.120 66.750 77.260 68.130 ;
        RECT 77.060 66.430 77.320 66.750 ;
        RECT 76.600 65.750 76.860 66.070 ;
        RECT 77.580 64.710 77.720 68.810 ;
        RECT 78.040 66.410 78.180 88.450 ;
        RECT 78.440 84.450 78.700 84.770 ;
        RECT 78.500 77.290 78.640 84.450 ;
        RECT 78.960 83.070 79.100 90.375 ;
        RECT 79.360 90.230 79.620 90.550 ;
        RECT 79.420 87.830 79.560 90.230 ;
        RECT 79.880 88.510 80.020 93.095 ;
        RECT 80.340 91.310 80.480 93.290 ;
        RECT 81.260 91.990 81.400 95.250 ;
        RECT 81.720 93.950 81.860 95.330 ;
        RECT 82.110 94.030 82.390 94.145 ;
        RECT 82.640 94.030 82.780 102.130 ;
        RECT 83.490 101.935 83.770 102.305 ;
        RECT 84.020 102.110 84.160 109.610 ;
        RECT 84.480 105.170 84.620 109.950 ;
        RECT 84.940 107.745 85.080 125.930 ;
        RECT 85.400 121.490 85.540 131.970 ;
        RECT 85.800 130.690 86.060 131.010 ;
        RECT 85.860 128.630 86.000 130.690 ;
        RECT 85.800 128.310 86.060 128.630 ;
        RECT 86.260 128.310 86.520 128.630 ;
        RECT 86.320 126.250 86.460 128.310 ;
        RECT 86.260 125.930 86.520 126.250 ;
        RECT 86.780 121.830 86.920 144.970 ;
        RECT 87.240 139.850 87.380 144.970 ;
        RECT 87.180 139.530 87.440 139.850 ;
        RECT 87.700 137.665 87.840 147.010 ;
        RECT 88.160 141.890 88.300 148.030 ;
        RECT 88.100 141.570 88.360 141.890 ;
        RECT 87.630 137.295 87.910 137.665 ;
        RECT 87.640 136.810 87.900 137.130 ;
        RECT 87.700 133.730 87.840 136.810 ;
        RECT 87.640 133.410 87.900 133.730 ;
        RECT 87.700 132.370 87.840 133.410 ;
        RECT 87.640 132.050 87.900 132.370 ;
        RECT 87.700 128.970 87.840 132.050 ;
        RECT 87.640 128.650 87.900 128.970 ;
        RECT 87.180 125.930 87.440 126.250 ;
        RECT 86.720 121.510 86.980 121.830 ;
        RECT 85.340 121.170 85.600 121.490 ;
        RECT 84.870 107.375 85.150 107.745 ;
        RECT 84.880 106.890 85.140 107.210 ;
        RECT 84.420 104.850 84.680 105.170 ;
        RECT 84.940 105.025 85.080 106.890 ;
        RECT 83.960 101.790 84.220 102.110 ;
        RECT 83.500 101.450 83.760 101.770 ;
        RECT 83.560 100.070 83.700 101.450 ;
        RECT 83.500 99.750 83.760 100.070 ;
        RECT 83.500 98.110 83.760 98.370 ;
        RECT 83.100 98.050 83.760 98.110 ;
        RECT 83.100 97.970 83.700 98.050 ;
        RECT 83.100 95.990 83.240 97.970 ;
        RECT 83.040 95.670 83.300 95.990 ;
        RECT 83.100 94.290 83.240 95.670 ;
        RECT 81.660 93.630 81.920 93.950 ;
        RECT 82.110 93.890 82.780 94.030 ;
        RECT 83.040 93.970 83.300 94.290 ;
        RECT 82.110 93.775 82.390 93.890 ;
        RECT 83.500 93.630 83.760 93.950 ;
        RECT 81.660 92.950 81.920 93.270 ;
        RECT 82.570 93.095 82.850 93.465 ;
        RECT 82.580 92.950 82.840 93.095 ;
        RECT 81.720 92.670 81.860 92.950 ;
        RECT 81.720 92.530 82.780 92.670 ;
        RECT 81.260 91.850 82.320 91.990 ;
        RECT 80.340 91.170 81.400 91.310 ;
        RECT 80.280 90.745 80.540 90.890 ;
        RECT 80.270 90.375 80.550 90.745 ;
        RECT 80.740 90.230 81.000 90.550 ;
        RECT 79.820 88.190 80.080 88.510 ;
        RECT 79.360 87.510 79.620 87.830 ;
        RECT 78.900 82.750 79.160 83.070 ;
        RECT 79.420 80.010 79.560 87.510 ;
        RECT 79.880 86.470 80.020 88.190 ;
        RECT 80.800 86.470 80.940 90.230 ;
        RECT 81.260 88.850 81.400 91.170 ;
        RECT 82.180 90.550 82.320 91.850 ;
        RECT 82.120 90.230 82.380 90.550 ;
        RECT 81.660 89.890 81.920 90.210 ;
        RECT 82.640 90.065 82.780 92.530 ;
        RECT 83.560 91.910 83.700 93.630 ;
        RECT 84.020 92.930 84.160 101.790 ;
        RECT 84.480 101.770 84.620 104.850 ;
        RECT 84.870 104.655 85.150 105.025 ;
        RECT 85.400 102.190 85.540 121.170 ;
        RECT 86.260 117.770 86.520 118.090 ;
        RECT 86.720 117.770 86.980 118.090 ;
        RECT 85.800 117.265 86.060 117.410 ;
        RECT 85.790 116.895 86.070 117.265 ;
        RECT 85.800 115.620 86.060 115.710 ;
        RECT 86.320 115.620 86.460 117.770 ;
        RECT 86.780 116.390 86.920 117.770 ;
        RECT 86.720 116.070 86.980 116.390 ;
        RECT 85.800 115.480 86.460 115.620 ;
        RECT 85.800 115.390 86.060 115.480 ;
        RECT 85.800 114.710 86.060 115.030 ;
        RECT 84.940 102.050 85.540 102.190 ;
        RECT 84.420 101.450 84.680 101.770 ;
        RECT 84.940 100.150 85.080 102.050 ;
        RECT 85.340 101.110 85.600 101.430 ;
        RECT 84.480 100.010 85.080 100.150 ;
        RECT 84.480 96.670 84.620 100.010 ;
        RECT 85.400 99.730 85.540 101.110 ;
        RECT 85.340 99.410 85.600 99.730 ;
        RECT 85.860 99.390 86.000 114.710 ;
        RECT 86.320 111.970 86.460 115.480 ;
        RECT 86.720 115.390 86.980 115.710 ;
        RECT 86.260 111.650 86.520 111.970 ;
        RECT 86.320 107.210 86.460 111.650 ;
        RECT 86.780 111.145 86.920 115.390 ;
        RECT 86.710 110.775 86.990 111.145 ;
        RECT 87.240 110.860 87.380 125.930 ;
        RECT 88.160 121.150 88.300 141.570 ;
        RECT 88.620 128.630 88.760 167.070 ;
        RECT 88.560 128.310 88.820 128.630 ;
        RECT 89.080 126.930 89.220 173.190 ;
        RECT 89.020 126.610 89.280 126.930 ;
        RECT 89.080 121.490 89.220 126.610 ;
        RECT 89.020 121.170 89.280 121.490 ;
        RECT 88.100 120.830 88.360 121.150 ;
        RECT 87.640 117.090 87.900 117.410 ;
        RECT 87.700 113.865 87.840 117.090 ;
        RECT 89.080 115.370 89.220 121.170 ;
        RECT 89.020 115.050 89.280 115.370 ;
        RECT 88.100 114.370 88.360 114.690 ;
        RECT 87.630 113.495 87.910 113.865 ;
        RECT 86.780 110.270 86.920 110.775 ;
        RECT 87.240 110.720 87.840 110.860 ;
        RECT 86.720 109.950 86.980 110.270 ;
        RECT 87.180 109.950 87.440 110.270 ;
        RECT 87.240 108.230 87.380 109.950 ;
        RECT 87.180 107.910 87.440 108.230 ;
        RECT 87.700 107.210 87.840 110.720 ;
        RECT 88.160 110.465 88.300 114.370 ;
        RECT 88.090 110.095 88.370 110.465 ;
        RECT 88.100 109.610 88.360 109.930 ;
        RECT 88.160 107.550 88.300 109.610 ;
        RECT 88.100 107.230 88.360 107.550 ;
        RECT 88.550 107.375 88.830 107.745 ;
        RECT 86.260 106.890 86.520 107.210 ;
        RECT 87.640 106.890 87.900 107.210 ;
        RECT 86.720 106.210 86.980 106.530 ;
        RECT 86.260 103.490 86.520 103.810 ;
        RECT 86.320 101.430 86.460 103.490 ;
        RECT 86.780 101.430 86.920 106.210 ;
        RECT 87.180 101.680 87.440 101.770 ;
        RECT 87.700 101.680 87.840 106.890 ;
        RECT 87.180 101.540 87.840 101.680 ;
        RECT 88.100 101.625 88.360 101.770 ;
        RECT 87.180 101.450 87.440 101.540 ;
        RECT 86.260 101.110 86.520 101.430 ;
        RECT 86.720 101.110 86.980 101.430 ;
        RECT 88.090 101.255 88.370 101.625 ;
        RECT 84.880 99.070 85.140 99.390 ;
        RECT 85.800 99.070 86.060 99.390 ;
        RECT 84.420 96.350 84.680 96.670 ;
        RECT 84.940 95.990 85.080 99.070 ;
        RECT 86.780 96.070 86.920 101.110 ;
        RECT 87.640 96.350 87.900 96.670 ;
        RECT 88.090 96.495 88.370 96.865 ;
        RECT 84.880 95.670 85.140 95.990 ;
        RECT 85.800 95.670 86.060 95.990 ;
        RECT 86.780 95.930 87.380 96.070 ;
        RECT 84.420 93.290 84.680 93.610 ;
        RECT 83.960 92.610 84.220 92.930 ;
        RECT 83.500 91.590 83.760 91.910 ;
        RECT 84.020 91.230 84.160 92.610 ;
        RECT 84.480 92.105 84.620 93.290 ;
        RECT 84.410 91.735 84.690 92.105 ;
        RECT 83.960 90.910 84.220 91.230 ;
        RECT 81.200 88.530 81.460 88.850 ;
        RECT 79.820 86.150 80.080 86.470 ;
        RECT 80.740 86.380 81.000 86.470 ;
        RECT 80.340 86.240 81.000 86.380 ;
        RECT 79.880 84.770 80.020 86.150 ;
        RECT 79.820 84.450 80.080 84.770 ;
        RECT 79.810 82.895 80.090 83.265 ;
        RECT 80.340 83.070 80.480 86.240 ;
        RECT 80.740 86.150 81.000 86.240 ;
        RECT 81.260 85.450 81.400 88.530 ;
        RECT 81.720 85.790 81.860 89.890 ;
        RECT 82.570 89.695 82.850 90.065 ;
        RECT 84.420 89.890 84.680 90.210 ;
        RECT 82.110 89.015 82.390 89.385 ;
        RECT 81.660 85.470 81.920 85.790 ;
        RECT 81.200 85.130 81.460 85.450 ;
        RECT 79.360 79.690 79.620 80.010 ;
        RECT 79.420 77.290 79.560 79.690 ;
        RECT 78.440 76.970 78.700 77.290 ;
        RECT 79.360 76.970 79.620 77.290 ;
        RECT 78.500 74.990 78.640 76.970 ;
        RECT 78.500 74.910 79.100 74.990 ;
        RECT 78.440 74.850 79.100 74.910 ;
        RECT 78.440 74.590 78.700 74.850 ;
        RECT 78.440 71.870 78.700 72.190 ;
        RECT 78.500 67.510 78.640 71.870 ;
        RECT 78.960 68.305 79.100 74.850 ;
        RECT 79.420 68.790 79.560 76.970 ;
        RECT 79.880 73.890 80.020 82.895 ;
        RECT 80.280 82.750 80.540 83.070 ;
        RECT 80.740 82.070 81.000 82.390 ;
        RECT 80.280 81.730 80.540 82.050 ;
        RECT 80.340 80.010 80.480 81.730 ;
        RECT 80.280 79.690 80.540 80.010 ;
        RECT 80.280 73.910 80.540 74.230 ;
        RECT 79.820 73.570 80.080 73.890 ;
        RECT 80.340 71.850 80.480 73.910 ;
        RECT 79.820 71.530 80.080 71.850 ;
        RECT 80.280 71.530 80.540 71.850 ;
        RECT 79.880 69.810 80.020 71.530 ;
        RECT 79.820 69.490 80.080 69.810 ;
        RECT 79.360 68.470 79.620 68.790 ;
        RECT 80.340 68.450 80.480 71.530 ;
        RECT 80.800 71.170 80.940 82.070 ;
        RECT 81.260 79.330 81.400 85.130 ;
        RECT 81.660 82.980 81.920 83.070 ;
        RECT 82.180 82.980 82.320 89.015 ;
        RECT 83.040 88.870 83.300 89.190 ;
        RECT 83.100 86.665 83.240 88.870 ;
        RECT 84.480 88.850 84.620 89.890 ;
        RECT 84.420 88.530 84.680 88.850 ;
        RECT 84.940 88.510 85.080 95.670 ;
        RECT 85.340 93.630 85.600 93.950 ;
        RECT 85.400 91.425 85.540 93.630 ;
        RECT 85.330 91.055 85.610 91.425 ;
        RECT 85.340 90.230 85.600 90.550 ;
        RECT 85.400 89.385 85.540 90.230 ;
        RECT 85.330 89.015 85.610 89.385 ;
        RECT 84.880 88.190 85.140 88.510 ;
        RECT 85.860 87.490 86.000 95.670 ;
        RECT 86.720 95.330 86.980 95.650 ;
        RECT 86.780 90.890 86.920 95.330 ;
        RECT 86.720 90.570 86.980 90.890 ;
        RECT 85.800 87.170 86.060 87.490 ;
        RECT 86.720 87.170 86.980 87.490 ;
        RECT 83.030 86.295 83.310 86.665 ;
        RECT 83.030 85.615 83.310 85.985 ;
        RECT 83.100 85.450 83.240 85.615 ;
        RECT 86.780 85.450 86.920 87.170 ;
        RECT 87.240 85.450 87.380 95.930 ;
        RECT 83.040 85.130 83.300 85.450 ;
        RECT 84.420 85.130 84.680 85.450 ;
        RECT 86.720 85.130 86.980 85.450 ;
        RECT 87.180 85.130 87.440 85.450 ;
        RECT 81.660 82.840 82.320 82.980 ;
        RECT 81.660 82.750 81.920 82.840 ;
        RECT 81.720 82.390 81.860 82.750 ;
        RECT 81.660 82.070 81.920 82.390 ;
        RECT 82.120 81.730 82.380 82.050 ;
        RECT 81.200 79.010 81.460 79.330 ;
        RECT 81.260 72.190 81.400 79.010 ;
        RECT 82.180 77.970 82.320 81.730 ;
        RECT 82.580 80.710 82.840 81.030 ;
        RECT 82.640 79.070 82.780 80.710 ;
        RECT 83.100 79.670 83.240 85.130 ;
        RECT 83.490 83.575 83.770 83.945 ;
        RECT 83.560 83.070 83.700 83.575 ;
        RECT 83.500 82.750 83.760 83.070 ;
        RECT 83.040 79.350 83.300 79.670 ;
        RECT 82.640 78.930 83.240 79.070 ;
        RECT 82.580 77.990 82.840 78.310 ;
        RECT 82.120 77.650 82.380 77.970 ;
        RECT 82.120 75.270 82.380 75.590 ;
        RECT 82.180 72.870 82.320 75.270 ;
        RECT 82.640 74.570 82.780 77.990 ;
        RECT 83.100 74.910 83.240 78.930 ;
        RECT 83.560 77.030 83.700 82.750 ;
        RECT 83.560 76.890 84.160 77.030 ;
        RECT 83.490 76.095 83.770 76.465 ;
        RECT 83.560 75.590 83.700 76.095 ;
        RECT 83.500 75.270 83.760 75.590 ;
        RECT 83.040 74.590 83.300 74.910 ;
        RECT 82.580 74.250 82.840 74.570 ;
        RECT 83.040 73.910 83.300 74.230 ;
        RECT 82.120 72.550 82.380 72.870 ;
        RECT 81.200 71.870 81.460 72.190 ;
        RECT 80.740 70.850 81.000 71.170 ;
        RECT 81.260 69.550 81.400 71.870 ;
        RECT 82.580 71.530 82.840 71.850 ;
        RECT 81.660 69.830 81.920 70.150 ;
        RECT 82.640 70.110 82.780 71.530 ;
        RECT 82.180 69.970 82.780 70.110 ;
        RECT 81.720 69.665 81.860 69.830 ;
        RECT 80.800 69.410 81.400 69.550 ;
        RECT 78.890 67.935 79.170 68.305 ;
        RECT 80.280 68.130 80.540 68.450 ;
        RECT 78.500 67.370 79.560 67.510 ;
        RECT 78.430 66.575 78.710 66.945 ;
        RECT 78.440 66.430 78.700 66.575 ;
        RECT 77.980 66.090 78.240 66.410 ;
        RECT 77.520 64.390 77.780 64.710 ;
        RECT 76.140 63.710 76.400 64.030 ;
        RECT 75.680 63.370 75.940 63.690 ;
        RECT 75.740 56.210 75.880 63.370 ;
        RECT 78.040 63.350 78.180 66.090 ;
        RECT 78.440 65.410 78.700 65.730 ;
        RECT 79.420 65.470 79.560 67.370 ;
        RECT 76.140 63.030 76.400 63.350 ;
        RECT 77.980 63.030 78.240 63.350 ;
        RECT 75.680 55.890 75.940 56.210 ;
        RECT 75.680 52.720 75.940 52.810 ;
        RECT 76.200 52.720 76.340 63.030 ;
        RECT 77.060 62.690 77.320 63.010 ;
        RECT 77.120 61.310 77.260 62.690 ;
        RECT 78.500 61.310 78.640 65.410 ;
        RECT 78.960 65.330 79.560 65.470 ;
        RECT 78.960 63.690 79.100 65.330 ;
        RECT 79.360 64.390 79.620 64.710 ;
        RECT 79.420 63.690 79.560 64.390 ;
        RECT 78.900 63.370 79.160 63.690 ;
        RECT 79.360 63.370 79.620 63.690 ;
        RECT 78.960 61.310 79.100 63.370 ;
        RECT 77.060 60.990 77.320 61.310 ;
        RECT 78.440 60.990 78.700 61.310 ;
        RECT 78.900 60.990 79.160 61.310 ;
        RECT 76.600 59.970 76.860 60.290 ;
        RECT 76.660 58.250 76.800 59.970 ;
        RECT 77.060 58.670 77.320 58.930 ;
        RECT 78.960 58.670 79.100 60.990 ;
        RECT 77.060 58.610 79.100 58.670 ;
        RECT 77.120 58.530 79.100 58.610 ;
        RECT 76.600 57.930 76.860 58.250 ;
        RECT 75.680 52.580 76.340 52.720 ;
        RECT 75.680 52.490 75.940 52.580 ;
        RECT 75.220 50.790 75.480 51.110 ;
        RECT 75.220 50.340 75.480 50.430 ;
        RECT 74.820 50.200 75.480 50.340 ;
        RECT 75.220 50.110 75.480 50.200 ;
        RECT 74.300 47.050 74.560 47.370 ;
        RECT 74.760 47.050 75.020 47.370 ;
        RECT 75.220 47.050 75.480 47.370 ;
        RECT 74.820 45.670 74.960 47.050 ;
        RECT 74.760 45.350 75.020 45.670 ;
        RECT 75.280 41.930 75.420 47.050 ;
        RECT 72.920 41.610 73.180 41.930 ;
        RECT 73.380 41.610 73.640 41.930 ;
        RECT 74.300 41.610 74.560 41.930 ;
        RECT 75.220 41.610 75.480 41.930 ;
        RECT 72.460 40.930 72.720 41.250 ;
        RECT 73.440 41.105 73.580 41.610 ;
        RECT 72.000 39.910 72.260 40.230 ;
        RECT 71.080 39.570 71.340 39.890 ;
        RECT 72.520 39.745 72.660 40.930 ;
        RECT 73.370 40.735 73.650 41.105 ;
        RECT 72.450 39.375 72.730 39.745 ;
        RECT 70.160 38.210 70.420 38.530 ;
        RECT 70.620 38.210 70.880 38.530 ;
        RECT 70.610 37.335 70.890 37.705 ;
        RECT 70.680 36.490 70.820 37.335 ;
        RECT 67.860 36.170 68.120 36.490 ;
        RECT 70.620 36.170 70.880 36.490 ;
        RECT 72.000 35.830 72.260 36.150 ;
        RECT 68.320 35.665 68.580 35.810 ;
        RECT 68.310 35.295 68.590 35.665 ;
        RECT 70.160 34.470 70.420 34.790 ;
        RECT 71.530 34.615 71.810 34.985 ;
        RECT 66.940 33.450 67.200 33.770 ;
        RECT 67.400 33.450 67.660 33.770 ;
        RECT 65.100 32.770 65.360 33.090 ;
        RECT 65.160 31.050 65.300 32.770 ;
        RECT 65.100 30.730 65.360 31.050 ;
        RECT 64.640 30.390 64.900 30.710 ;
        RECT 64.700 29.545 64.840 30.390 ;
        RECT 67.000 30.370 67.140 33.450 ;
        RECT 66.940 30.050 67.200 30.370 ;
        RECT 64.630 29.175 64.910 29.545 ;
        RECT 64.640 29.030 64.900 29.175 ;
        RECT 67.460 26.630 67.600 33.450 ;
        RECT 68.780 32.770 69.040 33.090 ;
        RECT 67.400 26.310 67.660 26.630 ;
        RECT 66.480 25.630 66.740 25.950 ;
        RECT 64.180 24.950 64.440 25.270 ;
        RECT 62.800 23.590 63.060 23.910 ;
        RECT 66.540 23.570 66.680 25.630 ;
        RECT 68.840 25.270 68.980 32.770 ;
        RECT 70.220 32.070 70.360 34.470 ;
        RECT 71.070 33.935 71.350 34.305 ;
        RECT 71.080 33.790 71.340 33.935 ;
        RECT 71.600 33.770 71.740 34.615 ;
        RECT 71.540 33.450 71.800 33.770 ;
        RECT 71.080 33.110 71.340 33.430 ;
        RECT 70.160 31.750 70.420 32.070 ;
        RECT 71.140 31.390 71.280 33.110 ;
        RECT 71.080 31.070 71.340 31.390 ;
        RECT 71.080 30.050 71.340 30.370 ;
        RECT 71.140 29.010 71.280 30.050 ;
        RECT 71.080 28.690 71.340 29.010 ;
        RECT 72.060 25.610 72.200 35.830 ;
        RECT 73.440 34.450 73.580 40.735 ;
        RECT 74.360 40.230 74.500 41.610 ;
        RECT 74.760 40.930 75.020 41.250 ;
        RECT 74.300 39.910 74.560 40.230 ;
        RECT 74.820 39.630 74.960 40.930 ;
        RECT 74.360 39.550 74.960 39.630 ;
        RECT 74.300 39.490 74.960 39.550 ;
        RECT 74.300 39.230 74.560 39.490 ;
        RECT 75.740 39.460 75.880 52.490 ;
        RECT 76.140 51.810 76.400 52.130 ;
        RECT 76.200 50.430 76.340 51.810 ;
        RECT 76.660 50.430 76.800 57.930 ;
        RECT 77.520 55.890 77.780 56.210 ;
        RECT 76.140 50.110 76.400 50.430 ;
        RECT 76.600 50.110 76.860 50.430 ;
        RECT 76.660 47.370 76.800 50.110 ;
        RECT 76.600 47.050 76.860 47.370 ;
        RECT 76.600 43.650 76.860 43.970 ;
        RECT 76.660 41.930 76.800 43.650 ;
        RECT 77.580 41.930 77.720 55.890 ;
        RECT 78.960 55.270 79.100 58.530 ;
        RECT 79.420 56.550 79.560 63.370 ;
        RECT 79.360 56.230 79.620 56.550 ;
        RECT 80.340 55.870 80.480 68.130 ;
        RECT 80.800 67.090 80.940 69.410 ;
        RECT 81.650 69.295 81.930 69.665 ;
        RECT 81.200 68.470 81.460 68.790 ;
        RECT 80.740 66.770 81.000 67.090 ;
        RECT 81.260 66.750 81.400 68.470 ;
        RECT 82.180 67.430 82.320 69.970 ;
        RECT 83.100 69.470 83.240 73.910 ;
        RECT 84.020 70.110 84.160 76.890 ;
        RECT 84.480 75.590 84.620 85.130 ;
        RECT 84.880 82.750 85.140 83.070 ;
        RECT 86.260 82.750 86.520 83.070 ;
        RECT 86.720 82.750 86.980 83.070 ;
        RECT 84.940 81.030 85.080 82.750 ;
        RECT 86.320 82.390 86.460 82.750 ;
        RECT 86.260 82.070 86.520 82.390 ;
        RECT 84.880 80.710 85.140 81.030 ;
        RECT 84.880 79.690 85.140 80.010 ;
        RECT 84.940 76.610 85.080 79.690 ;
        RECT 84.880 76.290 85.140 76.610 ;
        RECT 84.420 75.270 84.680 75.590 ;
        RECT 84.940 72.190 85.080 76.290 ;
        RECT 85.340 73.570 85.600 73.890 ;
        RECT 85.400 72.190 85.540 73.570 ;
        RECT 84.880 71.870 85.140 72.190 ;
        RECT 85.340 71.870 85.600 72.190 ;
        RECT 85.800 71.870 86.060 72.190 ;
        RECT 85.860 71.025 86.000 71.870 ;
        RECT 85.790 70.655 86.070 71.025 ;
        RECT 86.320 70.230 86.460 82.070 ;
        RECT 86.780 79.330 86.920 82.750 ;
        RECT 87.240 80.690 87.380 85.130 ;
        RECT 87.700 83.410 87.840 96.350 ;
        RECT 88.160 96.330 88.300 96.495 ;
        RECT 88.100 96.010 88.360 96.330 ;
        RECT 88.100 95.330 88.360 95.650 ;
        RECT 88.160 90.890 88.300 95.330 ;
        RECT 88.620 93.610 88.760 107.375 ;
        RECT 95.400 100.035 95.645 217.375 ;
        RECT 96.145 100.700 96.445 216.925 ;
        RECT 96.825 101.360 97.110 217.555 ;
        RECT 97.505 101.930 97.770 216.935 ;
        RECT 98.170 102.480 98.440 217.670 ;
        RECT 99.205 217.340 99.465 217.660 ;
        RECT 98.755 216.765 99.015 217.085 ;
        RECT 98.780 102.970 98.990 216.765 ;
        RECT 99.225 103.390 99.440 217.340 ;
        RECT 99.700 216.790 99.960 217.110 ;
        RECT 99.710 103.900 99.945 216.790 ;
        RECT 110.010 206.150 110.150 218.060 ;
        RECT 111.010 206.600 111.150 218.690 ;
        RECT 110.920 206.340 111.240 206.600 ;
        RECT 109.920 205.890 110.240 206.150 ;
        RECT 111.420 206.120 111.560 219.040 ;
        RECT 111.330 205.860 111.650 206.120 ;
        RECT 101.480 205.335 105.480 205.405 ;
        RECT 111.810 205.335 111.950 219.350 ;
        RECT 121.210 218.215 121.530 218.275 ;
        RECT 125.435 218.215 125.805 218.285 ;
        RECT 121.210 218.075 125.805 218.215 ;
        RECT 121.210 218.015 121.530 218.075 ;
        RECT 125.435 218.005 125.805 218.075 ;
        RECT 128.010 218.215 128.330 218.275 ;
        RECT 132.235 218.215 132.605 218.285 ;
        RECT 139.035 218.275 139.405 218.285 ;
        RECT 128.010 218.075 132.605 218.215 ;
        RECT 128.010 218.015 128.330 218.075 ;
        RECT 132.235 218.005 132.605 218.075 ;
        RECT 138.890 218.015 139.405 218.275 ;
        RECT 139.035 218.005 139.405 218.015 ;
        RECT 116.450 217.755 116.770 217.815 ;
        RECT 119.850 217.755 120.170 217.815 ;
        RECT 121.550 217.755 121.870 217.815 ;
        RECT 116.450 217.615 121.870 217.755 ;
        RECT 116.450 217.555 116.770 217.615 ;
        RECT 119.850 217.555 120.170 217.615 ;
        RECT 121.550 217.555 121.870 217.615 ;
        RECT 124.610 217.755 124.930 217.815 ;
        RECT 126.650 217.755 126.970 217.815 ;
        RECT 124.610 217.615 126.970 217.755 ;
        RECT 124.610 217.555 124.930 217.615 ;
        RECT 126.650 217.555 126.970 217.615 ;
        RECT 127.330 217.755 127.650 217.815 ;
        RECT 130.050 217.755 130.370 217.815 ;
        RECT 131.750 217.755 132.070 217.815 ;
        RECT 127.330 217.615 132.070 217.755 ;
        RECT 127.330 217.555 127.650 217.615 ;
        RECT 130.050 217.555 130.370 217.615 ;
        RECT 131.750 217.555 132.070 217.615 ;
        RECT 133.110 217.755 133.430 217.815 ;
        RECT 134.470 217.755 134.790 217.815 ;
        RECT 133.110 217.615 134.790 217.755 ;
        RECT 133.110 217.555 133.430 217.615 ;
        RECT 134.470 217.555 134.790 217.615 ;
        RECT 138.890 215.915 139.210 215.975 ;
        RECT 140.250 215.915 140.570 215.975 ;
        RECT 138.890 215.775 140.570 215.915 ;
        RECT 138.890 215.715 139.210 215.775 ;
        RECT 140.250 215.715 140.570 215.775 ;
        RECT 123.930 215.455 124.250 215.515 ;
        RECT 126.310 215.455 126.630 215.515 ;
        RECT 123.930 215.315 126.630 215.455 ;
        RECT 123.930 215.255 124.250 215.315 ;
        RECT 126.310 215.255 126.630 215.315 ;
        RECT 135.490 215.455 135.810 215.515 ;
        RECT 137.530 215.455 137.850 215.515 ;
        RECT 135.490 215.315 137.850 215.455 ;
        RECT 135.490 215.255 135.810 215.315 ;
        RECT 137.530 215.255 137.850 215.315 ;
        RECT 117.130 214.995 117.450 215.055 ;
        RECT 118.490 214.995 118.810 215.055 ;
        RECT 117.130 214.855 118.810 214.995 ;
        RECT 117.130 214.795 117.450 214.855 ;
        RECT 118.490 214.795 118.810 214.855 ;
        RECT 144.330 213.615 144.650 213.675 ;
        RECT 146.030 213.615 146.350 213.675 ;
        RECT 144.330 213.475 146.350 213.615 ;
        RECT 144.330 213.415 144.650 213.475 ;
        RECT 146.030 213.415 146.350 213.475 ;
        RECT 117.130 213.155 117.450 213.215 ;
        RECT 120.870 213.155 121.190 213.215 ;
        RECT 117.130 213.015 121.190 213.155 ;
        RECT 117.130 212.955 117.450 213.015 ;
        RECT 120.870 212.955 121.190 213.015 ;
        RECT 130.730 213.155 131.050 213.215 ;
        RECT 134.470 213.155 134.790 213.215 ;
        RECT 130.730 213.015 134.790 213.155 ;
        RECT 130.730 212.955 131.050 213.015 ;
        RECT 134.470 212.955 134.790 213.015 ;
        RECT 117.130 212.695 117.450 212.755 ;
        RECT 121.210 212.695 121.530 212.755 ;
        RECT 126.990 212.695 127.310 212.755 ;
        RECT 117.130 212.555 127.310 212.695 ;
        RECT 117.130 212.495 117.450 212.555 ;
        RECT 121.210 212.495 121.530 212.555 ;
        RECT 126.990 212.495 127.310 212.555 ;
        RECT 128.010 212.695 128.330 212.755 ;
        RECT 129.030 212.695 129.350 212.755 ;
        RECT 128.010 212.555 129.350 212.695 ;
        RECT 128.010 212.495 128.330 212.555 ;
        RECT 129.030 212.495 129.350 212.555 ;
        RECT 126.990 212.235 127.310 212.295 ;
        RECT 134.810 212.235 135.130 212.295 ;
        RECT 137.870 212.235 138.190 212.295 ;
        RECT 126.990 212.095 138.190 212.235 ;
        RECT 126.990 212.035 127.310 212.095 ;
        RECT 134.810 212.035 135.130 212.095 ;
        RECT 137.870 212.035 138.190 212.095 ;
        RECT 119.170 210.855 119.490 210.915 ;
        RECT 124.270 210.855 124.590 210.915 ;
        RECT 119.170 210.715 124.590 210.855 ;
        RECT 119.170 210.655 119.490 210.715 ;
        RECT 124.270 210.655 124.590 210.715 ;
        RECT 132.770 210.855 133.090 210.915 ;
        RECT 135.150 210.855 135.470 210.915 ;
        RECT 132.770 210.715 135.470 210.855 ;
        RECT 132.770 210.655 133.090 210.715 ;
        RECT 135.150 210.655 135.470 210.715 ;
        RECT 138.210 210.855 138.530 210.915 ;
        RECT 139.910 210.855 140.230 210.915 ;
        RECT 138.210 210.715 140.230 210.855 ;
        RECT 138.210 210.655 138.530 210.715 ;
        RECT 139.910 210.655 140.230 210.715 ;
        RECT 117.130 210.395 117.450 210.455 ;
        RECT 121.550 210.395 121.870 210.455 ;
        RECT 117.130 210.255 121.870 210.395 ;
        RECT 117.130 210.195 117.450 210.255 ;
        RECT 121.550 210.195 121.870 210.255 ;
        RECT 138.890 210.395 139.210 210.455 ;
        RECT 139.910 210.395 140.230 210.455 ;
        RECT 138.890 210.255 140.230 210.395 ;
        RECT 138.890 210.195 139.210 210.255 ;
        RECT 139.910 210.195 140.230 210.255 ;
        RECT 121.890 209.935 122.210 209.995 ;
        RECT 125.290 209.935 125.610 209.995 ;
        RECT 129.710 209.935 130.030 209.995 ;
        RECT 121.890 209.795 130.030 209.935 ;
        RECT 121.890 209.735 122.210 209.795 ;
        RECT 125.290 209.735 125.610 209.795 ;
        RECT 129.710 209.735 130.030 209.795 ;
        RECT 144.330 209.015 144.650 209.075 ;
        RECT 146.030 209.015 146.350 209.075 ;
        RECT 144.330 208.875 146.350 209.015 ;
        RECT 144.330 208.815 144.650 208.875 ;
        RECT 146.030 208.815 146.350 208.875 ;
        RECT 143.795 208.555 144.165 208.625 ;
        RECT 146.030 208.555 146.350 208.615 ;
        RECT 143.795 208.415 146.350 208.555 ;
        RECT 143.795 208.345 144.165 208.415 ;
        RECT 146.030 208.355 146.350 208.415 ;
        RECT 113.390 208.095 113.710 208.155 ;
        RECT 117.130 208.095 117.450 208.155 ;
        RECT 113.390 207.955 117.450 208.095 ;
        RECT 113.390 207.895 113.710 207.955 ;
        RECT 117.130 207.895 117.450 207.955 ;
        RECT 135.150 208.095 135.470 208.155 ;
        RECT 138.890 208.095 139.210 208.155 ;
        RECT 140.590 208.095 140.910 208.155 ;
        RECT 142.630 208.095 142.950 208.155 ;
        RECT 135.150 207.955 142.950 208.095 ;
        RECT 135.150 207.895 135.470 207.955 ;
        RECT 138.890 207.895 139.210 207.955 ;
        RECT 140.590 207.895 140.910 207.955 ;
        RECT 142.630 207.895 142.950 207.955 ;
        RECT 133.110 207.175 133.430 207.235 ;
        RECT 142.435 207.175 142.805 207.245 ;
        RECT 133.110 207.035 142.805 207.175 ;
        RECT 133.110 206.975 133.430 207.035 ;
        RECT 142.435 206.965 142.805 207.035 ;
        RECT 143.990 206.715 144.310 206.775 ;
        RECT 145.350 206.715 145.670 206.775 ;
        RECT 143.990 206.575 145.670 206.715 ;
        RECT 143.990 206.515 144.310 206.575 ;
        RECT 145.350 206.515 145.670 206.575 ;
        RECT 116.110 206.255 116.430 206.315 ;
        RECT 121.550 206.255 121.870 206.315 ;
        RECT 127.670 206.255 127.990 206.315 ;
        RECT 116.110 206.115 127.990 206.255 ;
        RECT 116.110 206.055 116.430 206.115 ;
        RECT 121.550 206.055 121.870 206.115 ;
        RECT 127.670 206.055 127.990 206.115 ;
        RECT 135.490 205.795 135.810 205.855 ;
        RECT 138.890 205.795 139.210 205.855 ;
        RECT 135.490 205.655 139.210 205.795 ;
        RECT 135.490 205.595 135.810 205.655 ;
        RECT 138.890 205.595 139.210 205.655 ;
        RECT 141.610 205.795 141.930 205.855 ;
        RECT 143.650 205.795 143.970 205.855 ;
        RECT 141.610 205.655 143.970 205.795 ;
        RECT 141.610 205.595 141.930 205.655 ;
        RECT 143.650 205.595 143.970 205.655 ;
        RECT 112.710 205.335 113.030 205.395 ;
        RECT 101.480 205.195 113.030 205.335 ;
        RECT 101.480 205.125 105.480 205.195 ;
        RECT 112.710 205.135 113.030 205.195 ;
        RECT 147.050 205.335 147.370 205.395 ;
        RECT 149.680 205.335 150.000 205.430 ;
        RECT 155.245 205.335 159.245 205.405 ;
        RECT 147.050 205.195 159.245 205.335 ;
        RECT 147.050 205.135 147.370 205.195 ;
        RECT 149.680 205.100 150.000 205.195 ;
        RECT 155.245 205.125 159.245 205.195 ;
        RECT 123.930 204.875 124.250 204.935 ;
        RECT 126.650 204.875 126.970 204.935 ;
        RECT 123.930 204.735 126.970 204.875 ;
        RECT 123.930 204.675 124.250 204.735 ;
        RECT 126.650 204.675 126.970 204.735 ;
        RECT 127.670 204.875 127.990 204.935 ;
        RECT 130.730 204.875 131.050 204.935 ;
        RECT 136.170 204.875 136.490 204.935 ;
        RECT 138.890 204.875 139.210 204.935 ;
        RECT 127.670 204.735 139.210 204.875 ;
        RECT 127.670 204.675 127.990 204.735 ;
        RECT 130.730 204.675 131.050 204.735 ;
        RECT 136.170 204.675 136.490 204.735 ;
        RECT 138.890 204.675 139.210 204.735 ;
        RECT 128.010 204.415 128.330 204.475 ;
        RECT 129.710 204.415 130.030 204.475 ;
        RECT 128.010 204.275 130.030 204.415 ;
        RECT 128.010 204.215 128.330 204.275 ;
        RECT 129.710 204.215 130.030 204.275 ;
        RECT 130.730 204.415 131.050 204.475 ;
        RECT 143.795 204.415 144.165 204.485 ;
        RECT 130.730 204.275 144.165 204.415 ;
        RECT 130.730 204.215 131.050 204.275 ;
        RECT 143.795 204.205 144.165 204.275 ;
        RECT 113.390 202.835 113.710 203.095 ;
        RECT 111.360 202.575 111.620 202.665 ;
        RECT 112.710 202.575 113.030 202.635 ;
        RECT 107.190 202.435 113.030 202.575 ;
        RECT 101.480 202.115 105.480 202.185 ;
        RECT 107.190 202.115 107.330 202.435 ;
        RECT 111.360 202.345 111.620 202.435 ;
        RECT 112.710 202.375 113.030 202.435 ;
        RECT 101.480 201.975 107.330 202.115 ;
        RECT 101.480 201.905 105.480 201.975 ;
        RECT 113.480 201.655 113.620 202.835 ;
        RECT 114.895 202.205 115.265 203.745 ;
        RECT 120.335 202.205 120.705 203.745 ;
        RECT 125.775 202.205 126.145 203.745 ;
        RECT 131.215 202.205 131.585 203.745 ;
        RECT 136.655 202.205 137.025 203.745 ;
        RECT 142.095 202.205 142.465 203.745 ;
        RECT 147.535 202.205 147.905 203.745 ;
        RECT 155.245 202.115 159.245 202.185 ;
        RECT 148.670 201.975 159.245 202.115 ;
        RECT 117.130 201.655 117.450 201.715 ;
        RECT 120.870 201.655 121.190 201.715 ;
        RECT 113.480 201.515 116.850 201.655 ;
        RECT 116.710 200.795 116.850 201.515 ;
        RECT 117.130 201.515 121.190 201.655 ;
        RECT 117.130 201.455 117.450 201.515 ;
        RECT 120.870 201.455 121.190 201.515 ;
        RECT 129.710 201.655 130.030 201.715 ;
        RECT 139.910 201.655 140.230 201.715 ;
        RECT 129.710 201.515 140.230 201.655 ;
        RECT 129.710 201.455 130.030 201.515 ;
        RECT 139.910 201.455 140.230 201.515 ;
        RECT 140.590 201.655 140.910 201.715 ;
        RECT 145.350 201.655 145.670 201.715 ;
        RECT 140.590 201.515 145.670 201.655 ;
        RECT 140.590 201.455 140.910 201.515 ;
        RECT 145.350 201.455 145.670 201.515 ;
        RECT 118.830 201.195 119.150 201.255 ;
        RECT 131.750 201.195 132.070 201.255 ;
        RECT 138.210 201.195 138.530 201.255 ;
        RECT 118.830 201.055 138.530 201.195 ;
        RECT 118.830 200.995 119.150 201.055 ;
        RECT 131.750 200.995 132.070 201.055 ;
        RECT 138.210 200.995 138.530 201.055 ;
        RECT 138.890 201.195 139.210 201.255 ;
        RECT 140.590 201.195 140.910 201.255 ;
        RECT 138.890 201.055 140.910 201.195 ;
        RECT 138.890 200.995 139.210 201.055 ;
        RECT 140.590 200.995 140.910 201.055 ;
        RECT 142.970 201.195 143.290 201.255 ;
        RECT 148.110 201.195 148.440 201.290 ;
        RECT 148.670 201.195 148.810 201.975 ;
        RECT 155.245 201.905 159.245 201.975 ;
        RECT 142.970 201.055 148.810 201.195 ;
        RECT 142.970 200.995 143.290 201.055 ;
        RECT 148.110 200.960 148.440 201.055 ;
        RECT 113.050 200.735 113.370 200.795 ;
        RECT 115.430 200.735 115.750 200.795 ;
        RECT 113.050 200.595 115.750 200.735 ;
        RECT 116.710 200.735 117.110 200.795 ;
        RECT 119.850 200.735 120.170 200.795 ;
        RECT 121.890 200.735 122.210 200.795 ;
        RECT 123.590 200.735 123.910 200.795 ;
        RECT 116.710 200.595 123.910 200.735 ;
        RECT 113.050 200.535 113.370 200.595 ;
        RECT 115.430 200.535 115.750 200.595 ;
        RECT 116.790 200.535 117.110 200.595 ;
        RECT 119.850 200.535 120.170 200.595 ;
        RECT 121.890 200.535 122.210 200.595 ;
        RECT 123.590 200.535 123.910 200.595 ;
        RECT 129.710 200.735 130.030 200.795 ;
        RECT 132.430 200.735 132.750 200.795 ;
        RECT 137.190 200.735 137.510 200.795 ;
        RECT 129.710 200.595 132.750 200.735 ;
        RECT 129.710 200.535 130.030 200.595 ;
        RECT 132.430 200.535 132.750 200.595 ;
        RECT 133.030 200.595 137.510 200.735 ;
        RECT 101.480 198.895 105.480 198.965 ;
        RECT 112.175 198.905 112.545 200.445 ;
        RECT 117.615 198.905 117.985 200.445 ;
        RECT 123.055 198.905 123.425 200.445 ;
        RECT 128.495 198.905 128.865 200.445 ;
        RECT 130.390 200.275 130.710 200.335 ;
        RECT 133.030 200.275 133.170 200.595 ;
        RECT 137.190 200.535 137.510 200.595 ;
        RECT 141.610 200.735 141.930 200.795 ;
        RECT 146.710 200.735 147.030 200.795 ;
        RECT 141.610 200.595 147.030 200.735 ;
        RECT 141.610 200.535 141.930 200.595 ;
        RECT 146.710 200.535 147.030 200.595 ;
        RECT 130.390 200.135 133.170 200.275 ;
        RECT 130.390 200.075 130.710 200.135 ;
        RECT 133.935 198.905 134.305 200.445 ;
        RECT 139.375 198.905 139.745 200.445 ;
        RECT 140.590 200.275 140.910 200.335 ;
        RECT 143.310 200.275 143.630 200.335 ;
        RECT 140.590 200.135 143.630 200.275 ;
        RECT 140.590 200.075 140.910 200.135 ;
        RECT 143.310 200.075 143.630 200.135 ;
        RECT 144.815 198.905 145.185 200.445 ;
        RECT 147.050 198.895 147.370 198.955 ;
        RECT 148.660 198.895 148.920 198.985 ;
        RECT 155.245 198.895 159.245 198.965 ;
        RECT 101.480 198.755 107.330 198.895 ;
        RECT 101.480 198.685 105.480 198.755 ;
        RECT 107.190 198.435 107.330 198.755 ;
        RECT 147.050 198.755 159.245 198.895 ;
        RECT 147.050 198.695 147.370 198.755 ;
        RECT 148.660 198.665 148.920 198.755 ;
        RECT 155.245 198.685 159.245 198.755 ;
        RECT 111.410 198.435 111.740 198.530 ;
        RECT 112.710 198.435 113.030 198.495 ;
        RECT 107.190 198.295 113.030 198.435 ;
        RECT 111.410 198.200 111.740 198.295 ;
        RECT 112.710 198.235 113.030 198.295 ;
        RECT 126.990 198.435 127.310 198.495 ;
        RECT 134.470 198.435 134.790 198.495 ;
        RECT 136.170 198.435 136.490 198.495 ;
        RECT 140.590 198.435 140.910 198.495 ;
        RECT 126.990 198.295 135.890 198.435 ;
        RECT 126.990 198.235 127.310 198.295 ;
        RECT 134.470 198.235 134.790 198.295 ;
        RECT 114.410 197.975 114.730 198.035 ;
        RECT 123.590 197.975 123.910 198.035 ;
        RECT 126.990 197.975 127.310 198.035 ;
        RECT 114.410 197.835 127.310 197.975 ;
        RECT 114.410 197.775 114.730 197.835 ;
        RECT 123.590 197.775 123.910 197.835 ;
        RECT 126.990 197.775 127.310 197.835 ;
        RECT 133.450 197.975 133.770 198.035 ;
        RECT 134.810 197.975 135.130 198.035 ;
        RECT 133.450 197.835 135.130 197.975 ;
        RECT 135.750 197.975 135.890 198.295 ;
        RECT 136.170 198.295 140.910 198.435 ;
        RECT 136.170 198.235 136.490 198.295 ;
        RECT 140.590 198.235 140.910 198.295 ;
        RECT 144.330 198.435 144.650 198.495 ;
        RECT 146.030 198.435 146.350 198.495 ;
        RECT 144.330 198.295 146.350 198.435 ;
        RECT 144.330 198.235 144.650 198.295 ;
        RECT 146.030 198.235 146.350 198.295 ;
        RECT 140.590 197.975 140.910 198.035 ;
        RECT 135.750 197.835 140.910 197.975 ;
        RECT 133.450 197.775 133.770 197.835 ;
        RECT 134.810 197.775 135.130 197.835 ;
        RECT 140.590 197.775 140.910 197.835 ;
        RECT 143.990 197.975 144.310 198.035 ;
        RECT 145.350 197.975 145.670 198.035 ;
        RECT 143.990 197.835 145.670 197.975 ;
        RECT 143.990 197.775 144.310 197.835 ;
        RECT 145.350 197.775 145.670 197.835 ;
        RECT 124.610 197.515 124.930 197.575 ;
        RECT 124.610 197.315 125.010 197.515 ;
        RECT 128.010 197.315 128.330 197.575 ;
        RECT 135.150 197.515 135.470 197.575 ;
        RECT 137.870 197.515 138.190 197.575 ;
        RECT 135.150 197.375 138.190 197.515 ;
        RECT 135.150 197.315 135.470 197.375 ;
        RECT 137.870 197.315 138.190 197.375 ;
        RECT 140.930 197.515 141.250 197.575 ;
        RECT 142.630 197.515 142.950 197.575 ;
        RECT 140.930 197.375 142.950 197.515 ;
        RECT 140.930 197.315 141.250 197.375 ;
        RECT 142.630 197.315 142.950 197.375 ;
        RECT 124.870 197.055 125.010 197.315 ;
        RECT 128.100 197.055 128.240 197.315 ;
        RECT 130.050 197.055 130.370 197.115 ;
        RECT 135.830 197.055 136.150 197.115 ;
        RECT 124.870 196.915 136.150 197.055 ;
        RECT 130.050 196.855 130.370 196.915 ;
        RECT 135.830 196.855 136.150 196.915 ;
        RECT 140.590 197.055 140.910 197.115 ;
        RECT 143.650 197.055 143.970 197.115 ;
        RECT 140.590 196.915 143.970 197.055 ;
        RECT 140.590 196.855 140.910 196.915 ;
        RECT 143.650 196.855 143.970 196.915 ;
        RECT 124.950 196.595 125.270 196.655 ;
        RECT 134.810 196.595 135.130 196.655 ;
        RECT 124.950 196.455 135.130 196.595 ;
        RECT 124.950 196.395 125.270 196.455 ;
        RECT 134.810 196.395 135.130 196.455 ;
        RECT 117.130 196.135 117.450 196.195 ;
        RECT 122.230 196.135 122.550 196.195 ;
        RECT 126.650 196.135 126.970 196.195 ;
        RECT 117.130 195.995 126.970 196.135 ;
        RECT 117.130 195.935 117.450 195.995 ;
        RECT 122.230 195.935 122.550 195.995 ;
        RECT 126.650 195.935 126.970 195.995 ;
        RECT 130.390 196.135 130.710 196.195 ;
        RECT 131.750 196.135 132.070 196.195 ;
        RECT 138.550 196.135 138.870 196.195 ;
        RECT 143.310 196.135 143.630 196.195 ;
        RECT 130.390 195.995 143.630 196.135 ;
        RECT 130.390 195.935 130.710 195.995 ;
        RECT 131.750 195.935 132.070 195.995 ;
        RECT 138.550 195.935 138.870 195.995 ;
        RECT 143.310 195.935 143.630 195.995 ;
        RECT 133.450 195.675 133.770 195.735 ;
        RECT 137.530 195.675 137.850 195.735 ;
        RECT 140.250 195.675 140.570 195.735 ;
        RECT 141.610 195.675 141.930 195.735 ;
        RECT 143.650 195.675 143.970 195.735 ;
        RECT 133.450 195.535 140.570 195.675 ;
        RECT 133.450 195.475 133.770 195.535 ;
        RECT 137.530 195.475 137.850 195.535 ;
        RECT 140.250 195.475 140.570 195.535 ;
        RECT 141.190 195.535 143.970 195.675 ;
        RECT 116.110 195.215 116.430 195.275 ;
        RECT 121.890 195.215 122.210 195.275 ;
        RECT 125.290 195.215 125.610 195.275 ;
        RECT 141.190 195.215 141.330 195.535 ;
        RECT 141.610 195.475 141.930 195.535 ;
        RECT 143.650 195.475 143.970 195.535 ;
        RECT 146.030 195.675 146.350 195.735 ;
        RECT 148.050 195.675 148.470 195.800 ;
        RECT 155.245 195.675 159.245 195.745 ;
        RECT 146.030 195.535 159.245 195.675 ;
        RECT 146.030 195.475 146.350 195.535 ;
        RECT 148.050 195.410 148.470 195.535 ;
        RECT 155.245 195.465 159.245 195.535 ;
        RECT 116.110 195.075 141.330 195.215 ;
        RECT 116.110 195.015 116.430 195.075 ;
        RECT 121.890 195.015 122.210 195.075 ;
        RECT 125.290 195.015 125.610 195.075 ;
        RECT 113.390 194.755 113.710 194.815 ;
        RECT 114.070 194.755 114.390 194.815 ;
        RECT 116.110 194.755 116.430 194.815 ;
        RECT 113.390 194.615 116.430 194.755 ;
        RECT 113.390 194.555 113.710 194.615 ;
        RECT 114.070 194.555 114.390 194.615 ;
        RECT 116.110 194.555 116.430 194.615 ;
        RECT 140.590 194.755 140.910 194.815 ;
        RECT 142.630 194.755 142.950 194.815 ;
        RECT 140.590 194.615 142.950 194.755 ;
        RECT 140.590 194.555 140.910 194.615 ;
        RECT 142.630 194.555 142.950 194.615 ;
        RECT 120.870 194.295 121.190 194.355 ;
        RECT 121.550 194.295 121.870 194.355 ;
        RECT 129.030 194.295 129.350 194.355 ;
        RECT 120.870 194.155 129.350 194.295 ;
        RECT 120.870 194.095 121.190 194.155 ;
        RECT 121.550 194.095 121.870 194.155 ;
        RECT 129.030 194.095 129.350 194.155 ;
        RECT 115.235 193.835 115.605 193.905 ;
        RECT 118.830 193.835 119.150 193.895 ;
        RECT 115.235 193.695 119.150 193.835 ;
        RECT 115.235 193.625 115.605 193.695 ;
        RECT 118.830 193.635 119.150 193.695 ;
        RECT 127.330 193.835 127.650 193.895 ;
        RECT 130.730 193.835 131.050 193.895 ;
        RECT 137.190 193.835 137.510 193.895 ;
        RECT 127.330 193.695 137.510 193.835 ;
        RECT 127.330 193.635 127.650 193.695 ;
        RECT 130.730 193.635 131.050 193.695 ;
        RECT 137.190 193.635 137.510 193.695 ;
        RECT 143.650 193.835 143.970 193.895 ;
        RECT 146.710 193.835 147.030 193.895 ;
        RECT 143.650 193.695 147.030 193.835 ;
        RECT 143.650 193.635 143.970 193.695 ;
        RECT 146.710 193.635 147.030 193.695 ;
        RECT 132.770 192.915 133.090 192.975 ;
        RECT 134.470 192.915 134.790 192.975 ;
        RECT 132.770 192.775 134.790 192.915 ;
        RECT 132.770 192.715 133.090 192.775 ;
        RECT 134.470 192.715 134.790 192.775 ;
        RECT 101.480 192.455 105.480 192.525 ;
        RECT 109.920 192.455 110.240 192.515 ;
        RECT 112.710 192.455 113.030 192.515 ;
        RECT 101.480 192.315 113.030 192.455 ;
        RECT 101.480 192.245 105.480 192.315 ;
        RECT 109.920 192.255 110.240 192.315 ;
        RECT 112.710 192.255 113.030 192.315 ;
        RECT 118.830 192.455 119.150 192.515 ;
        RECT 125.435 192.455 125.805 192.525 ;
        RECT 118.830 192.315 125.805 192.455 ;
        RECT 118.830 192.255 119.150 192.315 ;
        RECT 125.435 192.245 125.805 192.315 ;
        RECT 147.050 192.455 147.370 192.515 ;
        RECT 148.570 192.455 148.900 192.550 ;
        RECT 155.245 192.455 159.245 192.525 ;
        RECT 147.050 192.315 159.245 192.455 ;
        RECT 147.050 192.255 147.370 192.315 ;
        RECT 148.570 192.220 148.900 192.315 ;
        RECT 155.245 192.245 159.245 192.315 ;
        RECT 113.390 191.995 113.710 192.055 ;
        RECT 120.870 191.995 121.190 192.055 ;
        RECT 124.270 191.995 124.590 192.055 ;
        RECT 113.390 191.855 124.590 191.995 ;
        RECT 113.390 191.795 113.710 191.855 ;
        RECT 120.870 191.795 121.190 191.855 ;
        RECT 124.270 191.795 124.590 191.855 ;
        RECT 132.770 191.995 133.090 192.055 ;
        RECT 138.210 191.995 138.530 192.055 ;
        RECT 145.350 191.995 145.670 192.055 ;
        RECT 132.770 191.855 145.670 191.995 ;
        RECT 132.770 191.795 133.090 191.855 ;
        RECT 138.210 191.795 138.530 191.855 ;
        RECT 145.350 191.795 145.670 191.855 ;
        RECT 127.330 191.535 127.650 191.595 ;
        RECT 129.030 191.535 129.350 191.595 ;
        RECT 127.330 191.395 129.350 191.535 ;
        RECT 127.330 191.335 127.650 191.395 ;
        RECT 129.030 191.335 129.350 191.395 ;
        RECT 138.550 191.535 138.870 191.595 ;
        RECT 138.550 191.395 143.880 191.535 ;
        RECT 138.550 191.335 138.870 191.395 ;
        RECT 143.740 191.145 143.880 191.395 ;
        RECT 118.635 191.135 119.005 191.145 ;
        RECT 143.740 191.135 144.165 191.145 ;
        RECT 118.635 190.875 119.150 191.135 ;
        RECT 122.570 191.075 122.890 191.135 ;
        RECT 123.590 191.075 123.910 191.135 ;
        RECT 122.570 190.935 123.910 191.075 ;
        RECT 122.570 190.875 122.890 190.935 ;
        RECT 123.590 190.875 123.910 190.935 ;
        RECT 129.710 191.075 130.030 191.135 ;
        RECT 135.150 191.075 135.470 191.135 ;
        RECT 137.530 191.075 137.850 191.135 ;
        RECT 138.550 191.075 138.870 191.135 ;
        RECT 129.710 190.935 130.450 191.075 ;
        RECT 129.710 190.875 130.030 190.935 ;
        RECT 118.635 190.865 119.005 190.875 ;
        RECT 128.835 190.155 129.205 190.225 ;
        RECT 129.710 190.155 130.030 190.215 ;
        RECT 128.835 190.015 130.030 190.155 ;
        RECT 130.310 190.155 130.450 190.935 ;
        RECT 135.150 190.935 138.870 191.075 ;
        RECT 135.150 190.875 135.470 190.935 ;
        RECT 137.530 190.875 137.850 190.935 ;
        RECT 138.550 190.875 138.870 190.935 ;
        RECT 143.650 190.875 144.165 191.135 ;
        RECT 143.795 190.865 144.165 190.875 ;
        RECT 141.610 190.615 141.930 190.675 ;
        RECT 142.970 190.615 143.290 190.675 ;
        RECT 146.030 190.615 146.350 190.675 ;
        RECT 141.610 190.475 146.350 190.615 ;
        RECT 141.610 190.415 141.930 190.475 ;
        RECT 142.970 190.415 143.290 190.475 ;
        RECT 146.030 190.415 146.350 190.475 ;
        RECT 135.830 190.155 136.150 190.215 ;
        RECT 130.310 190.015 136.150 190.155 ;
        RECT 128.835 189.945 129.205 190.015 ;
        RECT 129.710 189.955 130.030 190.015 ;
        RECT 135.830 189.955 136.150 190.015 ;
        RECT 113.730 189.695 114.050 189.755 ;
        RECT 116.110 189.695 116.430 189.755 ;
        RECT 118.150 189.695 118.470 189.755 ;
        RECT 113.730 189.555 118.470 189.695 ;
        RECT 113.730 189.495 114.050 189.555 ;
        RECT 116.110 189.495 116.430 189.555 ;
        RECT 118.150 189.495 118.470 189.555 ;
        RECT 124.610 189.695 124.930 189.755 ;
        RECT 127.670 189.695 127.990 189.755 ;
        RECT 129.370 189.695 129.690 189.755 ;
        RECT 131.750 189.695 132.070 189.755 ;
        RECT 124.610 189.555 132.070 189.695 ;
        RECT 124.610 189.495 124.930 189.555 ;
        RECT 127.670 189.495 127.990 189.555 ;
        RECT 129.370 189.495 129.690 189.555 ;
        RECT 131.750 189.495 132.070 189.555 ;
        RECT 111.835 189.235 112.205 189.305 ;
        RECT 113.390 189.235 113.710 189.295 ;
        RECT 111.835 189.095 113.710 189.235 ;
        RECT 111.835 189.025 112.205 189.095 ;
        RECT 113.390 189.035 113.710 189.095 ;
        RECT 116.450 189.235 116.770 189.295 ;
        RECT 118.150 189.235 118.470 189.295 ;
        RECT 116.450 189.095 118.470 189.235 ;
        RECT 116.450 189.035 116.770 189.095 ;
        RECT 118.150 189.035 118.470 189.095 ;
        RECT 119.850 189.235 120.170 189.295 ;
        RECT 121.550 189.235 121.870 189.295 ;
        RECT 124.270 189.235 124.590 189.295 ;
        RECT 119.850 189.095 124.590 189.235 ;
        RECT 119.850 189.035 120.170 189.095 ;
        RECT 121.550 189.035 121.870 189.095 ;
        RECT 124.270 189.035 124.590 189.095 ;
        RECT 125.290 189.235 125.610 189.295 ;
        RECT 135.490 189.235 135.810 189.295 ;
        RECT 125.290 189.095 135.810 189.235 ;
        RECT 125.290 189.035 125.610 189.095 ;
        RECT 135.490 189.035 135.810 189.095 ;
        RECT 122.035 188.835 122.405 188.845 ;
        RECT 114.070 188.775 114.390 188.835 ;
        RECT 119.510 188.775 119.830 188.835 ;
        RECT 114.070 188.635 119.830 188.775 ;
        RECT 114.070 188.575 114.390 188.635 ;
        RECT 119.510 188.575 119.830 188.635 ;
        RECT 121.890 188.575 122.405 188.835 ;
        RECT 140.590 188.775 140.910 188.835 ;
        RECT 142.630 188.775 142.950 188.835 ;
        RECT 140.590 188.635 142.950 188.775 ;
        RECT 140.590 188.575 140.910 188.635 ;
        RECT 142.630 188.575 142.950 188.635 ;
        RECT 122.035 188.565 122.405 188.575 ;
        RECT 114.410 188.315 114.730 188.375 ;
        RECT 118.830 188.315 119.150 188.375 ;
        RECT 120.870 188.315 121.190 188.375 ;
        RECT 127.330 188.315 127.650 188.375 ;
        RECT 114.410 188.175 127.650 188.315 ;
        RECT 114.410 188.115 114.730 188.175 ;
        RECT 118.830 188.115 119.150 188.175 ;
        RECT 120.870 188.115 121.190 188.175 ;
        RECT 127.330 188.115 127.650 188.175 ;
        RECT 135.150 188.315 135.470 188.375 ;
        RECT 138.210 188.315 138.530 188.375 ;
        RECT 138.890 188.315 139.210 188.375 ;
        RECT 145.350 188.315 145.670 188.375 ;
        RECT 135.150 188.175 145.670 188.315 ;
        RECT 135.150 188.115 135.470 188.175 ;
        RECT 138.210 188.115 138.530 188.175 ;
        RECT 138.890 188.115 139.210 188.175 ;
        RECT 145.350 188.115 145.670 188.175 ;
        RECT 119.850 187.855 120.170 187.915 ;
        RECT 127.330 187.855 127.650 187.915 ;
        RECT 119.850 187.715 127.650 187.855 ;
        RECT 119.850 187.655 120.170 187.715 ;
        RECT 127.330 187.655 127.650 187.715 ;
        RECT 128.010 187.855 128.330 187.915 ;
        RECT 129.710 187.855 130.030 187.915 ;
        RECT 128.010 187.715 130.030 187.855 ;
        RECT 128.010 187.655 128.330 187.715 ;
        RECT 129.710 187.655 130.030 187.715 ;
        RECT 130.390 187.855 130.710 187.915 ;
        RECT 135.150 187.855 135.470 187.915 ;
        RECT 141.610 187.855 141.930 187.915 ;
        RECT 143.650 187.855 143.970 187.915 ;
        RECT 130.390 187.715 141.330 187.855 ;
        RECT 130.390 187.655 130.710 187.715 ;
        RECT 135.150 187.655 135.470 187.715 ;
        RECT 118.830 187.395 119.150 187.455 ;
        RECT 121.890 187.395 122.210 187.455 ;
        RECT 118.830 187.255 122.210 187.395 ;
        RECT 118.830 187.195 119.150 187.255 ;
        RECT 121.890 187.195 122.210 187.255 ;
        RECT 122.570 187.395 122.890 187.455 ;
        RECT 126.990 187.395 127.310 187.455 ;
        RECT 122.570 187.255 127.310 187.395 ;
        RECT 122.570 187.195 122.890 187.255 ;
        RECT 126.990 187.195 127.310 187.255 ;
        RECT 129.710 187.395 130.030 187.455 ;
        RECT 132.770 187.395 133.090 187.455 ;
        RECT 129.710 187.255 133.090 187.395 ;
        RECT 129.710 187.195 130.030 187.255 ;
        RECT 132.770 187.195 133.090 187.255 ;
        RECT 135.635 187.395 136.005 187.465 ;
        RECT 140.590 187.395 140.910 187.455 ;
        RECT 135.635 187.255 140.910 187.395 ;
        RECT 141.190 187.395 141.330 187.715 ;
        RECT 141.610 187.715 143.970 187.855 ;
        RECT 141.610 187.655 141.930 187.715 ;
        RECT 143.650 187.655 143.970 187.715 ;
        RECT 146.030 187.855 146.350 187.915 ;
        RECT 149.235 187.855 149.605 187.925 ;
        RECT 146.030 187.715 149.605 187.855 ;
        RECT 146.030 187.655 146.350 187.715 ;
        RECT 149.235 187.645 149.605 187.715 ;
        RECT 142.970 187.395 143.290 187.455 ;
        RECT 141.190 187.255 143.290 187.395 ;
        RECT 135.635 187.185 136.005 187.255 ;
        RECT 140.590 187.195 140.910 187.255 ;
        RECT 142.970 187.195 143.290 187.255 ;
        RECT 122.230 186.935 122.550 186.995 ;
        RECT 124.270 186.935 124.590 186.995 ;
        RECT 129.370 186.935 129.690 186.995 ;
        RECT 122.230 186.795 129.690 186.935 ;
        RECT 122.230 186.735 122.550 186.795 ;
        RECT 124.270 186.735 124.590 186.795 ;
        RECT 129.370 186.735 129.690 186.795 ;
        RECT 136.170 186.935 136.490 186.995 ;
        RECT 138.210 186.935 138.530 186.995 ;
        RECT 136.170 186.795 138.530 186.935 ;
        RECT 136.170 186.735 136.490 186.795 ;
        RECT 138.210 186.735 138.530 186.795 ;
        RECT 145.835 186.535 146.205 186.545 ;
        RECT 117.130 186.475 117.450 186.535 ;
        RECT 124.270 186.475 124.590 186.535 ;
        RECT 117.130 186.335 124.590 186.475 ;
        RECT 117.130 186.275 117.450 186.335 ;
        RECT 124.270 186.275 124.590 186.335 ;
        RECT 130.730 186.475 131.050 186.535 ;
        RECT 135.150 186.475 135.470 186.535 ;
        RECT 139.910 186.475 140.230 186.535 ;
        RECT 130.730 186.335 135.470 186.475 ;
        RECT 130.730 186.275 131.050 186.335 ;
        RECT 135.150 186.275 135.470 186.335 ;
        RECT 135.750 186.335 140.230 186.475 ;
        RECT 114.410 186.015 114.730 186.075 ;
        RECT 118.830 186.015 119.150 186.075 ;
        RECT 114.410 185.875 119.150 186.015 ;
        RECT 114.410 185.815 114.730 185.875 ;
        RECT 118.830 185.815 119.150 185.875 ;
        RECT 121.550 186.015 121.870 186.075 ;
        RECT 127.330 186.015 127.650 186.075 ;
        RECT 121.550 185.875 127.650 186.015 ;
        RECT 121.550 185.815 121.870 185.875 ;
        RECT 127.330 185.815 127.650 185.875 ;
        RECT 132.770 186.015 133.090 186.075 ;
        RECT 135.150 186.015 135.470 186.075 ;
        RECT 135.750 186.015 135.890 186.335 ;
        RECT 139.910 186.275 140.230 186.335 ;
        RECT 145.835 186.275 146.350 186.535 ;
        RECT 145.835 186.265 146.205 186.275 ;
        RECT 132.770 185.875 135.890 186.015 ;
        RECT 138.890 186.015 139.210 186.075 ;
        RECT 139.910 186.015 140.230 186.075 ;
        RECT 138.890 185.875 140.230 186.015 ;
        RECT 132.770 185.815 133.090 185.875 ;
        RECT 135.150 185.815 135.470 185.875 ;
        RECT 138.890 185.815 139.210 185.875 ;
        RECT 139.910 185.815 140.230 185.875 ;
        RECT 108.435 185.555 108.805 185.625 ;
        RECT 119.170 185.555 119.490 185.615 ;
        RECT 108.435 185.415 119.490 185.555 ;
        RECT 108.435 185.345 108.805 185.415 ;
        RECT 119.170 185.355 119.490 185.415 ;
        RECT 135.830 185.555 136.150 185.615 ;
        RECT 138.210 185.555 138.530 185.615 ;
        RECT 145.350 185.555 145.670 185.615 ;
        RECT 135.830 185.415 145.670 185.555 ;
        RECT 135.830 185.355 136.150 185.415 ;
        RECT 138.210 185.355 138.530 185.415 ;
        RECT 145.350 185.355 145.670 185.415 ;
        RECT 116.110 185.095 116.430 185.155 ;
        RECT 118.830 185.095 119.150 185.155 ;
        RECT 121.210 185.095 121.530 185.155 ;
        RECT 116.110 184.955 121.530 185.095 ;
        RECT 116.110 184.895 116.430 184.955 ;
        RECT 118.830 184.895 119.150 184.955 ;
        RECT 121.210 184.895 121.530 184.955 ;
        RECT 132.235 185.095 132.605 185.165 ;
        RECT 132.770 185.095 133.090 185.155 ;
        RECT 132.235 184.955 133.090 185.095 ;
        RECT 132.235 184.885 132.605 184.955 ;
        RECT 132.770 184.895 133.090 184.955 ;
        RECT 139.035 185.095 139.405 185.165 ;
        RECT 140.590 185.095 140.910 185.155 ;
        RECT 139.035 184.955 140.910 185.095 ;
        RECT 139.035 184.885 139.405 184.955 ;
        RECT 140.590 184.895 140.910 184.955 ;
        RECT 142.435 185.095 142.805 185.165 ;
        RECT 143.650 185.095 143.970 185.155 ;
        RECT 142.435 184.955 143.970 185.095 ;
        RECT 142.435 184.885 142.805 184.955 ;
        RECT 143.650 184.895 143.970 184.955 ;
        RECT 146.030 185.095 146.350 185.155 ;
        RECT 152.635 185.095 153.005 185.165 ;
        RECT 146.030 184.955 153.005 185.095 ;
        RECT 146.030 184.895 146.350 184.955 ;
        RECT 152.635 184.885 153.005 184.955 ;
        RECT 100.970 182.410 102.630 184.070 ;
        RECT 123.240 180.480 125.770 180.490 ;
        RECT 100.360 180.380 108.770 180.390 ;
        RECT 100.360 180.100 108.805 180.380 ;
        RECT 123.240 180.200 125.805 180.480 ;
        RECT 123.240 180.190 125.770 180.200 ;
        RECT 100.360 180.090 108.770 180.100 ;
        RECT 100.360 105.820 100.660 180.090 ;
        RECT 100.860 179.630 118.970 179.640 ;
        RECT 100.860 179.350 119.005 179.630 ;
        RECT 100.860 179.340 118.970 179.350 ;
        RECT 100.860 120.760 101.160 179.340 ;
        RECT 101.580 178.940 122.370 178.950 ;
        RECT 101.580 178.660 122.405 178.940 ;
        RECT 101.580 178.650 122.370 178.660 ;
        RECT 101.580 135.760 101.880 178.650 ;
        RECT 102.210 178.350 115.570 178.360 ;
        RECT 102.210 178.070 115.605 178.350 ;
        RECT 102.210 178.060 115.570 178.070 ;
        RECT 102.210 150.840 102.510 178.060 ;
        RECT 102.770 177.660 112.170 177.670 ;
        RECT 102.770 177.380 112.205 177.660 ;
        RECT 102.770 177.370 112.170 177.380 ;
        RECT 102.790 165.570 103.090 177.370 ;
        RECT 106.840 176.770 107.540 176.780 ;
        RECT 106.500 176.030 107.850 176.770 ;
        RECT 106.840 166.600 107.540 176.030 ;
        RECT 117.980 174.620 118.880 176.640 ;
        RECT 116.255 172.705 116.575 172.760 ;
        RECT 116.255 172.550 118.860 172.705 ;
        RECT 116.255 172.500 116.575 172.550 ;
        RECT 108.890 171.080 116.880 171.470 ;
        RECT 108.820 168.770 109.400 169.400 ;
        RECT 111.430 168.020 114.090 171.080 ;
        RECT 108.930 167.570 116.870 168.020 ;
        RECT 106.750 165.810 107.610 166.600 ;
        RECT 106.840 161.770 107.540 161.780 ;
        RECT 106.500 161.030 107.850 161.770 ;
        RECT 106.840 151.600 107.540 161.030 ;
        RECT 116.160 157.690 116.480 157.750 ;
        RECT 116.160 157.550 118.510 157.690 ;
        RECT 116.160 157.490 116.480 157.550 ;
        RECT 108.890 156.080 116.880 156.470 ;
        RECT 108.790 153.690 109.370 154.320 ;
        RECT 111.430 153.020 114.090 156.080 ;
        RECT 108.930 152.570 116.870 153.020 ;
        RECT 102.210 150.540 103.050 150.840 ;
        RECT 106.750 150.810 107.610 151.600 ;
        RECT 106.840 146.720 107.540 146.730 ;
        RECT 106.500 145.980 107.850 146.720 ;
        RECT 106.840 136.550 107.540 145.980 ;
        RECT 116.400 142.635 116.720 142.690 ;
        RECT 116.400 142.485 118.115 142.635 ;
        RECT 116.400 142.430 116.720 142.485 ;
        RECT 108.890 141.030 116.880 141.420 ;
        RECT 108.790 138.740 109.370 139.370 ;
        RECT 111.430 137.970 114.090 141.030 ;
        RECT 108.930 137.520 116.870 137.970 ;
        RECT 106.750 135.760 107.610 136.550 ;
        RECT 101.580 135.460 103.130 135.760 ;
        RECT 106.840 131.720 107.540 131.730 ;
        RECT 106.500 130.980 107.850 131.720 ;
        RECT 106.840 121.550 107.540 130.980 ;
        RECT 116.290 127.640 116.610 127.680 ;
        RECT 116.290 127.460 117.690 127.640 ;
        RECT 116.290 127.420 116.610 127.460 ;
        RECT 108.890 126.030 116.880 126.420 ;
        RECT 108.790 123.740 109.370 124.370 ;
        RECT 111.430 122.970 114.090 126.030 ;
        RECT 108.930 122.520 116.870 122.970 ;
        RECT 106.750 120.760 107.610 121.550 ;
        RECT 100.860 120.460 103.170 120.760 ;
        RECT 106.790 116.780 107.490 116.790 ;
        RECT 106.450 116.040 107.800 116.780 ;
        RECT 106.790 106.610 107.490 116.040 ;
        RECT 116.510 112.675 116.830 112.720 ;
        RECT 116.510 112.505 117.195 112.675 ;
        RECT 116.510 112.460 116.830 112.505 ;
        RECT 108.840 111.090 116.830 111.480 ;
        RECT 108.750 108.700 109.330 109.330 ;
        RECT 111.380 108.030 114.040 111.090 ;
        RECT 108.880 107.580 116.820 108.030 ;
        RECT 106.700 105.820 107.560 106.610 ;
        RECT 100.360 105.520 103.080 105.820 ;
        RECT 99.710 103.665 112.290 103.900 ;
        RECT 99.225 103.175 110.620 103.390 ;
        RECT 98.780 102.760 109.045 102.970 ;
        RECT 98.170 102.210 107.455 102.480 ;
        RECT 97.505 101.665 105.905 101.930 ;
        RECT 96.825 101.075 104.305 101.360 ;
        RECT 96.145 100.400 102.800 100.700 ;
        RECT 95.400 99.790 101.275 100.035 ;
        RECT 88.560 93.290 88.820 93.610 ;
        RECT 101.030 92.875 101.275 99.790 ;
        RECT 102.500 92.925 102.800 100.400 ;
        RECT 104.020 92.925 104.305 101.075 ;
        RECT 105.640 92.955 105.905 101.665 ;
        RECT 100.620 92.615 101.680 92.875 ;
        RECT 102.120 92.625 103.180 92.925 ;
        RECT 103.630 92.640 104.690 92.925 ;
        RECT 105.240 92.690 106.300 92.955 ;
        RECT 107.185 92.925 107.455 102.210 ;
        RECT 108.835 92.955 109.045 102.760 ;
        RECT 106.790 92.655 107.850 92.925 ;
        RECT 108.410 92.695 109.470 92.955 ;
        RECT 110.405 92.925 110.620 103.175 ;
        RECT 112.055 92.945 112.290 103.665 ;
        RECT 117.025 101.605 117.195 112.505 ;
        RECT 117.510 102.010 117.690 127.460 ;
        RECT 117.965 102.335 118.115 142.485 ;
        RECT 118.370 102.640 118.510 157.550 ;
        RECT 118.705 102.965 118.860 172.550 ;
        RECT 123.240 169.890 123.540 180.190 ;
        RECT 120.480 169.590 123.540 169.890 ;
        RECT 123.830 179.710 129.170 179.720 ;
        RECT 123.830 179.430 129.205 179.710 ;
        RECT 152.680 179.480 152.960 179.515 ;
        RECT 123.830 179.420 129.170 179.430 ;
        RECT 120.480 105.740 120.780 169.590 ;
        RECT 123.830 168.770 124.130 179.420 ;
        RECT 143.320 179.180 152.970 179.480 ;
        RECT 121.150 168.470 124.130 168.770 ;
        RECT 124.430 179.000 132.570 179.010 ;
        RECT 124.430 178.720 132.605 179.000 ;
        RECT 124.430 178.710 132.570 178.720 ;
        RECT 121.150 120.900 121.450 168.470 ;
        RECT 124.430 167.820 124.730 178.710 ;
        RECT 121.750 167.520 124.730 167.820 ;
        RECT 124.920 178.280 135.970 178.290 ;
        RECT 124.920 178.000 136.005 178.280 ;
        RECT 124.920 177.990 135.970 178.000 ;
        RECT 121.750 135.710 122.050 167.520 ;
        RECT 124.920 166.810 125.220 177.990 ;
        RECT 122.310 166.510 125.220 166.810 ;
        RECT 125.540 177.560 142.770 177.570 ;
        RECT 125.540 177.280 142.805 177.560 ;
        RECT 125.540 177.270 142.770 177.280 ;
        RECT 122.310 150.820 122.610 166.510 ;
        RECT 125.540 166.000 125.840 177.270 ;
        RECT 126.720 176.720 127.420 176.730 ;
        RECT 126.380 175.980 127.730 176.720 ;
        RECT 126.720 166.550 127.420 175.980 ;
        RECT 137.800 174.600 138.700 176.620 ;
        RECT 136.460 172.635 136.780 172.690 ;
        RECT 136.460 172.485 138.465 172.635 ;
        RECT 136.460 172.430 136.780 172.485 ;
        RECT 128.770 171.030 136.760 171.420 ;
        RECT 128.680 168.760 129.260 169.390 ;
        RECT 131.310 167.970 133.970 171.030 ;
        RECT 128.810 167.520 136.750 167.970 ;
        RECT 122.900 165.700 125.840 166.000 ;
        RECT 126.630 165.760 127.490 166.550 ;
        RECT 126.720 161.770 127.420 161.780 ;
        RECT 126.380 161.030 127.730 161.770 ;
        RECT 126.720 151.600 127.420 161.030 ;
        RECT 136.270 157.695 136.590 157.720 ;
        RECT 136.270 157.485 138.095 157.695 ;
        RECT 136.270 157.460 136.590 157.485 ;
        RECT 128.770 156.080 136.760 156.470 ;
        RECT 128.680 153.800 129.260 154.430 ;
        RECT 131.310 153.020 133.970 156.080 ;
        RECT 128.810 152.570 136.750 153.020 ;
        RECT 122.310 150.520 122.980 150.820 ;
        RECT 126.630 150.810 127.490 151.600 ;
        RECT 126.720 146.720 127.420 146.730 ;
        RECT 126.380 145.980 127.730 146.720 ;
        RECT 126.720 136.550 127.420 145.980 ;
        RECT 136.150 142.705 136.470 142.750 ;
        RECT 136.150 142.535 137.715 142.705 ;
        RECT 136.150 142.490 136.470 142.535 ;
        RECT 128.770 141.030 136.760 141.420 ;
        RECT 128.680 138.730 129.260 139.360 ;
        RECT 131.310 137.970 133.970 141.030 ;
        RECT 128.810 137.520 136.750 137.970 ;
        RECT 126.630 135.760 127.490 136.550 ;
        RECT 121.750 135.410 122.980 135.710 ;
        RECT 126.720 131.780 127.420 131.790 ;
        RECT 126.380 131.040 127.730 131.780 ;
        RECT 126.720 121.610 127.420 131.040 ;
        RECT 136.335 127.700 136.655 127.760 ;
        RECT 136.335 127.555 137.375 127.700 ;
        RECT 136.335 127.500 136.655 127.555 ;
        RECT 128.770 126.090 136.760 126.480 ;
        RECT 128.610 123.790 129.190 124.420 ;
        RECT 131.310 123.030 133.970 126.090 ;
        RECT 128.810 122.580 136.750 123.030 ;
        RECT 121.150 120.600 123.010 120.900 ;
        RECT 126.630 120.820 127.490 121.610 ;
        RECT 126.720 116.780 127.420 116.790 ;
        RECT 126.380 116.040 127.730 116.780 ;
        RECT 126.720 106.610 127.420 116.040 ;
        RECT 136.160 112.690 136.480 112.750 ;
        RECT 136.160 112.550 137.090 112.690 ;
        RECT 136.160 112.490 136.480 112.550 ;
        RECT 128.770 111.090 136.760 111.480 ;
        RECT 128.730 108.760 129.310 109.390 ;
        RECT 131.310 108.030 133.970 111.090 ;
        RECT 128.810 107.580 136.750 108.030 ;
        RECT 126.630 105.820 127.490 106.610 ;
        RECT 120.480 105.440 123.040 105.740 ;
        RECT 136.950 103.450 137.090 112.550 ;
        RECT 137.230 103.740 137.375 127.555 ;
        RECT 137.545 104.065 137.715 142.535 ;
        RECT 137.885 104.455 138.095 157.485 ;
        RECT 138.315 104.825 138.465 172.485 ;
        RECT 143.320 169.390 143.620 179.180 ;
        RECT 152.680 179.145 152.960 179.180 ;
        RECT 140.280 169.090 143.620 169.390 ;
        RECT 144.050 178.740 146.170 178.750 ;
        RECT 144.050 178.460 146.205 178.740 ;
        RECT 144.050 178.450 146.170 178.460 ;
        RECT 140.280 105.820 140.580 169.090 ;
        RECT 144.050 168.490 144.350 178.450 ;
        RECT 145.290 178.030 149.570 178.040 ;
        RECT 145.290 177.750 149.605 178.030 ;
        RECT 145.290 177.740 149.570 177.750 ;
        RECT 144.680 176.850 144.960 176.885 ;
        RECT 140.940 168.190 144.350 168.490 ;
        RECT 140.940 120.830 141.240 168.190 ;
        RECT 144.670 167.700 144.970 176.850 ;
        RECT 141.710 167.400 144.970 167.700 ;
        RECT 141.710 135.850 142.010 167.400 ;
        RECT 145.290 166.930 145.590 177.740 ;
        RECT 142.350 166.630 145.590 166.930 ;
        RECT 145.960 177.370 148.420 177.380 ;
        RECT 145.960 177.090 148.455 177.370 ;
        RECT 145.960 177.080 148.420 177.090 ;
        RECT 142.350 150.730 142.650 166.630 ;
        RECT 145.960 166.020 146.260 177.080 ;
        RECT 146.750 176.770 147.450 176.780 ;
        RECT 146.410 176.030 147.760 176.770 ;
        RECT 146.750 166.600 147.450 176.030 ;
        RECT 157.570 174.580 158.470 176.600 ;
        RECT 156.415 172.650 156.735 172.710 ;
        RECT 156.415 172.505 158.350 172.650 ;
        RECT 156.415 172.450 156.735 172.505 ;
        RECT 148.800 171.080 156.790 171.470 ;
        RECT 148.880 168.740 149.460 169.370 ;
        RECT 151.340 168.020 154.000 171.080 ;
        RECT 148.840 167.570 156.780 168.020 ;
        RECT 142.960 165.720 146.260 166.020 ;
        RECT 146.660 165.810 147.520 166.600 ;
        RECT 146.800 161.720 147.500 161.730 ;
        RECT 146.460 160.980 147.810 161.720 ;
        RECT 146.800 151.550 147.500 160.980 ;
        RECT 156.500 157.640 156.820 157.700 ;
        RECT 156.500 157.500 158.030 157.640 ;
        RECT 156.500 157.440 156.820 157.500 ;
        RECT 148.850 156.030 156.840 156.420 ;
        RECT 148.920 153.710 149.500 154.340 ;
        RECT 151.390 152.970 154.050 156.030 ;
        RECT 148.890 152.520 156.830 152.970 ;
        RECT 146.710 150.760 147.570 151.550 ;
        RECT 142.350 150.430 142.970 150.730 ;
        RECT 146.750 146.720 147.450 146.730 ;
        RECT 146.410 145.980 147.760 146.720 ;
        RECT 146.750 136.550 147.450 145.980 ;
        RECT 156.330 142.625 156.590 142.710 ;
        RECT 156.330 142.475 157.705 142.625 ;
        RECT 156.330 142.390 156.590 142.475 ;
        RECT 148.800 141.030 156.790 141.420 ;
        RECT 148.830 138.670 149.410 139.300 ;
        RECT 151.340 137.970 154.000 141.030 ;
        RECT 148.840 137.520 156.780 137.970 ;
        RECT 141.710 135.550 143.010 135.850 ;
        RECT 146.660 135.760 147.520 136.550 ;
        RECT 146.750 131.780 147.450 131.790 ;
        RECT 146.410 131.040 147.760 131.780 ;
        RECT 146.750 121.610 147.450 131.040 ;
        RECT 156.410 127.660 156.730 127.720 ;
        RECT 156.410 127.520 157.410 127.660 ;
        RECT 156.410 127.460 156.730 127.520 ;
        RECT 148.800 126.090 156.790 126.480 ;
        RECT 148.950 123.750 149.530 124.380 ;
        RECT 151.340 123.030 154.000 126.090 ;
        RECT 148.840 122.580 156.780 123.030 ;
        RECT 140.940 120.530 142.990 120.830 ;
        RECT 146.660 120.820 147.520 121.610 ;
        RECT 146.750 116.780 147.450 116.790 ;
        RECT 146.410 116.040 147.760 116.780 ;
        RECT 146.750 106.610 147.450 116.040 ;
        RECT 156.000 112.715 156.320 112.770 ;
        RECT 156.000 112.565 157.115 112.715 ;
        RECT 156.000 112.510 156.320 112.565 ;
        RECT 148.800 111.090 156.790 111.480 ;
        RECT 148.910 108.790 149.490 109.420 ;
        RECT 151.340 108.030 154.000 111.090 ;
        RECT 148.840 107.580 156.780 108.030 ;
        RECT 146.660 105.820 147.520 106.610 ;
        RECT 140.280 105.520 143.020 105.820 ;
        RECT 138.315 104.675 149.650 104.825 ;
        RECT 137.885 104.245 147.750 104.455 ;
        RECT 137.545 103.895 146.220 104.065 ;
        RECT 137.230 103.595 144.785 103.740 ;
        RECT 136.950 103.310 143.320 103.450 ;
        RECT 118.705 102.810 141.785 102.965 ;
        RECT 118.370 102.500 140.290 102.640 ;
        RECT 117.965 102.185 138.860 102.335 ;
        RECT 117.510 101.970 137.340 102.010 ;
        RECT 117.510 101.830 137.730 101.970 ;
        RECT 137.160 101.620 137.730 101.830 ;
        RECT 117.025 101.435 135.840 101.605 ;
        RECT 137.210 101.500 137.730 101.620 ;
        RECT 135.670 99.200 135.840 101.435 ;
        RECT 138.710 99.390 138.860 102.185 ;
        RECT 140.150 101.990 140.290 102.500 ;
        RECT 140.150 101.620 140.700 101.990 ;
        RECT 140.180 101.520 140.700 101.620 ;
        RECT 135.670 98.995 136.300 99.200 ;
        RECT 138.710 99.015 139.270 99.390 ;
        RECT 135.690 98.720 136.300 98.995 ;
        RECT 138.750 98.920 139.270 99.015 ;
        RECT 141.630 99.310 141.785 102.810 ;
        RECT 143.180 102.050 143.320 103.310 ;
        RECT 143.180 101.580 143.700 102.050 ;
        RECT 144.640 99.340 144.785 103.595 ;
        RECT 146.050 102.080 146.220 103.895 ;
        RECT 146.050 101.950 146.610 102.080 ;
        RECT 146.090 101.610 146.610 101.950 ;
        RECT 147.540 99.390 147.750 104.245 ;
        RECT 149.500 101.940 149.650 104.675 ;
        RECT 156.965 103.015 157.115 112.565 ;
        RECT 149.120 101.705 149.650 101.940 ;
        RECT 150.960 102.865 157.115 103.015 ;
        RECT 149.120 101.470 149.640 101.705 ;
        RECT 141.630 98.955 142.180 99.310 ;
        RECT 141.660 98.840 142.180 98.955 ;
        RECT 144.640 98.870 145.160 99.340 ;
        RECT 147.540 99.075 148.230 99.390 ;
        RECT 150.960 99.310 151.110 102.865 ;
        RECT 157.270 102.720 157.410 127.520 ;
        RECT 152.470 102.580 157.410 102.720 ;
        RECT 152.470 102.060 152.610 102.580 ;
        RECT 157.555 102.375 157.705 142.475 ;
        RECT 152.090 101.590 152.610 102.060 ;
        RECT 153.960 102.225 157.705 102.375 ;
        RECT 147.560 98.860 148.230 99.075 ;
        RECT 150.570 99.055 151.110 99.310 ;
        RECT 153.960 99.280 154.110 102.225 ;
        RECT 155.040 101.990 155.560 102.050 ;
        RECT 157.890 101.990 158.030 157.500 ;
        RECT 155.040 101.850 158.030 101.990 ;
        RECT 155.040 101.580 155.560 101.850 ;
        RECT 158.205 99.285 158.350 172.505 ;
        RECT 153.580 99.115 154.110 99.280 ;
        RECT 156.480 99.140 158.350 99.285 ;
        RECT 150.570 98.840 151.090 99.055 ;
        RECT 153.580 98.810 154.100 99.115 ;
        RECT 156.510 98.780 157.030 99.140 ;
        RECT 109.980 92.665 111.040 92.925 ;
        RECT 111.640 92.685 112.700 92.945 ;
        RECT 88.100 90.570 88.360 90.890 ;
        RECT 100.150 90.045 100.470 90.915 ;
        RECT 100.140 89.015 100.470 90.045 ;
        RECT 101.820 90.025 102.140 90.905 ;
        RECT 100.140 87.255 100.450 89.015 ;
        RECT 101.800 89.005 102.140 90.025 ;
        RECT 103.380 89.005 103.700 90.905 ;
        RECT 104.920 90.015 105.240 90.915 ;
        RECT 104.900 89.015 105.240 90.015 ;
        RECT 106.510 89.825 106.830 90.935 ;
        RECT 101.800 87.365 102.110 89.005 ;
        RECT 100.140 87.095 100.360 87.255 ;
        RECT 100.610 87.095 101.150 87.235 ;
        RECT 88.560 85.130 88.820 85.450 ;
        RECT 87.640 83.090 87.900 83.410 ;
        RECT 87.180 80.370 87.440 80.690 ;
        RECT 87.700 79.670 87.840 83.090 ;
        RECT 88.090 82.895 88.370 83.265 ;
        RECT 87.640 79.350 87.900 79.670 ;
        RECT 86.720 79.070 86.980 79.330 ;
        RECT 86.720 79.010 87.380 79.070 ;
        RECT 86.780 78.930 87.380 79.010 ;
        RECT 86.720 77.310 86.980 77.630 ;
        RECT 86.780 72.870 86.920 77.310 ;
        RECT 87.240 74.570 87.380 78.930 ;
        RECT 87.640 77.990 87.900 78.310 ;
        RECT 87.180 74.250 87.440 74.570 ;
        RECT 86.720 72.550 86.980 72.870 ;
        RECT 83.560 69.970 84.160 70.110 ;
        RECT 85.860 70.090 86.460 70.230 ;
        RECT 83.040 69.150 83.300 69.470 ;
        RECT 82.580 68.130 82.840 68.450 ;
        RECT 82.120 67.110 82.380 67.430 ;
        RECT 81.200 66.430 81.460 66.750 ;
        RECT 80.740 66.090 81.000 66.410 ;
        RECT 80.800 64.710 80.940 66.090 ;
        RECT 80.740 64.390 81.000 64.710 ;
        RECT 81.260 64.030 81.400 66.430 ;
        RECT 82.120 65.470 82.380 65.730 ;
        RECT 81.720 65.410 82.380 65.470 ;
        RECT 81.720 65.330 82.320 65.410 ;
        RECT 81.200 63.710 81.460 64.030 ;
        RECT 81.260 60.970 81.400 63.710 ;
        RECT 81.720 61.990 81.860 65.330 ;
        RECT 82.640 63.690 82.780 68.130 ;
        RECT 82.580 63.370 82.840 63.690 ;
        RECT 83.040 63.030 83.300 63.350 ;
        RECT 83.100 61.990 83.240 63.030 ;
        RECT 81.660 61.670 81.920 61.990 ;
        RECT 83.040 61.670 83.300 61.990 ;
        RECT 83.560 61.220 83.700 69.970 ;
        RECT 83.960 68.985 84.220 69.130 ;
        RECT 83.950 68.615 84.230 68.985 ;
        RECT 84.880 68.810 85.140 69.130 ;
        RECT 85.340 69.040 85.600 69.130 ;
        RECT 85.860 69.040 86.000 70.090 ;
        RECT 86.260 69.150 86.520 69.470 ;
        RECT 85.340 68.900 86.000 69.040 ;
        RECT 85.340 68.810 85.600 68.900 ;
        RECT 84.420 68.130 84.680 68.450 ;
        RECT 84.480 66.945 84.620 68.130 ;
        RECT 84.410 66.575 84.690 66.945 ;
        RECT 83.960 61.220 84.220 61.310 ;
        RECT 83.560 61.080 84.220 61.220 ;
        RECT 83.960 60.990 84.220 61.080 ;
        RECT 80.740 60.650 81.000 60.970 ;
        RECT 81.200 60.650 81.460 60.970 ;
        RECT 80.800 57.570 80.940 60.650 ;
        RECT 82.580 59.970 82.840 60.290 ;
        RECT 82.640 59.465 82.780 59.970 ;
        RECT 82.570 59.095 82.850 59.465 ;
        RECT 83.040 58.950 83.300 59.270 ;
        RECT 80.740 57.250 81.000 57.570 ;
        RECT 80.800 56.210 80.940 57.250 ;
        RECT 80.740 55.890 81.000 56.210 ;
        RECT 80.280 55.550 80.540 55.870 ;
        RECT 81.660 55.550 81.920 55.870 ;
        RECT 78.500 55.130 79.100 55.270 ;
        RECT 78.500 49.750 78.640 55.130 ;
        RECT 79.350 55.015 79.630 55.385 ;
        RECT 79.360 54.870 79.620 55.015 ;
        RECT 78.900 54.530 79.160 54.850 ;
        RECT 79.820 54.530 80.080 54.850 ;
        RECT 78.960 53.490 79.100 54.530 ;
        RECT 78.900 53.170 79.160 53.490 ;
        RECT 79.880 50.770 80.020 54.530 ;
        RECT 79.820 50.450 80.080 50.770 ;
        RECT 78.440 49.430 78.700 49.750 ;
        RECT 78.500 47.370 78.640 49.430 ;
        RECT 77.980 47.050 78.240 47.370 ;
        RECT 78.440 47.050 78.700 47.370 ;
        RECT 78.900 47.225 79.160 47.370 ;
        RECT 76.600 41.610 76.860 41.930 ;
        RECT 77.520 41.610 77.780 41.930 ;
        RECT 76.140 39.460 76.400 39.550 ;
        RECT 75.740 39.320 76.400 39.460 ;
        RECT 76.140 39.230 76.400 39.320 ;
        RECT 74.360 36.150 74.500 39.230 ;
        RECT 74.760 38.950 75.020 39.210 ;
        RECT 74.760 38.890 75.880 38.950 ;
        RECT 74.820 38.810 75.880 38.890 ;
        RECT 75.740 38.530 75.880 38.810 ;
        RECT 75.220 38.210 75.480 38.530 ;
        RECT 75.680 38.210 75.940 38.530 ;
        RECT 74.300 35.830 74.560 36.150 ;
        RECT 74.760 35.490 75.020 35.810 ;
        RECT 73.380 34.130 73.640 34.450 ;
        RECT 74.820 33.430 74.960 35.490 ;
        RECT 75.280 34.190 75.420 38.210 ;
        RECT 76.200 36.830 76.340 39.230 ;
        RECT 76.660 39.210 76.800 41.610 ;
        RECT 76.600 38.890 76.860 39.210 ;
        RECT 77.060 38.890 77.320 39.210 ;
        RECT 76.140 36.510 76.400 36.830 ;
        RECT 75.680 35.830 75.940 36.150 ;
        RECT 75.740 34.985 75.880 35.830 ;
        RECT 75.670 34.615 75.950 34.985 ;
        RECT 75.680 34.190 75.940 34.450 ;
        RECT 75.280 34.130 75.940 34.190 ;
        RECT 75.280 34.050 75.880 34.130 ;
        RECT 76.140 33.790 76.400 34.110 ;
        RECT 76.200 33.430 76.340 33.790 ;
        RECT 74.760 33.110 75.020 33.430 ;
        RECT 76.140 33.110 76.400 33.430 ;
        RECT 73.380 32.770 73.640 33.090 ;
        RECT 73.440 28.670 73.580 32.770 ;
        RECT 75.680 28.690 75.940 29.010 ;
        RECT 73.380 28.350 73.640 28.670 ;
        RECT 72.000 25.290 72.260 25.610 ;
        RECT 68.780 24.950 69.040 25.270 ;
        RECT 75.740 23.570 75.880 28.690 ;
        RECT 76.200 26.290 76.340 33.110 ;
        RECT 76.140 25.970 76.400 26.290 ;
        RECT 76.140 24.950 76.400 25.270 ;
        RECT 76.200 23.910 76.340 24.950 ;
        RECT 76.140 23.590 76.400 23.910 ;
        RECT 66.480 23.250 66.740 23.570 ;
        RECT 75.680 23.250 75.940 23.570 ;
        RECT 60.960 22.570 61.220 22.890 ;
        RECT 61.420 22.570 61.680 22.890 ;
        RECT 61.020 20.850 61.160 22.570 ;
        RECT 75.680 22.230 75.940 22.550 ;
        RECT 60.960 20.530 61.220 20.850 ;
        RECT 53.140 20.190 53.400 20.510 ;
        RECT 75.740 20.170 75.880 22.230 ;
        RECT 76.200 20.170 76.340 23.590 ;
        RECT 76.660 20.170 76.800 38.890 ;
        RECT 77.120 37.510 77.260 38.890 ;
        RECT 77.060 37.190 77.320 37.510 ;
        RECT 77.580 37.170 77.720 41.610 ;
        RECT 78.040 40.230 78.180 47.050 ;
        RECT 78.890 46.855 79.170 47.225 ;
        RECT 80.340 47.110 80.480 55.550 ;
        RECT 81.200 52.490 81.460 52.810 ;
        RECT 80.740 51.810 81.000 52.130 ;
        RECT 81.260 51.870 81.400 52.490 ;
        RECT 81.720 52.470 81.860 55.550 ;
        RECT 82.580 52.550 82.840 52.810 ;
        RECT 83.100 52.665 83.240 58.950 ;
        RECT 82.180 52.490 82.840 52.550 ;
        RECT 81.660 52.150 81.920 52.470 ;
        RECT 82.180 52.410 82.780 52.490 ;
        RECT 80.800 50.770 80.940 51.810 ;
        RECT 81.260 51.730 81.860 51.870 ;
        RECT 80.740 50.450 81.000 50.770 ;
        RECT 81.200 49.770 81.460 50.090 ;
        RECT 80.740 47.730 81.000 48.050 ;
        RECT 79.880 46.970 80.480 47.110 ;
        RECT 79.360 43.650 79.620 43.970 ;
        RECT 78.900 42.630 79.160 42.950 ;
        RECT 78.960 42.465 79.100 42.630 ;
        RECT 78.890 42.095 79.170 42.465 ;
        RECT 79.420 41.590 79.560 43.650 ;
        RECT 79.880 41.930 80.020 46.970 ;
        RECT 80.800 46.690 80.940 47.730 ;
        RECT 81.260 47.710 81.400 49.770 ;
        RECT 81.200 47.390 81.460 47.710 ;
        RECT 80.280 46.370 80.540 46.690 ;
        RECT 80.740 46.370 81.000 46.690 ;
        RECT 80.340 44.990 80.480 46.370 ;
        RECT 81.260 45.330 81.400 47.390 ;
        RECT 81.720 46.690 81.860 51.730 ;
        RECT 82.180 47.030 82.320 52.410 ;
        RECT 83.030 52.295 83.310 52.665 ;
        RECT 83.500 52.490 83.760 52.810 ;
        RECT 82.580 49.090 82.840 49.410 ;
        RECT 82.640 47.370 82.780 49.090 ;
        RECT 82.580 47.050 82.840 47.370 ;
        RECT 82.120 46.710 82.380 47.030 ;
        RECT 81.660 46.370 81.920 46.690 ;
        RECT 81.200 45.010 81.460 45.330 ;
        RECT 80.280 44.670 80.540 44.990 ;
        RECT 81.260 42.270 81.400 45.010 ;
        RECT 81.200 41.950 81.460 42.270 ;
        RECT 79.820 41.610 80.080 41.930 ;
        RECT 78.440 41.270 78.700 41.590 ;
        RECT 79.360 41.270 79.620 41.590 ;
        RECT 77.980 39.910 78.240 40.230 ;
        RECT 78.500 39.550 78.640 41.270 ;
        RECT 78.900 40.930 79.160 41.250 ;
        RECT 78.960 39.890 79.100 40.930 ;
        RECT 79.880 39.890 80.020 41.610 ;
        RECT 78.900 39.570 79.160 39.890 ;
        RECT 79.820 39.570 80.080 39.890 ;
        RECT 78.440 39.230 78.700 39.550 ;
        RECT 79.360 39.230 79.620 39.550 ;
        RECT 77.520 36.850 77.780 37.170 ;
        RECT 77.520 36.400 77.780 36.490 ;
        RECT 77.520 36.260 79.100 36.400 ;
        RECT 77.520 36.170 77.780 36.260 ;
        RECT 77.520 35.720 77.780 35.810 ;
        RECT 78.440 35.720 78.700 35.810 ;
        RECT 77.520 35.580 78.700 35.720 ;
        RECT 77.520 35.490 77.780 35.580 ;
        RECT 77.520 33.450 77.780 33.770 ;
        RECT 77.580 26.630 77.720 33.450 ;
        RECT 78.040 32.070 78.180 35.580 ;
        RECT 78.440 35.490 78.700 35.580 ;
        RECT 78.440 33.790 78.700 34.110 ;
        RECT 78.500 33.090 78.640 33.790 ;
        RECT 78.440 32.770 78.700 33.090 ;
        RECT 77.980 31.750 78.240 32.070 ;
        RECT 78.440 30.730 78.700 31.050 ;
        RECT 77.520 26.310 77.780 26.630 ;
        RECT 77.060 24.610 77.320 24.930 ;
        RECT 77.120 23.230 77.260 24.610 ;
        RECT 77.580 23.230 77.720 26.310 ;
        RECT 78.500 25.610 78.640 30.730 ;
        RECT 78.960 27.650 79.100 36.260 ;
        RECT 79.420 36.150 79.560 39.230 ;
        RECT 79.880 36.490 80.020 39.570 ;
        RECT 80.270 38.015 80.550 38.385 ;
        RECT 80.340 37.170 80.480 38.015 ;
        RECT 80.280 36.850 80.540 37.170 ;
        RECT 79.820 36.170 80.080 36.490 ;
        RECT 79.360 35.830 79.620 36.150 ;
        RECT 80.270 35.975 80.550 36.345 ;
        RECT 80.280 35.830 80.540 35.975 ;
        RECT 80.740 35.490 81.000 35.810 ;
        RECT 80.800 34.190 80.940 35.490 ;
        RECT 79.420 34.050 80.940 34.190 ;
        RECT 78.900 27.330 79.160 27.650 ;
        RECT 77.980 25.290 78.240 25.610 ;
        RECT 78.440 25.290 78.700 25.610 ;
        RECT 78.040 23.230 78.180 25.290 ;
        RECT 77.060 22.910 77.320 23.230 ;
        RECT 77.520 22.910 77.780 23.230 ;
        RECT 77.980 22.910 78.240 23.230 ;
        RECT 78.960 22.550 79.100 27.330 ;
        RECT 79.420 23.910 79.560 34.050 ;
        RECT 79.820 33.450 80.080 33.770 ;
        RECT 79.880 31.050 80.020 33.450 ;
        RECT 80.280 32.770 80.540 33.090 ;
        RECT 79.820 30.730 80.080 31.050 ;
        RECT 80.340 30.710 80.480 32.770 ;
        RECT 81.260 31.050 81.400 41.950 ;
        RECT 81.650 39.375 81.930 39.745 ;
        RECT 81.660 39.220 81.920 39.375 ;
        RECT 81.660 38.210 81.920 38.530 ;
        RECT 81.720 36.150 81.860 38.210 ;
        RECT 81.660 35.830 81.920 36.150 ;
        RECT 81.200 30.730 81.460 31.050 ;
        RECT 80.280 30.390 80.540 30.710 ;
        RECT 81.260 29.010 81.400 30.730 ;
        RECT 81.200 28.690 81.460 29.010 ;
        RECT 80.270 27.815 80.550 28.185 ;
        RECT 79.360 23.590 79.620 23.910 ;
        RECT 80.340 23.570 80.480 27.815 ;
        RECT 81.260 25.950 81.400 28.690 ;
        RECT 81.720 27.990 81.860 35.830 ;
        RECT 82.180 34.110 82.320 46.710 ;
        RECT 82.570 42.095 82.850 42.465 ;
        RECT 82.640 40.230 82.780 42.095 ;
        RECT 83.030 40.735 83.310 41.105 ;
        RECT 82.580 39.910 82.840 40.230 ;
        RECT 82.625 39.460 82.885 39.550 ;
        RECT 83.100 39.460 83.240 40.735 ;
        RECT 83.560 39.745 83.700 52.490 ;
        RECT 82.625 39.320 83.240 39.460 ;
        RECT 83.490 39.375 83.770 39.745 ;
        RECT 82.625 39.230 82.885 39.320 ;
        RECT 82.570 38.695 82.850 39.065 ;
        RECT 82.580 38.550 82.840 38.695 ;
        RECT 83.100 37.170 83.240 39.320 ;
        RECT 83.040 36.850 83.300 37.170 ;
        RECT 83.040 35.490 83.300 35.810 ;
        RECT 82.570 34.615 82.850 34.985 ;
        RECT 82.640 34.110 82.780 34.615 ;
        RECT 82.120 33.790 82.380 34.110 ;
        RECT 82.580 33.790 82.840 34.110 ;
        RECT 82.180 33.430 82.320 33.790 ;
        RECT 82.120 33.110 82.380 33.430 ;
        RECT 82.570 28.495 82.850 28.865 ;
        RECT 81.660 27.670 81.920 27.990 ;
        RECT 81.200 25.630 81.460 25.950 ;
        RECT 80.730 25.095 81.010 25.465 ;
        RECT 80.280 23.250 80.540 23.570 ;
        RECT 79.360 22.910 79.620 23.230 ;
        RECT 78.900 22.230 79.160 22.550 ;
        RECT 79.420 20.850 79.560 22.910 ;
        RECT 80.340 22.210 80.480 23.250 ;
        RECT 79.820 21.890 80.080 22.210 ;
        RECT 80.280 21.890 80.540 22.210 ;
        RECT 79.360 20.530 79.620 20.850 ;
        RECT 79.880 20.170 80.020 21.890 ;
        RECT 80.340 20.170 80.480 21.890 ;
        RECT 80.800 21.190 80.940 25.095 ;
        RECT 81.260 23.230 81.400 25.630 ;
        RECT 81.200 22.910 81.460 23.230 ;
        RECT 82.640 21.190 82.780 28.495 ;
        RECT 83.100 23.570 83.240 35.490 ;
        RECT 83.560 34.790 83.700 39.375 ;
        RECT 84.020 37.025 84.160 60.990 ;
        RECT 84.480 57.570 84.620 66.575 ;
        RECT 84.420 57.250 84.680 57.570 ;
        RECT 84.940 56.210 85.080 68.810 ;
        RECT 85.400 63.010 85.540 68.810 ;
        RECT 86.320 64.370 86.460 69.150 ;
        RECT 86.720 68.470 86.980 68.790 ;
        RECT 86.780 65.730 86.920 68.470 ;
        RECT 86.720 65.410 86.980 65.730 ;
        RECT 86.260 64.050 86.520 64.370 ;
        RECT 85.340 62.690 85.600 63.010 ;
        RECT 85.800 61.670 86.060 61.990 ;
        RECT 85.330 58.415 85.610 58.785 ;
        RECT 84.880 55.890 85.140 56.210 ;
        RECT 85.400 52.810 85.540 58.415 ;
        RECT 85.860 52.810 86.000 61.670 ;
        RECT 86.320 55.530 86.460 64.050 ;
        RECT 87.240 58.250 87.380 74.250 ;
        RECT 87.700 73.065 87.840 77.990 ;
        RECT 87.630 72.695 87.910 73.065 ;
        RECT 87.640 68.130 87.900 68.450 ;
        RECT 87.700 64.710 87.840 68.130 ;
        RECT 87.640 64.390 87.900 64.710 ;
        RECT 87.630 62.495 87.910 62.865 ;
        RECT 87.180 57.930 87.440 58.250 ;
        RECT 87.180 57.250 87.440 57.570 ;
        RECT 87.240 56.210 87.380 57.250 ;
        RECT 87.180 55.890 87.440 56.210 ;
        RECT 86.720 55.550 86.980 55.870 ;
        RECT 86.260 55.210 86.520 55.530 ;
        RECT 85.340 52.490 85.600 52.810 ;
        RECT 85.800 52.490 86.060 52.810 ;
        RECT 85.400 51.110 85.540 52.490 ;
        RECT 86.260 52.150 86.520 52.470 ;
        RECT 85.340 50.790 85.600 51.110 ;
        RECT 85.340 50.110 85.600 50.430 ;
        RECT 84.420 41.270 84.680 41.590 ;
        RECT 84.480 40.230 84.620 41.270 ;
        RECT 84.420 39.910 84.680 40.230 ;
        RECT 84.870 40.055 85.150 40.425 ;
        RECT 84.880 39.910 85.140 40.055 ;
        RECT 85.400 39.550 85.540 50.110 ;
        RECT 86.320 41.250 86.460 52.150 ;
        RECT 86.780 48.390 86.920 55.550 ;
        RECT 87.240 52.470 87.380 55.890 ;
        RECT 87.700 53.830 87.840 62.495 ;
        RECT 88.160 59.270 88.300 82.895 ;
        RECT 88.620 68.790 88.760 85.130 ;
        RECT 100.140 85.005 101.150 87.095 ;
        RECT 100.180 84.985 101.150 85.005 ;
        RECT 101.800 87.045 102.610 87.365 ;
        RECT 103.380 87.235 103.690 89.005 ;
        RECT 101.800 84.985 102.530 87.045 ;
        RECT 100.540 84.895 101.150 84.985 ;
        RECT 102.080 84.955 102.530 84.985 ;
        RECT 102.110 84.925 102.480 84.955 ;
        RECT 103.380 84.945 104.050 87.235 ;
        RECT 104.900 87.215 105.210 89.015 ;
        RECT 106.470 87.245 106.840 89.825 ;
        RECT 108.070 89.815 108.390 90.905 ;
        RECT 109.660 89.855 109.980 90.925 ;
        RECT 111.260 90.165 111.540 90.915 ;
        RECT 108.050 87.275 108.420 89.815 ;
        RECT 104.900 84.975 105.560 87.215 ;
        RECT 103.500 84.885 104.050 84.945 ;
        RECT 105.010 84.865 105.560 84.975 ;
        RECT 106.470 84.895 107.020 87.245 ;
        RECT 107.950 84.925 108.500 87.275 ;
        RECT 109.660 87.265 110.010 89.855 ;
        RECT 111.240 87.275 111.540 90.165 ;
        RECT 109.400 85.015 110.010 87.265 ;
        RECT 109.400 84.915 109.950 85.015 ;
        RECT 110.900 84.985 111.540 87.275 ;
        RECT 110.900 84.925 111.450 84.985 ;
        RECT 88.560 68.470 88.820 68.790 ;
        RECT 88.100 58.950 88.360 59.270 ;
        RECT 87.640 53.510 87.900 53.830 ;
        RECT 87.180 52.150 87.440 52.470 ;
        RECT 87.630 48.895 87.910 49.265 ;
        RECT 86.720 48.070 86.980 48.390 ;
        RECT 86.780 44.990 86.920 48.070 ;
        RECT 87.700 45.670 87.840 48.895 ;
        RECT 88.100 46.370 88.360 46.690 ;
        RECT 87.640 45.350 87.900 45.670 ;
        RECT 86.720 44.670 86.980 44.990 ;
        RECT 86.260 40.930 86.520 41.250 ;
        RECT 86.780 40.230 86.920 44.670 ;
        RECT 87.640 40.930 87.900 41.250 ;
        RECT 86.720 39.910 86.980 40.230 ;
        RECT 87.700 39.550 87.840 40.930 ;
        RECT 85.340 39.230 85.600 39.550 ;
        RECT 86.720 39.230 86.980 39.550 ;
        RECT 87.640 39.230 87.900 39.550 ;
        RECT 86.780 37.510 86.920 39.230 ;
        RECT 87.700 37.705 87.840 39.230 ;
        RECT 86.720 37.190 86.980 37.510 ;
        RECT 87.630 37.335 87.910 37.705 ;
        RECT 83.950 36.655 84.230 37.025 ;
        RECT 84.870 36.655 85.150 37.025 ;
        RECT 84.940 36.490 85.080 36.655 ;
        RECT 84.880 36.170 85.140 36.490 ;
        RECT 85.800 36.170 86.060 36.490 ;
        RECT 86.260 36.170 86.520 36.490 ;
        RECT 87.180 36.170 87.440 36.490 ;
        RECT 83.500 34.470 83.760 34.790 ;
        RECT 83.560 34.110 83.700 34.470 ;
        RECT 83.500 33.790 83.760 34.110 ;
        RECT 83.560 33.090 83.700 33.790 ;
        RECT 83.500 32.770 83.760 33.090 ;
        RECT 83.960 32.770 84.220 33.090 ;
        RECT 84.020 28.670 84.160 32.770 ;
        RECT 85.860 31.730 86.000 36.170 ;
        RECT 85.800 31.410 86.060 31.730 ;
        RECT 84.420 30.050 84.680 30.370 ;
        RECT 83.960 28.350 84.220 28.670 ;
        RECT 84.480 25.610 84.620 30.050 ;
        RECT 84.870 27.815 85.150 28.185 ;
        RECT 84.940 26.630 85.080 27.815 ;
        RECT 84.880 26.310 85.140 26.630 ;
        RECT 84.420 25.290 84.680 25.610 ;
        RECT 83.040 23.250 83.300 23.570 ;
        RECT 80.740 20.870 81.000 21.190 ;
        RECT 82.580 20.870 82.840 21.190 ;
        RECT 84.940 20.170 85.080 26.310 ;
        RECT 85.860 25.270 86.000 31.410 ;
        RECT 85.800 24.950 86.060 25.270 ;
        RECT 86.320 23.910 86.460 36.170 ;
        RECT 87.240 34.110 87.380 36.170 ;
        RECT 87.180 33.790 87.440 34.110 ;
        RECT 87.240 31.050 87.380 33.790 ;
        RECT 87.630 31.895 87.910 32.265 ;
        RECT 86.720 30.730 86.980 31.050 ;
        RECT 87.180 30.730 87.440 31.050 ;
        RECT 86.260 23.590 86.520 23.910 ;
        RECT 86.780 21.190 86.920 30.730 ;
        RECT 87.700 21.190 87.840 31.895 ;
        RECT 88.160 30.710 88.300 46.370 ;
        RECT 88.100 30.390 88.360 30.710 ;
        RECT 86.720 20.870 86.980 21.190 ;
        RECT 87.640 20.870 87.900 21.190 ;
        RECT 42.100 19.850 42.360 20.170 ;
        RECT 50.380 19.850 50.640 20.170 ;
        RECT 52.680 19.850 52.940 20.170 ;
        RECT 75.680 19.850 75.940 20.170 ;
        RECT 76.140 19.850 76.400 20.170 ;
        RECT 76.600 19.850 76.860 20.170 ;
        RECT 79.820 19.850 80.080 20.170 ;
        RECT 80.280 19.850 80.540 20.170 ;
        RECT 84.880 19.850 85.140 20.170 ;
        RECT 30.950 18.635 32.490 19.005 ;
        RECT 42.160 11.940 42.300 19.850 ;
        RECT 45.320 19.510 45.580 19.830 ;
        RECT 54.980 19.510 55.240 19.830 ;
        RECT 45.380 11.940 45.520 19.510 ;
        RECT 48.540 19.170 48.800 19.490 ;
        RECT 51.760 19.170 52.020 19.490 ;
        RECT 48.600 11.940 48.740 19.170 ;
        RECT 51.820 11.940 51.960 19.170 ;
        RECT 55.040 11.940 55.180 19.510 ;
        RECT 71.080 19.170 71.340 19.490 ;
        RECT 74.300 19.170 74.560 19.490 ;
        RECT 77.520 19.170 77.780 19.490 ;
        RECT 71.140 11.940 71.280 19.170 ;
        RECT 74.360 11.940 74.500 19.170 ;
        RECT 77.580 11.940 77.720 19.170 ;
        RECT 42.090 7.940 42.370 11.940 ;
        RECT 45.310 7.940 45.590 11.940 ;
        RECT 48.530 7.940 48.810 11.940 ;
        RECT 51.750 7.940 52.030 11.940 ;
        RECT 54.970 7.940 55.250 11.940 ;
        RECT 71.070 7.940 71.350 11.940 ;
        RECT 74.290 7.940 74.570 11.940 ;
        RECT 77.510 7.940 77.790 11.940 ;
      LAYER met3 ;
        RECT 63.690 224.960 64.010 225.340 ;
        RECT 63.700 218.305 64.000 224.960 ;
        RECT 66.520 224.940 66.840 225.320 ;
        RECT 69.240 224.980 69.560 225.360 ;
        RECT 72.110 225.020 72.430 225.400 ;
        RECT 66.530 218.835 66.830 224.940 ;
        RECT 69.250 222.665 69.550 224.980 ;
        RECT 69.225 222.315 69.575 222.665 ;
        RECT 72.120 222.195 72.420 225.020 ;
        RECT 74.805 224.950 75.125 225.330 ;
        RECT 77.570 224.970 77.890 225.350 ;
        RECT 72.095 221.845 72.445 222.195 ;
        RECT 74.815 221.810 75.115 224.950 ;
        RECT 74.790 221.460 75.140 221.810 ;
        RECT 77.580 219.195 77.880 224.970 ;
        RECT 80.310 224.890 80.630 225.270 ;
        RECT 83.120 224.920 83.440 225.300 ;
        RECT 85.820 225.000 86.140 225.380 ;
        RECT 80.320 221.330 80.620 224.890 ;
        RECT 80.295 220.980 80.645 221.330 ;
        RECT 83.130 221.005 83.430 224.920 ;
        RECT 83.105 220.655 83.455 221.005 ;
        RECT 85.830 220.620 86.130 225.000 ;
        RECT 88.590 224.930 88.910 225.310 ;
        RECT 91.315 224.960 91.635 225.340 ;
        RECT 93.990 224.990 94.310 225.370 ;
        RECT 85.805 220.270 86.155 220.620 ;
        RECT 88.600 219.595 88.900 224.930 ;
        RECT 91.325 220.245 91.625 224.960 ;
        RECT 91.300 219.895 91.650 220.245 ;
        RECT 94.000 219.905 94.300 224.990 ;
        RECT 115.120 220.825 115.720 224.815 ;
        RECT 118.795 224.565 119.455 225.215 ;
        RECT 121.530 224.805 122.190 225.455 ;
        RECT 124.275 224.945 124.935 225.595 ;
        RECT 127.145 224.965 127.805 225.615 ;
        RECT 129.605 224.960 130.265 225.610 ;
        RECT 132.985 225.100 133.645 225.595 ;
        RECT 133.055 224.945 133.645 225.100 ;
        RECT 134.915 225.075 135.575 225.725 ;
        RECT 137.630 224.895 138.410 225.575 ;
        RECT 142.460 225.130 142.780 225.440 ;
        RECT 142.400 224.815 142.840 225.130 ;
        RECT 115.120 220.815 116.250 220.825 ;
        RECT 125.320 220.815 125.920 224.815 ;
        RECT 132.120 220.815 132.720 224.815 ;
        RECT 138.920 220.815 139.520 224.815 ;
        RECT 142.320 220.815 142.920 224.815 ;
        RECT 115.270 220.610 116.250 220.815 ;
        RECT 115.270 220.525 116.265 220.610 ;
        RECT 115.935 220.280 116.265 220.525 ;
        RECT 88.575 219.245 88.925 219.595 ;
        RECT 93.975 219.555 94.325 219.905 ;
        RECT 77.555 218.845 77.905 219.195 ;
        RECT 66.505 218.485 66.855 218.835 ;
        RECT 125.470 218.310 125.770 220.815 ;
        RECT 132.270 220.455 132.570 220.815 ;
        RECT 132.255 220.125 132.585 220.455 ;
        RECT 132.270 218.310 132.570 220.125 ;
        RECT 139.070 218.310 139.370 220.815 ;
        RECT 63.675 217.955 64.025 218.305 ;
        RECT 125.455 217.980 125.785 218.310 ;
        RECT 132.255 217.980 132.585 218.310 ;
        RECT 139.055 217.980 139.385 218.310 ;
        RECT 142.470 207.270 142.770 220.815 ;
        RECT 143.815 208.320 144.145 208.650 ;
        RECT 142.455 206.940 142.785 207.270 ;
        RECT 143.830 204.510 144.130 208.320 ;
        RECT 143.815 204.180 144.145 204.510 ;
        RECT 8.180 203.770 9.760 203.795 ;
        RECT 1.125 202.180 9.765 203.770 ;
        RECT 103.875 203.765 105.465 203.770 ;
        RECT 103.850 202.185 105.490 203.765 ;
        RECT 114.915 202.185 115.245 203.765 ;
        RECT 120.355 202.185 120.685 203.765 ;
        RECT 125.795 202.185 126.125 203.765 ;
        RECT 131.235 202.185 131.565 203.765 ;
        RECT 136.675 202.185 137.005 203.765 ;
        RECT 142.115 202.185 142.445 203.765 ;
        RECT 8.180 202.155 9.760 202.180 ;
        RECT 100.980 199.740 102.620 200.510 ;
        RECT 101.005 184.070 102.595 199.740 ;
        RECT 100.970 182.410 102.630 184.070 ;
        RECT 103.875 176.485 105.465 202.185 ;
        RECT 109.840 198.890 113.500 200.480 ;
        RECT 112.195 198.885 112.525 198.890 ;
        RECT 117.635 198.885 117.965 200.465 ;
        RECT 123.075 198.885 123.405 200.465 ;
        RECT 128.515 198.885 128.845 200.465 ;
        RECT 133.955 198.885 134.285 200.465 ;
        RECT 139.395 198.885 139.725 200.465 ;
        RECT 115.255 193.600 115.585 193.930 ;
        RECT 111.855 189.000 112.185 189.330 ;
        RECT 108.455 185.320 108.785 185.650 ;
        RECT 108.470 181.770 108.770 185.320 ;
        RECT 111.870 181.770 112.170 189.000 ;
        RECT 115.270 181.770 115.570 193.600 ;
        RECT 125.455 192.220 125.785 192.550 ;
        RECT 118.655 190.840 118.985 191.170 ;
        RECT 118.670 181.770 118.970 190.840 ;
        RECT 122.055 188.540 122.385 188.870 ;
        RECT 122.070 181.770 122.370 188.540 ;
        RECT 125.470 181.770 125.770 192.220 ;
        RECT 143.830 191.170 144.130 204.180 ;
        RECT 147.555 202.185 147.885 203.765 ;
        RECT 144.835 198.885 145.165 200.465 ;
        RECT 148.095 195.430 148.445 195.780 ;
        RECT 143.815 190.840 144.145 191.170 ;
        RECT 128.855 189.920 129.185 190.250 ;
        RECT 128.870 181.770 129.170 189.920 ;
        RECT 135.655 187.160 135.985 187.490 ;
        RECT 132.255 184.860 132.585 185.190 ;
        RECT 132.270 181.770 132.570 184.860 ;
        RECT 135.670 181.770 135.970 187.160 ;
        RECT 145.855 186.240 146.185 186.570 ;
        RECT 139.055 184.860 139.385 185.190 ;
        RECT 142.455 184.860 142.785 185.190 ;
        RECT 139.070 181.770 139.370 184.860 ;
        RECT 142.470 181.770 142.770 184.860 ;
        RECT 145.870 181.770 146.170 186.240 ;
        RECT 108.320 177.770 108.920 181.770 ;
        RECT 111.720 177.770 112.320 181.770 ;
        RECT 115.120 177.770 115.720 181.770 ;
        RECT 118.520 177.770 119.120 181.770 ;
        RECT 121.920 177.770 122.520 181.770 ;
        RECT 125.320 177.770 125.920 181.770 ;
        RECT 128.720 177.770 129.320 181.770 ;
        RECT 132.120 177.770 132.720 181.770 ;
        RECT 135.520 177.770 136.120 181.770 ;
        RECT 138.920 177.770 139.520 181.770 ;
        RECT 142.320 177.770 142.920 181.770 ;
        RECT 145.720 177.770 146.320 181.770 ;
        RECT 111.850 177.430 112.190 177.770 ;
        RECT 111.855 177.355 112.185 177.430 ;
        RECT 139.070 176.850 139.370 177.770 ;
        RECT 142.450 177.440 142.790 177.770 ;
        RECT 142.455 177.255 142.785 177.440 ;
        RECT 148.120 177.395 148.420 195.430 ;
        RECT 149.255 187.620 149.585 187.950 ;
        RECT 149.270 181.770 149.570 187.620 ;
        RECT 152.655 184.860 152.985 185.190 ;
        RECT 152.670 181.770 152.970 184.860 ;
        RECT 149.120 177.770 149.720 181.770 ;
        RECT 152.520 177.770 153.120 181.770 ;
        RECT 149.255 177.725 149.585 177.770 ;
        RECT 148.105 177.065 148.435 177.395 ;
        RECT 144.655 176.850 144.985 176.865 ;
        RECT 117.980 176.485 118.880 176.640 ;
        RECT 137.800 176.485 138.700 176.620 ;
        RECT 139.070 176.550 144.985 176.850 ;
        RECT 144.655 176.535 144.985 176.550 ;
        RECT 103.865 176.250 138.700 176.485 ;
        RECT 157.570 176.250 158.470 176.600 ;
        RECT 103.865 176.230 144.350 176.250 ;
        RECT 145.300 176.230 158.470 176.250 ;
        RECT 103.865 175.110 158.470 176.230 ;
        RECT 103.865 174.875 138.700 175.110 ;
        RECT 117.980 174.620 118.880 174.875 ;
        RECT 137.800 174.600 138.700 174.875 ;
        RECT 157.570 174.580 158.470 175.110 ;
        RECT 27.630 173.695 29.210 174.025 ;
        RECT 70.585 172.310 70.915 172.325 ;
        RECT 83.005 172.310 83.335 172.325 ;
        RECT 70.585 172.010 83.335 172.310 ;
        RECT 70.585 171.995 70.915 172.010 ;
        RECT 83.005 171.995 83.335 172.010 ;
        RECT 69.205 171.630 69.535 171.645 ;
        RECT 85.765 171.630 86.095 171.645 ;
        RECT 69.205 171.330 86.095 171.630 ;
        RECT 69.205 171.315 69.535 171.330 ;
        RECT 85.765 171.315 86.095 171.330 ;
        RECT 30.930 170.975 32.510 171.305 ;
        RECT 78.405 169.590 78.735 169.605 ;
        RECT 79.325 169.590 79.655 169.605 ;
        RECT 81.165 169.590 81.495 169.605 ;
        RECT 78.405 169.290 81.495 169.590 ;
        RECT 108.820 169.350 109.400 169.400 ;
        RECT 128.680 169.350 129.260 169.390 ;
        RECT 148.880 169.350 149.460 169.370 ;
        RECT 78.405 169.275 78.735 169.290 ;
        RECT 79.325 169.275 79.655 169.290 ;
        RECT 81.165 169.275 81.495 169.290 ;
        RECT 66.445 168.910 66.775 168.925 ;
        RECT 84.845 168.910 85.175 168.925 ;
        RECT 87.145 168.910 87.475 168.925 ;
        RECT 66.445 168.610 87.475 168.910 ;
        RECT 108.800 168.720 149.480 169.350 ;
        RECT 66.445 168.595 66.775 168.610 ;
        RECT 84.845 168.595 85.175 168.610 ;
        RECT 87.145 168.595 87.475 168.610 ;
        RECT 27.630 168.255 29.210 168.585 ;
        RECT 84.385 168.230 84.715 168.245 ;
        RECT 68.530 167.930 84.715 168.230 ;
        RECT 41.605 167.550 41.935 167.565 ;
        RECT 47.330 167.550 47.710 167.560 ;
        RECT 41.605 167.250 47.710 167.550 ;
        RECT 41.605 167.235 41.935 167.250 ;
        RECT 47.330 167.240 47.710 167.250 ;
        RECT 65.065 167.550 65.395 167.565 ;
        RECT 68.530 167.550 68.830 167.930 ;
        RECT 84.385 167.915 84.715 167.930 ;
        RECT 65.065 167.250 68.830 167.550 ;
        RECT 75.645 167.560 75.975 167.565 ;
        RECT 75.645 167.550 76.230 167.560 ;
        RECT 77.945 167.550 78.275 167.565 ;
        RECT 79.325 167.550 79.655 167.565 ;
        RECT 75.645 167.250 76.430 167.550 ;
        RECT 77.945 167.250 79.655 167.550 ;
        RECT 65.065 167.235 65.395 167.250 ;
        RECT 75.645 167.240 76.230 167.250 ;
        RECT 75.645 167.235 75.975 167.240 ;
        RECT 77.945 167.235 78.275 167.250 ;
        RECT 79.325 167.235 79.655 167.250 ;
        RECT 42.525 166.870 42.855 166.885 ;
        RECT 45.490 166.870 45.870 166.880 ;
        RECT 42.525 166.570 45.870 166.870 ;
        RECT 42.525 166.555 42.855 166.570 ;
        RECT 45.490 166.560 45.870 166.570 ;
        RECT 30.930 165.535 32.510 165.865 ;
        RECT 74.010 165.510 74.390 165.520 ;
        RECT 74.725 165.510 75.055 165.525 ;
        RECT 74.010 165.210 75.055 165.510 ;
        RECT 74.010 165.200 74.390 165.210 ;
        RECT 74.725 165.195 75.055 165.210 ;
        RECT 6.580 164.840 10.580 164.980 ;
        RECT 6.580 164.520 10.910 164.840 ;
        RECT 88.065 164.830 88.395 164.845 ;
        RECT 91.525 164.830 95.525 164.980 ;
        RECT 88.065 164.530 95.525 164.830 ;
        RECT 6.580 164.380 10.580 164.520 ;
        RECT 88.065 164.515 88.395 164.530 ;
        RECT 91.525 164.380 95.525 164.530 ;
        RECT 27.630 162.815 29.210 163.145 ;
        RECT 59.085 161.430 59.415 161.445 ;
        RECT 91.525 161.430 95.525 161.580 ;
        RECT 59.085 161.130 95.525 161.430 ;
        RECT 59.085 161.115 59.415 161.130 ;
        RECT 91.525 160.980 95.525 161.130 ;
        RECT 77.690 160.750 78.070 160.760 ;
        RECT 83.465 160.750 83.795 160.765 ;
        RECT 77.690 160.450 83.795 160.750 ;
        RECT 77.690 160.440 78.070 160.450 ;
        RECT 83.465 160.435 83.795 160.450 ;
        RECT 30.930 160.095 32.510 160.425 ;
        RECT 60.465 160.080 60.795 160.085 ;
        RECT 60.210 160.070 60.795 160.080 ;
        RECT 60.010 159.770 82.630 160.070 ;
        RECT 60.210 159.760 60.795 159.770 ;
        RECT 60.465 159.755 60.795 159.760 ;
        RECT 82.330 159.390 82.630 159.770 ;
        RECT 86.225 159.390 86.555 159.405 ;
        RECT 82.330 159.090 86.555 159.390 ;
        RECT 86.225 159.075 86.555 159.090 ;
        RECT 7.105 158.710 7.435 158.725 ;
        RECT 77.025 158.720 77.355 158.725 ;
        RECT 10.530 158.710 10.910 158.720 ;
        RECT 7.105 158.410 10.910 158.710 ;
        RECT 7.105 158.395 7.435 158.410 ;
        RECT 10.530 158.400 10.910 158.410 ;
        RECT 76.770 158.710 77.355 158.720 ;
        RECT 76.770 158.410 77.580 158.710 ;
        RECT 76.770 158.400 77.355 158.410 ;
        RECT 77.025 158.395 77.355 158.400 ;
        RECT 83.465 158.030 83.795 158.045 ;
        RECT 91.525 158.030 95.525 158.180 ;
        RECT 83.465 157.730 95.525 158.030 ;
        RECT 83.465 157.715 83.795 157.730 ;
        RECT 27.630 157.375 29.210 157.705 ;
        RECT 91.525 157.580 95.525 157.730 ;
        RECT 41.145 156.670 41.475 156.685 ;
        RECT 42.985 156.670 43.315 156.685 ;
        RECT 47.125 156.670 47.455 156.685 ;
        RECT 41.145 156.370 47.455 156.670 ;
        RECT 41.145 156.355 41.475 156.370 ;
        RECT 42.985 156.355 43.315 156.370 ;
        RECT 47.125 156.355 47.455 156.370 ;
        RECT 64.605 155.310 64.935 155.325 ;
        RECT 66.650 155.310 67.030 155.320 ;
        RECT 64.605 155.010 67.030 155.310 ;
        RECT 64.605 154.995 64.935 155.010 ;
        RECT 66.650 155.000 67.030 155.010 ;
        RECT 30.930 154.655 32.510 154.985 ;
        RECT 88.065 154.630 88.395 154.645 ;
        RECT 91.525 154.630 95.525 154.780 ;
        RECT 88.065 154.330 95.525 154.630 ;
        RECT 128.680 154.340 129.260 154.430 ;
        RECT 139.065 154.340 139.695 168.720 ;
        RECT 88.065 154.315 88.395 154.330 ;
        RECT 91.525 154.180 95.525 154.330 ;
        RECT 53.770 153.950 54.150 153.960 ;
        RECT 86.225 153.950 86.555 153.965 ;
        RECT 53.770 153.650 86.555 153.950 ;
        RECT 108.740 153.710 149.500 154.340 ;
        RECT 108.790 153.690 109.370 153.710 ;
        RECT 53.770 153.640 54.150 153.650 ;
        RECT 86.225 153.635 86.555 153.650 ;
        RECT 65.730 153.270 66.110 153.280 ;
        RECT 81.625 153.270 81.955 153.285 ;
        RECT 65.730 152.970 81.955 153.270 ;
        RECT 65.730 152.960 66.110 152.970 ;
        RECT 81.625 152.955 81.955 152.970 ;
        RECT 27.630 151.935 29.210 152.265 ;
        RECT 62.765 151.230 63.095 151.245 ;
        RECT 91.525 151.230 95.525 151.380 ;
        RECT 62.765 150.930 95.525 151.230 ;
        RECT 62.765 150.915 63.095 150.930 ;
        RECT 91.525 150.780 95.525 150.930 ;
        RECT 30.930 149.215 32.510 149.545 ;
        RECT 83.465 147.830 83.795 147.845 ;
        RECT 91.525 147.830 95.525 147.980 ;
        RECT 83.465 147.530 95.525 147.830 ;
        RECT 83.465 147.515 83.795 147.530 ;
        RECT 91.525 147.380 95.525 147.530 ;
        RECT 27.630 146.495 29.210 146.825 ;
        RECT 69.410 146.470 69.790 146.480 ;
        RECT 71.505 146.470 71.835 146.485 ;
        RECT 69.410 146.170 71.835 146.470 ;
        RECT 69.410 146.160 69.790 146.170 ;
        RECT 71.505 146.155 71.835 146.170 ;
        RECT 75.850 144.430 76.230 144.440 ;
        RECT 91.525 144.430 95.525 144.580 ;
        RECT 75.850 144.130 95.525 144.430 ;
        RECT 75.850 144.120 76.230 144.130 ;
        RECT 30.930 143.775 32.510 144.105 ;
        RECT 91.525 143.980 95.525 144.130 ;
        RECT 20.445 143.070 20.775 143.085 ;
        RECT 30.565 143.070 30.895 143.085 ;
        RECT 36.085 143.070 36.415 143.085 ;
        RECT 20.445 142.770 36.415 143.070 ;
        RECT 20.445 142.755 20.775 142.770 ;
        RECT 30.565 142.755 30.895 142.770 ;
        RECT 36.085 142.755 36.415 142.770 ;
        RECT 20.905 142.390 21.235 142.405 ;
        RECT 31.945 142.390 32.275 142.405 ;
        RECT 73.805 142.400 74.135 142.405 ;
        RECT 73.805 142.390 74.390 142.400 ;
        RECT 20.905 142.090 32.275 142.390 ;
        RECT 73.580 142.090 74.390 142.390 ;
        RECT 20.905 142.075 21.235 142.090 ;
        RECT 31.945 142.075 32.275 142.090 ;
        RECT 73.805 142.080 74.390 142.090 ;
        RECT 73.805 142.075 74.135 142.080 ;
        RECT 21.825 141.710 22.155 141.725 ;
        RECT 24.125 141.710 24.455 141.725 ;
        RECT 21.825 141.410 24.455 141.710 ;
        RECT 21.825 141.395 22.155 141.410 ;
        RECT 24.125 141.395 24.455 141.410 ;
        RECT 27.630 141.055 29.210 141.385 ;
        RECT 61.845 141.030 62.175 141.045 ;
        RECT 91.525 141.030 95.525 141.180 ;
        RECT 61.845 140.730 95.525 141.030 ;
        RECT 61.845 140.715 62.175 140.730 ;
        RECT 91.525 140.580 95.525 140.730 ;
        RECT 19.525 140.350 19.855 140.365 ;
        RECT 20.445 140.350 20.775 140.365 ;
        RECT 19.525 140.050 20.775 140.350 ;
        RECT 19.525 140.035 19.855 140.050 ;
        RECT 20.445 140.035 20.775 140.050 ;
        RECT 70.585 140.350 70.915 140.365 ;
        RECT 77.690 140.350 78.070 140.360 ;
        RECT 70.585 140.050 78.070 140.350 ;
        RECT 70.585 140.035 70.915 140.050 ;
        RECT 77.690 140.040 78.070 140.050 ;
        RECT 65.525 139.670 65.855 139.685 ;
        RECT 68.745 139.670 69.075 139.685 ;
        RECT 75.645 139.670 75.975 139.685 ;
        RECT 65.525 139.370 75.975 139.670 ;
        RECT 65.525 139.355 65.855 139.370 ;
        RECT 68.745 139.355 69.075 139.370 ;
        RECT 75.645 139.355 75.975 139.370 ;
        RECT 80.450 139.670 80.830 139.680 ;
        RECT 85.765 139.670 86.095 139.685 ;
        RECT 80.450 139.370 86.095 139.670 ;
        RECT 80.450 139.360 80.830 139.370 ;
        RECT 85.765 139.355 86.095 139.370 ;
        RECT 108.790 139.340 109.370 139.370 ;
        RECT 128.680 139.340 129.260 139.360 ;
        RECT 139.065 139.340 139.695 153.710 ;
        RECT 108.790 138.740 149.490 139.340 ;
        RECT 108.810 138.710 149.490 138.740 ;
        RECT 30.930 138.335 32.510 138.665 ;
        RECT 87.605 137.630 87.935 137.645 ;
        RECT 91.525 137.630 95.525 137.780 ;
        RECT 87.605 137.330 95.525 137.630 ;
        RECT 87.605 137.315 87.935 137.330 ;
        RECT 91.525 137.180 95.525 137.330 ;
        RECT 27.630 135.615 29.210 135.945 ;
        RECT 44.825 135.590 45.155 135.605 ;
        RECT 47.125 135.600 47.455 135.605 ;
        RECT 45.490 135.590 45.870 135.600 ;
        RECT 47.125 135.590 47.710 135.600 ;
        RECT 44.825 135.290 45.870 135.590 ;
        RECT 46.900 135.290 47.710 135.590 ;
        RECT 44.825 135.275 45.155 135.290 ;
        RECT 45.490 135.280 45.870 135.290 ;
        RECT 47.125 135.280 47.710 135.290 ;
        RECT 47.125 135.275 47.455 135.280 ;
        RECT 10.785 134.910 11.115 134.925 ;
        RECT 10.570 134.595 11.115 134.910 ;
        RECT 79.530 134.910 79.910 134.920 ;
        RECT 84.385 134.910 84.715 134.925 ;
        RECT 79.530 134.610 84.715 134.910 ;
        RECT 79.530 134.600 79.910 134.610 ;
        RECT 84.385 134.595 84.715 134.610 ;
        RECT 10.570 134.380 10.870 134.595 ;
        RECT 6.580 133.930 10.870 134.380 ;
        RECT 76.105 134.230 76.435 134.245 ;
        RECT 91.525 134.230 95.525 134.380 ;
        RECT 76.105 133.930 95.525 134.230 ;
        RECT 6.580 133.780 10.580 133.930 ;
        RECT 76.105 133.915 76.435 133.930 ;
        RECT 91.525 133.780 95.525 133.930 ;
        RECT 30.930 132.895 32.510 133.225 ;
        RECT 61.385 132.880 61.715 132.885 ;
        RECT 61.130 132.870 61.715 132.880 ;
        RECT 60.930 132.570 61.715 132.870 ;
        RECT 61.130 132.560 61.715 132.570 ;
        RECT 67.570 132.870 67.950 132.880 ;
        RECT 76.770 132.870 77.150 132.880 ;
        RECT 67.570 132.570 77.150 132.870 ;
        RECT 67.570 132.560 67.950 132.570 ;
        RECT 76.770 132.560 77.150 132.570 ;
        RECT 61.385 132.555 61.715 132.560 ;
        RECT 67.365 130.830 67.695 130.845 ;
        RECT 91.525 130.830 95.525 130.980 ;
        RECT 67.365 130.530 95.525 130.830 ;
        RECT 67.365 130.515 67.695 130.530 ;
        RECT 27.630 130.175 29.210 130.505 ;
        RECT 91.525 130.380 95.525 130.530 ;
        RECT 79.785 130.150 80.115 130.165 ;
        RECT 82.085 130.150 82.415 130.165 ;
        RECT 79.785 129.850 82.415 130.150 ;
        RECT 79.785 129.835 80.115 129.850 ;
        RECT 82.085 129.835 82.415 129.850 ;
        RECT 26.425 129.480 26.755 129.485 ;
        RECT 26.170 129.470 26.755 129.480 ;
        RECT 25.970 129.170 26.755 129.470 ;
        RECT 26.170 129.160 26.755 129.170 ;
        RECT 26.425 129.155 26.755 129.160 ;
        RECT 22.490 128.790 22.870 128.800 ;
        RECT 23.665 128.790 23.995 128.805 ;
        RECT 22.490 128.490 23.995 128.790 ;
        RECT 22.490 128.480 22.870 128.490 ;
        RECT 23.665 128.475 23.995 128.490 ;
        RECT 66.445 128.790 66.775 128.805 ;
        RECT 67.365 128.790 67.695 128.805 ;
        RECT 66.445 128.490 67.695 128.790 ;
        RECT 66.445 128.475 66.775 128.490 ;
        RECT 67.365 128.475 67.695 128.490 ;
        RECT 30.930 127.455 32.510 127.785 ;
        RECT 82.545 127.430 82.875 127.445 ;
        RECT 91.525 127.430 95.525 127.580 ;
        RECT 82.545 127.130 95.525 127.430 ;
        RECT 82.545 127.115 82.875 127.130 ;
        RECT 91.525 126.980 95.525 127.130 ;
        RECT 70.585 126.070 70.915 126.085 ;
        RECT 71.250 126.070 71.630 126.080 ;
        RECT 70.585 125.770 71.630 126.070 ;
        RECT 70.585 125.755 70.915 125.770 ;
        RECT 71.250 125.760 71.630 125.770 ;
        RECT 62.765 125.390 63.095 125.405 ;
        RECT 65.065 125.390 65.395 125.405 ;
        RECT 62.765 125.090 65.395 125.390 ;
        RECT 62.765 125.075 63.095 125.090 ;
        RECT 65.065 125.075 65.395 125.090 ;
        RECT 27.630 124.735 29.210 125.065 ;
        RECT 58.165 124.710 58.495 124.725 ;
        RECT 65.525 124.710 65.855 124.725 ;
        RECT 75.645 124.710 75.975 124.725 ;
        RECT 58.165 124.410 75.975 124.710 ;
        RECT 58.165 124.395 58.495 124.410 ;
        RECT 65.525 124.395 65.855 124.410 ;
        RECT 75.645 124.395 75.975 124.410 ;
        RECT 128.610 124.380 129.190 124.420 ;
        RECT 139.065 124.380 139.695 138.710 ;
        RECT 148.830 138.670 149.410 138.710 ;
        RECT 108.800 124.370 149.530 124.380 ;
        RECT 78.865 124.030 79.195 124.045 ;
        RECT 80.450 124.030 80.830 124.040 ;
        RECT 78.865 123.730 80.830 124.030 ;
        RECT 78.865 123.715 79.195 123.730 ;
        RECT 80.450 123.720 80.830 123.730 ;
        RECT 82.545 124.030 82.875 124.045 ;
        RECT 91.525 124.030 95.525 124.180 ;
        RECT 82.545 123.730 95.525 124.030 ;
        RECT 108.790 123.750 149.530 124.370 ;
        RECT 108.790 123.740 109.370 123.750 ;
        RECT 82.545 123.715 82.875 123.730 ;
        RECT 91.525 123.580 95.525 123.730 ;
        RECT 51.930 123.350 52.310 123.360 ;
        RECT 54.025 123.350 54.355 123.365 ;
        RECT 51.930 123.050 54.355 123.350 ;
        RECT 51.930 123.040 52.310 123.050 ;
        RECT 54.025 123.035 54.355 123.050 ;
        RECT 64.810 123.350 65.190 123.360 ;
        RECT 67.825 123.350 68.155 123.365 ;
        RECT 64.810 123.050 68.155 123.350 ;
        RECT 64.810 123.040 65.190 123.050 ;
        RECT 67.825 123.035 68.155 123.050 ;
        RECT 67.365 122.670 67.695 122.685 ;
        RECT 69.205 122.670 69.535 122.685 ;
        RECT 67.365 122.370 69.535 122.670 ;
        RECT 67.365 122.355 67.695 122.370 ;
        RECT 69.205 122.355 69.535 122.370 ;
        RECT 30.930 122.015 32.510 122.345 ;
        RECT 63.890 121.990 64.270 122.000 ;
        RECT 66.905 121.990 67.235 122.005 ;
        RECT 63.890 121.690 67.235 121.990 ;
        RECT 63.890 121.680 64.270 121.690 ;
        RECT 66.905 121.675 67.235 121.690 ;
        RECT 83.005 120.630 83.335 120.645 ;
        RECT 91.525 120.630 95.525 120.780 ;
        RECT 83.005 120.330 95.525 120.630 ;
        RECT 83.005 120.315 83.335 120.330 ;
        RECT 91.525 120.180 95.525 120.330 ;
        RECT 27.630 119.295 29.210 119.625 ;
        RECT 54.945 119.270 55.275 119.285 ;
        RECT 68.745 119.270 69.075 119.285 ;
        RECT 54.945 118.970 69.075 119.270 ;
        RECT 54.945 118.955 55.275 118.970 ;
        RECT 68.745 118.955 69.075 118.970 ;
        RECT 65.730 118.590 66.110 118.600 ;
        RECT 80.450 118.590 80.830 118.600 ;
        RECT 65.730 118.290 80.830 118.590 ;
        RECT 65.730 118.280 66.110 118.290 ;
        RECT 80.450 118.280 80.830 118.290 ;
        RECT 71.505 117.910 71.835 117.925 ;
        RECT 72.170 117.910 72.550 117.920 ;
        RECT 71.505 117.610 72.550 117.910 ;
        RECT 71.505 117.595 71.835 117.610 ;
        RECT 72.170 117.600 72.550 117.610 ;
        RECT 85.765 117.230 86.095 117.245 ;
        RECT 91.525 117.230 95.525 117.380 ;
        RECT 85.765 116.930 95.525 117.230 ;
        RECT 85.765 116.915 86.095 116.930 ;
        RECT 30.930 116.575 32.510 116.905 ;
        RECT 91.525 116.780 95.525 116.930 ;
        RECT 66.650 115.190 67.030 115.200 ;
        RECT 74.010 115.190 74.390 115.200 ;
        RECT 66.650 114.890 74.390 115.190 ;
        RECT 66.650 114.880 67.030 114.890 ;
        RECT 74.010 114.880 74.390 114.890 ;
        RECT 10.785 114.510 11.115 114.525 ;
        RECT 10.570 114.195 11.115 114.510 ;
        RECT 10.570 113.980 10.870 114.195 ;
        RECT 6.580 113.530 10.870 113.980 ;
        RECT 27.630 113.855 29.210 114.185 ;
        RECT 68.285 113.830 68.615 113.845 ;
        RECT 69.410 113.830 69.790 113.840 ;
        RECT 68.285 113.530 69.790 113.830 ;
        RECT 6.580 113.380 10.580 113.530 ;
        RECT 68.285 113.515 68.615 113.530 ;
        RECT 69.410 113.520 69.790 113.530 ;
        RECT 87.605 113.830 87.935 113.845 ;
        RECT 91.525 113.830 95.525 113.980 ;
        RECT 87.605 113.530 95.525 113.830 ;
        RECT 87.605 113.515 87.935 113.530 ;
        RECT 91.525 113.380 95.525 113.530 ;
        RECT 17.685 112.470 18.015 112.485 ;
        RECT 20.905 112.470 21.235 112.485 ;
        RECT 17.685 112.170 21.235 112.470 ;
        RECT 17.685 112.155 18.015 112.170 ;
        RECT 20.905 112.155 21.235 112.170 ;
        RECT 52.850 111.790 53.230 111.800 ;
        RECT 53.565 111.790 53.895 111.805 ;
        RECT 52.850 111.490 53.895 111.790 ;
        RECT 52.850 111.480 53.230 111.490 ;
        RECT 53.565 111.475 53.895 111.490 ;
        RECT 30.930 111.135 32.510 111.465 ;
        RECT 26.170 111.110 26.550 111.120 ;
        RECT 27.345 111.110 27.675 111.125 ;
        RECT 26.170 110.810 27.675 111.110 ;
        RECT 26.170 110.800 26.550 110.810 ;
        RECT 27.345 110.795 27.675 110.810 ;
        RECT 80.705 111.110 81.035 111.125 ;
        RECT 86.685 111.110 87.015 111.125 ;
        RECT 80.705 110.810 87.015 111.110 ;
        RECT 80.705 110.795 81.035 110.810 ;
        RECT 86.685 110.795 87.015 110.810 ;
        RECT 88.065 110.430 88.395 110.445 ;
        RECT 91.525 110.430 95.525 110.580 ;
        RECT 88.065 110.130 95.525 110.430 ;
        RECT 88.065 110.115 88.395 110.130 ;
        RECT 91.525 109.980 95.525 110.130 ;
        RECT 128.730 109.330 129.310 109.390 ;
        RECT 139.065 109.330 139.695 123.750 ;
        RECT 148.910 109.330 149.490 109.420 ;
        RECT 108.740 108.790 149.490 109.330 ;
        RECT 27.630 108.415 29.210 108.745 ;
        RECT 108.740 108.700 149.420 108.790 ;
        RECT 84.845 107.710 85.175 107.725 ;
        RECT 88.525 107.710 88.855 107.725 ;
        RECT 84.845 107.410 88.855 107.710 ;
        RECT 84.845 107.395 85.175 107.410 ;
        RECT 88.525 107.395 88.855 107.410 ;
        RECT 32.405 107.030 32.735 107.045 ;
        RECT 33.325 107.030 33.655 107.045 ;
        RECT 32.405 106.730 33.655 107.030 ;
        RECT 32.405 106.715 32.735 106.730 ;
        RECT 33.325 106.715 33.655 106.730 ;
        RECT 82.545 107.030 82.875 107.045 ;
        RECT 91.525 107.030 95.525 107.180 ;
        RECT 82.545 106.730 95.525 107.030 ;
        RECT 82.545 106.715 82.875 106.730 ;
        RECT 91.525 106.580 95.525 106.730 ;
        RECT 30.930 105.695 32.510 106.025 ;
        RECT 32.405 104.990 32.735 105.005 ;
        RECT 36.545 104.990 36.875 105.005 ;
        RECT 67.365 105.000 67.695 105.005 ;
        RECT 67.365 104.990 67.950 105.000 ;
        RECT 32.405 104.690 36.875 104.990 ;
        RECT 67.140 104.690 67.950 104.990 ;
        RECT 32.405 104.675 32.735 104.690 ;
        RECT 36.545 104.675 36.875 104.690 ;
        RECT 67.365 104.680 67.950 104.690 ;
        RECT 78.405 104.990 78.735 105.005 ;
        RECT 84.845 104.990 85.175 105.005 ;
        RECT 78.405 104.690 85.175 104.990 ;
        RECT 67.365 104.675 67.695 104.680 ;
        RECT 78.405 104.675 78.735 104.690 ;
        RECT 84.845 104.675 85.175 104.690 ;
        RECT 26.170 104.310 26.550 104.320 ;
        RECT 27.805 104.310 28.135 104.325 ;
        RECT 26.170 104.010 28.135 104.310 ;
        RECT 26.170 104.000 26.550 104.010 ;
        RECT 27.805 103.995 28.135 104.010 ;
        RECT 77.485 103.630 77.815 103.645 ;
        RECT 91.525 103.630 95.525 103.780 ;
        RECT 77.485 103.330 95.525 103.630 ;
        RECT 77.485 103.315 77.815 103.330 ;
        RECT 27.630 102.975 29.210 103.305 ;
        RECT 91.525 103.180 95.525 103.330 ;
        RECT 139.065 102.305 139.695 108.700 ;
        RECT 83.465 102.280 83.795 102.285 ;
        RECT 83.210 102.270 83.795 102.280 ;
        RECT 83.010 101.970 83.795 102.270 ;
        RECT 83.210 101.960 83.795 101.970 ;
        RECT 83.465 101.955 83.795 101.960 ;
        RECT 139.065 101.675 158.365 102.305 ;
        RECT 74.930 101.590 75.310 101.600 ;
        RECT 88.065 101.590 88.395 101.605 ;
        RECT 74.930 101.290 88.395 101.590 ;
        RECT 74.930 101.280 75.310 101.290 ;
        RECT 88.065 101.275 88.395 101.290 ;
        RECT 30.930 100.255 32.510 100.585 ;
        RECT 71.965 100.230 72.295 100.245 ;
        RECT 91.525 100.230 95.525 100.380 ;
        RECT 71.965 99.930 95.525 100.230 ;
        RECT 71.965 99.915 72.295 99.930 ;
        RECT 91.525 99.780 95.525 99.930 ;
        RECT 27.630 97.535 29.210 97.865 ;
        RECT 62.765 97.510 63.095 97.525 ;
        RECT 72.170 97.510 72.550 97.520 ;
        RECT 62.765 97.210 72.550 97.510 ;
        RECT 62.765 97.195 63.095 97.210 ;
        RECT 72.170 97.200 72.550 97.210 ;
        RECT 60.210 96.830 60.590 96.840 ;
        RECT 88.065 96.830 88.395 96.845 ;
        RECT 91.525 96.830 95.525 96.980 ;
        RECT 60.210 96.530 88.395 96.830 ;
        RECT 60.210 96.520 60.590 96.530 ;
        RECT 88.065 96.515 88.395 96.530 ;
        RECT 88.770 96.530 95.525 96.830 ;
        RECT 157.735 96.565 158.365 101.675 ;
        RECT 18.605 96.150 18.935 96.165 ;
        RECT 25.965 96.150 26.295 96.165 ;
        RECT 18.605 95.850 26.295 96.150 ;
        RECT 18.605 95.835 18.935 95.850 ;
        RECT 25.965 95.835 26.295 95.850 ;
        RECT 75.645 96.150 75.975 96.165 ;
        RECT 88.770 96.150 89.070 96.530 ;
        RECT 91.525 96.380 95.525 96.530 ;
        RECT 75.645 95.850 89.070 96.150 ;
        RECT 75.645 95.835 75.975 95.850 ;
        RECT 30.930 94.815 32.510 95.145 ;
        RECT 22.285 94.120 22.615 94.125 ;
        RECT 22.285 94.110 22.870 94.120 ;
        RECT 80.705 94.110 81.035 94.125 ;
        RECT 82.085 94.110 82.415 94.125 ;
        RECT 22.060 93.810 22.870 94.110 ;
        RECT 22.285 93.800 22.870 93.810 ;
        RECT 80.490 93.810 82.415 94.110 ;
        RECT 22.285 93.795 22.615 93.800 ;
        RECT 80.490 93.795 81.035 93.810 ;
        RECT 82.085 93.795 82.415 93.810 ;
        RECT 79.785 93.430 80.115 93.445 ;
        RECT 80.490 93.430 80.790 93.795 ;
        RECT 79.785 93.130 80.790 93.430 ;
        RECT 82.545 93.430 82.875 93.445 ;
        RECT 91.525 93.430 95.525 93.580 ;
        RECT 82.545 93.130 95.525 93.430 ;
        RECT 79.785 93.115 80.115 93.130 ;
        RECT 82.545 93.115 82.875 93.130 ;
        RECT 91.525 92.980 95.525 93.130 ;
        RECT 27.630 92.095 29.210 92.425 ;
        RECT 77.690 92.070 78.070 92.080 ;
        RECT 84.385 92.070 84.715 92.085 ;
        RECT 77.690 91.770 84.715 92.070 ;
        RECT 77.690 91.760 78.070 91.770 ;
        RECT 84.385 91.755 84.715 91.770 ;
        RECT 61.130 91.390 61.510 91.400 ;
        RECT 64.145 91.390 64.475 91.405 ;
        RECT 61.130 91.090 64.475 91.390 ;
        RECT 61.130 91.080 61.510 91.090 ;
        RECT 64.145 91.075 64.475 91.090 ;
        RECT 81.370 91.390 81.750 91.400 ;
        RECT 85.305 91.390 85.635 91.405 ;
        RECT 81.370 91.090 85.635 91.390 ;
        RECT 81.370 91.080 81.750 91.090 ;
        RECT 85.305 91.075 85.635 91.090 ;
        RECT 53.105 90.720 53.435 90.725 ;
        RECT 52.850 90.710 53.435 90.720 ;
        RECT 52.650 90.410 53.435 90.710 ;
        RECT 52.850 90.400 53.435 90.410 ;
        RECT 53.105 90.395 53.435 90.400 ;
        RECT 76.565 90.710 76.895 90.725 ;
        RECT 78.865 90.710 79.195 90.725 ;
        RECT 80.245 90.710 80.575 90.725 ;
        RECT 76.565 90.410 80.575 90.710 ;
        RECT 76.565 90.395 76.895 90.410 ;
        RECT 78.865 90.395 79.195 90.410 ;
        RECT 80.245 90.395 80.575 90.410 ;
        RECT 82.545 90.030 82.875 90.045 ;
        RECT 91.525 90.030 95.525 90.180 ;
        RECT 82.545 89.730 95.525 90.030 ;
        RECT 82.545 89.715 82.875 89.730 ;
        RECT 30.930 89.375 32.510 89.705 ;
        RECT 91.525 89.580 95.525 89.730 ;
        RECT 72.885 89.350 73.215 89.365 ;
        RECT 82.085 89.350 82.415 89.365 ;
        RECT 85.305 89.350 85.635 89.365 ;
        RECT 72.885 89.050 85.635 89.350 ;
        RECT 72.885 89.035 73.215 89.050 ;
        RECT 82.085 89.035 82.415 89.050 ;
        RECT 85.305 89.035 85.635 89.050 ;
        RECT 54.485 88.670 54.815 88.685 ;
        RECT 56.785 88.670 57.115 88.685 ;
        RECT 54.485 88.370 57.115 88.670 ;
        RECT 54.485 88.355 54.815 88.370 ;
        RECT 56.570 88.355 57.115 88.370 ;
        RECT 27.630 86.655 29.210 86.985 ;
        RECT 20.905 86.630 21.235 86.645 ;
        RECT 22.490 86.630 22.870 86.640 ;
        RECT 20.905 86.330 22.870 86.630 ;
        RECT 20.905 86.315 21.235 86.330 ;
        RECT 22.490 86.320 22.870 86.330 ;
        RECT 56.570 85.965 56.870 88.355 ;
        RECT 83.005 86.630 83.335 86.645 ;
        RECT 91.525 86.630 95.525 86.780 ;
        RECT 83.005 86.330 95.525 86.630 ;
        RECT 83.005 86.315 83.335 86.330 ;
        RECT 91.525 86.180 95.525 86.330 ;
        RECT 19.985 85.950 20.315 85.965 ;
        RECT 22.745 85.950 23.075 85.965 ;
        RECT 32.405 85.950 32.735 85.965 ;
        RECT 19.985 85.650 32.735 85.950 ;
        RECT 19.985 85.635 20.315 85.650 ;
        RECT 22.745 85.635 23.075 85.650 ;
        RECT 32.405 85.635 32.735 85.650 ;
        RECT 50.805 85.950 51.135 85.965 ;
        RECT 56.325 85.950 56.870 85.965 ;
        RECT 50.805 85.650 56.870 85.950 ;
        RECT 67.825 85.950 68.155 85.965 ;
        RECT 83.005 85.960 83.335 85.965 ;
        RECT 83.005 85.950 83.590 85.960 ;
        RECT 67.825 85.650 83.590 85.950 ;
        RECT 50.805 85.635 51.135 85.650 ;
        RECT 56.325 85.635 56.655 85.650 ;
        RECT 67.825 85.635 68.155 85.650 ;
        RECT 83.005 85.640 83.590 85.650 ;
        RECT 83.005 85.635 83.335 85.640 ;
        RECT 22.285 85.270 22.615 85.285 ;
        RECT 26.885 85.270 27.215 85.285 ;
        RECT 22.285 84.970 27.215 85.270 ;
        RECT 22.285 84.955 22.615 84.970 ;
        RECT 26.885 84.955 27.215 84.970 ;
        RECT 29.850 85.270 30.230 85.280 ;
        RECT 31.025 85.270 31.355 85.285 ;
        RECT 29.850 84.970 31.355 85.270 ;
        RECT 29.850 84.960 30.230 84.970 ;
        RECT 31.025 84.955 31.355 84.970 ;
        RECT 31.945 85.270 32.275 85.285 ;
        RECT 55.405 85.270 55.735 85.285 ;
        RECT 61.845 85.270 62.175 85.285 ;
        RECT 31.945 84.970 35.710 85.270 ;
        RECT 31.945 84.955 32.275 84.970 ;
        RECT 35.410 84.605 35.710 84.970 ;
        RECT 55.405 84.970 62.175 85.270 ;
        RECT 55.405 84.955 55.735 84.970 ;
        RECT 61.845 84.955 62.175 84.970 ;
        RECT 35.410 84.600 35.955 84.605 ;
        RECT 35.370 84.590 35.955 84.600 ;
        RECT 50.345 84.590 50.675 84.605 ;
        RECT 59.545 84.590 59.875 84.605 ;
        RECT 35.370 84.290 36.180 84.590 ;
        RECT 50.345 84.290 59.875 84.590 ;
        RECT 35.370 84.280 35.955 84.290 ;
        RECT 35.625 84.275 35.955 84.280 ;
        RECT 50.345 84.275 50.675 84.290 ;
        RECT 59.545 84.275 59.875 84.290 ;
        RECT 69.205 84.590 69.535 84.605 ;
        RECT 70.330 84.590 70.710 84.600 ;
        RECT 69.205 84.290 70.710 84.590 ;
        RECT 69.205 84.275 69.535 84.290 ;
        RECT 70.330 84.280 70.710 84.290 ;
        RECT 30.930 83.935 32.510 84.265 ;
        RECT 67.570 83.910 67.950 83.920 ;
        RECT 83.465 83.910 83.795 83.925 ;
        RECT 67.570 83.610 83.795 83.910 ;
        RECT 67.570 83.600 67.950 83.610 ;
        RECT 83.465 83.595 83.795 83.610 ;
        RECT 65.525 83.230 65.855 83.245 ;
        RECT 66.650 83.230 67.030 83.240 ;
        RECT 65.525 82.930 67.030 83.230 ;
        RECT 65.525 82.915 65.855 82.930 ;
        RECT 66.650 82.920 67.030 82.930 ;
        RECT 77.025 83.230 77.355 83.245 ;
        RECT 77.690 83.230 78.070 83.240 ;
        RECT 79.785 83.230 80.115 83.245 ;
        RECT 77.025 82.930 80.115 83.230 ;
        RECT 77.025 82.915 77.355 82.930 ;
        RECT 77.690 82.920 78.070 82.930 ;
        RECT 79.785 82.915 80.115 82.930 ;
        RECT 88.065 83.230 88.395 83.245 ;
        RECT 91.525 83.230 95.525 83.380 ;
        RECT 88.065 82.930 95.525 83.230 ;
        RECT 88.065 82.915 88.395 82.930 ;
        RECT 91.525 82.780 95.525 82.930 ;
        RECT 27.630 81.215 29.210 81.545 ;
        RECT 23.410 79.830 23.790 79.840 ;
        RECT 38.385 79.830 38.715 79.845 ;
        RECT 40.225 79.830 40.555 79.845 ;
        RECT 23.410 79.530 40.555 79.830 ;
        RECT 23.410 79.520 23.790 79.530 ;
        RECT 38.385 79.515 38.715 79.530 ;
        RECT 40.225 79.515 40.555 79.530 ;
        RECT 55.405 79.830 55.735 79.845 ;
        RECT 64.605 79.830 64.935 79.845 ;
        RECT 91.525 79.830 95.525 79.980 ;
        RECT 55.405 79.530 64.935 79.830 ;
        RECT 55.405 79.515 55.735 79.530 ;
        RECT 64.605 79.515 64.935 79.530 ;
        RECT 76.120 79.530 95.525 79.830 ;
        RECT 30.930 78.495 32.510 78.825 ;
        RECT 24.585 77.790 24.915 77.805 ;
        RECT 25.250 77.790 25.630 77.800 ;
        RECT 30.565 77.790 30.895 77.805 ;
        RECT 24.585 77.490 30.895 77.790 ;
        RECT 24.585 77.475 24.915 77.490 ;
        RECT 25.250 77.480 25.630 77.490 ;
        RECT 30.565 77.475 30.895 77.490 ;
        RECT 75.185 77.790 75.515 77.805 ;
        RECT 76.120 77.790 76.420 79.530 ;
        RECT 91.525 79.380 95.525 79.530 ;
        RECT 75.185 77.490 76.420 77.790 ;
        RECT 75.185 77.475 75.515 77.490 ;
        RECT 24.585 76.430 24.915 76.445 ;
        RECT 26.170 76.430 26.550 76.440 ;
        RECT 24.585 76.130 26.550 76.430 ;
        RECT 24.585 76.115 24.915 76.130 ;
        RECT 26.170 76.120 26.550 76.130 ;
        RECT 83.465 76.430 83.795 76.445 ;
        RECT 91.525 76.430 95.525 76.580 ;
        RECT 83.465 76.130 95.525 76.430 ;
        RECT 83.465 76.115 83.795 76.130 ;
        RECT 27.630 75.775 29.210 76.105 ;
        RECT 91.525 75.980 95.525 76.130 ;
        RECT 23.665 74.755 23.995 75.085 ;
        RECT 25.965 75.070 26.295 75.085 ;
        RECT 27.805 75.070 28.135 75.085 ;
        RECT 25.965 74.770 28.135 75.070 ;
        RECT 25.965 74.755 26.295 74.770 ;
        RECT 27.805 74.755 28.135 74.770 ;
        RECT 55.865 75.070 56.195 75.085 ;
        RECT 64.810 75.070 65.190 75.080 ;
        RECT 55.865 74.770 65.190 75.070 ;
        RECT 55.865 74.755 56.195 74.770 ;
        RECT 64.810 74.760 65.190 74.770 ;
        RECT 23.680 74.390 23.980 74.755 ;
        RECT 27.805 74.390 28.135 74.405 ;
        RECT 23.680 74.090 28.135 74.390 ;
        RECT 27.805 74.075 28.135 74.090 ;
        RECT 30.930 73.055 32.510 73.385 ;
        RECT 87.605 73.030 87.935 73.045 ;
        RECT 91.525 73.030 95.525 73.180 ;
        RECT 87.605 72.730 95.525 73.030 ;
        RECT 87.605 72.715 87.935 72.730 ;
        RECT 91.525 72.580 95.525 72.730 ;
        RECT 31.025 72.350 31.355 72.365 ;
        RECT 35.370 72.350 35.750 72.360 ;
        RECT 31.025 72.050 35.750 72.350 ;
        RECT 31.025 72.035 31.355 72.050 ;
        RECT 35.370 72.040 35.750 72.050 ;
        RECT 78.610 70.990 78.990 71.000 ;
        RECT 85.765 70.990 86.095 71.005 ;
        RECT 78.610 70.690 86.095 70.990 ;
        RECT 78.610 70.680 78.990 70.690 ;
        RECT 85.765 70.675 86.095 70.690 ;
        RECT 27.630 70.335 29.210 70.665 ;
        RECT 31.485 70.310 31.815 70.325 ;
        RECT 38.845 70.310 39.175 70.325 ;
        RECT 31.485 70.010 39.175 70.310 ;
        RECT 31.485 69.995 31.815 70.010 ;
        RECT 38.845 69.995 39.175 70.010 ;
        RECT 23.665 69.640 23.995 69.645 ;
        RECT 52.185 69.640 52.515 69.645 ;
        RECT 23.410 69.630 23.995 69.640 ;
        RECT 51.930 69.630 52.515 69.640 ;
        RECT 55.865 69.630 56.195 69.645 ;
        RECT 23.410 69.330 24.220 69.630 ;
        RECT 51.730 69.330 56.195 69.630 ;
        RECT 23.410 69.320 23.995 69.330 ;
        RECT 51.930 69.320 52.515 69.330 ;
        RECT 23.665 69.315 23.995 69.320 ;
        RECT 52.185 69.315 52.515 69.320 ;
        RECT 55.865 69.315 56.195 69.330 ;
        RECT 81.625 69.630 81.955 69.645 ;
        RECT 91.525 69.630 95.525 69.780 ;
        RECT 81.625 69.330 95.525 69.630 ;
        RECT 81.625 69.315 81.955 69.330 ;
        RECT 91.525 69.180 95.525 69.330 ;
        RECT 70.125 68.950 70.455 68.965 ;
        RECT 68.530 68.650 70.455 68.950 ;
        RECT 20.905 68.270 21.235 68.285 ;
        RECT 27.345 68.270 27.675 68.285 ;
        RECT 20.905 67.970 27.675 68.270 ;
        RECT 20.905 67.955 21.235 67.970 ;
        RECT 27.345 67.955 27.675 67.970 ;
        RECT 67.825 68.270 68.155 68.285 ;
        RECT 68.530 68.270 68.830 68.650 ;
        RECT 70.125 68.635 70.455 68.650 ;
        RECT 73.805 68.950 74.135 68.965 ;
        RECT 83.925 68.950 84.255 68.965 ;
        RECT 73.805 68.650 84.255 68.950 ;
        RECT 73.805 68.635 74.135 68.650 ;
        RECT 83.925 68.635 84.255 68.650 ;
        RECT 67.825 67.970 68.830 68.270 ;
        RECT 76.565 68.270 76.895 68.285 ;
        RECT 78.865 68.270 79.195 68.285 ;
        RECT 76.565 67.970 79.195 68.270 ;
        RECT 67.825 67.955 68.155 67.970 ;
        RECT 76.565 67.955 76.895 67.970 ;
        RECT 78.865 67.955 79.195 67.970 ;
        RECT 30.930 67.615 32.510 67.945 ;
        RECT 78.405 66.910 78.735 66.925 ;
        RECT 84.385 66.910 84.715 66.925 ;
        RECT 78.405 66.610 84.715 66.910 ;
        RECT 78.405 66.595 78.735 66.610 ;
        RECT 84.385 66.595 84.715 66.610 ;
        RECT 74.725 66.230 75.055 66.245 ;
        RECT 91.525 66.230 95.525 66.380 ;
        RECT 74.725 65.930 95.525 66.230 ;
        RECT 74.725 65.915 75.055 65.930 ;
        RECT 91.525 65.780 95.525 65.930 ;
        RECT 51.930 65.550 52.310 65.560 ;
        RECT 52.645 65.550 52.975 65.565 ;
        RECT 51.930 65.250 52.975 65.550 ;
        RECT 51.930 65.240 52.310 65.250 ;
        RECT 52.645 65.235 52.975 65.250 ;
        RECT 27.630 64.895 29.210 65.225 ;
        RECT 25.250 64.190 25.630 64.200 ;
        RECT 29.185 64.190 29.515 64.205 ;
        RECT 25.250 63.890 29.515 64.190 ;
        RECT 25.250 63.880 25.630 63.890 ;
        RECT 29.185 63.875 29.515 63.890 ;
        RECT 61.385 62.830 61.715 62.845 ;
        RECT 69.410 62.830 69.790 62.840 ;
        RECT 61.385 62.530 69.790 62.830 ;
        RECT 61.385 62.515 61.715 62.530 ;
        RECT 69.410 62.520 69.790 62.530 ;
        RECT 87.605 62.830 87.935 62.845 ;
        RECT 91.525 62.830 95.525 62.980 ;
        RECT 87.605 62.530 95.525 62.830 ;
        RECT 87.605 62.515 87.935 62.530 ;
        RECT 30.930 62.175 32.510 62.505 ;
        RECT 91.525 62.380 95.525 62.530 ;
        RECT 29.850 61.470 30.230 61.480 ;
        RECT 31.485 61.470 31.815 61.485 ;
        RECT 29.850 61.170 31.815 61.470 ;
        RECT 29.850 61.160 30.230 61.170 ;
        RECT 31.485 61.155 31.815 61.170 ;
        RECT 27.630 59.455 29.210 59.785 ;
        RECT 82.545 59.430 82.875 59.445 ;
        RECT 91.525 59.430 95.525 59.580 ;
        RECT 82.545 59.130 95.525 59.430 ;
        RECT 82.545 59.115 82.875 59.130 ;
        RECT 91.525 58.980 95.525 59.130 ;
        RECT 72.425 58.750 72.755 58.765 ;
        RECT 74.930 58.750 75.310 58.760 ;
        RECT 85.305 58.750 85.635 58.765 ;
        RECT 72.425 58.450 85.635 58.750 ;
        RECT 72.425 58.435 72.755 58.450 ;
        RECT 74.930 58.440 75.310 58.450 ;
        RECT 85.305 58.435 85.635 58.450 ;
        RECT 30.930 56.735 32.510 57.065 ;
        RECT 71.045 56.720 71.375 56.725 ;
        RECT 71.045 56.710 71.630 56.720 ;
        RECT 70.820 56.410 71.630 56.710 ;
        RECT 71.045 56.400 71.630 56.410 ;
        RECT 71.045 56.395 71.375 56.400 ;
        RECT 66.905 56.030 67.235 56.045 ;
        RECT 91.525 56.030 95.525 56.180 ;
        RECT 66.905 55.730 95.525 56.030 ;
        RECT 66.905 55.715 67.235 55.730 ;
        RECT 91.525 55.580 95.525 55.730 ;
        RECT 74.010 55.350 74.390 55.360 ;
        RECT 79.325 55.350 79.655 55.365 ;
        RECT 74.010 55.050 79.655 55.350 ;
        RECT 74.010 55.040 74.390 55.050 ;
        RECT 79.325 55.035 79.655 55.050 ;
        RECT 27.630 54.015 29.210 54.345 ;
        RECT 83.005 52.630 83.335 52.645 ;
        RECT 91.525 52.630 95.525 52.780 ;
        RECT 83.005 52.330 95.525 52.630 ;
        RECT 83.005 52.315 83.335 52.330 ;
        RECT 91.525 52.180 95.525 52.330 ;
        RECT 30.930 51.295 32.510 51.625 ;
        RECT 87.605 49.230 87.935 49.245 ;
        RECT 91.525 49.230 95.525 49.380 ;
        RECT 87.605 48.930 95.525 49.230 ;
        RECT 87.605 48.915 87.935 48.930 ;
        RECT 27.630 48.575 29.210 48.905 ;
        RECT 91.525 48.780 95.525 48.930 ;
        RECT 32.865 47.190 33.195 47.205 ;
        RECT 72.885 47.190 73.215 47.205 ;
        RECT 78.865 47.190 79.195 47.205 ;
        RECT 32.865 46.890 33.870 47.190 ;
        RECT 32.865 46.875 33.195 46.890 ;
        RECT 30.930 45.855 32.510 46.185 ;
        RECT 26.885 45.150 27.215 45.165 ;
        RECT 32.405 45.150 32.735 45.165 ;
        RECT 33.570 45.150 33.870 46.890 ;
        RECT 72.885 46.890 79.195 47.190 ;
        RECT 72.885 46.875 73.215 46.890 ;
        RECT 78.865 46.875 79.195 46.890 ;
        RECT 70.585 45.830 70.915 45.845 ;
        RECT 91.525 45.830 95.525 45.980 ;
        RECT 70.585 45.530 95.525 45.830 ;
        RECT 70.585 45.515 70.915 45.530 ;
        RECT 91.525 45.380 95.525 45.530 ;
        RECT 26.885 44.850 33.870 45.150 ;
        RECT 26.885 44.835 27.215 44.850 ;
        RECT 32.405 44.835 32.735 44.850 ;
        RECT 27.630 43.135 29.210 43.465 ;
        RECT 78.865 42.430 79.195 42.445 ;
        RECT 79.530 42.430 79.910 42.440 ;
        RECT 78.865 42.130 79.910 42.430 ;
        RECT 78.865 42.115 79.195 42.130 ;
        RECT 79.530 42.120 79.910 42.130 ;
        RECT 82.545 42.430 82.875 42.445 ;
        RECT 91.525 42.430 95.525 42.580 ;
        RECT 82.545 42.130 95.525 42.430 ;
        RECT 82.545 42.115 82.875 42.130 ;
        RECT 91.525 41.980 95.525 42.130 ;
        RECT 21.365 41.750 21.695 41.765 ;
        RECT 33.325 41.750 33.655 41.765 ;
        RECT 21.365 41.450 33.655 41.750 ;
        RECT 21.365 41.435 21.695 41.450 ;
        RECT 33.325 41.435 33.655 41.450 ;
        RECT 73.345 41.070 73.675 41.085 ;
        RECT 83.005 41.070 83.335 41.085 ;
        RECT 73.345 40.770 83.335 41.070 ;
        RECT 73.345 40.755 73.675 40.770 ;
        RECT 83.005 40.755 83.335 40.770 ;
        RECT 30.930 40.415 32.510 40.745 ;
        RECT 53.770 40.390 54.150 40.400 ;
        RECT 84.845 40.390 85.175 40.405 ;
        RECT 53.770 40.090 85.175 40.390 ;
        RECT 53.770 40.080 54.150 40.090 ;
        RECT 84.845 40.075 85.175 40.090 ;
        RECT 72.425 39.710 72.755 39.725 ;
        RECT 81.625 39.710 81.955 39.725 ;
        RECT 83.465 39.710 83.795 39.725 ;
        RECT 72.425 39.410 83.795 39.710 ;
        RECT 72.425 39.395 72.755 39.410 ;
        RECT 81.625 39.395 81.955 39.410 ;
        RECT 83.465 39.395 83.795 39.410 ;
        RECT 82.545 39.030 82.875 39.045 ;
        RECT 91.525 39.030 95.525 39.180 ;
        RECT 82.545 38.730 95.525 39.030 ;
        RECT 82.545 38.715 82.875 38.730 ;
        RECT 91.525 38.580 95.525 38.730 ;
        RECT 45.285 38.350 45.615 38.365 ;
        RECT 80.245 38.350 80.575 38.365 ;
        RECT 45.285 38.050 80.575 38.350 ;
        RECT 45.285 38.035 45.615 38.050 ;
        RECT 80.245 38.035 80.575 38.050 ;
        RECT 27.630 37.695 29.210 38.025 ;
        RECT 70.585 37.670 70.915 37.685 ;
        RECT 87.605 37.670 87.935 37.685 ;
        RECT 70.585 37.370 87.935 37.670 ;
        RECT 70.585 37.355 70.915 37.370 ;
        RECT 87.605 37.355 87.935 37.370 ;
        RECT 62.765 36.990 63.095 37.005 ;
        RECT 83.925 36.990 84.255 37.005 ;
        RECT 84.845 36.990 85.175 37.005 ;
        RECT 62.765 36.690 85.175 36.990 ;
        RECT 62.765 36.675 63.095 36.690 ;
        RECT 83.925 36.675 84.255 36.690 ;
        RECT 84.845 36.675 85.175 36.690 ;
        RECT 80.245 36.320 80.575 36.325 ;
        RECT 80.245 36.310 80.830 36.320 ;
        RECT 80.020 36.010 80.830 36.310 ;
        RECT 80.245 36.000 80.830 36.010 ;
        RECT 80.245 35.995 80.575 36.000 ;
        RECT 68.285 35.630 68.615 35.645 ;
        RECT 91.525 35.630 95.525 35.780 ;
        RECT 68.285 35.330 95.525 35.630 ;
        RECT 68.285 35.315 68.615 35.330 ;
        RECT 30.930 34.975 32.510 35.305 ;
        RECT 91.525 35.180 95.525 35.330 ;
        RECT 66.445 34.960 66.775 34.965 ;
        RECT 66.445 34.950 67.030 34.960 ;
        RECT 66.220 34.650 67.030 34.950 ;
        RECT 66.445 34.640 67.030 34.650 ;
        RECT 69.410 34.950 69.790 34.960 ;
        RECT 71.505 34.950 71.835 34.965 ;
        RECT 69.410 34.650 71.835 34.950 ;
        RECT 69.410 34.640 69.790 34.650 ;
        RECT 66.445 34.635 66.775 34.640 ;
        RECT 71.505 34.635 71.835 34.650 ;
        RECT 75.645 34.950 75.975 34.965 ;
        RECT 82.545 34.950 82.875 34.965 ;
        RECT 75.645 34.650 82.875 34.950 ;
        RECT 75.645 34.635 75.975 34.650 ;
        RECT 82.545 34.635 82.875 34.650 ;
        RECT 70.330 34.270 70.710 34.280 ;
        RECT 71.045 34.270 71.375 34.285 ;
        RECT 70.330 33.970 71.375 34.270 ;
        RECT 70.330 33.960 70.710 33.970 ;
        RECT 71.045 33.955 71.375 33.970 ;
        RECT 27.630 32.255 29.210 32.585 ;
        RECT 87.605 32.230 87.935 32.245 ;
        RECT 91.525 32.230 95.525 32.380 ;
        RECT 87.605 31.930 95.525 32.230 ;
        RECT 87.605 31.915 87.935 31.930 ;
        RECT 91.525 31.780 95.525 31.930 ;
        RECT 30.930 29.535 32.510 29.865 ;
        RECT 63.890 29.510 64.270 29.520 ;
        RECT 64.605 29.510 64.935 29.525 ;
        RECT 63.890 29.210 64.935 29.510 ;
        RECT 63.890 29.200 64.270 29.210 ;
        RECT 64.605 29.195 64.935 29.210 ;
        RECT 82.545 28.830 82.875 28.845 ;
        RECT 91.525 28.830 95.525 28.980 ;
        RECT 82.545 28.530 95.525 28.830 ;
        RECT 82.545 28.515 82.875 28.530 ;
        RECT 91.525 28.380 95.525 28.530 ;
        RECT 50.345 28.150 50.675 28.165 ;
        RECT 51.930 28.150 52.310 28.160 ;
        RECT 50.345 27.850 52.310 28.150 ;
        RECT 50.345 27.835 50.675 27.850 ;
        RECT 51.930 27.840 52.310 27.850 ;
        RECT 78.610 28.150 78.990 28.160 ;
        RECT 80.245 28.150 80.575 28.165 ;
        RECT 78.610 27.850 80.575 28.150 ;
        RECT 78.610 27.840 78.990 27.850 ;
        RECT 80.245 27.835 80.575 27.850 ;
        RECT 81.370 28.150 81.750 28.160 ;
        RECT 84.845 28.150 85.175 28.165 ;
        RECT 81.370 27.850 85.175 28.150 ;
        RECT 81.370 27.840 81.750 27.850 ;
        RECT 84.845 27.835 85.175 27.850 ;
        RECT 27.630 26.815 29.210 27.145 ;
        RECT 80.705 25.430 81.035 25.445 ;
        RECT 91.525 25.430 95.525 25.580 ;
        RECT 80.705 25.130 95.525 25.430 ;
        RECT 80.705 25.115 81.035 25.130 ;
        RECT 91.525 24.980 95.525 25.130 ;
        RECT 30.930 24.095 32.510 24.425 ;
        RECT 27.630 21.375 29.210 21.705 ;
        RECT 30.930 18.655 32.510 18.985 ;
      LAYER met4 ;
        RECT 63.685 224.985 63.790 225.315 ;
        RECT 66.515 224.965 66.550 225.295 ;
        RECT 69.235 225.005 69.310 225.335 ;
        RECT 72.370 225.045 72.435 225.375 ;
        RECT 74.800 224.975 74.830 225.305 ;
        RECT 77.565 224.995 77.590 225.325 ;
        RECT 77.890 224.995 77.895 225.325 ;
        RECT 80.305 224.915 80.350 225.245 ;
        RECT 83.410 224.945 83.445 225.275 ;
        RECT 85.815 225.025 85.870 225.355 ;
        RECT 88.585 224.955 88.630 225.285 ;
        RECT 91.310 224.985 91.390 225.315 ;
        RECT 93.985 225.015 94.150 225.345 ;
        RECT 118.795 224.760 118.990 225.215 ;
        RECT 119.290 224.760 119.455 225.215 ;
        RECT 121.530 224.805 121.750 225.455 ;
        RECT 122.050 224.805 122.190 225.455 ;
        RECT 124.275 224.945 124.510 225.595 ;
        RECT 124.810 224.945 124.935 225.595 ;
        RECT 127.145 224.965 127.270 225.615 ;
        RECT 127.570 224.965 127.805 225.615 ;
        RECT 129.605 224.960 130.030 225.610 ;
        RECT 133.090 224.945 133.645 225.595 ;
        RECT 134.915 225.075 135.550 225.725 ;
        RECT 137.630 224.895 138.310 225.575 ;
        RECT 142.455 225.400 142.785 225.415 ;
        RECT 142.455 225.100 143.830 225.400 ;
        RECT 142.455 225.085 142.785 225.100 ;
        RECT 118.795 224.565 119.455 224.760 ;
        RECT 112.120 203.770 147.960 203.775 ;
        RECT 8.175 202.180 147.960 203.770 ;
        RECT 112.120 202.175 147.960 202.180 ;
        RECT 6.000 200.475 113.500 200.480 ;
        RECT 6.000 198.890 147.960 200.475 ;
        RECT 112.120 198.875 147.960 198.890 ;
        RECT 10.555 164.515 10.885 164.845 ;
        RECT 10.570 158.725 10.870 164.515 ;
        RECT 10.555 158.395 10.885 158.725 ;
        RECT 26.195 129.155 26.525 129.485 ;
        RECT 22.515 128.475 22.845 128.805 ;
        RECT 22.530 94.125 22.830 128.475 ;
        RECT 26.210 111.125 26.510 129.155 ;
        RECT 26.195 110.795 26.525 111.125 ;
        RECT 26.195 103.995 26.525 104.325 ;
        RECT 22.515 93.795 22.845 94.125 ;
        RECT 22.530 86.645 22.830 93.795 ;
        RECT 22.515 86.315 22.845 86.645 ;
        RECT 22.530 84.590 22.830 86.315 ;
        RECT 22.530 84.290 23.750 84.590 ;
        RECT 23.450 79.845 23.750 84.290 ;
        RECT 23.435 79.515 23.765 79.845 ;
        RECT 23.450 69.645 23.750 79.515 ;
        RECT 25.275 77.475 25.605 77.805 ;
        RECT 23.435 69.315 23.765 69.645 ;
        RECT 25.290 64.205 25.590 77.475 ;
        RECT 26.210 76.445 26.510 103.995 ;
        RECT 26.195 76.115 26.525 76.445 ;
        RECT 25.275 63.875 25.605 64.205 ;
        RECT 27.620 18.580 29.220 174.100 ;
        RECT 29.875 84.955 30.205 85.285 ;
        RECT 29.890 61.485 30.190 84.955 ;
        RECT 29.875 61.155 30.205 61.485 ;
        RECT 30.920 18.580 32.520 174.100 ;
        RECT 47.355 167.235 47.685 167.565 ;
        RECT 75.875 167.235 76.205 167.565 ;
        RECT 45.515 166.555 45.845 166.885 ;
        RECT 45.530 135.605 45.830 166.555 ;
        RECT 47.370 135.605 47.670 167.235 ;
        RECT 74.035 165.195 74.365 165.525 ;
        RECT 60.235 159.755 60.565 160.085 ;
        RECT 53.795 153.635 54.125 153.965 ;
        RECT 45.515 135.275 45.845 135.605 ;
        RECT 47.355 135.275 47.685 135.605 ;
        RECT 51.955 123.035 52.285 123.365 ;
        RECT 35.395 84.275 35.725 84.605 ;
        RECT 35.410 72.365 35.710 84.275 ;
        RECT 35.395 72.035 35.725 72.365 ;
        RECT 51.970 69.645 52.270 123.035 ;
        RECT 52.875 111.475 53.205 111.805 ;
        RECT 52.890 90.725 53.190 111.475 ;
        RECT 52.875 90.395 53.205 90.725 ;
        RECT 51.955 69.315 52.285 69.645 ;
        RECT 51.955 65.235 52.285 65.565 ;
        RECT 51.970 28.165 52.270 65.235 ;
        RECT 53.810 40.405 54.110 153.635 ;
        RECT 60.250 96.845 60.550 159.755 ;
        RECT 66.675 154.995 67.005 155.325 ;
        RECT 65.755 152.955 66.085 153.285 ;
        RECT 61.155 132.555 61.485 132.885 ;
        RECT 60.235 96.515 60.565 96.845 ;
        RECT 61.170 91.405 61.470 132.555 ;
        RECT 64.835 123.035 65.165 123.365 ;
        RECT 63.915 121.675 64.245 122.005 ;
        RECT 61.155 91.075 61.485 91.405 ;
        RECT 53.795 40.075 54.125 40.405 ;
        RECT 63.930 29.525 64.230 121.675 ;
        RECT 64.850 75.085 65.150 123.035 ;
        RECT 65.770 118.605 66.070 152.955 ;
        RECT 65.755 118.275 66.085 118.605 ;
        RECT 66.690 115.205 66.990 154.995 ;
        RECT 69.435 146.155 69.765 146.485 ;
        RECT 67.595 132.555 67.925 132.885 ;
        RECT 66.675 114.875 67.005 115.205 ;
        RECT 67.610 108.390 67.910 132.555 ;
        RECT 69.450 113.845 69.750 146.155 ;
        RECT 74.050 142.405 74.350 165.195 ;
        RECT 75.890 144.445 76.190 167.235 ;
        RECT 77.715 160.435 78.045 160.765 ;
        RECT 76.795 158.395 77.125 158.725 ;
        RECT 75.875 144.115 76.205 144.445 ;
        RECT 74.035 142.075 74.365 142.405 ;
        RECT 76.810 132.885 77.110 158.395 ;
        RECT 77.730 140.365 78.030 160.435 ;
        RECT 77.715 140.035 78.045 140.365 ;
        RECT 80.475 139.355 80.805 139.685 ;
        RECT 79.555 134.595 79.885 134.925 ;
        RECT 76.795 132.555 77.125 132.885 ;
        RECT 71.275 125.755 71.605 126.085 ;
        RECT 69.435 113.515 69.765 113.845 ;
        RECT 66.690 108.090 67.910 108.390 ;
        RECT 66.690 83.245 66.990 108.090 ;
        RECT 67.595 104.675 67.925 105.005 ;
        RECT 67.610 83.925 67.910 104.675 ;
        RECT 70.355 84.275 70.685 84.605 ;
        RECT 67.595 83.595 67.925 83.925 ;
        RECT 66.675 82.915 67.005 83.245 ;
        RECT 64.835 74.755 65.165 75.085 ;
        RECT 66.690 34.965 66.990 82.915 ;
        RECT 69.435 62.515 69.765 62.845 ;
        RECT 69.450 34.965 69.750 62.515 ;
        RECT 66.675 34.635 67.005 34.965 ;
        RECT 69.435 34.635 69.765 34.965 ;
        RECT 70.370 34.285 70.670 84.275 ;
        RECT 71.290 56.725 71.590 125.755 ;
        RECT 72.195 117.595 72.525 117.925 ;
        RECT 72.210 97.525 72.510 117.595 ;
        RECT 74.035 114.875 74.365 115.205 ;
        RECT 72.195 97.195 72.525 97.525 ;
        RECT 71.275 56.395 71.605 56.725 ;
        RECT 74.050 55.365 74.350 114.875 ;
        RECT 74.955 101.275 75.285 101.605 ;
        RECT 74.970 58.765 75.270 101.275 ;
        RECT 77.715 91.755 78.045 92.085 ;
        RECT 77.730 83.245 78.030 91.755 ;
        RECT 77.715 82.915 78.045 83.245 ;
        RECT 78.635 70.675 78.965 71.005 ;
        RECT 74.955 58.435 75.285 58.765 ;
        RECT 74.035 55.035 74.365 55.365 ;
        RECT 70.355 33.955 70.685 34.285 ;
        RECT 63.915 29.195 64.245 29.525 ;
        RECT 78.650 28.165 78.950 70.675 ;
        RECT 79.570 42.445 79.870 134.595 ;
        RECT 80.490 124.045 80.790 139.355 ;
        RECT 80.475 123.715 80.805 124.045 ;
        RECT 80.475 118.275 80.805 118.605 ;
        RECT 79.555 42.115 79.885 42.445 ;
        RECT 80.490 36.325 80.790 118.275 ;
        RECT 83.235 101.955 83.565 102.285 ;
        RECT 81.395 91.075 81.725 91.405 ;
        RECT 80.475 35.995 80.805 36.325 ;
        RECT 81.410 28.165 81.710 91.075 ;
        RECT 83.250 85.965 83.550 101.955 ;
        RECT 157.730 96.590 158.370 97.230 ;
        RECT 83.235 85.635 83.565 85.965 ;
        RECT 51.955 27.835 52.285 28.165 ;
        RECT 78.635 27.835 78.965 28.165 ;
        RECT 81.395 27.835 81.725 28.165 ;
        RECT 157.735 1.065 158.365 96.590 ;
        RECT 16.570 1.000 17.470 1.040 ;
        RECT 35.890 1.000 36.790 1.040 ;
        RECT 55.210 1.000 56.110 1.020 ;
        RECT 152.045 1.000 158.365 1.065 ;
        RECT 152.710 0.435 158.365 1.000 ;
  END
END tt_um_tim2305_adc_dac
END LIBRARY

