* SPICE3 file created from tt_um_tim2305_adc_dac.ext - technology: sky130A

.subckt sky130_fd_pr__res_xhigh_po_0p35_MGD972 a_n35_n486# a_n165_n616# a_n35_54#
X0 a_n35_54# a_n35_n486# a_n165_n616# sky130_fd_pr__res_xhigh_po_0p35 l=0.7
.ends

.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
X0 Q a_1059_315# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_891_413# a_193_47# a_634_159# VNB sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2 a_561_413# a_27_47# a_466_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X3 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4 Q a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 VGND a_634_159# a_592_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X7 VPWR a_891_413# a_1059_315# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8 a_466_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X9 VPWR a_634_159# a_561_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X10 a_634_159# a_466_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X11 a_634_159# a_466_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X12 a_975_413# a_193_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 VGND a_1059_315# a_1017_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X14 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15 a_891_413# a_27_47# a_634_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X16 a_592_47# a_193_47# a_466_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X17 a_1017_47# a_27_47# a_891_413# VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X18 VPWR a_1059_315# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X19 a_466_413# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X20 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X21 VGND a_891_413# a_1059_315# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X22 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X23 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
X0 a_222_93# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X1 VPWR A1 a_544_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.105 ps=1.21 w=1 l=0.15
X2 VGND a_79_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_222_93# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.18575 ps=1.415 w=0.42 l=0.15
X4 VGND A2 a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X5 a_448_47# a_222_93# a_79_199# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X6 a_79_199# a_222_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.3 ps=2.6 w=1 l=0.15
X7 a_544_297# A2 a_79_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X8 a_448_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VPWR a_79_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18575 pd=1.415 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
X0 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X1 a_109_53# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_215_297# a_109_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.101875 ps=0.99 w=0.65 l=0.15
X4 a_392_297# C a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.04515 pd=0.635 as=0.06825 ps=0.745 w=0.42 l=0.15
X5 a_465_297# B a_392_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06405 pd=0.725 as=0.04515 ps=0.635 w=0.42 l=0.15
X6 a_215_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 VPWR A a_465_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06405 ps=0.725 w=0.42 l=0.15
X8 a_297_297# a_109_53# a_215_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 a_109_53# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X10 VGND C a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06405 ps=0.725 w=0.42 l=0.15
X11 VGND A a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=0.59
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=0.59
.ends

.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
X0 VPWR a_505_21# a_535_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_505_21# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_218_374# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X3 VGND a_505_21# a_439_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_76_199# A0 a_218_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X5 a_505_21# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X6 a_439_47# A0 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X7 a_535_374# A1 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X8 a_76_199# A1 a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_218_47# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=1.05
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=1.05
.ends

.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=2.89
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=2.89
.ends

.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X1 a_209_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X2 a_303_47# A2 a_209_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X3 a_209_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X5 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X6 a_80_21# A1 a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X7 VPWR A2 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X8 a_80_21# B1 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X9 a_209_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
X0 VPWR A a_49_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 VGND a_285_47# a_391_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.5
X2 X a_391_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X3 VGND A a_49_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 VPWR a_285_47# a_391_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.5
X5 a_285_47# a_49_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X6 a_285_47# a_49_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X7 X a_391_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.101875 ps=0.99 w=0.65 l=0.15
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.14825 ps=1.34 w=1 l=0.15
X7 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
X0 VPWR B a_207_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X1 X a_207_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X2 a_297_47# a_27_413# a_207_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 X a_207_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X4 a_207_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 VGND B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X7 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
X0 X a_29_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.14825 ps=1.34 w=1 l=0.15
X1 a_111_297# C a_29_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 X a_29_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.101875 ps=0.99 w=0.65 l=0.15
X3 a_183_297# B a_111_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 VPWR A a_183_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_29_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VGND C a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 VGND A a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
X0 VPWR a_212_413# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_297_47# a_27_413# a_212_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 X a_212_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.22895 ps=1.745 w=1 l=0.15
X3 X a_212_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.101875 ps=0.99 w=0.65 l=0.15
X4 a_212_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.07665 ps=0.785 w=0.42 l=0.15
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 VPWR B a_212_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.22895 pd=1.745 as=0.0609 ps=0.71 w=0.42 l=0.15
X7 VGND B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VGND a_212_413# X VNB sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=1.97
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=1.97
.ends

.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X6 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X7 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X14 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X16 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X17 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X18 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X19 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X20 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X21 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X22 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X23 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X24 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X25 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X26 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X27 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X28 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X29 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X30 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X31 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X32 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X33 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X34 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X35 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X36 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X37 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X38 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X39 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
.ends

.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
X0 a_103_199# B1 a_253_47# VNB sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X1 VPWR a_103_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.36 ps=2.72 w=1 l=0.15
X2 a_337_297# A2 a_253_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3 a_103_199# A3 a_337_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2125 pd=1.425 as=0.165 ps=1.33 w=1 l=0.15
X4 a_253_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.195 ps=1.39 w=1 l=0.15
X5 VPWR B1 a_103_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.345 pd=2.69 as=0.2125 ps=1.425 w=1 l=0.15
X6 VGND a_103_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.234 ps=2.02 w=0.65 l=0.15
X7 a_253_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12675 ps=1.04 w=0.65 l=0.15
X8 a_253_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X9 VGND A2 a_253_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
X0 VPWR A a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_109_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
X0 VGND A4 a_321_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_321_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.1235 ps=1.03 w=0.65 l=0.15
X2 a_103_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=1.52 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR a_103_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.425 ps=2.85 w=1 l=0.15
X4 VGND a_103_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.247 ps=2.06 w=0.65 l=0.15
X5 VGND A2 a_321_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X6 a_321_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.12675 ps=1.04 w=0.65 l=0.15
X7 a_511_297# A3 a_393_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.22 ps=1.44 w=1 l=0.15
X8 a_619_297# A2 a_511_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X9 a_321_47# B1 a_103_21# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10 a_393_297# A4 a_103_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.26 ps=1.52 w=1 l=0.15
X11 VPWR A1 a_619_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.195 ps=1.39 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
X0 VGND A a_68_297# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_68_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 X a_68_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X3 VPWR A a_150_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 X a_68_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X5 a_150_297# B a_68_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=4.73
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=4.73
.ends

.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
X0 VPWR A1 a_382_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X1 a_297_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X2 a_297_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VGND A2 a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3275 pd=1.655 as=0.28 ps=2.56 w=1 l=0.15
X5 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.3275 ps=1.655 w=1 l=0.15
X6 a_382_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.195 ps=1.39 w=1 l=0.15
X7 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt bit4_encoder VPWR bus0[0] bus0[1] bus0[2] bus0[3] bus1[0] bus1[1] bus1[2]
+ bus1[3] bus2[0] bus2[1] bus2[2] bus2[3] clk compr[0] compr[12] compr[14] compr[1]
+ compr[2] compr[3] compr[4] compr[5] compr[8] compr[11] compr[7] compr[13] compr[9]
+ compr[10] VGND compr[6]
X_83_ clknet_1_0__leaf_clk _05_ VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__dfxtp_1
X_49_ net2 _21_ net3 VGND VGND VPWR VPWR _22_ sky130_fd_sc_hd__o21ba_1
X_66_ net15 _33_ net2 _27_ VGND VGND VPWR VPWR _36_ sky130_fd_sc_hd__or4b_1
XPHY_EDGE_ROW_12_Left_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput20 net20 VGND VGND VPWR VPWR bus1[0] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_0_Left_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_82_ clknet_1_0__leaf_clk _04_ VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__dfxtp_1
X_65_ net28 _35_ _15_ VGND VGND VPWR VPWR _04_ sky130_fd_sc_hd__mux2_1
X_48_ net14 _20_ net15 VGND VGND VPWR VPWR _21_ sky130_fd_sc_hd__o21ba_1
Xoutput21 net21 VGND VGND VPWR VPWR bus1[1] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_81_ clknet_1_1__leaf_clk _03_ VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__dfxtp_1
XFILLER_3_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_47_ net12 _19_ net13 VGND VGND VPWR VPWR _20_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_64_ _27_ _29_ _34_ _33_ VGND VGND VPWR VPWR _35_ sky130_fd_sc_hd__a31o_1
Xhold10 net20 VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__dlygate4sd3_1
Xoutput22 net22 VGND VGND VPWR VPWR bus1[2] sky130_fd_sc_hd__buf_2
X_80_ clknet_1_1__leaf_clk _02_ VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__dfxtp_1
X_63_ net9 net10 net11 net12 VGND VGND VPWR VPWR _34_ sky130_fd_sc_hd__or4_1
XFILLER_9_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_46_ net10 _18_ net11 VGND VGND VPWR VPWR _19_ sky130_fd_sc_hd__o21ba_1
Xhold11 net24 VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__dlygate4sd3_1
Xoutput23 net23 VGND VGND VPWR VPWR bus1[3] sky130_fd_sc_hd__buf_2
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_62_ net3 net4 net5 net6 VGND VGND VPWR VPWR _33_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_4_Left_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold12 bus_count\[1\] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__dlygate4sd3_1
X_45_ net8 _17_ net9 VGND VGND VPWR VPWR _18_ sky130_fd_sc_hd__o21ba_1
XPHY_EDGE_ROW_7_Left_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput24 net24 VGND VGND VPWR VPWR bus2[0] sky130_fd_sc_hd__buf_2
XFILLER_6_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_61_ net33 _32_ _15_ VGND VGND VPWR VPWR _03_ sky130_fd_sc_hd__mux2_1
XFILLER_9_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_44_ net7 net1 VGND VGND VPWR VPWR _17_ sky130_fd_sc_hd__and2b_1
Xhold13 _10_ VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__dlygate4sd3_1
Xoutput25 net25 VGND VGND VPWR VPWR bus2[1] sky130_fd_sc_hd__buf_2
X_60_ net5 net6 _31_ VGND VGND VPWR VPWR _32_ sky130_fd_sc_hd__or3_1
X_43_ _15_ VGND VGND VPWR VPWR _16_ sky130_fd_sc_hd__inv_2
Xhold14 bus_count\[0\] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__dlygate4sd3_1
Xoutput26 net26 VGND VGND VPWR VPWR bus2[2] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_42_ bus_count\[0\] bus_count\[1\] VGND VGND VPWR VPWR _15_ sky130_fd_sc_hd__and2b_2
Xoutput16 net16 VGND VGND VPWR VPWR bus0[0] sky130_fd_sc_hd__buf_2
XFILLER_7_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
Xoutput27 net27 VGND VGND VPWR VPWR bus2[3] sky130_fd_sc_hd__buf_2
XFILLER_4_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_41_ _01_ VGND VGND VPWR VPWR _14_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_11_Left_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput17 net17 VGND VGND VPWR VPWR bus0[1] sky130_fd_sc_hd__buf_2
X_40_ bus_count\[1\] bus_count\[0\] VGND VGND VPWR VPWR _01_ sky130_fd_sc_hd__and2b_2
Xoutput18 net18 VGND VGND VPWR VPWR bus0[2] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput19 net19 VGND VGND VPWR VPWR bus0[3] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_3_Left_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput1 compr[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput2 compr[10] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__buf_1
X_79_ clknet_1_1__leaf_clk _01_ VGND VGND VPWR VPWR bus_count\[1\] sky130_fd_sc_hd__dfxtp_1
Xinput3 compr[11] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
XFILLER_1_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_78_ clknet_1_0__leaf_clk _00_ VGND VGND VPWR VPWR bus_count\[0\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput4 compr[12] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_1
X_77_ net30 _36_ _00_ VGND VGND VPWR VPWR _13_ sky130_fd_sc_hd__mux2_1
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput5 compr[13] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_1
X_76_ net35 _35_ _00_ VGND VGND VPWR VPWR _12_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_10_Left_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_59_ net15 net2 _28_ _30_ VGND VGND VPWR VPWR _31_ sky130_fd_sc_hd__o31a_1
XFILLER_1_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput6 compr[14] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__buf_1
X_58_ net3 net4 VGND VGND VPWR VPWR _30_ sky130_fd_sc_hd__nor2_1
X_75_ net32 _32_ _00_ VGND VGND VPWR VPWR _11_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_91_ clknet_1_0__leaf_clk _13_ VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__dfxtp_1
X_74_ bus_count\[0\] net39 net6 _23_ _38_ VGND VGND VPWR VPWR _10_ sky130_fd_sc_hd__o41a_1
Xinput7 compr[1] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_1
XFILLER_5_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_57_ net15 net2 VGND VGND VPWR VPWR _29_ sky130_fd_sc_hd__nor2_1
Xinput10 compr[4] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__buf_1
XFILLER_4_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_90_ clknet_1_0__leaf_clk _12_ VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__dfxtp_1
X_73_ net16 _00_ VGND VGND VPWR VPWR _38_ sky130_fd_sc_hd__or2_1
Xinput8 compr[2] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_1
X_56_ net11 net12 _26_ _27_ VGND VGND VPWR VPWR _28_ sky130_fd_sc_hd__o31a_1
X_39_ net41 net39 VGND VGND VPWR VPWR _00_ sky130_fd_sc_hd__nor2_1
Xclkbuf_1_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
Xinput11 compr[5] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_2_Left_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput9 compr[3] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_1
X_72_ net31 _36_ _01_ VGND VGND VPWR VPWR _09_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput12 compr[6] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__buf_1
X_55_ net13 net14 VGND VGND VPWR VPWR _27_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1 net26 VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__dlygate4sd3_1
X_54_ net7 net8 _25_ VGND VGND VPWR VPWR _26_ sky130_fd_sc_hd__o21a_1
X_71_ net36 _35_ _01_ VGND VGND VPWR VPWR _08_ sky130_fd_sc_hd__mux2_1
Xinput13 compr[7] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_1
Xhold2 net21 VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__dlygate4sd3_1
X_70_ net29 _32_ _01_ VGND VGND VPWR VPWR _07_ sky130_fd_sc_hd__mux2_1
Xinput14 compr[8] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_1
X_53_ net9 net10 VGND VGND VPWR VPWR _25_ sky130_fd_sc_hd__nor2_1
Xhold3 net19 VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__dlygate4sd3_1
X_52_ net6 _16_ _23_ _24_ VGND VGND VPWR VPWR _02_ sky130_fd_sc_hd__o31a_1
Xinput15 compr[9] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_6_Left_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_9_Left_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold4 net23 VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__dlygate4sd3_1
X_51_ net38 _15_ VGND VGND VPWR VPWR _24_ sky130_fd_sc_hd__or2_1
XFILLER_0_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold5 net17 VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__dlygate4sd3_1
X_50_ net4 _22_ net5 VGND VGND VPWR VPWR _23_ sky130_fd_sc_hd__o21ba_1
Xhold6 net25 VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold7 net27 VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold8 net18 VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_1_Left_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold9 net22 VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_89_ clknet_1_1__leaf_clk _11_ VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__dfxtp_1
XFILLER_2_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_88_ clknet_1_1__leaf_clk net40 VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__dfxtp_1
X_87_ clknet_1_0__leaf_clk _09_ VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_5_Left_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_8_Left_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_86_ clknet_1_0__leaf_clk _08_ VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__dfxtp_1
X_69_ net6 _14_ _23_ _37_ VGND VGND VPWR VPWR _06_ sky130_fd_sc_hd__o31a_1
XFILLER_12_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_85_ clknet_1_1__leaf_clk _07_ VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__dfxtp_1
X_68_ net37 _01_ VGND VGND VPWR VPWR _37_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_84_ clknet_1_1__leaf_clk _06_ VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__dfxtp_1
X_67_ net34 _36_ _15_ VGND VGND VPWR VPWR _05_ sky130_fd_sc_hd__mux2_1
XFILLER_6_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
C0 VPWR _36_ 2.108505f
C1 VPWR clknet_1_1__leaf_clk 2.109072f
C2 VPWR clknet_1_0__leaf_clk 2.060224f
C3 VPWR _00_ 2.496267f
C4 _01_ VGND 3.226816f
C5 _00_ VGND 2.658476f
C6 VPWR VGND 92.371376f
C7 _15_ VGND 2.114687f
C8 clknet_1_0__leaf_clk VGND 3.388226f
.ends

.subckt sky130_fd_pr__nfet_01v8_64Z3AY a_15_n131# a_n175_n243# a_n33_91# a_n73_n131#
X0 a_15_n131# a_n33_91# a_n73_n131# a_n175_n243# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_3H2EVM a_n100_n897# a_100_n800# w_n296_n1019# a_n158_n800#
+ VSUBS
X0 a_100_n800# a_n100_n897# a_n158_n800# w_n296_n1019# sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=1
C0 w_n296_n1019# VSUBS 4.82082f
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_AHMAL2 a_n260_n574# a_100_n400# a_n158_n400# a_n100_n488#
X0 a_100_n400# a_n100_n488# a_n158_n400# a_n260_n574# sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_AHRV9L a_n258_n400# a_n200_n488# a_n360_n574#
+ a_200_n400#
X0 a_200_n400# a_n200_n488# a_n258_n400# a_n360_n574# sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_GWPMZG a_n200_n897# a_200_n800# w_n396_n1019#
+ a_n258_n800# VSUBS
X0 a_200_n800# a_n200_n897# a_n258_n800# w_n396_n1019# sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=2
C0 w_n396_n1019# VSUBS 6.14037f
.ends

.subckt sky130_fd_pr__pfet_01v8_MGSNAN a_n73_n336# a_n33_295# w_n211_n484# VSUBS
X0 a_15_n336# a_n33_295# a_n73_n336# w_n211_n484# sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
.ends

.subckt compr out vdd in+ in- vss
XXM1 out vss m1_2518_1378# vss sky130_fd_pr__nfet_01v8_64Z3AY
XXM3 m1_1460_732# vdd vdd m1_1264_902# vss sky130_fd_pr__pfet_01v8_3H2EVM
XXM4 vss vss m1_1264_902# m1_1460_732# sky130_fd_pr__nfet_01v8_lvt_AHMAL2
XXM5 m1_1824_498# m1_1824_498# vss vss sky130_fd_pr__nfet_01v8_lvt_AHRV9L
XXM6 m1_2518_1378# m1_2518_1378# vss vss sky130_fd_pr__nfet_01v8_lvt_AHRV9L
XXM7 in- m1_2324_1380# vdd m1_1824_498# vss sky130_fd_pr__pfet_01v8_lvt_GWPMZG
XXM8 m1_1264_902# vdd vdd m1_2324_1380# vss sky130_fd_pr__pfet_01v8_3H2EVM
XXM9 in+ m1_2324_1380# vdd m1_2518_1378# vss sky130_fd_pr__pfet_01v8_lvt_GWPMZG
XXM21 out m1_2518_1378# vdd vss sky130_fd_pr__pfet_01v8_MGSNAN
R0 m1_1264_902# m1_1264_902# sky130_fd_pr__res_generic_m1 w=0.42 l=7.37
C0 m1_2518_1378# vss 3.214547f
C1 vdd vss 21.48598f
C2 m1_1824_498# vss 2.487121f
.ends

.subckt flash_adc out VSUBS
XXR1 compr_13/in- VSUBS compr_14/in- sky130_fd_pr__res_xhigh_po_0p35_MGD972
XXR2 compr_5/in- VSUBS compr_6/in- sky130_fd_pr__res_xhigh_po_0p35_MGD972
XXR10 compr_6/in- VSUBS compr_7/in- sky130_fd_pr__res_xhigh_po_0p35_MGD972
XXR3 compr_11/in- VSUBS compr_12/in- sky130_fd_pr__res_xhigh_po_0p35_MGD972
XXR11 compr_10/in- VSUBS compr_11/in- sky130_fd_pr__res_xhigh_po_0p35_MGD972
Xbit4_encoder_0 bit4_encoder_0/VPWR bit4_encoder_0/bus0[0] bit4_encoder_0/bus0[1]
+ bit4_encoder_0/bus0[2] bit4_encoder_0/bus0[3] bit4_encoder_0/bus1[0] bit4_encoder_0/bus1[1]
+ bit4_encoder_0/bus1[2] bit4_encoder_0/bus1[3] bit4_encoder_0/bus2[0] bit4_encoder_0/bus2[1]
+ bit4_encoder_0/bus2[2] bit4_encoder_0/bus2[3] bit4_encoder_0/clk compr_0/out compr_12/out
+ compr_14/out compr_1/out compr_2/out compr_3/out compr_4/out compr_5/out compr_8/out
+ compr_11/out compr_7/out compr_13/out compr_9/out compr_10/out VSUBS compr_6/out
+ bit4_encoder
XXR4 compr_14/in- VSUBS compr_14/vdd sky130_fd_pr__res_xhigh_po_0p35_MGD972
XXR5 compr_7/in- VSUBS compr_8/in- sky130_fd_pr__res_xhigh_po_0p35_MGD972
XXR12 compr_8/in- VSUBS compr_9/in- sky130_fd_pr__res_xhigh_po_0p35_MGD972
XXR6 compr_0/in- VSUBS compr_1/in- sky130_fd_pr__res_xhigh_po_0p35_MGD972
XXR13 VSUBS VSUBS compr_0/in- sky130_fd_pr__res_xhigh_po_0p35_MGD972
XXR14 compr_1/in- VSUBS compr_2/in- sky130_fd_pr__res_xhigh_po_0p35_MGD972
XXR7 compr_9/in- VSUBS compr_10/in- sky130_fd_pr__res_xhigh_po_0p35_MGD972
XXR15 compr_3/in- VSUBS compr_4/in- sky130_fd_pr__res_xhigh_po_0p35_MGD972
XXR8 compr_4/in- VSUBS compr_5/in- sky130_fd_pr__res_xhigh_po_0p35_MGD972
XXR16 compr_2/in- VSUBS compr_3/in- sky130_fd_pr__res_xhigh_po_0p35_MGD972
XXR9 compr_12/in- VSUBS compr_13/in- sky130_fd_pr__res_xhigh_po_0p35_MGD972
Xcompr_0 compr_0/out compr_4/vdd out compr_0/in- VSUBS compr
Xcompr_1 compr_1/out compr_4/vdd out compr_1/in- VSUBS compr
Xcompr_2 compr_2/out compr_4/vdd out compr_2/in- VSUBS compr
Xcompr_3 compr_3/out compr_4/vdd out compr_3/in- VSUBS compr
Xcompr_4 compr_4/out compr_4/vdd out compr_4/in- VSUBS compr
Xcompr_5 compr_5/out compr_9/vdd out compr_5/in- VSUBS compr
Xcompr_6 compr_6/out compr_9/vdd out compr_6/in- VSUBS compr
Xcompr_7 compr_7/out compr_9/vdd out compr_7/in- VSUBS compr
Xcompr_10 compr_10/out compr_14/vdd out compr_10/in- VSUBS compr
Xcompr_8 compr_8/out compr_9/vdd out compr_8/in- VSUBS compr
Xcompr_11 compr_11/out compr_14/vdd out compr_11/in- VSUBS compr
Xcompr_9 compr_9/out compr_9/vdd out compr_9/in- VSUBS compr
Xcompr_13 compr_13/out compr_14/vdd out compr_13/in- VSUBS compr
Xcompr_12 compr_12/out compr_14/vdd out compr_12/in- VSUBS compr
Xcompr_14 compr_14/out compr_14/vdd out compr_14/in- VSUBS compr
C0 compr_5/out compr_4/in- 6.637179f
C1 compr_1/in- out 2.212074f
C2 compr_14/vdd compr_14/in- 3.817381f
C3 compr_7/out compr_8/out 3.990631f
C4 compr_4/vdd compr_2/in- 4.728872f
C5 compr_11/out compr_12/out 3.951141f
C6 compr_13/in- compr_14/in- 6.444436f
C7 compr_6/out compr_7/out 5.567697f
C8 compr_7/in- compr_8/in- 4.873167f
C9 compr_8/out compr_9/out 3.030994f
C10 compr_9/vdd compr_7/in- 2.60179f
C11 compr_11/out compr_10/out 7.344403f
C12 compr_4/vdd compr_3/in- 3.604922f
C13 compr_11/in- compr_14/vdd 2.383896f
C14 compr_6/in- compr_5/in- 2.207374f
C15 compr_2/in- compr_3/in- 3.707407f
C16 compr_12/in- compr_11/in- 3.861109f
C17 compr_4/out compr_3/out 2.196932f
C18 compr_1/out compr_0/out 6.062403f
C19 compr_13/in- compr_14/vdd 3.767509f
C20 compr_12/in- compr_14/vdd 3.328351f
C21 compr_14/out compr_13/out 2.960663f
C22 out compr_9/vdd 2.042017f
C23 compr_1/out compr_2/out 5.785456f
C24 compr_4/in- compr_3/in- 6.431217f
C25 compr_12/in- compr_13/in- 5.007227f
C26 compr_9/vdd compr_6/in- 3.191535f
C27 compr_9/in- compr_10/out 6.166734f
C28 compr_7/in- compr_6/in- 3.808161f
C29 compr_3/out compr_2/out 3.621265f
C30 compr_13/out compr_12/out 2.705792f
C31 compr_6/out compr_5/out 6.042858f
C32 compr_9/in- compr_8/in- 6.294752f
C33 compr_14/m1_2518_1378# VSUBS 2.251797f
C34 compr_14/vdd VSUBS 0.104742p
C35 compr_14/in- VSUBS 2.919514f
C36 compr_12/m1_2518_1378# VSUBS 2.251923f
C37 compr_13/m1_2518_1378# VSUBS 2.251823f
C38 compr_9/m1_2518_1378# VSUBS 2.252194f
C39 compr_9/vdd VSUBS 0.106776p
C40 compr_11/out VSUBS 2.551758f
C41 compr_11/m1_2518_1378# VSUBS 2.251958f
C42 compr_8/m1_2518_1378# VSUBS 2.252175f
C43 compr_10/out VSUBS 5.61895f
C44 compr_10/m1_2518_1378# VSUBS 2.248816f
C45 compr_7/out VSUBS 3.429728f
C46 compr_7/m1_2518_1378# VSUBS 2.251962f
C47 compr_6/m1_2518_1378# VSUBS 2.25198f
C48 compr_5/m1_2518_1378# VSUBS 2.248871f
C49 compr_4/m1_2518_1378# VSUBS 2.252f
C50 compr_4/vdd VSUBS 0.106607p
C51 out VSUBS 11.112763f
C52 compr_4/in- VSUBS 3.311688f
C53 compr_3/m1_2518_1378# VSUBS 2.252004f
C54 compr_3/in- VSUBS 2.123285f
C55 compr_2/out VSUBS 2.544032f
C56 compr_2/m1_2518_1378# VSUBS 2.251982f
C57 compr_1/out VSUBS 2.914421f
C58 compr_1/m1_2518_1378# VSUBS 2.252f
C59 compr_0/out VSUBS 7.89841f
C60 compr_0/m1_2518_1378# VSUBS 2.253713f
C61 compr_0/in- VSUBS 2.051001f
C62 compr_12/in- VSUBS 2.12567f
C63 compr_13/in- VSUBS 2.125113f
C64 compr_2/in- VSUBS 2.024528f
C65 compr_5/in- VSUBS 2.088458f
C66 compr_8/in- VSUBS 3.977413f
C67 compr_9/in- VSUBS 6.995159f
C68 compr_6/out VSUBS 4.979608f
C69 compr_5/out VSUBS 5.536202f
C70 bit4_encoder_0/VPWR VSUBS 94.88836f
C71 compr_12/out VSUBS 2.188971f
C72 compr_10/in- VSUBS 2.024571f
C73 compr_11/in- VSUBS 2.107752f
C74 compr_7/in- VSUBS 2.354412f
.ends

.subckt tt_um_tim2305_adc_dac clk ena rst_n ua[0] ua[1] ua[2] ua[3] ua[4] ua[5] ua[6]
+ ua[7] ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0]
+ uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7] uio_oe[0]
+ uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0]
+ uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7] uo_out[0]
+ uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7] VDPWR VGND
Xflash_adc_0 ua[0] VSUBS flash_adc
C0 VGND VDPWR 12.918099f
C1 VGND VSUBS 12.5347f
C2 VDPWR VSUBS 12.5347f
C3 flash_adc_0/compr_14/m1_2518_1378# VSUBS 2.24793f
C4 flash_adc_0/compr_14/vdd VSUBS 0.103907p
C5 flash_adc_0/compr_14/in- VSUBS 2.830427f
C6 flash_adc_0/compr_12/m1_2518_1378# VSUBS 2.24793f
C7 flash_adc_0/compr_13/m1_2518_1378# VSUBS 2.24793f
C8 flash_adc_0/compr_9/m1_2518_1378# VSUBS 2.24793f
C9 flash_adc_0/compr_9/vdd VSUBS 99.35699f
C10 flash_adc_0/compr_11/m1_2518_1378# VSUBS 2.24793f
C11 flash_adc_0/compr_8/m1_2518_1378# VSUBS 2.24793f
C12 flash_adc_0/compr_10/m1_2518_1378# VSUBS 2.24793f
C13 flash_adc_0/compr_7/m1_2518_1378# VSUBS 2.24793f
C14 flash_adc_0/compr_6/m1_2518_1378# VSUBS 2.24793f
C15 flash_adc_0/compr_5/m1_2518_1378# VSUBS 2.24793f
C16 flash_adc_0/compr_4/m1_2518_1378# VSUBS 2.24793f
C17 flash_adc_0/compr_4/vdd VSUBS 99.06754f
C18 ua[0] VSUBS 19.831497f
C19 flash_adc_0/compr_3/m1_2518_1378# VSUBS 2.24793f
C20 flash_adc_0/compr_2/m1_2518_1378# VSUBS 2.24793f
C21 flash_adc_0/compr_1/m1_2518_1378# VSUBS 2.24793f
C22 flash_adc_0/compr_0/out VSUBS 2.16099f
C23 flash_adc_0/compr_0/m1_2518_1378# VSUBS 2.24793f
C24 flash_adc_0/compr_13/in- VSUBS 2.017837f
C25 flash_adc_0/compr_8/in- VSUBS 2.135297f
C26 flash_adc_0/bit4_encoder_0/VPWR VSUBS 94.88836f
C27 flash_adc_0/compr_7/in- VSUBS 2.004427f
.ends

